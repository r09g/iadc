magic
tech sky130A
magscale 1 2
timestamp 1654728500
<< nwell >>
rect -64 1502 3554 3096
<< pwell >>
rect -34 -64 3524 1452
<< mvnmos >>
rect 194 194 294 1194
rect 352 194 452 1194
rect 510 194 610 1194
rect 668 194 768 1194
rect 826 194 926 1194
rect 984 194 1084 1194
rect 1142 194 1242 1194
rect 1300 194 1400 1194
rect 1458 194 1558 1194
rect 1616 194 1716 1194
rect 1774 194 1874 1194
rect 1932 194 2032 1194
rect 2090 194 2190 1194
rect 2248 194 2348 1194
rect 2406 194 2506 1194
rect 2564 194 2664 1194
rect 2722 194 2822 1194
rect 2880 194 2980 1194
rect 3038 194 3138 1194
rect 3196 194 3296 1194
<< mvpmos >>
rect 194 1799 294 2799
rect 352 1799 452 2799
rect 510 1799 610 2799
rect 668 1799 768 2799
rect 826 1799 926 2799
rect 984 1799 1084 2799
rect 1142 1799 1242 2799
rect 1300 1799 1400 2799
rect 1458 1799 1558 2799
rect 1616 1799 1716 2799
rect 1774 1799 1874 2799
rect 1932 1799 2032 2799
rect 2090 1799 2190 2799
rect 2248 1799 2348 2799
rect 2406 1799 2506 2799
rect 2564 1799 2664 2799
rect 2722 1799 2822 2799
rect 2880 1799 2980 2799
rect 3038 1799 3138 2799
rect 3196 1799 3296 2799
<< mvndiff >>
rect 136 1182 194 1194
rect 136 206 148 1182
rect 182 206 194 1182
rect 136 194 194 206
rect 294 1182 352 1194
rect 294 206 306 1182
rect 340 206 352 1182
rect 294 194 352 206
rect 452 1182 510 1194
rect 452 206 464 1182
rect 498 206 510 1182
rect 452 194 510 206
rect 610 1182 668 1194
rect 610 206 622 1182
rect 656 206 668 1182
rect 610 194 668 206
rect 768 1182 826 1194
rect 768 206 780 1182
rect 814 206 826 1182
rect 768 194 826 206
rect 926 1182 984 1194
rect 926 206 938 1182
rect 972 206 984 1182
rect 926 194 984 206
rect 1084 1182 1142 1194
rect 1084 206 1096 1182
rect 1130 206 1142 1182
rect 1084 194 1142 206
rect 1242 1182 1300 1194
rect 1242 206 1254 1182
rect 1288 206 1300 1182
rect 1242 194 1300 206
rect 1400 1182 1458 1194
rect 1400 206 1412 1182
rect 1446 206 1458 1182
rect 1400 194 1458 206
rect 1558 1182 1616 1194
rect 1558 206 1570 1182
rect 1604 206 1616 1182
rect 1558 194 1616 206
rect 1716 1182 1774 1194
rect 1716 206 1728 1182
rect 1762 206 1774 1182
rect 1716 194 1774 206
rect 1874 1182 1932 1194
rect 1874 206 1886 1182
rect 1920 206 1932 1182
rect 1874 194 1932 206
rect 2032 1182 2090 1194
rect 2032 206 2044 1182
rect 2078 206 2090 1182
rect 2032 194 2090 206
rect 2190 1182 2248 1194
rect 2190 206 2202 1182
rect 2236 206 2248 1182
rect 2190 194 2248 206
rect 2348 1182 2406 1194
rect 2348 206 2360 1182
rect 2394 206 2406 1182
rect 2348 194 2406 206
rect 2506 1182 2564 1194
rect 2506 206 2518 1182
rect 2552 206 2564 1182
rect 2506 194 2564 206
rect 2664 1182 2722 1194
rect 2664 206 2676 1182
rect 2710 206 2722 1182
rect 2664 194 2722 206
rect 2822 1182 2880 1194
rect 2822 206 2834 1182
rect 2868 206 2880 1182
rect 2822 194 2880 206
rect 2980 1182 3038 1194
rect 2980 206 2992 1182
rect 3026 206 3038 1182
rect 2980 194 3038 206
rect 3138 1182 3196 1194
rect 3138 206 3150 1182
rect 3184 206 3196 1182
rect 3138 194 3196 206
rect 3296 1182 3354 1194
rect 3296 206 3308 1182
rect 3342 206 3354 1182
rect 3296 194 3354 206
<< mvpdiff >>
rect 136 2787 194 2799
rect 136 1811 148 2787
rect 182 1811 194 2787
rect 136 1799 194 1811
rect 294 2787 352 2799
rect 294 1811 306 2787
rect 340 1811 352 2787
rect 294 1799 352 1811
rect 452 2787 510 2799
rect 452 1811 464 2787
rect 498 1811 510 2787
rect 452 1799 510 1811
rect 610 2787 668 2799
rect 610 1811 622 2787
rect 656 1811 668 2787
rect 610 1799 668 1811
rect 768 2787 826 2799
rect 768 1811 780 2787
rect 814 1811 826 2787
rect 768 1799 826 1811
rect 926 2787 984 2799
rect 926 1811 938 2787
rect 972 1811 984 2787
rect 926 1799 984 1811
rect 1084 2787 1142 2799
rect 1084 1811 1096 2787
rect 1130 1811 1142 2787
rect 1084 1799 1142 1811
rect 1242 2787 1300 2799
rect 1242 1811 1254 2787
rect 1288 1811 1300 2787
rect 1242 1799 1300 1811
rect 1400 2787 1458 2799
rect 1400 1811 1412 2787
rect 1446 1811 1458 2787
rect 1400 1799 1458 1811
rect 1558 2787 1616 2799
rect 1558 1811 1570 2787
rect 1604 1811 1616 2787
rect 1558 1799 1616 1811
rect 1716 2787 1774 2799
rect 1716 1811 1728 2787
rect 1762 1811 1774 2787
rect 1716 1799 1774 1811
rect 1874 2787 1932 2799
rect 1874 1811 1886 2787
rect 1920 1811 1932 2787
rect 1874 1799 1932 1811
rect 2032 2787 2090 2799
rect 2032 1811 2044 2787
rect 2078 1811 2090 2787
rect 2032 1799 2090 1811
rect 2190 2787 2248 2799
rect 2190 1811 2202 2787
rect 2236 1811 2248 2787
rect 2190 1799 2248 1811
rect 2348 2787 2406 2799
rect 2348 1811 2360 2787
rect 2394 1811 2406 2787
rect 2348 1799 2406 1811
rect 2506 2787 2564 2799
rect 2506 1811 2518 2787
rect 2552 1811 2564 2787
rect 2506 1799 2564 1811
rect 2664 2787 2722 2799
rect 2664 1811 2676 2787
rect 2710 1811 2722 2787
rect 2664 1799 2722 1811
rect 2822 2787 2880 2799
rect 2822 1811 2834 2787
rect 2868 1811 2880 2787
rect 2822 1799 2880 1811
rect 2980 2787 3038 2799
rect 2980 1811 2992 2787
rect 3026 1811 3038 2787
rect 2980 1799 3038 1811
rect 3138 2787 3196 2799
rect 3138 1811 3150 2787
rect 3184 1811 3196 2787
rect 3138 1799 3196 1811
rect 3296 2787 3354 2799
rect 3296 1811 3308 2787
rect 3342 1811 3354 2787
rect 3296 1799 3354 1811
<< mvndiffc >>
rect 148 206 182 1182
rect 306 206 340 1182
rect 464 206 498 1182
rect 622 206 656 1182
rect 780 206 814 1182
rect 938 206 972 1182
rect 1096 206 1130 1182
rect 1254 206 1288 1182
rect 1412 206 1446 1182
rect 1570 206 1604 1182
rect 1728 206 1762 1182
rect 1886 206 1920 1182
rect 2044 206 2078 1182
rect 2202 206 2236 1182
rect 2360 206 2394 1182
rect 2518 206 2552 1182
rect 2676 206 2710 1182
rect 2834 206 2868 1182
rect 2992 206 3026 1182
rect 3150 206 3184 1182
rect 3308 206 3342 1182
<< mvpdiffc >>
rect 148 1811 182 2787
rect 306 1811 340 2787
rect 464 1811 498 2787
rect 622 1811 656 2787
rect 780 1811 814 2787
rect 938 1811 972 2787
rect 1096 1811 1130 2787
rect 1254 1811 1288 2787
rect 1412 1811 1446 2787
rect 1570 1811 1604 2787
rect 1728 1811 1762 2787
rect 1886 1811 1920 2787
rect 2044 1811 2078 2787
rect 2202 1811 2236 2787
rect 2360 1811 2394 2787
rect 2518 1811 2552 2787
rect 2676 1811 2710 2787
rect 2834 1811 2868 2787
rect 2992 1811 3026 2787
rect 3150 1811 3184 2787
rect 3308 1811 3342 2787
<< mvpsubdiff >>
rect 2 1404 3488 1416
rect 2 1370 110 1404
rect 3380 1370 3488 1404
rect 2 1358 3488 1370
rect 2 1308 60 1358
rect 2 80 14 1308
rect 48 80 60 1308
rect 3430 1308 3488 1358
rect 2 30 60 80
rect 3430 80 3442 1308
rect 3476 80 3488 1308
rect 3430 30 3488 80
rect 2 18 3488 30
rect 2 -16 110 18
rect 3380 -16 3488 18
rect 2 -28 3488 -16
<< mvnsubdiff >>
rect 2 3018 3488 3030
rect 2 2984 110 3018
rect 3380 2984 3488 3018
rect 2 2972 3488 2984
rect 2 2922 60 2972
rect 2 1676 14 2922
rect 48 1676 60 2922
rect 3430 2922 3488 2972
rect 2 1626 60 1676
rect 3430 1676 3442 2922
rect 3476 1676 3488 2922
rect 3430 1626 3488 1676
rect 2 1614 3488 1626
rect 2 1580 110 1614
rect 3380 1580 3488 1614
rect 2 1568 3488 1580
<< mvpsubdiffcont >>
rect 110 1370 3380 1404
rect 14 80 48 1308
rect 3442 80 3476 1308
rect 110 -16 3380 18
<< mvnsubdiffcont >>
rect 110 2984 3380 3018
rect 14 1676 48 2922
rect 3442 1676 3476 2922
rect 110 1580 3380 1614
<< poly >>
rect 194 2880 294 2896
rect 194 2846 210 2880
rect 278 2846 294 2880
rect 194 2799 294 2846
rect 352 2880 452 2896
rect 352 2846 368 2880
rect 436 2846 452 2880
rect 352 2799 452 2846
rect 510 2880 610 2896
rect 510 2846 526 2880
rect 594 2846 610 2880
rect 510 2799 610 2846
rect 668 2880 768 2896
rect 668 2846 684 2880
rect 752 2846 768 2880
rect 668 2799 768 2846
rect 826 2880 926 2896
rect 826 2846 842 2880
rect 910 2846 926 2880
rect 826 2799 926 2846
rect 984 2880 1084 2896
rect 984 2846 1000 2880
rect 1068 2846 1084 2880
rect 984 2799 1084 2846
rect 1142 2880 1242 2896
rect 1142 2846 1158 2880
rect 1226 2846 1242 2880
rect 1142 2799 1242 2846
rect 1300 2880 1400 2896
rect 1300 2846 1316 2880
rect 1384 2846 1400 2880
rect 1300 2799 1400 2846
rect 1458 2880 1558 2896
rect 1458 2846 1474 2880
rect 1542 2846 1558 2880
rect 1458 2799 1558 2846
rect 1616 2880 1716 2896
rect 1616 2846 1632 2880
rect 1700 2846 1716 2880
rect 1616 2799 1716 2846
rect 1774 2880 1874 2896
rect 1774 2846 1790 2880
rect 1858 2846 1874 2880
rect 1774 2799 1874 2846
rect 1932 2880 2032 2896
rect 1932 2846 1948 2880
rect 2016 2846 2032 2880
rect 1932 2799 2032 2846
rect 2090 2880 2190 2896
rect 2090 2846 2106 2880
rect 2174 2846 2190 2880
rect 2090 2799 2190 2846
rect 2248 2880 2348 2896
rect 2248 2846 2264 2880
rect 2332 2846 2348 2880
rect 2248 2799 2348 2846
rect 2406 2880 2506 2896
rect 2406 2846 2422 2880
rect 2490 2846 2506 2880
rect 2406 2799 2506 2846
rect 2564 2880 2664 2896
rect 2564 2846 2580 2880
rect 2648 2846 2664 2880
rect 2564 2799 2664 2846
rect 2722 2880 2822 2896
rect 2722 2846 2738 2880
rect 2806 2846 2822 2880
rect 2722 2799 2822 2846
rect 2880 2880 2980 2896
rect 2880 2846 2896 2880
rect 2964 2846 2980 2880
rect 2880 2799 2980 2846
rect 3038 2880 3138 2896
rect 3038 2846 3054 2880
rect 3122 2846 3138 2880
rect 3038 2799 3138 2846
rect 3196 2880 3296 2896
rect 3196 2846 3212 2880
rect 3280 2846 3296 2880
rect 3196 2799 3296 2846
rect 194 1752 294 1799
rect 194 1718 210 1752
rect 278 1718 294 1752
rect 194 1702 294 1718
rect 352 1752 452 1799
rect 352 1718 368 1752
rect 436 1718 452 1752
rect 352 1702 452 1718
rect 510 1752 610 1799
rect 510 1718 526 1752
rect 594 1718 610 1752
rect 510 1702 610 1718
rect 668 1752 768 1799
rect 668 1718 684 1752
rect 752 1718 768 1752
rect 668 1702 768 1718
rect 826 1752 926 1799
rect 826 1718 842 1752
rect 910 1718 926 1752
rect 826 1702 926 1718
rect 984 1752 1084 1799
rect 984 1718 1000 1752
rect 1068 1718 1084 1752
rect 984 1702 1084 1718
rect 1142 1752 1242 1799
rect 1142 1718 1158 1752
rect 1226 1718 1242 1752
rect 1142 1702 1242 1718
rect 1300 1752 1400 1799
rect 1300 1718 1316 1752
rect 1384 1718 1400 1752
rect 1300 1702 1400 1718
rect 1458 1752 1558 1799
rect 1458 1718 1474 1752
rect 1542 1718 1558 1752
rect 1458 1702 1558 1718
rect 1616 1752 1716 1799
rect 1616 1718 1632 1752
rect 1700 1718 1716 1752
rect 1616 1702 1716 1718
rect 1774 1752 1874 1799
rect 1774 1718 1790 1752
rect 1858 1718 1874 1752
rect 1774 1702 1874 1718
rect 1932 1752 2032 1799
rect 1932 1718 1948 1752
rect 2016 1718 2032 1752
rect 1932 1702 2032 1718
rect 2090 1752 2190 1799
rect 2090 1718 2106 1752
rect 2174 1718 2190 1752
rect 2090 1702 2190 1718
rect 2248 1752 2348 1799
rect 2248 1718 2264 1752
rect 2332 1718 2348 1752
rect 2248 1702 2348 1718
rect 2406 1752 2506 1799
rect 2406 1718 2422 1752
rect 2490 1718 2506 1752
rect 2406 1702 2506 1718
rect 2564 1752 2664 1799
rect 2564 1718 2580 1752
rect 2648 1718 2664 1752
rect 2564 1702 2664 1718
rect 2722 1752 2822 1799
rect 2722 1718 2738 1752
rect 2806 1718 2822 1752
rect 2722 1702 2822 1718
rect 2880 1752 2980 1799
rect 2880 1718 2896 1752
rect 2964 1718 2980 1752
rect 2880 1702 2980 1718
rect 3038 1752 3138 1799
rect 3038 1718 3054 1752
rect 3122 1718 3138 1752
rect 3038 1702 3138 1718
rect 3196 1752 3296 1799
rect 3196 1718 3212 1752
rect 3280 1718 3296 1752
rect 3196 1702 3296 1718
rect 194 1266 294 1282
rect 194 1232 210 1266
rect 278 1232 294 1266
rect 194 1194 294 1232
rect 352 1266 452 1282
rect 352 1232 368 1266
rect 436 1232 452 1266
rect 352 1194 452 1232
rect 510 1266 610 1282
rect 510 1232 526 1266
rect 594 1232 610 1266
rect 510 1194 610 1232
rect 668 1266 768 1282
rect 668 1232 684 1266
rect 752 1232 768 1266
rect 668 1194 768 1232
rect 826 1266 926 1282
rect 826 1232 842 1266
rect 910 1232 926 1266
rect 826 1194 926 1232
rect 984 1266 1084 1282
rect 984 1232 1000 1266
rect 1068 1232 1084 1266
rect 984 1194 1084 1232
rect 1142 1266 1242 1282
rect 1142 1232 1158 1266
rect 1226 1232 1242 1266
rect 1142 1194 1242 1232
rect 1300 1266 1400 1282
rect 1300 1232 1316 1266
rect 1384 1232 1400 1266
rect 1300 1194 1400 1232
rect 1458 1266 1558 1282
rect 1458 1232 1474 1266
rect 1542 1232 1558 1266
rect 1458 1194 1558 1232
rect 1616 1266 1716 1282
rect 1616 1232 1632 1266
rect 1700 1232 1716 1266
rect 1616 1194 1716 1232
rect 1774 1266 1874 1282
rect 1774 1232 1790 1266
rect 1858 1232 1874 1266
rect 1774 1194 1874 1232
rect 1932 1266 2032 1282
rect 1932 1232 1948 1266
rect 2016 1232 2032 1266
rect 1932 1194 2032 1232
rect 2090 1266 2190 1282
rect 2090 1232 2106 1266
rect 2174 1232 2190 1266
rect 2090 1194 2190 1232
rect 2248 1266 2348 1282
rect 2248 1232 2264 1266
rect 2332 1232 2348 1266
rect 2248 1194 2348 1232
rect 2406 1266 2506 1282
rect 2406 1232 2422 1266
rect 2490 1232 2506 1266
rect 2406 1194 2506 1232
rect 2564 1266 2664 1282
rect 2564 1232 2580 1266
rect 2648 1232 2664 1266
rect 2564 1194 2664 1232
rect 2722 1266 2822 1282
rect 2722 1232 2738 1266
rect 2806 1232 2822 1266
rect 2722 1194 2822 1232
rect 2880 1266 2980 1282
rect 2880 1232 2896 1266
rect 2964 1232 2980 1266
rect 2880 1194 2980 1232
rect 3038 1266 3138 1282
rect 3038 1232 3054 1266
rect 3122 1232 3138 1266
rect 3038 1194 3138 1232
rect 3196 1266 3296 1282
rect 3196 1232 3212 1266
rect 3280 1232 3296 1266
rect 3196 1194 3296 1232
rect 194 156 294 194
rect 194 122 210 156
rect 278 122 294 156
rect 194 106 294 122
rect 352 156 452 194
rect 352 122 368 156
rect 436 122 452 156
rect 352 106 452 122
rect 510 156 610 194
rect 510 122 526 156
rect 594 122 610 156
rect 510 106 610 122
rect 668 156 768 194
rect 668 122 684 156
rect 752 122 768 156
rect 668 106 768 122
rect 826 156 926 194
rect 826 122 842 156
rect 910 122 926 156
rect 826 106 926 122
rect 984 156 1084 194
rect 984 122 1000 156
rect 1068 122 1084 156
rect 984 106 1084 122
rect 1142 156 1242 194
rect 1142 122 1158 156
rect 1226 122 1242 156
rect 1142 106 1242 122
rect 1300 156 1400 194
rect 1300 122 1316 156
rect 1384 122 1400 156
rect 1300 106 1400 122
rect 1458 156 1558 194
rect 1458 122 1474 156
rect 1542 122 1558 156
rect 1458 106 1558 122
rect 1616 156 1716 194
rect 1616 122 1632 156
rect 1700 122 1716 156
rect 1616 106 1716 122
rect 1774 156 1874 194
rect 1774 122 1790 156
rect 1858 122 1874 156
rect 1774 106 1874 122
rect 1932 156 2032 194
rect 1932 122 1948 156
rect 2016 122 2032 156
rect 1932 106 2032 122
rect 2090 156 2190 194
rect 2090 122 2106 156
rect 2174 122 2190 156
rect 2090 106 2190 122
rect 2248 156 2348 194
rect 2248 122 2264 156
rect 2332 122 2348 156
rect 2248 106 2348 122
rect 2406 156 2506 194
rect 2406 122 2422 156
rect 2490 122 2506 156
rect 2406 106 2506 122
rect 2564 156 2664 194
rect 2564 122 2580 156
rect 2648 122 2664 156
rect 2564 106 2664 122
rect 2722 156 2822 194
rect 2722 122 2738 156
rect 2806 122 2822 156
rect 2722 106 2822 122
rect 2880 156 2980 194
rect 2880 122 2896 156
rect 2964 122 2980 156
rect 2880 106 2980 122
rect 3038 156 3138 194
rect 3038 122 3054 156
rect 3122 122 3138 156
rect 3038 106 3138 122
rect 3196 156 3296 194
rect 3196 122 3212 156
rect 3280 122 3296 156
rect 3196 106 3296 122
<< polycont >>
rect 210 2846 278 2880
rect 368 2846 436 2880
rect 526 2846 594 2880
rect 684 2846 752 2880
rect 842 2846 910 2880
rect 1000 2846 1068 2880
rect 1158 2846 1226 2880
rect 1316 2846 1384 2880
rect 1474 2846 1542 2880
rect 1632 2846 1700 2880
rect 1790 2846 1858 2880
rect 1948 2846 2016 2880
rect 2106 2846 2174 2880
rect 2264 2846 2332 2880
rect 2422 2846 2490 2880
rect 2580 2846 2648 2880
rect 2738 2846 2806 2880
rect 2896 2846 2964 2880
rect 3054 2846 3122 2880
rect 3212 2846 3280 2880
rect 210 1718 278 1752
rect 368 1718 436 1752
rect 526 1718 594 1752
rect 684 1718 752 1752
rect 842 1718 910 1752
rect 1000 1718 1068 1752
rect 1158 1718 1226 1752
rect 1316 1718 1384 1752
rect 1474 1718 1542 1752
rect 1632 1718 1700 1752
rect 1790 1718 1858 1752
rect 1948 1718 2016 1752
rect 2106 1718 2174 1752
rect 2264 1718 2332 1752
rect 2422 1718 2490 1752
rect 2580 1718 2648 1752
rect 2738 1718 2806 1752
rect 2896 1718 2964 1752
rect 3054 1718 3122 1752
rect 3212 1718 3280 1752
rect 210 1232 278 1266
rect 368 1232 436 1266
rect 526 1232 594 1266
rect 684 1232 752 1266
rect 842 1232 910 1266
rect 1000 1232 1068 1266
rect 1158 1232 1226 1266
rect 1316 1232 1384 1266
rect 1474 1232 1542 1266
rect 1632 1232 1700 1266
rect 1790 1232 1858 1266
rect 1948 1232 2016 1266
rect 2106 1232 2174 1266
rect 2264 1232 2332 1266
rect 2422 1232 2490 1266
rect 2580 1232 2648 1266
rect 2738 1232 2806 1266
rect 2896 1232 2964 1266
rect 3054 1232 3122 1266
rect 3212 1232 3280 1266
rect 210 122 278 156
rect 368 122 436 156
rect 526 122 594 156
rect 684 122 752 156
rect 842 122 910 156
rect 1000 122 1068 156
rect 1158 122 1226 156
rect 1316 122 1384 156
rect 1474 122 1542 156
rect 1632 122 1700 156
rect 1790 122 1858 156
rect 1948 122 2016 156
rect 2106 122 2174 156
rect 2264 122 2332 156
rect 2422 122 2490 156
rect 2580 122 2648 156
rect 2738 122 2806 156
rect 2896 122 2964 156
rect 3054 122 3122 156
rect 3212 122 3280 156
<< locali >>
rect 14 2984 110 3018
rect 3380 2984 3476 3018
rect 14 2922 48 2984
rect 3442 2922 3476 2984
rect 194 2846 210 2880
rect 278 2846 294 2880
rect 352 2846 368 2880
rect 436 2846 452 2880
rect 510 2846 526 2880
rect 594 2846 610 2880
rect 668 2846 684 2880
rect 752 2846 768 2880
rect 826 2846 842 2880
rect 910 2846 926 2880
rect 984 2846 1000 2880
rect 1068 2846 1084 2880
rect 1142 2846 1158 2880
rect 1226 2846 1242 2880
rect 1300 2846 1316 2880
rect 1384 2846 1400 2880
rect 1458 2846 1474 2880
rect 1542 2846 1558 2880
rect 1616 2846 1632 2880
rect 1700 2846 1716 2880
rect 1774 2846 1790 2880
rect 1858 2846 1874 2880
rect 1932 2846 1948 2880
rect 2016 2846 2032 2880
rect 2090 2846 2106 2880
rect 2174 2846 2190 2880
rect 2248 2846 2264 2880
rect 2332 2846 2348 2880
rect 2406 2846 2422 2880
rect 2490 2846 2506 2880
rect 2564 2846 2580 2880
rect 2648 2846 2664 2880
rect 2722 2846 2738 2880
rect 2806 2846 2822 2880
rect 2880 2846 2896 2880
rect 2964 2846 2980 2880
rect 3038 2846 3054 2880
rect 3122 2846 3138 2880
rect 3196 2846 3212 2880
rect 3280 2846 3296 2880
rect 148 2787 182 2803
rect 148 1795 182 1811
rect 306 2787 340 2803
rect 306 1795 340 1811
rect 464 2787 498 2803
rect 464 1795 498 1811
rect 622 2787 656 2803
rect 622 1795 656 1811
rect 780 2787 814 2803
rect 780 1795 814 1811
rect 938 2787 972 2803
rect 938 1795 972 1811
rect 1096 2787 1130 2803
rect 1096 1795 1130 1811
rect 1254 2787 1288 2803
rect 1254 1795 1288 1811
rect 1412 2787 1446 2803
rect 1412 1795 1446 1811
rect 1570 2787 1604 2803
rect 1570 1795 1604 1811
rect 1728 2787 1762 2803
rect 1728 1795 1762 1811
rect 1886 2787 1920 2803
rect 1886 1795 1920 1811
rect 2044 2787 2078 2803
rect 2044 1795 2078 1811
rect 2202 2787 2236 2803
rect 2202 1795 2236 1811
rect 2360 2787 2394 2803
rect 2360 1795 2394 1811
rect 2518 2787 2552 2803
rect 2518 1795 2552 1811
rect 2676 2787 2710 2803
rect 2676 1795 2710 1811
rect 2834 2787 2868 2803
rect 2834 1795 2868 1811
rect 2992 2787 3026 2803
rect 2992 1795 3026 1811
rect 3150 2787 3184 2803
rect 3150 1795 3184 1811
rect 3308 2787 3342 2803
rect 3308 1795 3342 1811
rect 194 1718 210 1752
rect 278 1718 294 1752
rect 352 1718 368 1752
rect 436 1718 452 1752
rect 510 1718 526 1752
rect 594 1718 610 1752
rect 668 1718 684 1752
rect 752 1718 768 1752
rect 826 1718 842 1752
rect 910 1718 926 1752
rect 984 1718 1000 1752
rect 1068 1718 1084 1752
rect 1142 1718 1158 1752
rect 1226 1718 1242 1752
rect 1300 1718 1316 1752
rect 1384 1718 1400 1752
rect 1458 1718 1474 1752
rect 1542 1718 1558 1752
rect 1616 1718 1632 1752
rect 1700 1718 1716 1752
rect 1774 1718 1790 1752
rect 1858 1718 1874 1752
rect 1932 1718 1948 1752
rect 2016 1718 2032 1752
rect 2090 1718 2106 1752
rect 2174 1718 2190 1752
rect 2248 1718 2264 1752
rect 2332 1718 2348 1752
rect 2406 1718 2422 1752
rect 2490 1718 2506 1752
rect 2564 1718 2580 1752
rect 2648 1718 2664 1752
rect 2722 1718 2738 1752
rect 2806 1718 2822 1752
rect 2880 1718 2896 1752
rect 2964 1718 2980 1752
rect 3038 1718 3054 1752
rect 3122 1718 3138 1752
rect 3196 1718 3212 1752
rect 3280 1718 3296 1752
rect 14 1614 48 1676
rect 3442 1614 3476 1676
rect 14 1580 110 1614
rect 3380 1580 3476 1614
rect 14 1370 110 1404
rect 3380 1370 3476 1404
rect 14 1308 48 1370
rect 3442 1308 3476 1370
rect 194 1232 210 1266
rect 278 1232 294 1266
rect 352 1232 368 1266
rect 436 1232 452 1266
rect 510 1232 526 1266
rect 594 1232 610 1266
rect 668 1232 684 1266
rect 752 1232 768 1266
rect 826 1232 842 1266
rect 910 1232 926 1266
rect 984 1232 1000 1266
rect 1068 1232 1084 1266
rect 1142 1232 1158 1266
rect 1226 1232 1242 1266
rect 1300 1232 1316 1266
rect 1384 1232 1400 1266
rect 1458 1232 1474 1266
rect 1542 1232 1558 1266
rect 1616 1232 1632 1266
rect 1700 1232 1716 1266
rect 1774 1232 1790 1266
rect 1858 1232 1874 1266
rect 1932 1232 1948 1266
rect 2016 1232 2032 1266
rect 2090 1232 2106 1266
rect 2174 1232 2190 1266
rect 2248 1232 2264 1266
rect 2332 1232 2348 1266
rect 2406 1232 2422 1266
rect 2490 1232 2506 1266
rect 2564 1232 2580 1266
rect 2648 1232 2664 1266
rect 2722 1232 2738 1266
rect 2806 1232 2822 1266
rect 2880 1232 2896 1266
rect 2964 1232 2980 1266
rect 3038 1232 3054 1266
rect 3122 1232 3138 1266
rect 3196 1232 3212 1266
rect 3280 1232 3296 1266
rect 148 1182 182 1198
rect 148 190 182 206
rect 306 1182 340 1198
rect 306 190 340 206
rect 464 1182 498 1198
rect 464 190 498 206
rect 622 1182 656 1198
rect 622 190 656 206
rect 780 1182 814 1198
rect 780 190 814 206
rect 938 1182 972 1198
rect 938 190 972 206
rect 1096 1182 1130 1198
rect 1096 190 1130 206
rect 1254 1182 1288 1198
rect 1254 190 1288 206
rect 1412 1182 1446 1198
rect 1412 190 1446 206
rect 1570 1182 1604 1198
rect 1570 190 1604 206
rect 1728 1182 1762 1198
rect 1728 190 1762 206
rect 1886 1182 1920 1198
rect 1886 190 1920 206
rect 2044 1182 2078 1198
rect 2044 190 2078 206
rect 2202 1182 2236 1198
rect 2202 190 2236 206
rect 2360 1182 2394 1198
rect 2360 190 2394 206
rect 2518 1182 2552 1198
rect 2518 190 2552 206
rect 2676 1182 2710 1198
rect 2676 190 2710 206
rect 2834 1182 2868 1198
rect 2834 190 2868 206
rect 2992 1182 3026 1198
rect 2992 190 3026 206
rect 3150 1182 3184 1198
rect 3150 190 3184 206
rect 3308 1182 3342 1198
rect 3308 190 3342 206
rect 194 122 210 156
rect 278 122 294 156
rect 352 122 368 156
rect 436 122 452 156
rect 510 122 526 156
rect 594 122 610 156
rect 668 122 684 156
rect 752 122 768 156
rect 826 122 842 156
rect 910 122 926 156
rect 984 122 1000 156
rect 1068 122 1084 156
rect 1142 122 1158 156
rect 1226 122 1242 156
rect 1300 122 1316 156
rect 1384 122 1400 156
rect 1458 122 1474 156
rect 1542 122 1558 156
rect 1616 122 1632 156
rect 1700 122 1716 156
rect 1774 122 1790 156
rect 1858 122 1874 156
rect 1932 122 1948 156
rect 2016 122 2032 156
rect 2090 122 2106 156
rect 2174 122 2190 156
rect 2248 122 2264 156
rect 2332 122 2348 156
rect 2406 122 2422 156
rect 2490 122 2506 156
rect 2564 122 2580 156
rect 2648 122 2664 156
rect 2722 122 2738 156
rect 2806 122 2822 156
rect 2880 122 2896 156
rect 2964 122 2980 156
rect 3038 122 3054 156
rect 3122 122 3138 156
rect 3196 122 3212 156
rect 3280 122 3296 156
rect 14 18 48 80
rect 3442 18 3476 80
rect 14 -16 110 18
rect 3380 -16 3476 18
<< viali >>
rect 110 2984 3380 3018
rect 14 1676 48 2922
rect 226 2846 260 2880
rect 384 2846 418 2880
rect 542 2846 576 2880
rect 700 2846 734 2880
rect 858 2846 892 2880
rect 1016 2846 1050 2880
rect 1174 2846 1208 2880
rect 1332 2846 1366 2880
rect 1490 2846 1524 2880
rect 1648 2846 1682 2880
rect 1808 2846 1842 2880
rect 1966 2846 2000 2880
rect 2124 2846 2158 2880
rect 2282 2846 2316 2880
rect 2440 2846 2474 2880
rect 2598 2846 2632 2880
rect 2756 2846 2790 2880
rect 2914 2846 2948 2880
rect 3072 2846 3106 2880
rect 3230 2846 3264 2880
rect 148 1811 182 2787
rect 306 1811 340 2787
rect 464 1811 498 2787
rect 622 1811 656 2787
rect 780 1811 814 2787
rect 938 1811 972 2787
rect 1096 1811 1130 2787
rect 1254 1811 1288 2787
rect 1412 1811 1446 2787
rect 1570 1811 1604 2787
rect 1728 1811 1762 2787
rect 1886 1811 1920 2787
rect 2044 1811 2078 2787
rect 2202 1811 2236 2787
rect 2360 1811 2394 2787
rect 2518 1811 2552 2787
rect 2676 1811 2710 2787
rect 2834 1811 2868 2787
rect 2992 1811 3026 2787
rect 3150 1811 3184 2787
rect 3308 1811 3342 2787
rect 226 1718 260 1752
rect 384 1718 418 1752
rect 542 1718 576 1752
rect 700 1718 734 1752
rect 858 1718 892 1752
rect 1016 1718 1050 1752
rect 1174 1718 1208 1752
rect 1332 1718 1366 1752
rect 1490 1718 1524 1752
rect 1648 1718 1682 1752
rect 1808 1718 1842 1752
rect 1966 1718 2000 1752
rect 2124 1718 2158 1752
rect 2282 1718 2316 1752
rect 2440 1718 2474 1752
rect 2598 1718 2632 1752
rect 2756 1718 2790 1752
rect 2914 1718 2948 1752
rect 3072 1718 3106 1752
rect 3230 1718 3264 1752
rect 3442 1676 3476 2922
rect 14 80 48 1308
rect 226 1232 260 1266
rect 384 1232 418 1266
rect 542 1232 576 1266
rect 700 1232 734 1266
rect 858 1232 892 1266
rect 1016 1232 1050 1266
rect 1174 1232 1208 1266
rect 1332 1232 1366 1266
rect 1490 1232 1524 1266
rect 1648 1232 1682 1266
rect 1808 1232 1842 1266
rect 1966 1232 2000 1266
rect 2124 1232 2158 1266
rect 2282 1232 2316 1266
rect 2440 1232 2474 1266
rect 2598 1232 2632 1266
rect 2756 1232 2790 1266
rect 2914 1232 2948 1266
rect 3072 1232 3106 1266
rect 3230 1232 3264 1266
rect 148 206 182 1182
rect 306 206 340 1182
rect 464 206 498 1182
rect 622 206 656 1182
rect 780 206 814 1182
rect 938 206 972 1182
rect 1096 206 1130 1182
rect 1254 206 1288 1182
rect 1412 206 1446 1182
rect 1570 206 1604 1182
rect 1728 206 1762 1182
rect 1886 206 1920 1182
rect 2044 206 2078 1182
rect 2202 206 2236 1182
rect 2360 206 2394 1182
rect 2518 206 2552 1182
rect 2676 206 2710 1182
rect 2834 206 2868 1182
rect 2992 206 3026 1182
rect 3150 206 3184 1182
rect 3308 206 3342 1182
rect 226 122 260 156
rect 384 122 418 156
rect 542 122 576 156
rect 700 122 734 156
rect 858 122 892 156
rect 1016 122 1050 156
rect 1174 122 1208 156
rect 1332 122 1366 156
rect 1490 122 1524 156
rect 1648 122 1682 156
rect 1808 122 1842 156
rect 1966 122 2000 156
rect 2124 122 2158 156
rect 2282 122 2316 156
rect 2440 122 2474 156
rect 2598 122 2632 156
rect 2756 122 2790 156
rect 2914 122 2948 156
rect 3072 122 3106 156
rect 3230 122 3264 156
rect 3442 80 3476 1308
rect 110 -16 3380 18
<< metal1 >>
rect 8 3018 3482 3024
rect 8 2984 110 3018
rect 3380 2984 3482 3018
rect 8 2922 3482 2984
rect 8 1676 14 2922
rect 48 2880 3442 2922
rect 48 2846 226 2880
rect 260 2846 384 2880
rect 418 2846 542 2880
rect 576 2846 700 2880
rect 734 2846 858 2880
rect 892 2846 1016 2880
rect 1050 2846 1174 2880
rect 1208 2846 1332 2880
rect 1366 2846 1490 2880
rect 1524 2846 1648 2880
rect 1682 2846 1808 2880
rect 1842 2846 1966 2880
rect 2000 2846 2124 2880
rect 2158 2846 2282 2880
rect 2316 2846 2440 2880
rect 2474 2846 2598 2880
rect 2632 2846 2756 2880
rect 2790 2846 2914 2880
rect 2948 2846 3072 2880
rect 3106 2846 3230 2880
rect 3264 2846 3442 2880
rect 48 2840 3442 2846
rect 48 1758 60 2840
rect 142 2787 188 2840
rect 300 2787 346 2799
rect 458 2787 504 2840
rect 616 2787 662 2799
rect 774 2787 820 2840
rect 932 2787 978 2799
rect 1090 2787 1136 2840
rect 1248 2787 1294 2799
rect 1406 2787 1452 2840
rect 1564 2787 1610 2799
rect 1722 2787 1768 2840
rect 1880 2787 1926 2799
rect 2038 2787 2084 2840
rect 2196 2787 2242 2799
rect 2354 2787 2400 2840
rect 2512 2787 2558 2799
rect 2670 2787 2716 2840
rect 2828 2787 2874 2799
rect 2986 2787 3032 2840
rect 3144 2787 3190 2799
rect 3302 2787 3348 2840
rect 142 1811 148 2787
rect 182 1811 188 2787
rect 287 1811 297 2787
rect 349 1811 359 2787
rect 458 1811 464 2787
rect 498 1811 504 2787
rect 603 1811 613 2787
rect 665 1811 675 2787
rect 774 1811 780 2787
rect 814 1811 820 2787
rect 919 1811 929 2787
rect 981 1811 991 2787
rect 1090 1811 1096 2787
rect 1130 1811 1136 2787
rect 1235 1811 1245 2787
rect 1297 1811 1307 2787
rect 1406 1811 1412 2787
rect 1446 1811 1452 2787
rect 1551 1811 1561 2787
rect 1613 1811 1623 2787
rect 1722 1811 1728 2787
rect 1762 1811 1768 2787
rect 1867 1811 1877 2787
rect 1929 1811 1939 2787
rect 2038 1811 2044 2787
rect 2078 1811 2084 2787
rect 2183 1811 2193 2787
rect 2245 1811 2255 2787
rect 2354 1811 2360 2787
rect 2394 1811 2400 2787
rect 2499 1811 2509 2787
rect 2561 1811 2571 2787
rect 2670 1811 2676 2787
rect 2710 1811 2716 2787
rect 2815 1811 2825 2787
rect 2877 1811 2887 2787
rect 2986 1811 2992 2787
rect 3026 1811 3032 2787
rect 3131 1811 3141 2787
rect 3193 1811 3203 2787
rect 3302 1811 3308 2787
rect 3342 1811 3348 2787
rect 142 1758 188 1811
rect 300 1799 346 1811
rect 458 1799 504 1811
rect 616 1799 662 1811
rect 774 1799 820 1811
rect 932 1799 978 1811
rect 1090 1799 1136 1811
rect 1248 1799 1294 1811
rect 1406 1799 1452 1811
rect 1564 1799 1610 1811
rect 1722 1799 1768 1811
rect 1880 1799 1926 1811
rect 2038 1799 2084 1811
rect 2196 1799 2242 1811
rect 2354 1799 2400 1811
rect 2512 1799 2558 1811
rect 2670 1799 2716 1811
rect 2828 1799 2874 1811
rect 2986 1799 3032 1811
rect 3144 1799 3190 1811
rect 3302 1758 3348 1811
rect 3430 1758 3442 2840
rect 48 1752 3442 1758
rect 48 1718 226 1752
rect 260 1718 384 1752
rect 418 1718 542 1752
rect 576 1718 700 1752
rect 734 1718 858 1752
rect 892 1718 1016 1752
rect 1050 1718 1174 1752
rect 1208 1718 1332 1752
rect 1366 1718 1490 1752
rect 1524 1718 1648 1752
rect 1682 1718 1808 1752
rect 1842 1718 1966 1752
rect 2000 1718 2124 1752
rect 2158 1718 2282 1752
rect 2316 1718 2440 1752
rect 2474 1718 2598 1752
rect 2632 1718 2756 1752
rect 2790 1718 2914 1752
rect 2948 1718 3072 1752
rect 3106 1718 3230 1752
rect 3264 1718 3442 1752
rect 48 1712 3442 1718
rect 48 1676 54 1712
rect 8 1664 54 1676
rect 3436 1676 3442 1712
rect 3476 1676 3482 2922
rect 3436 1664 3482 1676
rect -64 1545 3554 1556
rect -64 1441 297 1545
rect 349 1441 613 1545
rect 665 1441 929 1545
rect 981 1441 1245 1545
rect 1297 1441 1561 1545
rect 1613 1441 1877 1545
rect 1929 1441 2193 1545
rect 2245 1441 2509 1545
rect 2561 1441 2825 1545
rect 2877 1441 3141 1545
rect 3193 1441 3554 1545
rect -64 1428 3554 1441
rect 8 1308 54 1320
rect 8 80 14 1308
rect 48 1272 54 1308
rect 3436 1308 3482 1320
rect 3436 1272 3442 1308
rect 48 1266 3442 1272
rect 48 1232 226 1266
rect 260 1232 384 1266
rect 418 1232 542 1266
rect 576 1232 700 1266
rect 734 1232 858 1266
rect 892 1232 1016 1266
rect 1050 1232 1174 1266
rect 1208 1232 1332 1266
rect 1366 1232 1490 1266
rect 1524 1232 1648 1266
rect 1682 1232 1808 1266
rect 1842 1232 1966 1266
rect 2000 1232 2124 1266
rect 2158 1232 2282 1266
rect 2316 1232 2440 1266
rect 2474 1232 2598 1266
rect 2632 1232 2756 1266
rect 2790 1232 2914 1266
rect 2948 1232 3072 1266
rect 3106 1232 3230 1266
rect 3264 1232 3442 1266
rect 48 1226 3442 1232
rect 48 162 54 1226
rect 142 1182 188 1194
rect 300 1182 346 1194
rect 458 1182 504 1194
rect 616 1182 662 1194
rect 774 1182 820 1194
rect 932 1182 978 1194
rect 1090 1182 1136 1194
rect 1248 1182 1294 1194
rect 1406 1182 1452 1194
rect 1564 1182 1610 1194
rect 1722 1182 1768 1194
rect 1880 1182 1926 1194
rect 2038 1182 2084 1194
rect 2196 1182 2242 1194
rect 2354 1182 2400 1194
rect 2512 1182 2558 1194
rect 2670 1182 2716 1194
rect 2828 1182 2874 1194
rect 2986 1182 3032 1194
rect 3144 1182 3190 1194
rect 3302 1182 3348 1226
rect 142 206 148 1182
rect 182 206 188 1182
rect 287 206 297 1182
rect 349 206 359 1182
rect 458 206 464 1182
rect 498 206 504 1182
rect 603 206 613 1182
rect 665 206 675 1182
rect 774 206 780 1182
rect 814 206 820 1182
rect 919 206 929 1182
rect 981 206 991 1182
rect 1090 206 1096 1182
rect 1130 206 1136 1182
rect 1235 206 1245 1182
rect 1297 206 1307 1182
rect 1406 206 1412 1182
rect 1446 206 1452 1182
rect 1551 206 1561 1182
rect 1613 206 1623 1182
rect 1722 206 1728 1182
rect 1762 206 1768 1182
rect 1867 206 1877 1182
rect 1929 206 1939 1182
rect 2038 206 2044 1182
rect 2078 206 2084 1182
rect 2183 206 2193 1182
rect 2245 206 2255 1182
rect 2354 206 2360 1182
rect 2394 206 2400 1182
rect 2499 206 2509 1182
rect 2561 206 2571 1182
rect 2670 206 2676 1182
rect 2710 206 2716 1182
rect 2815 206 2825 1182
rect 2877 206 2887 1182
rect 2986 206 2992 1182
rect 3026 206 3032 1182
rect 3131 206 3141 1182
rect 3193 206 3203 1182
rect 3302 206 3308 1182
rect 3342 206 3348 1182
rect 142 162 188 206
rect 300 194 346 206
rect 458 162 504 206
rect 616 194 662 206
rect 774 162 820 206
rect 932 194 978 206
rect 1090 162 1136 206
rect 1248 194 1294 206
rect 1406 162 1452 206
rect 1564 194 1610 206
rect 1722 162 1768 206
rect 1880 194 1926 206
rect 2038 162 2084 206
rect 2196 194 2242 206
rect 2354 162 2400 206
rect 2512 194 2558 206
rect 2670 162 2716 206
rect 2828 194 2874 206
rect 2986 162 3032 206
rect 3144 194 3190 206
rect 3302 162 3348 206
rect 3436 162 3442 1226
rect 48 156 3442 162
rect 48 122 226 156
rect 260 122 384 156
rect 418 122 542 156
rect 576 122 700 156
rect 734 122 858 156
rect 892 122 1016 156
rect 1050 122 1174 156
rect 1208 122 1332 156
rect 1366 122 1490 156
rect 1524 122 1648 156
rect 1682 122 1808 156
rect 1842 122 1966 156
rect 2000 122 2124 156
rect 2158 122 2282 156
rect 2316 122 2440 156
rect 2474 122 2598 156
rect 2632 122 2756 156
rect 2790 122 2914 156
rect 2948 122 3072 156
rect 3106 122 3230 156
rect 3264 122 3442 156
rect 48 80 3442 122
rect 3476 80 3482 1308
rect 8 18 3482 80
rect 8 -16 110 18
rect 3380 -16 3482 18
rect 8 -22 3482 -16
<< via1 >>
rect 297 1811 306 2787
rect 306 1811 340 2787
rect 340 1811 349 2787
rect 613 1811 622 2787
rect 622 1811 656 2787
rect 656 1811 665 2787
rect 929 1811 938 2787
rect 938 1811 972 2787
rect 972 1811 981 2787
rect 1245 1811 1254 2787
rect 1254 1811 1288 2787
rect 1288 1811 1297 2787
rect 1561 1811 1570 2787
rect 1570 1811 1604 2787
rect 1604 1811 1613 2787
rect 1877 1811 1886 2787
rect 1886 1811 1920 2787
rect 1920 1811 1929 2787
rect 2193 1811 2202 2787
rect 2202 1811 2236 2787
rect 2236 1811 2245 2787
rect 2509 1811 2518 2787
rect 2518 1811 2552 2787
rect 2552 1811 2561 2787
rect 2825 1811 2834 2787
rect 2834 1811 2868 2787
rect 2868 1811 2877 2787
rect 3141 1811 3150 2787
rect 3150 1811 3184 2787
rect 3184 1811 3193 2787
rect 297 1441 349 1545
rect 613 1441 665 1545
rect 929 1441 981 1545
rect 1245 1441 1297 1545
rect 1561 1441 1613 1545
rect 1877 1441 1929 1545
rect 2193 1441 2245 1545
rect 2509 1441 2561 1545
rect 2825 1441 2877 1545
rect 3141 1441 3193 1545
rect 297 206 306 1182
rect 306 206 340 1182
rect 340 206 349 1182
rect 613 206 622 1182
rect 622 206 656 1182
rect 656 206 665 1182
rect 929 206 938 1182
rect 938 206 972 1182
rect 972 206 981 1182
rect 1245 206 1254 1182
rect 1254 206 1288 1182
rect 1288 206 1297 1182
rect 1561 206 1570 1182
rect 1570 206 1604 1182
rect 1604 206 1613 1182
rect 1877 206 1886 1182
rect 1886 206 1920 1182
rect 1920 206 1929 1182
rect 2193 206 2202 1182
rect 2202 206 2236 1182
rect 2236 206 2245 1182
rect 2509 206 2518 1182
rect 2518 206 2552 1182
rect 2552 206 2561 1182
rect 2825 206 2834 1182
rect 2834 206 2868 1182
rect 2868 206 2877 1182
rect 3141 206 3150 1182
rect 3150 206 3184 1182
rect 3184 206 3193 1182
<< metal2 >>
rect 297 2787 349 2797
rect 297 1545 349 1811
rect 297 1182 349 1441
rect 297 196 349 206
rect 613 2787 665 2797
rect 613 1545 665 1811
rect 613 1182 665 1441
rect 613 196 665 206
rect 929 2787 981 2797
rect 929 1545 981 1811
rect 929 1182 981 1441
rect 929 196 981 206
rect 1245 2787 1297 2797
rect 1245 1545 1297 1811
rect 1245 1182 1297 1441
rect 1245 196 1297 206
rect 1561 2787 1613 2797
rect 1561 1545 1613 1811
rect 1561 1182 1613 1441
rect 1561 196 1613 206
rect 1877 2787 1929 2797
rect 1877 1545 1929 1811
rect 1877 1182 1929 1441
rect 1877 196 1929 206
rect 2193 2787 2245 2797
rect 2193 1545 2245 1811
rect 2193 1182 2245 1441
rect 2193 196 2245 206
rect 2509 2787 2561 2797
rect 2509 1545 2561 1811
rect 2509 1182 2561 1441
rect 2509 196 2561 206
rect 2825 2787 2877 2797
rect 2825 1545 2877 1811
rect 2825 1182 2877 1441
rect 2825 196 2877 206
rect 3141 2787 3193 2797
rect 3141 1545 3193 1811
rect 3141 1182 3193 1441
rect 3141 196 3193 206
<< labels >>
flabel metal1 -53 1488 -53 1488 1 FreeSans 400 0 0 0 esd
port 1 n
flabel metal1 31 2928 31 2928 1 FreeSans 400 0 0 0 VDD
port 2 n power bidirectional
flabel metal1 31 72 31 72 1 FreeSans 400 0 0 0 VSS
port 3 n power bidirectional
<< end >>
