magic
tech sky130A
magscale 1 2
timestamp 1653995921
<< nwell >>
rect -3035 -295 16729 26
rect -3035 -1383 16729 -817
rect -3035 -2471 16729 -1905
rect -3035 -3559 16729 -2993
rect -3035 -4647 16729 -4081
rect -3035 -5735 16729 -5169
rect -3035 -6823 16729 -6257
rect -3035 -7911 16729 -7345
rect -3035 -8999 16729 -8433
rect -3035 -10087 16729 -9521
rect -3035 -11175 16729 -10609
rect -3035 -12263 16729 -11697
rect -3035 -13351 16729 -12785
rect -3035 -14194 16729 -13873
<< pwell >>
rect -968 -360 -698 -353
rect 2446 -360 2958 -353
rect 6954 -360 7466 -353
rect 8242 -360 8754 -353
rect 9530 -360 10042 -353
rect 10712 -360 11486 -353
rect -3035 -508 16728 -360
rect -2996 -535 -2262 -508
rect -2258 -518 -2172 -508
rect -1432 -535 -1066 -508
rect -1062 -518 -976 -508
rect -968 -535 -698 -508
rect -694 -518 -608 -508
rect -604 -535 -238 -508
rect -234 -518 -148 -508
rect -63 -535 422 -508
rect 502 -518 588 -508
rect 592 -535 958 -508
rect 962 -518 1048 -508
rect 1135 -535 1326 -508
rect 1330 -518 1416 -508
rect 1420 -535 1786 -508
rect 1790 -518 1876 -508
rect 1880 -535 2246 -508
rect 2250 -518 2336 -508
rect 2340 -535 3074 -508
rect 3078 -518 3164 -508
rect 3168 -535 3534 -508
rect 3538 -518 3624 -508
rect 4364 -535 5466 -508
rect 6298 -518 6384 -508
rect 6388 -535 6754 -508
rect 6758 -518 6844 -508
rect 6848 -535 7582 -508
rect 7586 -518 7672 -508
rect 7676 -535 8042 -508
rect 8046 -518 8132 -508
rect 8136 -535 8870 -508
rect 8874 -518 8960 -508
rect 8964 -535 9330 -508
rect 9334 -518 9420 -508
rect 9424 -535 10158 -508
rect 10162 -518 10248 -508
rect 10252 -535 10618 -508
rect 10622 -518 10708 -508
rect 10712 -535 11486 -508
rect 11542 -518 11628 -508
rect 11632 -535 11998 -508
rect 13474 -518 13560 -508
rect -2968 -573 -2934 -535
rect -2324 -577 -2290 -539
rect -2134 -568 -2112 -544
rect -1858 -568 -1836 -544
rect -1680 -568 -1648 -544
rect -1586 -566 -1554 -544
rect -1404 -573 -1370 -535
rect -945 -539 -911 -535
rect -945 -573 -910 -539
rect -576 -573 -542 -535
rect -944 -577 -910 -573
rect -208 -577 -174 -539
rect -116 -573 -82 -539
rect 252 -577 286 -539
rect 620 -573 654 -535
rect 1079 -573 1114 -539
rect 1448 -573 1482 -535
rect 1079 -577 1113 -573
rect 1540 -577 1574 -539
rect 1908 -573 1942 -535
rect 2369 -539 2403 -535
rect 2368 -573 2403 -539
rect 2368 -577 2402 -573
rect 2828 -577 2862 -539
rect 3196 -573 3230 -535
rect 3655 -546 3689 -539
rect 3653 -577 3697 -546
rect 4116 -577 4150 -539
rect 4392 -573 4426 -535
rect 4944 -577 4978 -539
rect 5404 -577 5438 -539
rect 5502 -568 5524 -544
rect 5863 -567 5887 -545
rect 5962 -568 5984 -544
rect 6231 -577 6265 -539
rect 6416 -573 6450 -535
rect 6692 -577 6726 -539
rect 6877 -573 6911 -535
rect 7520 -577 7554 -539
rect 7704 -573 7738 -535
rect 7980 -577 8014 -539
rect 8165 -573 8199 -535
rect 8807 -577 8841 -539
rect 8992 -573 9026 -535
rect 9268 -577 9302 -539
rect 9453 -573 9487 -535
rect 10096 -577 10130 -539
rect 10280 -545 10314 -535
rect 10648 -545 10682 -539
rect 10280 -567 10315 -545
rect 10648 -567 10683 -545
rect 10280 -573 10314 -567
rect 10648 -577 10682 -567
rect 10741 -573 10775 -535
rect 11383 -577 11417 -539
rect 11579 -567 11603 -545
rect 11660 -573 11694 -535
rect 11936 -577 11970 -539
rect -2996 -604 -2262 -577
rect -2258 -604 -2172 -594
rect -1616 -604 -882 -577
rect -880 -604 -146 -577
rect -142 -604 -56 -594
rect -52 -604 314 -577
rect 318 -604 404 -594
rect 408 -604 1142 -577
rect 1146 -604 1232 -594
rect 1236 -604 1602 -577
rect 1606 -604 1692 -594
rect 1696 -604 2430 -577
rect 2434 -604 2520 -594
rect 2524 -604 2890 -577
rect 2894 -604 2980 -594
rect 2984 -604 3718 -577
rect 3722 -604 3808 -594
rect 3812 -604 4178 -577
rect 4182 -604 4268 -594
rect 4272 -604 5006 -577
rect 5010 -604 5096 -594
rect 5100 -604 5466 -577
rect 5470 -604 5556 -594
rect 5560 -604 6294 -577
rect 6298 -604 6384 -594
rect 6388 -604 6754 -577
rect 6758 -604 6844 -594
rect 6848 -604 7582 -577
rect 7586 -604 7672 -594
rect 7676 -604 8042 -577
rect 8046 -604 8132 -594
rect 8136 -604 8870 -577
rect 8874 -604 8960 -594
rect 8964 -604 9330 -577
rect 9334 -604 9420 -594
rect 9424 -604 10158 -577
rect 10162 -604 10248 -594
rect 10344 -604 10710 -577
rect 10712 -604 11446 -577
rect 11450 -604 11536 -594
rect 11632 -604 11998 -577
rect 12025 -580 12069 -546
rect 12665 -566 12709 -532
rect 12761 -580 12805 -546
rect 13401 -566 13445 -532
rect 13564 -535 14666 -508
rect 14670 -518 14756 -508
rect 14760 -535 15862 -508
rect 15866 -518 15952 -508
rect 15956 -535 16690 -508
rect 13511 -567 13535 -545
rect 13592 -573 13626 -535
rect 13684 -577 13718 -539
rect 14788 -573 14822 -535
rect 15984 -573 16018 -535
rect 16628 -577 16662 -539
rect 13566 -604 13652 -594
rect 13656 -604 15477 -577
rect 15498 -604 15584 -594
rect 15588 -604 16690 -577
rect -3034 -752 16729 -604
rect 524 -759 1036 -752
rect 3100 -759 3612 -752
rect 5676 -759 6188 -752
rect 8252 -759 8764 -752
rect 10828 -759 11340 -752
rect 514 -1448 1026 -1441
rect 3090 -1448 3602 -1441
rect 5666 -1448 6178 -1441
rect 8242 -1448 8754 -1441
rect 10818 -1448 11330 -1441
rect -3035 -1596 16728 -1448
rect -2996 -1623 -2262 -1596
rect -2258 -1606 -2172 -1596
rect -1616 -1623 -882 -1596
rect -880 -1623 -146 -1596
rect -142 -1606 -56 -1596
rect -52 -1623 314 -1596
rect 318 -1606 404 -1596
rect 408 -1623 1142 -1596
rect 1146 -1606 1232 -1596
rect 1236 -1623 1602 -1596
rect 1606 -1606 1692 -1596
rect 1696 -1623 2430 -1596
rect 2434 -1606 2520 -1596
rect 2524 -1623 2890 -1596
rect 2894 -1606 2980 -1596
rect 2984 -1623 3718 -1596
rect 3722 -1606 3808 -1596
rect 3812 -1623 4178 -1596
rect 4182 -1606 4268 -1596
rect 4272 -1623 5006 -1596
rect 5010 -1606 5096 -1596
rect 5100 -1623 5466 -1596
rect 5470 -1606 5556 -1596
rect 5560 -1623 6294 -1596
rect 6298 -1606 6384 -1596
rect 6388 -1623 6754 -1596
rect 6758 -1606 6844 -1596
rect 6848 -1623 7582 -1596
rect 7586 -1606 7672 -1596
rect 7676 -1623 8042 -1596
rect 8046 -1606 8132 -1596
rect 8136 -1623 8870 -1596
rect 8874 -1606 8960 -1596
rect 8964 -1623 9330 -1596
rect 9334 -1606 9420 -1596
rect 9424 -1623 10158 -1596
rect 10162 -1606 10248 -1596
rect 10344 -1623 10710 -1596
rect 10712 -1623 11446 -1596
rect 11450 -1606 11536 -1596
rect 11632 -1623 11998 -1596
rect 12370 -1606 12456 -1596
rect 12541 -1623 13026 -1596
rect 13106 -1606 13192 -1596
rect 13196 -1623 13562 -1596
rect 13566 -1606 13652 -1596
rect 13656 -1623 15477 -1596
rect 15498 -1606 15584 -1596
rect 15588 -1623 16690 -1596
rect -2968 -1661 -2934 -1623
rect -2324 -1665 -2290 -1627
rect -2134 -1656 -2112 -1632
rect -1858 -1656 -1836 -1632
rect -1770 -1654 -1738 -1632
rect -1680 -1656 -1648 -1634
rect -1588 -1661 -1554 -1623
rect -944 -1665 -910 -1627
rect -852 -1661 -818 -1623
rect -209 -1665 -175 -1627
rect 252 -1665 286 -1623
rect 437 -1661 471 -1623
rect 1079 -1665 1113 -1627
rect 1540 -1665 1574 -1623
rect 1724 -1661 1758 -1623
rect 2368 -1665 2402 -1627
rect 2828 -1665 2862 -1623
rect 3013 -1661 3047 -1623
rect 3655 -1665 3689 -1627
rect 4116 -1665 4150 -1623
rect 4300 -1661 4334 -1623
rect 4944 -1665 4978 -1627
rect 5404 -1665 5438 -1623
rect 5589 -1661 5623 -1623
rect 6231 -1665 6265 -1627
rect 6692 -1665 6726 -1623
rect 6876 -1661 6910 -1623
rect 7520 -1665 7554 -1627
rect 7980 -1665 8014 -1623
rect 8165 -1661 8199 -1623
rect 8807 -1665 8841 -1627
rect 9268 -1665 9302 -1623
rect 9452 -1661 9486 -1623
rect 10096 -1665 10130 -1627
rect 10648 -1633 10682 -1623
rect 10291 -1655 10315 -1633
rect 10648 -1655 10683 -1633
rect 10648 -1665 10682 -1655
rect 10741 -1661 10775 -1623
rect 11383 -1665 11417 -1627
rect 11579 -1655 11603 -1633
rect 11936 -1665 11970 -1623
rect 12034 -1656 12056 -1632
rect 12488 -1661 12522 -1627
rect 12665 -1654 12709 -1623
rect 13224 -1661 13258 -1623
rect 13401 -1654 13445 -1623
rect 13511 -1655 13535 -1633
rect 13684 -1665 13718 -1623
rect 15616 -1661 15650 -1623
rect 16628 -1665 16662 -1627
rect -2996 -1692 -2262 -1665
rect -2258 -1692 -2172 -1682
rect -1616 -1692 -882 -1665
rect -880 -1692 -146 -1665
rect -142 -1692 -56 -1682
rect -52 -1692 314 -1665
rect 318 -1692 404 -1682
rect 408 -1692 1142 -1665
rect 1146 -1692 1232 -1682
rect 1236 -1692 1602 -1665
rect 1606 -1692 1692 -1682
rect 1696 -1692 2430 -1665
rect 2434 -1692 2520 -1682
rect 2524 -1692 2890 -1665
rect 2894 -1692 2980 -1682
rect 2984 -1692 3718 -1665
rect 3722 -1692 3808 -1682
rect 3812 -1692 4178 -1665
rect 4182 -1692 4268 -1682
rect 4272 -1692 5006 -1665
rect 5010 -1692 5096 -1682
rect 5100 -1692 5466 -1665
rect 5470 -1692 5556 -1682
rect 5560 -1692 6294 -1665
rect 6298 -1692 6384 -1682
rect 6388 -1692 6754 -1665
rect 6758 -1692 6844 -1682
rect 6848 -1692 7582 -1665
rect 7586 -1692 7672 -1682
rect 7676 -1692 8042 -1665
rect 8046 -1692 8132 -1682
rect 8136 -1692 8870 -1665
rect 8874 -1692 8960 -1682
rect 8964 -1692 9330 -1665
rect 9334 -1692 9420 -1682
rect 9424 -1692 10158 -1665
rect 10162 -1692 10248 -1682
rect 10344 -1692 10710 -1665
rect 10712 -1692 11446 -1665
rect 11450 -1692 11536 -1682
rect 11632 -1692 11998 -1665
rect 13566 -1692 13652 -1682
rect 13656 -1692 15477 -1665
rect 15498 -1692 15584 -1682
rect 15588 -1692 16690 -1665
rect -3034 -1840 16729 -1692
rect -764 -1847 -252 -1840
rect 524 -1847 1036 -1840
rect 3100 -1847 3612 -1840
rect 5676 -1847 6188 -1840
rect 8252 -1847 8764 -1840
rect 10828 -1847 11340 -1840
rect 514 -2536 1026 -2529
rect 3090 -2536 3602 -2529
rect 5666 -2536 6178 -2529
rect 8242 -2536 8754 -2529
rect 10818 -2536 11330 -2529
rect -3035 -2684 16728 -2536
rect -2996 -2711 -2262 -2684
rect -2258 -2694 -2172 -2684
rect -1616 -2711 -882 -2684
rect -880 -2711 -146 -2684
rect -142 -2694 -56 -2684
rect -52 -2711 314 -2684
rect 318 -2694 404 -2684
rect 408 -2711 1142 -2684
rect 1146 -2694 1232 -2684
rect 1236 -2711 1602 -2684
rect 1606 -2694 1692 -2684
rect 1696 -2711 2430 -2684
rect 2434 -2694 2520 -2684
rect 2524 -2711 2890 -2684
rect 2894 -2694 2980 -2684
rect 2984 -2711 3718 -2684
rect 3722 -2694 3808 -2684
rect 3812 -2711 4178 -2684
rect 4182 -2694 4268 -2684
rect 4272 -2711 5006 -2684
rect 5010 -2694 5096 -2684
rect 5100 -2711 5466 -2684
rect 5470 -2694 5556 -2684
rect 5560 -2711 6294 -2684
rect 6298 -2694 6384 -2684
rect 6388 -2711 6754 -2684
rect 6758 -2694 6844 -2684
rect 6848 -2711 7582 -2684
rect 7586 -2694 7672 -2684
rect 7676 -2711 8042 -2684
rect 8046 -2694 8132 -2684
rect 8136 -2711 8870 -2684
rect 8874 -2694 8960 -2684
rect 8964 -2711 9330 -2684
rect 9334 -2694 9420 -2684
rect 9424 -2711 10158 -2684
rect 10162 -2694 10248 -2684
rect 10344 -2711 10710 -2684
rect 10712 -2711 11446 -2684
rect 11450 -2694 11536 -2684
rect 11632 -2711 11998 -2684
rect 12370 -2694 12456 -2684
rect 12541 -2711 13026 -2684
rect 13106 -2694 13192 -2684
rect 13196 -2711 13562 -2684
rect 13566 -2694 13652 -2684
rect 13656 -2711 15477 -2684
rect 15498 -2694 15584 -2684
rect 15588 -2711 16690 -2684
rect -2968 -2749 -2934 -2711
rect -2324 -2753 -2290 -2715
rect -2134 -2744 -2112 -2720
rect -2048 -2744 -2016 -2722
rect -1956 -2749 -1922 -2715
rect -1770 -2742 -1738 -2720
rect -1588 -2749 -1554 -2711
rect -944 -2753 -910 -2715
rect -852 -2749 -818 -2711
rect -208 -2753 -174 -2715
rect 252 -2753 286 -2711
rect 437 -2749 471 -2711
rect 1079 -2753 1113 -2715
rect 1540 -2753 1574 -2711
rect 1724 -2749 1758 -2711
rect 2368 -2753 2402 -2715
rect 2828 -2753 2862 -2711
rect 3013 -2749 3047 -2711
rect 3655 -2753 3689 -2715
rect 4116 -2753 4150 -2711
rect 4300 -2749 4334 -2711
rect 4944 -2753 4978 -2715
rect 5404 -2753 5438 -2711
rect 5589 -2749 5623 -2711
rect 6231 -2753 6265 -2715
rect 6692 -2753 6726 -2711
rect 6876 -2749 6910 -2711
rect 7520 -2753 7554 -2715
rect 7980 -2753 8014 -2711
rect 8165 -2749 8199 -2711
rect 8807 -2753 8841 -2715
rect 9268 -2753 9302 -2711
rect 9452 -2749 9486 -2711
rect 10096 -2753 10130 -2715
rect 10648 -2721 10682 -2711
rect 10291 -2743 10315 -2721
rect 10648 -2743 10683 -2721
rect 10648 -2753 10682 -2743
rect 10741 -2749 10775 -2711
rect 11383 -2753 11417 -2715
rect 11579 -2743 11603 -2721
rect 11936 -2753 11970 -2711
rect 12034 -2744 12056 -2720
rect 12488 -2749 12522 -2715
rect 12665 -2742 12709 -2711
rect 13224 -2749 13258 -2711
rect 13401 -2742 13445 -2711
rect 13684 -2749 13718 -2711
rect 14604 -2753 14638 -2715
rect 15616 -2749 15650 -2711
rect 15800 -2753 15834 -2715
rect 16628 -2753 16662 -2715
rect -2996 -2780 -2262 -2753
rect -2258 -2780 -2172 -2770
rect -1901 -2780 -1710 -2753
rect -1706 -2780 -1620 -2770
rect -1616 -2780 -882 -2753
rect -880 -2780 -146 -2753
rect -142 -2780 -56 -2770
rect -52 -2780 314 -2753
rect 318 -2780 404 -2770
rect 408 -2780 1142 -2753
rect 1146 -2780 1232 -2770
rect 1236 -2780 1602 -2753
rect 1606 -2780 1692 -2770
rect 1696 -2780 2430 -2753
rect 2434 -2780 2520 -2770
rect 2524 -2780 2890 -2753
rect 2894 -2780 2980 -2770
rect 2984 -2780 3718 -2753
rect 3722 -2780 3808 -2770
rect 3812 -2780 4178 -2753
rect 4182 -2780 4268 -2770
rect 4272 -2780 5006 -2753
rect 5010 -2780 5096 -2770
rect 5100 -2780 5466 -2753
rect 5470 -2780 5556 -2770
rect 5560 -2780 6294 -2753
rect 6298 -2780 6384 -2770
rect 6388 -2780 6754 -2753
rect 6758 -2780 6844 -2770
rect 6848 -2780 7582 -2753
rect 7586 -2780 7672 -2770
rect 7676 -2780 8042 -2753
rect 8046 -2780 8132 -2770
rect 8136 -2780 8870 -2753
rect 8874 -2780 8960 -2770
rect 8964 -2780 9330 -2753
rect 9334 -2780 9420 -2770
rect 9424 -2780 10158 -2753
rect 10162 -2780 10248 -2770
rect 10344 -2780 10710 -2753
rect 10712 -2780 11446 -2753
rect 11450 -2780 11536 -2770
rect 11632 -2780 11998 -2753
rect 13474 -2780 13560 -2770
rect 13564 -2780 14666 -2753
rect 14670 -2780 14756 -2770
rect 14760 -2780 15862 -2753
rect 15866 -2780 15952 -2770
rect 15956 -2780 16690 -2753
rect -3034 -2928 16729 -2780
rect 524 -2935 1036 -2928
rect 3100 -2935 3612 -2928
rect 5676 -2935 6188 -2928
rect 8252 -2935 8764 -2928
rect 10828 -2935 11340 -2928
rect 524 -3624 1036 -3617
rect 3100 -3624 3612 -3617
rect 5676 -3624 6188 -3617
rect 8252 -3624 8764 -3617
rect 10828 -3624 11340 -3617
rect -3035 -3772 16728 -3624
rect -2996 -3799 -2262 -3772
rect -2258 -3782 -2172 -3772
rect -1616 -3799 -882 -3772
rect -880 -3799 -146 -3772
rect -142 -3782 -56 -3772
rect -52 -3799 314 -3772
rect 318 -3782 404 -3772
rect 408 -3799 1142 -3772
rect 1146 -3782 1232 -3772
rect 1236 -3799 1602 -3772
rect 1606 -3782 1692 -3772
rect 1696 -3799 2430 -3772
rect 2434 -3782 2520 -3772
rect 2524 -3799 2890 -3772
rect 2894 -3782 2980 -3772
rect 2984 -3799 3718 -3772
rect 3722 -3782 3808 -3772
rect 3812 -3799 4178 -3772
rect 4182 -3782 4268 -3772
rect 4272 -3799 5006 -3772
rect 5010 -3782 5096 -3772
rect 5100 -3799 5466 -3772
rect 5470 -3782 5556 -3772
rect 5560 -3799 6294 -3772
rect 6298 -3782 6384 -3772
rect 6388 -3799 6754 -3772
rect 6758 -3782 6844 -3772
rect 6848 -3799 7582 -3772
rect 7586 -3782 7672 -3772
rect 7676 -3799 8042 -3772
rect 8046 -3782 8132 -3772
rect 8136 -3799 8870 -3772
rect 8874 -3782 8960 -3772
rect 8964 -3799 9330 -3772
rect 9334 -3782 9420 -3772
rect 9424 -3799 10158 -3772
rect 10162 -3782 10248 -3772
rect 10344 -3799 10710 -3772
rect 10712 -3799 11446 -3772
rect 11450 -3782 11536 -3772
rect 11632 -3799 11998 -3772
rect 13474 -3782 13560 -3772
rect 13564 -3799 14666 -3772
rect 14670 -3782 14756 -3772
rect 14760 -3799 15862 -3772
rect 15866 -3782 15952 -3772
rect 15956 -3799 16690 -3772
rect -2968 -3837 -2934 -3799
rect -2324 -3841 -2290 -3803
rect -2134 -3832 -2112 -3808
rect -1858 -3832 -1836 -3808
rect -1770 -3830 -1738 -3808
rect -1680 -3832 -1648 -3810
rect -1588 -3841 -1554 -3803
rect -944 -3837 -910 -3799
rect -852 -3841 -818 -3803
rect -208 -3837 -174 -3799
rect 252 -3841 286 -3799
rect 437 -3841 471 -3803
rect 1079 -3837 1113 -3799
rect 1540 -3841 1574 -3799
rect 1724 -3837 1758 -3799
rect 2368 -3841 2402 -3803
rect 2828 -3841 2862 -3799
rect 3013 -3841 3047 -3803
rect 3655 -3837 3689 -3799
rect 4116 -3841 4150 -3799
rect 4300 -3837 4334 -3799
rect 4944 -3841 4978 -3803
rect 5404 -3841 5438 -3799
rect 5589 -3841 5623 -3803
rect 6231 -3837 6265 -3799
rect 6692 -3841 6726 -3799
rect 6876 -3837 6910 -3799
rect 7520 -3841 7554 -3803
rect 7980 -3841 8014 -3799
rect 8165 -3841 8199 -3803
rect 8807 -3837 8841 -3799
rect 9268 -3841 9302 -3799
rect 9452 -3837 9486 -3799
rect 10096 -3841 10130 -3803
rect 10648 -3809 10682 -3799
rect 10291 -3831 10315 -3809
rect 10648 -3831 10683 -3809
rect 10648 -3841 10682 -3831
rect 10741 -3841 10775 -3803
rect 11383 -3837 11417 -3799
rect 11579 -3831 11603 -3809
rect 11936 -3841 11970 -3799
rect 12034 -3832 12056 -3808
rect 12488 -3837 12522 -3803
rect 12665 -3841 12709 -3810
rect 13224 -3841 13258 -3803
rect 13401 -3841 13445 -3810
rect 13684 -3841 13718 -3803
rect 14604 -3837 14638 -3799
rect 15616 -3841 15650 -3803
rect 15800 -3837 15834 -3799
rect 16628 -3837 16662 -3799
rect -2996 -3868 -2262 -3841
rect -2258 -3868 -2172 -3858
rect -1616 -3868 -882 -3841
rect -880 -3868 -146 -3841
rect -142 -3868 -56 -3858
rect -52 -3868 314 -3841
rect 318 -3868 404 -3858
rect 408 -3868 1142 -3841
rect 1146 -3868 1232 -3858
rect 1236 -3868 1602 -3841
rect 1606 -3868 1692 -3858
rect 1696 -3868 2430 -3841
rect 2434 -3868 2520 -3858
rect 2524 -3868 2890 -3841
rect 2894 -3868 2980 -3858
rect 2984 -3868 3718 -3841
rect 3722 -3868 3808 -3858
rect 3812 -3868 4178 -3841
rect 4182 -3868 4268 -3858
rect 4272 -3868 5006 -3841
rect 5010 -3868 5096 -3858
rect 5100 -3868 5466 -3841
rect 5470 -3868 5556 -3858
rect 5560 -3868 6294 -3841
rect 6298 -3868 6384 -3858
rect 6388 -3868 6754 -3841
rect 6758 -3868 6844 -3858
rect 6848 -3868 7582 -3841
rect 7586 -3868 7672 -3858
rect 7676 -3868 8042 -3841
rect 8046 -3868 8132 -3858
rect 8136 -3868 8870 -3841
rect 8874 -3868 8960 -3858
rect 8964 -3868 9330 -3841
rect 9334 -3868 9420 -3858
rect 9424 -3868 10158 -3841
rect 10162 -3868 10248 -3858
rect 10344 -3868 10710 -3841
rect 10712 -3868 11446 -3841
rect 11450 -3868 11536 -3858
rect 11632 -3868 11998 -3841
rect 12370 -3868 12456 -3858
rect 12541 -3868 13026 -3841
rect 13106 -3868 13192 -3858
rect 13196 -3868 13562 -3841
rect 13566 -3868 13652 -3858
rect 13656 -3868 15477 -3841
rect 15498 -3868 15584 -3858
rect 15588 -3868 16690 -3841
rect -3034 -4016 16729 -3868
rect 514 -4023 1026 -4016
rect 3090 -4023 3602 -4016
rect 5666 -4023 6178 -4016
rect 8242 -4023 8754 -4016
rect 10818 -4023 11330 -4016
rect -764 -4712 -252 -4705
rect 524 -4712 1036 -4705
rect 3100 -4712 3612 -4705
rect 5676 -4712 6188 -4705
rect 8252 -4712 8764 -4705
rect 10828 -4712 11340 -4705
rect -3035 -4860 16728 -4712
rect -2996 -4887 -2262 -4860
rect -2258 -4870 -2172 -4860
rect -1616 -4887 -882 -4860
rect -880 -4887 -146 -4860
rect -142 -4870 -56 -4860
rect -52 -4887 314 -4860
rect 318 -4870 404 -4860
rect 408 -4887 1142 -4860
rect 1146 -4870 1232 -4860
rect 1236 -4887 1602 -4860
rect 1606 -4870 1692 -4860
rect 1696 -4887 2430 -4860
rect 2434 -4870 2520 -4860
rect 2524 -4887 2890 -4860
rect 2894 -4870 2980 -4860
rect 2984 -4887 3718 -4860
rect 3722 -4870 3808 -4860
rect 3812 -4887 4178 -4860
rect 4182 -4870 4268 -4860
rect 4272 -4887 5006 -4860
rect 5010 -4870 5096 -4860
rect 5100 -4887 5466 -4860
rect 5470 -4870 5556 -4860
rect 5560 -4887 6294 -4860
rect 6298 -4870 6384 -4860
rect 6388 -4887 6754 -4860
rect 6758 -4870 6844 -4860
rect 6848 -4887 7582 -4860
rect 7586 -4870 7672 -4860
rect 7676 -4887 8042 -4860
rect 8046 -4870 8132 -4860
rect 8136 -4887 8870 -4860
rect 8874 -4870 8960 -4860
rect 8964 -4887 9330 -4860
rect 9334 -4870 9420 -4860
rect 9424 -4887 10158 -4860
rect 10162 -4870 10248 -4860
rect 10344 -4887 10710 -4860
rect 10712 -4887 11446 -4860
rect 11450 -4870 11536 -4860
rect 11632 -4887 11998 -4860
rect 13566 -4870 13652 -4860
rect 13656 -4887 15477 -4860
rect 15498 -4870 15584 -4860
rect 15588 -4887 16690 -4860
rect -2968 -4925 -2934 -4887
rect -2324 -4929 -2290 -4891
rect -2134 -4920 -2112 -4896
rect -1858 -4920 -1836 -4896
rect -1770 -4918 -1738 -4896
rect -1680 -4920 -1648 -4898
rect -1588 -4929 -1554 -4891
rect -944 -4925 -910 -4887
rect -852 -4929 -818 -4891
rect -209 -4925 -175 -4887
rect 252 -4929 286 -4887
rect 437 -4929 471 -4891
rect 1079 -4925 1113 -4887
rect 1540 -4929 1574 -4887
rect 1724 -4925 1758 -4887
rect 2368 -4929 2402 -4891
rect 2828 -4929 2862 -4887
rect 3013 -4929 3047 -4891
rect 3655 -4925 3689 -4887
rect 4116 -4929 4150 -4887
rect 4300 -4925 4334 -4887
rect 4944 -4929 4978 -4891
rect 5404 -4929 5438 -4887
rect 5589 -4929 5623 -4891
rect 6231 -4925 6265 -4887
rect 6692 -4929 6726 -4887
rect 6876 -4925 6910 -4887
rect 7520 -4929 7554 -4891
rect 7980 -4929 8014 -4887
rect 8165 -4929 8199 -4891
rect 8807 -4925 8841 -4887
rect 9268 -4929 9302 -4887
rect 9452 -4925 9486 -4887
rect 10096 -4929 10130 -4891
rect 10648 -4897 10682 -4887
rect 10291 -4919 10315 -4897
rect 10648 -4919 10683 -4897
rect 10648 -4929 10682 -4919
rect 10741 -4929 10775 -4891
rect 11383 -4925 11417 -4887
rect 11579 -4919 11603 -4897
rect 11936 -4929 11970 -4887
rect 12034 -4920 12056 -4896
rect 12488 -4925 12522 -4891
rect 12665 -4929 12709 -4898
rect 13224 -4929 13258 -4891
rect 13401 -4929 13445 -4898
rect 13511 -4919 13535 -4897
rect 13684 -4929 13718 -4887
rect 15616 -4929 15650 -4891
rect 16628 -4925 16662 -4887
rect -2996 -4956 -2262 -4929
rect -2258 -4956 -2172 -4946
rect -1616 -4956 -882 -4929
rect -880 -4956 -146 -4929
rect -142 -4956 -56 -4946
rect -52 -4956 314 -4929
rect 318 -4956 404 -4946
rect 408 -4956 1142 -4929
rect 1146 -4956 1232 -4946
rect 1236 -4956 1602 -4929
rect 1606 -4956 1692 -4946
rect 1696 -4956 2430 -4929
rect 2434 -4956 2520 -4946
rect 2524 -4956 2890 -4929
rect 2894 -4956 2980 -4946
rect 2984 -4956 3718 -4929
rect 3722 -4956 3808 -4946
rect 3812 -4956 4178 -4929
rect 4182 -4956 4268 -4946
rect 4272 -4956 5006 -4929
rect 5010 -4956 5096 -4946
rect 5100 -4956 5466 -4929
rect 5470 -4956 5556 -4946
rect 5560 -4956 6294 -4929
rect 6298 -4956 6384 -4946
rect 6388 -4956 6754 -4929
rect 6758 -4956 6844 -4946
rect 6848 -4956 7582 -4929
rect 7586 -4956 7672 -4946
rect 7676 -4956 8042 -4929
rect 8046 -4956 8132 -4946
rect 8136 -4956 8870 -4929
rect 8874 -4956 8960 -4946
rect 8964 -4956 9330 -4929
rect 9334 -4956 9420 -4946
rect 9424 -4956 10158 -4929
rect 10162 -4956 10248 -4946
rect 10344 -4956 10710 -4929
rect 10712 -4956 11446 -4929
rect 11450 -4956 11536 -4946
rect 11632 -4956 11998 -4929
rect 12370 -4956 12456 -4946
rect 12541 -4956 13026 -4929
rect 13106 -4956 13192 -4946
rect 13196 -4956 13562 -4929
rect 13566 -4956 13652 -4946
rect 13656 -4956 15477 -4929
rect 15498 -4956 15584 -4946
rect 15588 -4956 16690 -4929
rect -3034 -5104 16729 -4956
rect 514 -5111 1026 -5104
rect 3090 -5111 3602 -5104
rect 5666 -5111 6178 -5104
rect 8242 -5111 8754 -5104
rect 10818 -5111 11330 -5104
rect -948 -5793 -896 -5780
rect 524 -5800 1036 -5793
rect 3100 -5800 3612 -5793
rect 5676 -5800 6188 -5793
rect 8252 -5800 8764 -5793
rect 10828 -5800 11340 -5793
rect -3035 -5948 16728 -5800
rect -2996 -5975 -2262 -5948
rect -2258 -5958 -2172 -5948
rect -1616 -5975 -882 -5948
rect -880 -5975 -146 -5948
rect -142 -5958 -56 -5948
rect -52 -5975 314 -5948
rect 318 -5958 404 -5948
rect 408 -5975 1142 -5948
rect 1146 -5958 1232 -5948
rect 1236 -5975 1602 -5948
rect 1606 -5958 1692 -5948
rect 1696 -5975 2430 -5948
rect 2434 -5958 2520 -5948
rect 2524 -5975 2890 -5948
rect 2894 -5958 2980 -5948
rect 2984 -5975 3718 -5948
rect 3722 -5958 3808 -5948
rect 3812 -5975 4178 -5948
rect 4182 -5958 4268 -5948
rect 4272 -5975 5006 -5948
rect 5010 -5958 5096 -5948
rect 5100 -5975 5466 -5948
rect 5470 -5958 5556 -5948
rect 5560 -5975 6294 -5948
rect 6298 -5958 6384 -5948
rect 6388 -5975 6754 -5948
rect 6758 -5958 6844 -5948
rect 6848 -5975 7582 -5948
rect 7586 -5958 7672 -5948
rect 7676 -5975 8042 -5948
rect 8046 -5958 8132 -5948
rect 8136 -5975 8870 -5948
rect 8874 -5958 8960 -5948
rect 8964 -5975 9330 -5948
rect 9334 -5958 9420 -5948
rect 9424 -5975 10158 -5948
rect 10162 -5958 10248 -5948
rect 10344 -5975 10710 -5948
rect 10712 -5975 11446 -5948
rect 11450 -5958 11536 -5948
rect 11632 -5975 11998 -5948
rect 13566 -5958 13652 -5948
rect -2968 -6013 -2934 -5975
rect -944 -5979 -910 -5975
rect -2324 -6017 -2290 -5979
rect -2134 -6008 -2112 -5984
rect -1858 -6008 -1836 -5984
rect -1770 -6006 -1738 -5984
rect -1680 -6008 -1648 -5986
rect -1586 -6008 -1554 -5986
rect -1404 -6017 -1370 -5979
rect -945 -6013 -910 -5979
rect -945 -6017 -911 -6013
rect -576 -6017 -542 -5979
rect -208 -6013 -174 -5975
rect -116 -6013 -82 -5979
rect 252 -6013 286 -5975
rect 1079 -5979 1113 -5975
rect 620 -6017 654 -5979
rect 1079 -6013 1114 -5979
rect 1448 -6017 1482 -5979
rect 1540 -6013 1574 -5975
rect 1724 -6013 1758 -5975
rect 1908 -6017 1942 -5979
rect 2369 -6017 2403 -5979
rect 2828 -6013 2862 -5975
rect 3196 -6017 3230 -5979
rect 3653 -6006 3697 -5975
rect 3655 -6013 3689 -6006
rect 4116 -6013 4150 -5975
rect 4300 -6013 4334 -5975
rect 4392 -6017 4426 -5979
rect 5404 -6013 5438 -5975
rect 5502 -6008 5524 -5984
rect 5863 -6007 5887 -5985
rect 5962 -6008 5984 -5984
rect 6231 -6013 6265 -5975
rect 6416 -6017 6450 -5979
rect 6692 -6013 6726 -5975
rect 6876 -5979 6910 -5975
rect 6876 -6013 6911 -5979
rect 6877 -6017 6911 -6013
rect 7704 -6017 7738 -5979
rect 7980 -6013 8014 -5975
rect 8165 -6017 8199 -5979
rect 8807 -6013 8841 -5975
rect 8992 -6017 9026 -5979
rect 9268 -6013 9302 -5975
rect 9452 -5979 9486 -5975
rect 9452 -6013 9487 -5979
rect 9453 -6017 9487 -6013
rect 10280 -5985 10314 -5979
rect 10648 -5985 10682 -5975
rect 10280 -6007 10315 -5985
rect 10648 -6007 10683 -5985
rect 10280 -6017 10314 -6007
rect 10648 -6013 10682 -6007
rect 10741 -6017 10775 -5979
rect 11383 -6013 11417 -5975
rect 11579 -6007 11603 -5985
rect 11660 -6017 11694 -5979
rect 11936 -6013 11970 -5975
rect 12025 -6006 12069 -5972
rect -2996 -6044 -2262 -6017
rect -2258 -6044 -2172 -6034
rect -1432 -6044 -1066 -6017
rect -1062 -6044 -976 -6034
rect -968 -6044 -698 -6017
rect -694 -6044 -608 -6034
rect -604 -6044 -238 -6017
rect -234 -6044 -148 -6034
rect -63 -6044 422 -6017
rect 502 -6044 588 -6034
rect 592 -6044 958 -6017
rect 962 -6044 1048 -6034
rect 1135 -6044 1326 -6017
rect 1330 -6044 1416 -6034
rect 1420 -6044 1786 -6017
rect 1790 -6044 1876 -6034
rect 1880 -6044 2246 -6017
rect 2250 -6044 2336 -6034
rect 2340 -6044 3074 -6017
rect 3078 -6044 3164 -6034
rect 3168 -6044 3534 -6017
rect 3538 -6044 3624 -6034
rect 4364 -6044 5466 -6017
rect 6298 -6044 6384 -6034
rect 6388 -6044 6754 -6017
rect 6758 -6044 6844 -6034
rect 6848 -6044 7582 -6017
rect 7586 -6044 7672 -6034
rect 7676 -6044 8042 -6017
rect 8046 -6044 8132 -6034
rect 8136 -6044 8870 -6017
rect 8874 -6044 8960 -6034
rect 8964 -6044 9330 -6017
rect 9334 -6044 9420 -6034
rect 9424 -6044 10158 -6017
rect 10162 -6044 10248 -6034
rect 10252 -6044 10618 -6017
rect 10622 -6044 10708 -6034
rect 10712 -6044 11486 -6017
rect 11542 -6044 11628 -6034
rect 11632 -6044 11998 -6017
rect 12665 -6020 12709 -5986
rect 12761 -6006 12805 -5972
rect 13656 -5975 15477 -5948
rect 15498 -5958 15584 -5948
rect 15588 -5975 16690 -5948
rect 13401 -6020 13445 -5986
rect 13511 -6007 13535 -5985
rect 13592 -6017 13626 -5979
rect 13684 -6013 13718 -5975
rect 14788 -6017 14822 -5979
rect 15984 -6017 16018 -5979
rect 16628 -6013 16662 -5975
rect 13474 -6044 13560 -6034
rect 13564 -6044 14666 -6017
rect 14670 -6044 14756 -6034
rect 14760 -6044 15862 -6017
rect 15866 -6044 15952 -6034
rect 15956 -6044 16690 -6017
rect -3034 -6192 16729 -6044
rect -968 -6199 -698 -6192
rect 2446 -6199 2958 -6192
rect 6954 -6199 7466 -6192
rect 8242 -6199 8754 -6192
rect 9530 -6199 10042 -6192
rect 10712 -6199 11486 -6192
rect -1925 -6888 -1743 -6883
rect -1435 -6888 -882 -6881
rect -3035 -7036 16728 -6888
rect -2996 -7063 -2722 -7036
rect -2718 -7046 -2632 -7036
rect -2628 -7063 -882 -7036
rect -880 -7063 -146 -7036
rect -142 -7046 -56 -7036
rect -52 -7063 682 -7036
rect 684 -7063 1418 -7036
rect 1422 -7046 1508 -7036
rect 1512 -7063 2246 -7036
rect 2248 -7063 2982 -7036
rect 2986 -7046 3072 -7036
rect 3076 -7063 3810 -7036
rect 3812 -7063 4546 -7036
rect 4550 -7046 4636 -7036
rect 4640 -7063 5374 -7036
rect 5376 -7063 6110 -7036
rect 6114 -7046 6200 -7036
rect 6204 -7063 6938 -7036
rect 6940 -7063 7674 -7036
rect 7678 -7046 7764 -7036
rect 7768 -7063 8502 -7036
rect 8504 -7063 9238 -7036
rect 9242 -7046 9328 -7036
rect 15866 -7046 15952 -7036
rect -2968 -7101 -2934 -7063
rect -2600 -7101 -2566 -7063
rect -2324 -7105 -2290 -7067
rect -1858 -7096 -1836 -7072
rect -1680 -7096 -1648 -7074
rect -1588 -7105 -1554 -7067
rect -852 -7105 -818 -7067
rect -208 -7101 -174 -7063
rect -24 -7105 10 -7067
rect 620 -7101 654 -7063
rect 712 -7105 746 -7067
rect 1356 -7101 1390 -7063
rect 1540 -7105 1574 -7067
rect 2184 -7101 2218 -7063
rect 2552 -7105 2586 -7067
rect 2736 -7096 2768 -7074
rect 2920 -7101 2954 -7063
rect 3748 -7067 3782 -7063
rect 3104 -7101 3138 -7067
rect 3564 -7105 3598 -7067
rect 3747 -7101 3782 -7067
rect 3747 -7105 3781 -7101
rect 4392 -7105 4426 -7067
rect 4484 -7101 4518 -7063
rect 4631 -7105 4665 -7067
rect 5312 -7101 5346 -7063
rect 5772 -7105 5806 -7067
rect 6048 -7101 6082 -7063
rect 6876 -7101 6910 -7063
rect 7612 -7105 7646 -7063
rect 7796 -7105 7830 -7067
rect 8440 -7101 8474 -7063
rect 8532 -7105 8566 -7067
rect 9176 -7101 9210 -7063
rect -2996 -7132 -2262 -7105
rect -2258 -7132 -2172 -7122
rect -1616 -7132 -882 -7105
rect -880 -7132 -146 -7105
rect -142 -7132 -56 -7122
rect -52 -7132 682 -7105
rect 684 -7132 1418 -7105
rect 1422 -7132 1508 -7122
rect 1512 -7132 2246 -7105
rect 2248 -7132 2614 -7105
rect 2802 -7132 2888 -7122
rect 2892 -7132 3083 -7105
rect 3170 -7132 3256 -7122
rect 3260 -7132 3626 -7105
rect 3630 -7132 3716 -7122
rect 3724 -7132 3994 -7105
rect 3998 -7132 4084 -7122
rect 4088 -7132 4454 -7105
rect 4458 -7132 4544 -7122
rect 4548 -7132 5328 -7105
rect 5378 -7132 5464 -7122
rect 5468 -7132 5834 -7105
rect 5838 -7132 5924 -7122
rect 5928 -7132 7674 -7105
rect 7678 -7132 7764 -7122
rect 7768 -7132 8502 -7105
rect 8504 -7132 9238 -7105
rect 9357 -7108 9401 -7074
rect 9997 -7094 10041 -7060
rect 10093 -7108 10137 -7074
rect 10733 -7094 10777 -7060
rect 10829 -7108 10873 -7074
rect 11469 -7094 11513 -7060
rect 11565 -7108 11609 -7074
rect 12205 -7094 12249 -7060
rect 12301 -7108 12345 -7074
rect 12941 -7094 12985 -7060
rect 13037 -7108 13081 -7074
rect 13677 -7094 13721 -7060
rect 13773 -7108 13817 -7074
rect 14413 -7094 14457 -7060
rect 14509 -7108 14553 -7074
rect 15149 -7094 15193 -7060
rect 15245 -7108 15289 -7074
rect 15885 -7094 15929 -7060
rect 15956 -7063 16690 -7036
rect 15984 -7105 16018 -7067
rect 16628 -7101 16662 -7063
rect 9242 -7132 9328 -7122
rect 15866 -7132 15952 -7122
rect 15956 -7132 16690 -7105
rect -3034 -7280 16729 -7132
rect 3724 -7287 3994 -7280
rect 4548 -7287 4734 -7280
rect 5928 -7287 6481 -7280
rect 6789 -7285 6971 -7280
rect -968 -7976 -698 -7969
rect 2446 -7976 2958 -7969
rect 6954 -7976 7466 -7969
rect 8242 -7976 8754 -7969
rect 9530 -7976 10042 -7969
rect 10712 -7976 11486 -7969
rect -3035 -8124 16728 -7976
rect -2996 -8151 -2262 -8124
rect -2258 -8134 -2172 -8124
rect -1432 -8151 -1066 -8124
rect -1062 -8134 -976 -8124
rect -968 -8151 -698 -8124
rect -694 -8134 -608 -8124
rect -604 -8151 -238 -8124
rect -234 -8134 -148 -8124
rect -63 -8151 422 -8124
rect 502 -8134 588 -8124
rect 592 -8151 958 -8124
rect 962 -8134 1048 -8124
rect 1135 -8151 1326 -8124
rect 1330 -8134 1416 -8124
rect 1420 -8151 1786 -8124
rect 1790 -8134 1876 -8124
rect 1880 -8151 2246 -8124
rect 2250 -8134 2336 -8124
rect 2340 -8151 3074 -8124
rect 3078 -8134 3164 -8124
rect 3168 -8151 3534 -8124
rect 3538 -8134 3624 -8124
rect 4364 -8151 5466 -8124
rect 6298 -8134 6384 -8124
rect 6388 -8151 6754 -8124
rect 6758 -8134 6844 -8124
rect 6848 -8151 7582 -8124
rect 7586 -8134 7672 -8124
rect 7676 -8151 8042 -8124
rect 8046 -8134 8132 -8124
rect 8136 -8151 8870 -8124
rect 8874 -8134 8960 -8124
rect 8964 -8151 9330 -8124
rect 9334 -8134 9420 -8124
rect 9424 -8151 10158 -8124
rect 10162 -8134 10248 -8124
rect 10252 -8151 10618 -8124
rect 10622 -8134 10708 -8124
rect 10712 -8151 11486 -8124
rect 11542 -8134 11628 -8124
rect 11632 -8151 11998 -8124
rect 13474 -8134 13560 -8124
rect -2968 -8189 -2934 -8151
rect -2324 -8193 -2290 -8155
rect -2134 -8184 -2112 -8160
rect -1858 -8184 -1836 -8160
rect -1770 -8182 -1738 -8160
rect -1680 -8184 -1648 -8162
rect -1586 -8182 -1554 -8160
rect -1404 -8189 -1370 -8151
rect -945 -8155 -911 -8151
rect -945 -8189 -910 -8155
rect -576 -8189 -542 -8151
rect -944 -8193 -910 -8189
rect -208 -8193 -174 -8155
rect -116 -8189 -82 -8155
rect 252 -8193 286 -8155
rect 620 -8189 654 -8151
rect 1079 -8189 1114 -8155
rect 1448 -8189 1482 -8151
rect 1079 -8193 1113 -8189
rect 1540 -8193 1574 -8155
rect 1908 -8189 1942 -8151
rect 2369 -8155 2403 -8151
rect 2368 -8189 2403 -8155
rect 2368 -8193 2402 -8189
rect 2828 -8193 2862 -8155
rect 3196 -8189 3230 -8151
rect 3655 -8162 3689 -8155
rect 3653 -8193 3697 -8162
rect 4116 -8193 4150 -8155
rect 4392 -8189 4426 -8151
rect 4944 -8193 4978 -8155
rect 5404 -8193 5438 -8155
rect 5502 -8184 5524 -8160
rect 5863 -8183 5887 -8161
rect 5962 -8184 5984 -8160
rect 6231 -8193 6265 -8155
rect 6416 -8189 6450 -8151
rect 6692 -8193 6726 -8155
rect 6877 -8189 6911 -8151
rect 7520 -8193 7554 -8155
rect 7704 -8189 7738 -8151
rect 7980 -8193 8014 -8155
rect 8165 -8189 8199 -8151
rect 8807 -8193 8841 -8155
rect 8992 -8189 9026 -8151
rect 9268 -8193 9302 -8155
rect 9453 -8189 9487 -8151
rect 10096 -8193 10130 -8155
rect 10280 -8161 10314 -8151
rect 10648 -8161 10682 -8155
rect 10280 -8183 10315 -8161
rect 10648 -8183 10683 -8161
rect 10280 -8189 10314 -8183
rect 10648 -8193 10682 -8183
rect 10741 -8189 10775 -8151
rect 11383 -8193 11417 -8155
rect 11579 -8183 11603 -8161
rect 11660 -8189 11694 -8151
rect 11936 -8193 11970 -8155
rect -2996 -8220 -2262 -8193
rect -2258 -8220 -2172 -8210
rect -1616 -8220 -882 -8193
rect -880 -8220 -146 -8193
rect -142 -8220 -56 -8210
rect -52 -8220 314 -8193
rect 318 -8220 404 -8210
rect 408 -8220 1142 -8193
rect 1146 -8220 1232 -8210
rect 1236 -8220 1602 -8193
rect 1606 -8220 1692 -8210
rect 1696 -8220 2430 -8193
rect 2434 -8220 2520 -8210
rect 2524 -8220 2890 -8193
rect 2894 -8220 2980 -8210
rect 2984 -8220 3718 -8193
rect 3722 -8220 3808 -8210
rect 3812 -8220 4178 -8193
rect 4182 -8220 4268 -8210
rect 4272 -8220 5006 -8193
rect 5010 -8220 5096 -8210
rect 5100 -8220 5466 -8193
rect 5470 -8220 5556 -8210
rect 5560 -8220 6294 -8193
rect 6298 -8220 6384 -8210
rect 6388 -8220 6754 -8193
rect 6758 -8220 6844 -8210
rect 6848 -8220 7582 -8193
rect 7586 -8220 7672 -8210
rect 7676 -8220 8042 -8193
rect 8046 -8220 8132 -8210
rect 8136 -8220 8870 -8193
rect 8874 -8220 8960 -8210
rect 8964 -8220 9330 -8193
rect 9334 -8220 9420 -8210
rect 9424 -8220 10158 -8193
rect 10162 -8220 10248 -8210
rect 10344 -8220 10710 -8193
rect 10712 -8220 11446 -8193
rect 11450 -8220 11536 -8210
rect 11632 -8220 11998 -8193
rect 12025 -8196 12069 -8162
rect 12665 -8182 12709 -8148
rect 12761 -8196 12805 -8162
rect 13401 -8182 13445 -8148
rect 13564 -8151 14666 -8124
rect 14670 -8134 14756 -8124
rect 14760 -8151 15862 -8124
rect 15866 -8134 15952 -8124
rect 15956 -8151 16690 -8124
rect 13511 -8183 13535 -8161
rect 13592 -8189 13626 -8151
rect 13684 -8193 13718 -8155
rect 14788 -8189 14822 -8151
rect 15984 -8189 16018 -8151
rect 16628 -8193 16662 -8155
rect 13566 -8220 13652 -8210
rect 13656 -8220 15477 -8193
rect 15498 -8220 15584 -8210
rect 15588 -8220 16690 -8193
rect -3034 -8368 16729 -8220
rect 524 -8375 1036 -8368
rect 3100 -8375 3612 -8368
rect 5676 -8375 6188 -8368
rect 8252 -8375 8764 -8368
rect 10828 -8375 11340 -8368
rect 514 -9064 1026 -9057
rect 3090 -9064 3602 -9057
rect 5666 -9064 6178 -9057
rect 8242 -9064 8754 -9057
rect 10818 -9064 11330 -9057
rect -3035 -9212 16728 -9064
rect -2996 -9239 -2262 -9212
rect -2258 -9222 -2172 -9212
rect -1616 -9239 -882 -9212
rect -880 -9239 -146 -9212
rect -142 -9222 -56 -9212
rect -52 -9239 314 -9212
rect 318 -9222 404 -9212
rect 408 -9239 1142 -9212
rect 1146 -9222 1232 -9212
rect 1236 -9239 1602 -9212
rect 1606 -9222 1692 -9212
rect 1696 -9239 2430 -9212
rect 2434 -9222 2520 -9212
rect 2524 -9239 2890 -9212
rect 2894 -9222 2980 -9212
rect 2984 -9239 3718 -9212
rect 3722 -9222 3808 -9212
rect 3812 -9239 4178 -9212
rect 4182 -9222 4268 -9212
rect 4272 -9239 5006 -9212
rect 5010 -9222 5096 -9212
rect 5100 -9239 5466 -9212
rect 5470 -9222 5556 -9212
rect 5560 -9239 6294 -9212
rect 6298 -9222 6384 -9212
rect 6388 -9239 6754 -9212
rect 6758 -9222 6844 -9212
rect 6848 -9239 7582 -9212
rect 7586 -9222 7672 -9212
rect 7676 -9239 8042 -9212
rect 8046 -9222 8132 -9212
rect 8136 -9239 8870 -9212
rect 8874 -9222 8960 -9212
rect 8964 -9239 9330 -9212
rect 9334 -9222 9420 -9212
rect 9424 -9239 10158 -9212
rect 10162 -9222 10248 -9212
rect 10344 -9239 10710 -9212
rect 10712 -9239 11446 -9212
rect 11450 -9222 11536 -9212
rect 11632 -9239 11998 -9212
rect 12370 -9222 12456 -9212
rect 12541 -9239 13026 -9212
rect 13106 -9222 13192 -9212
rect 13196 -9239 13562 -9212
rect 13566 -9222 13652 -9212
rect 13656 -9239 15477 -9212
rect 15498 -9222 15584 -9212
rect 15588 -9239 16690 -9212
rect -2968 -9277 -2934 -9239
rect -2324 -9281 -2290 -9243
rect -2134 -9272 -2112 -9248
rect -1858 -9272 -1836 -9248
rect -1770 -9270 -1738 -9248
rect -1680 -9272 -1648 -9250
rect -1588 -9277 -1554 -9239
rect -944 -9281 -910 -9243
rect -852 -9277 -818 -9239
rect -209 -9281 -175 -9243
rect 252 -9281 286 -9239
rect 437 -9277 471 -9239
rect 1079 -9281 1113 -9243
rect 1540 -9281 1574 -9239
rect 1724 -9277 1758 -9239
rect 2368 -9281 2402 -9243
rect 2828 -9281 2862 -9239
rect 3013 -9277 3047 -9239
rect 3655 -9281 3689 -9243
rect 4116 -9281 4150 -9239
rect 4300 -9277 4334 -9239
rect 4944 -9281 4978 -9243
rect 5404 -9281 5438 -9239
rect 5589 -9277 5623 -9239
rect 6231 -9281 6265 -9243
rect 6692 -9281 6726 -9239
rect 6876 -9277 6910 -9239
rect 7520 -9281 7554 -9243
rect 7980 -9281 8014 -9239
rect 8165 -9277 8199 -9239
rect 8807 -9281 8841 -9243
rect 9268 -9281 9302 -9239
rect 9452 -9277 9486 -9239
rect 10096 -9281 10130 -9243
rect 10648 -9249 10682 -9239
rect 10291 -9271 10315 -9249
rect 10648 -9271 10683 -9249
rect 10648 -9281 10682 -9271
rect 10741 -9277 10775 -9239
rect 11383 -9281 11417 -9243
rect 11579 -9271 11603 -9249
rect 11936 -9281 11970 -9239
rect 12034 -9272 12056 -9248
rect 12488 -9277 12522 -9243
rect 12665 -9270 12709 -9239
rect 13224 -9277 13258 -9239
rect 13401 -9270 13445 -9239
rect 13511 -9271 13535 -9249
rect 13684 -9281 13718 -9239
rect 15616 -9277 15650 -9239
rect 16628 -9281 16662 -9243
rect -2996 -9308 -2262 -9281
rect -2258 -9308 -2172 -9298
rect -1616 -9308 -882 -9281
rect -880 -9308 -146 -9281
rect -142 -9308 -56 -9298
rect -52 -9308 314 -9281
rect 318 -9308 404 -9298
rect 408 -9308 1142 -9281
rect 1146 -9308 1232 -9298
rect 1236 -9308 1602 -9281
rect 1606 -9308 1692 -9298
rect 1696 -9308 2430 -9281
rect 2434 -9308 2520 -9298
rect 2524 -9308 2890 -9281
rect 2894 -9308 2980 -9298
rect 2984 -9308 3718 -9281
rect 3722 -9308 3808 -9298
rect 3812 -9308 4178 -9281
rect 4182 -9308 4268 -9298
rect 4272 -9308 5006 -9281
rect 5010 -9308 5096 -9298
rect 5100 -9308 5466 -9281
rect 5470 -9308 5556 -9298
rect 5560 -9308 6294 -9281
rect 6298 -9308 6384 -9298
rect 6388 -9308 6754 -9281
rect 6758 -9308 6844 -9298
rect 6848 -9308 7582 -9281
rect 7586 -9308 7672 -9298
rect 7676 -9308 8042 -9281
rect 8046 -9308 8132 -9298
rect 8136 -9308 8870 -9281
rect 8874 -9308 8960 -9298
rect 8964 -9308 9330 -9281
rect 9334 -9308 9420 -9298
rect 9424 -9308 10158 -9281
rect 10162 -9308 10248 -9298
rect 10344 -9308 10710 -9281
rect 10712 -9308 11446 -9281
rect 11450 -9308 11536 -9298
rect 11632 -9308 11998 -9281
rect 13566 -9308 13652 -9298
rect 13656 -9308 15477 -9281
rect 15498 -9308 15584 -9298
rect 15588 -9308 16690 -9281
rect -3034 -9456 16729 -9308
rect -764 -9463 -252 -9456
rect 524 -9463 1036 -9456
rect 3100 -9463 3612 -9456
rect 5676 -9463 6188 -9456
rect 8252 -9463 8764 -9456
rect 10828 -9463 11340 -9456
rect 514 -10152 1026 -10145
rect 3090 -10152 3602 -10145
rect 5666 -10152 6178 -10145
rect 8242 -10152 8754 -10145
rect 10818 -10152 11330 -10145
rect -3035 -10300 16728 -10152
rect -2996 -10327 -2262 -10300
rect -2258 -10310 -2172 -10300
rect -1616 -10327 -882 -10300
rect -880 -10327 -146 -10300
rect -142 -10310 -56 -10300
rect -52 -10327 314 -10300
rect 318 -10310 404 -10300
rect 408 -10327 1142 -10300
rect 1146 -10310 1232 -10300
rect 1236 -10327 1602 -10300
rect 1606 -10310 1692 -10300
rect 1696 -10327 2430 -10300
rect 2434 -10310 2520 -10300
rect 2524 -10327 2890 -10300
rect 2894 -10310 2980 -10300
rect 2984 -10327 3718 -10300
rect 3722 -10310 3808 -10300
rect 3812 -10327 4178 -10300
rect 4182 -10310 4268 -10300
rect 4272 -10327 5006 -10300
rect 5010 -10310 5096 -10300
rect 5100 -10327 5466 -10300
rect 5470 -10310 5556 -10300
rect 5560 -10327 6294 -10300
rect 6298 -10310 6384 -10300
rect 6388 -10327 6754 -10300
rect 6758 -10310 6844 -10300
rect 6848 -10327 7582 -10300
rect 7586 -10310 7672 -10300
rect 7676 -10327 8042 -10300
rect 8046 -10310 8132 -10300
rect 8136 -10327 8870 -10300
rect 8874 -10310 8960 -10300
rect 8964 -10327 9330 -10300
rect 9334 -10310 9420 -10300
rect 9424 -10327 10158 -10300
rect 10162 -10310 10248 -10300
rect 10344 -10327 10710 -10300
rect 10712 -10327 11446 -10300
rect 11450 -10310 11536 -10300
rect 11632 -10327 11998 -10300
rect 12370 -10310 12456 -10300
rect 12541 -10327 13026 -10300
rect 13106 -10310 13192 -10300
rect 13196 -10327 13562 -10300
rect 13566 -10310 13652 -10300
rect 13656 -10327 15477 -10300
rect 15498 -10310 15584 -10300
rect 15588 -10327 16690 -10300
rect -2968 -10365 -2934 -10327
rect -2324 -10369 -2290 -10331
rect -2134 -10360 -2112 -10336
rect -2048 -10360 -2016 -10338
rect -1956 -10365 -1922 -10331
rect -1770 -10358 -1738 -10336
rect -1588 -10365 -1554 -10327
rect -944 -10369 -910 -10331
rect -852 -10365 -818 -10327
rect -208 -10369 -174 -10331
rect 252 -10369 286 -10327
rect 437 -10365 471 -10327
rect 1079 -10369 1113 -10331
rect 1540 -10369 1574 -10327
rect 1724 -10365 1758 -10327
rect 2368 -10369 2402 -10331
rect 2828 -10369 2862 -10327
rect 3013 -10365 3047 -10327
rect 3655 -10369 3689 -10331
rect 4116 -10369 4150 -10327
rect 4300 -10365 4334 -10327
rect 4944 -10369 4978 -10331
rect 5404 -10369 5438 -10327
rect 5589 -10365 5623 -10327
rect 6231 -10369 6265 -10331
rect 6692 -10369 6726 -10327
rect 6876 -10365 6910 -10327
rect 7520 -10369 7554 -10331
rect 7980 -10369 8014 -10327
rect 8165 -10365 8199 -10327
rect 8807 -10369 8841 -10331
rect 9268 -10369 9302 -10327
rect 9452 -10365 9486 -10327
rect 10096 -10369 10130 -10331
rect 10648 -10337 10682 -10327
rect 10291 -10359 10315 -10337
rect 10648 -10359 10683 -10337
rect 10648 -10369 10682 -10359
rect 10741 -10365 10775 -10327
rect 11383 -10369 11417 -10331
rect 11579 -10359 11603 -10337
rect 11936 -10369 11970 -10327
rect 12034 -10360 12056 -10336
rect 12488 -10365 12522 -10331
rect 12665 -10358 12709 -10327
rect 13224 -10365 13258 -10327
rect 13401 -10358 13445 -10327
rect 13684 -10365 13718 -10327
rect 14604 -10369 14638 -10331
rect 15616 -10365 15650 -10327
rect 15800 -10369 15834 -10331
rect 16628 -10369 16662 -10331
rect -2996 -10396 -2262 -10369
rect -2258 -10396 -2172 -10386
rect -1901 -10396 -1710 -10369
rect -1706 -10396 -1620 -10386
rect -1616 -10396 -882 -10369
rect -880 -10396 -146 -10369
rect -142 -10396 -56 -10386
rect -52 -10396 314 -10369
rect 318 -10396 404 -10386
rect 408 -10396 1142 -10369
rect 1146 -10396 1232 -10386
rect 1236 -10396 1602 -10369
rect 1606 -10396 1692 -10386
rect 1696 -10396 2430 -10369
rect 2434 -10396 2520 -10386
rect 2524 -10396 2890 -10369
rect 2894 -10396 2980 -10386
rect 2984 -10396 3718 -10369
rect 3722 -10396 3808 -10386
rect 3812 -10396 4178 -10369
rect 4182 -10396 4268 -10386
rect 4272 -10396 5006 -10369
rect 5010 -10396 5096 -10386
rect 5100 -10396 5466 -10369
rect 5470 -10396 5556 -10386
rect 5560 -10396 6294 -10369
rect 6298 -10396 6384 -10386
rect 6388 -10396 6754 -10369
rect 6758 -10396 6844 -10386
rect 6848 -10396 7582 -10369
rect 7586 -10396 7672 -10386
rect 7676 -10396 8042 -10369
rect 8046 -10396 8132 -10386
rect 8136 -10396 8870 -10369
rect 8874 -10396 8960 -10386
rect 8964 -10396 9330 -10369
rect 9334 -10396 9420 -10386
rect 9424 -10396 10158 -10369
rect 10162 -10396 10248 -10386
rect 10344 -10396 10710 -10369
rect 10712 -10396 11446 -10369
rect 11450 -10396 11536 -10386
rect 11632 -10396 11998 -10369
rect 13474 -10396 13560 -10386
rect 13564 -10396 14666 -10369
rect 14670 -10396 14756 -10386
rect 14760 -10396 15862 -10369
rect 15866 -10396 15952 -10386
rect 15956 -10396 16690 -10369
rect -3034 -10544 16729 -10396
rect 524 -10551 1036 -10544
rect 3100 -10551 3612 -10544
rect 5676 -10551 6188 -10544
rect 8252 -10551 8764 -10544
rect 10828 -10551 11340 -10544
rect 524 -11240 1036 -11233
rect 3100 -11240 3612 -11233
rect 5676 -11240 6188 -11233
rect 8252 -11240 8764 -11233
rect 10828 -11240 11340 -11233
rect -3035 -11388 16728 -11240
rect -2996 -11415 -2262 -11388
rect -2258 -11398 -2172 -11388
rect -1616 -11415 -882 -11388
rect -880 -11415 -146 -11388
rect -142 -11398 -56 -11388
rect -52 -11415 314 -11388
rect 318 -11398 404 -11388
rect 408 -11415 1142 -11388
rect 1146 -11398 1232 -11388
rect 1236 -11415 1602 -11388
rect 1606 -11398 1692 -11388
rect 1696 -11415 2430 -11388
rect 2434 -11398 2520 -11388
rect 2524 -11415 2890 -11388
rect 2894 -11398 2980 -11388
rect 2984 -11415 3718 -11388
rect 3722 -11398 3808 -11388
rect 3812 -11415 4178 -11388
rect 4182 -11398 4268 -11388
rect 4272 -11415 5006 -11388
rect 5010 -11398 5096 -11388
rect 5100 -11415 5466 -11388
rect 5470 -11398 5556 -11388
rect 5560 -11415 6294 -11388
rect 6298 -11398 6384 -11388
rect 6388 -11415 6754 -11388
rect 6758 -11398 6844 -11388
rect 6848 -11415 7582 -11388
rect 7586 -11398 7672 -11388
rect 7676 -11415 8042 -11388
rect 8046 -11398 8132 -11388
rect 8136 -11415 8870 -11388
rect 8874 -11398 8960 -11388
rect 8964 -11415 9330 -11388
rect 9334 -11398 9420 -11388
rect 9424 -11415 10158 -11388
rect 10162 -11398 10248 -11388
rect 10344 -11415 10710 -11388
rect 10712 -11415 11446 -11388
rect 11450 -11398 11536 -11388
rect 11632 -11415 11998 -11388
rect 13474 -11398 13560 -11388
rect 13564 -11415 14666 -11388
rect 14670 -11398 14756 -11388
rect 14760 -11415 15862 -11388
rect 15866 -11398 15952 -11388
rect 15956 -11415 16690 -11388
rect -2968 -11453 -2934 -11415
rect -2324 -11457 -2290 -11419
rect -2134 -11448 -2112 -11424
rect -1858 -11448 -1836 -11424
rect -1770 -11446 -1738 -11424
rect -1680 -11448 -1648 -11426
rect -1588 -11457 -1554 -11419
rect -944 -11453 -910 -11415
rect -852 -11457 -818 -11419
rect -208 -11453 -174 -11415
rect 252 -11457 286 -11415
rect 437 -11457 471 -11419
rect 1079 -11453 1113 -11415
rect 1540 -11457 1574 -11415
rect 1724 -11453 1758 -11415
rect 2368 -11457 2402 -11419
rect 2828 -11457 2862 -11415
rect 3013 -11457 3047 -11419
rect 3655 -11453 3689 -11415
rect 4116 -11457 4150 -11415
rect 4300 -11453 4334 -11415
rect 4944 -11457 4978 -11419
rect 5404 -11457 5438 -11415
rect 5589 -11457 5623 -11419
rect 6231 -11453 6265 -11415
rect 6692 -11457 6726 -11415
rect 6876 -11453 6910 -11415
rect 7520 -11457 7554 -11419
rect 7980 -11457 8014 -11415
rect 8165 -11457 8199 -11419
rect 8807 -11453 8841 -11415
rect 9268 -11457 9302 -11415
rect 9452 -11453 9486 -11415
rect 10096 -11457 10130 -11419
rect 10648 -11425 10682 -11415
rect 10291 -11447 10315 -11425
rect 10648 -11447 10683 -11425
rect 10648 -11457 10682 -11447
rect 10741 -11457 10775 -11419
rect 11383 -11453 11417 -11415
rect 11579 -11447 11603 -11425
rect 11936 -11457 11970 -11415
rect 12034 -11448 12056 -11424
rect 12488 -11453 12522 -11419
rect 12665 -11457 12709 -11426
rect 13224 -11457 13258 -11419
rect 13401 -11457 13445 -11426
rect 13684 -11457 13718 -11419
rect 14604 -11453 14638 -11415
rect 15616 -11457 15650 -11419
rect 15800 -11453 15834 -11415
rect 16628 -11453 16662 -11415
rect -2996 -11484 -2262 -11457
rect -2258 -11484 -2172 -11474
rect -1616 -11484 -882 -11457
rect -880 -11484 -146 -11457
rect -142 -11484 -56 -11474
rect -52 -11484 314 -11457
rect 318 -11484 404 -11474
rect 408 -11484 1142 -11457
rect 1146 -11484 1232 -11474
rect 1236 -11484 1602 -11457
rect 1606 -11484 1692 -11474
rect 1696 -11484 2430 -11457
rect 2434 -11484 2520 -11474
rect 2524 -11484 2890 -11457
rect 2894 -11484 2980 -11474
rect 2984 -11484 3718 -11457
rect 3722 -11484 3808 -11474
rect 3812 -11484 4178 -11457
rect 4182 -11484 4268 -11474
rect 4272 -11484 5006 -11457
rect 5010 -11484 5096 -11474
rect 5100 -11484 5466 -11457
rect 5470 -11484 5556 -11474
rect 5560 -11484 6294 -11457
rect 6298 -11484 6384 -11474
rect 6388 -11484 6754 -11457
rect 6758 -11484 6844 -11474
rect 6848 -11484 7582 -11457
rect 7586 -11484 7672 -11474
rect 7676 -11484 8042 -11457
rect 8046 -11484 8132 -11474
rect 8136 -11484 8870 -11457
rect 8874 -11484 8960 -11474
rect 8964 -11484 9330 -11457
rect 9334 -11484 9420 -11474
rect 9424 -11484 10158 -11457
rect 10162 -11484 10248 -11474
rect 10344 -11484 10710 -11457
rect 10712 -11484 11446 -11457
rect 11450 -11484 11536 -11474
rect 11632 -11484 11998 -11457
rect 12370 -11484 12456 -11474
rect 12541 -11484 13026 -11457
rect 13106 -11484 13192 -11474
rect 13196 -11484 13562 -11457
rect 13566 -11484 13652 -11474
rect 13656 -11484 15477 -11457
rect 15498 -11484 15584 -11474
rect 15588 -11484 16690 -11457
rect -3034 -11632 16729 -11484
rect 514 -11639 1026 -11632
rect 3090 -11639 3602 -11632
rect 5666 -11639 6178 -11632
rect 8242 -11639 8754 -11632
rect 10818 -11639 11330 -11632
rect -764 -12328 -252 -12321
rect 524 -12328 1036 -12321
rect 3100 -12328 3612 -12321
rect 5676 -12328 6188 -12321
rect 8252 -12328 8764 -12321
rect 10828 -12328 11340 -12321
rect -3035 -12476 16728 -12328
rect -2996 -12503 -2262 -12476
rect -2258 -12486 -2172 -12476
rect -1616 -12503 -882 -12476
rect -880 -12503 -146 -12476
rect -142 -12486 -56 -12476
rect -52 -12503 314 -12476
rect 318 -12486 404 -12476
rect 408 -12503 1142 -12476
rect 1146 -12486 1232 -12476
rect 1236 -12503 1602 -12476
rect 1606 -12486 1692 -12476
rect 1696 -12503 2430 -12476
rect 2434 -12486 2520 -12476
rect 2524 -12503 2890 -12476
rect 2894 -12486 2980 -12476
rect 2984 -12503 3718 -12476
rect 3722 -12486 3808 -12476
rect 3812 -12503 4178 -12476
rect 4182 -12486 4268 -12476
rect 4272 -12503 5006 -12476
rect 5010 -12486 5096 -12476
rect 5100 -12503 5466 -12476
rect 5470 -12486 5556 -12476
rect 5560 -12503 6294 -12476
rect 6298 -12486 6384 -12476
rect 6388 -12503 6754 -12476
rect 6758 -12486 6844 -12476
rect 6848 -12503 7582 -12476
rect 7586 -12486 7672 -12476
rect 7676 -12503 8042 -12476
rect 8046 -12486 8132 -12476
rect 8136 -12503 8870 -12476
rect 8874 -12486 8960 -12476
rect 8964 -12503 9330 -12476
rect 9334 -12486 9420 -12476
rect 9424 -12503 10158 -12476
rect 10162 -12486 10248 -12476
rect 10344 -12503 10710 -12476
rect 10712 -12503 11446 -12476
rect 11450 -12486 11536 -12476
rect 11632 -12503 11998 -12476
rect 13566 -12486 13652 -12476
rect 13656 -12503 15477 -12476
rect 15498 -12486 15584 -12476
rect 15588 -12503 16690 -12476
rect -2968 -12541 -2934 -12503
rect -2324 -12545 -2290 -12507
rect -2134 -12536 -2112 -12512
rect -1858 -12536 -1836 -12512
rect -1770 -12534 -1738 -12512
rect -1680 -12536 -1648 -12514
rect -1588 -12545 -1554 -12507
rect -944 -12541 -910 -12503
rect -852 -12545 -818 -12507
rect -209 -12541 -175 -12503
rect 252 -12545 286 -12503
rect 437 -12545 471 -12507
rect 1079 -12541 1113 -12503
rect 1540 -12545 1574 -12503
rect 1724 -12541 1758 -12503
rect 2368 -12545 2402 -12507
rect 2828 -12545 2862 -12503
rect 3013 -12545 3047 -12507
rect 3655 -12541 3689 -12503
rect 4116 -12545 4150 -12503
rect 4300 -12541 4334 -12503
rect 4944 -12545 4978 -12507
rect 5404 -12545 5438 -12503
rect 5589 -12545 5623 -12507
rect 6231 -12541 6265 -12503
rect 6692 -12545 6726 -12503
rect 6876 -12541 6910 -12503
rect 7520 -12545 7554 -12507
rect 7980 -12545 8014 -12503
rect 8165 -12545 8199 -12507
rect 8807 -12541 8841 -12503
rect 9268 -12545 9302 -12503
rect 9452 -12541 9486 -12503
rect 10096 -12545 10130 -12507
rect 10648 -12513 10682 -12503
rect 10291 -12535 10315 -12513
rect 10648 -12535 10683 -12513
rect 10648 -12545 10682 -12535
rect 10741 -12545 10775 -12507
rect 11383 -12541 11417 -12503
rect 11579 -12535 11603 -12513
rect 11936 -12545 11970 -12503
rect 12034 -12536 12056 -12512
rect 12488 -12541 12522 -12507
rect 12665 -12545 12709 -12514
rect 13224 -12545 13258 -12507
rect 13401 -12545 13445 -12514
rect 13511 -12535 13535 -12513
rect 13684 -12545 13718 -12503
rect 15616 -12545 15650 -12507
rect 16628 -12541 16662 -12503
rect -2996 -12572 -2262 -12545
rect -2258 -12572 -2172 -12562
rect -1616 -12572 -882 -12545
rect -880 -12572 -146 -12545
rect -142 -12572 -56 -12562
rect -52 -12572 314 -12545
rect 318 -12572 404 -12562
rect 408 -12572 1142 -12545
rect 1146 -12572 1232 -12562
rect 1236 -12572 1602 -12545
rect 1606 -12572 1692 -12562
rect 1696 -12572 2430 -12545
rect 2434 -12572 2520 -12562
rect 2524 -12572 2890 -12545
rect 2894 -12572 2980 -12562
rect 2984 -12572 3718 -12545
rect 3722 -12572 3808 -12562
rect 3812 -12572 4178 -12545
rect 4182 -12572 4268 -12562
rect 4272 -12572 5006 -12545
rect 5010 -12572 5096 -12562
rect 5100 -12572 5466 -12545
rect 5470 -12572 5556 -12562
rect 5560 -12572 6294 -12545
rect 6298 -12572 6384 -12562
rect 6388 -12572 6754 -12545
rect 6758 -12572 6844 -12562
rect 6848 -12572 7582 -12545
rect 7586 -12572 7672 -12562
rect 7676 -12572 8042 -12545
rect 8046 -12572 8132 -12562
rect 8136 -12572 8870 -12545
rect 8874 -12572 8960 -12562
rect 8964 -12572 9330 -12545
rect 9334 -12572 9420 -12562
rect 9424 -12572 10158 -12545
rect 10162 -12572 10248 -12562
rect 10344 -12572 10710 -12545
rect 10712 -12572 11446 -12545
rect 11450 -12572 11536 -12562
rect 11632 -12572 11998 -12545
rect 12370 -12572 12456 -12562
rect 12541 -12572 13026 -12545
rect 13106 -12572 13192 -12562
rect 13196 -12572 13562 -12545
rect 13566 -12572 13652 -12562
rect 13656 -12572 15477 -12545
rect 15498 -12572 15584 -12562
rect 15588 -12572 16690 -12545
rect -3034 -12720 16729 -12572
rect 514 -12727 1026 -12720
rect 3090 -12727 3602 -12720
rect 5666 -12727 6178 -12720
rect 8242 -12727 8754 -12720
rect 10818 -12727 11330 -12720
rect 524 -13416 1036 -13409
rect 3100 -13416 3612 -13409
rect 5676 -13416 6188 -13409
rect 8252 -13416 8764 -13409
rect 10828 -13416 11340 -13409
rect -3035 -13564 16728 -13416
rect -2996 -13591 -2262 -13564
rect -2258 -13574 -2172 -13564
rect -1616 -13591 -882 -13564
rect -880 -13591 -146 -13564
rect -142 -13574 -56 -13564
rect -52 -13591 314 -13564
rect 318 -13574 404 -13564
rect 408 -13591 1142 -13564
rect 1146 -13574 1232 -13564
rect 1236 -13591 1602 -13564
rect 1606 -13574 1692 -13564
rect 1696 -13591 2430 -13564
rect 2434 -13574 2520 -13564
rect 2524 -13591 2890 -13564
rect 2894 -13574 2980 -13564
rect 2984 -13591 3718 -13564
rect 3722 -13574 3808 -13564
rect 3812 -13591 4178 -13564
rect 4182 -13574 4268 -13564
rect 4272 -13591 5006 -13564
rect 5010 -13574 5096 -13564
rect 5100 -13591 5466 -13564
rect 5470 -13574 5556 -13564
rect 5560 -13591 6294 -13564
rect 6298 -13574 6384 -13564
rect 6388 -13591 6754 -13564
rect 6758 -13574 6844 -13564
rect 6848 -13591 7582 -13564
rect 7586 -13574 7672 -13564
rect 7676 -13591 8042 -13564
rect 8046 -13574 8132 -13564
rect 8136 -13591 8870 -13564
rect 8874 -13574 8960 -13564
rect 8964 -13591 9330 -13564
rect 9334 -13574 9420 -13564
rect 9424 -13591 10158 -13564
rect 10162 -13574 10248 -13564
rect 10344 -13591 10710 -13564
rect 10712 -13591 11446 -13564
rect 11450 -13574 11536 -13564
rect 11632 -13591 11998 -13564
rect 13566 -13574 13652 -13564
rect -2968 -13629 -2934 -13591
rect -944 -13595 -910 -13591
rect -2324 -13633 -2290 -13595
rect -2134 -13624 -2112 -13600
rect -1858 -13624 -1836 -13600
rect -1770 -13622 -1738 -13600
rect -1680 -13624 -1648 -13602
rect -1586 -13624 -1554 -13602
rect -1404 -13633 -1370 -13595
rect -945 -13629 -910 -13595
rect -945 -13633 -911 -13629
rect -576 -13633 -542 -13595
rect -208 -13629 -174 -13591
rect -116 -13629 -82 -13595
rect 252 -13629 286 -13591
rect 1079 -13595 1113 -13591
rect 620 -13633 654 -13595
rect 1079 -13629 1114 -13595
rect 1448 -13633 1482 -13595
rect 1540 -13629 1574 -13591
rect 1724 -13629 1758 -13591
rect 1908 -13633 1942 -13595
rect 2369 -13633 2403 -13595
rect 2828 -13629 2862 -13591
rect 3196 -13633 3230 -13595
rect 3653 -13622 3697 -13591
rect 3655 -13629 3689 -13622
rect 4116 -13629 4150 -13591
rect 4300 -13629 4334 -13591
rect 4392 -13633 4426 -13595
rect 5404 -13629 5438 -13591
rect 5502 -13624 5524 -13600
rect 5863 -13623 5887 -13601
rect 5962 -13624 5984 -13600
rect 6231 -13629 6265 -13591
rect 6416 -13633 6450 -13595
rect 6692 -13629 6726 -13591
rect 6876 -13595 6910 -13591
rect 6876 -13629 6911 -13595
rect 6877 -13633 6911 -13629
rect 7704 -13633 7738 -13595
rect 7980 -13629 8014 -13591
rect 8165 -13633 8199 -13595
rect 8807 -13629 8841 -13591
rect 8992 -13633 9026 -13595
rect 9268 -13629 9302 -13591
rect 9452 -13595 9486 -13591
rect 9452 -13629 9487 -13595
rect 9453 -13633 9487 -13629
rect 10280 -13601 10314 -13595
rect 10648 -13601 10682 -13591
rect 10280 -13623 10315 -13601
rect 10648 -13623 10683 -13601
rect 10280 -13633 10314 -13623
rect 10648 -13629 10682 -13623
rect 10741 -13633 10775 -13595
rect 11383 -13629 11417 -13591
rect 11579 -13623 11603 -13601
rect 11660 -13633 11694 -13595
rect 11936 -13629 11970 -13591
rect 12025 -13622 12069 -13588
rect -2996 -13660 -2262 -13633
rect -2258 -13660 -2172 -13650
rect -1432 -13660 -1066 -13633
rect -1062 -13660 -976 -13650
rect -968 -13660 -698 -13633
rect -694 -13660 -608 -13650
rect -604 -13660 -238 -13633
rect -234 -13660 -148 -13650
rect -63 -13660 422 -13633
rect 502 -13660 588 -13650
rect 592 -13660 958 -13633
rect 962 -13660 1048 -13650
rect 1135 -13660 1326 -13633
rect 1330 -13660 1416 -13650
rect 1420 -13660 1786 -13633
rect 1790 -13660 1876 -13650
rect 1880 -13660 2246 -13633
rect 2250 -13660 2336 -13650
rect 2340 -13660 3074 -13633
rect 3078 -13660 3164 -13650
rect 3168 -13660 3534 -13633
rect 3538 -13660 3624 -13650
rect 4364 -13660 5466 -13633
rect 6298 -13660 6384 -13650
rect 6388 -13660 6754 -13633
rect 6758 -13660 6844 -13650
rect 6848 -13660 7582 -13633
rect 7586 -13660 7672 -13650
rect 7676 -13660 8042 -13633
rect 8046 -13660 8132 -13650
rect 8136 -13660 8870 -13633
rect 8874 -13660 8960 -13650
rect 8964 -13660 9330 -13633
rect 9334 -13660 9420 -13650
rect 9424 -13660 10158 -13633
rect 10162 -13660 10248 -13650
rect 10252 -13660 10618 -13633
rect 10622 -13660 10708 -13650
rect 10712 -13660 11486 -13633
rect 11542 -13660 11628 -13650
rect 11632 -13660 11998 -13633
rect 12665 -13636 12709 -13602
rect 12761 -13622 12805 -13588
rect 13656 -13591 15477 -13564
rect 15498 -13574 15584 -13564
rect 15588 -13591 16690 -13564
rect 13401 -13636 13445 -13602
rect 13511 -13623 13535 -13601
rect 13592 -13633 13626 -13595
rect 13684 -13629 13718 -13591
rect 14788 -13633 14822 -13595
rect 15984 -13633 16018 -13595
rect 16628 -13629 16662 -13591
rect 13474 -13660 13560 -13650
rect 13564 -13660 14666 -13633
rect 14670 -13660 14756 -13650
rect 14760 -13660 15862 -13633
rect 15866 -13660 15952 -13650
rect 15956 -13660 16690 -13633
rect -3034 -13808 16729 -13660
rect -968 -13815 -698 -13808
rect 2446 -13815 2958 -13808
rect 6954 -13815 7466 -13808
rect 8242 -13815 8754 -13808
rect 9530 -13815 10042 -13808
rect 10712 -13815 11486 -13808
<< scnmos >>
rect -2918 -509 -2340 -399
rect -1354 -509 -1144 -399
rect -890 -509 -860 -379
rect -806 -509 -776 -379
rect -526 -509 -316 -399
rect 29 -509 59 -425
rect 115 -509 145 -425
rect 201 -509 231 -425
rect 287 -509 317 -425
rect 670 -509 880 -399
rect 1213 -509 1243 -425
rect 1498 -509 1708 -399
rect 1958 -509 2168 -399
rect 2420 -509 2450 -425
rect 2522 -509 2622 -379
rect 2782 -509 2882 -379
rect 2947 -509 2977 -425
rect 3246 -509 3456 -399
rect 4442 -509 5388 -399
rect 6466 -509 6676 -399
rect 6928 -509 6958 -425
rect 7030 -509 7130 -379
rect 7290 -509 7390 -379
rect 7455 -509 7485 -425
rect 7754 -509 7964 -399
rect 8216 -509 8246 -425
rect 8318 -509 8418 -379
rect 8578 -509 8678 -379
rect 8743 -509 8773 -425
rect 9042 -509 9252 -399
rect 9504 -509 9534 -425
rect 9606 -509 9706 -379
rect 9866 -509 9966 -379
rect 10031 -509 10061 -425
rect 10330 -509 10540 -399
rect 10790 -509 10820 -379
rect 10874 -509 10904 -379
rect 10958 -509 10988 -379
rect 11042 -509 11072 -379
rect 11126 -509 11156 -379
rect 11210 -509 11240 -379
rect 11294 -509 11324 -379
rect 11378 -509 11408 -379
rect 11710 -509 11920 -399
rect 13642 -509 14588 -399
rect 14838 -509 15784 -399
rect 16034 -509 16612 -399
rect -2918 -713 -2340 -603
rect -1538 -713 -960 -603
rect -802 -713 -224 -603
rect 26 -713 236 -603
rect 505 -687 535 -603
rect 600 -733 700 -603
rect 860 -733 960 -603
rect 1032 -687 1062 -603
rect 1314 -713 1524 -603
rect 1774 -713 2352 -603
rect 2602 -713 2812 -603
rect 3081 -687 3111 -603
rect 3176 -733 3276 -603
rect 3436 -733 3536 -603
rect 3608 -687 3638 -603
rect 3890 -713 4100 -603
rect 4350 -713 4928 -603
rect 5178 -713 5388 -603
rect 5657 -687 5687 -603
rect 5752 -733 5852 -603
rect 6012 -733 6112 -603
rect 6184 -687 6214 -603
rect 6466 -713 6676 -603
rect 6926 -713 7504 -603
rect 7754 -713 7964 -603
rect 8233 -687 8263 -603
rect 8328 -733 8428 -603
rect 8588 -733 8688 -603
rect 8760 -687 8790 -603
rect 9042 -713 9252 -603
rect 9502 -713 10080 -603
rect 10422 -713 10632 -603
rect 10809 -687 10839 -603
rect 10904 -733 11004 -603
rect 11164 -733 11264 -603
rect 11336 -687 11366 -603
rect 11710 -713 11920 -603
rect 13735 -687 13765 -603
rect 13821 -687 13851 -603
rect 13907 -687 13937 -603
rect 13993 -687 14023 -603
rect 14079 -687 14109 -603
rect 14165 -687 14195 -603
rect 14251 -687 14281 -603
rect 14337 -687 14367 -603
rect 14423 -687 14453 -603
rect 14509 -687 14539 -603
rect 14595 -687 14625 -603
rect 14681 -687 14711 -603
rect 14766 -687 14796 -603
rect 14852 -687 14882 -603
rect 14938 -687 14968 -603
rect 15024 -687 15054 -603
rect 15110 -687 15140 -603
rect 15196 -687 15226 -603
rect 15282 -687 15312 -603
rect 15368 -687 15398 -603
rect 15666 -713 16612 -603
rect -2918 -1597 -2340 -1487
rect -1538 -1597 -960 -1487
rect -802 -1597 -224 -1487
rect 26 -1597 236 -1487
rect 488 -1597 518 -1513
rect 590 -1597 690 -1467
rect 850 -1597 950 -1467
rect 1015 -1597 1045 -1513
rect 1314 -1597 1524 -1487
rect 1774 -1597 2352 -1487
rect 2602 -1597 2812 -1487
rect 3064 -1597 3094 -1513
rect 3166 -1597 3266 -1467
rect 3426 -1597 3526 -1467
rect 3591 -1597 3621 -1513
rect 3890 -1597 4100 -1487
rect 4350 -1597 4928 -1487
rect 5178 -1597 5388 -1487
rect 5640 -1597 5670 -1513
rect 5742 -1597 5842 -1467
rect 6002 -1597 6102 -1467
rect 6167 -1597 6197 -1513
rect 6466 -1597 6676 -1487
rect 6926 -1597 7504 -1487
rect 7754 -1597 7964 -1487
rect 8216 -1597 8246 -1513
rect 8318 -1597 8418 -1467
rect 8578 -1597 8678 -1467
rect 8743 -1597 8773 -1513
rect 9042 -1597 9252 -1487
rect 9502 -1597 10080 -1487
rect 10422 -1597 10632 -1487
rect 10792 -1597 10822 -1513
rect 10894 -1597 10994 -1467
rect 11154 -1597 11254 -1467
rect 11319 -1597 11349 -1513
rect 11710 -1597 11920 -1487
rect 12633 -1597 12663 -1513
rect 12719 -1597 12749 -1513
rect 12805 -1597 12835 -1513
rect 12891 -1597 12921 -1513
rect 13274 -1597 13484 -1487
rect 13735 -1597 13765 -1513
rect 13821 -1597 13851 -1513
rect 13907 -1597 13937 -1513
rect 13993 -1597 14023 -1513
rect 14079 -1597 14109 -1513
rect 14165 -1597 14195 -1513
rect 14251 -1597 14281 -1513
rect 14337 -1597 14367 -1513
rect 14423 -1597 14453 -1513
rect 14509 -1597 14539 -1513
rect 14595 -1597 14625 -1513
rect 14681 -1597 14711 -1513
rect 14766 -1597 14796 -1513
rect 14852 -1597 14882 -1513
rect 14938 -1597 14968 -1513
rect 15024 -1597 15054 -1513
rect 15110 -1597 15140 -1513
rect 15196 -1597 15226 -1513
rect 15282 -1597 15312 -1513
rect 15368 -1597 15398 -1513
rect 15666 -1597 16612 -1487
rect -2918 -1801 -2340 -1691
rect -1538 -1801 -960 -1691
rect -783 -1775 -753 -1691
rect -688 -1821 -588 -1691
rect -428 -1821 -328 -1691
rect -256 -1775 -226 -1691
rect 26 -1801 236 -1691
rect 505 -1775 535 -1691
rect 600 -1821 700 -1691
rect 860 -1821 960 -1691
rect 1032 -1775 1062 -1691
rect 1314 -1801 1524 -1691
rect 1774 -1801 2352 -1691
rect 2602 -1801 2812 -1691
rect 3081 -1775 3111 -1691
rect 3176 -1821 3276 -1691
rect 3436 -1821 3536 -1691
rect 3608 -1775 3638 -1691
rect 3890 -1801 4100 -1691
rect 4350 -1801 4928 -1691
rect 5178 -1801 5388 -1691
rect 5657 -1775 5687 -1691
rect 5752 -1821 5852 -1691
rect 6012 -1821 6112 -1691
rect 6184 -1775 6214 -1691
rect 6466 -1801 6676 -1691
rect 6926 -1801 7504 -1691
rect 7754 -1801 7964 -1691
rect 8233 -1775 8263 -1691
rect 8328 -1821 8428 -1691
rect 8588 -1821 8688 -1691
rect 8760 -1775 8790 -1691
rect 9042 -1801 9252 -1691
rect 9502 -1801 10080 -1691
rect 10422 -1801 10632 -1691
rect 10809 -1775 10839 -1691
rect 10904 -1821 11004 -1691
rect 11164 -1821 11264 -1691
rect 11336 -1775 11366 -1691
rect 11710 -1801 11920 -1691
rect 13735 -1775 13765 -1691
rect 13821 -1775 13851 -1691
rect 13907 -1775 13937 -1691
rect 13993 -1775 14023 -1691
rect 14079 -1775 14109 -1691
rect 14165 -1775 14195 -1691
rect 14251 -1775 14281 -1691
rect 14337 -1775 14367 -1691
rect 14423 -1775 14453 -1691
rect 14509 -1775 14539 -1691
rect 14595 -1775 14625 -1691
rect 14681 -1775 14711 -1691
rect 14766 -1775 14796 -1691
rect 14852 -1775 14882 -1691
rect 14938 -1775 14968 -1691
rect 15024 -1775 15054 -1691
rect 15110 -1775 15140 -1691
rect 15196 -1775 15226 -1691
rect 15282 -1775 15312 -1691
rect 15368 -1775 15398 -1691
rect 15666 -1801 16612 -1691
rect -2918 -2685 -2340 -2575
rect -1538 -2685 -960 -2575
rect -802 -2685 -224 -2575
rect 26 -2685 236 -2575
rect 488 -2685 518 -2601
rect 590 -2685 690 -2555
rect 850 -2685 950 -2555
rect 1015 -2685 1045 -2601
rect 1314 -2685 1524 -2575
rect 1774 -2685 2352 -2575
rect 2602 -2685 2812 -2575
rect 3064 -2685 3094 -2601
rect 3166 -2685 3266 -2555
rect 3426 -2685 3526 -2555
rect 3591 -2685 3621 -2601
rect 3890 -2685 4100 -2575
rect 4350 -2685 4928 -2575
rect 5178 -2685 5388 -2575
rect 5640 -2685 5670 -2601
rect 5742 -2685 5842 -2555
rect 6002 -2685 6102 -2555
rect 6167 -2685 6197 -2601
rect 6466 -2685 6676 -2575
rect 6926 -2685 7504 -2575
rect 7754 -2685 7964 -2575
rect 8216 -2685 8246 -2601
rect 8318 -2685 8418 -2555
rect 8578 -2685 8678 -2555
rect 8743 -2685 8773 -2601
rect 9042 -2685 9252 -2575
rect 9502 -2685 10080 -2575
rect 10422 -2685 10632 -2575
rect 10792 -2685 10822 -2601
rect 10894 -2685 10994 -2555
rect 11154 -2685 11254 -2555
rect 11319 -2685 11349 -2601
rect 11710 -2685 11920 -2575
rect 12633 -2685 12663 -2601
rect 12719 -2685 12749 -2601
rect 12805 -2685 12835 -2601
rect 12891 -2685 12921 -2601
rect 13274 -2685 13484 -2575
rect 13735 -2685 13765 -2601
rect 13821 -2685 13851 -2601
rect 13907 -2685 13937 -2601
rect 13993 -2685 14023 -2601
rect 14079 -2685 14109 -2601
rect 14165 -2685 14195 -2601
rect 14251 -2685 14281 -2601
rect 14337 -2685 14367 -2601
rect 14423 -2685 14453 -2601
rect 14509 -2685 14539 -2601
rect 14595 -2685 14625 -2601
rect 14681 -2685 14711 -2601
rect 14766 -2685 14796 -2601
rect 14852 -2685 14882 -2601
rect 14938 -2685 14968 -2601
rect 15024 -2685 15054 -2601
rect 15110 -2685 15140 -2601
rect 15196 -2685 15226 -2601
rect 15282 -2685 15312 -2601
rect 15368 -2685 15398 -2601
rect 15666 -2685 16612 -2575
rect -2918 -2889 -2340 -2779
rect -1823 -2863 -1793 -2779
rect -1538 -2889 -960 -2779
rect -802 -2889 -224 -2779
rect 26 -2889 236 -2779
rect 505 -2863 535 -2779
rect 600 -2909 700 -2779
rect 860 -2909 960 -2779
rect 1032 -2863 1062 -2779
rect 1314 -2889 1524 -2779
rect 1774 -2889 2352 -2779
rect 2602 -2889 2812 -2779
rect 3081 -2863 3111 -2779
rect 3176 -2909 3276 -2779
rect 3436 -2909 3536 -2779
rect 3608 -2863 3638 -2779
rect 3890 -2889 4100 -2779
rect 4350 -2889 4928 -2779
rect 5178 -2889 5388 -2779
rect 5657 -2863 5687 -2779
rect 5752 -2909 5852 -2779
rect 6012 -2909 6112 -2779
rect 6184 -2863 6214 -2779
rect 6466 -2889 6676 -2779
rect 6926 -2889 7504 -2779
rect 7754 -2889 7964 -2779
rect 8233 -2863 8263 -2779
rect 8328 -2909 8428 -2779
rect 8588 -2909 8688 -2779
rect 8760 -2863 8790 -2779
rect 9042 -2889 9252 -2779
rect 9502 -2889 10080 -2779
rect 10422 -2889 10632 -2779
rect 10809 -2863 10839 -2779
rect 10904 -2909 11004 -2779
rect 11164 -2909 11264 -2779
rect 11336 -2863 11366 -2779
rect 11710 -2889 11920 -2779
rect 13642 -2889 14588 -2779
rect 14838 -2889 15784 -2779
rect 16034 -2889 16612 -2779
rect -2918 -3773 -2340 -3663
rect -1538 -3773 -960 -3663
rect -802 -3773 -224 -3663
rect 26 -3773 236 -3663
rect 505 -3773 535 -3689
rect 600 -3773 700 -3643
rect 860 -3773 960 -3643
rect 1032 -3773 1062 -3689
rect 1314 -3773 1524 -3663
rect 1774 -3773 2352 -3663
rect 2602 -3773 2812 -3663
rect 3081 -3773 3111 -3689
rect 3176 -3773 3276 -3643
rect 3436 -3773 3536 -3643
rect 3608 -3773 3638 -3689
rect 3890 -3773 4100 -3663
rect 4350 -3773 4928 -3663
rect 5178 -3773 5388 -3663
rect 5657 -3773 5687 -3689
rect 5752 -3773 5852 -3643
rect 6012 -3773 6112 -3643
rect 6184 -3773 6214 -3689
rect 6466 -3773 6676 -3663
rect 6926 -3773 7504 -3663
rect 7754 -3773 7964 -3663
rect 8233 -3773 8263 -3689
rect 8328 -3773 8428 -3643
rect 8588 -3773 8688 -3643
rect 8760 -3773 8790 -3689
rect 9042 -3773 9252 -3663
rect 9502 -3773 10080 -3663
rect 10422 -3773 10632 -3663
rect 10809 -3773 10839 -3689
rect 10904 -3773 11004 -3643
rect 11164 -3773 11264 -3643
rect 11336 -3773 11366 -3689
rect 11710 -3773 11920 -3663
rect 13642 -3773 14588 -3663
rect 14838 -3773 15784 -3663
rect 16034 -3773 16612 -3663
rect -2918 -3977 -2340 -3867
rect -1538 -3977 -960 -3867
rect -802 -3977 -224 -3867
rect 26 -3977 236 -3867
rect 488 -3951 518 -3867
rect 590 -3997 690 -3867
rect 850 -3997 950 -3867
rect 1015 -3951 1045 -3867
rect 1314 -3977 1524 -3867
rect 1774 -3977 2352 -3867
rect 2602 -3977 2812 -3867
rect 3064 -3951 3094 -3867
rect 3166 -3997 3266 -3867
rect 3426 -3997 3526 -3867
rect 3591 -3951 3621 -3867
rect 3890 -3977 4100 -3867
rect 4350 -3977 4928 -3867
rect 5178 -3977 5388 -3867
rect 5640 -3951 5670 -3867
rect 5742 -3997 5842 -3867
rect 6002 -3997 6102 -3867
rect 6167 -3951 6197 -3867
rect 6466 -3977 6676 -3867
rect 6926 -3977 7504 -3867
rect 7754 -3977 7964 -3867
rect 8216 -3951 8246 -3867
rect 8318 -3997 8418 -3867
rect 8578 -3997 8678 -3867
rect 8743 -3951 8773 -3867
rect 9042 -3977 9252 -3867
rect 9502 -3977 10080 -3867
rect 10422 -3977 10632 -3867
rect 10792 -3951 10822 -3867
rect 10894 -3997 10994 -3867
rect 11154 -3997 11254 -3867
rect 11319 -3951 11349 -3867
rect 11710 -3977 11920 -3867
rect 12633 -3951 12663 -3867
rect 12719 -3951 12749 -3867
rect 12805 -3951 12835 -3867
rect 12891 -3951 12921 -3867
rect 13274 -3977 13484 -3867
rect 13735 -3951 13765 -3867
rect 13821 -3951 13851 -3867
rect 13907 -3951 13937 -3867
rect 13993 -3951 14023 -3867
rect 14079 -3951 14109 -3867
rect 14165 -3951 14195 -3867
rect 14251 -3951 14281 -3867
rect 14337 -3951 14367 -3867
rect 14423 -3951 14453 -3867
rect 14509 -3951 14539 -3867
rect 14595 -3951 14625 -3867
rect 14681 -3951 14711 -3867
rect 14766 -3951 14796 -3867
rect 14852 -3951 14882 -3867
rect 14938 -3951 14968 -3867
rect 15024 -3951 15054 -3867
rect 15110 -3951 15140 -3867
rect 15196 -3951 15226 -3867
rect 15282 -3951 15312 -3867
rect 15368 -3951 15398 -3867
rect 15666 -3977 16612 -3867
rect -2918 -4861 -2340 -4751
rect -1538 -4861 -960 -4751
rect -783 -4861 -753 -4777
rect -688 -4861 -588 -4731
rect -428 -4861 -328 -4731
rect -256 -4861 -226 -4777
rect 26 -4861 236 -4751
rect 505 -4861 535 -4777
rect 600 -4861 700 -4731
rect 860 -4861 960 -4731
rect 1032 -4861 1062 -4777
rect 1314 -4861 1524 -4751
rect 1774 -4861 2352 -4751
rect 2602 -4861 2812 -4751
rect 3081 -4861 3111 -4777
rect 3176 -4861 3276 -4731
rect 3436 -4861 3536 -4731
rect 3608 -4861 3638 -4777
rect 3890 -4861 4100 -4751
rect 4350 -4861 4928 -4751
rect 5178 -4861 5388 -4751
rect 5657 -4861 5687 -4777
rect 5752 -4861 5852 -4731
rect 6012 -4861 6112 -4731
rect 6184 -4861 6214 -4777
rect 6466 -4861 6676 -4751
rect 6926 -4861 7504 -4751
rect 7754 -4861 7964 -4751
rect 8233 -4861 8263 -4777
rect 8328 -4861 8428 -4731
rect 8588 -4861 8688 -4731
rect 8760 -4861 8790 -4777
rect 9042 -4861 9252 -4751
rect 9502 -4861 10080 -4751
rect 10422 -4861 10632 -4751
rect 10809 -4861 10839 -4777
rect 10904 -4861 11004 -4731
rect 11164 -4861 11264 -4731
rect 11336 -4861 11366 -4777
rect 11710 -4861 11920 -4751
rect 13735 -4861 13765 -4777
rect 13821 -4861 13851 -4777
rect 13907 -4861 13937 -4777
rect 13993 -4861 14023 -4777
rect 14079 -4861 14109 -4777
rect 14165 -4861 14195 -4777
rect 14251 -4861 14281 -4777
rect 14337 -4861 14367 -4777
rect 14423 -4861 14453 -4777
rect 14509 -4861 14539 -4777
rect 14595 -4861 14625 -4777
rect 14681 -4861 14711 -4777
rect 14766 -4861 14796 -4777
rect 14852 -4861 14882 -4777
rect 14938 -4861 14968 -4777
rect 15024 -4861 15054 -4777
rect 15110 -4861 15140 -4777
rect 15196 -4861 15226 -4777
rect 15282 -4861 15312 -4777
rect 15368 -4861 15398 -4777
rect 15666 -4861 16612 -4751
rect -2918 -5065 -2340 -4955
rect -1538 -5065 -960 -4955
rect -802 -5065 -224 -4955
rect 26 -5065 236 -4955
rect 488 -5039 518 -4955
rect 590 -5085 690 -4955
rect 850 -5085 950 -4955
rect 1015 -5039 1045 -4955
rect 1314 -5065 1524 -4955
rect 1774 -5065 2352 -4955
rect 2602 -5065 2812 -4955
rect 3064 -5039 3094 -4955
rect 3166 -5085 3266 -4955
rect 3426 -5085 3526 -4955
rect 3591 -5039 3621 -4955
rect 3890 -5065 4100 -4955
rect 4350 -5065 4928 -4955
rect 5178 -5065 5388 -4955
rect 5640 -5039 5670 -4955
rect 5742 -5085 5842 -4955
rect 6002 -5085 6102 -4955
rect 6167 -5039 6197 -4955
rect 6466 -5065 6676 -4955
rect 6926 -5065 7504 -4955
rect 7754 -5065 7964 -4955
rect 8216 -5039 8246 -4955
rect 8318 -5085 8418 -4955
rect 8578 -5085 8678 -4955
rect 8743 -5039 8773 -4955
rect 9042 -5065 9252 -4955
rect 9502 -5065 10080 -4955
rect 10422 -5065 10632 -4955
rect 10792 -5039 10822 -4955
rect 10894 -5085 10994 -4955
rect 11154 -5085 11254 -4955
rect 11319 -5039 11349 -4955
rect 11710 -5065 11920 -4955
rect 12633 -5039 12663 -4955
rect 12719 -5039 12749 -4955
rect 12805 -5039 12835 -4955
rect 12891 -5039 12921 -4955
rect 13274 -5065 13484 -4955
rect 13735 -5039 13765 -4955
rect 13821 -5039 13851 -4955
rect 13907 -5039 13937 -4955
rect 13993 -5039 14023 -4955
rect 14079 -5039 14109 -4955
rect 14165 -5039 14195 -4955
rect 14251 -5039 14281 -4955
rect 14337 -5039 14367 -4955
rect 14423 -5039 14453 -4955
rect 14509 -5039 14539 -4955
rect 14595 -5039 14625 -4955
rect 14681 -5039 14711 -4955
rect 14766 -5039 14796 -4955
rect 14852 -5039 14882 -4955
rect 14938 -5039 14968 -4955
rect 15024 -5039 15054 -4955
rect 15110 -5039 15140 -4955
rect 15196 -5039 15226 -4955
rect 15282 -5039 15312 -4955
rect 15368 -5039 15398 -4955
rect 15666 -5065 16612 -4955
rect -2918 -5949 -2340 -5839
rect -1538 -5949 -960 -5839
rect -802 -5949 -224 -5839
rect 26 -5949 236 -5839
rect 505 -5949 535 -5865
rect 600 -5949 700 -5819
rect 860 -5949 960 -5819
rect 1032 -5949 1062 -5865
rect 1314 -5949 1524 -5839
rect 1774 -5949 2352 -5839
rect 2602 -5949 2812 -5839
rect 3081 -5949 3111 -5865
rect 3176 -5949 3276 -5819
rect 3436 -5949 3536 -5819
rect 3608 -5949 3638 -5865
rect 3890 -5949 4100 -5839
rect 4350 -5949 4928 -5839
rect 5178 -5949 5388 -5839
rect 5657 -5949 5687 -5865
rect 5752 -5949 5852 -5819
rect 6012 -5949 6112 -5819
rect 6184 -5949 6214 -5865
rect 6466 -5949 6676 -5839
rect 6926 -5949 7504 -5839
rect 7754 -5949 7964 -5839
rect 8233 -5949 8263 -5865
rect 8328 -5949 8428 -5819
rect 8588 -5949 8688 -5819
rect 8760 -5949 8790 -5865
rect 9042 -5949 9252 -5839
rect 9502 -5949 10080 -5839
rect 10422 -5949 10632 -5839
rect 10809 -5949 10839 -5865
rect 10904 -5949 11004 -5819
rect 11164 -5949 11264 -5819
rect 11336 -5949 11366 -5865
rect 11710 -5949 11920 -5839
rect 13735 -5949 13765 -5865
rect 13821 -5949 13851 -5865
rect 13907 -5949 13937 -5865
rect 13993 -5949 14023 -5865
rect 14079 -5949 14109 -5865
rect 14165 -5949 14195 -5865
rect 14251 -5949 14281 -5865
rect 14337 -5949 14367 -5865
rect 14423 -5949 14453 -5865
rect 14509 -5949 14539 -5865
rect 14595 -5949 14625 -5865
rect 14681 -5949 14711 -5865
rect 14766 -5949 14796 -5865
rect 14852 -5949 14882 -5865
rect 14938 -5949 14968 -5865
rect 15024 -5949 15054 -5865
rect 15110 -5949 15140 -5865
rect 15196 -5949 15226 -5865
rect 15282 -5949 15312 -5865
rect 15368 -5949 15398 -5865
rect 15666 -5949 16612 -5839
rect -2918 -6153 -2340 -6043
rect -1354 -6153 -1144 -6043
rect -890 -6173 -860 -6043
rect -806 -6173 -776 -6043
rect -526 -6153 -316 -6043
rect 29 -6127 59 -6043
rect 115 -6127 145 -6043
rect 201 -6127 231 -6043
rect 287 -6127 317 -6043
rect 670 -6153 880 -6043
rect 1213 -6127 1243 -6043
rect 1498 -6153 1708 -6043
rect 1958 -6153 2168 -6043
rect 2420 -6127 2450 -6043
rect 2522 -6173 2622 -6043
rect 2782 -6173 2882 -6043
rect 2947 -6127 2977 -6043
rect 3246 -6153 3456 -6043
rect 4442 -6153 5388 -6043
rect 6466 -6153 6676 -6043
rect 6928 -6127 6958 -6043
rect 7030 -6173 7130 -6043
rect 7290 -6173 7390 -6043
rect 7455 -6127 7485 -6043
rect 7754 -6153 7964 -6043
rect 8216 -6127 8246 -6043
rect 8318 -6173 8418 -6043
rect 8578 -6173 8678 -6043
rect 8743 -6127 8773 -6043
rect 9042 -6153 9252 -6043
rect 9504 -6127 9534 -6043
rect 9606 -6173 9706 -6043
rect 9866 -6173 9966 -6043
rect 10031 -6127 10061 -6043
rect 10330 -6153 10540 -6043
rect 10790 -6173 10820 -6043
rect 10874 -6173 10904 -6043
rect 10958 -6173 10988 -6043
rect 11042 -6173 11072 -6043
rect 11126 -6173 11156 -6043
rect 11210 -6173 11240 -6043
rect 11294 -6173 11324 -6043
rect 11378 -6173 11408 -6043
rect 11710 -6153 11920 -6043
rect 13642 -6153 14588 -6043
rect 14838 -6153 15784 -6043
rect 16034 -6153 16612 -6043
rect -2918 -7037 -2800 -6927
rect -2550 -7037 -2520 -6953
rect -2466 -7037 -2436 -6953
rect -2278 -7037 -2248 -6953
rect -2166 -7037 -2136 -6965
rect -2067 -7037 -2037 -6965
rect -1968 -7037 -1938 -6953
rect -1849 -7037 -1819 -6909
rect -1748 -7037 -1718 -6965
rect -1642 -7037 -1612 -6965
rect -1547 -7037 -1517 -6953
rect -1357 -7037 -1327 -6907
rect -1273 -7037 -1243 -6907
rect -1085 -7037 -1055 -6953
rect -990 -7037 -960 -6907
rect -802 -7037 -224 -6927
rect 26 -7037 604 -6927
rect 762 -7037 1340 -6927
rect 1590 -7037 2168 -6927
rect 2326 -7037 2904 -6927
rect 3154 -7037 3732 -6927
rect 3890 -7037 4468 -6927
rect 4718 -7037 5296 -6927
rect 5454 -7037 6032 -6927
rect 6282 -7037 6860 -6927
rect 7018 -7037 7596 -6927
rect 7846 -7037 8424 -6927
rect 8582 -7037 9160 -6927
rect 16034 -7037 16612 -6927
rect -2918 -7241 -2340 -7131
rect -1538 -7241 -960 -7131
rect -802 -7241 -224 -7131
rect 26 -7241 604 -7131
rect 762 -7241 1340 -7131
rect 1590 -7241 2168 -7131
rect 2326 -7241 2536 -7131
rect 2975 -7215 3005 -7131
rect 3338 -7241 3548 -7131
rect 3802 -7261 3832 -7131
rect 3886 -7261 3916 -7131
rect 4166 -7241 4376 -7131
rect 4626 -7261 4656 -7131
rect 4735 -7215 4765 -7131
rect 4831 -7215 4861 -7131
rect 4956 -7215 4986 -7131
rect 5052 -7215 5082 -7131
rect 5220 -7215 5250 -7131
rect 5546 -7241 5756 -7131
rect 6006 -7261 6036 -7131
rect 6101 -7215 6131 -7131
rect 6289 -7261 6319 -7131
rect 6373 -7261 6403 -7131
rect 6563 -7215 6593 -7131
rect 6658 -7203 6688 -7131
rect 6764 -7203 6794 -7131
rect 6865 -7259 6895 -7131
rect 6984 -7215 7014 -7131
rect 7083 -7203 7113 -7131
rect 7182 -7203 7212 -7131
rect 7294 -7215 7324 -7131
rect 7482 -7215 7512 -7131
rect 7566 -7215 7596 -7131
rect 7846 -7241 8424 -7131
rect 8582 -7241 9160 -7131
rect 16034 -7241 16612 -7131
rect -2918 -8125 -2340 -8015
rect -1354 -8125 -1144 -8015
rect -890 -8125 -860 -7995
rect -806 -8125 -776 -7995
rect -526 -8125 -316 -8015
rect 29 -8125 59 -8041
rect 115 -8125 145 -8041
rect 201 -8125 231 -8041
rect 287 -8125 317 -8041
rect 670 -8125 880 -8015
rect 1213 -8125 1243 -8041
rect 1498 -8125 1708 -8015
rect 1958 -8125 2168 -8015
rect 2420 -8125 2450 -8041
rect 2522 -8125 2622 -7995
rect 2782 -8125 2882 -7995
rect 2947 -8125 2977 -8041
rect 3246 -8125 3456 -8015
rect 4442 -8125 5388 -8015
rect 6466 -8125 6676 -8015
rect 6928 -8125 6958 -8041
rect 7030 -8125 7130 -7995
rect 7290 -8125 7390 -7995
rect 7455 -8125 7485 -8041
rect 7754 -8125 7964 -8015
rect 8216 -8125 8246 -8041
rect 8318 -8125 8418 -7995
rect 8578 -8125 8678 -7995
rect 8743 -8125 8773 -8041
rect 9042 -8125 9252 -8015
rect 9504 -8125 9534 -8041
rect 9606 -8125 9706 -7995
rect 9866 -8125 9966 -7995
rect 10031 -8125 10061 -8041
rect 10330 -8125 10540 -8015
rect 10790 -8125 10820 -7995
rect 10874 -8125 10904 -7995
rect 10958 -8125 10988 -7995
rect 11042 -8125 11072 -7995
rect 11126 -8125 11156 -7995
rect 11210 -8125 11240 -7995
rect 11294 -8125 11324 -7995
rect 11378 -8125 11408 -7995
rect 11710 -8125 11920 -8015
rect 13642 -8125 14588 -8015
rect 14838 -8125 15784 -8015
rect 16034 -8125 16612 -8015
rect -2918 -8329 -2340 -8219
rect -1538 -8329 -960 -8219
rect -802 -8329 -224 -8219
rect 26 -8329 236 -8219
rect 505 -8303 535 -8219
rect 600 -8349 700 -8219
rect 860 -8349 960 -8219
rect 1032 -8303 1062 -8219
rect 1314 -8329 1524 -8219
rect 1774 -8329 2352 -8219
rect 2602 -8329 2812 -8219
rect 3081 -8303 3111 -8219
rect 3176 -8349 3276 -8219
rect 3436 -8349 3536 -8219
rect 3608 -8303 3638 -8219
rect 3890 -8329 4100 -8219
rect 4350 -8329 4928 -8219
rect 5178 -8329 5388 -8219
rect 5657 -8303 5687 -8219
rect 5752 -8349 5852 -8219
rect 6012 -8349 6112 -8219
rect 6184 -8303 6214 -8219
rect 6466 -8329 6676 -8219
rect 6926 -8329 7504 -8219
rect 7754 -8329 7964 -8219
rect 8233 -8303 8263 -8219
rect 8328 -8349 8428 -8219
rect 8588 -8349 8688 -8219
rect 8760 -8303 8790 -8219
rect 9042 -8329 9252 -8219
rect 9502 -8329 10080 -8219
rect 10422 -8329 10632 -8219
rect 10809 -8303 10839 -8219
rect 10904 -8349 11004 -8219
rect 11164 -8349 11264 -8219
rect 11336 -8303 11366 -8219
rect 11710 -8329 11920 -8219
rect 13735 -8303 13765 -8219
rect 13821 -8303 13851 -8219
rect 13907 -8303 13937 -8219
rect 13993 -8303 14023 -8219
rect 14079 -8303 14109 -8219
rect 14165 -8303 14195 -8219
rect 14251 -8303 14281 -8219
rect 14337 -8303 14367 -8219
rect 14423 -8303 14453 -8219
rect 14509 -8303 14539 -8219
rect 14595 -8303 14625 -8219
rect 14681 -8303 14711 -8219
rect 14766 -8303 14796 -8219
rect 14852 -8303 14882 -8219
rect 14938 -8303 14968 -8219
rect 15024 -8303 15054 -8219
rect 15110 -8303 15140 -8219
rect 15196 -8303 15226 -8219
rect 15282 -8303 15312 -8219
rect 15368 -8303 15398 -8219
rect 15666 -8329 16612 -8219
rect -2918 -9213 -2340 -9103
rect -1538 -9213 -960 -9103
rect -802 -9213 -224 -9103
rect 26 -9213 236 -9103
rect 488 -9213 518 -9129
rect 590 -9213 690 -9083
rect 850 -9213 950 -9083
rect 1015 -9213 1045 -9129
rect 1314 -9213 1524 -9103
rect 1774 -9213 2352 -9103
rect 2602 -9213 2812 -9103
rect 3064 -9213 3094 -9129
rect 3166 -9213 3266 -9083
rect 3426 -9213 3526 -9083
rect 3591 -9213 3621 -9129
rect 3890 -9213 4100 -9103
rect 4350 -9213 4928 -9103
rect 5178 -9213 5388 -9103
rect 5640 -9213 5670 -9129
rect 5742 -9213 5842 -9083
rect 6002 -9213 6102 -9083
rect 6167 -9213 6197 -9129
rect 6466 -9213 6676 -9103
rect 6926 -9213 7504 -9103
rect 7754 -9213 7964 -9103
rect 8216 -9213 8246 -9129
rect 8318 -9213 8418 -9083
rect 8578 -9213 8678 -9083
rect 8743 -9213 8773 -9129
rect 9042 -9213 9252 -9103
rect 9502 -9213 10080 -9103
rect 10422 -9213 10632 -9103
rect 10792 -9213 10822 -9129
rect 10894 -9213 10994 -9083
rect 11154 -9213 11254 -9083
rect 11319 -9213 11349 -9129
rect 11710 -9213 11920 -9103
rect 12633 -9213 12663 -9129
rect 12719 -9213 12749 -9129
rect 12805 -9213 12835 -9129
rect 12891 -9213 12921 -9129
rect 13274 -9213 13484 -9103
rect 13735 -9213 13765 -9129
rect 13821 -9213 13851 -9129
rect 13907 -9213 13937 -9129
rect 13993 -9213 14023 -9129
rect 14079 -9213 14109 -9129
rect 14165 -9213 14195 -9129
rect 14251 -9213 14281 -9129
rect 14337 -9213 14367 -9129
rect 14423 -9213 14453 -9129
rect 14509 -9213 14539 -9129
rect 14595 -9213 14625 -9129
rect 14681 -9213 14711 -9129
rect 14766 -9213 14796 -9129
rect 14852 -9213 14882 -9129
rect 14938 -9213 14968 -9129
rect 15024 -9213 15054 -9129
rect 15110 -9213 15140 -9129
rect 15196 -9213 15226 -9129
rect 15282 -9213 15312 -9129
rect 15368 -9213 15398 -9129
rect 15666 -9213 16612 -9103
rect -2918 -9417 -2340 -9307
rect -1538 -9417 -960 -9307
rect -783 -9391 -753 -9307
rect -688 -9437 -588 -9307
rect -428 -9437 -328 -9307
rect -256 -9391 -226 -9307
rect 26 -9417 236 -9307
rect 505 -9391 535 -9307
rect 600 -9437 700 -9307
rect 860 -9437 960 -9307
rect 1032 -9391 1062 -9307
rect 1314 -9417 1524 -9307
rect 1774 -9417 2352 -9307
rect 2602 -9417 2812 -9307
rect 3081 -9391 3111 -9307
rect 3176 -9437 3276 -9307
rect 3436 -9437 3536 -9307
rect 3608 -9391 3638 -9307
rect 3890 -9417 4100 -9307
rect 4350 -9417 4928 -9307
rect 5178 -9417 5388 -9307
rect 5657 -9391 5687 -9307
rect 5752 -9437 5852 -9307
rect 6012 -9437 6112 -9307
rect 6184 -9391 6214 -9307
rect 6466 -9417 6676 -9307
rect 6926 -9417 7504 -9307
rect 7754 -9417 7964 -9307
rect 8233 -9391 8263 -9307
rect 8328 -9437 8428 -9307
rect 8588 -9437 8688 -9307
rect 8760 -9391 8790 -9307
rect 9042 -9417 9252 -9307
rect 9502 -9417 10080 -9307
rect 10422 -9417 10632 -9307
rect 10809 -9391 10839 -9307
rect 10904 -9437 11004 -9307
rect 11164 -9437 11264 -9307
rect 11336 -9391 11366 -9307
rect 11710 -9417 11920 -9307
rect 13735 -9391 13765 -9307
rect 13821 -9391 13851 -9307
rect 13907 -9391 13937 -9307
rect 13993 -9391 14023 -9307
rect 14079 -9391 14109 -9307
rect 14165 -9391 14195 -9307
rect 14251 -9391 14281 -9307
rect 14337 -9391 14367 -9307
rect 14423 -9391 14453 -9307
rect 14509 -9391 14539 -9307
rect 14595 -9391 14625 -9307
rect 14681 -9391 14711 -9307
rect 14766 -9391 14796 -9307
rect 14852 -9391 14882 -9307
rect 14938 -9391 14968 -9307
rect 15024 -9391 15054 -9307
rect 15110 -9391 15140 -9307
rect 15196 -9391 15226 -9307
rect 15282 -9391 15312 -9307
rect 15368 -9391 15398 -9307
rect 15666 -9417 16612 -9307
rect -2918 -10301 -2340 -10191
rect -1538 -10301 -960 -10191
rect -802 -10301 -224 -10191
rect 26 -10301 236 -10191
rect 488 -10301 518 -10217
rect 590 -10301 690 -10171
rect 850 -10301 950 -10171
rect 1015 -10301 1045 -10217
rect 1314 -10301 1524 -10191
rect 1774 -10301 2352 -10191
rect 2602 -10301 2812 -10191
rect 3064 -10301 3094 -10217
rect 3166 -10301 3266 -10171
rect 3426 -10301 3526 -10171
rect 3591 -10301 3621 -10217
rect 3890 -10301 4100 -10191
rect 4350 -10301 4928 -10191
rect 5178 -10301 5388 -10191
rect 5640 -10301 5670 -10217
rect 5742 -10301 5842 -10171
rect 6002 -10301 6102 -10171
rect 6167 -10301 6197 -10217
rect 6466 -10301 6676 -10191
rect 6926 -10301 7504 -10191
rect 7754 -10301 7964 -10191
rect 8216 -10301 8246 -10217
rect 8318 -10301 8418 -10171
rect 8578 -10301 8678 -10171
rect 8743 -10301 8773 -10217
rect 9042 -10301 9252 -10191
rect 9502 -10301 10080 -10191
rect 10422 -10301 10632 -10191
rect 10792 -10301 10822 -10217
rect 10894 -10301 10994 -10171
rect 11154 -10301 11254 -10171
rect 11319 -10301 11349 -10217
rect 11710 -10301 11920 -10191
rect 12633 -10301 12663 -10217
rect 12719 -10301 12749 -10217
rect 12805 -10301 12835 -10217
rect 12891 -10301 12921 -10217
rect 13274 -10301 13484 -10191
rect 13735 -10301 13765 -10217
rect 13821 -10301 13851 -10217
rect 13907 -10301 13937 -10217
rect 13993 -10301 14023 -10217
rect 14079 -10301 14109 -10217
rect 14165 -10301 14195 -10217
rect 14251 -10301 14281 -10217
rect 14337 -10301 14367 -10217
rect 14423 -10301 14453 -10217
rect 14509 -10301 14539 -10217
rect 14595 -10301 14625 -10217
rect 14681 -10301 14711 -10217
rect 14766 -10301 14796 -10217
rect 14852 -10301 14882 -10217
rect 14938 -10301 14968 -10217
rect 15024 -10301 15054 -10217
rect 15110 -10301 15140 -10217
rect 15196 -10301 15226 -10217
rect 15282 -10301 15312 -10217
rect 15368 -10301 15398 -10217
rect 15666 -10301 16612 -10191
rect -2918 -10505 -2340 -10395
rect -1823 -10479 -1793 -10395
rect -1538 -10505 -960 -10395
rect -802 -10505 -224 -10395
rect 26 -10505 236 -10395
rect 505 -10479 535 -10395
rect 600 -10525 700 -10395
rect 860 -10525 960 -10395
rect 1032 -10479 1062 -10395
rect 1314 -10505 1524 -10395
rect 1774 -10505 2352 -10395
rect 2602 -10505 2812 -10395
rect 3081 -10479 3111 -10395
rect 3176 -10525 3276 -10395
rect 3436 -10525 3536 -10395
rect 3608 -10479 3638 -10395
rect 3890 -10505 4100 -10395
rect 4350 -10505 4928 -10395
rect 5178 -10505 5388 -10395
rect 5657 -10479 5687 -10395
rect 5752 -10525 5852 -10395
rect 6012 -10525 6112 -10395
rect 6184 -10479 6214 -10395
rect 6466 -10505 6676 -10395
rect 6926 -10505 7504 -10395
rect 7754 -10505 7964 -10395
rect 8233 -10479 8263 -10395
rect 8328 -10525 8428 -10395
rect 8588 -10525 8688 -10395
rect 8760 -10479 8790 -10395
rect 9042 -10505 9252 -10395
rect 9502 -10505 10080 -10395
rect 10422 -10505 10632 -10395
rect 10809 -10479 10839 -10395
rect 10904 -10525 11004 -10395
rect 11164 -10525 11264 -10395
rect 11336 -10479 11366 -10395
rect 11710 -10505 11920 -10395
rect 13642 -10505 14588 -10395
rect 14838 -10505 15784 -10395
rect 16034 -10505 16612 -10395
rect -2918 -11389 -2340 -11279
rect -1538 -11389 -960 -11279
rect -802 -11389 -224 -11279
rect 26 -11389 236 -11279
rect 505 -11389 535 -11305
rect 600 -11389 700 -11259
rect 860 -11389 960 -11259
rect 1032 -11389 1062 -11305
rect 1314 -11389 1524 -11279
rect 1774 -11389 2352 -11279
rect 2602 -11389 2812 -11279
rect 3081 -11389 3111 -11305
rect 3176 -11389 3276 -11259
rect 3436 -11389 3536 -11259
rect 3608 -11389 3638 -11305
rect 3890 -11389 4100 -11279
rect 4350 -11389 4928 -11279
rect 5178 -11389 5388 -11279
rect 5657 -11389 5687 -11305
rect 5752 -11389 5852 -11259
rect 6012 -11389 6112 -11259
rect 6184 -11389 6214 -11305
rect 6466 -11389 6676 -11279
rect 6926 -11389 7504 -11279
rect 7754 -11389 7964 -11279
rect 8233 -11389 8263 -11305
rect 8328 -11389 8428 -11259
rect 8588 -11389 8688 -11259
rect 8760 -11389 8790 -11305
rect 9042 -11389 9252 -11279
rect 9502 -11389 10080 -11279
rect 10422 -11389 10632 -11279
rect 10809 -11389 10839 -11305
rect 10904 -11389 11004 -11259
rect 11164 -11389 11264 -11259
rect 11336 -11389 11366 -11305
rect 11710 -11389 11920 -11279
rect 13642 -11389 14588 -11279
rect 14838 -11389 15784 -11279
rect 16034 -11389 16612 -11279
rect -2918 -11593 -2340 -11483
rect -1538 -11593 -960 -11483
rect -802 -11593 -224 -11483
rect 26 -11593 236 -11483
rect 488 -11567 518 -11483
rect 590 -11613 690 -11483
rect 850 -11613 950 -11483
rect 1015 -11567 1045 -11483
rect 1314 -11593 1524 -11483
rect 1774 -11593 2352 -11483
rect 2602 -11593 2812 -11483
rect 3064 -11567 3094 -11483
rect 3166 -11613 3266 -11483
rect 3426 -11613 3526 -11483
rect 3591 -11567 3621 -11483
rect 3890 -11593 4100 -11483
rect 4350 -11593 4928 -11483
rect 5178 -11593 5388 -11483
rect 5640 -11567 5670 -11483
rect 5742 -11613 5842 -11483
rect 6002 -11613 6102 -11483
rect 6167 -11567 6197 -11483
rect 6466 -11593 6676 -11483
rect 6926 -11593 7504 -11483
rect 7754 -11593 7964 -11483
rect 8216 -11567 8246 -11483
rect 8318 -11613 8418 -11483
rect 8578 -11613 8678 -11483
rect 8743 -11567 8773 -11483
rect 9042 -11593 9252 -11483
rect 9502 -11593 10080 -11483
rect 10422 -11593 10632 -11483
rect 10792 -11567 10822 -11483
rect 10894 -11613 10994 -11483
rect 11154 -11613 11254 -11483
rect 11319 -11567 11349 -11483
rect 11710 -11593 11920 -11483
rect 12633 -11567 12663 -11483
rect 12719 -11567 12749 -11483
rect 12805 -11567 12835 -11483
rect 12891 -11567 12921 -11483
rect 13274 -11593 13484 -11483
rect 13735 -11567 13765 -11483
rect 13821 -11567 13851 -11483
rect 13907 -11567 13937 -11483
rect 13993 -11567 14023 -11483
rect 14079 -11567 14109 -11483
rect 14165 -11567 14195 -11483
rect 14251 -11567 14281 -11483
rect 14337 -11567 14367 -11483
rect 14423 -11567 14453 -11483
rect 14509 -11567 14539 -11483
rect 14595 -11567 14625 -11483
rect 14681 -11567 14711 -11483
rect 14766 -11567 14796 -11483
rect 14852 -11567 14882 -11483
rect 14938 -11567 14968 -11483
rect 15024 -11567 15054 -11483
rect 15110 -11567 15140 -11483
rect 15196 -11567 15226 -11483
rect 15282 -11567 15312 -11483
rect 15368 -11567 15398 -11483
rect 15666 -11593 16612 -11483
rect -2918 -12477 -2340 -12367
rect -1538 -12477 -960 -12367
rect -783 -12477 -753 -12393
rect -688 -12477 -588 -12347
rect -428 -12477 -328 -12347
rect -256 -12477 -226 -12393
rect 26 -12477 236 -12367
rect 505 -12477 535 -12393
rect 600 -12477 700 -12347
rect 860 -12477 960 -12347
rect 1032 -12477 1062 -12393
rect 1314 -12477 1524 -12367
rect 1774 -12477 2352 -12367
rect 2602 -12477 2812 -12367
rect 3081 -12477 3111 -12393
rect 3176 -12477 3276 -12347
rect 3436 -12477 3536 -12347
rect 3608 -12477 3638 -12393
rect 3890 -12477 4100 -12367
rect 4350 -12477 4928 -12367
rect 5178 -12477 5388 -12367
rect 5657 -12477 5687 -12393
rect 5752 -12477 5852 -12347
rect 6012 -12477 6112 -12347
rect 6184 -12477 6214 -12393
rect 6466 -12477 6676 -12367
rect 6926 -12477 7504 -12367
rect 7754 -12477 7964 -12367
rect 8233 -12477 8263 -12393
rect 8328 -12477 8428 -12347
rect 8588 -12477 8688 -12347
rect 8760 -12477 8790 -12393
rect 9042 -12477 9252 -12367
rect 9502 -12477 10080 -12367
rect 10422 -12477 10632 -12367
rect 10809 -12477 10839 -12393
rect 10904 -12477 11004 -12347
rect 11164 -12477 11264 -12347
rect 11336 -12477 11366 -12393
rect 11710 -12477 11920 -12367
rect 13735 -12477 13765 -12393
rect 13821 -12477 13851 -12393
rect 13907 -12477 13937 -12393
rect 13993 -12477 14023 -12393
rect 14079 -12477 14109 -12393
rect 14165 -12477 14195 -12393
rect 14251 -12477 14281 -12393
rect 14337 -12477 14367 -12393
rect 14423 -12477 14453 -12393
rect 14509 -12477 14539 -12393
rect 14595 -12477 14625 -12393
rect 14681 -12477 14711 -12393
rect 14766 -12477 14796 -12393
rect 14852 -12477 14882 -12393
rect 14938 -12477 14968 -12393
rect 15024 -12477 15054 -12393
rect 15110 -12477 15140 -12393
rect 15196 -12477 15226 -12393
rect 15282 -12477 15312 -12393
rect 15368 -12477 15398 -12393
rect 15666 -12477 16612 -12367
rect -2918 -12681 -2340 -12571
rect -1538 -12681 -960 -12571
rect -802 -12681 -224 -12571
rect 26 -12681 236 -12571
rect 488 -12655 518 -12571
rect 590 -12701 690 -12571
rect 850 -12701 950 -12571
rect 1015 -12655 1045 -12571
rect 1314 -12681 1524 -12571
rect 1774 -12681 2352 -12571
rect 2602 -12681 2812 -12571
rect 3064 -12655 3094 -12571
rect 3166 -12701 3266 -12571
rect 3426 -12701 3526 -12571
rect 3591 -12655 3621 -12571
rect 3890 -12681 4100 -12571
rect 4350 -12681 4928 -12571
rect 5178 -12681 5388 -12571
rect 5640 -12655 5670 -12571
rect 5742 -12701 5842 -12571
rect 6002 -12701 6102 -12571
rect 6167 -12655 6197 -12571
rect 6466 -12681 6676 -12571
rect 6926 -12681 7504 -12571
rect 7754 -12681 7964 -12571
rect 8216 -12655 8246 -12571
rect 8318 -12701 8418 -12571
rect 8578 -12701 8678 -12571
rect 8743 -12655 8773 -12571
rect 9042 -12681 9252 -12571
rect 9502 -12681 10080 -12571
rect 10422 -12681 10632 -12571
rect 10792 -12655 10822 -12571
rect 10894 -12701 10994 -12571
rect 11154 -12701 11254 -12571
rect 11319 -12655 11349 -12571
rect 11710 -12681 11920 -12571
rect 12633 -12655 12663 -12571
rect 12719 -12655 12749 -12571
rect 12805 -12655 12835 -12571
rect 12891 -12655 12921 -12571
rect 13274 -12681 13484 -12571
rect 13735 -12655 13765 -12571
rect 13821 -12655 13851 -12571
rect 13907 -12655 13937 -12571
rect 13993 -12655 14023 -12571
rect 14079 -12655 14109 -12571
rect 14165 -12655 14195 -12571
rect 14251 -12655 14281 -12571
rect 14337 -12655 14367 -12571
rect 14423 -12655 14453 -12571
rect 14509 -12655 14539 -12571
rect 14595 -12655 14625 -12571
rect 14681 -12655 14711 -12571
rect 14766 -12655 14796 -12571
rect 14852 -12655 14882 -12571
rect 14938 -12655 14968 -12571
rect 15024 -12655 15054 -12571
rect 15110 -12655 15140 -12571
rect 15196 -12655 15226 -12571
rect 15282 -12655 15312 -12571
rect 15368 -12655 15398 -12571
rect 15666 -12681 16612 -12571
rect -2918 -13565 -2340 -13455
rect -1538 -13565 -960 -13455
rect -802 -13565 -224 -13455
rect 26 -13565 236 -13455
rect 505 -13565 535 -13481
rect 600 -13565 700 -13435
rect 860 -13565 960 -13435
rect 1032 -13565 1062 -13481
rect 1314 -13565 1524 -13455
rect 1774 -13565 2352 -13455
rect 2602 -13565 2812 -13455
rect 3081 -13565 3111 -13481
rect 3176 -13565 3276 -13435
rect 3436 -13565 3536 -13435
rect 3608 -13565 3638 -13481
rect 3890 -13565 4100 -13455
rect 4350 -13565 4928 -13455
rect 5178 -13565 5388 -13455
rect 5657 -13565 5687 -13481
rect 5752 -13565 5852 -13435
rect 6012 -13565 6112 -13435
rect 6184 -13565 6214 -13481
rect 6466 -13565 6676 -13455
rect 6926 -13565 7504 -13455
rect 7754 -13565 7964 -13455
rect 8233 -13565 8263 -13481
rect 8328 -13565 8428 -13435
rect 8588 -13565 8688 -13435
rect 8760 -13565 8790 -13481
rect 9042 -13565 9252 -13455
rect 9502 -13565 10080 -13455
rect 10422 -13565 10632 -13455
rect 10809 -13565 10839 -13481
rect 10904 -13565 11004 -13435
rect 11164 -13565 11264 -13435
rect 11336 -13565 11366 -13481
rect 11710 -13565 11920 -13455
rect 13735 -13565 13765 -13481
rect 13821 -13565 13851 -13481
rect 13907 -13565 13937 -13481
rect 13993 -13565 14023 -13481
rect 14079 -13565 14109 -13481
rect 14165 -13565 14195 -13481
rect 14251 -13565 14281 -13481
rect 14337 -13565 14367 -13481
rect 14423 -13565 14453 -13481
rect 14509 -13565 14539 -13481
rect 14595 -13565 14625 -13481
rect 14681 -13565 14711 -13481
rect 14766 -13565 14796 -13481
rect 14852 -13565 14882 -13481
rect 14938 -13565 14968 -13481
rect 15024 -13565 15054 -13481
rect 15110 -13565 15140 -13481
rect 15196 -13565 15226 -13481
rect 15282 -13565 15312 -13481
rect 15368 -13565 15398 -13481
rect 15666 -13565 16612 -13455
rect -2918 -13769 -2340 -13659
rect -1354 -13769 -1144 -13659
rect -890 -13789 -860 -13659
rect -806 -13789 -776 -13659
rect -526 -13769 -316 -13659
rect 29 -13743 59 -13659
rect 115 -13743 145 -13659
rect 201 -13743 231 -13659
rect 287 -13743 317 -13659
rect 670 -13769 880 -13659
rect 1213 -13743 1243 -13659
rect 1498 -13769 1708 -13659
rect 1958 -13769 2168 -13659
rect 2420 -13743 2450 -13659
rect 2522 -13789 2622 -13659
rect 2782 -13789 2882 -13659
rect 2947 -13743 2977 -13659
rect 3246 -13769 3456 -13659
rect 4442 -13769 5388 -13659
rect 6466 -13769 6676 -13659
rect 6928 -13743 6958 -13659
rect 7030 -13789 7130 -13659
rect 7290 -13789 7390 -13659
rect 7455 -13743 7485 -13659
rect 7754 -13769 7964 -13659
rect 8216 -13743 8246 -13659
rect 8318 -13789 8418 -13659
rect 8578 -13789 8678 -13659
rect 8743 -13743 8773 -13659
rect 9042 -13769 9252 -13659
rect 9504 -13743 9534 -13659
rect 9606 -13789 9706 -13659
rect 9866 -13789 9966 -13659
rect 10031 -13743 10061 -13659
rect 10330 -13769 10540 -13659
rect 10790 -13789 10820 -13659
rect 10874 -13789 10904 -13659
rect 10958 -13789 10988 -13659
rect 11042 -13789 11072 -13659
rect 11126 -13789 11156 -13659
rect 11210 -13789 11240 -13659
rect 11294 -13789 11324 -13659
rect 11378 -13789 11408 -13659
rect 11710 -13769 11920 -13659
rect 13642 -13769 14588 -13659
rect 14838 -13769 15784 -13659
rect 16034 -13769 16612 -13659
<< scpmoshvt >>
rect -2918 -233 -2340 -59
rect -1354 -233 -1144 -59
rect -890 -259 -860 -59
rect -806 -259 -776 -59
rect -526 -233 -316 -59
rect -57 -259 -27 -59
rect 29 -259 59 -59
rect 115 -259 145 -59
rect 201 -259 231 -59
rect 287 -259 317 -59
rect 373 -259 403 -59
rect 670 -233 880 -59
rect 1130 -227 1160 -59
rect 1214 -227 1244 -59
rect 1498 -233 1708 -59
rect 1958 -233 2168 -59
rect 2420 -259 2450 -59
rect 2522 -223 2622 -59
rect 2782 -223 2882 -59
rect 2947 -259 2977 -59
rect 3246 -233 3456 -59
rect 4442 -233 5388 -59
rect 6466 -233 6676 -59
rect 6928 -259 6958 -59
rect 7030 -223 7130 -59
rect 7290 -223 7390 -59
rect 7455 -259 7485 -59
rect 7754 -233 7964 -59
rect 8216 -259 8246 -59
rect 8318 -223 8418 -59
rect 8578 -223 8678 -59
rect 8743 -259 8773 -59
rect 9042 -233 9252 -59
rect 9504 -259 9534 -59
rect 9606 -223 9706 -59
rect 9866 -223 9966 -59
rect 10031 -259 10061 -59
rect 10330 -233 10540 -59
rect 10790 -259 10820 -59
rect 10874 -259 10904 -59
rect 10958 -259 10988 -59
rect 11042 -259 11072 -59
rect 11126 -259 11156 -59
rect 11210 -259 11240 -59
rect 11294 -259 11324 -59
rect 11378 -259 11408 -59
rect 11710 -233 11920 -59
rect 13642 -233 14588 -59
rect 14838 -233 15784 -59
rect 16034 -233 16612 -59
rect -2918 -1053 -2340 -879
rect -1538 -1053 -960 -879
rect -802 -1053 -224 -879
rect 26 -1053 236 -879
rect 505 -1053 535 -853
rect 600 -1053 700 -889
rect 860 -1053 960 -889
rect 1032 -1053 1062 -853
rect 1314 -1053 1524 -879
rect 1774 -1053 2352 -879
rect 2602 -1053 2812 -879
rect 3081 -1053 3111 -853
rect 3176 -1053 3276 -889
rect 3436 -1053 3536 -889
rect 3608 -1053 3638 -853
rect 3890 -1053 4100 -879
rect 4350 -1053 4928 -879
rect 5178 -1053 5388 -879
rect 5657 -1053 5687 -853
rect 5752 -1053 5852 -889
rect 6012 -1053 6112 -889
rect 6184 -1053 6214 -853
rect 6466 -1053 6676 -879
rect 6926 -1053 7504 -879
rect 7754 -1053 7964 -879
rect 8233 -1053 8263 -853
rect 8328 -1053 8428 -889
rect 8588 -1053 8688 -889
rect 8760 -1053 8790 -853
rect 9042 -1053 9252 -879
rect 9502 -1053 10080 -879
rect 10422 -1053 10632 -879
rect 10809 -1053 10839 -853
rect 10904 -1053 11004 -889
rect 11164 -1053 11264 -889
rect 11336 -1053 11366 -853
rect 11710 -1053 11920 -879
rect 13735 -1053 13765 -853
rect 13821 -1053 13851 -853
rect 13907 -1053 13937 -853
rect 13993 -1053 14023 -853
rect 14079 -1053 14109 -853
rect 14165 -1053 14195 -853
rect 14251 -1053 14281 -853
rect 14337 -1053 14367 -853
rect 14423 -1053 14453 -853
rect 14509 -1053 14539 -853
rect 14595 -1053 14625 -853
rect 14681 -1053 14711 -853
rect 14766 -1053 14796 -853
rect 14852 -1053 14882 -853
rect 14938 -1053 14968 -853
rect 15024 -1053 15054 -853
rect 15110 -1053 15140 -853
rect 15196 -1053 15226 -853
rect 15282 -1053 15312 -853
rect 15368 -1053 15398 -853
rect 15666 -1053 16612 -879
rect -2918 -1321 -2340 -1147
rect -1538 -1321 -960 -1147
rect -802 -1321 -224 -1147
rect 26 -1321 236 -1147
rect 488 -1347 518 -1147
rect 590 -1311 690 -1147
rect 850 -1311 950 -1147
rect 1015 -1347 1045 -1147
rect 1314 -1321 1524 -1147
rect 1774 -1321 2352 -1147
rect 2602 -1321 2812 -1147
rect 3064 -1347 3094 -1147
rect 3166 -1311 3266 -1147
rect 3426 -1311 3526 -1147
rect 3591 -1347 3621 -1147
rect 3890 -1321 4100 -1147
rect 4350 -1321 4928 -1147
rect 5178 -1321 5388 -1147
rect 5640 -1347 5670 -1147
rect 5742 -1311 5842 -1147
rect 6002 -1311 6102 -1147
rect 6167 -1347 6197 -1147
rect 6466 -1321 6676 -1147
rect 6926 -1321 7504 -1147
rect 7754 -1321 7964 -1147
rect 8216 -1347 8246 -1147
rect 8318 -1311 8418 -1147
rect 8578 -1311 8678 -1147
rect 8743 -1347 8773 -1147
rect 9042 -1321 9252 -1147
rect 9502 -1321 10080 -1147
rect 10422 -1321 10632 -1147
rect 10792 -1347 10822 -1147
rect 10894 -1311 10994 -1147
rect 11154 -1311 11254 -1147
rect 11319 -1347 11349 -1147
rect 11710 -1321 11920 -1147
rect 12547 -1347 12577 -1147
rect 12633 -1347 12663 -1147
rect 12719 -1347 12749 -1147
rect 12805 -1347 12835 -1147
rect 12891 -1347 12921 -1147
rect 12977 -1347 13007 -1147
rect 13274 -1321 13484 -1147
rect 13735 -1347 13765 -1147
rect 13821 -1347 13851 -1147
rect 13907 -1347 13937 -1147
rect 13993 -1347 14023 -1147
rect 14079 -1347 14109 -1147
rect 14165 -1347 14195 -1147
rect 14251 -1347 14281 -1147
rect 14337 -1347 14367 -1147
rect 14423 -1347 14453 -1147
rect 14509 -1347 14539 -1147
rect 14595 -1347 14625 -1147
rect 14681 -1347 14711 -1147
rect 14766 -1347 14796 -1147
rect 14852 -1347 14882 -1147
rect 14938 -1347 14968 -1147
rect 15024 -1347 15054 -1147
rect 15110 -1347 15140 -1147
rect 15196 -1347 15226 -1147
rect 15282 -1347 15312 -1147
rect 15368 -1347 15398 -1147
rect 15666 -1321 16612 -1147
rect -2918 -2141 -2340 -1967
rect -1538 -2141 -960 -1967
rect -783 -2141 -753 -1941
rect -688 -2141 -588 -1977
rect -428 -2141 -328 -1977
rect -256 -2141 -226 -1941
rect 26 -2141 236 -1967
rect 505 -2141 535 -1941
rect 600 -2141 700 -1977
rect 860 -2141 960 -1977
rect 1032 -2141 1062 -1941
rect 1314 -2141 1524 -1967
rect 1774 -2141 2352 -1967
rect 2602 -2141 2812 -1967
rect 3081 -2141 3111 -1941
rect 3176 -2141 3276 -1977
rect 3436 -2141 3536 -1977
rect 3608 -2141 3638 -1941
rect 3890 -2141 4100 -1967
rect 4350 -2141 4928 -1967
rect 5178 -2141 5388 -1967
rect 5657 -2141 5687 -1941
rect 5752 -2141 5852 -1977
rect 6012 -2141 6112 -1977
rect 6184 -2141 6214 -1941
rect 6466 -2141 6676 -1967
rect 6926 -2141 7504 -1967
rect 7754 -2141 7964 -1967
rect 8233 -2141 8263 -1941
rect 8328 -2141 8428 -1977
rect 8588 -2141 8688 -1977
rect 8760 -2141 8790 -1941
rect 9042 -2141 9252 -1967
rect 9502 -2141 10080 -1967
rect 10422 -2141 10632 -1967
rect 10809 -2141 10839 -1941
rect 10904 -2141 11004 -1977
rect 11164 -2141 11264 -1977
rect 11336 -2141 11366 -1941
rect 11710 -2141 11920 -1967
rect 13735 -2141 13765 -1941
rect 13821 -2141 13851 -1941
rect 13907 -2141 13937 -1941
rect 13993 -2141 14023 -1941
rect 14079 -2141 14109 -1941
rect 14165 -2141 14195 -1941
rect 14251 -2141 14281 -1941
rect 14337 -2141 14367 -1941
rect 14423 -2141 14453 -1941
rect 14509 -2141 14539 -1941
rect 14595 -2141 14625 -1941
rect 14681 -2141 14711 -1941
rect 14766 -2141 14796 -1941
rect 14852 -2141 14882 -1941
rect 14938 -2141 14968 -1941
rect 15024 -2141 15054 -1941
rect 15110 -2141 15140 -1941
rect 15196 -2141 15226 -1941
rect 15282 -2141 15312 -1941
rect 15368 -2141 15398 -1941
rect 15666 -2141 16612 -1967
rect -2918 -2409 -2340 -2235
rect -1538 -2409 -960 -2235
rect -802 -2409 -224 -2235
rect 26 -2409 236 -2235
rect 488 -2435 518 -2235
rect 590 -2399 690 -2235
rect 850 -2399 950 -2235
rect 1015 -2435 1045 -2235
rect 1314 -2409 1524 -2235
rect 1774 -2409 2352 -2235
rect 2602 -2409 2812 -2235
rect 3064 -2435 3094 -2235
rect 3166 -2399 3266 -2235
rect 3426 -2399 3526 -2235
rect 3591 -2435 3621 -2235
rect 3890 -2409 4100 -2235
rect 4350 -2409 4928 -2235
rect 5178 -2409 5388 -2235
rect 5640 -2435 5670 -2235
rect 5742 -2399 5842 -2235
rect 6002 -2399 6102 -2235
rect 6167 -2435 6197 -2235
rect 6466 -2409 6676 -2235
rect 6926 -2409 7504 -2235
rect 7754 -2409 7964 -2235
rect 8216 -2435 8246 -2235
rect 8318 -2399 8418 -2235
rect 8578 -2399 8678 -2235
rect 8743 -2435 8773 -2235
rect 9042 -2409 9252 -2235
rect 9502 -2409 10080 -2235
rect 10422 -2409 10632 -2235
rect 10792 -2435 10822 -2235
rect 10894 -2399 10994 -2235
rect 11154 -2399 11254 -2235
rect 11319 -2435 11349 -2235
rect 11710 -2409 11920 -2235
rect 12547 -2435 12577 -2235
rect 12633 -2435 12663 -2235
rect 12719 -2435 12749 -2235
rect 12805 -2435 12835 -2235
rect 12891 -2435 12921 -2235
rect 12977 -2435 13007 -2235
rect 13274 -2409 13484 -2235
rect 13735 -2435 13765 -2235
rect 13821 -2435 13851 -2235
rect 13907 -2435 13937 -2235
rect 13993 -2435 14023 -2235
rect 14079 -2435 14109 -2235
rect 14165 -2435 14195 -2235
rect 14251 -2435 14281 -2235
rect 14337 -2435 14367 -2235
rect 14423 -2435 14453 -2235
rect 14509 -2435 14539 -2235
rect 14595 -2435 14625 -2235
rect 14681 -2435 14711 -2235
rect 14766 -2435 14796 -2235
rect 14852 -2435 14882 -2235
rect 14938 -2435 14968 -2235
rect 15024 -2435 15054 -2235
rect 15110 -2435 15140 -2235
rect 15196 -2435 15226 -2235
rect 15282 -2435 15312 -2235
rect 15368 -2435 15398 -2235
rect 15666 -2409 16612 -2235
rect -2918 -3229 -2340 -3055
rect -1906 -3229 -1876 -3061
rect -1822 -3229 -1792 -3061
rect -1538 -3229 -960 -3055
rect -802 -3229 -224 -3055
rect 26 -3229 236 -3055
rect 505 -3229 535 -3029
rect 600 -3229 700 -3065
rect 860 -3229 960 -3065
rect 1032 -3229 1062 -3029
rect 1314 -3229 1524 -3055
rect 1774 -3229 2352 -3055
rect 2602 -3229 2812 -3055
rect 3081 -3229 3111 -3029
rect 3176 -3229 3276 -3065
rect 3436 -3229 3536 -3065
rect 3608 -3229 3638 -3029
rect 3890 -3229 4100 -3055
rect 4350 -3229 4928 -3055
rect 5178 -3229 5388 -3055
rect 5657 -3229 5687 -3029
rect 5752 -3229 5852 -3065
rect 6012 -3229 6112 -3065
rect 6184 -3229 6214 -3029
rect 6466 -3229 6676 -3055
rect 6926 -3229 7504 -3055
rect 7754 -3229 7964 -3055
rect 8233 -3229 8263 -3029
rect 8328 -3229 8428 -3065
rect 8588 -3229 8688 -3065
rect 8760 -3229 8790 -3029
rect 9042 -3229 9252 -3055
rect 9502 -3229 10080 -3055
rect 10422 -3229 10632 -3055
rect 10809 -3229 10839 -3029
rect 10904 -3229 11004 -3065
rect 11164 -3229 11264 -3065
rect 11336 -3229 11366 -3029
rect 11710 -3229 11920 -3055
rect 13642 -3229 14588 -3055
rect 14838 -3229 15784 -3055
rect 16034 -3229 16612 -3055
rect -2918 -3497 -2340 -3323
rect -1538 -3497 -960 -3323
rect -802 -3497 -224 -3323
rect 26 -3497 236 -3323
rect 505 -3523 535 -3323
rect 600 -3487 700 -3323
rect 860 -3487 960 -3323
rect 1032 -3523 1062 -3323
rect 1314 -3497 1524 -3323
rect 1774 -3497 2352 -3323
rect 2602 -3497 2812 -3323
rect 3081 -3523 3111 -3323
rect 3176 -3487 3276 -3323
rect 3436 -3487 3536 -3323
rect 3608 -3523 3638 -3323
rect 3890 -3497 4100 -3323
rect 4350 -3497 4928 -3323
rect 5178 -3497 5388 -3323
rect 5657 -3523 5687 -3323
rect 5752 -3487 5852 -3323
rect 6012 -3487 6112 -3323
rect 6184 -3523 6214 -3323
rect 6466 -3497 6676 -3323
rect 6926 -3497 7504 -3323
rect 7754 -3497 7964 -3323
rect 8233 -3523 8263 -3323
rect 8328 -3487 8428 -3323
rect 8588 -3487 8688 -3323
rect 8760 -3523 8790 -3323
rect 9042 -3497 9252 -3323
rect 9502 -3497 10080 -3323
rect 10422 -3497 10632 -3323
rect 10809 -3523 10839 -3323
rect 10904 -3487 11004 -3323
rect 11164 -3487 11264 -3323
rect 11336 -3523 11366 -3323
rect 11710 -3497 11920 -3323
rect 13642 -3497 14588 -3323
rect 14838 -3497 15784 -3323
rect 16034 -3497 16612 -3323
rect -2918 -4317 -2340 -4143
rect -1538 -4317 -960 -4143
rect -802 -4317 -224 -4143
rect 26 -4317 236 -4143
rect 488 -4317 518 -4117
rect 590 -4317 690 -4153
rect 850 -4317 950 -4153
rect 1015 -4317 1045 -4117
rect 1314 -4317 1524 -4143
rect 1774 -4317 2352 -4143
rect 2602 -4317 2812 -4143
rect 3064 -4317 3094 -4117
rect 3166 -4317 3266 -4153
rect 3426 -4317 3526 -4153
rect 3591 -4317 3621 -4117
rect 3890 -4317 4100 -4143
rect 4350 -4317 4928 -4143
rect 5178 -4317 5388 -4143
rect 5640 -4317 5670 -4117
rect 5742 -4317 5842 -4153
rect 6002 -4317 6102 -4153
rect 6167 -4317 6197 -4117
rect 6466 -4317 6676 -4143
rect 6926 -4317 7504 -4143
rect 7754 -4317 7964 -4143
rect 8216 -4317 8246 -4117
rect 8318 -4317 8418 -4153
rect 8578 -4317 8678 -4153
rect 8743 -4317 8773 -4117
rect 9042 -4317 9252 -4143
rect 9502 -4317 10080 -4143
rect 10422 -4317 10632 -4143
rect 10792 -4317 10822 -4117
rect 10894 -4317 10994 -4153
rect 11154 -4317 11254 -4153
rect 11319 -4317 11349 -4117
rect 11710 -4317 11920 -4143
rect 12547 -4317 12577 -4117
rect 12633 -4317 12663 -4117
rect 12719 -4317 12749 -4117
rect 12805 -4317 12835 -4117
rect 12891 -4317 12921 -4117
rect 12977 -4317 13007 -4117
rect 13274 -4317 13484 -4143
rect 13735 -4317 13765 -4117
rect 13821 -4317 13851 -4117
rect 13907 -4317 13937 -4117
rect 13993 -4317 14023 -4117
rect 14079 -4317 14109 -4117
rect 14165 -4317 14195 -4117
rect 14251 -4317 14281 -4117
rect 14337 -4317 14367 -4117
rect 14423 -4317 14453 -4117
rect 14509 -4317 14539 -4117
rect 14595 -4317 14625 -4117
rect 14681 -4317 14711 -4117
rect 14766 -4317 14796 -4117
rect 14852 -4317 14882 -4117
rect 14938 -4317 14968 -4117
rect 15024 -4317 15054 -4117
rect 15110 -4317 15140 -4117
rect 15196 -4317 15226 -4117
rect 15282 -4317 15312 -4117
rect 15368 -4317 15398 -4117
rect 15666 -4317 16612 -4143
rect -2918 -4585 -2340 -4411
rect -1538 -4585 -960 -4411
rect -783 -4611 -753 -4411
rect -688 -4575 -588 -4411
rect -428 -4575 -328 -4411
rect -256 -4611 -226 -4411
rect 26 -4585 236 -4411
rect 505 -4611 535 -4411
rect 600 -4575 700 -4411
rect 860 -4575 960 -4411
rect 1032 -4611 1062 -4411
rect 1314 -4585 1524 -4411
rect 1774 -4585 2352 -4411
rect 2602 -4585 2812 -4411
rect 3081 -4611 3111 -4411
rect 3176 -4575 3276 -4411
rect 3436 -4575 3536 -4411
rect 3608 -4611 3638 -4411
rect 3890 -4585 4100 -4411
rect 4350 -4585 4928 -4411
rect 5178 -4585 5388 -4411
rect 5657 -4611 5687 -4411
rect 5752 -4575 5852 -4411
rect 6012 -4575 6112 -4411
rect 6184 -4611 6214 -4411
rect 6466 -4585 6676 -4411
rect 6926 -4585 7504 -4411
rect 7754 -4585 7964 -4411
rect 8233 -4611 8263 -4411
rect 8328 -4575 8428 -4411
rect 8588 -4575 8688 -4411
rect 8760 -4611 8790 -4411
rect 9042 -4585 9252 -4411
rect 9502 -4585 10080 -4411
rect 10422 -4585 10632 -4411
rect 10809 -4611 10839 -4411
rect 10904 -4575 11004 -4411
rect 11164 -4575 11264 -4411
rect 11336 -4611 11366 -4411
rect 11710 -4585 11920 -4411
rect 13735 -4611 13765 -4411
rect 13821 -4611 13851 -4411
rect 13907 -4611 13937 -4411
rect 13993 -4611 14023 -4411
rect 14079 -4611 14109 -4411
rect 14165 -4611 14195 -4411
rect 14251 -4611 14281 -4411
rect 14337 -4611 14367 -4411
rect 14423 -4611 14453 -4411
rect 14509 -4611 14539 -4411
rect 14595 -4611 14625 -4411
rect 14681 -4611 14711 -4411
rect 14766 -4611 14796 -4411
rect 14852 -4611 14882 -4411
rect 14938 -4611 14968 -4411
rect 15024 -4611 15054 -4411
rect 15110 -4611 15140 -4411
rect 15196 -4611 15226 -4411
rect 15282 -4611 15312 -4411
rect 15368 -4611 15398 -4411
rect 15666 -4585 16612 -4411
rect -2918 -5405 -2340 -5231
rect -1538 -5405 -960 -5231
rect -802 -5405 -224 -5231
rect 26 -5405 236 -5231
rect 488 -5405 518 -5205
rect 590 -5405 690 -5241
rect 850 -5405 950 -5241
rect 1015 -5405 1045 -5205
rect 1314 -5405 1524 -5231
rect 1774 -5405 2352 -5231
rect 2602 -5405 2812 -5231
rect 3064 -5405 3094 -5205
rect 3166 -5405 3266 -5241
rect 3426 -5405 3526 -5241
rect 3591 -5405 3621 -5205
rect 3890 -5405 4100 -5231
rect 4350 -5405 4928 -5231
rect 5178 -5405 5388 -5231
rect 5640 -5405 5670 -5205
rect 5742 -5405 5842 -5241
rect 6002 -5405 6102 -5241
rect 6167 -5405 6197 -5205
rect 6466 -5405 6676 -5231
rect 6926 -5405 7504 -5231
rect 7754 -5405 7964 -5231
rect 8216 -5405 8246 -5205
rect 8318 -5405 8418 -5241
rect 8578 -5405 8678 -5241
rect 8743 -5405 8773 -5205
rect 9042 -5405 9252 -5231
rect 9502 -5405 10080 -5231
rect 10422 -5405 10632 -5231
rect 10792 -5405 10822 -5205
rect 10894 -5405 10994 -5241
rect 11154 -5405 11254 -5241
rect 11319 -5405 11349 -5205
rect 11710 -5405 11920 -5231
rect 12547 -5405 12577 -5205
rect 12633 -5405 12663 -5205
rect 12719 -5405 12749 -5205
rect 12805 -5405 12835 -5205
rect 12891 -5405 12921 -5205
rect 12977 -5405 13007 -5205
rect 13274 -5405 13484 -5231
rect 13735 -5405 13765 -5205
rect 13821 -5405 13851 -5205
rect 13907 -5405 13937 -5205
rect 13993 -5405 14023 -5205
rect 14079 -5405 14109 -5205
rect 14165 -5405 14195 -5205
rect 14251 -5405 14281 -5205
rect 14337 -5405 14367 -5205
rect 14423 -5405 14453 -5205
rect 14509 -5405 14539 -5205
rect 14595 -5405 14625 -5205
rect 14681 -5405 14711 -5205
rect 14766 -5405 14796 -5205
rect 14852 -5405 14882 -5205
rect 14938 -5405 14968 -5205
rect 15024 -5405 15054 -5205
rect 15110 -5405 15140 -5205
rect 15196 -5405 15226 -5205
rect 15282 -5405 15312 -5205
rect 15368 -5405 15398 -5205
rect 15666 -5405 16612 -5231
rect -2918 -5673 -2340 -5499
rect -1538 -5673 -960 -5499
rect -802 -5673 -224 -5499
rect 26 -5673 236 -5499
rect 505 -5699 535 -5499
rect 600 -5663 700 -5499
rect 860 -5663 960 -5499
rect 1032 -5699 1062 -5499
rect 1314 -5673 1524 -5499
rect 1774 -5673 2352 -5499
rect 2602 -5673 2812 -5499
rect 3081 -5699 3111 -5499
rect 3176 -5663 3276 -5499
rect 3436 -5663 3536 -5499
rect 3608 -5699 3638 -5499
rect 3890 -5673 4100 -5499
rect 4350 -5673 4928 -5499
rect 5178 -5673 5388 -5499
rect 5657 -5699 5687 -5499
rect 5752 -5663 5852 -5499
rect 6012 -5663 6112 -5499
rect 6184 -5699 6214 -5499
rect 6466 -5673 6676 -5499
rect 6926 -5673 7504 -5499
rect 7754 -5673 7964 -5499
rect 8233 -5699 8263 -5499
rect 8328 -5663 8428 -5499
rect 8588 -5663 8688 -5499
rect 8760 -5699 8790 -5499
rect 9042 -5673 9252 -5499
rect 9502 -5673 10080 -5499
rect 10422 -5673 10632 -5499
rect 10809 -5699 10839 -5499
rect 10904 -5663 11004 -5499
rect 11164 -5663 11264 -5499
rect 11336 -5699 11366 -5499
rect 11710 -5673 11920 -5499
rect 13735 -5699 13765 -5499
rect 13821 -5699 13851 -5499
rect 13907 -5699 13937 -5499
rect 13993 -5699 14023 -5499
rect 14079 -5699 14109 -5499
rect 14165 -5699 14195 -5499
rect 14251 -5699 14281 -5499
rect 14337 -5699 14367 -5499
rect 14423 -5699 14453 -5499
rect 14509 -5699 14539 -5499
rect 14595 -5699 14625 -5499
rect 14681 -5699 14711 -5499
rect 14766 -5699 14796 -5499
rect 14852 -5699 14882 -5499
rect 14938 -5699 14968 -5499
rect 15024 -5699 15054 -5499
rect 15110 -5699 15140 -5499
rect 15196 -5699 15226 -5499
rect 15282 -5699 15312 -5499
rect 15368 -5699 15398 -5499
rect 15666 -5673 16612 -5499
rect -2918 -6493 -2340 -6319
rect -1354 -6493 -1144 -6319
rect -890 -6493 -860 -6293
rect -806 -6493 -776 -6293
rect -526 -6493 -316 -6319
rect -57 -6493 -27 -6293
rect 29 -6493 59 -6293
rect 115 -6493 145 -6293
rect 201 -6493 231 -6293
rect 287 -6493 317 -6293
rect 373 -6493 403 -6293
rect 670 -6493 880 -6319
rect 1130 -6493 1160 -6325
rect 1214 -6493 1244 -6325
rect 1498 -6493 1708 -6319
rect 1958 -6493 2168 -6319
rect 2420 -6493 2450 -6293
rect 2522 -6493 2622 -6329
rect 2782 -6493 2882 -6329
rect 2947 -6493 2977 -6293
rect 3246 -6493 3456 -6319
rect 4442 -6493 5388 -6319
rect 6466 -6493 6676 -6319
rect 6928 -6493 6958 -6293
rect 7030 -6493 7130 -6329
rect 7290 -6493 7390 -6329
rect 7455 -6493 7485 -6293
rect 7754 -6493 7964 -6319
rect 8216 -6493 8246 -6293
rect 8318 -6493 8418 -6329
rect 8578 -6493 8678 -6329
rect 8743 -6493 8773 -6293
rect 9042 -6493 9252 -6319
rect 9504 -6493 9534 -6293
rect 9606 -6493 9706 -6329
rect 9866 -6493 9966 -6329
rect 10031 -6493 10061 -6293
rect 10330 -6493 10540 -6319
rect 10790 -6493 10820 -6293
rect 10874 -6493 10904 -6293
rect 10958 -6493 10988 -6293
rect 11042 -6493 11072 -6293
rect 11126 -6493 11156 -6293
rect 11210 -6493 11240 -6293
rect 11294 -6493 11324 -6293
rect 11378 -6493 11408 -6293
rect 11710 -6493 11920 -6319
rect 13642 -6493 14588 -6319
rect 14838 -6493 15784 -6319
rect 16034 -6493 16612 -6319
rect -2918 -6761 -2800 -6587
rect -2550 -6721 -2520 -6593
rect -2466 -6721 -2436 -6593
rect -2278 -6671 -2248 -6587
rect -2193 -6671 -2163 -6587
rect -2098 -6671 -2068 -6587
rect -1995 -6671 -1965 -6587
rect -1863 -6737 -1833 -6587
rect -1768 -6671 -1738 -6587
rect -1684 -6671 -1654 -6587
rect -1570 -6671 -1540 -6587
rect -1359 -6787 -1329 -6587
rect -1275 -6787 -1245 -6587
rect -1087 -6715 -1057 -6587
rect -990 -6787 -960 -6587
rect -802 -6761 -224 -6587
rect 26 -6761 604 -6587
rect 762 -6761 1340 -6587
rect 1590 -6761 2168 -6587
rect 2326 -6761 2904 -6587
rect 3154 -6761 3732 -6587
rect 3890 -6761 4468 -6587
rect 4718 -6761 5296 -6587
rect 5454 -6761 6032 -6587
rect 6282 -6761 6860 -6587
rect 7018 -6761 7596 -6587
rect 7846 -6761 8424 -6587
rect 8582 -6761 9160 -6587
rect 16034 -6761 16612 -6587
rect -2918 -7581 -2340 -7407
rect -1538 -7581 -960 -7407
rect -802 -7581 -224 -7407
rect 26 -7581 604 -7407
rect 762 -7581 1340 -7407
rect 1590 -7581 2168 -7407
rect 2326 -7581 2536 -7407
rect 2974 -7581 3004 -7413
rect 3058 -7581 3088 -7413
rect 3338 -7581 3548 -7407
rect 3802 -7581 3832 -7381
rect 3886 -7581 3916 -7381
rect 4166 -7581 4376 -7407
rect 4626 -7581 4656 -7381
rect 4735 -7542 4765 -7458
rect 4838 -7542 4868 -7458
rect 5052 -7542 5082 -7458
rect 5124 -7542 5154 -7458
rect 5220 -7542 5250 -7458
rect 5546 -7581 5756 -7407
rect 6006 -7581 6036 -7381
rect 6103 -7581 6133 -7453
rect 6291 -7581 6321 -7381
rect 6375 -7581 6405 -7381
rect 6586 -7581 6616 -7497
rect 6700 -7581 6730 -7497
rect 6784 -7581 6814 -7497
rect 6879 -7581 6909 -7431
rect 7011 -7581 7041 -7497
rect 7114 -7581 7144 -7497
rect 7209 -7581 7239 -7497
rect 7294 -7581 7324 -7497
rect 7482 -7575 7512 -7447
rect 7566 -7575 7596 -7447
rect 7846 -7581 8424 -7407
rect 8582 -7581 9160 -7407
rect 16034 -7581 16612 -7407
rect -2918 -7849 -2340 -7675
rect -1354 -7849 -1144 -7675
rect -890 -7875 -860 -7675
rect -806 -7875 -776 -7675
rect -526 -7849 -316 -7675
rect -57 -7875 -27 -7675
rect 29 -7875 59 -7675
rect 115 -7875 145 -7675
rect 201 -7875 231 -7675
rect 287 -7875 317 -7675
rect 373 -7875 403 -7675
rect 670 -7849 880 -7675
rect 1130 -7843 1160 -7675
rect 1214 -7843 1244 -7675
rect 1498 -7849 1708 -7675
rect 1958 -7849 2168 -7675
rect 2420 -7875 2450 -7675
rect 2522 -7839 2622 -7675
rect 2782 -7839 2882 -7675
rect 2947 -7875 2977 -7675
rect 3246 -7849 3456 -7675
rect 4442 -7849 5388 -7675
rect 6466 -7849 6676 -7675
rect 6928 -7875 6958 -7675
rect 7030 -7839 7130 -7675
rect 7290 -7839 7390 -7675
rect 7455 -7875 7485 -7675
rect 7754 -7849 7964 -7675
rect 8216 -7875 8246 -7675
rect 8318 -7839 8418 -7675
rect 8578 -7839 8678 -7675
rect 8743 -7875 8773 -7675
rect 9042 -7849 9252 -7675
rect 9504 -7875 9534 -7675
rect 9606 -7839 9706 -7675
rect 9866 -7839 9966 -7675
rect 10031 -7875 10061 -7675
rect 10330 -7849 10540 -7675
rect 10790 -7875 10820 -7675
rect 10874 -7875 10904 -7675
rect 10958 -7875 10988 -7675
rect 11042 -7875 11072 -7675
rect 11126 -7875 11156 -7675
rect 11210 -7875 11240 -7675
rect 11294 -7875 11324 -7675
rect 11378 -7875 11408 -7675
rect 11710 -7849 11920 -7675
rect 13642 -7849 14588 -7675
rect 14838 -7849 15784 -7675
rect 16034 -7849 16612 -7675
rect -2918 -8669 -2340 -8495
rect -1538 -8669 -960 -8495
rect -802 -8669 -224 -8495
rect 26 -8669 236 -8495
rect 505 -8669 535 -8469
rect 600 -8669 700 -8505
rect 860 -8669 960 -8505
rect 1032 -8669 1062 -8469
rect 1314 -8669 1524 -8495
rect 1774 -8669 2352 -8495
rect 2602 -8669 2812 -8495
rect 3081 -8669 3111 -8469
rect 3176 -8669 3276 -8505
rect 3436 -8669 3536 -8505
rect 3608 -8669 3638 -8469
rect 3890 -8669 4100 -8495
rect 4350 -8669 4928 -8495
rect 5178 -8669 5388 -8495
rect 5657 -8669 5687 -8469
rect 5752 -8669 5852 -8505
rect 6012 -8669 6112 -8505
rect 6184 -8669 6214 -8469
rect 6466 -8669 6676 -8495
rect 6926 -8669 7504 -8495
rect 7754 -8669 7964 -8495
rect 8233 -8669 8263 -8469
rect 8328 -8669 8428 -8505
rect 8588 -8669 8688 -8505
rect 8760 -8669 8790 -8469
rect 9042 -8669 9252 -8495
rect 9502 -8669 10080 -8495
rect 10422 -8669 10632 -8495
rect 10809 -8669 10839 -8469
rect 10904 -8669 11004 -8505
rect 11164 -8669 11264 -8505
rect 11336 -8669 11366 -8469
rect 11710 -8669 11920 -8495
rect 13735 -8669 13765 -8469
rect 13821 -8669 13851 -8469
rect 13907 -8669 13937 -8469
rect 13993 -8669 14023 -8469
rect 14079 -8669 14109 -8469
rect 14165 -8669 14195 -8469
rect 14251 -8669 14281 -8469
rect 14337 -8669 14367 -8469
rect 14423 -8669 14453 -8469
rect 14509 -8669 14539 -8469
rect 14595 -8669 14625 -8469
rect 14681 -8669 14711 -8469
rect 14766 -8669 14796 -8469
rect 14852 -8669 14882 -8469
rect 14938 -8669 14968 -8469
rect 15024 -8669 15054 -8469
rect 15110 -8669 15140 -8469
rect 15196 -8669 15226 -8469
rect 15282 -8669 15312 -8469
rect 15368 -8669 15398 -8469
rect 15666 -8669 16612 -8495
rect -2918 -8937 -2340 -8763
rect -1538 -8937 -960 -8763
rect -802 -8937 -224 -8763
rect 26 -8937 236 -8763
rect 488 -8963 518 -8763
rect 590 -8927 690 -8763
rect 850 -8927 950 -8763
rect 1015 -8963 1045 -8763
rect 1314 -8937 1524 -8763
rect 1774 -8937 2352 -8763
rect 2602 -8937 2812 -8763
rect 3064 -8963 3094 -8763
rect 3166 -8927 3266 -8763
rect 3426 -8927 3526 -8763
rect 3591 -8963 3621 -8763
rect 3890 -8937 4100 -8763
rect 4350 -8937 4928 -8763
rect 5178 -8937 5388 -8763
rect 5640 -8963 5670 -8763
rect 5742 -8927 5842 -8763
rect 6002 -8927 6102 -8763
rect 6167 -8963 6197 -8763
rect 6466 -8937 6676 -8763
rect 6926 -8937 7504 -8763
rect 7754 -8937 7964 -8763
rect 8216 -8963 8246 -8763
rect 8318 -8927 8418 -8763
rect 8578 -8927 8678 -8763
rect 8743 -8963 8773 -8763
rect 9042 -8937 9252 -8763
rect 9502 -8937 10080 -8763
rect 10422 -8937 10632 -8763
rect 10792 -8963 10822 -8763
rect 10894 -8927 10994 -8763
rect 11154 -8927 11254 -8763
rect 11319 -8963 11349 -8763
rect 11710 -8937 11920 -8763
rect 12547 -8963 12577 -8763
rect 12633 -8963 12663 -8763
rect 12719 -8963 12749 -8763
rect 12805 -8963 12835 -8763
rect 12891 -8963 12921 -8763
rect 12977 -8963 13007 -8763
rect 13274 -8937 13484 -8763
rect 13735 -8963 13765 -8763
rect 13821 -8963 13851 -8763
rect 13907 -8963 13937 -8763
rect 13993 -8963 14023 -8763
rect 14079 -8963 14109 -8763
rect 14165 -8963 14195 -8763
rect 14251 -8963 14281 -8763
rect 14337 -8963 14367 -8763
rect 14423 -8963 14453 -8763
rect 14509 -8963 14539 -8763
rect 14595 -8963 14625 -8763
rect 14681 -8963 14711 -8763
rect 14766 -8963 14796 -8763
rect 14852 -8963 14882 -8763
rect 14938 -8963 14968 -8763
rect 15024 -8963 15054 -8763
rect 15110 -8963 15140 -8763
rect 15196 -8963 15226 -8763
rect 15282 -8963 15312 -8763
rect 15368 -8963 15398 -8763
rect 15666 -8937 16612 -8763
rect -2918 -9757 -2340 -9583
rect -1538 -9757 -960 -9583
rect -783 -9757 -753 -9557
rect -688 -9757 -588 -9593
rect -428 -9757 -328 -9593
rect -256 -9757 -226 -9557
rect 26 -9757 236 -9583
rect 505 -9757 535 -9557
rect 600 -9757 700 -9593
rect 860 -9757 960 -9593
rect 1032 -9757 1062 -9557
rect 1314 -9757 1524 -9583
rect 1774 -9757 2352 -9583
rect 2602 -9757 2812 -9583
rect 3081 -9757 3111 -9557
rect 3176 -9757 3276 -9593
rect 3436 -9757 3536 -9593
rect 3608 -9757 3638 -9557
rect 3890 -9757 4100 -9583
rect 4350 -9757 4928 -9583
rect 5178 -9757 5388 -9583
rect 5657 -9757 5687 -9557
rect 5752 -9757 5852 -9593
rect 6012 -9757 6112 -9593
rect 6184 -9757 6214 -9557
rect 6466 -9757 6676 -9583
rect 6926 -9757 7504 -9583
rect 7754 -9757 7964 -9583
rect 8233 -9757 8263 -9557
rect 8328 -9757 8428 -9593
rect 8588 -9757 8688 -9593
rect 8760 -9757 8790 -9557
rect 9042 -9757 9252 -9583
rect 9502 -9757 10080 -9583
rect 10422 -9757 10632 -9583
rect 10809 -9757 10839 -9557
rect 10904 -9757 11004 -9593
rect 11164 -9757 11264 -9593
rect 11336 -9757 11366 -9557
rect 11710 -9757 11920 -9583
rect 13735 -9757 13765 -9557
rect 13821 -9757 13851 -9557
rect 13907 -9757 13937 -9557
rect 13993 -9757 14023 -9557
rect 14079 -9757 14109 -9557
rect 14165 -9757 14195 -9557
rect 14251 -9757 14281 -9557
rect 14337 -9757 14367 -9557
rect 14423 -9757 14453 -9557
rect 14509 -9757 14539 -9557
rect 14595 -9757 14625 -9557
rect 14681 -9757 14711 -9557
rect 14766 -9757 14796 -9557
rect 14852 -9757 14882 -9557
rect 14938 -9757 14968 -9557
rect 15024 -9757 15054 -9557
rect 15110 -9757 15140 -9557
rect 15196 -9757 15226 -9557
rect 15282 -9757 15312 -9557
rect 15368 -9757 15398 -9557
rect 15666 -9757 16612 -9583
rect -2918 -10025 -2340 -9851
rect -1538 -10025 -960 -9851
rect -802 -10025 -224 -9851
rect 26 -10025 236 -9851
rect 488 -10051 518 -9851
rect 590 -10015 690 -9851
rect 850 -10015 950 -9851
rect 1015 -10051 1045 -9851
rect 1314 -10025 1524 -9851
rect 1774 -10025 2352 -9851
rect 2602 -10025 2812 -9851
rect 3064 -10051 3094 -9851
rect 3166 -10015 3266 -9851
rect 3426 -10015 3526 -9851
rect 3591 -10051 3621 -9851
rect 3890 -10025 4100 -9851
rect 4350 -10025 4928 -9851
rect 5178 -10025 5388 -9851
rect 5640 -10051 5670 -9851
rect 5742 -10015 5842 -9851
rect 6002 -10015 6102 -9851
rect 6167 -10051 6197 -9851
rect 6466 -10025 6676 -9851
rect 6926 -10025 7504 -9851
rect 7754 -10025 7964 -9851
rect 8216 -10051 8246 -9851
rect 8318 -10015 8418 -9851
rect 8578 -10015 8678 -9851
rect 8743 -10051 8773 -9851
rect 9042 -10025 9252 -9851
rect 9502 -10025 10080 -9851
rect 10422 -10025 10632 -9851
rect 10792 -10051 10822 -9851
rect 10894 -10015 10994 -9851
rect 11154 -10015 11254 -9851
rect 11319 -10051 11349 -9851
rect 11710 -10025 11920 -9851
rect 12547 -10051 12577 -9851
rect 12633 -10051 12663 -9851
rect 12719 -10051 12749 -9851
rect 12805 -10051 12835 -9851
rect 12891 -10051 12921 -9851
rect 12977 -10051 13007 -9851
rect 13274 -10025 13484 -9851
rect 13735 -10051 13765 -9851
rect 13821 -10051 13851 -9851
rect 13907 -10051 13937 -9851
rect 13993 -10051 14023 -9851
rect 14079 -10051 14109 -9851
rect 14165 -10051 14195 -9851
rect 14251 -10051 14281 -9851
rect 14337 -10051 14367 -9851
rect 14423 -10051 14453 -9851
rect 14509 -10051 14539 -9851
rect 14595 -10051 14625 -9851
rect 14681 -10051 14711 -9851
rect 14766 -10051 14796 -9851
rect 14852 -10051 14882 -9851
rect 14938 -10051 14968 -9851
rect 15024 -10051 15054 -9851
rect 15110 -10051 15140 -9851
rect 15196 -10051 15226 -9851
rect 15282 -10051 15312 -9851
rect 15368 -10051 15398 -9851
rect 15666 -10025 16612 -9851
rect -2918 -10845 -2340 -10671
rect -1906 -10845 -1876 -10677
rect -1822 -10845 -1792 -10677
rect -1538 -10845 -960 -10671
rect -802 -10845 -224 -10671
rect 26 -10845 236 -10671
rect 505 -10845 535 -10645
rect 600 -10845 700 -10681
rect 860 -10845 960 -10681
rect 1032 -10845 1062 -10645
rect 1314 -10845 1524 -10671
rect 1774 -10845 2352 -10671
rect 2602 -10845 2812 -10671
rect 3081 -10845 3111 -10645
rect 3176 -10845 3276 -10681
rect 3436 -10845 3536 -10681
rect 3608 -10845 3638 -10645
rect 3890 -10845 4100 -10671
rect 4350 -10845 4928 -10671
rect 5178 -10845 5388 -10671
rect 5657 -10845 5687 -10645
rect 5752 -10845 5852 -10681
rect 6012 -10845 6112 -10681
rect 6184 -10845 6214 -10645
rect 6466 -10845 6676 -10671
rect 6926 -10845 7504 -10671
rect 7754 -10845 7964 -10671
rect 8233 -10845 8263 -10645
rect 8328 -10845 8428 -10681
rect 8588 -10845 8688 -10681
rect 8760 -10845 8790 -10645
rect 9042 -10845 9252 -10671
rect 9502 -10845 10080 -10671
rect 10422 -10845 10632 -10671
rect 10809 -10845 10839 -10645
rect 10904 -10845 11004 -10681
rect 11164 -10845 11264 -10681
rect 11336 -10845 11366 -10645
rect 11710 -10845 11920 -10671
rect 13642 -10845 14588 -10671
rect 14838 -10845 15784 -10671
rect 16034 -10845 16612 -10671
rect -2918 -11113 -2340 -10939
rect -1538 -11113 -960 -10939
rect -802 -11113 -224 -10939
rect 26 -11113 236 -10939
rect 505 -11139 535 -10939
rect 600 -11103 700 -10939
rect 860 -11103 960 -10939
rect 1032 -11139 1062 -10939
rect 1314 -11113 1524 -10939
rect 1774 -11113 2352 -10939
rect 2602 -11113 2812 -10939
rect 3081 -11139 3111 -10939
rect 3176 -11103 3276 -10939
rect 3436 -11103 3536 -10939
rect 3608 -11139 3638 -10939
rect 3890 -11113 4100 -10939
rect 4350 -11113 4928 -10939
rect 5178 -11113 5388 -10939
rect 5657 -11139 5687 -10939
rect 5752 -11103 5852 -10939
rect 6012 -11103 6112 -10939
rect 6184 -11139 6214 -10939
rect 6466 -11113 6676 -10939
rect 6926 -11113 7504 -10939
rect 7754 -11113 7964 -10939
rect 8233 -11139 8263 -10939
rect 8328 -11103 8428 -10939
rect 8588 -11103 8688 -10939
rect 8760 -11139 8790 -10939
rect 9042 -11113 9252 -10939
rect 9502 -11113 10080 -10939
rect 10422 -11113 10632 -10939
rect 10809 -11139 10839 -10939
rect 10904 -11103 11004 -10939
rect 11164 -11103 11264 -10939
rect 11336 -11139 11366 -10939
rect 11710 -11113 11920 -10939
rect 13642 -11113 14588 -10939
rect 14838 -11113 15784 -10939
rect 16034 -11113 16612 -10939
rect -2918 -11933 -2340 -11759
rect -1538 -11933 -960 -11759
rect -802 -11933 -224 -11759
rect 26 -11933 236 -11759
rect 488 -11933 518 -11733
rect 590 -11933 690 -11769
rect 850 -11933 950 -11769
rect 1015 -11933 1045 -11733
rect 1314 -11933 1524 -11759
rect 1774 -11933 2352 -11759
rect 2602 -11933 2812 -11759
rect 3064 -11933 3094 -11733
rect 3166 -11933 3266 -11769
rect 3426 -11933 3526 -11769
rect 3591 -11933 3621 -11733
rect 3890 -11933 4100 -11759
rect 4350 -11933 4928 -11759
rect 5178 -11933 5388 -11759
rect 5640 -11933 5670 -11733
rect 5742 -11933 5842 -11769
rect 6002 -11933 6102 -11769
rect 6167 -11933 6197 -11733
rect 6466 -11933 6676 -11759
rect 6926 -11933 7504 -11759
rect 7754 -11933 7964 -11759
rect 8216 -11933 8246 -11733
rect 8318 -11933 8418 -11769
rect 8578 -11933 8678 -11769
rect 8743 -11933 8773 -11733
rect 9042 -11933 9252 -11759
rect 9502 -11933 10080 -11759
rect 10422 -11933 10632 -11759
rect 10792 -11933 10822 -11733
rect 10894 -11933 10994 -11769
rect 11154 -11933 11254 -11769
rect 11319 -11933 11349 -11733
rect 11710 -11933 11920 -11759
rect 12547 -11933 12577 -11733
rect 12633 -11933 12663 -11733
rect 12719 -11933 12749 -11733
rect 12805 -11933 12835 -11733
rect 12891 -11933 12921 -11733
rect 12977 -11933 13007 -11733
rect 13274 -11933 13484 -11759
rect 13735 -11933 13765 -11733
rect 13821 -11933 13851 -11733
rect 13907 -11933 13937 -11733
rect 13993 -11933 14023 -11733
rect 14079 -11933 14109 -11733
rect 14165 -11933 14195 -11733
rect 14251 -11933 14281 -11733
rect 14337 -11933 14367 -11733
rect 14423 -11933 14453 -11733
rect 14509 -11933 14539 -11733
rect 14595 -11933 14625 -11733
rect 14681 -11933 14711 -11733
rect 14766 -11933 14796 -11733
rect 14852 -11933 14882 -11733
rect 14938 -11933 14968 -11733
rect 15024 -11933 15054 -11733
rect 15110 -11933 15140 -11733
rect 15196 -11933 15226 -11733
rect 15282 -11933 15312 -11733
rect 15368 -11933 15398 -11733
rect 15666 -11933 16612 -11759
rect -2918 -12201 -2340 -12027
rect -1538 -12201 -960 -12027
rect -783 -12227 -753 -12027
rect -688 -12191 -588 -12027
rect -428 -12191 -328 -12027
rect -256 -12227 -226 -12027
rect 26 -12201 236 -12027
rect 505 -12227 535 -12027
rect 600 -12191 700 -12027
rect 860 -12191 960 -12027
rect 1032 -12227 1062 -12027
rect 1314 -12201 1524 -12027
rect 1774 -12201 2352 -12027
rect 2602 -12201 2812 -12027
rect 3081 -12227 3111 -12027
rect 3176 -12191 3276 -12027
rect 3436 -12191 3536 -12027
rect 3608 -12227 3638 -12027
rect 3890 -12201 4100 -12027
rect 4350 -12201 4928 -12027
rect 5178 -12201 5388 -12027
rect 5657 -12227 5687 -12027
rect 5752 -12191 5852 -12027
rect 6012 -12191 6112 -12027
rect 6184 -12227 6214 -12027
rect 6466 -12201 6676 -12027
rect 6926 -12201 7504 -12027
rect 7754 -12201 7964 -12027
rect 8233 -12227 8263 -12027
rect 8328 -12191 8428 -12027
rect 8588 -12191 8688 -12027
rect 8760 -12227 8790 -12027
rect 9042 -12201 9252 -12027
rect 9502 -12201 10080 -12027
rect 10422 -12201 10632 -12027
rect 10809 -12227 10839 -12027
rect 10904 -12191 11004 -12027
rect 11164 -12191 11264 -12027
rect 11336 -12227 11366 -12027
rect 11710 -12201 11920 -12027
rect 13735 -12227 13765 -12027
rect 13821 -12227 13851 -12027
rect 13907 -12227 13937 -12027
rect 13993 -12227 14023 -12027
rect 14079 -12227 14109 -12027
rect 14165 -12227 14195 -12027
rect 14251 -12227 14281 -12027
rect 14337 -12227 14367 -12027
rect 14423 -12227 14453 -12027
rect 14509 -12227 14539 -12027
rect 14595 -12227 14625 -12027
rect 14681 -12227 14711 -12027
rect 14766 -12227 14796 -12027
rect 14852 -12227 14882 -12027
rect 14938 -12227 14968 -12027
rect 15024 -12227 15054 -12027
rect 15110 -12227 15140 -12027
rect 15196 -12227 15226 -12027
rect 15282 -12227 15312 -12027
rect 15368 -12227 15398 -12027
rect 15666 -12201 16612 -12027
rect -2918 -13021 -2340 -12847
rect -1538 -13021 -960 -12847
rect -802 -13021 -224 -12847
rect 26 -13021 236 -12847
rect 488 -13021 518 -12821
rect 590 -13021 690 -12857
rect 850 -13021 950 -12857
rect 1015 -13021 1045 -12821
rect 1314 -13021 1524 -12847
rect 1774 -13021 2352 -12847
rect 2602 -13021 2812 -12847
rect 3064 -13021 3094 -12821
rect 3166 -13021 3266 -12857
rect 3426 -13021 3526 -12857
rect 3591 -13021 3621 -12821
rect 3890 -13021 4100 -12847
rect 4350 -13021 4928 -12847
rect 5178 -13021 5388 -12847
rect 5640 -13021 5670 -12821
rect 5742 -13021 5842 -12857
rect 6002 -13021 6102 -12857
rect 6167 -13021 6197 -12821
rect 6466 -13021 6676 -12847
rect 6926 -13021 7504 -12847
rect 7754 -13021 7964 -12847
rect 8216 -13021 8246 -12821
rect 8318 -13021 8418 -12857
rect 8578 -13021 8678 -12857
rect 8743 -13021 8773 -12821
rect 9042 -13021 9252 -12847
rect 9502 -13021 10080 -12847
rect 10422 -13021 10632 -12847
rect 10792 -13021 10822 -12821
rect 10894 -13021 10994 -12857
rect 11154 -13021 11254 -12857
rect 11319 -13021 11349 -12821
rect 11710 -13021 11920 -12847
rect 12547 -13021 12577 -12821
rect 12633 -13021 12663 -12821
rect 12719 -13021 12749 -12821
rect 12805 -13021 12835 -12821
rect 12891 -13021 12921 -12821
rect 12977 -13021 13007 -12821
rect 13274 -13021 13484 -12847
rect 13735 -13021 13765 -12821
rect 13821 -13021 13851 -12821
rect 13907 -13021 13937 -12821
rect 13993 -13021 14023 -12821
rect 14079 -13021 14109 -12821
rect 14165 -13021 14195 -12821
rect 14251 -13021 14281 -12821
rect 14337 -13021 14367 -12821
rect 14423 -13021 14453 -12821
rect 14509 -13021 14539 -12821
rect 14595 -13021 14625 -12821
rect 14681 -13021 14711 -12821
rect 14766 -13021 14796 -12821
rect 14852 -13021 14882 -12821
rect 14938 -13021 14968 -12821
rect 15024 -13021 15054 -12821
rect 15110 -13021 15140 -12821
rect 15196 -13021 15226 -12821
rect 15282 -13021 15312 -12821
rect 15368 -13021 15398 -12821
rect 15666 -13021 16612 -12847
rect -2918 -13289 -2340 -13115
rect -1538 -13289 -960 -13115
rect -802 -13289 -224 -13115
rect 26 -13289 236 -13115
rect 505 -13315 535 -13115
rect 600 -13279 700 -13115
rect 860 -13279 960 -13115
rect 1032 -13315 1062 -13115
rect 1314 -13289 1524 -13115
rect 1774 -13289 2352 -13115
rect 2602 -13289 2812 -13115
rect 3081 -13315 3111 -13115
rect 3176 -13279 3276 -13115
rect 3436 -13279 3536 -13115
rect 3608 -13315 3638 -13115
rect 3890 -13289 4100 -13115
rect 4350 -13289 4928 -13115
rect 5178 -13289 5388 -13115
rect 5657 -13315 5687 -13115
rect 5752 -13279 5852 -13115
rect 6012 -13279 6112 -13115
rect 6184 -13315 6214 -13115
rect 6466 -13289 6676 -13115
rect 6926 -13289 7504 -13115
rect 7754 -13289 7964 -13115
rect 8233 -13315 8263 -13115
rect 8328 -13279 8428 -13115
rect 8588 -13279 8688 -13115
rect 8760 -13315 8790 -13115
rect 9042 -13289 9252 -13115
rect 9502 -13289 10080 -13115
rect 10422 -13289 10632 -13115
rect 10809 -13315 10839 -13115
rect 10904 -13279 11004 -13115
rect 11164 -13279 11264 -13115
rect 11336 -13315 11366 -13115
rect 11710 -13289 11920 -13115
rect 13735 -13315 13765 -13115
rect 13821 -13315 13851 -13115
rect 13907 -13315 13937 -13115
rect 13993 -13315 14023 -13115
rect 14079 -13315 14109 -13115
rect 14165 -13315 14195 -13115
rect 14251 -13315 14281 -13115
rect 14337 -13315 14367 -13115
rect 14423 -13315 14453 -13115
rect 14509 -13315 14539 -13115
rect 14595 -13315 14625 -13115
rect 14681 -13315 14711 -13115
rect 14766 -13315 14796 -13115
rect 14852 -13315 14882 -13115
rect 14938 -13315 14968 -13115
rect 15024 -13315 15054 -13115
rect 15110 -13315 15140 -13115
rect 15196 -13315 15226 -13115
rect 15282 -13315 15312 -13115
rect 15368 -13315 15398 -13115
rect 15666 -13289 16612 -13115
rect -2918 -14109 -2340 -13935
rect -1354 -14109 -1144 -13935
rect -890 -14109 -860 -13909
rect -806 -14109 -776 -13909
rect -526 -14109 -316 -13935
rect -57 -14109 -27 -13909
rect 29 -14109 59 -13909
rect 115 -14109 145 -13909
rect 201 -14109 231 -13909
rect 287 -14109 317 -13909
rect 373 -14109 403 -13909
rect 670 -14109 880 -13935
rect 1130 -14109 1160 -13941
rect 1214 -14109 1244 -13941
rect 1498 -14109 1708 -13935
rect 1958 -14109 2168 -13935
rect 2420 -14109 2450 -13909
rect 2522 -14109 2622 -13945
rect 2782 -14109 2882 -13945
rect 2947 -14109 2977 -13909
rect 3246 -14109 3456 -13935
rect 4442 -14109 5388 -13935
rect 6466 -14109 6676 -13935
rect 6928 -14109 6958 -13909
rect 7030 -14109 7130 -13945
rect 7290 -14109 7390 -13945
rect 7455 -14109 7485 -13909
rect 7754 -14109 7964 -13935
rect 8216 -14109 8246 -13909
rect 8318 -14109 8418 -13945
rect 8578 -14109 8678 -13945
rect 8743 -14109 8773 -13909
rect 9042 -14109 9252 -13935
rect 9504 -14109 9534 -13909
rect 9606 -14109 9706 -13945
rect 9866 -14109 9966 -13945
rect 10031 -14109 10061 -13909
rect 10330 -14109 10540 -13935
rect 10790 -14109 10820 -13909
rect 10874 -14109 10904 -13909
rect 10958 -14109 10988 -13909
rect 11042 -14109 11072 -13909
rect 11126 -14109 11156 -13909
rect 11210 -14109 11240 -13909
rect 11294 -14109 11324 -13909
rect 11378 -14109 11408 -13909
rect 11710 -14109 11920 -13935
rect 13642 -14109 14588 -13935
rect 14838 -14109 15784 -13935
rect 16034 -14109 16612 -13935
<< ndiff >>
rect -2970 -444 -2918 -399
rect -2970 -478 -2962 -444
rect -2928 -478 -2918 -444
rect -2970 -509 -2918 -478
rect -2340 -444 -2288 -399
rect -2340 -478 -2330 -444
rect -2296 -478 -2288 -444
rect -2340 -509 -2288 -478
rect -1406 -437 -1354 -399
rect -1406 -471 -1398 -437
rect -1364 -471 -1354 -437
rect -1406 -509 -1354 -471
rect -1144 -437 -1092 -399
rect -1144 -471 -1134 -437
rect -1100 -471 -1092 -437
rect -1144 -509 -1092 -471
rect -942 -395 -890 -379
rect -942 -429 -934 -395
rect -900 -429 -890 -395
rect -942 -463 -890 -429
rect -942 -497 -934 -463
rect -900 -497 -890 -463
rect -942 -509 -890 -497
rect -860 -509 -806 -379
rect -776 -395 -724 -379
rect -776 -429 -766 -395
rect -732 -429 -724 -395
rect -776 -463 -724 -429
rect -776 -497 -766 -463
rect -732 -497 -724 -463
rect -578 -437 -526 -399
rect -578 -471 -570 -437
rect -536 -471 -526 -437
rect -776 -509 -724 -497
rect -578 -509 -526 -471
rect -316 -437 -264 -399
rect -316 -471 -306 -437
rect -272 -471 -264 -437
rect -316 -509 -264 -471
rect -37 -461 29 -425
rect -37 -495 -16 -461
rect 18 -495 29 -461
rect -37 -509 29 -495
rect 59 -450 115 -425
rect 59 -484 70 -450
rect 104 -484 115 -450
rect 59 -509 115 -484
rect 145 -461 201 -425
rect 145 -495 156 -461
rect 190 -495 201 -461
rect 145 -509 201 -495
rect 231 -450 287 -425
rect 231 -484 242 -450
rect 276 -484 287 -450
rect 231 -509 287 -484
rect 317 -461 396 -425
rect 317 -495 328 -461
rect 362 -495 396 -461
rect 618 -437 670 -399
rect 618 -471 626 -437
rect 660 -471 670 -437
rect 317 -509 396 -495
rect 618 -509 670 -471
rect 880 -437 932 -399
rect 880 -471 890 -437
rect 924 -471 932 -437
rect 880 -509 932 -471
rect 1161 -452 1213 -425
rect 1161 -486 1169 -452
rect 1203 -486 1213 -452
rect 1161 -509 1213 -486
rect 1243 -454 1300 -425
rect 1243 -488 1253 -454
rect 1287 -488 1300 -454
rect 1243 -509 1300 -488
rect 1446 -437 1498 -399
rect 1446 -471 1454 -437
rect 1488 -471 1498 -437
rect 1446 -509 1498 -471
rect 1708 -437 1760 -399
rect 1708 -471 1718 -437
rect 1752 -471 1760 -437
rect 1708 -509 1760 -471
rect 1906 -437 1958 -399
rect 1906 -471 1914 -437
rect 1948 -471 1958 -437
rect 1906 -509 1958 -471
rect 2168 -437 2220 -399
rect 2168 -471 2178 -437
rect 2212 -471 2220 -437
rect 2168 -509 2220 -471
rect 2472 -425 2522 -379
rect 2366 -452 2420 -425
rect 2366 -486 2375 -452
rect 2409 -486 2420 -452
rect 2366 -509 2420 -486
rect 2450 -452 2522 -425
rect 2450 -486 2472 -452
rect 2506 -486 2522 -452
rect 2450 -509 2522 -486
rect 2622 -452 2674 -379
rect 2622 -486 2632 -452
rect 2666 -486 2674 -452
rect 2622 -509 2674 -486
rect 2729 -452 2782 -379
rect 2729 -486 2737 -452
rect 2771 -486 2782 -452
rect 2729 -509 2782 -486
rect 2882 -425 2932 -379
rect 2882 -452 2947 -425
rect 2882 -486 2893 -452
rect 2927 -486 2947 -452
rect 2882 -509 2947 -486
rect 2977 -452 3048 -425
rect 2977 -486 2991 -452
rect 3025 -486 3048 -452
rect 2977 -509 3048 -486
rect 3194 -437 3246 -399
rect 3194 -471 3202 -437
rect 3236 -471 3246 -437
rect 3194 -509 3246 -471
rect 3456 -437 3508 -399
rect 3456 -471 3466 -437
rect 3500 -471 3508 -437
rect 3456 -509 3508 -471
rect 4390 -444 4442 -399
rect 4390 -478 4398 -444
rect 4432 -478 4442 -444
rect 4390 -509 4442 -478
rect 5388 -444 5440 -399
rect 5388 -478 5398 -444
rect 5432 -478 5440 -444
rect 5388 -509 5440 -478
rect 6414 -437 6466 -399
rect 6414 -471 6422 -437
rect 6456 -471 6466 -437
rect 6414 -509 6466 -471
rect 6676 -437 6728 -399
rect 6676 -471 6686 -437
rect 6720 -471 6728 -437
rect 6676 -509 6728 -471
rect 6980 -425 7030 -379
rect 6874 -452 6928 -425
rect 6874 -486 6883 -452
rect 6917 -486 6928 -452
rect 6874 -509 6928 -486
rect 6958 -452 7030 -425
rect 6958 -486 6980 -452
rect 7014 -486 7030 -452
rect 6958 -509 7030 -486
rect 7130 -452 7182 -379
rect 7130 -486 7140 -452
rect 7174 -486 7182 -452
rect 7130 -509 7182 -486
rect 7237 -452 7290 -379
rect 7237 -486 7245 -452
rect 7279 -486 7290 -452
rect 7237 -509 7290 -486
rect 7390 -425 7440 -379
rect 7390 -452 7455 -425
rect 7390 -486 7401 -452
rect 7435 -486 7455 -452
rect 7390 -509 7455 -486
rect 7485 -452 7556 -425
rect 7485 -486 7499 -452
rect 7533 -486 7556 -452
rect 7485 -509 7556 -486
rect 7702 -437 7754 -399
rect 7702 -471 7710 -437
rect 7744 -471 7754 -437
rect 7702 -509 7754 -471
rect 7964 -437 8016 -399
rect 7964 -471 7974 -437
rect 8008 -471 8016 -437
rect 7964 -509 8016 -471
rect 8268 -425 8318 -379
rect 8162 -452 8216 -425
rect 8162 -486 8171 -452
rect 8205 -486 8216 -452
rect 8162 -509 8216 -486
rect 8246 -452 8318 -425
rect 8246 -486 8268 -452
rect 8302 -486 8318 -452
rect 8246 -509 8318 -486
rect 8418 -452 8470 -379
rect 8418 -486 8428 -452
rect 8462 -486 8470 -452
rect 8418 -509 8470 -486
rect 8525 -452 8578 -379
rect 8525 -486 8533 -452
rect 8567 -486 8578 -452
rect 8525 -509 8578 -486
rect 8678 -425 8728 -379
rect 8678 -452 8743 -425
rect 8678 -486 8689 -452
rect 8723 -486 8743 -452
rect 8678 -509 8743 -486
rect 8773 -452 8844 -425
rect 8773 -486 8787 -452
rect 8821 -486 8844 -452
rect 8773 -509 8844 -486
rect 8990 -437 9042 -399
rect 8990 -471 8998 -437
rect 9032 -471 9042 -437
rect 8990 -509 9042 -471
rect 9252 -437 9304 -399
rect 9252 -471 9262 -437
rect 9296 -471 9304 -437
rect 9252 -509 9304 -471
rect 9556 -425 9606 -379
rect 9450 -452 9504 -425
rect 9450 -486 9459 -452
rect 9493 -486 9504 -452
rect 9450 -509 9504 -486
rect 9534 -452 9606 -425
rect 9534 -486 9556 -452
rect 9590 -486 9606 -452
rect 9534 -509 9606 -486
rect 9706 -452 9758 -379
rect 9706 -486 9716 -452
rect 9750 -486 9758 -452
rect 9706 -509 9758 -486
rect 9813 -452 9866 -379
rect 9813 -486 9821 -452
rect 9855 -486 9866 -452
rect 9813 -509 9866 -486
rect 9966 -425 10016 -379
rect 9966 -452 10031 -425
rect 9966 -486 9977 -452
rect 10011 -486 10031 -452
rect 9966 -509 10031 -486
rect 10061 -452 10132 -425
rect 10061 -486 10075 -452
rect 10109 -486 10132 -452
rect 10061 -509 10132 -486
rect 10278 -437 10330 -399
rect 10278 -471 10286 -437
rect 10320 -471 10330 -437
rect 10278 -509 10330 -471
rect 10540 -437 10592 -399
rect 10540 -471 10550 -437
rect 10584 -471 10592 -437
rect 10540 -509 10592 -471
rect 10738 -395 10790 -379
rect 10738 -429 10746 -395
rect 10780 -429 10790 -395
rect 10738 -463 10790 -429
rect 10738 -497 10746 -463
rect 10780 -497 10790 -463
rect 10738 -509 10790 -497
rect 10820 -463 10874 -379
rect 10820 -497 10830 -463
rect 10864 -497 10874 -463
rect 10820 -509 10874 -497
rect 10904 -395 10958 -379
rect 10904 -429 10914 -395
rect 10948 -429 10958 -395
rect 10904 -463 10958 -429
rect 10904 -497 10914 -463
rect 10948 -497 10958 -463
rect 10904 -509 10958 -497
rect 10988 -463 11042 -379
rect 10988 -497 10998 -463
rect 11032 -497 11042 -463
rect 10988 -509 11042 -497
rect 11072 -395 11126 -379
rect 11072 -429 11082 -395
rect 11116 -429 11126 -395
rect 11072 -463 11126 -429
rect 11072 -497 11082 -463
rect 11116 -497 11126 -463
rect 11072 -509 11126 -497
rect 11156 -395 11210 -379
rect 11156 -429 11166 -395
rect 11200 -429 11210 -395
rect 11156 -509 11210 -429
rect 11240 -463 11294 -379
rect 11240 -497 11250 -463
rect 11284 -497 11294 -463
rect 11240 -509 11294 -497
rect 11324 -395 11378 -379
rect 11324 -429 11334 -395
rect 11368 -429 11378 -395
rect 11324 -509 11378 -429
rect 11408 -395 11460 -379
rect 11408 -429 11418 -395
rect 11452 -429 11460 -395
rect 11408 -463 11460 -429
rect 11408 -497 11418 -463
rect 11452 -497 11460 -463
rect 11658 -437 11710 -399
rect 11658 -471 11666 -437
rect 11700 -471 11710 -437
rect 11408 -509 11460 -497
rect 11658 -509 11710 -471
rect 11920 -437 11972 -399
rect 11920 -471 11930 -437
rect 11964 -471 11972 -437
rect 11920 -509 11972 -471
rect 13590 -444 13642 -399
rect 13590 -478 13598 -444
rect 13632 -478 13642 -444
rect 13590 -509 13642 -478
rect 14588 -444 14640 -399
rect 14588 -478 14598 -444
rect 14632 -478 14640 -444
rect 14588 -509 14640 -478
rect 14786 -444 14838 -399
rect 14786 -478 14794 -444
rect 14828 -478 14838 -444
rect 14786 -509 14838 -478
rect 15784 -444 15836 -399
rect 15784 -478 15794 -444
rect 15828 -478 15836 -444
rect 15784 -509 15836 -478
rect 15982 -444 16034 -399
rect 15982 -478 15990 -444
rect 16024 -478 16034 -444
rect 15982 -509 16034 -478
rect 16612 -444 16664 -399
rect 16612 -478 16622 -444
rect 16656 -478 16664 -444
rect 16612 -509 16664 -478
rect -2970 -634 -2918 -603
rect -2970 -668 -2962 -634
rect -2928 -668 -2918 -634
rect -2970 -713 -2918 -668
rect -2340 -634 -2288 -603
rect -2340 -668 -2330 -634
rect -2296 -668 -2288 -634
rect -2340 -713 -2288 -668
rect -1590 -634 -1538 -603
rect -1590 -668 -1582 -634
rect -1548 -668 -1538 -634
rect -1590 -713 -1538 -668
rect -960 -634 -908 -603
rect -960 -668 -950 -634
rect -916 -668 -908 -634
rect -960 -713 -908 -668
rect -854 -634 -802 -603
rect -854 -668 -846 -634
rect -812 -668 -802 -634
rect -854 -713 -802 -668
rect -224 -634 -172 -603
rect -224 -668 -214 -634
rect -180 -668 -172 -634
rect -224 -713 -172 -668
rect -26 -641 26 -603
rect -26 -675 -18 -641
rect 16 -675 26 -641
rect -26 -713 26 -675
rect 236 -641 288 -603
rect 236 -675 246 -641
rect 280 -675 288 -641
rect 236 -713 288 -675
rect 434 -626 505 -603
rect 434 -660 457 -626
rect 491 -660 505 -626
rect 434 -687 505 -660
rect 535 -626 600 -603
rect 535 -660 555 -626
rect 589 -660 600 -626
rect 535 -687 600 -660
rect 550 -733 600 -687
rect 700 -626 753 -603
rect 700 -660 711 -626
rect 745 -660 753 -626
rect 700 -733 753 -660
rect 808 -626 860 -603
rect 808 -660 816 -626
rect 850 -660 860 -626
rect 808 -733 860 -660
rect 960 -626 1032 -603
rect 960 -660 976 -626
rect 1010 -660 1032 -626
rect 960 -687 1032 -660
rect 1062 -626 1116 -603
rect 1062 -660 1073 -626
rect 1107 -660 1116 -626
rect 1062 -687 1116 -660
rect 960 -733 1010 -687
rect 1262 -641 1314 -603
rect 1262 -675 1270 -641
rect 1304 -675 1314 -641
rect 1262 -713 1314 -675
rect 1524 -641 1576 -603
rect 1524 -675 1534 -641
rect 1568 -675 1576 -641
rect 1524 -713 1576 -675
rect 1722 -634 1774 -603
rect 1722 -668 1730 -634
rect 1764 -668 1774 -634
rect 1722 -713 1774 -668
rect 2352 -634 2404 -603
rect 2352 -668 2362 -634
rect 2396 -668 2404 -634
rect 2352 -713 2404 -668
rect 2550 -641 2602 -603
rect 2550 -675 2558 -641
rect 2592 -675 2602 -641
rect 2550 -713 2602 -675
rect 2812 -641 2864 -603
rect 2812 -675 2822 -641
rect 2856 -675 2864 -641
rect 2812 -713 2864 -675
rect 3010 -626 3081 -603
rect 3010 -660 3033 -626
rect 3067 -660 3081 -626
rect 3010 -687 3081 -660
rect 3111 -626 3176 -603
rect 3111 -660 3131 -626
rect 3165 -660 3176 -626
rect 3111 -687 3176 -660
rect 3126 -733 3176 -687
rect 3276 -626 3329 -603
rect 3276 -660 3287 -626
rect 3321 -660 3329 -626
rect 3276 -733 3329 -660
rect 3384 -626 3436 -603
rect 3384 -660 3392 -626
rect 3426 -660 3436 -626
rect 3384 -733 3436 -660
rect 3536 -626 3608 -603
rect 3536 -660 3552 -626
rect 3586 -660 3608 -626
rect 3536 -687 3608 -660
rect 3638 -626 3692 -603
rect 3638 -660 3649 -626
rect 3683 -660 3692 -626
rect 3638 -687 3692 -660
rect 3536 -733 3586 -687
rect 3838 -641 3890 -603
rect 3838 -675 3846 -641
rect 3880 -675 3890 -641
rect 3838 -713 3890 -675
rect 4100 -641 4152 -603
rect 4100 -675 4110 -641
rect 4144 -675 4152 -641
rect 4100 -713 4152 -675
rect 4298 -634 4350 -603
rect 4298 -668 4306 -634
rect 4340 -668 4350 -634
rect 4298 -713 4350 -668
rect 4928 -634 4980 -603
rect 4928 -668 4938 -634
rect 4972 -668 4980 -634
rect 4928 -713 4980 -668
rect 5126 -641 5178 -603
rect 5126 -675 5134 -641
rect 5168 -675 5178 -641
rect 5126 -713 5178 -675
rect 5388 -641 5440 -603
rect 5388 -675 5398 -641
rect 5432 -675 5440 -641
rect 5388 -713 5440 -675
rect 5586 -626 5657 -603
rect 5586 -660 5609 -626
rect 5643 -660 5657 -626
rect 5586 -687 5657 -660
rect 5687 -626 5752 -603
rect 5687 -660 5707 -626
rect 5741 -660 5752 -626
rect 5687 -687 5752 -660
rect 5702 -733 5752 -687
rect 5852 -626 5905 -603
rect 5852 -660 5863 -626
rect 5897 -660 5905 -626
rect 5852 -733 5905 -660
rect 5960 -626 6012 -603
rect 5960 -660 5968 -626
rect 6002 -660 6012 -626
rect 5960 -733 6012 -660
rect 6112 -626 6184 -603
rect 6112 -660 6128 -626
rect 6162 -660 6184 -626
rect 6112 -687 6184 -660
rect 6214 -626 6268 -603
rect 6214 -660 6225 -626
rect 6259 -660 6268 -626
rect 6214 -687 6268 -660
rect 6112 -733 6162 -687
rect 6414 -641 6466 -603
rect 6414 -675 6422 -641
rect 6456 -675 6466 -641
rect 6414 -713 6466 -675
rect 6676 -641 6728 -603
rect 6676 -675 6686 -641
rect 6720 -675 6728 -641
rect 6676 -713 6728 -675
rect 6874 -634 6926 -603
rect 6874 -668 6882 -634
rect 6916 -668 6926 -634
rect 6874 -713 6926 -668
rect 7504 -634 7556 -603
rect 7504 -668 7514 -634
rect 7548 -668 7556 -634
rect 7504 -713 7556 -668
rect 7702 -641 7754 -603
rect 7702 -675 7710 -641
rect 7744 -675 7754 -641
rect 7702 -713 7754 -675
rect 7964 -641 8016 -603
rect 7964 -675 7974 -641
rect 8008 -675 8016 -641
rect 7964 -713 8016 -675
rect 8162 -626 8233 -603
rect 8162 -660 8185 -626
rect 8219 -660 8233 -626
rect 8162 -687 8233 -660
rect 8263 -626 8328 -603
rect 8263 -660 8283 -626
rect 8317 -660 8328 -626
rect 8263 -687 8328 -660
rect 8278 -733 8328 -687
rect 8428 -626 8481 -603
rect 8428 -660 8439 -626
rect 8473 -660 8481 -626
rect 8428 -733 8481 -660
rect 8536 -626 8588 -603
rect 8536 -660 8544 -626
rect 8578 -660 8588 -626
rect 8536 -733 8588 -660
rect 8688 -626 8760 -603
rect 8688 -660 8704 -626
rect 8738 -660 8760 -626
rect 8688 -687 8760 -660
rect 8790 -626 8844 -603
rect 8790 -660 8801 -626
rect 8835 -660 8844 -626
rect 8790 -687 8844 -660
rect 8688 -733 8738 -687
rect 8990 -641 9042 -603
rect 8990 -675 8998 -641
rect 9032 -675 9042 -641
rect 8990 -713 9042 -675
rect 9252 -641 9304 -603
rect 9252 -675 9262 -641
rect 9296 -675 9304 -641
rect 9252 -713 9304 -675
rect 9450 -634 9502 -603
rect 9450 -668 9458 -634
rect 9492 -668 9502 -634
rect 9450 -713 9502 -668
rect 10080 -634 10132 -603
rect 10080 -668 10090 -634
rect 10124 -668 10132 -634
rect 10080 -713 10132 -668
rect 10370 -641 10422 -603
rect 10370 -675 10378 -641
rect 10412 -675 10422 -641
rect 10370 -713 10422 -675
rect 10632 -641 10684 -603
rect 10632 -675 10642 -641
rect 10676 -675 10684 -641
rect 10632 -713 10684 -675
rect 10738 -626 10809 -603
rect 10738 -660 10761 -626
rect 10795 -660 10809 -626
rect 10738 -687 10809 -660
rect 10839 -626 10904 -603
rect 10839 -660 10859 -626
rect 10893 -660 10904 -626
rect 10839 -687 10904 -660
rect 10854 -733 10904 -687
rect 11004 -626 11057 -603
rect 11004 -660 11015 -626
rect 11049 -660 11057 -626
rect 11004 -733 11057 -660
rect 11112 -626 11164 -603
rect 11112 -660 11120 -626
rect 11154 -660 11164 -626
rect 11112 -733 11164 -660
rect 11264 -626 11336 -603
rect 11264 -660 11280 -626
rect 11314 -660 11336 -626
rect 11264 -687 11336 -660
rect 11366 -626 11420 -603
rect 11366 -660 11377 -626
rect 11411 -660 11420 -626
rect 11366 -687 11420 -660
rect 11264 -733 11314 -687
rect 11658 -641 11710 -603
rect 11658 -675 11666 -641
rect 11700 -675 11710 -641
rect 11658 -713 11710 -675
rect 11920 -641 11972 -603
rect 13682 -615 13735 -603
rect 11920 -675 11930 -641
rect 11964 -675 11972 -641
rect 11920 -713 11972 -675
rect 13682 -649 13690 -615
rect 13724 -649 13735 -615
rect 13682 -687 13735 -649
rect 13765 -628 13821 -603
rect 13765 -662 13776 -628
rect 13810 -662 13821 -628
rect 13765 -687 13821 -662
rect 13851 -628 13907 -603
rect 13851 -662 13862 -628
rect 13896 -662 13907 -628
rect 13851 -687 13907 -662
rect 13937 -628 13993 -603
rect 13937 -662 13948 -628
rect 13982 -662 13993 -628
rect 13937 -687 13993 -662
rect 14023 -628 14079 -603
rect 14023 -662 14034 -628
rect 14068 -662 14079 -628
rect 14023 -687 14079 -662
rect 14109 -628 14165 -603
rect 14109 -662 14120 -628
rect 14154 -662 14165 -628
rect 14109 -687 14165 -662
rect 14195 -619 14251 -603
rect 14195 -653 14206 -619
rect 14240 -653 14251 -619
rect 14195 -687 14251 -653
rect 14281 -628 14337 -603
rect 14281 -662 14292 -628
rect 14326 -662 14337 -628
rect 14281 -687 14337 -662
rect 14367 -619 14423 -603
rect 14367 -653 14378 -619
rect 14412 -653 14423 -619
rect 14367 -687 14423 -653
rect 14453 -628 14509 -603
rect 14453 -662 14464 -628
rect 14498 -662 14509 -628
rect 14453 -687 14509 -662
rect 14539 -619 14595 -603
rect 14539 -653 14550 -619
rect 14584 -653 14595 -619
rect 14539 -687 14595 -653
rect 14625 -628 14681 -603
rect 14625 -662 14636 -628
rect 14670 -662 14681 -628
rect 14625 -687 14681 -662
rect 14711 -619 14766 -603
rect 14711 -653 14722 -619
rect 14756 -653 14766 -619
rect 14711 -687 14766 -653
rect 14796 -628 14852 -603
rect 14796 -662 14807 -628
rect 14841 -662 14852 -628
rect 14796 -687 14852 -662
rect 14882 -619 14938 -603
rect 14882 -653 14893 -619
rect 14927 -653 14938 -619
rect 14882 -687 14938 -653
rect 14968 -628 15024 -603
rect 14968 -662 14979 -628
rect 15013 -662 15024 -628
rect 14968 -687 15024 -662
rect 15054 -619 15110 -603
rect 15054 -653 15065 -619
rect 15099 -653 15110 -619
rect 15054 -687 15110 -653
rect 15140 -628 15196 -603
rect 15140 -662 15151 -628
rect 15185 -662 15196 -628
rect 15140 -687 15196 -662
rect 15226 -619 15282 -603
rect 15226 -653 15237 -619
rect 15271 -653 15282 -619
rect 15226 -687 15282 -653
rect 15312 -628 15368 -603
rect 15312 -662 15323 -628
rect 15357 -662 15368 -628
rect 15312 -687 15368 -662
rect 15398 -619 15451 -603
rect 15398 -653 15409 -619
rect 15443 -653 15451 -619
rect 15398 -687 15451 -653
rect 15614 -634 15666 -603
rect 15614 -668 15622 -634
rect 15656 -668 15666 -634
rect 15614 -713 15666 -668
rect 16612 -634 16664 -603
rect 16612 -668 16622 -634
rect 16656 -668 16664 -634
rect 16612 -713 16664 -668
rect -2970 -1532 -2918 -1487
rect -2970 -1566 -2962 -1532
rect -2928 -1566 -2918 -1532
rect -2970 -1597 -2918 -1566
rect -2340 -1532 -2288 -1487
rect -2340 -1566 -2330 -1532
rect -2296 -1566 -2288 -1532
rect -2340 -1597 -2288 -1566
rect -1590 -1532 -1538 -1487
rect -1590 -1566 -1582 -1532
rect -1548 -1566 -1538 -1532
rect -1590 -1597 -1538 -1566
rect -960 -1532 -908 -1487
rect -960 -1566 -950 -1532
rect -916 -1566 -908 -1532
rect -960 -1597 -908 -1566
rect -854 -1532 -802 -1487
rect -854 -1566 -846 -1532
rect -812 -1566 -802 -1532
rect -854 -1597 -802 -1566
rect -224 -1532 -172 -1487
rect -224 -1566 -214 -1532
rect -180 -1566 -172 -1532
rect -224 -1597 -172 -1566
rect -26 -1525 26 -1487
rect -26 -1559 -18 -1525
rect 16 -1559 26 -1525
rect -26 -1597 26 -1559
rect 236 -1525 288 -1487
rect 236 -1559 246 -1525
rect 280 -1559 288 -1525
rect 236 -1597 288 -1559
rect 540 -1513 590 -1467
rect 434 -1540 488 -1513
rect 434 -1574 443 -1540
rect 477 -1574 488 -1540
rect 434 -1597 488 -1574
rect 518 -1540 590 -1513
rect 518 -1574 540 -1540
rect 574 -1574 590 -1540
rect 518 -1597 590 -1574
rect 690 -1540 742 -1467
rect 690 -1574 700 -1540
rect 734 -1574 742 -1540
rect 690 -1597 742 -1574
rect 797 -1540 850 -1467
rect 797 -1574 805 -1540
rect 839 -1574 850 -1540
rect 797 -1597 850 -1574
rect 950 -1513 1000 -1467
rect 950 -1540 1015 -1513
rect 950 -1574 961 -1540
rect 995 -1574 1015 -1540
rect 950 -1597 1015 -1574
rect 1045 -1540 1116 -1513
rect 1045 -1574 1059 -1540
rect 1093 -1574 1116 -1540
rect 1045 -1597 1116 -1574
rect 1262 -1525 1314 -1487
rect 1262 -1559 1270 -1525
rect 1304 -1559 1314 -1525
rect 1262 -1597 1314 -1559
rect 1524 -1525 1576 -1487
rect 1524 -1559 1534 -1525
rect 1568 -1559 1576 -1525
rect 1524 -1597 1576 -1559
rect 1722 -1532 1774 -1487
rect 1722 -1566 1730 -1532
rect 1764 -1566 1774 -1532
rect 1722 -1597 1774 -1566
rect 2352 -1532 2404 -1487
rect 2352 -1566 2362 -1532
rect 2396 -1566 2404 -1532
rect 2352 -1597 2404 -1566
rect 2550 -1525 2602 -1487
rect 2550 -1559 2558 -1525
rect 2592 -1559 2602 -1525
rect 2550 -1597 2602 -1559
rect 2812 -1525 2864 -1487
rect 2812 -1559 2822 -1525
rect 2856 -1559 2864 -1525
rect 2812 -1597 2864 -1559
rect 3116 -1513 3166 -1467
rect 3010 -1540 3064 -1513
rect 3010 -1574 3019 -1540
rect 3053 -1574 3064 -1540
rect 3010 -1597 3064 -1574
rect 3094 -1540 3166 -1513
rect 3094 -1574 3116 -1540
rect 3150 -1574 3166 -1540
rect 3094 -1597 3166 -1574
rect 3266 -1540 3318 -1467
rect 3266 -1574 3276 -1540
rect 3310 -1574 3318 -1540
rect 3266 -1597 3318 -1574
rect 3373 -1540 3426 -1467
rect 3373 -1574 3381 -1540
rect 3415 -1574 3426 -1540
rect 3373 -1597 3426 -1574
rect 3526 -1513 3576 -1467
rect 3526 -1540 3591 -1513
rect 3526 -1574 3537 -1540
rect 3571 -1574 3591 -1540
rect 3526 -1597 3591 -1574
rect 3621 -1540 3692 -1513
rect 3621 -1574 3635 -1540
rect 3669 -1574 3692 -1540
rect 3621 -1597 3692 -1574
rect 3838 -1525 3890 -1487
rect 3838 -1559 3846 -1525
rect 3880 -1559 3890 -1525
rect 3838 -1597 3890 -1559
rect 4100 -1525 4152 -1487
rect 4100 -1559 4110 -1525
rect 4144 -1559 4152 -1525
rect 4100 -1597 4152 -1559
rect 4298 -1532 4350 -1487
rect 4298 -1566 4306 -1532
rect 4340 -1566 4350 -1532
rect 4298 -1597 4350 -1566
rect 4928 -1532 4980 -1487
rect 4928 -1566 4938 -1532
rect 4972 -1566 4980 -1532
rect 4928 -1597 4980 -1566
rect 5126 -1525 5178 -1487
rect 5126 -1559 5134 -1525
rect 5168 -1559 5178 -1525
rect 5126 -1597 5178 -1559
rect 5388 -1525 5440 -1487
rect 5388 -1559 5398 -1525
rect 5432 -1559 5440 -1525
rect 5388 -1597 5440 -1559
rect 5692 -1513 5742 -1467
rect 5586 -1540 5640 -1513
rect 5586 -1574 5595 -1540
rect 5629 -1574 5640 -1540
rect 5586 -1597 5640 -1574
rect 5670 -1540 5742 -1513
rect 5670 -1574 5692 -1540
rect 5726 -1574 5742 -1540
rect 5670 -1597 5742 -1574
rect 5842 -1540 5894 -1467
rect 5842 -1574 5852 -1540
rect 5886 -1574 5894 -1540
rect 5842 -1597 5894 -1574
rect 5949 -1540 6002 -1467
rect 5949 -1574 5957 -1540
rect 5991 -1574 6002 -1540
rect 5949 -1597 6002 -1574
rect 6102 -1513 6152 -1467
rect 6102 -1540 6167 -1513
rect 6102 -1574 6113 -1540
rect 6147 -1574 6167 -1540
rect 6102 -1597 6167 -1574
rect 6197 -1540 6268 -1513
rect 6197 -1574 6211 -1540
rect 6245 -1574 6268 -1540
rect 6197 -1597 6268 -1574
rect 6414 -1525 6466 -1487
rect 6414 -1559 6422 -1525
rect 6456 -1559 6466 -1525
rect 6414 -1597 6466 -1559
rect 6676 -1525 6728 -1487
rect 6676 -1559 6686 -1525
rect 6720 -1559 6728 -1525
rect 6676 -1597 6728 -1559
rect 6874 -1532 6926 -1487
rect 6874 -1566 6882 -1532
rect 6916 -1566 6926 -1532
rect 6874 -1597 6926 -1566
rect 7504 -1532 7556 -1487
rect 7504 -1566 7514 -1532
rect 7548 -1566 7556 -1532
rect 7504 -1597 7556 -1566
rect 7702 -1525 7754 -1487
rect 7702 -1559 7710 -1525
rect 7744 -1559 7754 -1525
rect 7702 -1597 7754 -1559
rect 7964 -1525 8016 -1487
rect 7964 -1559 7974 -1525
rect 8008 -1559 8016 -1525
rect 7964 -1597 8016 -1559
rect 8268 -1513 8318 -1467
rect 8162 -1540 8216 -1513
rect 8162 -1574 8171 -1540
rect 8205 -1574 8216 -1540
rect 8162 -1597 8216 -1574
rect 8246 -1540 8318 -1513
rect 8246 -1574 8268 -1540
rect 8302 -1574 8318 -1540
rect 8246 -1597 8318 -1574
rect 8418 -1540 8470 -1467
rect 8418 -1574 8428 -1540
rect 8462 -1574 8470 -1540
rect 8418 -1597 8470 -1574
rect 8525 -1540 8578 -1467
rect 8525 -1574 8533 -1540
rect 8567 -1574 8578 -1540
rect 8525 -1597 8578 -1574
rect 8678 -1513 8728 -1467
rect 8678 -1540 8743 -1513
rect 8678 -1574 8689 -1540
rect 8723 -1574 8743 -1540
rect 8678 -1597 8743 -1574
rect 8773 -1540 8844 -1513
rect 8773 -1574 8787 -1540
rect 8821 -1574 8844 -1540
rect 8773 -1597 8844 -1574
rect 8990 -1525 9042 -1487
rect 8990 -1559 8998 -1525
rect 9032 -1559 9042 -1525
rect 8990 -1597 9042 -1559
rect 9252 -1525 9304 -1487
rect 9252 -1559 9262 -1525
rect 9296 -1559 9304 -1525
rect 9252 -1597 9304 -1559
rect 9450 -1532 9502 -1487
rect 9450 -1566 9458 -1532
rect 9492 -1566 9502 -1532
rect 9450 -1597 9502 -1566
rect 10080 -1532 10132 -1487
rect 10080 -1566 10090 -1532
rect 10124 -1566 10132 -1532
rect 10080 -1597 10132 -1566
rect 10370 -1525 10422 -1487
rect 10370 -1559 10378 -1525
rect 10412 -1559 10422 -1525
rect 10370 -1597 10422 -1559
rect 10632 -1525 10684 -1487
rect 10844 -1513 10894 -1467
rect 10632 -1559 10642 -1525
rect 10676 -1559 10684 -1525
rect 10632 -1597 10684 -1559
rect 10738 -1540 10792 -1513
rect 10738 -1574 10747 -1540
rect 10781 -1574 10792 -1540
rect 10738 -1597 10792 -1574
rect 10822 -1540 10894 -1513
rect 10822 -1574 10844 -1540
rect 10878 -1574 10894 -1540
rect 10822 -1597 10894 -1574
rect 10994 -1540 11046 -1467
rect 10994 -1574 11004 -1540
rect 11038 -1574 11046 -1540
rect 10994 -1597 11046 -1574
rect 11101 -1540 11154 -1467
rect 11101 -1574 11109 -1540
rect 11143 -1574 11154 -1540
rect 11101 -1597 11154 -1574
rect 11254 -1513 11304 -1467
rect 11254 -1540 11319 -1513
rect 11254 -1574 11265 -1540
rect 11299 -1574 11319 -1540
rect 11254 -1597 11319 -1574
rect 11349 -1540 11420 -1513
rect 11349 -1574 11363 -1540
rect 11397 -1574 11420 -1540
rect 11349 -1597 11420 -1574
rect 11658 -1525 11710 -1487
rect 11658 -1559 11666 -1525
rect 11700 -1559 11710 -1525
rect 11658 -1597 11710 -1559
rect 11920 -1525 11972 -1487
rect 11920 -1559 11930 -1525
rect 11964 -1559 11972 -1525
rect 11920 -1597 11972 -1559
rect 12567 -1549 12633 -1513
rect 12567 -1583 12588 -1549
rect 12622 -1583 12633 -1549
rect 12567 -1597 12633 -1583
rect 12663 -1538 12719 -1513
rect 12663 -1572 12674 -1538
rect 12708 -1572 12719 -1538
rect 12663 -1597 12719 -1572
rect 12749 -1549 12805 -1513
rect 12749 -1583 12760 -1549
rect 12794 -1583 12805 -1549
rect 12749 -1597 12805 -1583
rect 12835 -1538 12891 -1513
rect 12835 -1572 12846 -1538
rect 12880 -1572 12891 -1538
rect 12835 -1597 12891 -1572
rect 12921 -1549 13000 -1513
rect 12921 -1583 12932 -1549
rect 12966 -1583 13000 -1549
rect 13222 -1525 13274 -1487
rect 13222 -1559 13230 -1525
rect 13264 -1559 13274 -1525
rect 12921 -1597 13000 -1583
rect 13222 -1597 13274 -1559
rect 13484 -1525 13536 -1487
rect 13484 -1559 13494 -1525
rect 13528 -1559 13536 -1525
rect 13484 -1597 13536 -1559
rect 13682 -1551 13735 -1513
rect 13682 -1585 13690 -1551
rect 13724 -1585 13735 -1551
rect 13682 -1597 13735 -1585
rect 13765 -1538 13821 -1513
rect 13765 -1572 13776 -1538
rect 13810 -1572 13821 -1538
rect 13765 -1597 13821 -1572
rect 13851 -1538 13907 -1513
rect 13851 -1572 13862 -1538
rect 13896 -1572 13907 -1538
rect 13851 -1597 13907 -1572
rect 13937 -1538 13993 -1513
rect 13937 -1572 13948 -1538
rect 13982 -1572 13993 -1538
rect 13937 -1597 13993 -1572
rect 14023 -1538 14079 -1513
rect 14023 -1572 14034 -1538
rect 14068 -1572 14079 -1538
rect 14023 -1597 14079 -1572
rect 14109 -1538 14165 -1513
rect 14109 -1572 14120 -1538
rect 14154 -1572 14165 -1538
rect 14109 -1597 14165 -1572
rect 14195 -1547 14251 -1513
rect 14195 -1581 14206 -1547
rect 14240 -1581 14251 -1547
rect 14195 -1597 14251 -1581
rect 14281 -1538 14337 -1513
rect 14281 -1572 14292 -1538
rect 14326 -1572 14337 -1538
rect 14281 -1597 14337 -1572
rect 14367 -1547 14423 -1513
rect 14367 -1581 14378 -1547
rect 14412 -1581 14423 -1547
rect 14367 -1597 14423 -1581
rect 14453 -1538 14509 -1513
rect 14453 -1572 14464 -1538
rect 14498 -1572 14509 -1538
rect 14453 -1597 14509 -1572
rect 14539 -1547 14595 -1513
rect 14539 -1581 14550 -1547
rect 14584 -1581 14595 -1547
rect 14539 -1597 14595 -1581
rect 14625 -1538 14681 -1513
rect 14625 -1572 14636 -1538
rect 14670 -1572 14681 -1538
rect 14625 -1597 14681 -1572
rect 14711 -1547 14766 -1513
rect 14711 -1581 14722 -1547
rect 14756 -1581 14766 -1547
rect 14711 -1597 14766 -1581
rect 14796 -1538 14852 -1513
rect 14796 -1572 14807 -1538
rect 14841 -1572 14852 -1538
rect 14796 -1597 14852 -1572
rect 14882 -1547 14938 -1513
rect 14882 -1581 14893 -1547
rect 14927 -1581 14938 -1547
rect 14882 -1597 14938 -1581
rect 14968 -1538 15024 -1513
rect 14968 -1572 14979 -1538
rect 15013 -1572 15024 -1538
rect 14968 -1597 15024 -1572
rect 15054 -1547 15110 -1513
rect 15054 -1581 15065 -1547
rect 15099 -1581 15110 -1547
rect 15054 -1597 15110 -1581
rect 15140 -1538 15196 -1513
rect 15140 -1572 15151 -1538
rect 15185 -1572 15196 -1538
rect 15140 -1597 15196 -1572
rect 15226 -1547 15282 -1513
rect 15226 -1581 15237 -1547
rect 15271 -1581 15282 -1547
rect 15226 -1597 15282 -1581
rect 15312 -1538 15368 -1513
rect 15312 -1572 15323 -1538
rect 15357 -1572 15368 -1538
rect 15312 -1597 15368 -1572
rect 15398 -1547 15451 -1513
rect 15398 -1581 15409 -1547
rect 15443 -1581 15451 -1547
rect 15614 -1532 15666 -1487
rect 15614 -1566 15622 -1532
rect 15656 -1566 15666 -1532
rect 15398 -1597 15451 -1581
rect 15614 -1597 15666 -1566
rect 16612 -1532 16664 -1487
rect 16612 -1566 16622 -1532
rect 16656 -1566 16664 -1532
rect 16612 -1597 16664 -1566
rect -2970 -1722 -2918 -1691
rect -2970 -1756 -2962 -1722
rect -2928 -1756 -2918 -1722
rect -2970 -1801 -2918 -1756
rect -2340 -1722 -2288 -1691
rect -2340 -1756 -2330 -1722
rect -2296 -1756 -2288 -1722
rect -2340 -1801 -2288 -1756
rect -1590 -1722 -1538 -1691
rect -1590 -1756 -1582 -1722
rect -1548 -1756 -1538 -1722
rect -1590 -1801 -1538 -1756
rect -960 -1722 -908 -1691
rect -960 -1756 -950 -1722
rect -916 -1756 -908 -1722
rect -960 -1801 -908 -1756
rect -854 -1714 -783 -1691
rect -854 -1748 -831 -1714
rect -797 -1748 -783 -1714
rect -854 -1775 -783 -1748
rect -753 -1714 -688 -1691
rect -753 -1748 -733 -1714
rect -699 -1748 -688 -1714
rect -753 -1775 -688 -1748
rect -738 -1821 -688 -1775
rect -588 -1714 -535 -1691
rect -588 -1748 -577 -1714
rect -543 -1748 -535 -1714
rect -588 -1821 -535 -1748
rect -480 -1714 -428 -1691
rect -480 -1748 -472 -1714
rect -438 -1748 -428 -1714
rect -480 -1821 -428 -1748
rect -328 -1714 -256 -1691
rect -328 -1748 -312 -1714
rect -278 -1748 -256 -1714
rect -328 -1775 -256 -1748
rect -226 -1714 -172 -1691
rect -226 -1748 -215 -1714
rect -181 -1748 -172 -1714
rect -226 -1775 -172 -1748
rect -328 -1821 -278 -1775
rect -26 -1729 26 -1691
rect -26 -1763 -18 -1729
rect 16 -1763 26 -1729
rect -26 -1801 26 -1763
rect 236 -1729 288 -1691
rect 236 -1763 246 -1729
rect 280 -1763 288 -1729
rect 236 -1801 288 -1763
rect 434 -1714 505 -1691
rect 434 -1748 457 -1714
rect 491 -1748 505 -1714
rect 434 -1775 505 -1748
rect 535 -1714 600 -1691
rect 535 -1748 555 -1714
rect 589 -1748 600 -1714
rect 535 -1775 600 -1748
rect 550 -1821 600 -1775
rect 700 -1714 753 -1691
rect 700 -1748 711 -1714
rect 745 -1748 753 -1714
rect 700 -1821 753 -1748
rect 808 -1714 860 -1691
rect 808 -1748 816 -1714
rect 850 -1748 860 -1714
rect 808 -1821 860 -1748
rect 960 -1714 1032 -1691
rect 960 -1748 976 -1714
rect 1010 -1748 1032 -1714
rect 960 -1775 1032 -1748
rect 1062 -1714 1116 -1691
rect 1062 -1748 1073 -1714
rect 1107 -1748 1116 -1714
rect 1062 -1775 1116 -1748
rect 960 -1821 1010 -1775
rect 1262 -1729 1314 -1691
rect 1262 -1763 1270 -1729
rect 1304 -1763 1314 -1729
rect 1262 -1801 1314 -1763
rect 1524 -1729 1576 -1691
rect 1524 -1763 1534 -1729
rect 1568 -1763 1576 -1729
rect 1524 -1801 1576 -1763
rect 1722 -1722 1774 -1691
rect 1722 -1756 1730 -1722
rect 1764 -1756 1774 -1722
rect 1722 -1801 1774 -1756
rect 2352 -1722 2404 -1691
rect 2352 -1756 2362 -1722
rect 2396 -1756 2404 -1722
rect 2352 -1801 2404 -1756
rect 2550 -1729 2602 -1691
rect 2550 -1763 2558 -1729
rect 2592 -1763 2602 -1729
rect 2550 -1801 2602 -1763
rect 2812 -1729 2864 -1691
rect 2812 -1763 2822 -1729
rect 2856 -1763 2864 -1729
rect 2812 -1801 2864 -1763
rect 3010 -1714 3081 -1691
rect 3010 -1748 3033 -1714
rect 3067 -1748 3081 -1714
rect 3010 -1775 3081 -1748
rect 3111 -1714 3176 -1691
rect 3111 -1748 3131 -1714
rect 3165 -1748 3176 -1714
rect 3111 -1775 3176 -1748
rect 3126 -1821 3176 -1775
rect 3276 -1714 3329 -1691
rect 3276 -1748 3287 -1714
rect 3321 -1748 3329 -1714
rect 3276 -1821 3329 -1748
rect 3384 -1714 3436 -1691
rect 3384 -1748 3392 -1714
rect 3426 -1748 3436 -1714
rect 3384 -1821 3436 -1748
rect 3536 -1714 3608 -1691
rect 3536 -1748 3552 -1714
rect 3586 -1748 3608 -1714
rect 3536 -1775 3608 -1748
rect 3638 -1714 3692 -1691
rect 3638 -1748 3649 -1714
rect 3683 -1748 3692 -1714
rect 3638 -1775 3692 -1748
rect 3536 -1821 3586 -1775
rect 3838 -1729 3890 -1691
rect 3838 -1763 3846 -1729
rect 3880 -1763 3890 -1729
rect 3838 -1801 3890 -1763
rect 4100 -1729 4152 -1691
rect 4100 -1763 4110 -1729
rect 4144 -1763 4152 -1729
rect 4100 -1801 4152 -1763
rect 4298 -1722 4350 -1691
rect 4298 -1756 4306 -1722
rect 4340 -1756 4350 -1722
rect 4298 -1801 4350 -1756
rect 4928 -1722 4980 -1691
rect 4928 -1756 4938 -1722
rect 4972 -1756 4980 -1722
rect 4928 -1801 4980 -1756
rect 5126 -1729 5178 -1691
rect 5126 -1763 5134 -1729
rect 5168 -1763 5178 -1729
rect 5126 -1801 5178 -1763
rect 5388 -1729 5440 -1691
rect 5388 -1763 5398 -1729
rect 5432 -1763 5440 -1729
rect 5388 -1801 5440 -1763
rect 5586 -1714 5657 -1691
rect 5586 -1748 5609 -1714
rect 5643 -1748 5657 -1714
rect 5586 -1775 5657 -1748
rect 5687 -1714 5752 -1691
rect 5687 -1748 5707 -1714
rect 5741 -1748 5752 -1714
rect 5687 -1775 5752 -1748
rect 5702 -1821 5752 -1775
rect 5852 -1714 5905 -1691
rect 5852 -1748 5863 -1714
rect 5897 -1748 5905 -1714
rect 5852 -1821 5905 -1748
rect 5960 -1714 6012 -1691
rect 5960 -1748 5968 -1714
rect 6002 -1748 6012 -1714
rect 5960 -1821 6012 -1748
rect 6112 -1714 6184 -1691
rect 6112 -1748 6128 -1714
rect 6162 -1748 6184 -1714
rect 6112 -1775 6184 -1748
rect 6214 -1714 6268 -1691
rect 6214 -1748 6225 -1714
rect 6259 -1748 6268 -1714
rect 6214 -1775 6268 -1748
rect 6112 -1821 6162 -1775
rect 6414 -1729 6466 -1691
rect 6414 -1763 6422 -1729
rect 6456 -1763 6466 -1729
rect 6414 -1801 6466 -1763
rect 6676 -1729 6728 -1691
rect 6676 -1763 6686 -1729
rect 6720 -1763 6728 -1729
rect 6676 -1801 6728 -1763
rect 6874 -1722 6926 -1691
rect 6874 -1756 6882 -1722
rect 6916 -1756 6926 -1722
rect 6874 -1801 6926 -1756
rect 7504 -1722 7556 -1691
rect 7504 -1756 7514 -1722
rect 7548 -1756 7556 -1722
rect 7504 -1801 7556 -1756
rect 7702 -1729 7754 -1691
rect 7702 -1763 7710 -1729
rect 7744 -1763 7754 -1729
rect 7702 -1801 7754 -1763
rect 7964 -1729 8016 -1691
rect 7964 -1763 7974 -1729
rect 8008 -1763 8016 -1729
rect 7964 -1801 8016 -1763
rect 8162 -1714 8233 -1691
rect 8162 -1748 8185 -1714
rect 8219 -1748 8233 -1714
rect 8162 -1775 8233 -1748
rect 8263 -1714 8328 -1691
rect 8263 -1748 8283 -1714
rect 8317 -1748 8328 -1714
rect 8263 -1775 8328 -1748
rect 8278 -1821 8328 -1775
rect 8428 -1714 8481 -1691
rect 8428 -1748 8439 -1714
rect 8473 -1748 8481 -1714
rect 8428 -1821 8481 -1748
rect 8536 -1714 8588 -1691
rect 8536 -1748 8544 -1714
rect 8578 -1748 8588 -1714
rect 8536 -1821 8588 -1748
rect 8688 -1714 8760 -1691
rect 8688 -1748 8704 -1714
rect 8738 -1748 8760 -1714
rect 8688 -1775 8760 -1748
rect 8790 -1714 8844 -1691
rect 8790 -1748 8801 -1714
rect 8835 -1748 8844 -1714
rect 8790 -1775 8844 -1748
rect 8688 -1821 8738 -1775
rect 8990 -1729 9042 -1691
rect 8990 -1763 8998 -1729
rect 9032 -1763 9042 -1729
rect 8990 -1801 9042 -1763
rect 9252 -1729 9304 -1691
rect 9252 -1763 9262 -1729
rect 9296 -1763 9304 -1729
rect 9252 -1801 9304 -1763
rect 9450 -1722 9502 -1691
rect 9450 -1756 9458 -1722
rect 9492 -1756 9502 -1722
rect 9450 -1801 9502 -1756
rect 10080 -1722 10132 -1691
rect 10080 -1756 10090 -1722
rect 10124 -1756 10132 -1722
rect 10080 -1801 10132 -1756
rect 10370 -1729 10422 -1691
rect 10370 -1763 10378 -1729
rect 10412 -1763 10422 -1729
rect 10370 -1801 10422 -1763
rect 10632 -1729 10684 -1691
rect 10632 -1763 10642 -1729
rect 10676 -1763 10684 -1729
rect 10632 -1801 10684 -1763
rect 10738 -1714 10809 -1691
rect 10738 -1748 10761 -1714
rect 10795 -1748 10809 -1714
rect 10738 -1775 10809 -1748
rect 10839 -1714 10904 -1691
rect 10839 -1748 10859 -1714
rect 10893 -1748 10904 -1714
rect 10839 -1775 10904 -1748
rect 10854 -1821 10904 -1775
rect 11004 -1714 11057 -1691
rect 11004 -1748 11015 -1714
rect 11049 -1748 11057 -1714
rect 11004 -1821 11057 -1748
rect 11112 -1714 11164 -1691
rect 11112 -1748 11120 -1714
rect 11154 -1748 11164 -1714
rect 11112 -1821 11164 -1748
rect 11264 -1714 11336 -1691
rect 11264 -1748 11280 -1714
rect 11314 -1748 11336 -1714
rect 11264 -1775 11336 -1748
rect 11366 -1714 11420 -1691
rect 11366 -1748 11377 -1714
rect 11411 -1748 11420 -1714
rect 11366 -1775 11420 -1748
rect 11264 -1821 11314 -1775
rect 11658 -1729 11710 -1691
rect 11658 -1763 11666 -1729
rect 11700 -1763 11710 -1729
rect 11658 -1801 11710 -1763
rect 11920 -1729 11972 -1691
rect 13682 -1703 13735 -1691
rect 11920 -1763 11930 -1729
rect 11964 -1763 11972 -1729
rect 11920 -1801 11972 -1763
rect 13682 -1737 13690 -1703
rect 13724 -1737 13735 -1703
rect 13682 -1775 13735 -1737
rect 13765 -1716 13821 -1691
rect 13765 -1750 13776 -1716
rect 13810 -1750 13821 -1716
rect 13765 -1775 13821 -1750
rect 13851 -1716 13907 -1691
rect 13851 -1750 13862 -1716
rect 13896 -1750 13907 -1716
rect 13851 -1775 13907 -1750
rect 13937 -1716 13993 -1691
rect 13937 -1750 13948 -1716
rect 13982 -1750 13993 -1716
rect 13937 -1775 13993 -1750
rect 14023 -1716 14079 -1691
rect 14023 -1750 14034 -1716
rect 14068 -1750 14079 -1716
rect 14023 -1775 14079 -1750
rect 14109 -1716 14165 -1691
rect 14109 -1750 14120 -1716
rect 14154 -1750 14165 -1716
rect 14109 -1775 14165 -1750
rect 14195 -1707 14251 -1691
rect 14195 -1741 14206 -1707
rect 14240 -1741 14251 -1707
rect 14195 -1775 14251 -1741
rect 14281 -1716 14337 -1691
rect 14281 -1750 14292 -1716
rect 14326 -1750 14337 -1716
rect 14281 -1775 14337 -1750
rect 14367 -1707 14423 -1691
rect 14367 -1741 14378 -1707
rect 14412 -1741 14423 -1707
rect 14367 -1775 14423 -1741
rect 14453 -1716 14509 -1691
rect 14453 -1750 14464 -1716
rect 14498 -1750 14509 -1716
rect 14453 -1775 14509 -1750
rect 14539 -1707 14595 -1691
rect 14539 -1741 14550 -1707
rect 14584 -1741 14595 -1707
rect 14539 -1775 14595 -1741
rect 14625 -1716 14681 -1691
rect 14625 -1750 14636 -1716
rect 14670 -1750 14681 -1716
rect 14625 -1775 14681 -1750
rect 14711 -1707 14766 -1691
rect 14711 -1741 14722 -1707
rect 14756 -1741 14766 -1707
rect 14711 -1775 14766 -1741
rect 14796 -1716 14852 -1691
rect 14796 -1750 14807 -1716
rect 14841 -1750 14852 -1716
rect 14796 -1775 14852 -1750
rect 14882 -1707 14938 -1691
rect 14882 -1741 14893 -1707
rect 14927 -1741 14938 -1707
rect 14882 -1775 14938 -1741
rect 14968 -1716 15024 -1691
rect 14968 -1750 14979 -1716
rect 15013 -1750 15024 -1716
rect 14968 -1775 15024 -1750
rect 15054 -1707 15110 -1691
rect 15054 -1741 15065 -1707
rect 15099 -1741 15110 -1707
rect 15054 -1775 15110 -1741
rect 15140 -1716 15196 -1691
rect 15140 -1750 15151 -1716
rect 15185 -1750 15196 -1716
rect 15140 -1775 15196 -1750
rect 15226 -1707 15282 -1691
rect 15226 -1741 15237 -1707
rect 15271 -1741 15282 -1707
rect 15226 -1775 15282 -1741
rect 15312 -1716 15368 -1691
rect 15312 -1750 15323 -1716
rect 15357 -1750 15368 -1716
rect 15312 -1775 15368 -1750
rect 15398 -1707 15451 -1691
rect 15398 -1741 15409 -1707
rect 15443 -1741 15451 -1707
rect 15398 -1775 15451 -1741
rect 15614 -1722 15666 -1691
rect 15614 -1756 15622 -1722
rect 15656 -1756 15666 -1722
rect 15614 -1801 15666 -1756
rect 16612 -1722 16664 -1691
rect 16612 -1756 16622 -1722
rect 16656 -1756 16664 -1722
rect 16612 -1801 16664 -1756
rect -2970 -2620 -2918 -2575
rect -2970 -2654 -2962 -2620
rect -2928 -2654 -2918 -2620
rect -2970 -2685 -2918 -2654
rect -2340 -2620 -2288 -2575
rect -2340 -2654 -2330 -2620
rect -2296 -2654 -2288 -2620
rect -2340 -2685 -2288 -2654
rect -1590 -2620 -1538 -2575
rect -1590 -2654 -1582 -2620
rect -1548 -2654 -1538 -2620
rect -1590 -2685 -1538 -2654
rect -960 -2620 -908 -2575
rect -960 -2654 -950 -2620
rect -916 -2654 -908 -2620
rect -960 -2685 -908 -2654
rect -854 -2620 -802 -2575
rect -854 -2654 -846 -2620
rect -812 -2654 -802 -2620
rect -854 -2685 -802 -2654
rect -224 -2620 -172 -2575
rect -224 -2654 -214 -2620
rect -180 -2654 -172 -2620
rect -224 -2685 -172 -2654
rect -26 -2613 26 -2575
rect -26 -2647 -18 -2613
rect 16 -2647 26 -2613
rect -26 -2685 26 -2647
rect 236 -2613 288 -2575
rect 236 -2647 246 -2613
rect 280 -2647 288 -2613
rect 236 -2685 288 -2647
rect 540 -2601 590 -2555
rect 434 -2628 488 -2601
rect 434 -2662 443 -2628
rect 477 -2662 488 -2628
rect 434 -2685 488 -2662
rect 518 -2628 590 -2601
rect 518 -2662 540 -2628
rect 574 -2662 590 -2628
rect 518 -2685 590 -2662
rect 690 -2628 742 -2555
rect 690 -2662 700 -2628
rect 734 -2662 742 -2628
rect 690 -2685 742 -2662
rect 797 -2628 850 -2555
rect 797 -2662 805 -2628
rect 839 -2662 850 -2628
rect 797 -2685 850 -2662
rect 950 -2601 1000 -2555
rect 950 -2628 1015 -2601
rect 950 -2662 961 -2628
rect 995 -2662 1015 -2628
rect 950 -2685 1015 -2662
rect 1045 -2628 1116 -2601
rect 1045 -2662 1059 -2628
rect 1093 -2662 1116 -2628
rect 1045 -2685 1116 -2662
rect 1262 -2613 1314 -2575
rect 1262 -2647 1270 -2613
rect 1304 -2647 1314 -2613
rect 1262 -2685 1314 -2647
rect 1524 -2613 1576 -2575
rect 1524 -2647 1534 -2613
rect 1568 -2647 1576 -2613
rect 1524 -2685 1576 -2647
rect 1722 -2620 1774 -2575
rect 1722 -2654 1730 -2620
rect 1764 -2654 1774 -2620
rect 1722 -2685 1774 -2654
rect 2352 -2620 2404 -2575
rect 2352 -2654 2362 -2620
rect 2396 -2654 2404 -2620
rect 2352 -2685 2404 -2654
rect 2550 -2613 2602 -2575
rect 2550 -2647 2558 -2613
rect 2592 -2647 2602 -2613
rect 2550 -2685 2602 -2647
rect 2812 -2613 2864 -2575
rect 2812 -2647 2822 -2613
rect 2856 -2647 2864 -2613
rect 2812 -2685 2864 -2647
rect 3116 -2601 3166 -2555
rect 3010 -2628 3064 -2601
rect 3010 -2662 3019 -2628
rect 3053 -2662 3064 -2628
rect 3010 -2685 3064 -2662
rect 3094 -2628 3166 -2601
rect 3094 -2662 3116 -2628
rect 3150 -2662 3166 -2628
rect 3094 -2685 3166 -2662
rect 3266 -2628 3318 -2555
rect 3266 -2662 3276 -2628
rect 3310 -2662 3318 -2628
rect 3266 -2685 3318 -2662
rect 3373 -2628 3426 -2555
rect 3373 -2662 3381 -2628
rect 3415 -2662 3426 -2628
rect 3373 -2685 3426 -2662
rect 3526 -2601 3576 -2555
rect 3526 -2628 3591 -2601
rect 3526 -2662 3537 -2628
rect 3571 -2662 3591 -2628
rect 3526 -2685 3591 -2662
rect 3621 -2628 3692 -2601
rect 3621 -2662 3635 -2628
rect 3669 -2662 3692 -2628
rect 3621 -2685 3692 -2662
rect 3838 -2613 3890 -2575
rect 3838 -2647 3846 -2613
rect 3880 -2647 3890 -2613
rect 3838 -2685 3890 -2647
rect 4100 -2613 4152 -2575
rect 4100 -2647 4110 -2613
rect 4144 -2647 4152 -2613
rect 4100 -2685 4152 -2647
rect 4298 -2620 4350 -2575
rect 4298 -2654 4306 -2620
rect 4340 -2654 4350 -2620
rect 4298 -2685 4350 -2654
rect 4928 -2620 4980 -2575
rect 4928 -2654 4938 -2620
rect 4972 -2654 4980 -2620
rect 4928 -2685 4980 -2654
rect 5126 -2613 5178 -2575
rect 5126 -2647 5134 -2613
rect 5168 -2647 5178 -2613
rect 5126 -2685 5178 -2647
rect 5388 -2613 5440 -2575
rect 5388 -2647 5398 -2613
rect 5432 -2647 5440 -2613
rect 5388 -2685 5440 -2647
rect 5692 -2601 5742 -2555
rect 5586 -2628 5640 -2601
rect 5586 -2662 5595 -2628
rect 5629 -2662 5640 -2628
rect 5586 -2685 5640 -2662
rect 5670 -2628 5742 -2601
rect 5670 -2662 5692 -2628
rect 5726 -2662 5742 -2628
rect 5670 -2685 5742 -2662
rect 5842 -2628 5894 -2555
rect 5842 -2662 5852 -2628
rect 5886 -2662 5894 -2628
rect 5842 -2685 5894 -2662
rect 5949 -2628 6002 -2555
rect 5949 -2662 5957 -2628
rect 5991 -2662 6002 -2628
rect 5949 -2685 6002 -2662
rect 6102 -2601 6152 -2555
rect 6102 -2628 6167 -2601
rect 6102 -2662 6113 -2628
rect 6147 -2662 6167 -2628
rect 6102 -2685 6167 -2662
rect 6197 -2628 6268 -2601
rect 6197 -2662 6211 -2628
rect 6245 -2662 6268 -2628
rect 6197 -2685 6268 -2662
rect 6414 -2613 6466 -2575
rect 6414 -2647 6422 -2613
rect 6456 -2647 6466 -2613
rect 6414 -2685 6466 -2647
rect 6676 -2613 6728 -2575
rect 6676 -2647 6686 -2613
rect 6720 -2647 6728 -2613
rect 6676 -2685 6728 -2647
rect 6874 -2620 6926 -2575
rect 6874 -2654 6882 -2620
rect 6916 -2654 6926 -2620
rect 6874 -2685 6926 -2654
rect 7504 -2620 7556 -2575
rect 7504 -2654 7514 -2620
rect 7548 -2654 7556 -2620
rect 7504 -2685 7556 -2654
rect 7702 -2613 7754 -2575
rect 7702 -2647 7710 -2613
rect 7744 -2647 7754 -2613
rect 7702 -2685 7754 -2647
rect 7964 -2613 8016 -2575
rect 7964 -2647 7974 -2613
rect 8008 -2647 8016 -2613
rect 7964 -2685 8016 -2647
rect 8268 -2601 8318 -2555
rect 8162 -2628 8216 -2601
rect 8162 -2662 8171 -2628
rect 8205 -2662 8216 -2628
rect 8162 -2685 8216 -2662
rect 8246 -2628 8318 -2601
rect 8246 -2662 8268 -2628
rect 8302 -2662 8318 -2628
rect 8246 -2685 8318 -2662
rect 8418 -2628 8470 -2555
rect 8418 -2662 8428 -2628
rect 8462 -2662 8470 -2628
rect 8418 -2685 8470 -2662
rect 8525 -2628 8578 -2555
rect 8525 -2662 8533 -2628
rect 8567 -2662 8578 -2628
rect 8525 -2685 8578 -2662
rect 8678 -2601 8728 -2555
rect 8678 -2628 8743 -2601
rect 8678 -2662 8689 -2628
rect 8723 -2662 8743 -2628
rect 8678 -2685 8743 -2662
rect 8773 -2628 8844 -2601
rect 8773 -2662 8787 -2628
rect 8821 -2662 8844 -2628
rect 8773 -2685 8844 -2662
rect 8990 -2613 9042 -2575
rect 8990 -2647 8998 -2613
rect 9032 -2647 9042 -2613
rect 8990 -2685 9042 -2647
rect 9252 -2613 9304 -2575
rect 9252 -2647 9262 -2613
rect 9296 -2647 9304 -2613
rect 9252 -2685 9304 -2647
rect 9450 -2620 9502 -2575
rect 9450 -2654 9458 -2620
rect 9492 -2654 9502 -2620
rect 9450 -2685 9502 -2654
rect 10080 -2620 10132 -2575
rect 10080 -2654 10090 -2620
rect 10124 -2654 10132 -2620
rect 10080 -2685 10132 -2654
rect 10370 -2613 10422 -2575
rect 10370 -2647 10378 -2613
rect 10412 -2647 10422 -2613
rect 10370 -2685 10422 -2647
rect 10632 -2613 10684 -2575
rect 10844 -2601 10894 -2555
rect 10632 -2647 10642 -2613
rect 10676 -2647 10684 -2613
rect 10632 -2685 10684 -2647
rect 10738 -2628 10792 -2601
rect 10738 -2662 10747 -2628
rect 10781 -2662 10792 -2628
rect 10738 -2685 10792 -2662
rect 10822 -2628 10894 -2601
rect 10822 -2662 10844 -2628
rect 10878 -2662 10894 -2628
rect 10822 -2685 10894 -2662
rect 10994 -2628 11046 -2555
rect 10994 -2662 11004 -2628
rect 11038 -2662 11046 -2628
rect 10994 -2685 11046 -2662
rect 11101 -2628 11154 -2555
rect 11101 -2662 11109 -2628
rect 11143 -2662 11154 -2628
rect 11101 -2685 11154 -2662
rect 11254 -2601 11304 -2555
rect 11254 -2628 11319 -2601
rect 11254 -2662 11265 -2628
rect 11299 -2662 11319 -2628
rect 11254 -2685 11319 -2662
rect 11349 -2628 11420 -2601
rect 11349 -2662 11363 -2628
rect 11397 -2662 11420 -2628
rect 11349 -2685 11420 -2662
rect 11658 -2613 11710 -2575
rect 11658 -2647 11666 -2613
rect 11700 -2647 11710 -2613
rect 11658 -2685 11710 -2647
rect 11920 -2613 11972 -2575
rect 11920 -2647 11930 -2613
rect 11964 -2647 11972 -2613
rect 11920 -2685 11972 -2647
rect 12567 -2637 12633 -2601
rect 12567 -2671 12588 -2637
rect 12622 -2671 12633 -2637
rect 12567 -2685 12633 -2671
rect 12663 -2626 12719 -2601
rect 12663 -2660 12674 -2626
rect 12708 -2660 12719 -2626
rect 12663 -2685 12719 -2660
rect 12749 -2637 12805 -2601
rect 12749 -2671 12760 -2637
rect 12794 -2671 12805 -2637
rect 12749 -2685 12805 -2671
rect 12835 -2626 12891 -2601
rect 12835 -2660 12846 -2626
rect 12880 -2660 12891 -2626
rect 12835 -2685 12891 -2660
rect 12921 -2637 13000 -2601
rect 12921 -2671 12932 -2637
rect 12966 -2671 13000 -2637
rect 13222 -2613 13274 -2575
rect 13222 -2647 13230 -2613
rect 13264 -2647 13274 -2613
rect 12921 -2685 13000 -2671
rect 13222 -2685 13274 -2647
rect 13484 -2613 13536 -2575
rect 13484 -2647 13494 -2613
rect 13528 -2647 13536 -2613
rect 13484 -2685 13536 -2647
rect 13682 -2639 13735 -2601
rect 13682 -2673 13690 -2639
rect 13724 -2673 13735 -2639
rect 13682 -2685 13735 -2673
rect 13765 -2626 13821 -2601
rect 13765 -2660 13776 -2626
rect 13810 -2660 13821 -2626
rect 13765 -2685 13821 -2660
rect 13851 -2626 13907 -2601
rect 13851 -2660 13862 -2626
rect 13896 -2660 13907 -2626
rect 13851 -2685 13907 -2660
rect 13937 -2626 13993 -2601
rect 13937 -2660 13948 -2626
rect 13982 -2660 13993 -2626
rect 13937 -2685 13993 -2660
rect 14023 -2626 14079 -2601
rect 14023 -2660 14034 -2626
rect 14068 -2660 14079 -2626
rect 14023 -2685 14079 -2660
rect 14109 -2626 14165 -2601
rect 14109 -2660 14120 -2626
rect 14154 -2660 14165 -2626
rect 14109 -2685 14165 -2660
rect 14195 -2635 14251 -2601
rect 14195 -2669 14206 -2635
rect 14240 -2669 14251 -2635
rect 14195 -2685 14251 -2669
rect 14281 -2626 14337 -2601
rect 14281 -2660 14292 -2626
rect 14326 -2660 14337 -2626
rect 14281 -2685 14337 -2660
rect 14367 -2635 14423 -2601
rect 14367 -2669 14378 -2635
rect 14412 -2669 14423 -2635
rect 14367 -2685 14423 -2669
rect 14453 -2626 14509 -2601
rect 14453 -2660 14464 -2626
rect 14498 -2660 14509 -2626
rect 14453 -2685 14509 -2660
rect 14539 -2635 14595 -2601
rect 14539 -2669 14550 -2635
rect 14584 -2669 14595 -2635
rect 14539 -2685 14595 -2669
rect 14625 -2626 14681 -2601
rect 14625 -2660 14636 -2626
rect 14670 -2660 14681 -2626
rect 14625 -2685 14681 -2660
rect 14711 -2635 14766 -2601
rect 14711 -2669 14722 -2635
rect 14756 -2669 14766 -2635
rect 14711 -2685 14766 -2669
rect 14796 -2626 14852 -2601
rect 14796 -2660 14807 -2626
rect 14841 -2660 14852 -2626
rect 14796 -2685 14852 -2660
rect 14882 -2635 14938 -2601
rect 14882 -2669 14893 -2635
rect 14927 -2669 14938 -2635
rect 14882 -2685 14938 -2669
rect 14968 -2626 15024 -2601
rect 14968 -2660 14979 -2626
rect 15013 -2660 15024 -2626
rect 14968 -2685 15024 -2660
rect 15054 -2635 15110 -2601
rect 15054 -2669 15065 -2635
rect 15099 -2669 15110 -2635
rect 15054 -2685 15110 -2669
rect 15140 -2626 15196 -2601
rect 15140 -2660 15151 -2626
rect 15185 -2660 15196 -2626
rect 15140 -2685 15196 -2660
rect 15226 -2635 15282 -2601
rect 15226 -2669 15237 -2635
rect 15271 -2669 15282 -2635
rect 15226 -2685 15282 -2669
rect 15312 -2626 15368 -2601
rect 15312 -2660 15323 -2626
rect 15357 -2660 15368 -2626
rect 15312 -2685 15368 -2660
rect 15398 -2635 15451 -2601
rect 15398 -2669 15409 -2635
rect 15443 -2669 15451 -2635
rect 15614 -2620 15666 -2575
rect 15614 -2654 15622 -2620
rect 15656 -2654 15666 -2620
rect 15398 -2685 15451 -2669
rect 15614 -2685 15666 -2654
rect 16612 -2620 16664 -2575
rect 16612 -2654 16622 -2620
rect 16656 -2654 16664 -2620
rect 16612 -2685 16664 -2654
rect -2970 -2810 -2918 -2779
rect -2970 -2844 -2962 -2810
rect -2928 -2844 -2918 -2810
rect -2970 -2889 -2918 -2844
rect -2340 -2810 -2288 -2779
rect -2340 -2844 -2330 -2810
rect -2296 -2844 -2288 -2810
rect -2340 -2889 -2288 -2844
rect -1875 -2802 -1823 -2779
rect -1875 -2836 -1867 -2802
rect -1833 -2836 -1823 -2802
rect -1875 -2863 -1823 -2836
rect -1793 -2800 -1736 -2779
rect -1793 -2834 -1783 -2800
rect -1749 -2834 -1736 -2800
rect -1793 -2863 -1736 -2834
rect -1590 -2810 -1538 -2779
rect -1590 -2844 -1582 -2810
rect -1548 -2844 -1538 -2810
rect -1590 -2889 -1538 -2844
rect -960 -2810 -908 -2779
rect -960 -2844 -950 -2810
rect -916 -2844 -908 -2810
rect -960 -2889 -908 -2844
rect -854 -2810 -802 -2779
rect -854 -2844 -846 -2810
rect -812 -2844 -802 -2810
rect -854 -2889 -802 -2844
rect -224 -2810 -172 -2779
rect -224 -2844 -214 -2810
rect -180 -2844 -172 -2810
rect -224 -2889 -172 -2844
rect -26 -2817 26 -2779
rect -26 -2851 -18 -2817
rect 16 -2851 26 -2817
rect -26 -2889 26 -2851
rect 236 -2817 288 -2779
rect 236 -2851 246 -2817
rect 280 -2851 288 -2817
rect 236 -2889 288 -2851
rect 434 -2802 505 -2779
rect 434 -2836 457 -2802
rect 491 -2836 505 -2802
rect 434 -2863 505 -2836
rect 535 -2802 600 -2779
rect 535 -2836 555 -2802
rect 589 -2836 600 -2802
rect 535 -2863 600 -2836
rect 550 -2909 600 -2863
rect 700 -2802 753 -2779
rect 700 -2836 711 -2802
rect 745 -2836 753 -2802
rect 700 -2909 753 -2836
rect 808 -2802 860 -2779
rect 808 -2836 816 -2802
rect 850 -2836 860 -2802
rect 808 -2909 860 -2836
rect 960 -2802 1032 -2779
rect 960 -2836 976 -2802
rect 1010 -2836 1032 -2802
rect 960 -2863 1032 -2836
rect 1062 -2802 1116 -2779
rect 1062 -2836 1073 -2802
rect 1107 -2836 1116 -2802
rect 1062 -2863 1116 -2836
rect 960 -2909 1010 -2863
rect 1262 -2817 1314 -2779
rect 1262 -2851 1270 -2817
rect 1304 -2851 1314 -2817
rect 1262 -2889 1314 -2851
rect 1524 -2817 1576 -2779
rect 1524 -2851 1534 -2817
rect 1568 -2851 1576 -2817
rect 1524 -2889 1576 -2851
rect 1722 -2810 1774 -2779
rect 1722 -2844 1730 -2810
rect 1764 -2844 1774 -2810
rect 1722 -2889 1774 -2844
rect 2352 -2810 2404 -2779
rect 2352 -2844 2362 -2810
rect 2396 -2844 2404 -2810
rect 2352 -2889 2404 -2844
rect 2550 -2817 2602 -2779
rect 2550 -2851 2558 -2817
rect 2592 -2851 2602 -2817
rect 2550 -2889 2602 -2851
rect 2812 -2817 2864 -2779
rect 2812 -2851 2822 -2817
rect 2856 -2851 2864 -2817
rect 2812 -2889 2864 -2851
rect 3010 -2802 3081 -2779
rect 3010 -2836 3033 -2802
rect 3067 -2836 3081 -2802
rect 3010 -2863 3081 -2836
rect 3111 -2802 3176 -2779
rect 3111 -2836 3131 -2802
rect 3165 -2836 3176 -2802
rect 3111 -2863 3176 -2836
rect 3126 -2909 3176 -2863
rect 3276 -2802 3329 -2779
rect 3276 -2836 3287 -2802
rect 3321 -2836 3329 -2802
rect 3276 -2909 3329 -2836
rect 3384 -2802 3436 -2779
rect 3384 -2836 3392 -2802
rect 3426 -2836 3436 -2802
rect 3384 -2909 3436 -2836
rect 3536 -2802 3608 -2779
rect 3536 -2836 3552 -2802
rect 3586 -2836 3608 -2802
rect 3536 -2863 3608 -2836
rect 3638 -2802 3692 -2779
rect 3638 -2836 3649 -2802
rect 3683 -2836 3692 -2802
rect 3638 -2863 3692 -2836
rect 3536 -2909 3586 -2863
rect 3838 -2817 3890 -2779
rect 3838 -2851 3846 -2817
rect 3880 -2851 3890 -2817
rect 3838 -2889 3890 -2851
rect 4100 -2817 4152 -2779
rect 4100 -2851 4110 -2817
rect 4144 -2851 4152 -2817
rect 4100 -2889 4152 -2851
rect 4298 -2810 4350 -2779
rect 4298 -2844 4306 -2810
rect 4340 -2844 4350 -2810
rect 4298 -2889 4350 -2844
rect 4928 -2810 4980 -2779
rect 4928 -2844 4938 -2810
rect 4972 -2844 4980 -2810
rect 4928 -2889 4980 -2844
rect 5126 -2817 5178 -2779
rect 5126 -2851 5134 -2817
rect 5168 -2851 5178 -2817
rect 5126 -2889 5178 -2851
rect 5388 -2817 5440 -2779
rect 5388 -2851 5398 -2817
rect 5432 -2851 5440 -2817
rect 5388 -2889 5440 -2851
rect 5586 -2802 5657 -2779
rect 5586 -2836 5609 -2802
rect 5643 -2836 5657 -2802
rect 5586 -2863 5657 -2836
rect 5687 -2802 5752 -2779
rect 5687 -2836 5707 -2802
rect 5741 -2836 5752 -2802
rect 5687 -2863 5752 -2836
rect 5702 -2909 5752 -2863
rect 5852 -2802 5905 -2779
rect 5852 -2836 5863 -2802
rect 5897 -2836 5905 -2802
rect 5852 -2909 5905 -2836
rect 5960 -2802 6012 -2779
rect 5960 -2836 5968 -2802
rect 6002 -2836 6012 -2802
rect 5960 -2909 6012 -2836
rect 6112 -2802 6184 -2779
rect 6112 -2836 6128 -2802
rect 6162 -2836 6184 -2802
rect 6112 -2863 6184 -2836
rect 6214 -2802 6268 -2779
rect 6214 -2836 6225 -2802
rect 6259 -2836 6268 -2802
rect 6214 -2863 6268 -2836
rect 6112 -2909 6162 -2863
rect 6414 -2817 6466 -2779
rect 6414 -2851 6422 -2817
rect 6456 -2851 6466 -2817
rect 6414 -2889 6466 -2851
rect 6676 -2817 6728 -2779
rect 6676 -2851 6686 -2817
rect 6720 -2851 6728 -2817
rect 6676 -2889 6728 -2851
rect 6874 -2810 6926 -2779
rect 6874 -2844 6882 -2810
rect 6916 -2844 6926 -2810
rect 6874 -2889 6926 -2844
rect 7504 -2810 7556 -2779
rect 7504 -2844 7514 -2810
rect 7548 -2844 7556 -2810
rect 7504 -2889 7556 -2844
rect 7702 -2817 7754 -2779
rect 7702 -2851 7710 -2817
rect 7744 -2851 7754 -2817
rect 7702 -2889 7754 -2851
rect 7964 -2817 8016 -2779
rect 7964 -2851 7974 -2817
rect 8008 -2851 8016 -2817
rect 7964 -2889 8016 -2851
rect 8162 -2802 8233 -2779
rect 8162 -2836 8185 -2802
rect 8219 -2836 8233 -2802
rect 8162 -2863 8233 -2836
rect 8263 -2802 8328 -2779
rect 8263 -2836 8283 -2802
rect 8317 -2836 8328 -2802
rect 8263 -2863 8328 -2836
rect 8278 -2909 8328 -2863
rect 8428 -2802 8481 -2779
rect 8428 -2836 8439 -2802
rect 8473 -2836 8481 -2802
rect 8428 -2909 8481 -2836
rect 8536 -2802 8588 -2779
rect 8536 -2836 8544 -2802
rect 8578 -2836 8588 -2802
rect 8536 -2909 8588 -2836
rect 8688 -2802 8760 -2779
rect 8688 -2836 8704 -2802
rect 8738 -2836 8760 -2802
rect 8688 -2863 8760 -2836
rect 8790 -2802 8844 -2779
rect 8790 -2836 8801 -2802
rect 8835 -2836 8844 -2802
rect 8790 -2863 8844 -2836
rect 8688 -2909 8738 -2863
rect 8990 -2817 9042 -2779
rect 8990 -2851 8998 -2817
rect 9032 -2851 9042 -2817
rect 8990 -2889 9042 -2851
rect 9252 -2817 9304 -2779
rect 9252 -2851 9262 -2817
rect 9296 -2851 9304 -2817
rect 9252 -2889 9304 -2851
rect 9450 -2810 9502 -2779
rect 9450 -2844 9458 -2810
rect 9492 -2844 9502 -2810
rect 9450 -2889 9502 -2844
rect 10080 -2810 10132 -2779
rect 10080 -2844 10090 -2810
rect 10124 -2844 10132 -2810
rect 10080 -2889 10132 -2844
rect 10370 -2817 10422 -2779
rect 10370 -2851 10378 -2817
rect 10412 -2851 10422 -2817
rect 10370 -2889 10422 -2851
rect 10632 -2817 10684 -2779
rect 10632 -2851 10642 -2817
rect 10676 -2851 10684 -2817
rect 10632 -2889 10684 -2851
rect 10738 -2802 10809 -2779
rect 10738 -2836 10761 -2802
rect 10795 -2836 10809 -2802
rect 10738 -2863 10809 -2836
rect 10839 -2802 10904 -2779
rect 10839 -2836 10859 -2802
rect 10893 -2836 10904 -2802
rect 10839 -2863 10904 -2836
rect 10854 -2909 10904 -2863
rect 11004 -2802 11057 -2779
rect 11004 -2836 11015 -2802
rect 11049 -2836 11057 -2802
rect 11004 -2909 11057 -2836
rect 11112 -2802 11164 -2779
rect 11112 -2836 11120 -2802
rect 11154 -2836 11164 -2802
rect 11112 -2909 11164 -2836
rect 11264 -2802 11336 -2779
rect 11264 -2836 11280 -2802
rect 11314 -2836 11336 -2802
rect 11264 -2863 11336 -2836
rect 11366 -2802 11420 -2779
rect 11366 -2836 11377 -2802
rect 11411 -2836 11420 -2802
rect 11366 -2863 11420 -2836
rect 11264 -2909 11314 -2863
rect 11658 -2817 11710 -2779
rect 11658 -2851 11666 -2817
rect 11700 -2851 11710 -2817
rect 11658 -2889 11710 -2851
rect 11920 -2817 11972 -2779
rect 11920 -2851 11930 -2817
rect 11964 -2851 11972 -2817
rect 11920 -2889 11972 -2851
rect 13590 -2810 13642 -2779
rect 13590 -2844 13598 -2810
rect 13632 -2844 13642 -2810
rect 13590 -2889 13642 -2844
rect 14588 -2810 14640 -2779
rect 14588 -2844 14598 -2810
rect 14632 -2844 14640 -2810
rect 14588 -2889 14640 -2844
rect 14786 -2810 14838 -2779
rect 14786 -2844 14794 -2810
rect 14828 -2844 14838 -2810
rect 14786 -2889 14838 -2844
rect 15784 -2810 15836 -2779
rect 15784 -2844 15794 -2810
rect 15828 -2844 15836 -2810
rect 15784 -2889 15836 -2844
rect 15982 -2810 16034 -2779
rect 15982 -2844 15990 -2810
rect 16024 -2844 16034 -2810
rect 15982 -2889 16034 -2844
rect 16612 -2810 16664 -2779
rect 16612 -2844 16622 -2810
rect 16656 -2844 16664 -2810
rect 16612 -2889 16664 -2844
rect -2970 -3708 -2918 -3663
rect -2970 -3742 -2962 -3708
rect -2928 -3742 -2918 -3708
rect -2970 -3773 -2918 -3742
rect -2340 -3708 -2288 -3663
rect -2340 -3742 -2330 -3708
rect -2296 -3742 -2288 -3708
rect -2340 -3773 -2288 -3742
rect -1590 -3708 -1538 -3663
rect -1590 -3742 -1582 -3708
rect -1548 -3742 -1538 -3708
rect -1590 -3773 -1538 -3742
rect -960 -3708 -908 -3663
rect -960 -3742 -950 -3708
rect -916 -3742 -908 -3708
rect -960 -3773 -908 -3742
rect -854 -3708 -802 -3663
rect -854 -3742 -846 -3708
rect -812 -3742 -802 -3708
rect -854 -3773 -802 -3742
rect -224 -3708 -172 -3663
rect -224 -3742 -214 -3708
rect -180 -3742 -172 -3708
rect -224 -3773 -172 -3742
rect -26 -3701 26 -3663
rect -26 -3735 -18 -3701
rect 16 -3735 26 -3701
rect -26 -3773 26 -3735
rect 236 -3701 288 -3663
rect 236 -3735 246 -3701
rect 280 -3735 288 -3701
rect 236 -3773 288 -3735
rect 550 -3689 600 -3643
rect 434 -3716 505 -3689
rect 434 -3750 457 -3716
rect 491 -3750 505 -3716
rect 434 -3773 505 -3750
rect 535 -3716 600 -3689
rect 535 -3750 555 -3716
rect 589 -3750 600 -3716
rect 535 -3773 600 -3750
rect 700 -3716 753 -3643
rect 700 -3750 711 -3716
rect 745 -3750 753 -3716
rect 700 -3773 753 -3750
rect 808 -3716 860 -3643
rect 808 -3750 816 -3716
rect 850 -3750 860 -3716
rect 808 -3773 860 -3750
rect 960 -3689 1010 -3643
rect 960 -3716 1032 -3689
rect 960 -3750 976 -3716
rect 1010 -3750 1032 -3716
rect 960 -3773 1032 -3750
rect 1062 -3716 1116 -3689
rect 1062 -3750 1073 -3716
rect 1107 -3750 1116 -3716
rect 1062 -3773 1116 -3750
rect 1262 -3701 1314 -3663
rect 1262 -3735 1270 -3701
rect 1304 -3735 1314 -3701
rect 1262 -3773 1314 -3735
rect 1524 -3701 1576 -3663
rect 1524 -3735 1534 -3701
rect 1568 -3735 1576 -3701
rect 1524 -3773 1576 -3735
rect 1722 -3708 1774 -3663
rect 1722 -3742 1730 -3708
rect 1764 -3742 1774 -3708
rect 1722 -3773 1774 -3742
rect 2352 -3708 2404 -3663
rect 2352 -3742 2362 -3708
rect 2396 -3742 2404 -3708
rect 2352 -3773 2404 -3742
rect 2550 -3701 2602 -3663
rect 2550 -3735 2558 -3701
rect 2592 -3735 2602 -3701
rect 2550 -3773 2602 -3735
rect 2812 -3701 2864 -3663
rect 2812 -3735 2822 -3701
rect 2856 -3735 2864 -3701
rect 2812 -3773 2864 -3735
rect 3126 -3689 3176 -3643
rect 3010 -3716 3081 -3689
rect 3010 -3750 3033 -3716
rect 3067 -3750 3081 -3716
rect 3010 -3773 3081 -3750
rect 3111 -3716 3176 -3689
rect 3111 -3750 3131 -3716
rect 3165 -3750 3176 -3716
rect 3111 -3773 3176 -3750
rect 3276 -3716 3329 -3643
rect 3276 -3750 3287 -3716
rect 3321 -3750 3329 -3716
rect 3276 -3773 3329 -3750
rect 3384 -3716 3436 -3643
rect 3384 -3750 3392 -3716
rect 3426 -3750 3436 -3716
rect 3384 -3773 3436 -3750
rect 3536 -3689 3586 -3643
rect 3536 -3716 3608 -3689
rect 3536 -3750 3552 -3716
rect 3586 -3750 3608 -3716
rect 3536 -3773 3608 -3750
rect 3638 -3716 3692 -3689
rect 3638 -3750 3649 -3716
rect 3683 -3750 3692 -3716
rect 3638 -3773 3692 -3750
rect 3838 -3701 3890 -3663
rect 3838 -3735 3846 -3701
rect 3880 -3735 3890 -3701
rect 3838 -3773 3890 -3735
rect 4100 -3701 4152 -3663
rect 4100 -3735 4110 -3701
rect 4144 -3735 4152 -3701
rect 4100 -3773 4152 -3735
rect 4298 -3708 4350 -3663
rect 4298 -3742 4306 -3708
rect 4340 -3742 4350 -3708
rect 4298 -3773 4350 -3742
rect 4928 -3708 4980 -3663
rect 4928 -3742 4938 -3708
rect 4972 -3742 4980 -3708
rect 4928 -3773 4980 -3742
rect 5126 -3701 5178 -3663
rect 5126 -3735 5134 -3701
rect 5168 -3735 5178 -3701
rect 5126 -3773 5178 -3735
rect 5388 -3701 5440 -3663
rect 5388 -3735 5398 -3701
rect 5432 -3735 5440 -3701
rect 5388 -3773 5440 -3735
rect 5702 -3689 5752 -3643
rect 5586 -3716 5657 -3689
rect 5586 -3750 5609 -3716
rect 5643 -3750 5657 -3716
rect 5586 -3773 5657 -3750
rect 5687 -3716 5752 -3689
rect 5687 -3750 5707 -3716
rect 5741 -3750 5752 -3716
rect 5687 -3773 5752 -3750
rect 5852 -3716 5905 -3643
rect 5852 -3750 5863 -3716
rect 5897 -3750 5905 -3716
rect 5852 -3773 5905 -3750
rect 5960 -3716 6012 -3643
rect 5960 -3750 5968 -3716
rect 6002 -3750 6012 -3716
rect 5960 -3773 6012 -3750
rect 6112 -3689 6162 -3643
rect 6112 -3716 6184 -3689
rect 6112 -3750 6128 -3716
rect 6162 -3750 6184 -3716
rect 6112 -3773 6184 -3750
rect 6214 -3716 6268 -3689
rect 6214 -3750 6225 -3716
rect 6259 -3750 6268 -3716
rect 6214 -3773 6268 -3750
rect 6414 -3701 6466 -3663
rect 6414 -3735 6422 -3701
rect 6456 -3735 6466 -3701
rect 6414 -3773 6466 -3735
rect 6676 -3701 6728 -3663
rect 6676 -3735 6686 -3701
rect 6720 -3735 6728 -3701
rect 6676 -3773 6728 -3735
rect 6874 -3708 6926 -3663
rect 6874 -3742 6882 -3708
rect 6916 -3742 6926 -3708
rect 6874 -3773 6926 -3742
rect 7504 -3708 7556 -3663
rect 7504 -3742 7514 -3708
rect 7548 -3742 7556 -3708
rect 7504 -3773 7556 -3742
rect 7702 -3701 7754 -3663
rect 7702 -3735 7710 -3701
rect 7744 -3735 7754 -3701
rect 7702 -3773 7754 -3735
rect 7964 -3701 8016 -3663
rect 7964 -3735 7974 -3701
rect 8008 -3735 8016 -3701
rect 7964 -3773 8016 -3735
rect 8278 -3689 8328 -3643
rect 8162 -3716 8233 -3689
rect 8162 -3750 8185 -3716
rect 8219 -3750 8233 -3716
rect 8162 -3773 8233 -3750
rect 8263 -3716 8328 -3689
rect 8263 -3750 8283 -3716
rect 8317 -3750 8328 -3716
rect 8263 -3773 8328 -3750
rect 8428 -3716 8481 -3643
rect 8428 -3750 8439 -3716
rect 8473 -3750 8481 -3716
rect 8428 -3773 8481 -3750
rect 8536 -3716 8588 -3643
rect 8536 -3750 8544 -3716
rect 8578 -3750 8588 -3716
rect 8536 -3773 8588 -3750
rect 8688 -3689 8738 -3643
rect 8688 -3716 8760 -3689
rect 8688 -3750 8704 -3716
rect 8738 -3750 8760 -3716
rect 8688 -3773 8760 -3750
rect 8790 -3716 8844 -3689
rect 8790 -3750 8801 -3716
rect 8835 -3750 8844 -3716
rect 8790 -3773 8844 -3750
rect 8990 -3701 9042 -3663
rect 8990 -3735 8998 -3701
rect 9032 -3735 9042 -3701
rect 8990 -3773 9042 -3735
rect 9252 -3701 9304 -3663
rect 9252 -3735 9262 -3701
rect 9296 -3735 9304 -3701
rect 9252 -3773 9304 -3735
rect 9450 -3708 9502 -3663
rect 9450 -3742 9458 -3708
rect 9492 -3742 9502 -3708
rect 9450 -3773 9502 -3742
rect 10080 -3708 10132 -3663
rect 10080 -3742 10090 -3708
rect 10124 -3742 10132 -3708
rect 10080 -3773 10132 -3742
rect 10370 -3701 10422 -3663
rect 10370 -3735 10378 -3701
rect 10412 -3735 10422 -3701
rect 10370 -3773 10422 -3735
rect 10632 -3701 10684 -3663
rect 10854 -3689 10904 -3643
rect 10632 -3735 10642 -3701
rect 10676 -3735 10684 -3701
rect 10632 -3773 10684 -3735
rect 10738 -3716 10809 -3689
rect 10738 -3750 10761 -3716
rect 10795 -3750 10809 -3716
rect 10738 -3773 10809 -3750
rect 10839 -3716 10904 -3689
rect 10839 -3750 10859 -3716
rect 10893 -3750 10904 -3716
rect 10839 -3773 10904 -3750
rect 11004 -3716 11057 -3643
rect 11004 -3750 11015 -3716
rect 11049 -3750 11057 -3716
rect 11004 -3773 11057 -3750
rect 11112 -3716 11164 -3643
rect 11112 -3750 11120 -3716
rect 11154 -3750 11164 -3716
rect 11112 -3773 11164 -3750
rect 11264 -3689 11314 -3643
rect 11264 -3716 11336 -3689
rect 11264 -3750 11280 -3716
rect 11314 -3750 11336 -3716
rect 11264 -3773 11336 -3750
rect 11366 -3716 11420 -3689
rect 11366 -3750 11377 -3716
rect 11411 -3750 11420 -3716
rect 11366 -3773 11420 -3750
rect 11658 -3701 11710 -3663
rect 11658 -3735 11666 -3701
rect 11700 -3735 11710 -3701
rect 11658 -3773 11710 -3735
rect 11920 -3701 11972 -3663
rect 11920 -3735 11930 -3701
rect 11964 -3735 11972 -3701
rect 11920 -3773 11972 -3735
rect 13590 -3708 13642 -3663
rect 13590 -3742 13598 -3708
rect 13632 -3742 13642 -3708
rect 13590 -3773 13642 -3742
rect 14588 -3708 14640 -3663
rect 14588 -3742 14598 -3708
rect 14632 -3742 14640 -3708
rect 14588 -3773 14640 -3742
rect 14786 -3708 14838 -3663
rect 14786 -3742 14794 -3708
rect 14828 -3742 14838 -3708
rect 14786 -3773 14838 -3742
rect 15784 -3708 15836 -3663
rect 15784 -3742 15794 -3708
rect 15828 -3742 15836 -3708
rect 15784 -3773 15836 -3742
rect 15982 -3708 16034 -3663
rect 15982 -3742 15990 -3708
rect 16024 -3742 16034 -3708
rect 15982 -3773 16034 -3742
rect 16612 -3708 16664 -3663
rect 16612 -3742 16622 -3708
rect 16656 -3742 16664 -3708
rect 16612 -3773 16664 -3742
rect -2970 -3898 -2918 -3867
rect -2970 -3932 -2962 -3898
rect -2928 -3932 -2918 -3898
rect -2970 -3977 -2918 -3932
rect -2340 -3898 -2288 -3867
rect -2340 -3932 -2330 -3898
rect -2296 -3932 -2288 -3898
rect -2340 -3977 -2288 -3932
rect -1590 -3898 -1538 -3867
rect -1590 -3932 -1582 -3898
rect -1548 -3932 -1538 -3898
rect -1590 -3977 -1538 -3932
rect -960 -3898 -908 -3867
rect -960 -3932 -950 -3898
rect -916 -3932 -908 -3898
rect -960 -3977 -908 -3932
rect -854 -3898 -802 -3867
rect -854 -3932 -846 -3898
rect -812 -3932 -802 -3898
rect -854 -3977 -802 -3932
rect -224 -3898 -172 -3867
rect -224 -3932 -214 -3898
rect -180 -3932 -172 -3898
rect -224 -3977 -172 -3932
rect -26 -3905 26 -3867
rect -26 -3939 -18 -3905
rect 16 -3939 26 -3905
rect -26 -3977 26 -3939
rect 236 -3905 288 -3867
rect 236 -3939 246 -3905
rect 280 -3939 288 -3905
rect 236 -3977 288 -3939
rect 434 -3890 488 -3867
rect 434 -3924 443 -3890
rect 477 -3924 488 -3890
rect 434 -3951 488 -3924
rect 518 -3890 590 -3867
rect 518 -3924 540 -3890
rect 574 -3924 590 -3890
rect 518 -3951 590 -3924
rect 540 -3997 590 -3951
rect 690 -3890 742 -3867
rect 690 -3924 700 -3890
rect 734 -3924 742 -3890
rect 690 -3997 742 -3924
rect 797 -3890 850 -3867
rect 797 -3924 805 -3890
rect 839 -3924 850 -3890
rect 797 -3997 850 -3924
rect 950 -3890 1015 -3867
rect 950 -3924 961 -3890
rect 995 -3924 1015 -3890
rect 950 -3951 1015 -3924
rect 1045 -3890 1116 -3867
rect 1045 -3924 1059 -3890
rect 1093 -3924 1116 -3890
rect 1045 -3951 1116 -3924
rect 950 -3997 1000 -3951
rect 1262 -3905 1314 -3867
rect 1262 -3939 1270 -3905
rect 1304 -3939 1314 -3905
rect 1262 -3977 1314 -3939
rect 1524 -3905 1576 -3867
rect 1524 -3939 1534 -3905
rect 1568 -3939 1576 -3905
rect 1524 -3977 1576 -3939
rect 1722 -3898 1774 -3867
rect 1722 -3932 1730 -3898
rect 1764 -3932 1774 -3898
rect 1722 -3977 1774 -3932
rect 2352 -3898 2404 -3867
rect 2352 -3932 2362 -3898
rect 2396 -3932 2404 -3898
rect 2352 -3977 2404 -3932
rect 2550 -3905 2602 -3867
rect 2550 -3939 2558 -3905
rect 2592 -3939 2602 -3905
rect 2550 -3977 2602 -3939
rect 2812 -3905 2864 -3867
rect 2812 -3939 2822 -3905
rect 2856 -3939 2864 -3905
rect 2812 -3977 2864 -3939
rect 3010 -3890 3064 -3867
rect 3010 -3924 3019 -3890
rect 3053 -3924 3064 -3890
rect 3010 -3951 3064 -3924
rect 3094 -3890 3166 -3867
rect 3094 -3924 3116 -3890
rect 3150 -3924 3166 -3890
rect 3094 -3951 3166 -3924
rect 3116 -3997 3166 -3951
rect 3266 -3890 3318 -3867
rect 3266 -3924 3276 -3890
rect 3310 -3924 3318 -3890
rect 3266 -3997 3318 -3924
rect 3373 -3890 3426 -3867
rect 3373 -3924 3381 -3890
rect 3415 -3924 3426 -3890
rect 3373 -3997 3426 -3924
rect 3526 -3890 3591 -3867
rect 3526 -3924 3537 -3890
rect 3571 -3924 3591 -3890
rect 3526 -3951 3591 -3924
rect 3621 -3890 3692 -3867
rect 3621 -3924 3635 -3890
rect 3669 -3924 3692 -3890
rect 3621 -3951 3692 -3924
rect 3526 -3997 3576 -3951
rect 3838 -3905 3890 -3867
rect 3838 -3939 3846 -3905
rect 3880 -3939 3890 -3905
rect 3838 -3977 3890 -3939
rect 4100 -3905 4152 -3867
rect 4100 -3939 4110 -3905
rect 4144 -3939 4152 -3905
rect 4100 -3977 4152 -3939
rect 4298 -3898 4350 -3867
rect 4298 -3932 4306 -3898
rect 4340 -3932 4350 -3898
rect 4298 -3977 4350 -3932
rect 4928 -3898 4980 -3867
rect 4928 -3932 4938 -3898
rect 4972 -3932 4980 -3898
rect 4928 -3977 4980 -3932
rect 5126 -3905 5178 -3867
rect 5126 -3939 5134 -3905
rect 5168 -3939 5178 -3905
rect 5126 -3977 5178 -3939
rect 5388 -3905 5440 -3867
rect 5388 -3939 5398 -3905
rect 5432 -3939 5440 -3905
rect 5388 -3977 5440 -3939
rect 5586 -3890 5640 -3867
rect 5586 -3924 5595 -3890
rect 5629 -3924 5640 -3890
rect 5586 -3951 5640 -3924
rect 5670 -3890 5742 -3867
rect 5670 -3924 5692 -3890
rect 5726 -3924 5742 -3890
rect 5670 -3951 5742 -3924
rect 5692 -3997 5742 -3951
rect 5842 -3890 5894 -3867
rect 5842 -3924 5852 -3890
rect 5886 -3924 5894 -3890
rect 5842 -3997 5894 -3924
rect 5949 -3890 6002 -3867
rect 5949 -3924 5957 -3890
rect 5991 -3924 6002 -3890
rect 5949 -3997 6002 -3924
rect 6102 -3890 6167 -3867
rect 6102 -3924 6113 -3890
rect 6147 -3924 6167 -3890
rect 6102 -3951 6167 -3924
rect 6197 -3890 6268 -3867
rect 6197 -3924 6211 -3890
rect 6245 -3924 6268 -3890
rect 6197 -3951 6268 -3924
rect 6102 -3997 6152 -3951
rect 6414 -3905 6466 -3867
rect 6414 -3939 6422 -3905
rect 6456 -3939 6466 -3905
rect 6414 -3977 6466 -3939
rect 6676 -3905 6728 -3867
rect 6676 -3939 6686 -3905
rect 6720 -3939 6728 -3905
rect 6676 -3977 6728 -3939
rect 6874 -3898 6926 -3867
rect 6874 -3932 6882 -3898
rect 6916 -3932 6926 -3898
rect 6874 -3977 6926 -3932
rect 7504 -3898 7556 -3867
rect 7504 -3932 7514 -3898
rect 7548 -3932 7556 -3898
rect 7504 -3977 7556 -3932
rect 7702 -3905 7754 -3867
rect 7702 -3939 7710 -3905
rect 7744 -3939 7754 -3905
rect 7702 -3977 7754 -3939
rect 7964 -3905 8016 -3867
rect 7964 -3939 7974 -3905
rect 8008 -3939 8016 -3905
rect 7964 -3977 8016 -3939
rect 8162 -3890 8216 -3867
rect 8162 -3924 8171 -3890
rect 8205 -3924 8216 -3890
rect 8162 -3951 8216 -3924
rect 8246 -3890 8318 -3867
rect 8246 -3924 8268 -3890
rect 8302 -3924 8318 -3890
rect 8246 -3951 8318 -3924
rect 8268 -3997 8318 -3951
rect 8418 -3890 8470 -3867
rect 8418 -3924 8428 -3890
rect 8462 -3924 8470 -3890
rect 8418 -3997 8470 -3924
rect 8525 -3890 8578 -3867
rect 8525 -3924 8533 -3890
rect 8567 -3924 8578 -3890
rect 8525 -3997 8578 -3924
rect 8678 -3890 8743 -3867
rect 8678 -3924 8689 -3890
rect 8723 -3924 8743 -3890
rect 8678 -3951 8743 -3924
rect 8773 -3890 8844 -3867
rect 8773 -3924 8787 -3890
rect 8821 -3924 8844 -3890
rect 8773 -3951 8844 -3924
rect 8678 -3997 8728 -3951
rect 8990 -3905 9042 -3867
rect 8990 -3939 8998 -3905
rect 9032 -3939 9042 -3905
rect 8990 -3977 9042 -3939
rect 9252 -3905 9304 -3867
rect 9252 -3939 9262 -3905
rect 9296 -3939 9304 -3905
rect 9252 -3977 9304 -3939
rect 9450 -3898 9502 -3867
rect 9450 -3932 9458 -3898
rect 9492 -3932 9502 -3898
rect 9450 -3977 9502 -3932
rect 10080 -3898 10132 -3867
rect 10080 -3932 10090 -3898
rect 10124 -3932 10132 -3898
rect 10080 -3977 10132 -3932
rect 10370 -3905 10422 -3867
rect 10370 -3939 10378 -3905
rect 10412 -3939 10422 -3905
rect 10370 -3977 10422 -3939
rect 10632 -3905 10684 -3867
rect 10632 -3939 10642 -3905
rect 10676 -3939 10684 -3905
rect 10632 -3977 10684 -3939
rect 10738 -3890 10792 -3867
rect 10738 -3924 10747 -3890
rect 10781 -3924 10792 -3890
rect 10738 -3951 10792 -3924
rect 10822 -3890 10894 -3867
rect 10822 -3924 10844 -3890
rect 10878 -3924 10894 -3890
rect 10822 -3951 10894 -3924
rect 10844 -3997 10894 -3951
rect 10994 -3890 11046 -3867
rect 10994 -3924 11004 -3890
rect 11038 -3924 11046 -3890
rect 10994 -3997 11046 -3924
rect 11101 -3890 11154 -3867
rect 11101 -3924 11109 -3890
rect 11143 -3924 11154 -3890
rect 11101 -3997 11154 -3924
rect 11254 -3890 11319 -3867
rect 11254 -3924 11265 -3890
rect 11299 -3924 11319 -3890
rect 11254 -3951 11319 -3924
rect 11349 -3890 11420 -3867
rect 11349 -3924 11363 -3890
rect 11397 -3924 11420 -3890
rect 11349 -3951 11420 -3924
rect 11254 -3997 11304 -3951
rect 11658 -3905 11710 -3867
rect 11658 -3939 11666 -3905
rect 11700 -3939 11710 -3905
rect 11658 -3977 11710 -3939
rect 11920 -3905 11972 -3867
rect 12567 -3881 12633 -3867
rect 11920 -3939 11930 -3905
rect 11964 -3939 11972 -3905
rect 11920 -3977 11972 -3939
rect 12567 -3915 12588 -3881
rect 12622 -3915 12633 -3881
rect 12567 -3951 12633 -3915
rect 12663 -3892 12719 -3867
rect 12663 -3926 12674 -3892
rect 12708 -3926 12719 -3892
rect 12663 -3951 12719 -3926
rect 12749 -3881 12805 -3867
rect 12749 -3915 12760 -3881
rect 12794 -3915 12805 -3881
rect 12749 -3951 12805 -3915
rect 12835 -3892 12891 -3867
rect 12835 -3926 12846 -3892
rect 12880 -3926 12891 -3892
rect 12835 -3951 12891 -3926
rect 12921 -3881 13000 -3867
rect 12921 -3915 12932 -3881
rect 12966 -3915 13000 -3881
rect 12921 -3951 13000 -3915
rect 13222 -3905 13274 -3867
rect 13222 -3939 13230 -3905
rect 13264 -3939 13274 -3905
rect 13222 -3977 13274 -3939
rect 13484 -3905 13536 -3867
rect 13682 -3879 13735 -3867
rect 13484 -3939 13494 -3905
rect 13528 -3939 13536 -3905
rect 13484 -3977 13536 -3939
rect 13682 -3913 13690 -3879
rect 13724 -3913 13735 -3879
rect 13682 -3951 13735 -3913
rect 13765 -3892 13821 -3867
rect 13765 -3926 13776 -3892
rect 13810 -3926 13821 -3892
rect 13765 -3951 13821 -3926
rect 13851 -3892 13907 -3867
rect 13851 -3926 13862 -3892
rect 13896 -3926 13907 -3892
rect 13851 -3951 13907 -3926
rect 13937 -3892 13993 -3867
rect 13937 -3926 13948 -3892
rect 13982 -3926 13993 -3892
rect 13937 -3951 13993 -3926
rect 14023 -3892 14079 -3867
rect 14023 -3926 14034 -3892
rect 14068 -3926 14079 -3892
rect 14023 -3951 14079 -3926
rect 14109 -3892 14165 -3867
rect 14109 -3926 14120 -3892
rect 14154 -3926 14165 -3892
rect 14109 -3951 14165 -3926
rect 14195 -3883 14251 -3867
rect 14195 -3917 14206 -3883
rect 14240 -3917 14251 -3883
rect 14195 -3951 14251 -3917
rect 14281 -3892 14337 -3867
rect 14281 -3926 14292 -3892
rect 14326 -3926 14337 -3892
rect 14281 -3951 14337 -3926
rect 14367 -3883 14423 -3867
rect 14367 -3917 14378 -3883
rect 14412 -3917 14423 -3883
rect 14367 -3951 14423 -3917
rect 14453 -3892 14509 -3867
rect 14453 -3926 14464 -3892
rect 14498 -3926 14509 -3892
rect 14453 -3951 14509 -3926
rect 14539 -3883 14595 -3867
rect 14539 -3917 14550 -3883
rect 14584 -3917 14595 -3883
rect 14539 -3951 14595 -3917
rect 14625 -3892 14681 -3867
rect 14625 -3926 14636 -3892
rect 14670 -3926 14681 -3892
rect 14625 -3951 14681 -3926
rect 14711 -3883 14766 -3867
rect 14711 -3917 14722 -3883
rect 14756 -3917 14766 -3883
rect 14711 -3951 14766 -3917
rect 14796 -3892 14852 -3867
rect 14796 -3926 14807 -3892
rect 14841 -3926 14852 -3892
rect 14796 -3951 14852 -3926
rect 14882 -3883 14938 -3867
rect 14882 -3917 14893 -3883
rect 14927 -3917 14938 -3883
rect 14882 -3951 14938 -3917
rect 14968 -3892 15024 -3867
rect 14968 -3926 14979 -3892
rect 15013 -3926 15024 -3892
rect 14968 -3951 15024 -3926
rect 15054 -3883 15110 -3867
rect 15054 -3917 15065 -3883
rect 15099 -3917 15110 -3883
rect 15054 -3951 15110 -3917
rect 15140 -3892 15196 -3867
rect 15140 -3926 15151 -3892
rect 15185 -3926 15196 -3892
rect 15140 -3951 15196 -3926
rect 15226 -3883 15282 -3867
rect 15226 -3917 15237 -3883
rect 15271 -3917 15282 -3883
rect 15226 -3951 15282 -3917
rect 15312 -3892 15368 -3867
rect 15312 -3926 15323 -3892
rect 15357 -3926 15368 -3892
rect 15312 -3951 15368 -3926
rect 15398 -3883 15451 -3867
rect 15398 -3917 15409 -3883
rect 15443 -3917 15451 -3883
rect 15398 -3951 15451 -3917
rect 15614 -3898 15666 -3867
rect 15614 -3932 15622 -3898
rect 15656 -3932 15666 -3898
rect 15614 -3977 15666 -3932
rect 16612 -3898 16664 -3867
rect 16612 -3932 16622 -3898
rect 16656 -3932 16664 -3898
rect 16612 -3977 16664 -3932
rect -2970 -4796 -2918 -4751
rect -2970 -4830 -2962 -4796
rect -2928 -4830 -2918 -4796
rect -2970 -4861 -2918 -4830
rect -2340 -4796 -2288 -4751
rect -2340 -4830 -2330 -4796
rect -2296 -4830 -2288 -4796
rect -2340 -4861 -2288 -4830
rect -1590 -4796 -1538 -4751
rect -1590 -4830 -1582 -4796
rect -1548 -4830 -1538 -4796
rect -1590 -4861 -1538 -4830
rect -960 -4796 -908 -4751
rect -738 -4777 -688 -4731
rect -960 -4830 -950 -4796
rect -916 -4830 -908 -4796
rect -960 -4861 -908 -4830
rect -854 -4804 -783 -4777
rect -854 -4838 -831 -4804
rect -797 -4838 -783 -4804
rect -854 -4861 -783 -4838
rect -753 -4804 -688 -4777
rect -753 -4838 -733 -4804
rect -699 -4838 -688 -4804
rect -753 -4861 -688 -4838
rect -588 -4804 -535 -4731
rect -588 -4838 -577 -4804
rect -543 -4838 -535 -4804
rect -588 -4861 -535 -4838
rect -480 -4804 -428 -4731
rect -480 -4838 -472 -4804
rect -438 -4838 -428 -4804
rect -480 -4861 -428 -4838
rect -328 -4777 -278 -4731
rect -328 -4804 -256 -4777
rect -328 -4838 -312 -4804
rect -278 -4838 -256 -4804
rect -328 -4861 -256 -4838
rect -226 -4804 -172 -4777
rect -226 -4838 -215 -4804
rect -181 -4838 -172 -4804
rect -226 -4861 -172 -4838
rect -26 -4789 26 -4751
rect -26 -4823 -18 -4789
rect 16 -4823 26 -4789
rect -26 -4861 26 -4823
rect 236 -4789 288 -4751
rect 236 -4823 246 -4789
rect 280 -4823 288 -4789
rect 236 -4861 288 -4823
rect 550 -4777 600 -4731
rect 434 -4804 505 -4777
rect 434 -4838 457 -4804
rect 491 -4838 505 -4804
rect 434 -4861 505 -4838
rect 535 -4804 600 -4777
rect 535 -4838 555 -4804
rect 589 -4838 600 -4804
rect 535 -4861 600 -4838
rect 700 -4804 753 -4731
rect 700 -4838 711 -4804
rect 745 -4838 753 -4804
rect 700 -4861 753 -4838
rect 808 -4804 860 -4731
rect 808 -4838 816 -4804
rect 850 -4838 860 -4804
rect 808 -4861 860 -4838
rect 960 -4777 1010 -4731
rect 960 -4804 1032 -4777
rect 960 -4838 976 -4804
rect 1010 -4838 1032 -4804
rect 960 -4861 1032 -4838
rect 1062 -4804 1116 -4777
rect 1062 -4838 1073 -4804
rect 1107 -4838 1116 -4804
rect 1062 -4861 1116 -4838
rect 1262 -4789 1314 -4751
rect 1262 -4823 1270 -4789
rect 1304 -4823 1314 -4789
rect 1262 -4861 1314 -4823
rect 1524 -4789 1576 -4751
rect 1524 -4823 1534 -4789
rect 1568 -4823 1576 -4789
rect 1524 -4861 1576 -4823
rect 1722 -4796 1774 -4751
rect 1722 -4830 1730 -4796
rect 1764 -4830 1774 -4796
rect 1722 -4861 1774 -4830
rect 2352 -4796 2404 -4751
rect 2352 -4830 2362 -4796
rect 2396 -4830 2404 -4796
rect 2352 -4861 2404 -4830
rect 2550 -4789 2602 -4751
rect 2550 -4823 2558 -4789
rect 2592 -4823 2602 -4789
rect 2550 -4861 2602 -4823
rect 2812 -4789 2864 -4751
rect 2812 -4823 2822 -4789
rect 2856 -4823 2864 -4789
rect 2812 -4861 2864 -4823
rect 3126 -4777 3176 -4731
rect 3010 -4804 3081 -4777
rect 3010 -4838 3033 -4804
rect 3067 -4838 3081 -4804
rect 3010 -4861 3081 -4838
rect 3111 -4804 3176 -4777
rect 3111 -4838 3131 -4804
rect 3165 -4838 3176 -4804
rect 3111 -4861 3176 -4838
rect 3276 -4804 3329 -4731
rect 3276 -4838 3287 -4804
rect 3321 -4838 3329 -4804
rect 3276 -4861 3329 -4838
rect 3384 -4804 3436 -4731
rect 3384 -4838 3392 -4804
rect 3426 -4838 3436 -4804
rect 3384 -4861 3436 -4838
rect 3536 -4777 3586 -4731
rect 3536 -4804 3608 -4777
rect 3536 -4838 3552 -4804
rect 3586 -4838 3608 -4804
rect 3536 -4861 3608 -4838
rect 3638 -4804 3692 -4777
rect 3638 -4838 3649 -4804
rect 3683 -4838 3692 -4804
rect 3638 -4861 3692 -4838
rect 3838 -4789 3890 -4751
rect 3838 -4823 3846 -4789
rect 3880 -4823 3890 -4789
rect 3838 -4861 3890 -4823
rect 4100 -4789 4152 -4751
rect 4100 -4823 4110 -4789
rect 4144 -4823 4152 -4789
rect 4100 -4861 4152 -4823
rect 4298 -4796 4350 -4751
rect 4298 -4830 4306 -4796
rect 4340 -4830 4350 -4796
rect 4298 -4861 4350 -4830
rect 4928 -4796 4980 -4751
rect 4928 -4830 4938 -4796
rect 4972 -4830 4980 -4796
rect 4928 -4861 4980 -4830
rect 5126 -4789 5178 -4751
rect 5126 -4823 5134 -4789
rect 5168 -4823 5178 -4789
rect 5126 -4861 5178 -4823
rect 5388 -4789 5440 -4751
rect 5388 -4823 5398 -4789
rect 5432 -4823 5440 -4789
rect 5388 -4861 5440 -4823
rect 5702 -4777 5752 -4731
rect 5586 -4804 5657 -4777
rect 5586 -4838 5609 -4804
rect 5643 -4838 5657 -4804
rect 5586 -4861 5657 -4838
rect 5687 -4804 5752 -4777
rect 5687 -4838 5707 -4804
rect 5741 -4838 5752 -4804
rect 5687 -4861 5752 -4838
rect 5852 -4804 5905 -4731
rect 5852 -4838 5863 -4804
rect 5897 -4838 5905 -4804
rect 5852 -4861 5905 -4838
rect 5960 -4804 6012 -4731
rect 5960 -4838 5968 -4804
rect 6002 -4838 6012 -4804
rect 5960 -4861 6012 -4838
rect 6112 -4777 6162 -4731
rect 6112 -4804 6184 -4777
rect 6112 -4838 6128 -4804
rect 6162 -4838 6184 -4804
rect 6112 -4861 6184 -4838
rect 6214 -4804 6268 -4777
rect 6214 -4838 6225 -4804
rect 6259 -4838 6268 -4804
rect 6214 -4861 6268 -4838
rect 6414 -4789 6466 -4751
rect 6414 -4823 6422 -4789
rect 6456 -4823 6466 -4789
rect 6414 -4861 6466 -4823
rect 6676 -4789 6728 -4751
rect 6676 -4823 6686 -4789
rect 6720 -4823 6728 -4789
rect 6676 -4861 6728 -4823
rect 6874 -4796 6926 -4751
rect 6874 -4830 6882 -4796
rect 6916 -4830 6926 -4796
rect 6874 -4861 6926 -4830
rect 7504 -4796 7556 -4751
rect 7504 -4830 7514 -4796
rect 7548 -4830 7556 -4796
rect 7504 -4861 7556 -4830
rect 7702 -4789 7754 -4751
rect 7702 -4823 7710 -4789
rect 7744 -4823 7754 -4789
rect 7702 -4861 7754 -4823
rect 7964 -4789 8016 -4751
rect 7964 -4823 7974 -4789
rect 8008 -4823 8016 -4789
rect 7964 -4861 8016 -4823
rect 8278 -4777 8328 -4731
rect 8162 -4804 8233 -4777
rect 8162 -4838 8185 -4804
rect 8219 -4838 8233 -4804
rect 8162 -4861 8233 -4838
rect 8263 -4804 8328 -4777
rect 8263 -4838 8283 -4804
rect 8317 -4838 8328 -4804
rect 8263 -4861 8328 -4838
rect 8428 -4804 8481 -4731
rect 8428 -4838 8439 -4804
rect 8473 -4838 8481 -4804
rect 8428 -4861 8481 -4838
rect 8536 -4804 8588 -4731
rect 8536 -4838 8544 -4804
rect 8578 -4838 8588 -4804
rect 8536 -4861 8588 -4838
rect 8688 -4777 8738 -4731
rect 8688 -4804 8760 -4777
rect 8688 -4838 8704 -4804
rect 8738 -4838 8760 -4804
rect 8688 -4861 8760 -4838
rect 8790 -4804 8844 -4777
rect 8790 -4838 8801 -4804
rect 8835 -4838 8844 -4804
rect 8790 -4861 8844 -4838
rect 8990 -4789 9042 -4751
rect 8990 -4823 8998 -4789
rect 9032 -4823 9042 -4789
rect 8990 -4861 9042 -4823
rect 9252 -4789 9304 -4751
rect 9252 -4823 9262 -4789
rect 9296 -4823 9304 -4789
rect 9252 -4861 9304 -4823
rect 9450 -4796 9502 -4751
rect 9450 -4830 9458 -4796
rect 9492 -4830 9502 -4796
rect 9450 -4861 9502 -4830
rect 10080 -4796 10132 -4751
rect 10080 -4830 10090 -4796
rect 10124 -4830 10132 -4796
rect 10080 -4861 10132 -4830
rect 10370 -4789 10422 -4751
rect 10370 -4823 10378 -4789
rect 10412 -4823 10422 -4789
rect 10370 -4861 10422 -4823
rect 10632 -4789 10684 -4751
rect 10854 -4777 10904 -4731
rect 10632 -4823 10642 -4789
rect 10676 -4823 10684 -4789
rect 10632 -4861 10684 -4823
rect 10738 -4804 10809 -4777
rect 10738 -4838 10761 -4804
rect 10795 -4838 10809 -4804
rect 10738 -4861 10809 -4838
rect 10839 -4804 10904 -4777
rect 10839 -4838 10859 -4804
rect 10893 -4838 10904 -4804
rect 10839 -4861 10904 -4838
rect 11004 -4804 11057 -4731
rect 11004 -4838 11015 -4804
rect 11049 -4838 11057 -4804
rect 11004 -4861 11057 -4838
rect 11112 -4804 11164 -4731
rect 11112 -4838 11120 -4804
rect 11154 -4838 11164 -4804
rect 11112 -4861 11164 -4838
rect 11264 -4777 11314 -4731
rect 11264 -4804 11336 -4777
rect 11264 -4838 11280 -4804
rect 11314 -4838 11336 -4804
rect 11264 -4861 11336 -4838
rect 11366 -4804 11420 -4777
rect 11366 -4838 11377 -4804
rect 11411 -4838 11420 -4804
rect 11366 -4861 11420 -4838
rect 11658 -4789 11710 -4751
rect 11658 -4823 11666 -4789
rect 11700 -4823 11710 -4789
rect 11658 -4861 11710 -4823
rect 11920 -4789 11972 -4751
rect 11920 -4823 11930 -4789
rect 11964 -4823 11972 -4789
rect 11920 -4861 11972 -4823
rect 13682 -4815 13735 -4777
rect 13682 -4849 13690 -4815
rect 13724 -4849 13735 -4815
rect 13682 -4861 13735 -4849
rect 13765 -4802 13821 -4777
rect 13765 -4836 13776 -4802
rect 13810 -4836 13821 -4802
rect 13765 -4861 13821 -4836
rect 13851 -4802 13907 -4777
rect 13851 -4836 13862 -4802
rect 13896 -4836 13907 -4802
rect 13851 -4861 13907 -4836
rect 13937 -4802 13993 -4777
rect 13937 -4836 13948 -4802
rect 13982 -4836 13993 -4802
rect 13937 -4861 13993 -4836
rect 14023 -4802 14079 -4777
rect 14023 -4836 14034 -4802
rect 14068 -4836 14079 -4802
rect 14023 -4861 14079 -4836
rect 14109 -4802 14165 -4777
rect 14109 -4836 14120 -4802
rect 14154 -4836 14165 -4802
rect 14109 -4861 14165 -4836
rect 14195 -4811 14251 -4777
rect 14195 -4845 14206 -4811
rect 14240 -4845 14251 -4811
rect 14195 -4861 14251 -4845
rect 14281 -4802 14337 -4777
rect 14281 -4836 14292 -4802
rect 14326 -4836 14337 -4802
rect 14281 -4861 14337 -4836
rect 14367 -4811 14423 -4777
rect 14367 -4845 14378 -4811
rect 14412 -4845 14423 -4811
rect 14367 -4861 14423 -4845
rect 14453 -4802 14509 -4777
rect 14453 -4836 14464 -4802
rect 14498 -4836 14509 -4802
rect 14453 -4861 14509 -4836
rect 14539 -4811 14595 -4777
rect 14539 -4845 14550 -4811
rect 14584 -4845 14595 -4811
rect 14539 -4861 14595 -4845
rect 14625 -4802 14681 -4777
rect 14625 -4836 14636 -4802
rect 14670 -4836 14681 -4802
rect 14625 -4861 14681 -4836
rect 14711 -4811 14766 -4777
rect 14711 -4845 14722 -4811
rect 14756 -4845 14766 -4811
rect 14711 -4861 14766 -4845
rect 14796 -4802 14852 -4777
rect 14796 -4836 14807 -4802
rect 14841 -4836 14852 -4802
rect 14796 -4861 14852 -4836
rect 14882 -4811 14938 -4777
rect 14882 -4845 14893 -4811
rect 14927 -4845 14938 -4811
rect 14882 -4861 14938 -4845
rect 14968 -4802 15024 -4777
rect 14968 -4836 14979 -4802
rect 15013 -4836 15024 -4802
rect 14968 -4861 15024 -4836
rect 15054 -4811 15110 -4777
rect 15054 -4845 15065 -4811
rect 15099 -4845 15110 -4811
rect 15054 -4861 15110 -4845
rect 15140 -4802 15196 -4777
rect 15140 -4836 15151 -4802
rect 15185 -4836 15196 -4802
rect 15140 -4861 15196 -4836
rect 15226 -4811 15282 -4777
rect 15226 -4845 15237 -4811
rect 15271 -4845 15282 -4811
rect 15226 -4861 15282 -4845
rect 15312 -4802 15368 -4777
rect 15312 -4836 15323 -4802
rect 15357 -4836 15368 -4802
rect 15312 -4861 15368 -4836
rect 15398 -4811 15451 -4777
rect 15398 -4845 15409 -4811
rect 15443 -4845 15451 -4811
rect 15614 -4796 15666 -4751
rect 15614 -4830 15622 -4796
rect 15656 -4830 15666 -4796
rect 15398 -4861 15451 -4845
rect 15614 -4861 15666 -4830
rect 16612 -4796 16664 -4751
rect 16612 -4830 16622 -4796
rect 16656 -4830 16664 -4796
rect 16612 -4861 16664 -4830
rect -2970 -4986 -2918 -4955
rect -2970 -5020 -2962 -4986
rect -2928 -5020 -2918 -4986
rect -2970 -5065 -2918 -5020
rect -2340 -4986 -2288 -4955
rect -2340 -5020 -2330 -4986
rect -2296 -5020 -2288 -4986
rect -2340 -5065 -2288 -5020
rect -1590 -4986 -1538 -4955
rect -1590 -5020 -1582 -4986
rect -1548 -5020 -1538 -4986
rect -1590 -5065 -1538 -5020
rect -960 -4986 -908 -4955
rect -960 -5020 -950 -4986
rect -916 -5020 -908 -4986
rect -960 -5065 -908 -5020
rect -854 -4986 -802 -4955
rect -854 -5020 -846 -4986
rect -812 -5020 -802 -4986
rect -854 -5065 -802 -5020
rect -224 -4986 -172 -4955
rect -224 -5020 -214 -4986
rect -180 -5020 -172 -4986
rect -224 -5065 -172 -5020
rect -26 -4993 26 -4955
rect -26 -5027 -18 -4993
rect 16 -5027 26 -4993
rect -26 -5065 26 -5027
rect 236 -4993 288 -4955
rect 236 -5027 246 -4993
rect 280 -5027 288 -4993
rect 236 -5065 288 -5027
rect 434 -4978 488 -4955
rect 434 -5012 443 -4978
rect 477 -5012 488 -4978
rect 434 -5039 488 -5012
rect 518 -4978 590 -4955
rect 518 -5012 540 -4978
rect 574 -5012 590 -4978
rect 518 -5039 590 -5012
rect 540 -5085 590 -5039
rect 690 -4978 742 -4955
rect 690 -5012 700 -4978
rect 734 -5012 742 -4978
rect 690 -5085 742 -5012
rect 797 -4978 850 -4955
rect 797 -5012 805 -4978
rect 839 -5012 850 -4978
rect 797 -5085 850 -5012
rect 950 -4978 1015 -4955
rect 950 -5012 961 -4978
rect 995 -5012 1015 -4978
rect 950 -5039 1015 -5012
rect 1045 -4978 1116 -4955
rect 1045 -5012 1059 -4978
rect 1093 -5012 1116 -4978
rect 1045 -5039 1116 -5012
rect 950 -5085 1000 -5039
rect 1262 -4993 1314 -4955
rect 1262 -5027 1270 -4993
rect 1304 -5027 1314 -4993
rect 1262 -5065 1314 -5027
rect 1524 -4993 1576 -4955
rect 1524 -5027 1534 -4993
rect 1568 -5027 1576 -4993
rect 1524 -5065 1576 -5027
rect 1722 -4986 1774 -4955
rect 1722 -5020 1730 -4986
rect 1764 -5020 1774 -4986
rect 1722 -5065 1774 -5020
rect 2352 -4986 2404 -4955
rect 2352 -5020 2362 -4986
rect 2396 -5020 2404 -4986
rect 2352 -5065 2404 -5020
rect 2550 -4993 2602 -4955
rect 2550 -5027 2558 -4993
rect 2592 -5027 2602 -4993
rect 2550 -5065 2602 -5027
rect 2812 -4993 2864 -4955
rect 2812 -5027 2822 -4993
rect 2856 -5027 2864 -4993
rect 2812 -5065 2864 -5027
rect 3010 -4978 3064 -4955
rect 3010 -5012 3019 -4978
rect 3053 -5012 3064 -4978
rect 3010 -5039 3064 -5012
rect 3094 -4978 3166 -4955
rect 3094 -5012 3116 -4978
rect 3150 -5012 3166 -4978
rect 3094 -5039 3166 -5012
rect 3116 -5085 3166 -5039
rect 3266 -4978 3318 -4955
rect 3266 -5012 3276 -4978
rect 3310 -5012 3318 -4978
rect 3266 -5085 3318 -5012
rect 3373 -4978 3426 -4955
rect 3373 -5012 3381 -4978
rect 3415 -5012 3426 -4978
rect 3373 -5085 3426 -5012
rect 3526 -4978 3591 -4955
rect 3526 -5012 3537 -4978
rect 3571 -5012 3591 -4978
rect 3526 -5039 3591 -5012
rect 3621 -4978 3692 -4955
rect 3621 -5012 3635 -4978
rect 3669 -5012 3692 -4978
rect 3621 -5039 3692 -5012
rect 3526 -5085 3576 -5039
rect 3838 -4993 3890 -4955
rect 3838 -5027 3846 -4993
rect 3880 -5027 3890 -4993
rect 3838 -5065 3890 -5027
rect 4100 -4993 4152 -4955
rect 4100 -5027 4110 -4993
rect 4144 -5027 4152 -4993
rect 4100 -5065 4152 -5027
rect 4298 -4986 4350 -4955
rect 4298 -5020 4306 -4986
rect 4340 -5020 4350 -4986
rect 4298 -5065 4350 -5020
rect 4928 -4986 4980 -4955
rect 4928 -5020 4938 -4986
rect 4972 -5020 4980 -4986
rect 4928 -5065 4980 -5020
rect 5126 -4993 5178 -4955
rect 5126 -5027 5134 -4993
rect 5168 -5027 5178 -4993
rect 5126 -5065 5178 -5027
rect 5388 -4993 5440 -4955
rect 5388 -5027 5398 -4993
rect 5432 -5027 5440 -4993
rect 5388 -5065 5440 -5027
rect 5586 -4978 5640 -4955
rect 5586 -5012 5595 -4978
rect 5629 -5012 5640 -4978
rect 5586 -5039 5640 -5012
rect 5670 -4978 5742 -4955
rect 5670 -5012 5692 -4978
rect 5726 -5012 5742 -4978
rect 5670 -5039 5742 -5012
rect 5692 -5085 5742 -5039
rect 5842 -4978 5894 -4955
rect 5842 -5012 5852 -4978
rect 5886 -5012 5894 -4978
rect 5842 -5085 5894 -5012
rect 5949 -4978 6002 -4955
rect 5949 -5012 5957 -4978
rect 5991 -5012 6002 -4978
rect 5949 -5085 6002 -5012
rect 6102 -4978 6167 -4955
rect 6102 -5012 6113 -4978
rect 6147 -5012 6167 -4978
rect 6102 -5039 6167 -5012
rect 6197 -4978 6268 -4955
rect 6197 -5012 6211 -4978
rect 6245 -5012 6268 -4978
rect 6197 -5039 6268 -5012
rect 6102 -5085 6152 -5039
rect 6414 -4993 6466 -4955
rect 6414 -5027 6422 -4993
rect 6456 -5027 6466 -4993
rect 6414 -5065 6466 -5027
rect 6676 -4993 6728 -4955
rect 6676 -5027 6686 -4993
rect 6720 -5027 6728 -4993
rect 6676 -5065 6728 -5027
rect 6874 -4986 6926 -4955
rect 6874 -5020 6882 -4986
rect 6916 -5020 6926 -4986
rect 6874 -5065 6926 -5020
rect 7504 -4986 7556 -4955
rect 7504 -5020 7514 -4986
rect 7548 -5020 7556 -4986
rect 7504 -5065 7556 -5020
rect 7702 -4993 7754 -4955
rect 7702 -5027 7710 -4993
rect 7744 -5027 7754 -4993
rect 7702 -5065 7754 -5027
rect 7964 -4993 8016 -4955
rect 7964 -5027 7974 -4993
rect 8008 -5027 8016 -4993
rect 7964 -5065 8016 -5027
rect 8162 -4978 8216 -4955
rect 8162 -5012 8171 -4978
rect 8205 -5012 8216 -4978
rect 8162 -5039 8216 -5012
rect 8246 -4978 8318 -4955
rect 8246 -5012 8268 -4978
rect 8302 -5012 8318 -4978
rect 8246 -5039 8318 -5012
rect 8268 -5085 8318 -5039
rect 8418 -4978 8470 -4955
rect 8418 -5012 8428 -4978
rect 8462 -5012 8470 -4978
rect 8418 -5085 8470 -5012
rect 8525 -4978 8578 -4955
rect 8525 -5012 8533 -4978
rect 8567 -5012 8578 -4978
rect 8525 -5085 8578 -5012
rect 8678 -4978 8743 -4955
rect 8678 -5012 8689 -4978
rect 8723 -5012 8743 -4978
rect 8678 -5039 8743 -5012
rect 8773 -4978 8844 -4955
rect 8773 -5012 8787 -4978
rect 8821 -5012 8844 -4978
rect 8773 -5039 8844 -5012
rect 8678 -5085 8728 -5039
rect 8990 -4993 9042 -4955
rect 8990 -5027 8998 -4993
rect 9032 -5027 9042 -4993
rect 8990 -5065 9042 -5027
rect 9252 -4993 9304 -4955
rect 9252 -5027 9262 -4993
rect 9296 -5027 9304 -4993
rect 9252 -5065 9304 -5027
rect 9450 -4986 9502 -4955
rect 9450 -5020 9458 -4986
rect 9492 -5020 9502 -4986
rect 9450 -5065 9502 -5020
rect 10080 -4986 10132 -4955
rect 10080 -5020 10090 -4986
rect 10124 -5020 10132 -4986
rect 10080 -5065 10132 -5020
rect 10370 -4993 10422 -4955
rect 10370 -5027 10378 -4993
rect 10412 -5027 10422 -4993
rect 10370 -5065 10422 -5027
rect 10632 -4993 10684 -4955
rect 10632 -5027 10642 -4993
rect 10676 -5027 10684 -4993
rect 10632 -5065 10684 -5027
rect 10738 -4978 10792 -4955
rect 10738 -5012 10747 -4978
rect 10781 -5012 10792 -4978
rect 10738 -5039 10792 -5012
rect 10822 -4978 10894 -4955
rect 10822 -5012 10844 -4978
rect 10878 -5012 10894 -4978
rect 10822 -5039 10894 -5012
rect 10844 -5085 10894 -5039
rect 10994 -4978 11046 -4955
rect 10994 -5012 11004 -4978
rect 11038 -5012 11046 -4978
rect 10994 -5085 11046 -5012
rect 11101 -4978 11154 -4955
rect 11101 -5012 11109 -4978
rect 11143 -5012 11154 -4978
rect 11101 -5085 11154 -5012
rect 11254 -4978 11319 -4955
rect 11254 -5012 11265 -4978
rect 11299 -5012 11319 -4978
rect 11254 -5039 11319 -5012
rect 11349 -4978 11420 -4955
rect 11349 -5012 11363 -4978
rect 11397 -5012 11420 -4978
rect 11349 -5039 11420 -5012
rect 11254 -5085 11304 -5039
rect 11658 -4993 11710 -4955
rect 11658 -5027 11666 -4993
rect 11700 -5027 11710 -4993
rect 11658 -5065 11710 -5027
rect 11920 -4993 11972 -4955
rect 12567 -4969 12633 -4955
rect 11920 -5027 11930 -4993
rect 11964 -5027 11972 -4993
rect 11920 -5065 11972 -5027
rect 12567 -5003 12588 -4969
rect 12622 -5003 12633 -4969
rect 12567 -5039 12633 -5003
rect 12663 -4980 12719 -4955
rect 12663 -5014 12674 -4980
rect 12708 -5014 12719 -4980
rect 12663 -5039 12719 -5014
rect 12749 -4969 12805 -4955
rect 12749 -5003 12760 -4969
rect 12794 -5003 12805 -4969
rect 12749 -5039 12805 -5003
rect 12835 -4980 12891 -4955
rect 12835 -5014 12846 -4980
rect 12880 -5014 12891 -4980
rect 12835 -5039 12891 -5014
rect 12921 -4969 13000 -4955
rect 12921 -5003 12932 -4969
rect 12966 -5003 13000 -4969
rect 12921 -5039 13000 -5003
rect 13222 -4993 13274 -4955
rect 13222 -5027 13230 -4993
rect 13264 -5027 13274 -4993
rect 13222 -5065 13274 -5027
rect 13484 -4993 13536 -4955
rect 13682 -4967 13735 -4955
rect 13484 -5027 13494 -4993
rect 13528 -5027 13536 -4993
rect 13484 -5065 13536 -5027
rect 13682 -5001 13690 -4967
rect 13724 -5001 13735 -4967
rect 13682 -5039 13735 -5001
rect 13765 -4980 13821 -4955
rect 13765 -5014 13776 -4980
rect 13810 -5014 13821 -4980
rect 13765 -5039 13821 -5014
rect 13851 -4980 13907 -4955
rect 13851 -5014 13862 -4980
rect 13896 -5014 13907 -4980
rect 13851 -5039 13907 -5014
rect 13937 -4980 13993 -4955
rect 13937 -5014 13948 -4980
rect 13982 -5014 13993 -4980
rect 13937 -5039 13993 -5014
rect 14023 -4980 14079 -4955
rect 14023 -5014 14034 -4980
rect 14068 -5014 14079 -4980
rect 14023 -5039 14079 -5014
rect 14109 -4980 14165 -4955
rect 14109 -5014 14120 -4980
rect 14154 -5014 14165 -4980
rect 14109 -5039 14165 -5014
rect 14195 -4971 14251 -4955
rect 14195 -5005 14206 -4971
rect 14240 -5005 14251 -4971
rect 14195 -5039 14251 -5005
rect 14281 -4980 14337 -4955
rect 14281 -5014 14292 -4980
rect 14326 -5014 14337 -4980
rect 14281 -5039 14337 -5014
rect 14367 -4971 14423 -4955
rect 14367 -5005 14378 -4971
rect 14412 -5005 14423 -4971
rect 14367 -5039 14423 -5005
rect 14453 -4980 14509 -4955
rect 14453 -5014 14464 -4980
rect 14498 -5014 14509 -4980
rect 14453 -5039 14509 -5014
rect 14539 -4971 14595 -4955
rect 14539 -5005 14550 -4971
rect 14584 -5005 14595 -4971
rect 14539 -5039 14595 -5005
rect 14625 -4980 14681 -4955
rect 14625 -5014 14636 -4980
rect 14670 -5014 14681 -4980
rect 14625 -5039 14681 -5014
rect 14711 -4971 14766 -4955
rect 14711 -5005 14722 -4971
rect 14756 -5005 14766 -4971
rect 14711 -5039 14766 -5005
rect 14796 -4980 14852 -4955
rect 14796 -5014 14807 -4980
rect 14841 -5014 14852 -4980
rect 14796 -5039 14852 -5014
rect 14882 -4971 14938 -4955
rect 14882 -5005 14893 -4971
rect 14927 -5005 14938 -4971
rect 14882 -5039 14938 -5005
rect 14968 -4980 15024 -4955
rect 14968 -5014 14979 -4980
rect 15013 -5014 15024 -4980
rect 14968 -5039 15024 -5014
rect 15054 -4971 15110 -4955
rect 15054 -5005 15065 -4971
rect 15099 -5005 15110 -4971
rect 15054 -5039 15110 -5005
rect 15140 -4980 15196 -4955
rect 15140 -5014 15151 -4980
rect 15185 -5014 15196 -4980
rect 15140 -5039 15196 -5014
rect 15226 -4971 15282 -4955
rect 15226 -5005 15237 -4971
rect 15271 -5005 15282 -4971
rect 15226 -5039 15282 -5005
rect 15312 -4980 15368 -4955
rect 15312 -5014 15323 -4980
rect 15357 -5014 15368 -4980
rect 15312 -5039 15368 -5014
rect 15398 -4971 15451 -4955
rect 15398 -5005 15409 -4971
rect 15443 -5005 15451 -4971
rect 15398 -5039 15451 -5005
rect 15614 -4986 15666 -4955
rect 15614 -5020 15622 -4986
rect 15656 -5020 15666 -4986
rect 15614 -5065 15666 -5020
rect 16612 -4986 16664 -4955
rect 16612 -5020 16622 -4986
rect 16656 -5020 16664 -4986
rect 16612 -5065 16664 -5020
rect -2970 -5884 -2918 -5839
rect -2970 -5918 -2962 -5884
rect -2928 -5918 -2918 -5884
rect -2970 -5949 -2918 -5918
rect -2340 -5884 -2288 -5839
rect -2340 -5918 -2330 -5884
rect -2296 -5918 -2288 -5884
rect -2340 -5949 -2288 -5918
rect -1590 -5884 -1538 -5839
rect -1590 -5918 -1582 -5884
rect -1548 -5918 -1538 -5884
rect -1590 -5949 -1538 -5918
rect -960 -5884 -908 -5839
rect -960 -5918 -950 -5884
rect -916 -5918 -908 -5884
rect -960 -5949 -908 -5918
rect -854 -5884 -802 -5839
rect -854 -5918 -846 -5884
rect -812 -5918 -802 -5884
rect -854 -5949 -802 -5918
rect -224 -5884 -172 -5839
rect -224 -5918 -214 -5884
rect -180 -5918 -172 -5884
rect -224 -5949 -172 -5918
rect -26 -5877 26 -5839
rect -26 -5911 -18 -5877
rect 16 -5911 26 -5877
rect -26 -5949 26 -5911
rect 236 -5877 288 -5839
rect 236 -5911 246 -5877
rect 280 -5911 288 -5877
rect 236 -5949 288 -5911
rect 550 -5865 600 -5819
rect 434 -5892 505 -5865
rect 434 -5926 457 -5892
rect 491 -5926 505 -5892
rect 434 -5949 505 -5926
rect 535 -5892 600 -5865
rect 535 -5926 555 -5892
rect 589 -5926 600 -5892
rect 535 -5949 600 -5926
rect 700 -5892 753 -5819
rect 700 -5926 711 -5892
rect 745 -5926 753 -5892
rect 700 -5949 753 -5926
rect 808 -5892 860 -5819
rect 808 -5926 816 -5892
rect 850 -5926 860 -5892
rect 808 -5949 860 -5926
rect 960 -5865 1010 -5819
rect 960 -5892 1032 -5865
rect 960 -5926 976 -5892
rect 1010 -5926 1032 -5892
rect 960 -5949 1032 -5926
rect 1062 -5892 1116 -5865
rect 1062 -5926 1073 -5892
rect 1107 -5926 1116 -5892
rect 1062 -5949 1116 -5926
rect 1262 -5877 1314 -5839
rect 1262 -5911 1270 -5877
rect 1304 -5911 1314 -5877
rect 1262 -5949 1314 -5911
rect 1524 -5877 1576 -5839
rect 1524 -5911 1534 -5877
rect 1568 -5911 1576 -5877
rect 1524 -5949 1576 -5911
rect 1722 -5884 1774 -5839
rect 1722 -5918 1730 -5884
rect 1764 -5918 1774 -5884
rect 1722 -5949 1774 -5918
rect 2352 -5884 2404 -5839
rect 2352 -5918 2362 -5884
rect 2396 -5918 2404 -5884
rect 2352 -5949 2404 -5918
rect 2550 -5877 2602 -5839
rect 2550 -5911 2558 -5877
rect 2592 -5911 2602 -5877
rect 2550 -5949 2602 -5911
rect 2812 -5877 2864 -5839
rect 2812 -5911 2822 -5877
rect 2856 -5911 2864 -5877
rect 2812 -5949 2864 -5911
rect 3126 -5865 3176 -5819
rect 3010 -5892 3081 -5865
rect 3010 -5926 3033 -5892
rect 3067 -5926 3081 -5892
rect 3010 -5949 3081 -5926
rect 3111 -5892 3176 -5865
rect 3111 -5926 3131 -5892
rect 3165 -5926 3176 -5892
rect 3111 -5949 3176 -5926
rect 3276 -5892 3329 -5819
rect 3276 -5926 3287 -5892
rect 3321 -5926 3329 -5892
rect 3276 -5949 3329 -5926
rect 3384 -5892 3436 -5819
rect 3384 -5926 3392 -5892
rect 3426 -5926 3436 -5892
rect 3384 -5949 3436 -5926
rect 3536 -5865 3586 -5819
rect 3536 -5892 3608 -5865
rect 3536 -5926 3552 -5892
rect 3586 -5926 3608 -5892
rect 3536 -5949 3608 -5926
rect 3638 -5892 3692 -5865
rect 3638 -5926 3649 -5892
rect 3683 -5926 3692 -5892
rect 3638 -5949 3692 -5926
rect 3838 -5877 3890 -5839
rect 3838 -5911 3846 -5877
rect 3880 -5911 3890 -5877
rect 3838 -5949 3890 -5911
rect 4100 -5877 4152 -5839
rect 4100 -5911 4110 -5877
rect 4144 -5911 4152 -5877
rect 4100 -5949 4152 -5911
rect 4298 -5884 4350 -5839
rect 4298 -5918 4306 -5884
rect 4340 -5918 4350 -5884
rect 4298 -5949 4350 -5918
rect 4928 -5884 4980 -5839
rect 4928 -5918 4938 -5884
rect 4972 -5918 4980 -5884
rect 4928 -5949 4980 -5918
rect 5126 -5877 5178 -5839
rect 5126 -5911 5134 -5877
rect 5168 -5911 5178 -5877
rect 5126 -5949 5178 -5911
rect 5388 -5877 5440 -5839
rect 5388 -5911 5398 -5877
rect 5432 -5911 5440 -5877
rect 5388 -5949 5440 -5911
rect 5702 -5865 5752 -5819
rect 5586 -5892 5657 -5865
rect 5586 -5926 5609 -5892
rect 5643 -5926 5657 -5892
rect 5586 -5949 5657 -5926
rect 5687 -5892 5752 -5865
rect 5687 -5926 5707 -5892
rect 5741 -5926 5752 -5892
rect 5687 -5949 5752 -5926
rect 5852 -5892 5905 -5819
rect 5852 -5926 5863 -5892
rect 5897 -5926 5905 -5892
rect 5852 -5949 5905 -5926
rect 5960 -5892 6012 -5819
rect 5960 -5926 5968 -5892
rect 6002 -5926 6012 -5892
rect 5960 -5949 6012 -5926
rect 6112 -5865 6162 -5819
rect 6112 -5892 6184 -5865
rect 6112 -5926 6128 -5892
rect 6162 -5926 6184 -5892
rect 6112 -5949 6184 -5926
rect 6214 -5892 6268 -5865
rect 6214 -5926 6225 -5892
rect 6259 -5926 6268 -5892
rect 6214 -5949 6268 -5926
rect 6414 -5877 6466 -5839
rect 6414 -5911 6422 -5877
rect 6456 -5911 6466 -5877
rect 6414 -5949 6466 -5911
rect 6676 -5877 6728 -5839
rect 6676 -5911 6686 -5877
rect 6720 -5911 6728 -5877
rect 6676 -5949 6728 -5911
rect 6874 -5884 6926 -5839
rect 6874 -5918 6882 -5884
rect 6916 -5918 6926 -5884
rect 6874 -5949 6926 -5918
rect 7504 -5884 7556 -5839
rect 7504 -5918 7514 -5884
rect 7548 -5918 7556 -5884
rect 7504 -5949 7556 -5918
rect 7702 -5877 7754 -5839
rect 7702 -5911 7710 -5877
rect 7744 -5911 7754 -5877
rect 7702 -5949 7754 -5911
rect 7964 -5877 8016 -5839
rect 7964 -5911 7974 -5877
rect 8008 -5911 8016 -5877
rect 7964 -5949 8016 -5911
rect 8278 -5865 8328 -5819
rect 8162 -5892 8233 -5865
rect 8162 -5926 8185 -5892
rect 8219 -5926 8233 -5892
rect 8162 -5949 8233 -5926
rect 8263 -5892 8328 -5865
rect 8263 -5926 8283 -5892
rect 8317 -5926 8328 -5892
rect 8263 -5949 8328 -5926
rect 8428 -5892 8481 -5819
rect 8428 -5926 8439 -5892
rect 8473 -5926 8481 -5892
rect 8428 -5949 8481 -5926
rect 8536 -5892 8588 -5819
rect 8536 -5926 8544 -5892
rect 8578 -5926 8588 -5892
rect 8536 -5949 8588 -5926
rect 8688 -5865 8738 -5819
rect 8688 -5892 8760 -5865
rect 8688 -5926 8704 -5892
rect 8738 -5926 8760 -5892
rect 8688 -5949 8760 -5926
rect 8790 -5892 8844 -5865
rect 8790 -5926 8801 -5892
rect 8835 -5926 8844 -5892
rect 8790 -5949 8844 -5926
rect 8990 -5877 9042 -5839
rect 8990 -5911 8998 -5877
rect 9032 -5911 9042 -5877
rect 8990 -5949 9042 -5911
rect 9252 -5877 9304 -5839
rect 9252 -5911 9262 -5877
rect 9296 -5911 9304 -5877
rect 9252 -5949 9304 -5911
rect 9450 -5884 9502 -5839
rect 9450 -5918 9458 -5884
rect 9492 -5918 9502 -5884
rect 9450 -5949 9502 -5918
rect 10080 -5884 10132 -5839
rect 10080 -5918 10090 -5884
rect 10124 -5918 10132 -5884
rect 10080 -5949 10132 -5918
rect 10370 -5877 10422 -5839
rect 10370 -5911 10378 -5877
rect 10412 -5911 10422 -5877
rect 10370 -5949 10422 -5911
rect 10632 -5877 10684 -5839
rect 10854 -5865 10904 -5819
rect 10632 -5911 10642 -5877
rect 10676 -5911 10684 -5877
rect 10632 -5949 10684 -5911
rect 10738 -5892 10809 -5865
rect 10738 -5926 10761 -5892
rect 10795 -5926 10809 -5892
rect 10738 -5949 10809 -5926
rect 10839 -5892 10904 -5865
rect 10839 -5926 10859 -5892
rect 10893 -5926 10904 -5892
rect 10839 -5949 10904 -5926
rect 11004 -5892 11057 -5819
rect 11004 -5926 11015 -5892
rect 11049 -5926 11057 -5892
rect 11004 -5949 11057 -5926
rect 11112 -5892 11164 -5819
rect 11112 -5926 11120 -5892
rect 11154 -5926 11164 -5892
rect 11112 -5949 11164 -5926
rect 11264 -5865 11314 -5819
rect 11264 -5892 11336 -5865
rect 11264 -5926 11280 -5892
rect 11314 -5926 11336 -5892
rect 11264 -5949 11336 -5926
rect 11366 -5892 11420 -5865
rect 11366 -5926 11377 -5892
rect 11411 -5926 11420 -5892
rect 11366 -5949 11420 -5926
rect 11658 -5877 11710 -5839
rect 11658 -5911 11666 -5877
rect 11700 -5911 11710 -5877
rect 11658 -5949 11710 -5911
rect 11920 -5877 11972 -5839
rect 11920 -5911 11930 -5877
rect 11964 -5911 11972 -5877
rect 11920 -5949 11972 -5911
rect 13682 -5903 13735 -5865
rect 13682 -5937 13690 -5903
rect 13724 -5937 13735 -5903
rect 13682 -5949 13735 -5937
rect 13765 -5890 13821 -5865
rect 13765 -5924 13776 -5890
rect 13810 -5924 13821 -5890
rect 13765 -5949 13821 -5924
rect 13851 -5890 13907 -5865
rect 13851 -5924 13862 -5890
rect 13896 -5924 13907 -5890
rect 13851 -5949 13907 -5924
rect 13937 -5890 13993 -5865
rect 13937 -5924 13948 -5890
rect 13982 -5924 13993 -5890
rect 13937 -5949 13993 -5924
rect 14023 -5890 14079 -5865
rect 14023 -5924 14034 -5890
rect 14068 -5924 14079 -5890
rect 14023 -5949 14079 -5924
rect 14109 -5890 14165 -5865
rect 14109 -5924 14120 -5890
rect 14154 -5924 14165 -5890
rect 14109 -5949 14165 -5924
rect 14195 -5899 14251 -5865
rect 14195 -5933 14206 -5899
rect 14240 -5933 14251 -5899
rect 14195 -5949 14251 -5933
rect 14281 -5890 14337 -5865
rect 14281 -5924 14292 -5890
rect 14326 -5924 14337 -5890
rect 14281 -5949 14337 -5924
rect 14367 -5899 14423 -5865
rect 14367 -5933 14378 -5899
rect 14412 -5933 14423 -5899
rect 14367 -5949 14423 -5933
rect 14453 -5890 14509 -5865
rect 14453 -5924 14464 -5890
rect 14498 -5924 14509 -5890
rect 14453 -5949 14509 -5924
rect 14539 -5899 14595 -5865
rect 14539 -5933 14550 -5899
rect 14584 -5933 14595 -5899
rect 14539 -5949 14595 -5933
rect 14625 -5890 14681 -5865
rect 14625 -5924 14636 -5890
rect 14670 -5924 14681 -5890
rect 14625 -5949 14681 -5924
rect 14711 -5899 14766 -5865
rect 14711 -5933 14722 -5899
rect 14756 -5933 14766 -5899
rect 14711 -5949 14766 -5933
rect 14796 -5890 14852 -5865
rect 14796 -5924 14807 -5890
rect 14841 -5924 14852 -5890
rect 14796 -5949 14852 -5924
rect 14882 -5899 14938 -5865
rect 14882 -5933 14893 -5899
rect 14927 -5933 14938 -5899
rect 14882 -5949 14938 -5933
rect 14968 -5890 15024 -5865
rect 14968 -5924 14979 -5890
rect 15013 -5924 15024 -5890
rect 14968 -5949 15024 -5924
rect 15054 -5899 15110 -5865
rect 15054 -5933 15065 -5899
rect 15099 -5933 15110 -5899
rect 15054 -5949 15110 -5933
rect 15140 -5890 15196 -5865
rect 15140 -5924 15151 -5890
rect 15185 -5924 15196 -5890
rect 15140 -5949 15196 -5924
rect 15226 -5899 15282 -5865
rect 15226 -5933 15237 -5899
rect 15271 -5933 15282 -5899
rect 15226 -5949 15282 -5933
rect 15312 -5890 15368 -5865
rect 15312 -5924 15323 -5890
rect 15357 -5924 15368 -5890
rect 15312 -5949 15368 -5924
rect 15398 -5899 15451 -5865
rect 15398 -5933 15409 -5899
rect 15443 -5933 15451 -5899
rect 15614 -5884 15666 -5839
rect 15614 -5918 15622 -5884
rect 15656 -5918 15666 -5884
rect 15398 -5949 15451 -5933
rect 15614 -5949 15666 -5918
rect 16612 -5884 16664 -5839
rect 16612 -5918 16622 -5884
rect 16656 -5918 16664 -5884
rect 16612 -5949 16664 -5918
rect -2970 -6074 -2918 -6043
rect -2970 -6108 -2962 -6074
rect -2928 -6108 -2918 -6074
rect -2970 -6153 -2918 -6108
rect -2340 -6074 -2288 -6043
rect -2340 -6108 -2330 -6074
rect -2296 -6108 -2288 -6074
rect -2340 -6153 -2288 -6108
rect -1406 -6081 -1354 -6043
rect -1406 -6115 -1398 -6081
rect -1364 -6115 -1354 -6081
rect -1406 -6153 -1354 -6115
rect -1144 -6081 -1092 -6043
rect -942 -6055 -890 -6043
rect -1144 -6115 -1134 -6081
rect -1100 -6115 -1092 -6081
rect -1144 -6153 -1092 -6115
rect -942 -6089 -934 -6055
rect -900 -6089 -890 -6055
rect -942 -6123 -890 -6089
rect -942 -6157 -934 -6123
rect -900 -6157 -890 -6123
rect -942 -6173 -890 -6157
rect -860 -6173 -806 -6043
rect -776 -6055 -724 -6043
rect -776 -6089 -766 -6055
rect -732 -6089 -724 -6055
rect -776 -6123 -724 -6089
rect -776 -6157 -766 -6123
rect -732 -6157 -724 -6123
rect -776 -6173 -724 -6157
rect -578 -6081 -526 -6043
rect -578 -6115 -570 -6081
rect -536 -6115 -526 -6081
rect -578 -6153 -526 -6115
rect -316 -6081 -264 -6043
rect -37 -6057 29 -6043
rect -316 -6115 -306 -6081
rect -272 -6115 -264 -6081
rect -316 -6153 -264 -6115
rect -37 -6091 -16 -6057
rect 18 -6091 29 -6057
rect -37 -6127 29 -6091
rect 59 -6068 115 -6043
rect 59 -6102 70 -6068
rect 104 -6102 115 -6068
rect 59 -6127 115 -6102
rect 145 -6057 201 -6043
rect 145 -6091 156 -6057
rect 190 -6091 201 -6057
rect 145 -6127 201 -6091
rect 231 -6068 287 -6043
rect 231 -6102 242 -6068
rect 276 -6102 287 -6068
rect 231 -6127 287 -6102
rect 317 -6057 396 -6043
rect 317 -6091 328 -6057
rect 362 -6091 396 -6057
rect 317 -6127 396 -6091
rect 618 -6081 670 -6043
rect 618 -6115 626 -6081
rect 660 -6115 670 -6081
rect 618 -6153 670 -6115
rect 880 -6081 932 -6043
rect 880 -6115 890 -6081
rect 924 -6115 932 -6081
rect 880 -6153 932 -6115
rect 1161 -6066 1213 -6043
rect 1161 -6100 1169 -6066
rect 1203 -6100 1213 -6066
rect 1161 -6127 1213 -6100
rect 1243 -6064 1300 -6043
rect 1243 -6098 1253 -6064
rect 1287 -6098 1300 -6064
rect 1243 -6127 1300 -6098
rect 1446 -6081 1498 -6043
rect 1446 -6115 1454 -6081
rect 1488 -6115 1498 -6081
rect 1446 -6153 1498 -6115
rect 1708 -6081 1760 -6043
rect 1708 -6115 1718 -6081
rect 1752 -6115 1760 -6081
rect 1708 -6153 1760 -6115
rect 1906 -6081 1958 -6043
rect 1906 -6115 1914 -6081
rect 1948 -6115 1958 -6081
rect 1906 -6153 1958 -6115
rect 2168 -6081 2220 -6043
rect 2168 -6115 2178 -6081
rect 2212 -6115 2220 -6081
rect 2168 -6153 2220 -6115
rect 2366 -6066 2420 -6043
rect 2366 -6100 2375 -6066
rect 2409 -6100 2420 -6066
rect 2366 -6127 2420 -6100
rect 2450 -6066 2522 -6043
rect 2450 -6100 2472 -6066
rect 2506 -6100 2522 -6066
rect 2450 -6127 2522 -6100
rect 2472 -6173 2522 -6127
rect 2622 -6066 2674 -6043
rect 2622 -6100 2632 -6066
rect 2666 -6100 2674 -6066
rect 2622 -6173 2674 -6100
rect 2729 -6066 2782 -6043
rect 2729 -6100 2737 -6066
rect 2771 -6100 2782 -6066
rect 2729 -6173 2782 -6100
rect 2882 -6066 2947 -6043
rect 2882 -6100 2893 -6066
rect 2927 -6100 2947 -6066
rect 2882 -6127 2947 -6100
rect 2977 -6066 3048 -6043
rect 2977 -6100 2991 -6066
rect 3025 -6100 3048 -6066
rect 2977 -6127 3048 -6100
rect 2882 -6173 2932 -6127
rect 3194 -6081 3246 -6043
rect 3194 -6115 3202 -6081
rect 3236 -6115 3246 -6081
rect 3194 -6153 3246 -6115
rect 3456 -6081 3508 -6043
rect 3456 -6115 3466 -6081
rect 3500 -6115 3508 -6081
rect 3456 -6153 3508 -6115
rect 4390 -6074 4442 -6043
rect 4390 -6108 4398 -6074
rect 4432 -6108 4442 -6074
rect 4390 -6153 4442 -6108
rect 5388 -6074 5440 -6043
rect 5388 -6108 5398 -6074
rect 5432 -6108 5440 -6074
rect 5388 -6153 5440 -6108
rect 6414 -6081 6466 -6043
rect 6414 -6115 6422 -6081
rect 6456 -6115 6466 -6081
rect 6414 -6153 6466 -6115
rect 6676 -6081 6728 -6043
rect 6676 -6115 6686 -6081
rect 6720 -6115 6728 -6081
rect 6676 -6153 6728 -6115
rect 6874 -6066 6928 -6043
rect 6874 -6100 6883 -6066
rect 6917 -6100 6928 -6066
rect 6874 -6127 6928 -6100
rect 6958 -6066 7030 -6043
rect 6958 -6100 6980 -6066
rect 7014 -6100 7030 -6066
rect 6958 -6127 7030 -6100
rect 6980 -6173 7030 -6127
rect 7130 -6066 7182 -6043
rect 7130 -6100 7140 -6066
rect 7174 -6100 7182 -6066
rect 7130 -6173 7182 -6100
rect 7237 -6066 7290 -6043
rect 7237 -6100 7245 -6066
rect 7279 -6100 7290 -6066
rect 7237 -6173 7290 -6100
rect 7390 -6066 7455 -6043
rect 7390 -6100 7401 -6066
rect 7435 -6100 7455 -6066
rect 7390 -6127 7455 -6100
rect 7485 -6066 7556 -6043
rect 7485 -6100 7499 -6066
rect 7533 -6100 7556 -6066
rect 7485 -6127 7556 -6100
rect 7390 -6173 7440 -6127
rect 7702 -6081 7754 -6043
rect 7702 -6115 7710 -6081
rect 7744 -6115 7754 -6081
rect 7702 -6153 7754 -6115
rect 7964 -6081 8016 -6043
rect 7964 -6115 7974 -6081
rect 8008 -6115 8016 -6081
rect 7964 -6153 8016 -6115
rect 8162 -6066 8216 -6043
rect 8162 -6100 8171 -6066
rect 8205 -6100 8216 -6066
rect 8162 -6127 8216 -6100
rect 8246 -6066 8318 -6043
rect 8246 -6100 8268 -6066
rect 8302 -6100 8318 -6066
rect 8246 -6127 8318 -6100
rect 8268 -6173 8318 -6127
rect 8418 -6066 8470 -6043
rect 8418 -6100 8428 -6066
rect 8462 -6100 8470 -6066
rect 8418 -6173 8470 -6100
rect 8525 -6066 8578 -6043
rect 8525 -6100 8533 -6066
rect 8567 -6100 8578 -6066
rect 8525 -6173 8578 -6100
rect 8678 -6066 8743 -6043
rect 8678 -6100 8689 -6066
rect 8723 -6100 8743 -6066
rect 8678 -6127 8743 -6100
rect 8773 -6066 8844 -6043
rect 8773 -6100 8787 -6066
rect 8821 -6100 8844 -6066
rect 8773 -6127 8844 -6100
rect 8678 -6173 8728 -6127
rect 8990 -6081 9042 -6043
rect 8990 -6115 8998 -6081
rect 9032 -6115 9042 -6081
rect 8990 -6153 9042 -6115
rect 9252 -6081 9304 -6043
rect 9252 -6115 9262 -6081
rect 9296 -6115 9304 -6081
rect 9252 -6153 9304 -6115
rect 9450 -6066 9504 -6043
rect 9450 -6100 9459 -6066
rect 9493 -6100 9504 -6066
rect 9450 -6127 9504 -6100
rect 9534 -6066 9606 -6043
rect 9534 -6100 9556 -6066
rect 9590 -6100 9606 -6066
rect 9534 -6127 9606 -6100
rect 9556 -6173 9606 -6127
rect 9706 -6066 9758 -6043
rect 9706 -6100 9716 -6066
rect 9750 -6100 9758 -6066
rect 9706 -6173 9758 -6100
rect 9813 -6066 9866 -6043
rect 9813 -6100 9821 -6066
rect 9855 -6100 9866 -6066
rect 9813 -6173 9866 -6100
rect 9966 -6066 10031 -6043
rect 9966 -6100 9977 -6066
rect 10011 -6100 10031 -6066
rect 9966 -6127 10031 -6100
rect 10061 -6066 10132 -6043
rect 10061 -6100 10075 -6066
rect 10109 -6100 10132 -6066
rect 10061 -6127 10132 -6100
rect 9966 -6173 10016 -6127
rect 10278 -6081 10330 -6043
rect 10278 -6115 10286 -6081
rect 10320 -6115 10330 -6081
rect 10278 -6153 10330 -6115
rect 10540 -6081 10592 -6043
rect 10738 -6055 10790 -6043
rect 10540 -6115 10550 -6081
rect 10584 -6115 10592 -6081
rect 10540 -6153 10592 -6115
rect 10738 -6089 10746 -6055
rect 10780 -6089 10790 -6055
rect 10738 -6123 10790 -6089
rect 10738 -6157 10746 -6123
rect 10780 -6157 10790 -6123
rect 10738 -6173 10790 -6157
rect 10820 -6055 10874 -6043
rect 10820 -6089 10830 -6055
rect 10864 -6089 10874 -6055
rect 10820 -6173 10874 -6089
rect 10904 -6055 10958 -6043
rect 10904 -6089 10914 -6055
rect 10948 -6089 10958 -6055
rect 10904 -6123 10958 -6089
rect 10904 -6157 10914 -6123
rect 10948 -6157 10958 -6123
rect 10904 -6173 10958 -6157
rect 10988 -6055 11042 -6043
rect 10988 -6089 10998 -6055
rect 11032 -6089 11042 -6055
rect 10988 -6173 11042 -6089
rect 11072 -6055 11126 -6043
rect 11072 -6089 11082 -6055
rect 11116 -6089 11126 -6055
rect 11072 -6123 11126 -6089
rect 11072 -6157 11082 -6123
rect 11116 -6157 11126 -6123
rect 11072 -6173 11126 -6157
rect 11156 -6123 11210 -6043
rect 11156 -6157 11166 -6123
rect 11200 -6157 11210 -6123
rect 11156 -6173 11210 -6157
rect 11240 -6055 11294 -6043
rect 11240 -6089 11250 -6055
rect 11284 -6089 11294 -6055
rect 11240 -6173 11294 -6089
rect 11324 -6123 11378 -6043
rect 11324 -6157 11334 -6123
rect 11368 -6157 11378 -6123
rect 11324 -6173 11378 -6157
rect 11408 -6055 11460 -6043
rect 11408 -6089 11418 -6055
rect 11452 -6089 11460 -6055
rect 11408 -6123 11460 -6089
rect 11408 -6157 11418 -6123
rect 11452 -6157 11460 -6123
rect 11408 -6173 11460 -6157
rect 11658 -6081 11710 -6043
rect 11658 -6115 11666 -6081
rect 11700 -6115 11710 -6081
rect 11658 -6153 11710 -6115
rect 11920 -6081 11972 -6043
rect 11920 -6115 11930 -6081
rect 11964 -6115 11972 -6081
rect 11920 -6153 11972 -6115
rect 13590 -6074 13642 -6043
rect 13590 -6108 13598 -6074
rect 13632 -6108 13642 -6074
rect 13590 -6153 13642 -6108
rect 14588 -6074 14640 -6043
rect 14588 -6108 14598 -6074
rect 14632 -6108 14640 -6074
rect 14588 -6153 14640 -6108
rect 14786 -6074 14838 -6043
rect 14786 -6108 14794 -6074
rect 14828 -6108 14838 -6074
rect 14786 -6153 14838 -6108
rect 15784 -6074 15836 -6043
rect 15784 -6108 15794 -6074
rect 15828 -6108 15836 -6074
rect 15784 -6153 15836 -6108
rect 15982 -6074 16034 -6043
rect 15982 -6108 15990 -6074
rect 16024 -6108 16034 -6074
rect 15982 -6153 16034 -6108
rect 16612 -6074 16664 -6043
rect 16612 -6108 16622 -6074
rect 16656 -6108 16664 -6074
rect 16612 -6153 16664 -6108
rect -2970 -6970 -2918 -6927
rect -2970 -7004 -2962 -6970
rect -2928 -7004 -2918 -6970
rect -2970 -7037 -2918 -7004
rect -2800 -6970 -2748 -6927
rect -2800 -7004 -2790 -6970
rect -2756 -7004 -2748 -6970
rect -2800 -7037 -2748 -7004
rect -2602 -6965 -2550 -6953
rect -2602 -6999 -2594 -6965
rect -2560 -6999 -2550 -6965
rect -2602 -7037 -2550 -6999
rect -2520 -6991 -2466 -6953
rect -2520 -7025 -2510 -6991
rect -2476 -7025 -2466 -6991
rect -2520 -7037 -2466 -7025
rect -2436 -6965 -2384 -6953
rect -2436 -6999 -2426 -6965
rect -2392 -6999 -2384 -6965
rect -2436 -7037 -2384 -6999
rect -2330 -6991 -2278 -6953
rect -2330 -7025 -2322 -6991
rect -2288 -7025 -2278 -6991
rect -2330 -7037 -2278 -7025
rect -2248 -6965 -2198 -6953
rect -1899 -6953 -1849 -6909
rect -2018 -6965 -1968 -6953
rect -2248 -6977 -2166 -6965
rect -2248 -7011 -2237 -6977
rect -2203 -7011 -2166 -6977
rect -2248 -7037 -2166 -7011
rect -2136 -6977 -2067 -6965
rect -2136 -7011 -2126 -6977
rect -2092 -7011 -2067 -6977
rect -2136 -7037 -2067 -7011
rect -2037 -7037 -1968 -6965
rect -1938 -6983 -1849 -6953
rect -1938 -7017 -1927 -6983
rect -1893 -7017 -1849 -6983
rect -1938 -7037 -1849 -7017
rect -1819 -6965 -1769 -6909
rect -1409 -6922 -1357 -6907
rect -1597 -6965 -1547 -6953
rect -1819 -6977 -1748 -6965
rect -1819 -7011 -1808 -6977
rect -1774 -7011 -1748 -6977
rect -1819 -7037 -1748 -7011
rect -1718 -6977 -1642 -6965
rect -1718 -7011 -1705 -6977
rect -1671 -7011 -1642 -6977
rect -1718 -7037 -1642 -7011
rect -1612 -7037 -1547 -6965
rect -1517 -6977 -1465 -6953
rect -1517 -7011 -1507 -6977
rect -1473 -7011 -1465 -6977
rect -1517 -7037 -1465 -7011
rect -1409 -6956 -1401 -6922
rect -1367 -6956 -1357 -6922
rect -1409 -6990 -1357 -6956
rect -1409 -7024 -1401 -6990
rect -1367 -7024 -1357 -6990
rect -1409 -7037 -1357 -7024
rect -1327 -6961 -1273 -6907
rect -1327 -6995 -1317 -6961
rect -1283 -6995 -1273 -6961
rect -1327 -7037 -1273 -6995
rect -1243 -6920 -1191 -6907
rect -1243 -6954 -1233 -6920
rect -1199 -6954 -1191 -6920
rect -1040 -6953 -990 -6907
rect -1243 -6988 -1191 -6954
rect -1243 -7022 -1233 -6988
rect -1199 -7022 -1191 -6988
rect -1243 -7037 -1191 -7022
rect -1137 -6965 -1085 -6953
rect -1137 -6999 -1129 -6965
rect -1095 -6999 -1085 -6965
rect -1137 -7037 -1085 -6999
rect -1055 -6991 -990 -6953
rect -1055 -7025 -1034 -6991
rect -1000 -7025 -990 -6991
rect -1055 -7037 -990 -7025
rect -960 -6953 -908 -6907
rect -960 -6987 -950 -6953
rect -916 -6987 -908 -6953
rect -960 -7037 -908 -6987
rect -854 -6972 -802 -6927
rect -854 -7006 -846 -6972
rect -812 -7006 -802 -6972
rect -854 -7037 -802 -7006
rect -224 -6972 -172 -6927
rect -224 -7006 -214 -6972
rect -180 -7006 -172 -6972
rect -224 -7037 -172 -7006
rect -26 -6972 26 -6927
rect -26 -7006 -18 -6972
rect 16 -7006 26 -6972
rect -26 -7037 26 -7006
rect 604 -6972 656 -6927
rect 604 -7006 614 -6972
rect 648 -7006 656 -6972
rect 604 -7037 656 -7006
rect 710 -6972 762 -6927
rect 710 -7006 718 -6972
rect 752 -7006 762 -6972
rect 710 -7037 762 -7006
rect 1340 -6972 1392 -6927
rect 1340 -7006 1350 -6972
rect 1384 -7006 1392 -6972
rect 1340 -7037 1392 -7006
rect 1538 -6972 1590 -6927
rect 1538 -7006 1546 -6972
rect 1580 -7006 1590 -6972
rect 1538 -7037 1590 -7006
rect 2168 -6972 2220 -6927
rect 2168 -7006 2178 -6972
rect 2212 -7006 2220 -6972
rect 2168 -7037 2220 -7006
rect 2274 -6972 2326 -6927
rect 2274 -7006 2282 -6972
rect 2316 -7006 2326 -6972
rect 2274 -7037 2326 -7006
rect 2904 -6972 2956 -6927
rect 2904 -7006 2914 -6972
rect 2948 -7006 2956 -6972
rect 2904 -7037 2956 -7006
rect 3102 -6972 3154 -6927
rect 3102 -7006 3110 -6972
rect 3144 -7006 3154 -6972
rect 3102 -7037 3154 -7006
rect 3732 -6972 3784 -6927
rect 3732 -7006 3742 -6972
rect 3776 -7006 3784 -6972
rect 3732 -7037 3784 -7006
rect 3838 -6972 3890 -6927
rect 3838 -7006 3846 -6972
rect 3880 -7006 3890 -6972
rect 3838 -7037 3890 -7006
rect 4468 -6972 4520 -6927
rect 4468 -7006 4478 -6972
rect 4512 -7006 4520 -6972
rect 4468 -7037 4520 -7006
rect 4666 -6972 4718 -6927
rect 4666 -7006 4674 -6972
rect 4708 -7006 4718 -6972
rect 4666 -7037 4718 -7006
rect 5296 -6972 5348 -6927
rect 5296 -7006 5306 -6972
rect 5340 -7006 5348 -6972
rect 5296 -7037 5348 -7006
rect 5402 -6972 5454 -6927
rect 5402 -7006 5410 -6972
rect 5444 -7006 5454 -6972
rect 5402 -7037 5454 -7006
rect 6032 -6972 6084 -6927
rect 6032 -7006 6042 -6972
rect 6076 -7006 6084 -6972
rect 6032 -7037 6084 -7006
rect 6230 -6972 6282 -6927
rect 6230 -7006 6238 -6972
rect 6272 -7006 6282 -6972
rect 6230 -7037 6282 -7006
rect 6860 -6972 6912 -6927
rect 6860 -7006 6870 -6972
rect 6904 -7006 6912 -6972
rect 6860 -7037 6912 -7006
rect 6966 -6972 7018 -6927
rect 6966 -7006 6974 -6972
rect 7008 -7006 7018 -6972
rect 6966 -7037 7018 -7006
rect 7596 -6972 7648 -6927
rect 7596 -7006 7606 -6972
rect 7640 -7006 7648 -6972
rect 7596 -7037 7648 -7006
rect 7794 -6972 7846 -6927
rect 7794 -7006 7802 -6972
rect 7836 -7006 7846 -6972
rect 7794 -7037 7846 -7006
rect 8424 -6972 8476 -6927
rect 8424 -7006 8434 -6972
rect 8468 -7006 8476 -6972
rect 8424 -7037 8476 -7006
rect 8530 -6972 8582 -6927
rect 8530 -7006 8538 -6972
rect 8572 -7006 8582 -6972
rect 8530 -7037 8582 -7006
rect 9160 -6972 9212 -6927
rect 9160 -7006 9170 -6972
rect 9204 -7006 9212 -6972
rect 9160 -7037 9212 -7006
rect 15982 -6972 16034 -6927
rect 15982 -7006 15990 -6972
rect 16024 -7006 16034 -6972
rect 15982 -7037 16034 -7006
rect 16612 -6972 16664 -6927
rect 16612 -7006 16622 -6972
rect 16656 -7006 16664 -6972
rect 16612 -7037 16664 -7006
rect -2970 -7162 -2918 -7131
rect -2970 -7196 -2962 -7162
rect -2928 -7196 -2918 -7162
rect -2970 -7241 -2918 -7196
rect -2340 -7162 -2288 -7131
rect -2340 -7196 -2330 -7162
rect -2296 -7196 -2288 -7162
rect -2340 -7241 -2288 -7196
rect -1590 -7162 -1538 -7131
rect -1590 -7196 -1582 -7162
rect -1548 -7196 -1538 -7162
rect -1590 -7241 -1538 -7196
rect -960 -7162 -908 -7131
rect -960 -7196 -950 -7162
rect -916 -7196 -908 -7162
rect -960 -7241 -908 -7196
rect -854 -7162 -802 -7131
rect -854 -7196 -846 -7162
rect -812 -7196 -802 -7162
rect -854 -7241 -802 -7196
rect -224 -7162 -172 -7131
rect -224 -7196 -214 -7162
rect -180 -7196 -172 -7162
rect -224 -7241 -172 -7196
rect -26 -7162 26 -7131
rect -26 -7196 -18 -7162
rect 16 -7196 26 -7162
rect -26 -7241 26 -7196
rect 604 -7162 656 -7131
rect 604 -7196 614 -7162
rect 648 -7196 656 -7162
rect 604 -7241 656 -7196
rect 710 -7162 762 -7131
rect 710 -7196 718 -7162
rect 752 -7196 762 -7162
rect 710 -7241 762 -7196
rect 1340 -7162 1392 -7131
rect 1340 -7196 1350 -7162
rect 1384 -7196 1392 -7162
rect 1340 -7241 1392 -7196
rect 1538 -7162 1590 -7131
rect 1538 -7196 1546 -7162
rect 1580 -7196 1590 -7162
rect 1538 -7241 1590 -7196
rect 2168 -7162 2220 -7131
rect 2168 -7196 2178 -7162
rect 2212 -7196 2220 -7162
rect 2168 -7241 2220 -7196
rect 2274 -7169 2326 -7131
rect 2274 -7203 2282 -7169
rect 2316 -7203 2326 -7169
rect 2274 -7241 2326 -7203
rect 2536 -7169 2588 -7131
rect 2536 -7203 2546 -7169
rect 2580 -7203 2588 -7169
rect 2536 -7241 2588 -7203
rect 2918 -7152 2975 -7131
rect 2918 -7186 2931 -7152
rect 2965 -7186 2975 -7152
rect 2918 -7215 2975 -7186
rect 3005 -7154 3057 -7131
rect 3005 -7188 3015 -7154
rect 3049 -7188 3057 -7154
rect 3005 -7215 3057 -7188
rect 3286 -7169 3338 -7131
rect 3286 -7203 3294 -7169
rect 3328 -7203 3338 -7169
rect 3286 -7241 3338 -7203
rect 3548 -7169 3600 -7131
rect 3750 -7143 3802 -7131
rect 3548 -7203 3558 -7169
rect 3592 -7203 3600 -7169
rect 3548 -7241 3600 -7203
rect 3750 -7177 3758 -7143
rect 3792 -7177 3802 -7143
rect 3750 -7211 3802 -7177
rect 3750 -7245 3758 -7211
rect 3792 -7245 3802 -7211
rect 3750 -7261 3802 -7245
rect 3832 -7261 3886 -7131
rect 3916 -7143 3968 -7131
rect 3916 -7177 3926 -7143
rect 3960 -7177 3968 -7143
rect 3916 -7211 3968 -7177
rect 3916 -7245 3926 -7211
rect 3960 -7245 3968 -7211
rect 3916 -7261 3968 -7245
rect 4114 -7169 4166 -7131
rect 4114 -7203 4122 -7169
rect 4156 -7203 4166 -7169
rect 4114 -7241 4166 -7203
rect 4376 -7169 4428 -7131
rect 4376 -7203 4386 -7169
rect 4420 -7203 4428 -7169
rect 4376 -7241 4428 -7203
rect 4574 -7162 4626 -7131
rect 4574 -7196 4582 -7162
rect 4616 -7196 4626 -7162
rect 4574 -7261 4626 -7196
rect 4656 -7143 4735 -7131
rect 4656 -7177 4666 -7143
rect 4700 -7177 4735 -7143
rect 4656 -7215 4735 -7177
rect 4765 -7215 4831 -7131
rect 4861 -7158 4956 -7131
rect 4861 -7192 4873 -7158
rect 4907 -7192 4956 -7158
rect 4861 -7215 4956 -7192
rect 4986 -7215 5052 -7131
rect 5082 -7158 5220 -7131
rect 5082 -7192 5108 -7158
rect 5142 -7192 5176 -7158
rect 5210 -7192 5220 -7158
rect 5082 -7215 5220 -7192
rect 5250 -7158 5302 -7131
rect 5250 -7192 5260 -7158
rect 5294 -7192 5302 -7158
rect 5250 -7215 5302 -7192
rect 4656 -7261 4708 -7215
rect 5494 -7169 5546 -7131
rect 5494 -7203 5502 -7169
rect 5536 -7203 5546 -7169
rect 5494 -7241 5546 -7203
rect 5756 -7169 5808 -7131
rect 5756 -7203 5766 -7169
rect 5800 -7203 5808 -7169
rect 5756 -7241 5808 -7203
rect 5954 -7181 6006 -7131
rect 5954 -7215 5962 -7181
rect 5996 -7215 6006 -7181
rect 5954 -7261 6006 -7215
rect 6036 -7143 6101 -7131
rect 6036 -7177 6046 -7143
rect 6080 -7177 6101 -7143
rect 6036 -7215 6101 -7177
rect 6131 -7169 6183 -7131
rect 6131 -7203 6141 -7169
rect 6175 -7203 6183 -7169
rect 6131 -7215 6183 -7203
rect 6237 -7146 6289 -7131
rect 6237 -7180 6245 -7146
rect 6279 -7180 6289 -7146
rect 6237 -7214 6289 -7180
rect 6036 -7261 6086 -7215
rect 6237 -7248 6245 -7214
rect 6279 -7248 6289 -7214
rect 6237 -7261 6289 -7248
rect 6319 -7173 6373 -7131
rect 6319 -7207 6329 -7173
rect 6363 -7207 6373 -7173
rect 6319 -7261 6373 -7207
rect 6403 -7144 6455 -7131
rect 6403 -7178 6413 -7144
rect 6447 -7178 6455 -7144
rect 6403 -7212 6455 -7178
rect 6403 -7246 6413 -7212
rect 6447 -7246 6455 -7212
rect 6511 -7157 6563 -7131
rect 6511 -7191 6519 -7157
rect 6553 -7191 6563 -7157
rect 6511 -7215 6563 -7191
rect 6593 -7203 6658 -7131
rect 6688 -7157 6764 -7131
rect 6688 -7191 6717 -7157
rect 6751 -7191 6764 -7157
rect 6688 -7203 6764 -7191
rect 6794 -7157 6865 -7131
rect 6794 -7191 6820 -7157
rect 6854 -7191 6865 -7157
rect 6794 -7203 6865 -7191
rect 6593 -7215 6643 -7203
rect 6403 -7261 6455 -7246
rect 6815 -7259 6865 -7203
rect 6895 -7151 6984 -7131
rect 6895 -7185 6939 -7151
rect 6973 -7185 6984 -7151
rect 6895 -7215 6984 -7185
rect 7014 -7203 7083 -7131
rect 7113 -7157 7182 -7131
rect 7113 -7191 7138 -7157
rect 7172 -7191 7182 -7157
rect 7113 -7203 7182 -7191
rect 7212 -7157 7294 -7131
rect 7212 -7191 7249 -7157
rect 7283 -7191 7294 -7157
rect 7212 -7203 7294 -7191
rect 7014 -7215 7064 -7203
rect 6895 -7259 6945 -7215
rect 7244 -7215 7294 -7203
rect 7324 -7143 7376 -7131
rect 7324 -7177 7334 -7143
rect 7368 -7177 7376 -7143
rect 7324 -7215 7376 -7177
rect 7430 -7169 7482 -7131
rect 7430 -7203 7438 -7169
rect 7472 -7203 7482 -7169
rect 7430 -7215 7482 -7203
rect 7512 -7143 7566 -7131
rect 7512 -7177 7522 -7143
rect 7556 -7177 7566 -7143
rect 7512 -7215 7566 -7177
rect 7596 -7169 7648 -7131
rect 7596 -7203 7606 -7169
rect 7640 -7203 7648 -7169
rect 7596 -7215 7648 -7203
rect 7794 -7162 7846 -7131
rect 7794 -7196 7802 -7162
rect 7836 -7196 7846 -7162
rect 7794 -7241 7846 -7196
rect 8424 -7162 8476 -7131
rect 8424 -7196 8434 -7162
rect 8468 -7196 8476 -7162
rect 8424 -7241 8476 -7196
rect 8530 -7162 8582 -7131
rect 8530 -7196 8538 -7162
rect 8572 -7196 8582 -7162
rect 8530 -7241 8582 -7196
rect 9160 -7162 9212 -7131
rect 9160 -7196 9170 -7162
rect 9204 -7196 9212 -7162
rect 9160 -7241 9212 -7196
rect 15982 -7162 16034 -7131
rect 15982 -7196 15990 -7162
rect 16024 -7196 16034 -7162
rect 15982 -7241 16034 -7196
rect 16612 -7162 16664 -7131
rect 16612 -7196 16622 -7162
rect 16656 -7196 16664 -7162
rect 16612 -7241 16664 -7196
rect -2970 -8060 -2918 -8015
rect -2970 -8094 -2962 -8060
rect -2928 -8094 -2918 -8060
rect -2970 -8125 -2918 -8094
rect -2340 -8060 -2288 -8015
rect -2340 -8094 -2330 -8060
rect -2296 -8094 -2288 -8060
rect -2340 -8125 -2288 -8094
rect -1406 -8053 -1354 -8015
rect -1406 -8087 -1398 -8053
rect -1364 -8087 -1354 -8053
rect -1406 -8125 -1354 -8087
rect -1144 -8053 -1092 -8015
rect -1144 -8087 -1134 -8053
rect -1100 -8087 -1092 -8053
rect -1144 -8125 -1092 -8087
rect -942 -8011 -890 -7995
rect -942 -8045 -934 -8011
rect -900 -8045 -890 -8011
rect -942 -8079 -890 -8045
rect -942 -8113 -934 -8079
rect -900 -8113 -890 -8079
rect -942 -8125 -890 -8113
rect -860 -8125 -806 -7995
rect -776 -8011 -724 -7995
rect -776 -8045 -766 -8011
rect -732 -8045 -724 -8011
rect -776 -8079 -724 -8045
rect -776 -8113 -766 -8079
rect -732 -8113 -724 -8079
rect -578 -8053 -526 -8015
rect -578 -8087 -570 -8053
rect -536 -8087 -526 -8053
rect -776 -8125 -724 -8113
rect -578 -8125 -526 -8087
rect -316 -8053 -264 -8015
rect -316 -8087 -306 -8053
rect -272 -8087 -264 -8053
rect -316 -8125 -264 -8087
rect -37 -8077 29 -8041
rect -37 -8111 -16 -8077
rect 18 -8111 29 -8077
rect -37 -8125 29 -8111
rect 59 -8066 115 -8041
rect 59 -8100 70 -8066
rect 104 -8100 115 -8066
rect 59 -8125 115 -8100
rect 145 -8077 201 -8041
rect 145 -8111 156 -8077
rect 190 -8111 201 -8077
rect 145 -8125 201 -8111
rect 231 -8066 287 -8041
rect 231 -8100 242 -8066
rect 276 -8100 287 -8066
rect 231 -8125 287 -8100
rect 317 -8077 396 -8041
rect 317 -8111 328 -8077
rect 362 -8111 396 -8077
rect 618 -8053 670 -8015
rect 618 -8087 626 -8053
rect 660 -8087 670 -8053
rect 317 -8125 396 -8111
rect 618 -8125 670 -8087
rect 880 -8053 932 -8015
rect 880 -8087 890 -8053
rect 924 -8087 932 -8053
rect 880 -8125 932 -8087
rect 1161 -8068 1213 -8041
rect 1161 -8102 1169 -8068
rect 1203 -8102 1213 -8068
rect 1161 -8125 1213 -8102
rect 1243 -8070 1300 -8041
rect 1243 -8104 1253 -8070
rect 1287 -8104 1300 -8070
rect 1243 -8125 1300 -8104
rect 1446 -8053 1498 -8015
rect 1446 -8087 1454 -8053
rect 1488 -8087 1498 -8053
rect 1446 -8125 1498 -8087
rect 1708 -8053 1760 -8015
rect 1708 -8087 1718 -8053
rect 1752 -8087 1760 -8053
rect 1708 -8125 1760 -8087
rect 1906 -8053 1958 -8015
rect 1906 -8087 1914 -8053
rect 1948 -8087 1958 -8053
rect 1906 -8125 1958 -8087
rect 2168 -8053 2220 -8015
rect 2168 -8087 2178 -8053
rect 2212 -8087 2220 -8053
rect 2168 -8125 2220 -8087
rect 2472 -8041 2522 -7995
rect 2366 -8068 2420 -8041
rect 2366 -8102 2375 -8068
rect 2409 -8102 2420 -8068
rect 2366 -8125 2420 -8102
rect 2450 -8068 2522 -8041
rect 2450 -8102 2472 -8068
rect 2506 -8102 2522 -8068
rect 2450 -8125 2522 -8102
rect 2622 -8068 2674 -7995
rect 2622 -8102 2632 -8068
rect 2666 -8102 2674 -8068
rect 2622 -8125 2674 -8102
rect 2729 -8068 2782 -7995
rect 2729 -8102 2737 -8068
rect 2771 -8102 2782 -8068
rect 2729 -8125 2782 -8102
rect 2882 -8041 2932 -7995
rect 2882 -8068 2947 -8041
rect 2882 -8102 2893 -8068
rect 2927 -8102 2947 -8068
rect 2882 -8125 2947 -8102
rect 2977 -8068 3048 -8041
rect 2977 -8102 2991 -8068
rect 3025 -8102 3048 -8068
rect 2977 -8125 3048 -8102
rect 3194 -8053 3246 -8015
rect 3194 -8087 3202 -8053
rect 3236 -8087 3246 -8053
rect 3194 -8125 3246 -8087
rect 3456 -8053 3508 -8015
rect 3456 -8087 3466 -8053
rect 3500 -8087 3508 -8053
rect 3456 -8125 3508 -8087
rect 4390 -8060 4442 -8015
rect 4390 -8094 4398 -8060
rect 4432 -8094 4442 -8060
rect 4390 -8125 4442 -8094
rect 5388 -8060 5440 -8015
rect 5388 -8094 5398 -8060
rect 5432 -8094 5440 -8060
rect 5388 -8125 5440 -8094
rect 6414 -8053 6466 -8015
rect 6414 -8087 6422 -8053
rect 6456 -8087 6466 -8053
rect 6414 -8125 6466 -8087
rect 6676 -8053 6728 -8015
rect 6676 -8087 6686 -8053
rect 6720 -8087 6728 -8053
rect 6676 -8125 6728 -8087
rect 6980 -8041 7030 -7995
rect 6874 -8068 6928 -8041
rect 6874 -8102 6883 -8068
rect 6917 -8102 6928 -8068
rect 6874 -8125 6928 -8102
rect 6958 -8068 7030 -8041
rect 6958 -8102 6980 -8068
rect 7014 -8102 7030 -8068
rect 6958 -8125 7030 -8102
rect 7130 -8068 7182 -7995
rect 7130 -8102 7140 -8068
rect 7174 -8102 7182 -8068
rect 7130 -8125 7182 -8102
rect 7237 -8068 7290 -7995
rect 7237 -8102 7245 -8068
rect 7279 -8102 7290 -8068
rect 7237 -8125 7290 -8102
rect 7390 -8041 7440 -7995
rect 7390 -8068 7455 -8041
rect 7390 -8102 7401 -8068
rect 7435 -8102 7455 -8068
rect 7390 -8125 7455 -8102
rect 7485 -8068 7556 -8041
rect 7485 -8102 7499 -8068
rect 7533 -8102 7556 -8068
rect 7485 -8125 7556 -8102
rect 7702 -8053 7754 -8015
rect 7702 -8087 7710 -8053
rect 7744 -8087 7754 -8053
rect 7702 -8125 7754 -8087
rect 7964 -8053 8016 -8015
rect 7964 -8087 7974 -8053
rect 8008 -8087 8016 -8053
rect 7964 -8125 8016 -8087
rect 8268 -8041 8318 -7995
rect 8162 -8068 8216 -8041
rect 8162 -8102 8171 -8068
rect 8205 -8102 8216 -8068
rect 8162 -8125 8216 -8102
rect 8246 -8068 8318 -8041
rect 8246 -8102 8268 -8068
rect 8302 -8102 8318 -8068
rect 8246 -8125 8318 -8102
rect 8418 -8068 8470 -7995
rect 8418 -8102 8428 -8068
rect 8462 -8102 8470 -8068
rect 8418 -8125 8470 -8102
rect 8525 -8068 8578 -7995
rect 8525 -8102 8533 -8068
rect 8567 -8102 8578 -8068
rect 8525 -8125 8578 -8102
rect 8678 -8041 8728 -7995
rect 8678 -8068 8743 -8041
rect 8678 -8102 8689 -8068
rect 8723 -8102 8743 -8068
rect 8678 -8125 8743 -8102
rect 8773 -8068 8844 -8041
rect 8773 -8102 8787 -8068
rect 8821 -8102 8844 -8068
rect 8773 -8125 8844 -8102
rect 8990 -8053 9042 -8015
rect 8990 -8087 8998 -8053
rect 9032 -8087 9042 -8053
rect 8990 -8125 9042 -8087
rect 9252 -8053 9304 -8015
rect 9252 -8087 9262 -8053
rect 9296 -8087 9304 -8053
rect 9252 -8125 9304 -8087
rect 9556 -8041 9606 -7995
rect 9450 -8068 9504 -8041
rect 9450 -8102 9459 -8068
rect 9493 -8102 9504 -8068
rect 9450 -8125 9504 -8102
rect 9534 -8068 9606 -8041
rect 9534 -8102 9556 -8068
rect 9590 -8102 9606 -8068
rect 9534 -8125 9606 -8102
rect 9706 -8068 9758 -7995
rect 9706 -8102 9716 -8068
rect 9750 -8102 9758 -8068
rect 9706 -8125 9758 -8102
rect 9813 -8068 9866 -7995
rect 9813 -8102 9821 -8068
rect 9855 -8102 9866 -8068
rect 9813 -8125 9866 -8102
rect 9966 -8041 10016 -7995
rect 9966 -8068 10031 -8041
rect 9966 -8102 9977 -8068
rect 10011 -8102 10031 -8068
rect 9966 -8125 10031 -8102
rect 10061 -8068 10132 -8041
rect 10061 -8102 10075 -8068
rect 10109 -8102 10132 -8068
rect 10061 -8125 10132 -8102
rect 10278 -8053 10330 -8015
rect 10278 -8087 10286 -8053
rect 10320 -8087 10330 -8053
rect 10278 -8125 10330 -8087
rect 10540 -8053 10592 -8015
rect 10540 -8087 10550 -8053
rect 10584 -8087 10592 -8053
rect 10540 -8125 10592 -8087
rect 10738 -8011 10790 -7995
rect 10738 -8045 10746 -8011
rect 10780 -8045 10790 -8011
rect 10738 -8079 10790 -8045
rect 10738 -8113 10746 -8079
rect 10780 -8113 10790 -8079
rect 10738 -8125 10790 -8113
rect 10820 -8079 10874 -7995
rect 10820 -8113 10830 -8079
rect 10864 -8113 10874 -8079
rect 10820 -8125 10874 -8113
rect 10904 -8011 10958 -7995
rect 10904 -8045 10914 -8011
rect 10948 -8045 10958 -8011
rect 10904 -8079 10958 -8045
rect 10904 -8113 10914 -8079
rect 10948 -8113 10958 -8079
rect 10904 -8125 10958 -8113
rect 10988 -8079 11042 -7995
rect 10988 -8113 10998 -8079
rect 11032 -8113 11042 -8079
rect 10988 -8125 11042 -8113
rect 11072 -8011 11126 -7995
rect 11072 -8045 11082 -8011
rect 11116 -8045 11126 -8011
rect 11072 -8079 11126 -8045
rect 11072 -8113 11082 -8079
rect 11116 -8113 11126 -8079
rect 11072 -8125 11126 -8113
rect 11156 -8011 11210 -7995
rect 11156 -8045 11166 -8011
rect 11200 -8045 11210 -8011
rect 11156 -8125 11210 -8045
rect 11240 -8079 11294 -7995
rect 11240 -8113 11250 -8079
rect 11284 -8113 11294 -8079
rect 11240 -8125 11294 -8113
rect 11324 -8011 11378 -7995
rect 11324 -8045 11334 -8011
rect 11368 -8045 11378 -8011
rect 11324 -8125 11378 -8045
rect 11408 -8011 11460 -7995
rect 11408 -8045 11418 -8011
rect 11452 -8045 11460 -8011
rect 11408 -8079 11460 -8045
rect 11408 -8113 11418 -8079
rect 11452 -8113 11460 -8079
rect 11658 -8053 11710 -8015
rect 11658 -8087 11666 -8053
rect 11700 -8087 11710 -8053
rect 11408 -8125 11460 -8113
rect 11658 -8125 11710 -8087
rect 11920 -8053 11972 -8015
rect 11920 -8087 11930 -8053
rect 11964 -8087 11972 -8053
rect 11920 -8125 11972 -8087
rect 13590 -8060 13642 -8015
rect 13590 -8094 13598 -8060
rect 13632 -8094 13642 -8060
rect 13590 -8125 13642 -8094
rect 14588 -8060 14640 -8015
rect 14588 -8094 14598 -8060
rect 14632 -8094 14640 -8060
rect 14588 -8125 14640 -8094
rect 14786 -8060 14838 -8015
rect 14786 -8094 14794 -8060
rect 14828 -8094 14838 -8060
rect 14786 -8125 14838 -8094
rect 15784 -8060 15836 -8015
rect 15784 -8094 15794 -8060
rect 15828 -8094 15836 -8060
rect 15784 -8125 15836 -8094
rect 15982 -8060 16034 -8015
rect 15982 -8094 15990 -8060
rect 16024 -8094 16034 -8060
rect 15982 -8125 16034 -8094
rect 16612 -8060 16664 -8015
rect 16612 -8094 16622 -8060
rect 16656 -8094 16664 -8060
rect 16612 -8125 16664 -8094
rect -2970 -8250 -2918 -8219
rect -2970 -8284 -2962 -8250
rect -2928 -8284 -2918 -8250
rect -2970 -8329 -2918 -8284
rect -2340 -8250 -2288 -8219
rect -2340 -8284 -2330 -8250
rect -2296 -8284 -2288 -8250
rect -2340 -8329 -2288 -8284
rect -1590 -8250 -1538 -8219
rect -1590 -8284 -1582 -8250
rect -1548 -8284 -1538 -8250
rect -1590 -8329 -1538 -8284
rect -960 -8250 -908 -8219
rect -960 -8284 -950 -8250
rect -916 -8284 -908 -8250
rect -960 -8329 -908 -8284
rect -854 -8250 -802 -8219
rect -854 -8284 -846 -8250
rect -812 -8284 -802 -8250
rect -854 -8329 -802 -8284
rect -224 -8250 -172 -8219
rect -224 -8284 -214 -8250
rect -180 -8284 -172 -8250
rect -224 -8329 -172 -8284
rect -26 -8257 26 -8219
rect -26 -8291 -18 -8257
rect 16 -8291 26 -8257
rect -26 -8329 26 -8291
rect 236 -8257 288 -8219
rect 236 -8291 246 -8257
rect 280 -8291 288 -8257
rect 236 -8329 288 -8291
rect 434 -8242 505 -8219
rect 434 -8276 457 -8242
rect 491 -8276 505 -8242
rect 434 -8303 505 -8276
rect 535 -8242 600 -8219
rect 535 -8276 555 -8242
rect 589 -8276 600 -8242
rect 535 -8303 600 -8276
rect 550 -8349 600 -8303
rect 700 -8242 753 -8219
rect 700 -8276 711 -8242
rect 745 -8276 753 -8242
rect 700 -8349 753 -8276
rect 808 -8242 860 -8219
rect 808 -8276 816 -8242
rect 850 -8276 860 -8242
rect 808 -8349 860 -8276
rect 960 -8242 1032 -8219
rect 960 -8276 976 -8242
rect 1010 -8276 1032 -8242
rect 960 -8303 1032 -8276
rect 1062 -8242 1116 -8219
rect 1062 -8276 1073 -8242
rect 1107 -8276 1116 -8242
rect 1062 -8303 1116 -8276
rect 960 -8349 1010 -8303
rect 1262 -8257 1314 -8219
rect 1262 -8291 1270 -8257
rect 1304 -8291 1314 -8257
rect 1262 -8329 1314 -8291
rect 1524 -8257 1576 -8219
rect 1524 -8291 1534 -8257
rect 1568 -8291 1576 -8257
rect 1524 -8329 1576 -8291
rect 1722 -8250 1774 -8219
rect 1722 -8284 1730 -8250
rect 1764 -8284 1774 -8250
rect 1722 -8329 1774 -8284
rect 2352 -8250 2404 -8219
rect 2352 -8284 2362 -8250
rect 2396 -8284 2404 -8250
rect 2352 -8329 2404 -8284
rect 2550 -8257 2602 -8219
rect 2550 -8291 2558 -8257
rect 2592 -8291 2602 -8257
rect 2550 -8329 2602 -8291
rect 2812 -8257 2864 -8219
rect 2812 -8291 2822 -8257
rect 2856 -8291 2864 -8257
rect 2812 -8329 2864 -8291
rect 3010 -8242 3081 -8219
rect 3010 -8276 3033 -8242
rect 3067 -8276 3081 -8242
rect 3010 -8303 3081 -8276
rect 3111 -8242 3176 -8219
rect 3111 -8276 3131 -8242
rect 3165 -8276 3176 -8242
rect 3111 -8303 3176 -8276
rect 3126 -8349 3176 -8303
rect 3276 -8242 3329 -8219
rect 3276 -8276 3287 -8242
rect 3321 -8276 3329 -8242
rect 3276 -8349 3329 -8276
rect 3384 -8242 3436 -8219
rect 3384 -8276 3392 -8242
rect 3426 -8276 3436 -8242
rect 3384 -8349 3436 -8276
rect 3536 -8242 3608 -8219
rect 3536 -8276 3552 -8242
rect 3586 -8276 3608 -8242
rect 3536 -8303 3608 -8276
rect 3638 -8242 3692 -8219
rect 3638 -8276 3649 -8242
rect 3683 -8276 3692 -8242
rect 3638 -8303 3692 -8276
rect 3536 -8349 3586 -8303
rect 3838 -8257 3890 -8219
rect 3838 -8291 3846 -8257
rect 3880 -8291 3890 -8257
rect 3838 -8329 3890 -8291
rect 4100 -8257 4152 -8219
rect 4100 -8291 4110 -8257
rect 4144 -8291 4152 -8257
rect 4100 -8329 4152 -8291
rect 4298 -8250 4350 -8219
rect 4298 -8284 4306 -8250
rect 4340 -8284 4350 -8250
rect 4298 -8329 4350 -8284
rect 4928 -8250 4980 -8219
rect 4928 -8284 4938 -8250
rect 4972 -8284 4980 -8250
rect 4928 -8329 4980 -8284
rect 5126 -8257 5178 -8219
rect 5126 -8291 5134 -8257
rect 5168 -8291 5178 -8257
rect 5126 -8329 5178 -8291
rect 5388 -8257 5440 -8219
rect 5388 -8291 5398 -8257
rect 5432 -8291 5440 -8257
rect 5388 -8329 5440 -8291
rect 5586 -8242 5657 -8219
rect 5586 -8276 5609 -8242
rect 5643 -8276 5657 -8242
rect 5586 -8303 5657 -8276
rect 5687 -8242 5752 -8219
rect 5687 -8276 5707 -8242
rect 5741 -8276 5752 -8242
rect 5687 -8303 5752 -8276
rect 5702 -8349 5752 -8303
rect 5852 -8242 5905 -8219
rect 5852 -8276 5863 -8242
rect 5897 -8276 5905 -8242
rect 5852 -8349 5905 -8276
rect 5960 -8242 6012 -8219
rect 5960 -8276 5968 -8242
rect 6002 -8276 6012 -8242
rect 5960 -8349 6012 -8276
rect 6112 -8242 6184 -8219
rect 6112 -8276 6128 -8242
rect 6162 -8276 6184 -8242
rect 6112 -8303 6184 -8276
rect 6214 -8242 6268 -8219
rect 6214 -8276 6225 -8242
rect 6259 -8276 6268 -8242
rect 6214 -8303 6268 -8276
rect 6112 -8349 6162 -8303
rect 6414 -8257 6466 -8219
rect 6414 -8291 6422 -8257
rect 6456 -8291 6466 -8257
rect 6414 -8329 6466 -8291
rect 6676 -8257 6728 -8219
rect 6676 -8291 6686 -8257
rect 6720 -8291 6728 -8257
rect 6676 -8329 6728 -8291
rect 6874 -8250 6926 -8219
rect 6874 -8284 6882 -8250
rect 6916 -8284 6926 -8250
rect 6874 -8329 6926 -8284
rect 7504 -8250 7556 -8219
rect 7504 -8284 7514 -8250
rect 7548 -8284 7556 -8250
rect 7504 -8329 7556 -8284
rect 7702 -8257 7754 -8219
rect 7702 -8291 7710 -8257
rect 7744 -8291 7754 -8257
rect 7702 -8329 7754 -8291
rect 7964 -8257 8016 -8219
rect 7964 -8291 7974 -8257
rect 8008 -8291 8016 -8257
rect 7964 -8329 8016 -8291
rect 8162 -8242 8233 -8219
rect 8162 -8276 8185 -8242
rect 8219 -8276 8233 -8242
rect 8162 -8303 8233 -8276
rect 8263 -8242 8328 -8219
rect 8263 -8276 8283 -8242
rect 8317 -8276 8328 -8242
rect 8263 -8303 8328 -8276
rect 8278 -8349 8328 -8303
rect 8428 -8242 8481 -8219
rect 8428 -8276 8439 -8242
rect 8473 -8276 8481 -8242
rect 8428 -8349 8481 -8276
rect 8536 -8242 8588 -8219
rect 8536 -8276 8544 -8242
rect 8578 -8276 8588 -8242
rect 8536 -8349 8588 -8276
rect 8688 -8242 8760 -8219
rect 8688 -8276 8704 -8242
rect 8738 -8276 8760 -8242
rect 8688 -8303 8760 -8276
rect 8790 -8242 8844 -8219
rect 8790 -8276 8801 -8242
rect 8835 -8276 8844 -8242
rect 8790 -8303 8844 -8276
rect 8688 -8349 8738 -8303
rect 8990 -8257 9042 -8219
rect 8990 -8291 8998 -8257
rect 9032 -8291 9042 -8257
rect 8990 -8329 9042 -8291
rect 9252 -8257 9304 -8219
rect 9252 -8291 9262 -8257
rect 9296 -8291 9304 -8257
rect 9252 -8329 9304 -8291
rect 9450 -8250 9502 -8219
rect 9450 -8284 9458 -8250
rect 9492 -8284 9502 -8250
rect 9450 -8329 9502 -8284
rect 10080 -8250 10132 -8219
rect 10080 -8284 10090 -8250
rect 10124 -8284 10132 -8250
rect 10080 -8329 10132 -8284
rect 10370 -8257 10422 -8219
rect 10370 -8291 10378 -8257
rect 10412 -8291 10422 -8257
rect 10370 -8329 10422 -8291
rect 10632 -8257 10684 -8219
rect 10632 -8291 10642 -8257
rect 10676 -8291 10684 -8257
rect 10632 -8329 10684 -8291
rect 10738 -8242 10809 -8219
rect 10738 -8276 10761 -8242
rect 10795 -8276 10809 -8242
rect 10738 -8303 10809 -8276
rect 10839 -8242 10904 -8219
rect 10839 -8276 10859 -8242
rect 10893 -8276 10904 -8242
rect 10839 -8303 10904 -8276
rect 10854 -8349 10904 -8303
rect 11004 -8242 11057 -8219
rect 11004 -8276 11015 -8242
rect 11049 -8276 11057 -8242
rect 11004 -8349 11057 -8276
rect 11112 -8242 11164 -8219
rect 11112 -8276 11120 -8242
rect 11154 -8276 11164 -8242
rect 11112 -8349 11164 -8276
rect 11264 -8242 11336 -8219
rect 11264 -8276 11280 -8242
rect 11314 -8276 11336 -8242
rect 11264 -8303 11336 -8276
rect 11366 -8242 11420 -8219
rect 11366 -8276 11377 -8242
rect 11411 -8276 11420 -8242
rect 11366 -8303 11420 -8276
rect 11264 -8349 11314 -8303
rect 11658 -8257 11710 -8219
rect 11658 -8291 11666 -8257
rect 11700 -8291 11710 -8257
rect 11658 -8329 11710 -8291
rect 11920 -8257 11972 -8219
rect 13682 -8231 13735 -8219
rect 11920 -8291 11930 -8257
rect 11964 -8291 11972 -8257
rect 11920 -8329 11972 -8291
rect 13682 -8265 13690 -8231
rect 13724 -8265 13735 -8231
rect 13682 -8303 13735 -8265
rect 13765 -8244 13821 -8219
rect 13765 -8278 13776 -8244
rect 13810 -8278 13821 -8244
rect 13765 -8303 13821 -8278
rect 13851 -8244 13907 -8219
rect 13851 -8278 13862 -8244
rect 13896 -8278 13907 -8244
rect 13851 -8303 13907 -8278
rect 13937 -8244 13993 -8219
rect 13937 -8278 13948 -8244
rect 13982 -8278 13993 -8244
rect 13937 -8303 13993 -8278
rect 14023 -8244 14079 -8219
rect 14023 -8278 14034 -8244
rect 14068 -8278 14079 -8244
rect 14023 -8303 14079 -8278
rect 14109 -8244 14165 -8219
rect 14109 -8278 14120 -8244
rect 14154 -8278 14165 -8244
rect 14109 -8303 14165 -8278
rect 14195 -8235 14251 -8219
rect 14195 -8269 14206 -8235
rect 14240 -8269 14251 -8235
rect 14195 -8303 14251 -8269
rect 14281 -8244 14337 -8219
rect 14281 -8278 14292 -8244
rect 14326 -8278 14337 -8244
rect 14281 -8303 14337 -8278
rect 14367 -8235 14423 -8219
rect 14367 -8269 14378 -8235
rect 14412 -8269 14423 -8235
rect 14367 -8303 14423 -8269
rect 14453 -8244 14509 -8219
rect 14453 -8278 14464 -8244
rect 14498 -8278 14509 -8244
rect 14453 -8303 14509 -8278
rect 14539 -8235 14595 -8219
rect 14539 -8269 14550 -8235
rect 14584 -8269 14595 -8235
rect 14539 -8303 14595 -8269
rect 14625 -8244 14681 -8219
rect 14625 -8278 14636 -8244
rect 14670 -8278 14681 -8244
rect 14625 -8303 14681 -8278
rect 14711 -8235 14766 -8219
rect 14711 -8269 14722 -8235
rect 14756 -8269 14766 -8235
rect 14711 -8303 14766 -8269
rect 14796 -8244 14852 -8219
rect 14796 -8278 14807 -8244
rect 14841 -8278 14852 -8244
rect 14796 -8303 14852 -8278
rect 14882 -8235 14938 -8219
rect 14882 -8269 14893 -8235
rect 14927 -8269 14938 -8235
rect 14882 -8303 14938 -8269
rect 14968 -8244 15024 -8219
rect 14968 -8278 14979 -8244
rect 15013 -8278 15024 -8244
rect 14968 -8303 15024 -8278
rect 15054 -8235 15110 -8219
rect 15054 -8269 15065 -8235
rect 15099 -8269 15110 -8235
rect 15054 -8303 15110 -8269
rect 15140 -8244 15196 -8219
rect 15140 -8278 15151 -8244
rect 15185 -8278 15196 -8244
rect 15140 -8303 15196 -8278
rect 15226 -8235 15282 -8219
rect 15226 -8269 15237 -8235
rect 15271 -8269 15282 -8235
rect 15226 -8303 15282 -8269
rect 15312 -8244 15368 -8219
rect 15312 -8278 15323 -8244
rect 15357 -8278 15368 -8244
rect 15312 -8303 15368 -8278
rect 15398 -8235 15451 -8219
rect 15398 -8269 15409 -8235
rect 15443 -8269 15451 -8235
rect 15398 -8303 15451 -8269
rect 15614 -8250 15666 -8219
rect 15614 -8284 15622 -8250
rect 15656 -8284 15666 -8250
rect 15614 -8329 15666 -8284
rect 16612 -8250 16664 -8219
rect 16612 -8284 16622 -8250
rect 16656 -8284 16664 -8250
rect 16612 -8329 16664 -8284
rect -2970 -9148 -2918 -9103
rect -2970 -9182 -2962 -9148
rect -2928 -9182 -2918 -9148
rect -2970 -9213 -2918 -9182
rect -2340 -9148 -2288 -9103
rect -2340 -9182 -2330 -9148
rect -2296 -9182 -2288 -9148
rect -2340 -9213 -2288 -9182
rect -1590 -9148 -1538 -9103
rect -1590 -9182 -1582 -9148
rect -1548 -9182 -1538 -9148
rect -1590 -9213 -1538 -9182
rect -960 -9148 -908 -9103
rect -960 -9182 -950 -9148
rect -916 -9182 -908 -9148
rect -960 -9213 -908 -9182
rect -854 -9148 -802 -9103
rect -854 -9182 -846 -9148
rect -812 -9182 -802 -9148
rect -854 -9213 -802 -9182
rect -224 -9148 -172 -9103
rect -224 -9182 -214 -9148
rect -180 -9182 -172 -9148
rect -224 -9213 -172 -9182
rect -26 -9141 26 -9103
rect -26 -9175 -18 -9141
rect 16 -9175 26 -9141
rect -26 -9213 26 -9175
rect 236 -9141 288 -9103
rect 236 -9175 246 -9141
rect 280 -9175 288 -9141
rect 236 -9213 288 -9175
rect 540 -9129 590 -9083
rect 434 -9156 488 -9129
rect 434 -9190 443 -9156
rect 477 -9190 488 -9156
rect 434 -9213 488 -9190
rect 518 -9156 590 -9129
rect 518 -9190 540 -9156
rect 574 -9190 590 -9156
rect 518 -9213 590 -9190
rect 690 -9156 742 -9083
rect 690 -9190 700 -9156
rect 734 -9190 742 -9156
rect 690 -9213 742 -9190
rect 797 -9156 850 -9083
rect 797 -9190 805 -9156
rect 839 -9190 850 -9156
rect 797 -9213 850 -9190
rect 950 -9129 1000 -9083
rect 950 -9156 1015 -9129
rect 950 -9190 961 -9156
rect 995 -9190 1015 -9156
rect 950 -9213 1015 -9190
rect 1045 -9156 1116 -9129
rect 1045 -9190 1059 -9156
rect 1093 -9190 1116 -9156
rect 1045 -9213 1116 -9190
rect 1262 -9141 1314 -9103
rect 1262 -9175 1270 -9141
rect 1304 -9175 1314 -9141
rect 1262 -9213 1314 -9175
rect 1524 -9141 1576 -9103
rect 1524 -9175 1534 -9141
rect 1568 -9175 1576 -9141
rect 1524 -9213 1576 -9175
rect 1722 -9148 1774 -9103
rect 1722 -9182 1730 -9148
rect 1764 -9182 1774 -9148
rect 1722 -9213 1774 -9182
rect 2352 -9148 2404 -9103
rect 2352 -9182 2362 -9148
rect 2396 -9182 2404 -9148
rect 2352 -9213 2404 -9182
rect 2550 -9141 2602 -9103
rect 2550 -9175 2558 -9141
rect 2592 -9175 2602 -9141
rect 2550 -9213 2602 -9175
rect 2812 -9141 2864 -9103
rect 2812 -9175 2822 -9141
rect 2856 -9175 2864 -9141
rect 2812 -9213 2864 -9175
rect 3116 -9129 3166 -9083
rect 3010 -9156 3064 -9129
rect 3010 -9190 3019 -9156
rect 3053 -9190 3064 -9156
rect 3010 -9213 3064 -9190
rect 3094 -9156 3166 -9129
rect 3094 -9190 3116 -9156
rect 3150 -9190 3166 -9156
rect 3094 -9213 3166 -9190
rect 3266 -9156 3318 -9083
rect 3266 -9190 3276 -9156
rect 3310 -9190 3318 -9156
rect 3266 -9213 3318 -9190
rect 3373 -9156 3426 -9083
rect 3373 -9190 3381 -9156
rect 3415 -9190 3426 -9156
rect 3373 -9213 3426 -9190
rect 3526 -9129 3576 -9083
rect 3526 -9156 3591 -9129
rect 3526 -9190 3537 -9156
rect 3571 -9190 3591 -9156
rect 3526 -9213 3591 -9190
rect 3621 -9156 3692 -9129
rect 3621 -9190 3635 -9156
rect 3669 -9190 3692 -9156
rect 3621 -9213 3692 -9190
rect 3838 -9141 3890 -9103
rect 3838 -9175 3846 -9141
rect 3880 -9175 3890 -9141
rect 3838 -9213 3890 -9175
rect 4100 -9141 4152 -9103
rect 4100 -9175 4110 -9141
rect 4144 -9175 4152 -9141
rect 4100 -9213 4152 -9175
rect 4298 -9148 4350 -9103
rect 4298 -9182 4306 -9148
rect 4340 -9182 4350 -9148
rect 4298 -9213 4350 -9182
rect 4928 -9148 4980 -9103
rect 4928 -9182 4938 -9148
rect 4972 -9182 4980 -9148
rect 4928 -9213 4980 -9182
rect 5126 -9141 5178 -9103
rect 5126 -9175 5134 -9141
rect 5168 -9175 5178 -9141
rect 5126 -9213 5178 -9175
rect 5388 -9141 5440 -9103
rect 5388 -9175 5398 -9141
rect 5432 -9175 5440 -9141
rect 5388 -9213 5440 -9175
rect 5692 -9129 5742 -9083
rect 5586 -9156 5640 -9129
rect 5586 -9190 5595 -9156
rect 5629 -9190 5640 -9156
rect 5586 -9213 5640 -9190
rect 5670 -9156 5742 -9129
rect 5670 -9190 5692 -9156
rect 5726 -9190 5742 -9156
rect 5670 -9213 5742 -9190
rect 5842 -9156 5894 -9083
rect 5842 -9190 5852 -9156
rect 5886 -9190 5894 -9156
rect 5842 -9213 5894 -9190
rect 5949 -9156 6002 -9083
rect 5949 -9190 5957 -9156
rect 5991 -9190 6002 -9156
rect 5949 -9213 6002 -9190
rect 6102 -9129 6152 -9083
rect 6102 -9156 6167 -9129
rect 6102 -9190 6113 -9156
rect 6147 -9190 6167 -9156
rect 6102 -9213 6167 -9190
rect 6197 -9156 6268 -9129
rect 6197 -9190 6211 -9156
rect 6245 -9190 6268 -9156
rect 6197 -9213 6268 -9190
rect 6414 -9141 6466 -9103
rect 6414 -9175 6422 -9141
rect 6456 -9175 6466 -9141
rect 6414 -9213 6466 -9175
rect 6676 -9141 6728 -9103
rect 6676 -9175 6686 -9141
rect 6720 -9175 6728 -9141
rect 6676 -9213 6728 -9175
rect 6874 -9148 6926 -9103
rect 6874 -9182 6882 -9148
rect 6916 -9182 6926 -9148
rect 6874 -9213 6926 -9182
rect 7504 -9148 7556 -9103
rect 7504 -9182 7514 -9148
rect 7548 -9182 7556 -9148
rect 7504 -9213 7556 -9182
rect 7702 -9141 7754 -9103
rect 7702 -9175 7710 -9141
rect 7744 -9175 7754 -9141
rect 7702 -9213 7754 -9175
rect 7964 -9141 8016 -9103
rect 7964 -9175 7974 -9141
rect 8008 -9175 8016 -9141
rect 7964 -9213 8016 -9175
rect 8268 -9129 8318 -9083
rect 8162 -9156 8216 -9129
rect 8162 -9190 8171 -9156
rect 8205 -9190 8216 -9156
rect 8162 -9213 8216 -9190
rect 8246 -9156 8318 -9129
rect 8246 -9190 8268 -9156
rect 8302 -9190 8318 -9156
rect 8246 -9213 8318 -9190
rect 8418 -9156 8470 -9083
rect 8418 -9190 8428 -9156
rect 8462 -9190 8470 -9156
rect 8418 -9213 8470 -9190
rect 8525 -9156 8578 -9083
rect 8525 -9190 8533 -9156
rect 8567 -9190 8578 -9156
rect 8525 -9213 8578 -9190
rect 8678 -9129 8728 -9083
rect 8678 -9156 8743 -9129
rect 8678 -9190 8689 -9156
rect 8723 -9190 8743 -9156
rect 8678 -9213 8743 -9190
rect 8773 -9156 8844 -9129
rect 8773 -9190 8787 -9156
rect 8821 -9190 8844 -9156
rect 8773 -9213 8844 -9190
rect 8990 -9141 9042 -9103
rect 8990 -9175 8998 -9141
rect 9032 -9175 9042 -9141
rect 8990 -9213 9042 -9175
rect 9252 -9141 9304 -9103
rect 9252 -9175 9262 -9141
rect 9296 -9175 9304 -9141
rect 9252 -9213 9304 -9175
rect 9450 -9148 9502 -9103
rect 9450 -9182 9458 -9148
rect 9492 -9182 9502 -9148
rect 9450 -9213 9502 -9182
rect 10080 -9148 10132 -9103
rect 10080 -9182 10090 -9148
rect 10124 -9182 10132 -9148
rect 10080 -9213 10132 -9182
rect 10370 -9141 10422 -9103
rect 10370 -9175 10378 -9141
rect 10412 -9175 10422 -9141
rect 10370 -9213 10422 -9175
rect 10632 -9141 10684 -9103
rect 10844 -9129 10894 -9083
rect 10632 -9175 10642 -9141
rect 10676 -9175 10684 -9141
rect 10632 -9213 10684 -9175
rect 10738 -9156 10792 -9129
rect 10738 -9190 10747 -9156
rect 10781 -9190 10792 -9156
rect 10738 -9213 10792 -9190
rect 10822 -9156 10894 -9129
rect 10822 -9190 10844 -9156
rect 10878 -9190 10894 -9156
rect 10822 -9213 10894 -9190
rect 10994 -9156 11046 -9083
rect 10994 -9190 11004 -9156
rect 11038 -9190 11046 -9156
rect 10994 -9213 11046 -9190
rect 11101 -9156 11154 -9083
rect 11101 -9190 11109 -9156
rect 11143 -9190 11154 -9156
rect 11101 -9213 11154 -9190
rect 11254 -9129 11304 -9083
rect 11254 -9156 11319 -9129
rect 11254 -9190 11265 -9156
rect 11299 -9190 11319 -9156
rect 11254 -9213 11319 -9190
rect 11349 -9156 11420 -9129
rect 11349 -9190 11363 -9156
rect 11397 -9190 11420 -9156
rect 11349 -9213 11420 -9190
rect 11658 -9141 11710 -9103
rect 11658 -9175 11666 -9141
rect 11700 -9175 11710 -9141
rect 11658 -9213 11710 -9175
rect 11920 -9141 11972 -9103
rect 11920 -9175 11930 -9141
rect 11964 -9175 11972 -9141
rect 11920 -9213 11972 -9175
rect 12567 -9165 12633 -9129
rect 12567 -9199 12588 -9165
rect 12622 -9199 12633 -9165
rect 12567 -9213 12633 -9199
rect 12663 -9154 12719 -9129
rect 12663 -9188 12674 -9154
rect 12708 -9188 12719 -9154
rect 12663 -9213 12719 -9188
rect 12749 -9165 12805 -9129
rect 12749 -9199 12760 -9165
rect 12794 -9199 12805 -9165
rect 12749 -9213 12805 -9199
rect 12835 -9154 12891 -9129
rect 12835 -9188 12846 -9154
rect 12880 -9188 12891 -9154
rect 12835 -9213 12891 -9188
rect 12921 -9165 13000 -9129
rect 12921 -9199 12932 -9165
rect 12966 -9199 13000 -9165
rect 13222 -9141 13274 -9103
rect 13222 -9175 13230 -9141
rect 13264 -9175 13274 -9141
rect 12921 -9213 13000 -9199
rect 13222 -9213 13274 -9175
rect 13484 -9141 13536 -9103
rect 13484 -9175 13494 -9141
rect 13528 -9175 13536 -9141
rect 13484 -9213 13536 -9175
rect 13682 -9167 13735 -9129
rect 13682 -9201 13690 -9167
rect 13724 -9201 13735 -9167
rect 13682 -9213 13735 -9201
rect 13765 -9154 13821 -9129
rect 13765 -9188 13776 -9154
rect 13810 -9188 13821 -9154
rect 13765 -9213 13821 -9188
rect 13851 -9154 13907 -9129
rect 13851 -9188 13862 -9154
rect 13896 -9188 13907 -9154
rect 13851 -9213 13907 -9188
rect 13937 -9154 13993 -9129
rect 13937 -9188 13948 -9154
rect 13982 -9188 13993 -9154
rect 13937 -9213 13993 -9188
rect 14023 -9154 14079 -9129
rect 14023 -9188 14034 -9154
rect 14068 -9188 14079 -9154
rect 14023 -9213 14079 -9188
rect 14109 -9154 14165 -9129
rect 14109 -9188 14120 -9154
rect 14154 -9188 14165 -9154
rect 14109 -9213 14165 -9188
rect 14195 -9163 14251 -9129
rect 14195 -9197 14206 -9163
rect 14240 -9197 14251 -9163
rect 14195 -9213 14251 -9197
rect 14281 -9154 14337 -9129
rect 14281 -9188 14292 -9154
rect 14326 -9188 14337 -9154
rect 14281 -9213 14337 -9188
rect 14367 -9163 14423 -9129
rect 14367 -9197 14378 -9163
rect 14412 -9197 14423 -9163
rect 14367 -9213 14423 -9197
rect 14453 -9154 14509 -9129
rect 14453 -9188 14464 -9154
rect 14498 -9188 14509 -9154
rect 14453 -9213 14509 -9188
rect 14539 -9163 14595 -9129
rect 14539 -9197 14550 -9163
rect 14584 -9197 14595 -9163
rect 14539 -9213 14595 -9197
rect 14625 -9154 14681 -9129
rect 14625 -9188 14636 -9154
rect 14670 -9188 14681 -9154
rect 14625 -9213 14681 -9188
rect 14711 -9163 14766 -9129
rect 14711 -9197 14722 -9163
rect 14756 -9197 14766 -9163
rect 14711 -9213 14766 -9197
rect 14796 -9154 14852 -9129
rect 14796 -9188 14807 -9154
rect 14841 -9188 14852 -9154
rect 14796 -9213 14852 -9188
rect 14882 -9163 14938 -9129
rect 14882 -9197 14893 -9163
rect 14927 -9197 14938 -9163
rect 14882 -9213 14938 -9197
rect 14968 -9154 15024 -9129
rect 14968 -9188 14979 -9154
rect 15013 -9188 15024 -9154
rect 14968 -9213 15024 -9188
rect 15054 -9163 15110 -9129
rect 15054 -9197 15065 -9163
rect 15099 -9197 15110 -9163
rect 15054 -9213 15110 -9197
rect 15140 -9154 15196 -9129
rect 15140 -9188 15151 -9154
rect 15185 -9188 15196 -9154
rect 15140 -9213 15196 -9188
rect 15226 -9163 15282 -9129
rect 15226 -9197 15237 -9163
rect 15271 -9197 15282 -9163
rect 15226 -9213 15282 -9197
rect 15312 -9154 15368 -9129
rect 15312 -9188 15323 -9154
rect 15357 -9188 15368 -9154
rect 15312 -9213 15368 -9188
rect 15398 -9163 15451 -9129
rect 15398 -9197 15409 -9163
rect 15443 -9197 15451 -9163
rect 15614 -9148 15666 -9103
rect 15614 -9182 15622 -9148
rect 15656 -9182 15666 -9148
rect 15398 -9213 15451 -9197
rect 15614 -9213 15666 -9182
rect 16612 -9148 16664 -9103
rect 16612 -9182 16622 -9148
rect 16656 -9182 16664 -9148
rect 16612 -9213 16664 -9182
rect -2970 -9338 -2918 -9307
rect -2970 -9372 -2962 -9338
rect -2928 -9372 -2918 -9338
rect -2970 -9417 -2918 -9372
rect -2340 -9338 -2288 -9307
rect -2340 -9372 -2330 -9338
rect -2296 -9372 -2288 -9338
rect -2340 -9417 -2288 -9372
rect -1590 -9338 -1538 -9307
rect -1590 -9372 -1582 -9338
rect -1548 -9372 -1538 -9338
rect -1590 -9417 -1538 -9372
rect -960 -9338 -908 -9307
rect -960 -9372 -950 -9338
rect -916 -9372 -908 -9338
rect -960 -9417 -908 -9372
rect -854 -9330 -783 -9307
rect -854 -9364 -831 -9330
rect -797 -9364 -783 -9330
rect -854 -9391 -783 -9364
rect -753 -9330 -688 -9307
rect -753 -9364 -733 -9330
rect -699 -9364 -688 -9330
rect -753 -9391 -688 -9364
rect -738 -9437 -688 -9391
rect -588 -9330 -535 -9307
rect -588 -9364 -577 -9330
rect -543 -9364 -535 -9330
rect -588 -9437 -535 -9364
rect -480 -9330 -428 -9307
rect -480 -9364 -472 -9330
rect -438 -9364 -428 -9330
rect -480 -9437 -428 -9364
rect -328 -9330 -256 -9307
rect -328 -9364 -312 -9330
rect -278 -9364 -256 -9330
rect -328 -9391 -256 -9364
rect -226 -9330 -172 -9307
rect -226 -9364 -215 -9330
rect -181 -9364 -172 -9330
rect -226 -9391 -172 -9364
rect -328 -9437 -278 -9391
rect -26 -9345 26 -9307
rect -26 -9379 -18 -9345
rect 16 -9379 26 -9345
rect -26 -9417 26 -9379
rect 236 -9345 288 -9307
rect 236 -9379 246 -9345
rect 280 -9379 288 -9345
rect 236 -9417 288 -9379
rect 434 -9330 505 -9307
rect 434 -9364 457 -9330
rect 491 -9364 505 -9330
rect 434 -9391 505 -9364
rect 535 -9330 600 -9307
rect 535 -9364 555 -9330
rect 589 -9364 600 -9330
rect 535 -9391 600 -9364
rect 550 -9437 600 -9391
rect 700 -9330 753 -9307
rect 700 -9364 711 -9330
rect 745 -9364 753 -9330
rect 700 -9437 753 -9364
rect 808 -9330 860 -9307
rect 808 -9364 816 -9330
rect 850 -9364 860 -9330
rect 808 -9437 860 -9364
rect 960 -9330 1032 -9307
rect 960 -9364 976 -9330
rect 1010 -9364 1032 -9330
rect 960 -9391 1032 -9364
rect 1062 -9330 1116 -9307
rect 1062 -9364 1073 -9330
rect 1107 -9364 1116 -9330
rect 1062 -9391 1116 -9364
rect 960 -9437 1010 -9391
rect 1262 -9345 1314 -9307
rect 1262 -9379 1270 -9345
rect 1304 -9379 1314 -9345
rect 1262 -9417 1314 -9379
rect 1524 -9345 1576 -9307
rect 1524 -9379 1534 -9345
rect 1568 -9379 1576 -9345
rect 1524 -9417 1576 -9379
rect 1722 -9338 1774 -9307
rect 1722 -9372 1730 -9338
rect 1764 -9372 1774 -9338
rect 1722 -9417 1774 -9372
rect 2352 -9338 2404 -9307
rect 2352 -9372 2362 -9338
rect 2396 -9372 2404 -9338
rect 2352 -9417 2404 -9372
rect 2550 -9345 2602 -9307
rect 2550 -9379 2558 -9345
rect 2592 -9379 2602 -9345
rect 2550 -9417 2602 -9379
rect 2812 -9345 2864 -9307
rect 2812 -9379 2822 -9345
rect 2856 -9379 2864 -9345
rect 2812 -9417 2864 -9379
rect 3010 -9330 3081 -9307
rect 3010 -9364 3033 -9330
rect 3067 -9364 3081 -9330
rect 3010 -9391 3081 -9364
rect 3111 -9330 3176 -9307
rect 3111 -9364 3131 -9330
rect 3165 -9364 3176 -9330
rect 3111 -9391 3176 -9364
rect 3126 -9437 3176 -9391
rect 3276 -9330 3329 -9307
rect 3276 -9364 3287 -9330
rect 3321 -9364 3329 -9330
rect 3276 -9437 3329 -9364
rect 3384 -9330 3436 -9307
rect 3384 -9364 3392 -9330
rect 3426 -9364 3436 -9330
rect 3384 -9437 3436 -9364
rect 3536 -9330 3608 -9307
rect 3536 -9364 3552 -9330
rect 3586 -9364 3608 -9330
rect 3536 -9391 3608 -9364
rect 3638 -9330 3692 -9307
rect 3638 -9364 3649 -9330
rect 3683 -9364 3692 -9330
rect 3638 -9391 3692 -9364
rect 3536 -9437 3586 -9391
rect 3838 -9345 3890 -9307
rect 3838 -9379 3846 -9345
rect 3880 -9379 3890 -9345
rect 3838 -9417 3890 -9379
rect 4100 -9345 4152 -9307
rect 4100 -9379 4110 -9345
rect 4144 -9379 4152 -9345
rect 4100 -9417 4152 -9379
rect 4298 -9338 4350 -9307
rect 4298 -9372 4306 -9338
rect 4340 -9372 4350 -9338
rect 4298 -9417 4350 -9372
rect 4928 -9338 4980 -9307
rect 4928 -9372 4938 -9338
rect 4972 -9372 4980 -9338
rect 4928 -9417 4980 -9372
rect 5126 -9345 5178 -9307
rect 5126 -9379 5134 -9345
rect 5168 -9379 5178 -9345
rect 5126 -9417 5178 -9379
rect 5388 -9345 5440 -9307
rect 5388 -9379 5398 -9345
rect 5432 -9379 5440 -9345
rect 5388 -9417 5440 -9379
rect 5586 -9330 5657 -9307
rect 5586 -9364 5609 -9330
rect 5643 -9364 5657 -9330
rect 5586 -9391 5657 -9364
rect 5687 -9330 5752 -9307
rect 5687 -9364 5707 -9330
rect 5741 -9364 5752 -9330
rect 5687 -9391 5752 -9364
rect 5702 -9437 5752 -9391
rect 5852 -9330 5905 -9307
rect 5852 -9364 5863 -9330
rect 5897 -9364 5905 -9330
rect 5852 -9437 5905 -9364
rect 5960 -9330 6012 -9307
rect 5960 -9364 5968 -9330
rect 6002 -9364 6012 -9330
rect 5960 -9437 6012 -9364
rect 6112 -9330 6184 -9307
rect 6112 -9364 6128 -9330
rect 6162 -9364 6184 -9330
rect 6112 -9391 6184 -9364
rect 6214 -9330 6268 -9307
rect 6214 -9364 6225 -9330
rect 6259 -9364 6268 -9330
rect 6214 -9391 6268 -9364
rect 6112 -9437 6162 -9391
rect 6414 -9345 6466 -9307
rect 6414 -9379 6422 -9345
rect 6456 -9379 6466 -9345
rect 6414 -9417 6466 -9379
rect 6676 -9345 6728 -9307
rect 6676 -9379 6686 -9345
rect 6720 -9379 6728 -9345
rect 6676 -9417 6728 -9379
rect 6874 -9338 6926 -9307
rect 6874 -9372 6882 -9338
rect 6916 -9372 6926 -9338
rect 6874 -9417 6926 -9372
rect 7504 -9338 7556 -9307
rect 7504 -9372 7514 -9338
rect 7548 -9372 7556 -9338
rect 7504 -9417 7556 -9372
rect 7702 -9345 7754 -9307
rect 7702 -9379 7710 -9345
rect 7744 -9379 7754 -9345
rect 7702 -9417 7754 -9379
rect 7964 -9345 8016 -9307
rect 7964 -9379 7974 -9345
rect 8008 -9379 8016 -9345
rect 7964 -9417 8016 -9379
rect 8162 -9330 8233 -9307
rect 8162 -9364 8185 -9330
rect 8219 -9364 8233 -9330
rect 8162 -9391 8233 -9364
rect 8263 -9330 8328 -9307
rect 8263 -9364 8283 -9330
rect 8317 -9364 8328 -9330
rect 8263 -9391 8328 -9364
rect 8278 -9437 8328 -9391
rect 8428 -9330 8481 -9307
rect 8428 -9364 8439 -9330
rect 8473 -9364 8481 -9330
rect 8428 -9437 8481 -9364
rect 8536 -9330 8588 -9307
rect 8536 -9364 8544 -9330
rect 8578 -9364 8588 -9330
rect 8536 -9437 8588 -9364
rect 8688 -9330 8760 -9307
rect 8688 -9364 8704 -9330
rect 8738 -9364 8760 -9330
rect 8688 -9391 8760 -9364
rect 8790 -9330 8844 -9307
rect 8790 -9364 8801 -9330
rect 8835 -9364 8844 -9330
rect 8790 -9391 8844 -9364
rect 8688 -9437 8738 -9391
rect 8990 -9345 9042 -9307
rect 8990 -9379 8998 -9345
rect 9032 -9379 9042 -9345
rect 8990 -9417 9042 -9379
rect 9252 -9345 9304 -9307
rect 9252 -9379 9262 -9345
rect 9296 -9379 9304 -9345
rect 9252 -9417 9304 -9379
rect 9450 -9338 9502 -9307
rect 9450 -9372 9458 -9338
rect 9492 -9372 9502 -9338
rect 9450 -9417 9502 -9372
rect 10080 -9338 10132 -9307
rect 10080 -9372 10090 -9338
rect 10124 -9372 10132 -9338
rect 10080 -9417 10132 -9372
rect 10370 -9345 10422 -9307
rect 10370 -9379 10378 -9345
rect 10412 -9379 10422 -9345
rect 10370 -9417 10422 -9379
rect 10632 -9345 10684 -9307
rect 10632 -9379 10642 -9345
rect 10676 -9379 10684 -9345
rect 10632 -9417 10684 -9379
rect 10738 -9330 10809 -9307
rect 10738 -9364 10761 -9330
rect 10795 -9364 10809 -9330
rect 10738 -9391 10809 -9364
rect 10839 -9330 10904 -9307
rect 10839 -9364 10859 -9330
rect 10893 -9364 10904 -9330
rect 10839 -9391 10904 -9364
rect 10854 -9437 10904 -9391
rect 11004 -9330 11057 -9307
rect 11004 -9364 11015 -9330
rect 11049 -9364 11057 -9330
rect 11004 -9437 11057 -9364
rect 11112 -9330 11164 -9307
rect 11112 -9364 11120 -9330
rect 11154 -9364 11164 -9330
rect 11112 -9437 11164 -9364
rect 11264 -9330 11336 -9307
rect 11264 -9364 11280 -9330
rect 11314 -9364 11336 -9330
rect 11264 -9391 11336 -9364
rect 11366 -9330 11420 -9307
rect 11366 -9364 11377 -9330
rect 11411 -9364 11420 -9330
rect 11366 -9391 11420 -9364
rect 11264 -9437 11314 -9391
rect 11658 -9345 11710 -9307
rect 11658 -9379 11666 -9345
rect 11700 -9379 11710 -9345
rect 11658 -9417 11710 -9379
rect 11920 -9345 11972 -9307
rect 13682 -9319 13735 -9307
rect 11920 -9379 11930 -9345
rect 11964 -9379 11972 -9345
rect 11920 -9417 11972 -9379
rect 13682 -9353 13690 -9319
rect 13724 -9353 13735 -9319
rect 13682 -9391 13735 -9353
rect 13765 -9332 13821 -9307
rect 13765 -9366 13776 -9332
rect 13810 -9366 13821 -9332
rect 13765 -9391 13821 -9366
rect 13851 -9332 13907 -9307
rect 13851 -9366 13862 -9332
rect 13896 -9366 13907 -9332
rect 13851 -9391 13907 -9366
rect 13937 -9332 13993 -9307
rect 13937 -9366 13948 -9332
rect 13982 -9366 13993 -9332
rect 13937 -9391 13993 -9366
rect 14023 -9332 14079 -9307
rect 14023 -9366 14034 -9332
rect 14068 -9366 14079 -9332
rect 14023 -9391 14079 -9366
rect 14109 -9332 14165 -9307
rect 14109 -9366 14120 -9332
rect 14154 -9366 14165 -9332
rect 14109 -9391 14165 -9366
rect 14195 -9323 14251 -9307
rect 14195 -9357 14206 -9323
rect 14240 -9357 14251 -9323
rect 14195 -9391 14251 -9357
rect 14281 -9332 14337 -9307
rect 14281 -9366 14292 -9332
rect 14326 -9366 14337 -9332
rect 14281 -9391 14337 -9366
rect 14367 -9323 14423 -9307
rect 14367 -9357 14378 -9323
rect 14412 -9357 14423 -9323
rect 14367 -9391 14423 -9357
rect 14453 -9332 14509 -9307
rect 14453 -9366 14464 -9332
rect 14498 -9366 14509 -9332
rect 14453 -9391 14509 -9366
rect 14539 -9323 14595 -9307
rect 14539 -9357 14550 -9323
rect 14584 -9357 14595 -9323
rect 14539 -9391 14595 -9357
rect 14625 -9332 14681 -9307
rect 14625 -9366 14636 -9332
rect 14670 -9366 14681 -9332
rect 14625 -9391 14681 -9366
rect 14711 -9323 14766 -9307
rect 14711 -9357 14722 -9323
rect 14756 -9357 14766 -9323
rect 14711 -9391 14766 -9357
rect 14796 -9332 14852 -9307
rect 14796 -9366 14807 -9332
rect 14841 -9366 14852 -9332
rect 14796 -9391 14852 -9366
rect 14882 -9323 14938 -9307
rect 14882 -9357 14893 -9323
rect 14927 -9357 14938 -9323
rect 14882 -9391 14938 -9357
rect 14968 -9332 15024 -9307
rect 14968 -9366 14979 -9332
rect 15013 -9366 15024 -9332
rect 14968 -9391 15024 -9366
rect 15054 -9323 15110 -9307
rect 15054 -9357 15065 -9323
rect 15099 -9357 15110 -9323
rect 15054 -9391 15110 -9357
rect 15140 -9332 15196 -9307
rect 15140 -9366 15151 -9332
rect 15185 -9366 15196 -9332
rect 15140 -9391 15196 -9366
rect 15226 -9323 15282 -9307
rect 15226 -9357 15237 -9323
rect 15271 -9357 15282 -9323
rect 15226 -9391 15282 -9357
rect 15312 -9332 15368 -9307
rect 15312 -9366 15323 -9332
rect 15357 -9366 15368 -9332
rect 15312 -9391 15368 -9366
rect 15398 -9323 15451 -9307
rect 15398 -9357 15409 -9323
rect 15443 -9357 15451 -9323
rect 15398 -9391 15451 -9357
rect 15614 -9338 15666 -9307
rect 15614 -9372 15622 -9338
rect 15656 -9372 15666 -9338
rect 15614 -9417 15666 -9372
rect 16612 -9338 16664 -9307
rect 16612 -9372 16622 -9338
rect 16656 -9372 16664 -9338
rect 16612 -9417 16664 -9372
rect -2970 -10236 -2918 -10191
rect -2970 -10270 -2962 -10236
rect -2928 -10270 -2918 -10236
rect -2970 -10301 -2918 -10270
rect -2340 -10236 -2288 -10191
rect -2340 -10270 -2330 -10236
rect -2296 -10270 -2288 -10236
rect -2340 -10301 -2288 -10270
rect -1590 -10236 -1538 -10191
rect -1590 -10270 -1582 -10236
rect -1548 -10270 -1538 -10236
rect -1590 -10301 -1538 -10270
rect -960 -10236 -908 -10191
rect -960 -10270 -950 -10236
rect -916 -10270 -908 -10236
rect -960 -10301 -908 -10270
rect -854 -10236 -802 -10191
rect -854 -10270 -846 -10236
rect -812 -10270 -802 -10236
rect -854 -10301 -802 -10270
rect -224 -10236 -172 -10191
rect -224 -10270 -214 -10236
rect -180 -10270 -172 -10236
rect -224 -10301 -172 -10270
rect -26 -10229 26 -10191
rect -26 -10263 -18 -10229
rect 16 -10263 26 -10229
rect -26 -10301 26 -10263
rect 236 -10229 288 -10191
rect 236 -10263 246 -10229
rect 280 -10263 288 -10229
rect 236 -10301 288 -10263
rect 540 -10217 590 -10171
rect 434 -10244 488 -10217
rect 434 -10278 443 -10244
rect 477 -10278 488 -10244
rect 434 -10301 488 -10278
rect 518 -10244 590 -10217
rect 518 -10278 540 -10244
rect 574 -10278 590 -10244
rect 518 -10301 590 -10278
rect 690 -10244 742 -10171
rect 690 -10278 700 -10244
rect 734 -10278 742 -10244
rect 690 -10301 742 -10278
rect 797 -10244 850 -10171
rect 797 -10278 805 -10244
rect 839 -10278 850 -10244
rect 797 -10301 850 -10278
rect 950 -10217 1000 -10171
rect 950 -10244 1015 -10217
rect 950 -10278 961 -10244
rect 995 -10278 1015 -10244
rect 950 -10301 1015 -10278
rect 1045 -10244 1116 -10217
rect 1045 -10278 1059 -10244
rect 1093 -10278 1116 -10244
rect 1045 -10301 1116 -10278
rect 1262 -10229 1314 -10191
rect 1262 -10263 1270 -10229
rect 1304 -10263 1314 -10229
rect 1262 -10301 1314 -10263
rect 1524 -10229 1576 -10191
rect 1524 -10263 1534 -10229
rect 1568 -10263 1576 -10229
rect 1524 -10301 1576 -10263
rect 1722 -10236 1774 -10191
rect 1722 -10270 1730 -10236
rect 1764 -10270 1774 -10236
rect 1722 -10301 1774 -10270
rect 2352 -10236 2404 -10191
rect 2352 -10270 2362 -10236
rect 2396 -10270 2404 -10236
rect 2352 -10301 2404 -10270
rect 2550 -10229 2602 -10191
rect 2550 -10263 2558 -10229
rect 2592 -10263 2602 -10229
rect 2550 -10301 2602 -10263
rect 2812 -10229 2864 -10191
rect 2812 -10263 2822 -10229
rect 2856 -10263 2864 -10229
rect 2812 -10301 2864 -10263
rect 3116 -10217 3166 -10171
rect 3010 -10244 3064 -10217
rect 3010 -10278 3019 -10244
rect 3053 -10278 3064 -10244
rect 3010 -10301 3064 -10278
rect 3094 -10244 3166 -10217
rect 3094 -10278 3116 -10244
rect 3150 -10278 3166 -10244
rect 3094 -10301 3166 -10278
rect 3266 -10244 3318 -10171
rect 3266 -10278 3276 -10244
rect 3310 -10278 3318 -10244
rect 3266 -10301 3318 -10278
rect 3373 -10244 3426 -10171
rect 3373 -10278 3381 -10244
rect 3415 -10278 3426 -10244
rect 3373 -10301 3426 -10278
rect 3526 -10217 3576 -10171
rect 3526 -10244 3591 -10217
rect 3526 -10278 3537 -10244
rect 3571 -10278 3591 -10244
rect 3526 -10301 3591 -10278
rect 3621 -10244 3692 -10217
rect 3621 -10278 3635 -10244
rect 3669 -10278 3692 -10244
rect 3621 -10301 3692 -10278
rect 3838 -10229 3890 -10191
rect 3838 -10263 3846 -10229
rect 3880 -10263 3890 -10229
rect 3838 -10301 3890 -10263
rect 4100 -10229 4152 -10191
rect 4100 -10263 4110 -10229
rect 4144 -10263 4152 -10229
rect 4100 -10301 4152 -10263
rect 4298 -10236 4350 -10191
rect 4298 -10270 4306 -10236
rect 4340 -10270 4350 -10236
rect 4298 -10301 4350 -10270
rect 4928 -10236 4980 -10191
rect 4928 -10270 4938 -10236
rect 4972 -10270 4980 -10236
rect 4928 -10301 4980 -10270
rect 5126 -10229 5178 -10191
rect 5126 -10263 5134 -10229
rect 5168 -10263 5178 -10229
rect 5126 -10301 5178 -10263
rect 5388 -10229 5440 -10191
rect 5388 -10263 5398 -10229
rect 5432 -10263 5440 -10229
rect 5388 -10301 5440 -10263
rect 5692 -10217 5742 -10171
rect 5586 -10244 5640 -10217
rect 5586 -10278 5595 -10244
rect 5629 -10278 5640 -10244
rect 5586 -10301 5640 -10278
rect 5670 -10244 5742 -10217
rect 5670 -10278 5692 -10244
rect 5726 -10278 5742 -10244
rect 5670 -10301 5742 -10278
rect 5842 -10244 5894 -10171
rect 5842 -10278 5852 -10244
rect 5886 -10278 5894 -10244
rect 5842 -10301 5894 -10278
rect 5949 -10244 6002 -10171
rect 5949 -10278 5957 -10244
rect 5991 -10278 6002 -10244
rect 5949 -10301 6002 -10278
rect 6102 -10217 6152 -10171
rect 6102 -10244 6167 -10217
rect 6102 -10278 6113 -10244
rect 6147 -10278 6167 -10244
rect 6102 -10301 6167 -10278
rect 6197 -10244 6268 -10217
rect 6197 -10278 6211 -10244
rect 6245 -10278 6268 -10244
rect 6197 -10301 6268 -10278
rect 6414 -10229 6466 -10191
rect 6414 -10263 6422 -10229
rect 6456 -10263 6466 -10229
rect 6414 -10301 6466 -10263
rect 6676 -10229 6728 -10191
rect 6676 -10263 6686 -10229
rect 6720 -10263 6728 -10229
rect 6676 -10301 6728 -10263
rect 6874 -10236 6926 -10191
rect 6874 -10270 6882 -10236
rect 6916 -10270 6926 -10236
rect 6874 -10301 6926 -10270
rect 7504 -10236 7556 -10191
rect 7504 -10270 7514 -10236
rect 7548 -10270 7556 -10236
rect 7504 -10301 7556 -10270
rect 7702 -10229 7754 -10191
rect 7702 -10263 7710 -10229
rect 7744 -10263 7754 -10229
rect 7702 -10301 7754 -10263
rect 7964 -10229 8016 -10191
rect 7964 -10263 7974 -10229
rect 8008 -10263 8016 -10229
rect 7964 -10301 8016 -10263
rect 8268 -10217 8318 -10171
rect 8162 -10244 8216 -10217
rect 8162 -10278 8171 -10244
rect 8205 -10278 8216 -10244
rect 8162 -10301 8216 -10278
rect 8246 -10244 8318 -10217
rect 8246 -10278 8268 -10244
rect 8302 -10278 8318 -10244
rect 8246 -10301 8318 -10278
rect 8418 -10244 8470 -10171
rect 8418 -10278 8428 -10244
rect 8462 -10278 8470 -10244
rect 8418 -10301 8470 -10278
rect 8525 -10244 8578 -10171
rect 8525 -10278 8533 -10244
rect 8567 -10278 8578 -10244
rect 8525 -10301 8578 -10278
rect 8678 -10217 8728 -10171
rect 8678 -10244 8743 -10217
rect 8678 -10278 8689 -10244
rect 8723 -10278 8743 -10244
rect 8678 -10301 8743 -10278
rect 8773 -10244 8844 -10217
rect 8773 -10278 8787 -10244
rect 8821 -10278 8844 -10244
rect 8773 -10301 8844 -10278
rect 8990 -10229 9042 -10191
rect 8990 -10263 8998 -10229
rect 9032 -10263 9042 -10229
rect 8990 -10301 9042 -10263
rect 9252 -10229 9304 -10191
rect 9252 -10263 9262 -10229
rect 9296 -10263 9304 -10229
rect 9252 -10301 9304 -10263
rect 9450 -10236 9502 -10191
rect 9450 -10270 9458 -10236
rect 9492 -10270 9502 -10236
rect 9450 -10301 9502 -10270
rect 10080 -10236 10132 -10191
rect 10080 -10270 10090 -10236
rect 10124 -10270 10132 -10236
rect 10080 -10301 10132 -10270
rect 10370 -10229 10422 -10191
rect 10370 -10263 10378 -10229
rect 10412 -10263 10422 -10229
rect 10370 -10301 10422 -10263
rect 10632 -10229 10684 -10191
rect 10844 -10217 10894 -10171
rect 10632 -10263 10642 -10229
rect 10676 -10263 10684 -10229
rect 10632 -10301 10684 -10263
rect 10738 -10244 10792 -10217
rect 10738 -10278 10747 -10244
rect 10781 -10278 10792 -10244
rect 10738 -10301 10792 -10278
rect 10822 -10244 10894 -10217
rect 10822 -10278 10844 -10244
rect 10878 -10278 10894 -10244
rect 10822 -10301 10894 -10278
rect 10994 -10244 11046 -10171
rect 10994 -10278 11004 -10244
rect 11038 -10278 11046 -10244
rect 10994 -10301 11046 -10278
rect 11101 -10244 11154 -10171
rect 11101 -10278 11109 -10244
rect 11143 -10278 11154 -10244
rect 11101 -10301 11154 -10278
rect 11254 -10217 11304 -10171
rect 11254 -10244 11319 -10217
rect 11254 -10278 11265 -10244
rect 11299 -10278 11319 -10244
rect 11254 -10301 11319 -10278
rect 11349 -10244 11420 -10217
rect 11349 -10278 11363 -10244
rect 11397 -10278 11420 -10244
rect 11349 -10301 11420 -10278
rect 11658 -10229 11710 -10191
rect 11658 -10263 11666 -10229
rect 11700 -10263 11710 -10229
rect 11658 -10301 11710 -10263
rect 11920 -10229 11972 -10191
rect 11920 -10263 11930 -10229
rect 11964 -10263 11972 -10229
rect 11920 -10301 11972 -10263
rect 12567 -10253 12633 -10217
rect 12567 -10287 12588 -10253
rect 12622 -10287 12633 -10253
rect 12567 -10301 12633 -10287
rect 12663 -10242 12719 -10217
rect 12663 -10276 12674 -10242
rect 12708 -10276 12719 -10242
rect 12663 -10301 12719 -10276
rect 12749 -10253 12805 -10217
rect 12749 -10287 12760 -10253
rect 12794 -10287 12805 -10253
rect 12749 -10301 12805 -10287
rect 12835 -10242 12891 -10217
rect 12835 -10276 12846 -10242
rect 12880 -10276 12891 -10242
rect 12835 -10301 12891 -10276
rect 12921 -10253 13000 -10217
rect 12921 -10287 12932 -10253
rect 12966 -10287 13000 -10253
rect 13222 -10229 13274 -10191
rect 13222 -10263 13230 -10229
rect 13264 -10263 13274 -10229
rect 12921 -10301 13000 -10287
rect 13222 -10301 13274 -10263
rect 13484 -10229 13536 -10191
rect 13484 -10263 13494 -10229
rect 13528 -10263 13536 -10229
rect 13484 -10301 13536 -10263
rect 13682 -10255 13735 -10217
rect 13682 -10289 13690 -10255
rect 13724 -10289 13735 -10255
rect 13682 -10301 13735 -10289
rect 13765 -10242 13821 -10217
rect 13765 -10276 13776 -10242
rect 13810 -10276 13821 -10242
rect 13765 -10301 13821 -10276
rect 13851 -10242 13907 -10217
rect 13851 -10276 13862 -10242
rect 13896 -10276 13907 -10242
rect 13851 -10301 13907 -10276
rect 13937 -10242 13993 -10217
rect 13937 -10276 13948 -10242
rect 13982 -10276 13993 -10242
rect 13937 -10301 13993 -10276
rect 14023 -10242 14079 -10217
rect 14023 -10276 14034 -10242
rect 14068 -10276 14079 -10242
rect 14023 -10301 14079 -10276
rect 14109 -10242 14165 -10217
rect 14109 -10276 14120 -10242
rect 14154 -10276 14165 -10242
rect 14109 -10301 14165 -10276
rect 14195 -10251 14251 -10217
rect 14195 -10285 14206 -10251
rect 14240 -10285 14251 -10251
rect 14195 -10301 14251 -10285
rect 14281 -10242 14337 -10217
rect 14281 -10276 14292 -10242
rect 14326 -10276 14337 -10242
rect 14281 -10301 14337 -10276
rect 14367 -10251 14423 -10217
rect 14367 -10285 14378 -10251
rect 14412 -10285 14423 -10251
rect 14367 -10301 14423 -10285
rect 14453 -10242 14509 -10217
rect 14453 -10276 14464 -10242
rect 14498 -10276 14509 -10242
rect 14453 -10301 14509 -10276
rect 14539 -10251 14595 -10217
rect 14539 -10285 14550 -10251
rect 14584 -10285 14595 -10251
rect 14539 -10301 14595 -10285
rect 14625 -10242 14681 -10217
rect 14625 -10276 14636 -10242
rect 14670 -10276 14681 -10242
rect 14625 -10301 14681 -10276
rect 14711 -10251 14766 -10217
rect 14711 -10285 14722 -10251
rect 14756 -10285 14766 -10251
rect 14711 -10301 14766 -10285
rect 14796 -10242 14852 -10217
rect 14796 -10276 14807 -10242
rect 14841 -10276 14852 -10242
rect 14796 -10301 14852 -10276
rect 14882 -10251 14938 -10217
rect 14882 -10285 14893 -10251
rect 14927 -10285 14938 -10251
rect 14882 -10301 14938 -10285
rect 14968 -10242 15024 -10217
rect 14968 -10276 14979 -10242
rect 15013 -10276 15024 -10242
rect 14968 -10301 15024 -10276
rect 15054 -10251 15110 -10217
rect 15054 -10285 15065 -10251
rect 15099 -10285 15110 -10251
rect 15054 -10301 15110 -10285
rect 15140 -10242 15196 -10217
rect 15140 -10276 15151 -10242
rect 15185 -10276 15196 -10242
rect 15140 -10301 15196 -10276
rect 15226 -10251 15282 -10217
rect 15226 -10285 15237 -10251
rect 15271 -10285 15282 -10251
rect 15226 -10301 15282 -10285
rect 15312 -10242 15368 -10217
rect 15312 -10276 15323 -10242
rect 15357 -10276 15368 -10242
rect 15312 -10301 15368 -10276
rect 15398 -10251 15451 -10217
rect 15398 -10285 15409 -10251
rect 15443 -10285 15451 -10251
rect 15614 -10236 15666 -10191
rect 15614 -10270 15622 -10236
rect 15656 -10270 15666 -10236
rect 15398 -10301 15451 -10285
rect 15614 -10301 15666 -10270
rect 16612 -10236 16664 -10191
rect 16612 -10270 16622 -10236
rect 16656 -10270 16664 -10236
rect 16612 -10301 16664 -10270
rect -2970 -10426 -2918 -10395
rect -2970 -10460 -2962 -10426
rect -2928 -10460 -2918 -10426
rect -2970 -10505 -2918 -10460
rect -2340 -10426 -2288 -10395
rect -2340 -10460 -2330 -10426
rect -2296 -10460 -2288 -10426
rect -2340 -10505 -2288 -10460
rect -1875 -10418 -1823 -10395
rect -1875 -10452 -1867 -10418
rect -1833 -10452 -1823 -10418
rect -1875 -10479 -1823 -10452
rect -1793 -10416 -1736 -10395
rect -1793 -10450 -1783 -10416
rect -1749 -10450 -1736 -10416
rect -1793 -10479 -1736 -10450
rect -1590 -10426 -1538 -10395
rect -1590 -10460 -1582 -10426
rect -1548 -10460 -1538 -10426
rect -1590 -10505 -1538 -10460
rect -960 -10426 -908 -10395
rect -960 -10460 -950 -10426
rect -916 -10460 -908 -10426
rect -960 -10505 -908 -10460
rect -854 -10426 -802 -10395
rect -854 -10460 -846 -10426
rect -812 -10460 -802 -10426
rect -854 -10505 -802 -10460
rect -224 -10426 -172 -10395
rect -224 -10460 -214 -10426
rect -180 -10460 -172 -10426
rect -224 -10505 -172 -10460
rect -26 -10433 26 -10395
rect -26 -10467 -18 -10433
rect 16 -10467 26 -10433
rect -26 -10505 26 -10467
rect 236 -10433 288 -10395
rect 236 -10467 246 -10433
rect 280 -10467 288 -10433
rect 236 -10505 288 -10467
rect 434 -10418 505 -10395
rect 434 -10452 457 -10418
rect 491 -10452 505 -10418
rect 434 -10479 505 -10452
rect 535 -10418 600 -10395
rect 535 -10452 555 -10418
rect 589 -10452 600 -10418
rect 535 -10479 600 -10452
rect 550 -10525 600 -10479
rect 700 -10418 753 -10395
rect 700 -10452 711 -10418
rect 745 -10452 753 -10418
rect 700 -10525 753 -10452
rect 808 -10418 860 -10395
rect 808 -10452 816 -10418
rect 850 -10452 860 -10418
rect 808 -10525 860 -10452
rect 960 -10418 1032 -10395
rect 960 -10452 976 -10418
rect 1010 -10452 1032 -10418
rect 960 -10479 1032 -10452
rect 1062 -10418 1116 -10395
rect 1062 -10452 1073 -10418
rect 1107 -10452 1116 -10418
rect 1062 -10479 1116 -10452
rect 960 -10525 1010 -10479
rect 1262 -10433 1314 -10395
rect 1262 -10467 1270 -10433
rect 1304 -10467 1314 -10433
rect 1262 -10505 1314 -10467
rect 1524 -10433 1576 -10395
rect 1524 -10467 1534 -10433
rect 1568 -10467 1576 -10433
rect 1524 -10505 1576 -10467
rect 1722 -10426 1774 -10395
rect 1722 -10460 1730 -10426
rect 1764 -10460 1774 -10426
rect 1722 -10505 1774 -10460
rect 2352 -10426 2404 -10395
rect 2352 -10460 2362 -10426
rect 2396 -10460 2404 -10426
rect 2352 -10505 2404 -10460
rect 2550 -10433 2602 -10395
rect 2550 -10467 2558 -10433
rect 2592 -10467 2602 -10433
rect 2550 -10505 2602 -10467
rect 2812 -10433 2864 -10395
rect 2812 -10467 2822 -10433
rect 2856 -10467 2864 -10433
rect 2812 -10505 2864 -10467
rect 3010 -10418 3081 -10395
rect 3010 -10452 3033 -10418
rect 3067 -10452 3081 -10418
rect 3010 -10479 3081 -10452
rect 3111 -10418 3176 -10395
rect 3111 -10452 3131 -10418
rect 3165 -10452 3176 -10418
rect 3111 -10479 3176 -10452
rect 3126 -10525 3176 -10479
rect 3276 -10418 3329 -10395
rect 3276 -10452 3287 -10418
rect 3321 -10452 3329 -10418
rect 3276 -10525 3329 -10452
rect 3384 -10418 3436 -10395
rect 3384 -10452 3392 -10418
rect 3426 -10452 3436 -10418
rect 3384 -10525 3436 -10452
rect 3536 -10418 3608 -10395
rect 3536 -10452 3552 -10418
rect 3586 -10452 3608 -10418
rect 3536 -10479 3608 -10452
rect 3638 -10418 3692 -10395
rect 3638 -10452 3649 -10418
rect 3683 -10452 3692 -10418
rect 3638 -10479 3692 -10452
rect 3536 -10525 3586 -10479
rect 3838 -10433 3890 -10395
rect 3838 -10467 3846 -10433
rect 3880 -10467 3890 -10433
rect 3838 -10505 3890 -10467
rect 4100 -10433 4152 -10395
rect 4100 -10467 4110 -10433
rect 4144 -10467 4152 -10433
rect 4100 -10505 4152 -10467
rect 4298 -10426 4350 -10395
rect 4298 -10460 4306 -10426
rect 4340 -10460 4350 -10426
rect 4298 -10505 4350 -10460
rect 4928 -10426 4980 -10395
rect 4928 -10460 4938 -10426
rect 4972 -10460 4980 -10426
rect 4928 -10505 4980 -10460
rect 5126 -10433 5178 -10395
rect 5126 -10467 5134 -10433
rect 5168 -10467 5178 -10433
rect 5126 -10505 5178 -10467
rect 5388 -10433 5440 -10395
rect 5388 -10467 5398 -10433
rect 5432 -10467 5440 -10433
rect 5388 -10505 5440 -10467
rect 5586 -10418 5657 -10395
rect 5586 -10452 5609 -10418
rect 5643 -10452 5657 -10418
rect 5586 -10479 5657 -10452
rect 5687 -10418 5752 -10395
rect 5687 -10452 5707 -10418
rect 5741 -10452 5752 -10418
rect 5687 -10479 5752 -10452
rect 5702 -10525 5752 -10479
rect 5852 -10418 5905 -10395
rect 5852 -10452 5863 -10418
rect 5897 -10452 5905 -10418
rect 5852 -10525 5905 -10452
rect 5960 -10418 6012 -10395
rect 5960 -10452 5968 -10418
rect 6002 -10452 6012 -10418
rect 5960 -10525 6012 -10452
rect 6112 -10418 6184 -10395
rect 6112 -10452 6128 -10418
rect 6162 -10452 6184 -10418
rect 6112 -10479 6184 -10452
rect 6214 -10418 6268 -10395
rect 6214 -10452 6225 -10418
rect 6259 -10452 6268 -10418
rect 6214 -10479 6268 -10452
rect 6112 -10525 6162 -10479
rect 6414 -10433 6466 -10395
rect 6414 -10467 6422 -10433
rect 6456 -10467 6466 -10433
rect 6414 -10505 6466 -10467
rect 6676 -10433 6728 -10395
rect 6676 -10467 6686 -10433
rect 6720 -10467 6728 -10433
rect 6676 -10505 6728 -10467
rect 6874 -10426 6926 -10395
rect 6874 -10460 6882 -10426
rect 6916 -10460 6926 -10426
rect 6874 -10505 6926 -10460
rect 7504 -10426 7556 -10395
rect 7504 -10460 7514 -10426
rect 7548 -10460 7556 -10426
rect 7504 -10505 7556 -10460
rect 7702 -10433 7754 -10395
rect 7702 -10467 7710 -10433
rect 7744 -10467 7754 -10433
rect 7702 -10505 7754 -10467
rect 7964 -10433 8016 -10395
rect 7964 -10467 7974 -10433
rect 8008 -10467 8016 -10433
rect 7964 -10505 8016 -10467
rect 8162 -10418 8233 -10395
rect 8162 -10452 8185 -10418
rect 8219 -10452 8233 -10418
rect 8162 -10479 8233 -10452
rect 8263 -10418 8328 -10395
rect 8263 -10452 8283 -10418
rect 8317 -10452 8328 -10418
rect 8263 -10479 8328 -10452
rect 8278 -10525 8328 -10479
rect 8428 -10418 8481 -10395
rect 8428 -10452 8439 -10418
rect 8473 -10452 8481 -10418
rect 8428 -10525 8481 -10452
rect 8536 -10418 8588 -10395
rect 8536 -10452 8544 -10418
rect 8578 -10452 8588 -10418
rect 8536 -10525 8588 -10452
rect 8688 -10418 8760 -10395
rect 8688 -10452 8704 -10418
rect 8738 -10452 8760 -10418
rect 8688 -10479 8760 -10452
rect 8790 -10418 8844 -10395
rect 8790 -10452 8801 -10418
rect 8835 -10452 8844 -10418
rect 8790 -10479 8844 -10452
rect 8688 -10525 8738 -10479
rect 8990 -10433 9042 -10395
rect 8990 -10467 8998 -10433
rect 9032 -10467 9042 -10433
rect 8990 -10505 9042 -10467
rect 9252 -10433 9304 -10395
rect 9252 -10467 9262 -10433
rect 9296 -10467 9304 -10433
rect 9252 -10505 9304 -10467
rect 9450 -10426 9502 -10395
rect 9450 -10460 9458 -10426
rect 9492 -10460 9502 -10426
rect 9450 -10505 9502 -10460
rect 10080 -10426 10132 -10395
rect 10080 -10460 10090 -10426
rect 10124 -10460 10132 -10426
rect 10080 -10505 10132 -10460
rect 10370 -10433 10422 -10395
rect 10370 -10467 10378 -10433
rect 10412 -10467 10422 -10433
rect 10370 -10505 10422 -10467
rect 10632 -10433 10684 -10395
rect 10632 -10467 10642 -10433
rect 10676 -10467 10684 -10433
rect 10632 -10505 10684 -10467
rect 10738 -10418 10809 -10395
rect 10738 -10452 10761 -10418
rect 10795 -10452 10809 -10418
rect 10738 -10479 10809 -10452
rect 10839 -10418 10904 -10395
rect 10839 -10452 10859 -10418
rect 10893 -10452 10904 -10418
rect 10839 -10479 10904 -10452
rect 10854 -10525 10904 -10479
rect 11004 -10418 11057 -10395
rect 11004 -10452 11015 -10418
rect 11049 -10452 11057 -10418
rect 11004 -10525 11057 -10452
rect 11112 -10418 11164 -10395
rect 11112 -10452 11120 -10418
rect 11154 -10452 11164 -10418
rect 11112 -10525 11164 -10452
rect 11264 -10418 11336 -10395
rect 11264 -10452 11280 -10418
rect 11314 -10452 11336 -10418
rect 11264 -10479 11336 -10452
rect 11366 -10418 11420 -10395
rect 11366 -10452 11377 -10418
rect 11411 -10452 11420 -10418
rect 11366 -10479 11420 -10452
rect 11264 -10525 11314 -10479
rect 11658 -10433 11710 -10395
rect 11658 -10467 11666 -10433
rect 11700 -10467 11710 -10433
rect 11658 -10505 11710 -10467
rect 11920 -10433 11972 -10395
rect 11920 -10467 11930 -10433
rect 11964 -10467 11972 -10433
rect 11920 -10505 11972 -10467
rect 13590 -10426 13642 -10395
rect 13590 -10460 13598 -10426
rect 13632 -10460 13642 -10426
rect 13590 -10505 13642 -10460
rect 14588 -10426 14640 -10395
rect 14588 -10460 14598 -10426
rect 14632 -10460 14640 -10426
rect 14588 -10505 14640 -10460
rect 14786 -10426 14838 -10395
rect 14786 -10460 14794 -10426
rect 14828 -10460 14838 -10426
rect 14786 -10505 14838 -10460
rect 15784 -10426 15836 -10395
rect 15784 -10460 15794 -10426
rect 15828 -10460 15836 -10426
rect 15784 -10505 15836 -10460
rect 15982 -10426 16034 -10395
rect 15982 -10460 15990 -10426
rect 16024 -10460 16034 -10426
rect 15982 -10505 16034 -10460
rect 16612 -10426 16664 -10395
rect 16612 -10460 16622 -10426
rect 16656 -10460 16664 -10426
rect 16612 -10505 16664 -10460
rect -2970 -11324 -2918 -11279
rect -2970 -11358 -2962 -11324
rect -2928 -11358 -2918 -11324
rect -2970 -11389 -2918 -11358
rect -2340 -11324 -2288 -11279
rect -2340 -11358 -2330 -11324
rect -2296 -11358 -2288 -11324
rect -2340 -11389 -2288 -11358
rect -1590 -11324 -1538 -11279
rect -1590 -11358 -1582 -11324
rect -1548 -11358 -1538 -11324
rect -1590 -11389 -1538 -11358
rect -960 -11324 -908 -11279
rect -960 -11358 -950 -11324
rect -916 -11358 -908 -11324
rect -960 -11389 -908 -11358
rect -854 -11324 -802 -11279
rect -854 -11358 -846 -11324
rect -812 -11358 -802 -11324
rect -854 -11389 -802 -11358
rect -224 -11324 -172 -11279
rect -224 -11358 -214 -11324
rect -180 -11358 -172 -11324
rect -224 -11389 -172 -11358
rect -26 -11317 26 -11279
rect -26 -11351 -18 -11317
rect 16 -11351 26 -11317
rect -26 -11389 26 -11351
rect 236 -11317 288 -11279
rect 236 -11351 246 -11317
rect 280 -11351 288 -11317
rect 236 -11389 288 -11351
rect 550 -11305 600 -11259
rect 434 -11332 505 -11305
rect 434 -11366 457 -11332
rect 491 -11366 505 -11332
rect 434 -11389 505 -11366
rect 535 -11332 600 -11305
rect 535 -11366 555 -11332
rect 589 -11366 600 -11332
rect 535 -11389 600 -11366
rect 700 -11332 753 -11259
rect 700 -11366 711 -11332
rect 745 -11366 753 -11332
rect 700 -11389 753 -11366
rect 808 -11332 860 -11259
rect 808 -11366 816 -11332
rect 850 -11366 860 -11332
rect 808 -11389 860 -11366
rect 960 -11305 1010 -11259
rect 960 -11332 1032 -11305
rect 960 -11366 976 -11332
rect 1010 -11366 1032 -11332
rect 960 -11389 1032 -11366
rect 1062 -11332 1116 -11305
rect 1062 -11366 1073 -11332
rect 1107 -11366 1116 -11332
rect 1062 -11389 1116 -11366
rect 1262 -11317 1314 -11279
rect 1262 -11351 1270 -11317
rect 1304 -11351 1314 -11317
rect 1262 -11389 1314 -11351
rect 1524 -11317 1576 -11279
rect 1524 -11351 1534 -11317
rect 1568 -11351 1576 -11317
rect 1524 -11389 1576 -11351
rect 1722 -11324 1774 -11279
rect 1722 -11358 1730 -11324
rect 1764 -11358 1774 -11324
rect 1722 -11389 1774 -11358
rect 2352 -11324 2404 -11279
rect 2352 -11358 2362 -11324
rect 2396 -11358 2404 -11324
rect 2352 -11389 2404 -11358
rect 2550 -11317 2602 -11279
rect 2550 -11351 2558 -11317
rect 2592 -11351 2602 -11317
rect 2550 -11389 2602 -11351
rect 2812 -11317 2864 -11279
rect 2812 -11351 2822 -11317
rect 2856 -11351 2864 -11317
rect 2812 -11389 2864 -11351
rect 3126 -11305 3176 -11259
rect 3010 -11332 3081 -11305
rect 3010 -11366 3033 -11332
rect 3067 -11366 3081 -11332
rect 3010 -11389 3081 -11366
rect 3111 -11332 3176 -11305
rect 3111 -11366 3131 -11332
rect 3165 -11366 3176 -11332
rect 3111 -11389 3176 -11366
rect 3276 -11332 3329 -11259
rect 3276 -11366 3287 -11332
rect 3321 -11366 3329 -11332
rect 3276 -11389 3329 -11366
rect 3384 -11332 3436 -11259
rect 3384 -11366 3392 -11332
rect 3426 -11366 3436 -11332
rect 3384 -11389 3436 -11366
rect 3536 -11305 3586 -11259
rect 3536 -11332 3608 -11305
rect 3536 -11366 3552 -11332
rect 3586 -11366 3608 -11332
rect 3536 -11389 3608 -11366
rect 3638 -11332 3692 -11305
rect 3638 -11366 3649 -11332
rect 3683 -11366 3692 -11332
rect 3638 -11389 3692 -11366
rect 3838 -11317 3890 -11279
rect 3838 -11351 3846 -11317
rect 3880 -11351 3890 -11317
rect 3838 -11389 3890 -11351
rect 4100 -11317 4152 -11279
rect 4100 -11351 4110 -11317
rect 4144 -11351 4152 -11317
rect 4100 -11389 4152 -11351
rect 4298 -11324 4350 -11279
rect 4298 -11358 4306 -11324
rect 4340 -11358 4350 -11324
rect 4298 -11389 4350 -11358
rect 4928 -11324 4980 -11279
rect 4928 -11358 4938 -11324
rect 4972 -11358 4980 -11324
rect 4928 -11389 4980 -11358
rect 5126 -11317 5178 -11279
rect 5126 -11351 5134 -11317
rect 5168 -11351 5178 -11317
rect 5126 -11389 5178 -11351
rect 5388 -11317 5440 -11279
rect 5388 -11351 5398 -11317
rect 5432 -11351 5440 -11317
rect 5388 -11389 5440 -11351
rect 5702 -11305 5752 -11259
rect 5586 -11332 5657 -11305
rect 5586 -11366 5609 -11332
rect 5643 -11366 5657 -11332
rect 5586 -11389 5657 -11366
rect 5687 -11332 5752 -11305
rect 5687 -11366 5707 -11332
rect 5741 -11366 5752 -11332
rect 5687 -11389 5752 -11366
rect 5852 -11332 5905 -11259
rect 5852 -11366 5863 -11332
rect 5897 -11366 5905 -11332
rect 5852 -11389 5905 -11366
rect 5960 -11332 6012 -11259
rect 5960 -11366 5968 -11332
rect 6002 -11366 6012 -11332
rect 5960 -11389 6012 -11366
rect 6112 -11305 6162 -11259
rect 6112 -11332 6184 -11305
rect 6112 -11366 6128 -11332
rect 6162 -11366 6184 -11332
rect 6112 -11389 6184 -11366
rect 6214 -11332 6268 -11305
rect 6214 -11366 6225 -11332
rect 6259 -11366 6268 -11332
rect 6214 -11389 6268 -11366
rect 6414 -11317 6466 -11279
rect 6414 -11351 6422 -11317
rect 6456 -11351 6466 -11317
rect 6414 -11389 6466 -11351
rect 6676 -11317 6728 -11279
rect 6676 -11351 6686 -11317
rect 6720 -11351 6728 -11317
rect 6676 -11389 6728 -11351
rect 6874 -11324 6926 -11279
rect 6874 -11358 6882 -11324
rect 6916 -11358 6926 -11324
rect 6874 -11389 6926 -11358
rect 7504 -11324 7556 -11279
rect 7504 -11358 7514 -11324
rect 7548 -11358 7556 -11324
rect 7504 -11389 7556 -11358
rect 7702 -11317 7754 -11279
rect 7702 -11351 7710 -11317
rect 7744 -11351 7754 -11317
rect 7702 -11389 7754 -11351
rect 7964 -11317 8016 -11279
rect 7964 -11351 7974 -11317
rect 8008 -11351 8016 -11317
rect 7964 -11389 8016 -11351
rect 8278 -11305 8328 -11259
rect 8162 -11332 8233 -11305
rect 8162 -11366 8185 -11332
rect 8219 -11366 8233 -11332
rect 8162 -11389 8233 -11366
rect 8263 -11332 8328 -11305
rect 8263 -11366 8283 -11332
rect 8317 -11366 8328 -11332
rect 8263 -11389 8328 -11366
rect 8428 -11332 8481 -11259
rect 8428 -11366 8439 -11332
rect 8473 -11366 8481 -11332
rect 8428 -11389 8481 -11366
rect 8536 -11332 8588 -11259
rect 8536 -11366 8544 -11332
rect 8578 -11366 8588 -11332
rect 8536 -11389 8588 -11366
rect 8688 -11305 8738 -11259
rect 8688 -11332 8760 -11305
rect 8688 -11366 8704 -11332
rect 8738 -11366 8760 -11332
rect 8688 -11389 8760 -11366
rect 8790 -11332 8844 -11305
rect 8790 -11366 8801 -11332
rect 8835 -11366 8844 -11332
rect 8790 -11389 8844 -11366
rect 8990 -11317 9042 -11279
rect 8990 -11351 8998 -11317
rect 9032 -11351 9042 -11317
rect 8990 -11389 9042 -11351
rect 9252 -11317 9304 -11279
rect 9252 -11351 9262 -11317
rect 9296 -11351 9304 -11317
rect 9252 -11389 9304 -11351
rect 9450 -11324 9502 -11279
rect 9450 -11358 9458 -11324
rect 9492 -11358 9502 -11324
rect 9450 -11389 9502 -11358
rect 10080 -11324 10132 -11279
rect 10080 -11358 10090 -11324
rect 10124 -11358 10132 -11324
rect 10080 -11389 10132 -11358
rect 10370 -11317 10422 -11279
rect 10370 -11351 10378 -11317
rect 10412 -11351 10422 -11317
rect 10370 -11389 10422 -11351
rect 10632 -11317 10684 -11279
rect 10854 -11305 10904 -11259
rect 10632 -11351 10642 -11317
rect 10676 -11351 10684 -11317
rect 10632 -11389 10684 -11351
rect 10738 -11332 10809 -11305
rect 10738 -11366 10761 -11332
rect 10795 -11366 10809 -11332
rect 10738 -11389 10809 -11366
rect 10839 -11332 10904 -11305
rect 10839 -11366 10859 -11332
rect 10893 -11366 10904 -11332
rect 10839 -11389 10904 -11366
rect 11004 -11332 11057 -11259
rect 11004 -11366 11015 -11332
rect 11049 -11366 11057 -11332
rect 11004 -11389 11057 -11366
rect 11112 -11332 11164 -11259
rect 11112 -11366 11120 -11332
rect 11154 -11366 11164 -11332
rect 11112 -11389 11164 -11366
rect 11264 -11305 11314 -11259
rect 11264 -11332 11336 -11305
rect 11264 -11366 11280 -11332
rect 11314 -11366 11336 -11332
rect 11264 -11389 11336 -11366
rect 11366 -11332 11420 -11305
rect 11366 -11366 11377 -11332
rect 11411 -11366 11420 -11332
rect 11366 -11389 11420 -11366
rect 11658 -11317 11710 -11279
rect 11658 -11351 11666 -11317
rect 11700 -11351 11710 -11317
rect 11658 -11389 11710 -11351
rect 11920 -11317 11972 -11279
rect 11920 -11351 11930 -11317
rect 11964 -11351 11972 -11317
rect 11920 -11389 11972 -11351
rect 13590 -11324 13642 -11279
rect 13590 -11358 13598 -11324
rect 13632 -11358 13642 -11324
rect 13590 -11389 13642 -11358
rect 14588 -11324 14640 -11279
rect 14588 -11358 14598 -11324
rect 14632 -11358 14640 -11324
rect 14588 -11389 14640 -11358
rect 14786 -11324 14838 -11279
rect 14786 -11358 14794 -11324
rect 14828 -11358 14838 -11324
rect 14786 -11389 14838 -11358
rect 15784 -11324 15836 -11279
rect 15784 -11358 15794 -11324
rect 15828 -11358 15836 -11324
rect 15784 -11389 15836 -11358
rect 15982 -11324 16034 -11279
rect 15982 -11358 15990 -11324
rect 16024 -11358 16034 -11324
rect 15982 -11389 16034 -11358
rect 16612 -11324 16664 -11279
rect 16612 -11358 16622 -11324
rect 16656 -11358 16664 -11324
rect 16612 -11389 16664 -11358
rect -2970 -11514 -2918 -11483
rect -2970 -11548 -2962 -11514
rect -2928 -11548 -2918 -11514
rect -2970 -11593 -2918 -11548
rect -2340 -11514 -2288 -11483
rect -2340 -11548 -2330 -11514
rect -2296 -11548 -2288 -11514
rect -2340 -11593 -2288 -11548
rect -1590 -11514 -1538 -11483
rect -1590 -11548 -1582 -11514
rect -1548 -11548 -1538 -11514
rect -1590 -11593 -1538 -11548
rect -960 -11514 -908 -11483
rect -960 -11548 -950 -11514
rect -916 -11548 -908 -11514
rect -960 -11593 -908 -11548
rect -854 -11514 -802 -11483
rect -854 -11548 -846 -11514
rect -812 -11548 -802 -11514
rect -854 -11593 -802 -11548
rect -224 -11514 -172 -11483
rect -224 -11548 -214 -11514
rect -180 -11548 -172 -11514
rect -224 -11593 -172 -11548
rect -26 -11521 26 -11483
rect -26 -11555 -18 -11521
rect 16 -11555 26 -11521
rect -26 -11593 26 -11555
rect 236 -11521 288 -11483
rect 236 -11555 246 -11521
rect 280 -11555 288 -11521
rect 236 -11593 288 -11555
rect 434 -11506 488 -11483
rect 434 -11540 443 -11506
rect 477 -11540 488 -11506
rect 434 -11567 488 -11540
rect 518 -11506 590 -11483
rect 518 -11540 540 -11506
rect 574 -11540 590 -11506
rect 518 -11567 590 -11540
rect 540 -11613 590 -11567
rect 690 -11506 742 -11483
rect 690 -11540 700 -11506
rect 734 -11540 742 -11506
rect 690 -11613 742 -11540
rect 797 -11506 850 -11483
rect 797 -11540 805 -11506
rect 839 -11540 850 -11506
rect 797 -11613 850 -11540
rect 950 -11506 1015 -11483
rect 950 -11540 961 -11506
rect 995 -11540 1015 -11506
rect 950 -11567 1015 -11540
rect 1045 -11506 1116 -11483
rect 1045 -11540 1059 -11506
rect 1093 -11540 1116 -11506
rect 1045 -11567 1116 -11540
rect 950 -11613 1000 -11567
rect 1262 -11521 1314 -11483
rect 1262 -11555 1270 -11521
rect 1304 -11555 1314 -11521
rect 1262 -11593 1314 -11555
rect 1524 -11521 1576 -11483
rect 1524 -11555 1534 -11521
rect 1568 -11555 1576 -11521
rect 1524 -11593 1576 -11555
rect 1722 -11514 1774 -11483
rect 1722 -11548 1730 -11514
rect 1764 -11548 1774 -11514
rect 1722 -11593 1774 -11548
rect 2352 -11514 2404 -11483
rect 2352 -11548 2362 -11514
rect 2396 -11548 2404 -11514
rect 2352 -11593 2404 -11548
rect 2550 -11521 2602 -11483
rect 2550 -11555 2558 -11521
rect 2592 -11555 2602 -11521
rect 2550 -11593 2602 -11555
rect 2812 -11521 2864 -11483
rect 2812 -11555 2822 -11521
rect 2856 -11555 2864 -11521
rect 2812 -11593 2864 -11555
rect 3010 -11506 3064 -11483
rect 3010 -11540 3019 -11506
rect 3053 -11540 3064 -11506
rect 3010 -11567 3064 -11540
rect 3094 -11506 3166 -11483
rect 3094 -11540 3116 -11506
rect 3150 -11540 3166 -11506
rect 3094 -11567 3166 -11540
rect 3116 -11613 3166 -11567
rect 3266 -11506 3318 -11483
rect 3266 -11540 3276 -11506
rect 3310 -11540 3318 -11506
rect 3266 -11613 3318 -11540
rect 3373 -11506 3426 -11483
rect 3373 -11540 3381 -11506
rect 3415 -11540 3426 -11506
rect 3373 -11613 3426 -11540
rect 3526 -11506 3591 -11483
rect 3526 -11540 3537 -11506
rect 3571 -11540 3591 -11506
rect 3526 -11567 3591 -11540
rect 3621 -11506 3692 -11483
rect 3621 -11540 3635 -11506
rect 3669 -11540 3692 -11506
rect 3621 -11567 3692 -11540
rect 3526 -11613 3576 -11567
rect 3838 -11521 3890 -11483
rect 3838 -11555 3846 -11521
rect 3880 -11555 3890 -11521
rect 3838 -11593 3890 -11555
rect 4100 -11521 4152 -11483
rect 4100 -11555 4110 -11521
rect 4144 -11555 4152 -11521
rect 4100 -11593 4152 -11555
rect 4298 -11514 4350 -11483
rect 4298 -11548 4306 -11514
rect 4340 -11548 4350 -11514
rect 4298 -11593 4350 -11548
rect 4928 -11514 4980 -11483
rect 4928 -11548 4938 -11514
rect 4972 -11548 4980 -11514
rect 4928 -11593 4980 -11548
rect 5126 -11521 5178 -11483
rect 5126 -11555 5134 -11521
rect 5168 -11555 5178 -11521
rect 5126 -11593 5178 -11555
rect 5388 -11521 5440 -11483
rect 5388 -11555 5398 -11521
rect 5432 -11555 5440 -11521
rect 5388 -11593 5440 -11555
rect 5586 -11506 5640 -11483
rect 5586 -11540 5595 -11506
rect 5629 -11540 5640 -11506
rect 5586 -11567 5640 -11540
rect 5670 -11506 5742 -11483
rect 5670 -11540 5692 -11506
rect 5726 -11540 5742 -11506
rect 5670 -11567 5742 -11540
rect 5692 -11613 5742 -11567
rect 5842 -11506 5894 -11483
rect 5842 -11540 5852 -11506
rect 5886 -11540 5894 -11506
rect 5842 -11613 5894 -11540
rect 5949 -11506 6002 -11483
rect 5949 -11540 5957 -11506
rect 5991 -11540 6002 -11506
rect 5949 -11613 6002 -11540
rect 6102 -11506 6167 -11483
rect 6102 -11540 6113 -11506
rect 6147 -11540 6167 -11506
rect 6102 -11567 6167 -11540
rect 6197 -11506 6268 -11483
rect 6197 -11540 6211 -11506
rect 6245 -11540 6268 -11506
rect 6197 -11567 6268 -11540
rect 6102 -11613 6152 -11567
rect 6414 -11521 6466 -11483
rect 6414 -11555 6422 -11521
rect 6456 -11555 6466 -11521
rect 6414 -11593 6466 -11555
rect 6676 -11521 6728 -11483
rect 6676 -11555 6686 -11521
rect 6720 -11555 6728 -11521
rect 6676 -11593 6728 -11555
rect 6874 -11514 6926 -11483
rect 6874 -11548 6882 -11514
rect 6916 -11548 6926 -11514
rect 6874 -11593 6926 -11548
rect 7504 -11514 7556 -11483
rect 7504 -11548 7514 -11514
rect 7548 -11548 7556 -11514
rect 7504 -11593 7556 -11548
rect 7702 -11521 7754 -11483
rect 7702 -11555 7710 -11521
rect 7744 -11555 7754 -11521
rect 7702 -11593 7754 -11555
rect 7964 -11521 8016 -11483
rect 7964 -11555 7974 -11521
rect 8008 -11555 8016 -11521
rect 7964 -11593 8016 -11555
rect 8162 -11506 8216 -11483
rect 8162 -11540 8171 -11506
rect 8205 -11540 8216 -11506
rect 8162 -11567 8216 -11540
rect 8246 -11506 8318 -11483
rect 8246 -11540 8268 -11506
rect 8302 -11540 8318 -11506
rect 8246 -11567 8318 -11540
rect 8268 -11613 8318 -11567
rect 8418 -11506 8470 -11483
rect 8418 -11540 8428 -11506
rect 8462 -11540 8470 -11506
rect 8418 -11613 8470 -11540
rect 8525 -11506 8578 -11483
rect 8525 -11540 8533 -11506
rect 8567 -11540 8578 -11506
rect 8525 -11613 8578 -11540
rect 8678 -11506 8743 -11483
rect 8678 -11540 8689 -11506
rect 8723 -11540 8743 -11506
rect 8678 -11567 8743 -11540
rect 8773 -11506 8844 -11483
rect 8773 -11540 8787 -11506
rect 8821 -11540 8844 -11506
rect 8773 -11567 8844 -11540
rect 8678 -11613 8728 -11567
rect 8990 -11521 9042 -11483
rect 8990 -11555 8998 -11521
rect 9032 -11555 9042 -11521
rect 8990 -11593 9042 -11555
rect 9252 -11521 9304 -11483
rect 9252 -11555 9262 -11521
rect 9296 -11555 9304 -11521
rect 9252 -11593 9304 -11555
rect 9450 -11514 9502 -11483
rect 9450 -11548 9458 -11514
rect 9492 -11548 9502 -11514
rect 9450 -11593 9502 -11548
rect 10080 -11514 10132 -11483
rect 10080 -11548 10090 -11514
rect 10124 -11548 10132 -11514
rect 10080 -11593 10132 -11548
rect 10370 -11521 10422 -11483
rect 10370 -11555 10378 -11521
rect 10412 -11555 10422 -11521
rect 10370 -11593 10422 -11555
rect 10632 -11521 10684 -11483
rect 10632 -11555 10642 -11521
rect 10676 -11555 10684 -11521
rect 10632 -11593 10684 -11555
rect 10738 -11506 10792 -11483
rect 10738 -11540 10747 -11506
rect 10781 -11540 10792 -11506
rect 10738 -11567 10792 -11540
rect 10822 -11506 10894 -11483
rect 10822 -11540 10844 -11506
rect 10878 -11540 10894 -11506
rect 10822 -11567 10894 -11540
rect 10844 -11613 10894 -11567
rect 10994 -11506 11046 -11483
rect 10994 -11540 11004 -11506
rect 11038 -11540 11046 -11506
rect 10994 -11613 11046 -11540
rect 11101 -11506 11154 -11483
rect 11101 -11540 11109 -11506
rect 11143 -11540 11154 -11506
rect 11101 -11613 11154 -11540
rect 11254 -11506 11319 -11483
rect 11254 -11540 11265 -11506
rect 11299 -11540 11319 -11506
rect 11254 -11567 11319 -11540
rect 11349 -11506 11420 -11483
rect 11349 -11540 11363 -11506
rect 11397 -11540 11420 -11506
rect 11349 -11567 11420 -11540
rect 11254 -11613 11304 -11567
rect 11658 -11521 11710 -11483
rect 11658 -11555 11666 -11521
rect 11700 -11555 11710 -11521
rect 11658 -11593 11710 -11555
rect 11920 -11521 11972 -11483
rect 12567 -11497 12633 -11483
rect 11920 -11555 11930 -11521
rect 11964 -11555 11972 -11521
rect 11920 -11593 11972 -11555
rect 12567 -11531 12588 -11497
rect 12622 -11531 12633 -11497
rect 12567 -11567 12633 -11531
rect 12663 -11508 12719 -11483
rect 12663 -11542 12674 -11508
rect 12708 -11542 12719 -11508
rect 12663 -11567 12719 -11542
rect 12749 -11497 12805 -11483
rect 12749 -11531 12760 -11497
rect 12794 -11531 12805 -11497
rect 12749 -11567 12805 -11531
rect 12835 -11508 12891 -11483
rect 12835 -11542 12846 -11508
rect 12880 -11542 12891 -11508
rect 12835 -11567 12891 -11542
rect 12921 -11497 13000 -11483
rect 12921 -11531 12932 -11497
rect 12966 -11531 13000 -11497
rect 12921 -11567 13000 -11531
rect 13222 -11521 13274 -11483
rect 13222 -11555 13230 -11521
rect 13264 -11555 13274 -11521
rect 13222 -11593 13274 -11555
rect 13484 -11521 13536 -11483
rect 13682 -11495 13735 -11483
rect 13484 -11555 13494 -11521
rect 13528 -11555 13536 -11521
rect 13484 -11593 13536 -11555
rect 13682 -11529 13690 -11495
rect 13724 -11529 13735 -11495
rect 13682 -11567 13735 -11529
rect 13765 -11508 13821 -11483
rect 13765 -11542 13776 -11508
rect 13810 -11542 13821 -11508
rect 13765 -11567 13821 -11542
rect 13851 -11508 13907 -11483
rect 13851 -11542 13862 -11508
rect 13896 -11542 13907 -11508
rect 13851 -11567 13907 -11542
rect 13937 -11508 13993 -11483
rect 13937 -11542 13948 -11508
rect 13982 -11542 13993 -11508
rect 13937 -11567 13993 -11542
rect 14023 -11508 14079 -11483
rect 14023 -11542 14034 -11508
rect 14068 -11542 14079 -11508
rect 14023 -11567 14079 -11542
rect 14109 -11508 14165 -11483
rect 14109 -11542 14120 -11508
rect 14154 -11542 14165 -11508
rect 14109 -11567 14165 -11542
rect 14195 -11499 14251 -11483
rect 14195 -11533 14206 -11499
rect 14240 -11533 14251 -11499
rect 14195 -11567 14251 -11533
rect 14281 -11508 14337 -11483
rect 14281 -11542 14292 -11508
rect 14326 -11542 14337 -11508
rect 14281 -11567 14337 -11542
rect 14367 -11499 14423 -11483
rect 14367 -11533 14378 -11499
rect 14412 -11533 14423 -11499
rect 14367 -11567 14423 -11533
rect 14453 -11508 14509 -11483
rect 14453 -11542 14464 -11508
rect 14498 -11542 14509 -11508
rect 14453 -11567 14509 -11542
rect 14539 -11499 14595 -11483
rect 14539 -11533 14550 -11499
rect 14584 -11533 14595 -11499
rect 14539 -11567 14595 -11533
rect 14625 -11508 14681 -11483
rect 14625 -11542 14636 -11508
rect 14670 -11542 14681 -11508
rect 14625 -11567 14681 -11542
rect 14711 -11499 14766 -11483
rect 14711 -11533 14722 -11499
rect 14756 -11533 14766 -11499
rect 14711 -11567 14766 -11533
rect 14796 -11508 14852 -11483
rect 14796 -11542 14807 -11508
rect 14841 -11542 14852 -11508
rect 14796 -11567 14852 -11542
rect 14882 -11499 14938 -11483
rect 14882 -11533 14893 -11499
rect 14927 -11533 14938 -11499
rect 14882 -11567 14938 -11533
rect 14968 -11508 15024 -11483
rect 14968 -11542 14979 -11508
rect 15013 -11542 15024 -11508
rect 14968 -11567 15024 -11542
rect 15054 -11499 15110 -11483
rect 15054 -11533 15065 -11499
rect 15099 -11533 15110 -11499
rect 15054 -11567 15110 -11533
rect 15140 -11508 15196 -11483
rect 15140 -11542 15151 -11508
rect 15185 -11542 15196 -11508
rect 15140 -11567 15196 -11542
rect 15226 -11499 15282 -11483
rect 15226 -11533 15237 -11499
rect 15271 -11533 15282 -11499
rect 15226 -11567 15282 -11533
rect 15312 -11508 15368 -11483
rect 15312 -11542 15323 -11508
rect 15357 -11542 15368 -11508
rect 15312 -11567 15368 -11542
rect 15398 -11499 15451 -11483
rect 15398 -11533 15409 -11499
rect 15443 -11533 15451 -11499
rect 15398 -11567 15451 -11533
rect 15614 -11514 15666 -11483
rect 15614 -11548 15622 -11514
rect 15656 -11548 15666 -11514
rect 15614 -11593 15666 -11548
rect 16612 -11514 16664 -11483
rect 16612 -11548 16622 -11514
rect 16656 -11548 16664 -11514
rect 16612 -11593 16664 -11548
rect -2970 -12412 -2918 -12367
rect -2970 -12446 -2962 -12412
rect -2928 -12446 -2918 -12412
rect -2970 -12477 -2918 -12446
rect -2340 -12412 -2288 -12367
rect -2340 -12446 -2330 -12412
rect -2296 -12446 -2288 -12412
rect -2340 -12477 -2288 -12446
rect -1590 -12412 -1538 -12367
rect -1590 -12446 -1582 -12412
rect -1548 -12446 -1538 -12412
rect -1590 -12477 -1538 -12446
rect -960 -12412 -908 -12367
rect -738 -12393 -688 -12347
rect -960 -12446 -950 -12412
rect -916 -12446 -908 -12412
rect -960 -12477 -908 -12446
rect -854 -12420 -783 -12393
rect -854 -12454 -831 -12420
rect -797 -12454 -783 -12420
rect -854 -12477 -783 -12454
rect -753 -12420 -688 -12393
rect -753 -12454 -733 -12420
rect -699 -12454 -688 -12420
rect -753 -12477 -688 -12454
rect -588 -12420 -535 -12347
rect -588 -12454 -577 -12420
rect -543 -12454 -535 -12420
rect -588 -12477 -535 -12454
rect -480 -12420 -428 -12347
rect -480 -12454 -472 -12420
rect -438 -12454 -428 -12420
rect -480 -12477 -428 -12454
rect -328 -12393 -278 -12347
rect -328 -12420 -256 -12393
rect -328 -12454 -312 -12420
rect -278 -12454 -256 -12420
rect -328 -12477 -256 -12454
rect -226 -12420 -172 -12393
rect -226 -12454 -215 -12420
rect -181 -12454 -172 -12420
rect -226 -12477 -172 -12454
rect -26 -12405 26 -12367
rect -26 -12439 -18 -12405
rect 16 -12439 26 -12405
rect -26 -12477 26 -12439
rect 236 -12405 288 -12367
rect 236 -12439 246 -12405
rect 280 -12439 288 -12405
rect 236 -12477 288 -12439
rect 550 -12393 600 -12347
rect 434 -12420 505 -12393
rect 434 -12454 457 -12420
rect 491 -12454 505 -12420
rect 434 -12477 505 -12454
rect 535 -12420 600 -12393
rect 535 -12454 555 -12420
rect 589 -12454 600 -12420
rect 535 -12477 600 -12454
rect 700 -12420 753 -12347
rect 700 -12454 711 -12420
rect 745 -12454 753 -12420
rect 700 -12477 753 -12454
rect 808 -12420 860 -12347
rect 808 -12454 816 -12420
rect 850 -12454 860 -12420
rect 808 -12477 860 -12454
rect 960 -12393 1010 -12347
rect 960 -12420 1032 -12393
rect 960 -12454 976 -12420
rect 1010 -12454 1032 -12420
rect 960 -12477 1032 -12454
rect 1062 -12420 1116 -12393
rect 1062 -12454 1073 -12420
rect 1107 -12454 1116 -12420
rect 1062 -12477 1116 -12454
rect 1262 -12405 1314 -12367
rect 1262 -12439 1270 -12405
rect 1304 -12439 1314 -12405
rect 1262 -12477 1314 -12439
rect 1524 -12405 1576 -12367
rect 1524 -12439 1534 -12405
rect 1568 -12439 1576 -12405
rect 1524 -12477 1576 -12439
rect 1722 -12412 1774 -12367
rect 1722 -12446 1730 -12412
rect 1764 -12446 1774 -12412
rect 1722 -12477 1774 -12446
rect 2352 -12412 2404 -12367
rect 2352 -12446 2362 -12412
rect 2396 -12446 2404 -12412
rect 2352 -12477 2404 -12446
rect 2550 -12405 2602 -12367
rect 2550 -12439 2558 -12405
rect 2592 -12439 2602 -12405
rect 2550 -12477 2602 -12439
rect 2812 -12405 2864 -12367
rect 2812 -12439 2822 -12405
rect 2856 -12439 2864 -12405
rect 2812 -12477 2864 -12439
rect 3126 -12393 3176 -12347
rect 3010 -12420 3081 -12393
rect 3010 -12454 3033 -12420
rect 3067 -12454 3081 -12420
rect 3010 -12477 3081 -12454
rect 3111 -12420 3176 -12393
rect 3111 -12454 3131 -12420
rect 3165 -12454 3176 -12420
rect 3111 -12477 3176 -12454
rect 3276 -12420 3329 -12347
rect 3276 -12454 3287 -12420
rect 3321 -12454 3329 -12420
rect 3276 -12477 3329 -12454
rect 3384 -12420 3436 -12347
rect 3384 -12454 3392 -12420
rect 3426 -12454 3436 -12420
rect 3384 -12477 3436 -12454
rect 3536 -12393 3586 -12347
rect 3536 -12420 3608 -12393
rect 3536 -12454 3552 -12420
rect 3586 -12454 3608 -12420
rect 3536 -12477 3608 -12454
rect 3638 -12420 3692 -12393
rect 3638 -12454 3649 -12420
rect 3683 -12454 3692 -12420
rect 3638 -12477 3692 -12454
rect 3838 -12405 3890 -12367
rect 3838 -12439 3846 -12405
rect 3880 -12439 3890 -12405
rect 3838 -12477 3890 -12439
rect 4100 -12405 4152 -12367
rect 4100 -12439 4110 -12405
rect 4144 -12439 4152 -12405
rect 4100 -12477 4152 -12439
rect 4298 -12412 4350 -12367
rect 4298 -12446 4306 -12412
rect 4340 -12446 4350 -12412
rect 4298 -12477 4350 -12446
rect 4928 -12412 4980 -12367
rect 4928 -12446 4938 -12412
rect 4972 -12446 4980 -12412
rect 4928 -12477 4980 -12446
rect 5126 -12405 5178 -12367
rect 5126 -12439 5134 -12405
rect 5168 -12439 5178 -12405
rect 5126 -12477 5178 -12439
rect 5388 -12405 5440 -12367
rect 5388 -12439 5398 -12405
rect 5432 -12439 5440 -12405
rect 5388 -12477 5440 -12439
rect 5702 -12393 5752 -12347
rect 5586 -12420 5657 -12393
rect 5586 -12454 5609 -12420
rect 5643 -12454 5657 -12420
rect 5586 -12477 5657 -12454
rect 5687 -12420 5752 -12393
rect 5687 -12454 5707 -12420
rect 5741 -12454 5752 -12420
rect 5687 -12477 5752 -12454
rect 5852 -12420 5905 -12347
rect 5852 -12454 5863 -12420
rect 5897 -12454 5905 -12420
rect 5852 -12477 5905 -12454
rect 5960 -12420 6012 -12347
rect 5960 -12454 5968 -12420
rect 6002 -12454 6012 -12420
rect 5960 -12477 6012 -12454
rect 6112 -12393 6162 -12347
rect 6112 -12420 6184 -12393
rect 6112 -12454 6128 -12420
rect 6162 -12454 6184 -12420
rect 6112 -12477 6184 -12454
rect 6214 -12420 6268 -12393
rect 6214 -12454 6225 -12420
rect 6259 -12454 6268 -12420
rect 6214 -12477 6268 -12454
rect 6414 -12405 6466 -12367
rect 6414 -12439 6422 -12405
rect 6456 -12439 6466 -12405
rect 6414 -12477 6466 -12439
rect 6676 -12405 6728 -12367
rect 6676 -12439 6686 -12405
rect 6720 -12439 6728 -12405
rect 6676 -12477 6728 -12439
rect 6874 -12412 6926 -12367
rect 6874 -12446 6882 -12412
rect 6916 -12446 6926 -12412
rect 6874 -12477 6926 -12446
rect 7504 -12412 7556 -12367
rect 7504 -12446 7514 -12412
rect 7548 -12446 7556 -12412
rect 7504 -12477 7556 -12446
rect 7702 -12405 7754 -12367
rect 7702 -12439 7710 -12405
rect 7744 -12439 7754 -12405
rect 7702 -12477 7754 -12439
rect 7964 -12405 8016 -12367
rect 7964 -12439 7974 -12405
rect 8008 -12439 8016 -12405
rect 7964 -12477 8016 -12439
rect 8278 -12393 8328 -12347
rect 8162 -12420 8233 -12393
rect 8162 -12454 8185 -12420
rect 8219 -12454 8233 -12420
rect 8162 -12477 8233 -12454
rect 8263 -12420 8328 -12393
rect 8263 -12454 8283 -12420
rect 8317 -12454 8328 -12420
rect 8263 -12477 8328 -12454
rect 8428 -12420 8481 -12347
rect 8428 -12454 8439 -12420
rect 8473 -12454 8481 -12420
rect 8428 -12477 8481 -12454
rect 8536 -12420 8588 -12347
rect 8536 -12454 8544 -12420
rect 8578 -12454 8588 -12420
rect 8536 -12477 8588 -12454
rect 8688 -12393 8738 -12347
rect 8688 -12420 8760 -12393
rect 8688 -12454 8704 -12420
rect 8738 -12454 8760 -12420
rect 8688 -12477 8760 -12454
rect 8790 -12420 8844 -12393
rect 8790 -12454 8801 -12420
rect 8835 -12454 8844 -12420
rect 8790 -12477 8844 -12454
rect 8990 -12405 9042 -12367
rect 8990 -12439 8998 -12405
rect 9032 -12439 9042 -12405
rect 8990 -12477 9042 -12439
rect 9252 -12405 9304 -12367
rect 9252 -12439 9262 -12405
rect 9296 -12439 9304 -12405
rect 9252 -12477 9304 -12439
rect 9450 -12412 9502 -12367
rect 9450 -12446 9458 -12412
rect 9492 -12446 9502 -12412
rect 9450 -12477 9502 -12446
rect 10080 -12412 10132 -12367
rect 10080 -12446 10090 -12412
rect 10124 -12446 10132 -12412
rect 10080 -12477 10132 -12446
rect 10370 -12405 10422 -12367
rect 10370 -12439 10378 -12405
rect 10412 -12439 10422 -12405
rect 10370 -12477 10422 -12439
rect 10632 -12405 10684 -12367
rect 10854 -12393 10904 -12347
rect 10632 -12439 10642 -12405
rect 10676 -12439 10684 -12405
rect 10632 -12477 10684 -12439
rect 10738 -12420 10809 -12393
rect 10738 -12454 10761 -12420
rect 10795 -12454 10809 -12420
rect 10738 -12477 10809 -12454
rect 10839 -12420 10904 -12393
rect 10839 -12454 10859 -12420
rect 10893 -12454 10904 -12420
rect 10839 -12477 10904 -12454
rect 11004 -12420 11057 -12347
rect 11004 -12454 11015 -12420
rect 11049 -12454 11057 -12420
rect 11004 -12477 11057 -12454
rect 11112 -12420 11164 -12347
rect 11112 -12454 11120 -12420
rect 11154 -12454 11164 -12420
rect 11112 -12477 11164 -12454
rect 11264 -12393 11314 -12347
rect 11264 -12420 11336 -12393
rect 11264 -12454 11280 -12420
rect 11314 -12454 11336 -12420
rect 11264 -12477 11336 -12454
rect 11366 -12420 11420 -12393
rect 11366 -12454 11377 -12420
rect 11411 -12454 11420 -12420
rect 11366 -12477 11420 -12454
rect 11658 -12405 11710 -12367
rect 11658 -12439 11666 -12405
rect 11700 -12439 11710 -12405
rect 11658 -12477 11710 -12439
rect 11920 -12405 11972 -12367
rect 11920 -12439 11930 -12405
rect 11964 -12439 11972 -12405
rect 11920 -12477 11972 -12439
rect 13682 -12431 13735 -12393
rect 13682 -12465 13690 -12431
rect 13724 -12465 13735 -12431
rect 13682 -12477 13735 -12465
rect 13765 -12418 13821 -12393
rect 13765 -12452 13776 -12418
rect 13810 -12452 13821 -12418
rect 13765 -12477 13821 -12452
rect 13851 -12418 13907 -12393
rect 13851 -12452 13862 -12418
rect 13896 -12452 13907 -12418
rect 13851 -12477 13907 -12452
rect 13937 -12418 13993 -12393
rect 13937 -12452 13948 -12418
rect 13982 -12452 13993 -12418
rect 13937 -12477 13993 -12452
rect 14023 -12418 14079 -12393
rect 14023 -12452 14034 -12418
rect 14068 -12452 14079 -12418
rect 14023 -12477 14079 -12452
rect 14109 -12418 14165 -12393
rect 14109 -12452 14120 -12418
rect 14154 -12452 14165 -12418
rect 14109 -12477 14165 -12452
rect 14195 -12427 14251 -12393
rect 14195 -12461 14206 -12427
rect 14240 -12461 14251 -12427
rect 14195 -12477 14251 -12461
rect 14281 -12418 14337 -12393
rect 14281 -12452 14292 -12418
rect 14326 -12452 14337 -12418
rect 14281 -12477 14337 -12452
rect 14367 -12427 14423 -12393
rect 14367 -12461 14378 -12427
rect 14412 -12461 14423 -12427
rect 14367 -12477 14423 -12461
rect 14453 -12418 14509 -12393
rect 14453 -12452 14464 -12418
rect 14498 -12452 14509 -12418
rect 14453 -12477 14509 -12452
rect 14539 -12427 14595 -12393
rect 14539 -12461 14550 -12427
rect 14584 -12461 14595 -12427
rect 14539 -12477 14595 -12461
rect 14625 -12418 14681 -12393
rect 14625 -12452 14636 -12418
rect 14670 -12452 14681 -12418
rect 14625 -12477 14681 -12452
rect 14711 -12427 14766 -12393
rect 14711 -12461 14722 -12427
rect 14756 -12461 14766 -12427
rect 14711 -12477 14766 -12461
rect 14796 -12418 14852 -12393
rect 14796 -12452 14807 -12418
rect 14841 -12452 14852 -12418
rect 14796 -12477 14852 -12452
rect 14882 -12427 14938 -12393
rect 14882 -12461 14893 -12427
rect 14927 -12461 14938 -12427
rect 14882 -12477 14938 -12461
rect 14968 -12418 15024 -12393
rect 14968 -12452 14979 -12418
rect 15013 -12452 15024 -12418
rect 14968 -12477 15024 -12452
rect 15054 -12427 15110 -12393
rect 15054 -12461 15065 -12427
rect 15099 -12461 15110 -12427
rect 15054 -12477 15110 -12461
rect 15140 -12418 15196 -12393
rect 15140 -12452 15151 -12418
rect 15185 -12452 15196 -12418
rect 15140 -12477 15196 -12452
rect 15226 -12427 15282 -12393
rect 15226 -12461 15237 -12427
rect 15271 -12461 15282 -12427
rect 15226 -12477 15282 -12461
rect 15312 -12418 15368 -12393
rect 15312 -12452 15323 -12418
rect 15357 -12452 15368 -12418
rect 15312 -12477 15368 -12452
rect 15398 -12427 15451 -12393
rect 15398 -12461 15409 -12427
rect 15443 -12461 15451 -12427
rect 15614 -12412 15666 -12367
rect 15614 -12446 15622 -12412
rect 15656 -12446 15666 -12412
rect 15398 -12477 15451 -12461
rect 15614 -12477 15666 -12446
rect 16612 -12412 16664 -12367
rect 16612 -12446 16622 -12412
rect 16656 -12446 16664 -12412
rect 16612 -12477 16664 -12446
rect -2970 -12602 -2918 -12571
rect -2970 -12636 -2962 -12602
rect -2928 -12636 -2918 -12602
rect -2970 -12681 -2918 -12636
rect -2340 -12602 -2288 -12571
rect -2340 -12636 -2330 -12602
rect -2296 -12636 -2288 -12602
rect -2340 -12681 -2288 -12636
rect -1590 -12602 -1538 -12571
rect -1590 -12636 -1582 -12602
rect -1548 -12636 -1538 -12602
rect -1590 -12681 -1538 -12636
rect -960 -12602 -908 -12571
rect -960 -12636 -950 -12602
rect -916 -12636 -908 -12602
rect -960 -12681 -908 -12636
rect -854 -12602 -802 -12571
rect -854 -12636 -846 -12602
rect -812 -12636 -802 -12602
rect -854 -12681 -802 -12636
rect -224 -12602 -172 -12571
rect -224 -12636 -214 -12602
rect -180 -12636 -172 -12602
rect -224 -12681 -172 -12636
rect -26 -12609 26 -12571
rect -26 -12643 -18 -12609
rect 16 -12643 26 -12609
rect -26 -12681 26 -12643
rect 236 -12609 288 -12571
rect 236 -12643 246 -12609
rect 280 -12643 288 -12609
rect 236 -12681 288 -12643
rect 434 -12594 488 -12571
rect 434 -12628 443 -12594
rect 477 -12628 488 -12594
rect 434 -12655 488 -12628
rect 518 -12594 590 -12571
rect 518 -12628 540 -12594
rect 574 -12628 590 -12594
rect 518 -12655 590 -12628
rect 540 -12701 590 -12655
rect 690 -12594 742 -12571
rect 690 -12628 700 -12594
rect 734 -12628 742 -12594
rect 690 -12701 742 -12628
rect 797 -12594 850 -12571
rect 797 -12628 805 -12594
rect 839 -12628 850 -12594
rect 797 -12701 850 -12628
rect 950 -12594 1015 -12571
rect 950 -12628 961 -12594
rect 995 -12628 1015 -12594
rect 950 -12655 1015 -12628
rect 1045 -12594 1116 -12571
rect 1045 -12628 1059 -12594
rect 1093 -12628 1116 -12594
rect 1045 -12655 1116 -12628
rect 950 -12701 1000 -12655
rect 1262 -12609 1314 -12571
rect 1262 -12643 1270 -12609
rect 1304 -12643 1314 -12609
rect 1262 -12681 1314 -12643
rect 1524 -12609 1576 -12571
rect 1524 -12643 1534 -12609
rect 1568 -12643 1576 -12609
rect 1524 -12681 1576 -12643
rect 1722 -12602 1774 -12571
rect 1722 -12636 1730 -12602
rect 1764 -12636 1774 -12602
rect 1722 -12681 1774 -12636
rect 2352 -12602 2404 -12571
rect 2352 -12636 2362 -12602
rect 2396 -12636 2404 -12602
rect 2352 -12681 2404 -12636
rect 2550 -12609 2602 -12571
rect 2550 -12643 2558 -12609
rect 2592 -12643 2602 -12609
rect 2550 -12681 2602 -12643
rect 2812 -12609 2864 -12571
rect 2812 -12643 2822 -12609
rect 2856 -12643 2864 -12609
rect 2812 -12681 2864 -12643
rect 3010 -12594 3064 -12571
rect 3010 -12628 3019 -12594
rect 3053 -12628 3064 -12594
rect 3010 -12655 3064 -12628
rect 3094 -12594 3166 -12571
rect 3094 -12628 3116 -12594
rect 3150 -12628 3166 -12594
rect 3094 -12655 3166 -12628
rect 3116 -12701 3166 -12655
rect 3266 -12594 3318 -12571
rect 3266 -12628 3276 -12594
rect 3310 -12628 3318 -12594
rect 3266 -12701 3318 -12628
rect 3373 -12594 3426 -12571
rect 3373 -12628 3381 -12594
rect 3415 -12628 3426 -12594
rect 3373 -12701 3426 -12628
rect 3526 -12594 3591 -12571
rect 3526 -12628 3537 -12594
rect 3571 -12628 3591 -12594
rect 3526 -12655 3591 -12628
rect 3621 -12594 3692 -12571
rect 3621 -12628 3635 -12594
rect 3669 -12628 3692 -12594
rect 3621 -12655 3692 -12628
rect 3526 -12701 3576 -12655
rect 3838 -12609 3890 -12571
rect 3838 -12643 3846 -12609
rect 3880 -12643 3890 -12609
rect 3838 -12681 3890 -12643
rect 4100 -12609 4152 -12571
rect 4100 -12643 4110 -12609
rect 4144 -12643 4152 -12609
rect 4100 -12681 4152 -12643
rect 4298 -12602 4350 -12571
rect 4298 -12636 4306 -12602
rect 4340 -12636 4350 -12602
rect 4298 -12681 4350 -12636
rect 4928 -12602 4980 -12571
rect 4928 -12636 4938 -12602
rect 4972 -12636 4980 -12602
rect 4928 -12681 4980 -12636
rect 5126 -12609 5178 -12571
rect 5126 -12643 5134 -12609
rect 5168 -12643 5178 -12609
rect 5126 -12681 5178 -12643
rect 5388 -12609 5440 -12571
rect 5388 -12643 5398 -12609
rect 5432 -12643 5440 -12609
rect 5388 -12681 5440 -12643
rect 5586 -12594 5640 -12571
rect 5586 -12628 5595 -12594
rect 5629 -12628 5640 -12594
rect 5586 -12655 5640 -12628
rect 5670 -12594 5742 -12571
rect 5670 -12628 5692 -12594
rect 5726 -12628 5742 -12594
rect 5670 -12655 5742 -12628
rect 5692 -12701 5742 -12655
rect 5842 -12594 5894 -12571
rect 5842 -12628 5852 -12594
rect 5886 -12628 5894 -12594
rect 5842 -12701 5894 -12628
rect 5949 -12594 6002 -12571
rect 5949 -12628 5957 -12594
rect 5991 -12628 6002 -12594
rect 5949 -12701 6002 -12628
rect 6102 -12594 6167 -12571
rect 6102 -12628 6113 -12594
rect 6147 -12628 6167 -12594
rect 6102 -12655 6167 -12628
rect 6197 -12594 6268 -12571
rect 6197 -12628 6211 -12594
rect 6245 -12628 6268 -12594
rect 6197 -12655 6268 -12628
rect 6102 -12701 6152 -12655
rect 6414 -12609 6466 -12571
rect 6414 -12643 6422 -12609
rect 6456 -12643 6466 -12609
rect 6414 -12681 6466 -12643
rect 6676 -12609 6728 -12571
rect 6676 -12643 6686 -12609
rect 6720 -12643 6728 -12609
rect 6676 -12681 6728 -12643
rect 6874 -12602 6926 -12571
rect 6874 -12636 6882 -12602
rect 6916 -12636 6926 -12602
rect 6874 -12681 6926 -12636
rect 7504 -12602 7556 -12571
rect 7504 -12636 7514 -12602
rect 7548 -12636 7556 -12602
rect 7504 -12681 7556 -12636
rect 7702 -12609 7754 -12571
rect 7702 -12643 7710 -12609
rect 7744 -12643 7754 -12609
rect 7702 -12681 7754 -12643
rect 7964 -12609 8016 -12571
rect 7964 -12643 7974 -12609
rect 8008 -12643 8016 -12609
rect 7964 -12681 8016 -12643
rect 8162 -12594 8216 -12571
rect 8162 -12628 8171 -12594
rect 8205 -12628 8216 -12594
rect 8162 -12655 8216 -12628
rect 8246 -12594 8318 -12571
rect 8246 -12628 8268 -12594
rect 8302 -12628 8318 -12594
rect 8246 -12655 8318 -12628
rect 8268 -12701 8318 -12655
rect 8418 -12594 8470 -12571
rect 8418 -12628 8428 -12594
rect 8462 -12628 8470 -12594
rect 8418 -12701 8470 -12628
rect 8525 -12594 8578 -12571
rect 8525 -12628 8533 -12594
rect 8567 -12628 8578 -12594
rect 8525 -12701 8578 -12628
rect 8678 -12594 8743 -12571
rect 8678 -12628 8689 -12594
rect 8723 -12628 8743 -12594
rect 8678 -12655 8743 -12628
rect 8773 -12594 8844 -12571
rect 8773 -12628 8787 -12594
rect 8821 -12628 8844 -12594
rect 8773 -12655 8844 -12628
rect 8678 -12701 8728 -12655
rect 8990 -12609 9042 -12571
rect 8990 -12643 8998 -12609
rect 9032 -12643 9042 -12609
rect 8990 -12681 9042 -12643
rect 9252 -12609 9304 -12571
rect 9252 -12643 9262 -12609
rect 9296 -12643 9304 -12609
rect 9252 -12681 9304 -12643
rect 9450 -12602 9502 -12571
rect 9450 -12636 9458 -12602
rect 9492 -12636 9502 -12602
rect 9450 -12681 9502 -12636
rect 10080 -12602 10132 -12571
rect 10080 -12636 10090 -12602
rect 10124 -12636 10132 -12602
rect 10080 -12681 10132 -12636
rect 10370 -12609 10422 -12571
rect 10370 -12643 10378 -12609
rect 10412 -12643 10422 -12609
rect 10370 -12681 10422 -12643
rect 10632 -12609 10684 -12571
rect 10632 -12643 10642 -12609
rect 10676 -12643 10684 -12609
rect 10632 -12681 10684 -12643
rect 10738 -12594 10792 -12571
rect 10738 -12628 10747 -12594
rect 10781 -12628 10792 -12594
rect 10738 -12655 10792 -12628
rect 10822 -12594 10894 -12571
rect 10822 -12628 10844 -12594
rect 10878 -12628 10894 -12594
rect 10822 -12655 10894 -12628
rect 10844 -12701 10894 -12655
rect 10994 -12594 11046 -12571
rect 10994 -12628 11004 -12594
rect 11038 -12628 11046 -12594
rect 10994 -12701 11046 -12628
rect 11101 -12594 11154 -12571
rect 11101 -12628 11109 -12594
rect 11143 -12628 11154 -12594
rect 11101 -12701 11154 -12628
rect 11254 -12594 11319 -12571
rect 11254 -12628 11265 -12594
rect 11299 -12628 11319 -12594
rect 11254 -12655 11319 -12628
rect 11349 -12594 11420 -12571
rect 11349 -12628 11363 -12594
rect 11397 -12628 11420 -12594
rect 11349 -12655 11420 -12628
rect 11254 -12701 11304 -12655
rect 11658 -12609 11710 -12571
rect 11658 -12643 11666 -12609
rect 11700 -12643 11710 -12609
rect 11658 -12681 11710 -12643
rect 11920 -12609 11972 -12571
rect 12567 -12585 12633 -12571
rect 11920 -12643 11930 -12609
rect 11964 -12643 11972 -12609
rect 11920 -12681 11972 -12643
rect 12567 -12619 12588 -12585
rect 12622 -12619 12633 -12585
rect 12567 -12655 12633 -12619
rect 12663 -12596 12719 -12571
rect 12663 -12630 12674 -12596
rect 12708 -12630 12719 -12596
rect 12663 -12655 12719 -12630
rect 12749 -12585 12805 -12571
rect 12749 -12619 12760 -12585
rect 12794 -12619 12805 -12585
rect 12749 -12655 12805 -12619
rect 12835 -12596 12891 -12571
rect 12835 -12630 12846 -12596
rect 12880 -12630 12891 -12596
rect 12835 -12655 12891 -12630
rect 12921 -12585 13000 -12571
rect 12921 -12619 12932 -12585
rect 12966 -12619 13000 -12585
rect 12921 -12655 13000 -12619
rect 13222 -12609 13274 -12571
rect 13222 -12643 13230 -12609
rect 13264 -12643 13274 -12609
rect 13222 -12681 13274 -12643
rect 13484 -12609 13536 -12571
rect 13682 -12583 13735 -12571
rect 13484 -12643 13494 -12609
rect 13528 -12643 13536 -12609
rect 13484 -12681 13536 -12643
rect 13682 -12617 13690 -12583
rect 13724 -12617 13735 -12583
rect 13682 -12655 13735 -12617
rect 13765 -12596 13821 -12571
rect 13765 -12630 13776 -12596
rect 13810 -12630 13821 -12596
rect 13765 -12655 13821 -12630
rect 13851 -12596 13907 -12571
rect 13851 -12630 13862 -12596
rect 13896 -12630 13907 -12596
rect 13851 -12655 13907 -12630
rect 13937 -12596 13993 -12571
rect 13937 -12630 13948 -12596
rect 13982 -12630 13993 -12596
rect 13937 -12655 13993 -12630
rect 14023 -12596 14079 -12571
rect 14023 -12630 14034 -12596
rect 14068 -12630 14079 -12596
rect 14023 -12655 14079 -12630
rect 14109 -12596 14165 -12571
rect 14109 -12630 14120 -12596
rect 14154 -12630 14165 -12596
rect 14109 -12655 14165 -12630
rect 14195 -12587 14251 -12571
rect 14195 -12621 14206 -12587
rect 14240 -12621 14251 -12587
rect 14195 -12655 14251 -12621
rect 14281 -12596 14337 -12571
rect 14281 -12630 14292 -12596
rect 14326 -12630 14337 -12596
rect 14281 -12655 14337 -12630
rect 14367 -12587 14423 -12571
rect 14367 -12621 14378 -12587
rect 14412 -12621 14423 -12587
rect 14367 -12655 14423 -12621
rect 14453 -12596 14509 -12571
rect 14453 -12630 14464 -12596
rect 14498 -12630 14509 -12596
rect 14453 -12655 14509 -12630
rect 14539 -12587 14595 -12571
rect 14539 -12621 14550 -12587
rect 14584 -12621 14595 -12587
rect 14539 -12655 14595 -12621
rect 14625 -12596 14681 -12571
rect 14625 -12630 14636 -12596
rect 14670 -12630 14681 -12596
rect 14625 -12655 14681 -12630
rect 14711 -12587 14766 -12571
rect 14711 -12621 14722 -12587
rect 14756 -12621 14766 -12587
rect 14711 -12655 14766 -12621
rect 14796 -12596 14852 -12571
rect 14796 -12630 14807 -12596
rect 14841 -12630 14852 -12596
rect 14796 -12655 14852 -12630
rect 14882 -12587 14938 -12571
rect 14882 -12621 14893 -12587
rect 14927 -12621 14938 -12587
rect 14882 -12655 14938 -12621
rect 14968 -12596 15024 -12571
rect 14968 -12630 14979 -12596
rect 15013 -12630 15024 -12596
rect 14968 -12655 15024 -12630
rect 15054 -12587 15110 -12571
rect 15054 -12621 15065 -12587
rect 15099 -12621 15110 -12587
rect 15054 -12655 15110 -12621
rect 15140 -12596 15196 -12571
rect 15140 -12630 15151 -12596
rect 15185 -12630 15196 -12596
rect 15140 -12655 15196 -12630
rect 15226 -12587 15282 -12571
rect 15226 -12621 15237 -12587
rect 15271 -12621 15282 -12587
rect 15226 -12655 15282 -12621
rect 15312 -12596 15368 -12571
rect 15312 -12630 15323 -12596
rect 15357 -12630 15368 -12596
rect 15312 -12655 15368 -12630
rect 15398 -12587 15451 -12571
rect 15398 -12621 15409 -12587
rect 15443 -12621 15451 -12587
rect 15398 -12655 15451 -12621
rect 15614 -12602 15666 -12571
rect 15614 -12636 15622 -12602
rect 15656 -12636 15666 -12602
rect 15614 -12681 15666 -12636
rect 16612 -12602 16664 -12571
rect 16612 -12636 16622 -12602
rect 16656 -12636 16664 -12602
rect 16612 -12681 16664 -12636
rect -2970 -13500 -2918 -13455
rect -2970 -13534 -2962 -13500
rect -2928 -13534 -2918 -13500
rect -2970 -13565 -2918 -13534
rect -2340 -13500 -2288 -13455
rect -2340 -13534 -2330 -13500
rect -2296 -13534 -2288 -13500
rect -2340 -13565 -2288 -13534
rect -1590 -13500 -1538 -13455
rect -1590 -13534 -1582 -13500
rect -1548 -13534 -1538 -13500
rect -1590 -13565 -1538 -13534
rect -960 -13500 -908 -13455
rect -960 -13534 -950 -13500
rect -916 -13534 -908 -13500
rect -960 -13565 -908 -13534
rect -854 -13500 -802 -13455
rect -854 -13534 -846 -13500
rect -812 -13534 -802 -13500
rect -854 -13565 -802 -13534
rect -224 -13500 -172 -13455
rect -224 -13534 -214 -13500
rect -180 -13534 -172 -13500
rect -224 -13565 -172 -13534
rect -26 -13493 26 -13455
rect -26 -13527 -18 -13493
rect 16 -13527 26 -13493
rect -26 -13565 26 -13527
rect 236 -13493 288 -13455
rect 236 -13527 246 -13493
rect 280 -13527 288 -13493
rect 236 -13565 288 -13527
rect 550 -13481 600 -13435
rect 434 -13508 505 -13481
rect 434 -13542 457 -13508
rect 491 -13542 505 -13508
rect 434 -13565 505 -13542
rect 535 -13508 600 -13481
rect 535 -13542 555 -13508
rect 589 -13542 600 -13508
rect 535 -13565 600 -13542
rect 700 -13508 753 -13435
rect 700 -13542 711 -13508
rect 745 -13542 753 -13508
rect 700 -13565 753 -13542
rect 808 -13508 860 -13435
rect 808 -13542 816 -13508
rect 850 -13542 860 -13508
rect 808 -13565 860 -13542
rect 960 -13481 1010 -13435
rect 960 -13508 1032 -13481
rect 960 -13542 976 -13508
rect 1010 -13542 1032 -13508
rect 960 -13565 1032 -13542
rect 1062 -13508 1116 -13481
rect 1062 -13542 1073 -13508
rect 1107 -13542 1116 -13508
rect 1062 -13565 1116 -13542
rect 1262 -13493 1314 -13455
rect 1262 -13527 1270 -13493
rect 1304 -13527 1314 -13493
rect 1262 -13565 1314 -13527
rect 1524 -13493 1576 -13455
rect 1524 -13527 1534 -13493
rect 1568 -13527 1576 -13493
rect 1524 -13565 1576 -13527
rect 1722 -13500 1774 -13455
rect 1722 -13534 1730 -13500
rect 1764 -13534 1774 -13500
rect 1722 -13565 1774 -13534
rect 2352 -13500 2404 -13455
rect 2352 -13534 2362 -13500
rect 2396 -13534 2404 -13500
rect 2352 -13565 2404 -13534
rect 2550 -13493 2602 -13455
rect 2550 -13527 2558 -13493
rect 2592 -13527 2602 -13493
rect 2550 -13565 2602 -13527
rect 2812 -13493 2864 -13455
rect 2812 -13527 2822 -13493
rect 2856 -13527 2864 -13493
rect 2812 -13565 2864 -13527
rect 3126 -13481 3176 -13435
rect 3010 -13508 3081 -13481
rect 3010 -13542 3033 -13508
rect 3067 -13542 3081 -13508
rect 3010 -13565 3081 -13542
rect 3111 -13508 3176 -13481
rect 3111 -13542 3131 -13508
rect 3165 -13542 3176 -13508
rect 3111 -13565 3176 -13542
rect 3276 -13508 3329 -13435
rect 3276 -13542 3287 -13508
rect 3321 -13542 3329 -13508
rect 3276 -13565 3329 -13542
rect 3384 -13508 3436 -13435
rect 3384 -13542 3392 -13508
rect 3426 -13542 3436 -13508
rect 3384 -13565 3436 -13542
rect 3536 -13481 3586 -13435
rect 3536 -13508 3608 -13481
rect 3536 -13542 3552 -13508
rect 3586 -13542 3608 -13508
rect 3536 -13565 3608 -13542
rect 3638 -13508 3692 -13481
rect 3638 -13542 3649 -13508
rect 3683 -13542 3692 -13508
rect 3638 -13565 3692 -13542
rect 3838 -13493 3890 -13455
rect 3838 -13527 3846 -13493
rect 3880 -13527 3890 -13493
rect 3838 -13565 3890 -13527
rect 4100 -13493 4152 -13455
rect 4100 -13527 4110 -13493
rect 4144 -13527 4152 -13493
rect 4100 -13565 4152 -13527
rect 4298 -13500 4350 -13455
rect 4298 -13534 4306 -13500
rect 4340 -13534 4350 -13500
rect 4298 -13565 4350 -13534
rect 4928 -13500 4980 -13455
rect 4928 -13534 4938 -13500
rect 4972 -13534 4980 -13500
rect 4928 -13565 4980 -13534
rect 5126 -13493 5178 -13455
rect 5126 -13527 5134 -13493
rect 5168 -13527 5178 -13493
rect 5126 -13565 5178 -13527
rect 5388 -13493 5440 -13455
rect 5388 -13527 5398 -13493
rect 5432 -13527 5440 -13493
rect 5388 -13565 5440 -13527
rect 5702 -13481 5752 -13435
rect 5586 -13508 5657 -13481
rect 5586 -13542 5609 -13508
rect 5643 -13542 5657 -13508
rect 5586 -13565 5657 -13542
rect 5687 -13508 5752 -13481
rect 5687 -13542 5707 -13508
rect 5741 -13542 5752 -13508
rect 5687 -13565 5752 -13542
rect 5852 -13508 5905 -13435
rect 5852 -13542 5863 -13508
rect 5897 -13542 5905 -13508
rect 5852 -13565 5905 -13542
rect 5960 -13508 6012 -13435
rect 5960 -13542 5968 -13508
rect 6002 -13542 6012 -13508
rect 5960 -13565 6012 -13542
rect 6112 -13481 6162 -13435
rect 6112 -13508 6184 -13481
rect 6112 -13542 6128 -13508
rect 6162 -13542 6184 -13508
rect 6112 -13565 6184 -13542
rect 6214 -13508 6268 -13481
rect 6214 -13542 6225 -13508
rect 6259 -13542 6268 -13508
rect 6214 -13565 6268 -13542
rect 6414 -13493 6466 -13455
rect 6414 -13527 6422 -13493
rect 6456 -13527 6466 -13493
rect 6414 -13565 6466 -13527
rect 6676 -13493 6728 -13455
rect 6676 -13527 6686 -13493
rect 6720 -13527 6728 -13493
rect 6676 -13565 6728 -13527
rect 6874 -13500 6926 -13455
rect 6874 -13534 6882 -13500
rect 6916 -13534 6926 -13500
rect 6874 -13565 6926 -13534
rect 7504 -13500 7556 -13455
rect 7504 -13534 7514 -13500
rect 7548 -13534 7556 -13500
rect 7504 -13565 7556 -13534
rect 7702 -13493 7754 -13455
rect 7702 -13527 7710 -13493
rect 7744 -13527 7754 -13493
rect 7702 -13565 7754 -13527
rect 7964 -13493 8016 -13455
rect 7964 -13527 7974 -13493
rect 8008 -13527 8016 -13493
rect 7964 -13565 8016 -13527
rect 8278 -13481 8328 -13435
rect 8162 -13508 8233 -13481
rect 8162 -13542 8185 -13508
rect 8219 -13542 8233 -13508
rect 8162 -13565 8233 -13542
rect 8263 -13508 8328 -13481
rect 8263 -13542 8283 -13508
rect 8317 -13542 8328 -13508
rect 8263 -13565 8328 -13542
rect 8428 -13508 8481 -13435
rect 8428 -13542 8439 -13508
rect 8473 -13542 8481 -13508
rect 8428 -13565 8481 -13542
rect 8536 -13508 8588 -13435
rect 8536 -13542 8544 -13508
rect 8578 -13542 8588 -13508
rect 8536 -13565 8588 -13542
rect 8688 -13481 8738 -13435
rect 8688 -13508 8760 -13481
rect 8688 -13542 8704 -13508
rect 8738 -13542 8760 -13508
rect 8688 -13565 8760 -13542
rect 8790 -13508 8844 -13481
rect 8790 -13542 8801 -13508
rect 8835 -13542 8844 -13508
rect 8790 -13565 8844 -13542
rect 8990 -13493 9042 -13455
rect 8990 -13527 8998 -13493
rect 9032 -13527 9042 -13493
rect 8990 -13565 9042 -13527
rect 9252 -13493 9304 -13455
rect 9252 -13527 9262 -13493
rect 9296 -13527 9304 -13493
rect 9252 -13565 9304 -13527
rect 9450 -13500 9502 -13455
rect 9450 -13534 9458 -13500
rect 9492 -13534 9502 -13500
rect 9450 -13565 9502 -13534
rect 10080 -13500 10132 -13455
rect 10080 -13534 10090 -13500
rect 10124 -13534 10132 -13500
rect 10080 -13565 10132 -13534
rect 10370 -13493 10422 -13455
rect 10370 -13527 10378 -13493
rect 10412 -13527 10422 -13493
rect 10370 -13565 10422 -13527
rect 10632 -13493 10684 -13455
rect 10854 -13481 10904 -13435
rect 10632 -13527 10642 -13493
rect 10676 -13527 10684 -13493
rect 10632 -13565 10684 -13527
rect 10738 -13508 10809 -13481
rect 10738 -13542 10761 -13508
rect 10795 -13542 10809 -13508
rect 10738 -13565 10809 -13542
rect 10839 -13508 10904 -13481
rect 10839 -13542 10859 -13508
rect 10893 -13542 10904 -13508
rect 10839 -13565 10904 -13542
rect 11004 -13508 11057 -13435
rect 11004 -13542 11015 -13508
rect 11049 -13542 11057 -13508
rect 11004 -13565 11057 -13542
rect 11112 -13508 11164 -13435
rect 11112 -13542 11120 -13508
rect 11154 -13542 11164 -13508
rect 11112 -13565 11164 -13542
rect 11264 -13481 11314 -13435
rect 11264 -13508 11336 -13481
rect 11264 -13542 11280 -13508
rect 11314 -13542 11336 -13508
rect 11264 -13565 11336 -13542
rect 11366 -13508 11420 -13481
rect 11366 -13542 11377 -13508
rect 11411 -13542 11420 -13508
rect 11366 -13565 11420 -13542
rect 11658 -13493 11710 -13455
rect 11658 -13527 11666 -13493
rect 11700 -13527 11710 -13493
rect 11658 -13565 11710 -13527
rect 11920 -13493 11972 -13455
rect 11920 -13527 11930 -13493
rect 11964 -13527 11972 -13493
rect 11920 -13565 11972 -13527
rect 13682 -13519 13735 -13481
rect 13682 -13553 13690 -13519
rect 13724 -13553 13735 -13519
rect 13682 -13565 13735 -13553
rect 13765 -13506 13821 -13481
rect 13765 -13540 13776 -13506
rect 13810 -13540 13821 -13506
rect 13765 -13565 13821 -13540
rect 13851 -13506 13907 -13481
rect 13851 -13540 13862 -13506
rect 13896 -13540 13907 -13506
rect 13851 -13565 13907 -13540
rect 13937 -13506 13993 -13481
rect 13937 -13540 13948 -13506
rect 13982 -13540 13993 -13506
rect 13937 -13565 13993 -13540
rect 14023 -13506 14079 -13481
rect 14023 -13540 14034 -13506
rect 14068 -13540 14079 -13506
rect 14023 -13565 14079 -13540
rect 14109 -13506 14165 -13481
rect 14109 -13540 14120 -13506
rect 14154 -13540 14165 -13506
rect 14109 -13565 14165 -13540
rect 14195 -13515 14251 -13481
rect 14195 -13549 14206 -13515
rect 14240 -13549 14251 -13515
rect 14195 -13565 14251 -13549
rect 14281 -13506 14337 -13481
rect 14281 -13540 14292 -13506
rect 14326 -13540 14337 -13506
rect 14281 -13565 14337 -13540
rect 14367 -13515 14423 -13481
rect 14367 -13549 14378 -13515
rect 14412 -13549 14423 -13515
rect 14367 -13565 14423 -13549
rect 14453 -13506 14509 -13481
rect 14453 -13540 14464 -13506
rect 14498 -13540 14509 -13506
rect 14453 -13565 14509 -13540
rect 14539 -13515 14595 -13481
rect 14539 -13549 14550 -13515
rect 14584 -13549 14595 -13515
rect 14539 -13565 14595 -13549
rect 14625 -13506 14681 -13481
rect 14625 -13540 14636 -13506
rect 14670 -13540 14681 -13506
rect 14625 -13565 14681 -13540
rect 14711 -13515 14766 -13481
rect 14711 -13549 14722 -13515
rect 14756 -13549 14766 -13515
rect 14711 -13565 14766 -13549
rect 14796 -13506 14852 -13481
rect 14796 -13540 14807 -13506
rect 14841 -13540 14852 -13506
rect 14796 -13565 14852 -13540
rect 14882 -13515 14938 -13481
rect 14882 -13549 14893 -13515
rect 14927 -13549 14938 -13515
rect 14882 -13565 14938 -13549
rect 14968 -13506 15024 -13481
rect 14968 -13540 14979 -13506
rect 15013 -13540 15024 -13506
rect 14968 -13565 15024 -13540
rect 15054 -13515 15110 -13481
rect 15054 -13549 15065 -13515
rect 15099 -13549 15110 -13515
rect 15054 -13565 15110 -13549
rect 15140 -13506 15196 -13481
rect 15140 -13540 15151 -13506
rect 15185 -13540 15196 -13506
rect 15140 -13565 15196 -13540
rect 15226 -13515 15282 -13481
rect 15226 -13549 15237 -13515
rect 15271 -13549 15282 -13515
rect 15226 -13565 15282 -13549
rect 15312 -13506 15368 -13481
rect 15312 -13540 15323 -13506
rect 15357 -13540 15368 -13506
rect 15312 -13565 15368 -13540
rect 15398 -13515 15451 -13481
rect 15398 -13549 15409 -13515
rect 15443 -13549 15451 -13515
rect 15614 -13500 15666 -13455
rect 15614 -13534 15622 -13500
rect 15656 -13534 15666 -13500
rect 15398 -13565 15451 -13549
rect 15614 -13565 15666 -13534
rect 16612 -13500 16664 -13455
rect 16612 -13534 16622 -13500
rect 16656 -13534 16664 -13500
rect 16612 -13565 16664 -13534
rect -2970 -13690 -2918 -13659
rect -2970 -13724 -2962 -13690
rect -2928 -13724 -2918 -13690
rect -2970 -13769 -2918 -13724
rect -2340 -13690 -2288 -13659
rect -2340 -13724 -2330 -13690
rect -2296 -13724 -2288 -13690
rect -2340 -13769 -2288 -13724
rect -1406 -13697 -1354 -13659
rect -1406 -13731 -1398 -13697
rect -1364 -13731 -1354 -13697
rect -1406 -13769 -1354 -13731
rect -1144 -13697 -1092 -13659
rect -942 -13671 -890 -13659
rect -1144 -13731 -1134 -13697
rect -1100 -13731 -1092 -13697
rect -1144 -13769 -1092 -13731
rect -942 -13705 -934 -13671
rect -900 -13705 -890 -13671
rect -942 -13739 -890 -13705
rect -942 -13773 -934 -13739
rect -900 -13773 -890 -13739
rect -942 -13789 -890 -13773
rect -860 -13789 -806 -13659
rect -776 -13671 -724 -13659
rect -776 -13705 -766 -13671
rect -732 -13705 -724 -13671
rect -776 -13739 -724 -13705
rect -776 -13773 -766 -13739
rect -732 -13773 -724 -13739
rect -776 -13789 -724 -13773
rect -578 -13697 -526 -13659
rect -578 -13731 -570 -13697
rect -536 -13731 -526 -13697
rect -578 -13769 -526 -13731
rect -316 -13697 -264 -13659
rect -37 -13673 29 -13659
rect -316 -13731 -306 -13697
rect -272 -13731 -264 -13697
rect -316 -13769 -264 -13731
rect -37 -13707 -16 -13673
rect 18 -13707 29 -13673
rect -37 -13743 29 -13707
rect 59 -13684 115 -13659
rect 59 -13718 70 -13684
rect 104 -13718 115 -13684
rect 59 -13743 115 -13718
rect 145 -13673 201 -13659
rect 145 -13707 156 -13673
rect 190 -13707 201 -13673
rect 145 -13743 201 -13707
rect 231 -13684 287 -13659
rect 231 -13718 242 -13684
rect 276 -13718 287 -13684
rect 231 -13743 287 -13718
rect 317 -13673 396 -13659
rect 317 -13707 328 -13673
rect 362 -13707 396 -13673
rect 317 -13743 396 -13707
rect 618 -13697 670 -13659
rect 618 -13731 626 -13697
rect 660 -13731 670 -13697
rect 618 -13769 670 -13731
rect 880 -13697 932 -13659
rect 880 -13731 890 -13697
rect 924 -13731 932 -13697
rect 880 -13769 932 -13731
rect 1161 -13682 1213 -13659
rect 1161 -13716 1169 -13682
rect 1203 -13716 1213 -13682
rect 1161 -13743 1213 -13716
rect 1243 -13680 1300 -13659
rect 1243 -13714 1253 -13680
rect 1287 -13714 1300 -13680
rect 1243 -13743 1300 -13714
rect 1446 -13697 1498 -13659
rect 1446 -13731 1454 -13697
rect 1488 -13731 1498 -13697
rect 1446 -13769 1498 -13731
rect 1708 -13697 1760 -13659
rect 1708 -13731 1718 -13697
rect 1752 -13731 1760 -13697
rect 1708 -13769 1760 -13731
rect 1906 -13697 1958 -13659
rect 1906 -13731 1914 -13697
rect 1948 -13731 1958 -13697
rect 1906 -13769 1958 -13731
rect 2168 -13697 2220 -13659
rect 2168 -13731 2178 -13697
rect 2212 -13731 2220 -13697
rect 2168 -13769 2220 -13731
rect 2366 -13682 2420 -13659
rect 2366 -13716 2375 -13682
rect 2409 -13716 2420 -13682
rect 2366 -13743 2420 -13716
rect 2450 -13682 2522 -13659
rect 2450 -13716 2472 -13682
rect 2506 -13716 2522 -13682
rect 2450 -13743 2522 -13716
rect 2472 -13789 2522 -13743
rect 2622 -13682 2674 -13659
rect 2622 -13716 2632 -13682
rect 2666 -13716 2674 -13682
rect 2622 -13789 2674 -13716
rect 2729 -13682 2782 -13659
rect 2729 -13716 2737 -13682
rect 2771 -13716 2782 -13682
rect 2729 -13789 2782 -13716
rect 2882 -13682 2947 -13659
rect 2882 -13716 2893 -13682
rect 2927 -13716 2947 -13682
rect 2882 -13743 2947 -13716
rect 2977 -13682 3048 -13659
rect 2977 -13716 2991 -13682
rect 3025 -13716 3048 -13682
rect 2977 -13743 3048 -13716
rect 2882 -13789 2932 -13743
rect 3194 -13697 3246 -13659
rect 3194 -13731 3202 -13697
rect 3236 -13731 3246 -13697
rect 3194 -13769 3246 -13731
rect 3456 -13697 3508 -13659
rect 3456 -13731 3466 -13697
rect 3500 -13731 3508 -13697
rect 3456 -13769 3508 -13731
rect 4390 -13690 4442 -13659
rect 4390 -13724 4398 -13690
rect 4432 -13724 4442 -13690
rect 4390 -13769 4442 -13724
rect 5388 -13690 5440 -13659
rect 5388 -13724 5398 -13690
rect 5432 -13724 5440 -13690
rect 5388 -13769 5440 -13724
rect 6414 -13697 6466 -13659
rect 6414 -13731 6422 -13697
rect 6456 -13731 6466 -13697
rect 6414 -13769 6466 -13731
rect 6676 -13697 6728 -13659
rect 6676 -13731 6686 -13697
rect 6720 -13731 6728 -13697
rect 6676 -13769 6728 -13731
rect 6874 -13682 6928 -13659
rect 6874 -13716 6883 -13682
rect 6917 -13716 6928 -13682
rect 6874 -13743 6928 -13716
rect 6958 -13682 7030 -13659
rect 6958 -13716 6980 -13682
rect 7014 -13716 7030 -13682
rect 6958 -13743 7030 -13716
rect 6980 -13789 7030 -13743
rect 7130 -13682 7182 -13659
rect 7130 -13716 7140 -13682
rect 7174 -13716 7182 -13682
rect 7130 -13789 7182 -13716
rect 7237 -13682 7290 -13659
rect 7237 -13716 7245 -13682
rect 7279 -13716 7290 -13682
rect 7237 -13789 7290 -13716
rect 7390 -13682 7455 -13659
rect 7390 -13716 7401 -13682
rect 7435 -13716 7455 -13682
rect 7390 -13743 7455 -13716
rect 7485 -13682 7556 -13659
rect 7485 -13716 7499 -13682
rect 7533 -13716 7556 -13682
rect 7485 -13743 7556 -13716
rect 7390 -13789 7440 -13743
rect 7702 -13697 7754 -13659
rect 7702 -13731 7710 -13697
rect 7744 -13731 7754 -13697
rect 7702 -13769 7754 -13731
rect 7964 -13697 8016 -13659
rect 7964 -13731 7974 -13697
rect 8008 -13731 8016 -13697
rect 7964 -13769 8016 -13731
rect 8162 -13682 8216 -13659
rect 8162 -13716 8171 -13682
rect 8205 -13716 8216 -13682
rect 8162 -13743 8216 -13716
rect 8246 -13682 8318 -13659
rect 8246 -13716 8268 -13682
rect 8302 -13716 8318 -13682
rect 8246 -13743 8318 -13716
rect 8268 -13789 8318 -13743
rect 8418 -13682 8470 -13659
rect 8418 -13716 8428 -13682
rect 8462 -13716 8470 -13682
rect 8418 -13789 8470 -13716
rect 8525 -13682 8578 -13659
rect 8525 -13716 8533 -13682
rect 8567 -13716 8578 -13682
rect 8525 -13789 8578 -13716
rect 8678 -13682 8743 -13659
rect 8678 -13716 8689 -13682
rect 8723 -13716 8743 -13682
rect 8678 -13743 8743 -13716
rect 8773 -13682 8844 -13659
rect 8773 -13716 8787 -13682
rect 8821 -13716 8844 -13682
rect 8773 -13743 8844 -13716
rect 8678 -13789 8728 -13743
rect 8990 -13697 9042 -13659
rect 8990 -13731 8998 -13697
rect 9032 -13731 9042 -13697
rect 8990 -13769 9042 -13731
rect 9252 -13697 9304 -13659
rect 9252 -13731 9262 -13697
rect 9296 -13731 9304 -13697
rect 9252 -13769 9304 -13731
rect 9450 -13682 9504 -13659
rect 9450 -13716 9459 -13682
rect 9493 -13716 9504 -13682
rect 9450 -13743 9504 -13716
rect 9534 -13682 9606 -13659
rect 9534 -13716 9556 -13682
rect 9590 -13716 9606 -13682
rect 9534 -13743 9606 -13716
rect 9556 -13789 9606 -13743
rect 9706 -13682 9758 -13659
rect 9706 -13716 9716 -13682
rect 9750 -13716 9758 -13682
rect 9706 -13789 9758 -13716
rect 9813 -13682 9866 -13659
rect 9813 -13716 9821 -13682
rect 9855 -13716 9866 -13682
rect 9813 -13789 9866 -13716
rect 9966 -13682 10031 -13659
rect 9966 -13716 9977 -13682
rect 10011 -13716 10031 -13682
rect 9966 -13743 10031 -13716
rect 10061 -13682 10132 -13659
rect 10061 -13716 10075 -13682
rect 10109 -13716 10132 -13682
rect 10061 -13743 10132 -13716
rect 9966 -13789 10016 -13743
rect 10278 -13697 10330 -13659
rect 10278 -13731 10286 -13697
rect 10320 -13731 10330 -13697
rect 10278 -13769 10330 -13731
rect 10540 -13697 10592 -13659
rect 10738 -13671 10790 -13659
rect 10540 -13731 10550 -13697
rect 10584 -13731 10592 -13697
rect 10540 -13769 10592 -13731
rect 10738 -13705 10746 -13671
rect 10780 -13705 10790 -13671
rect 10738 -13739 10790 -13705
rect 10738 -13773 10746 -13739
rect 10780 -13773 10790 -13739
rect 10738 -13789 10790 -13773
rect 10820 -13671 10874 -13659
rect 10820 -13705 10830 -13671
rect 10864 -13705 10874 -13671
rect 10820 -13789 10874 -13705
rect 10904 -13671 10958 -13659
rect 10904 -13705 10914 -13671
rect 10948 -13705 10958 -13671
rect 10904 -13739 10958 -13705
rect 10904 -13773 10914 -13739
rect 10948 -13773 10958 -13739
rect 10904 -13789 10958 -13773
rect 10988 -13671 11042 -13659
rect 10988 -13705 10998 -13671
rect 11032 -13705 11042 -13671
rect 10988 -13789 11042 -13705
rect 11072 -13671 11126 -13659
rect 11072 -13705 11082 -13671
rect 11116 -13705 11126 -13671
rect 11072 -13739 11126 -13705
rect 11072 -13773 11082 -13739
rect 11116 -13773 11126 -13739
rect 11072 -13789 11126 -13773
rect 11156 -13739 11210 -13659
rect 11156 -13773 11166 -13739
rect 11200 -13773 11210 -13739
rect 11156 -13789 11210 -13773
rect 11240 -13671 11294 -13659
rect 11240 -13705 11250 -13671
rect 11284 -13705 11294 -13671
rect 11240 -13789 11294 -13705
rect 11324 -13739 11378 -13659
rect 11324 -13773 11334 -13739
rect 11368 -13773 11378 -13739
rect 11324 -13789 11378 -13773
rect 11408 -13671 11460 -13659
rect 11408 -13705 11418 -13671
rect 11452 -13705 11460 -13671
rect 11408 -13739 11460 -13705
rect 11408 -13773 11418 -13739
rect 11452 -13773 11460 -13739
rect 11408 -13789 11460 -13773
rect 11658 -13697 11710 -13659
rect 11658 -13731 11666 -13697
rect 11700 -13731 11710 -13697
rect 11658 -13769 11710 -13731
rect 11920 -13697 11972 -13659
rect 11920 -13731 11930 -13697
rect 11964 -13731 11972 -13697
rect 11920 -13769 11972 -13731
rect 13590 -13690 13642 -13659
rect 13590 -13724 13598 -13690
rect 13632 -13724 13642 -13690
rect 13590 -13769 13642 -13724
rect 14588 -13690 14640 -13659
rect 14588 -13724 14598 -13690
rect 14632 -13724 14640 -13690
rect 14588 -13769 14640 -13724
rect 14786 -13690 14838 -13659
rect 14786 -13724 14794 -13690
rect 14828 -13724 14838 -13690
rect 14786 -13769 14838 -13724
rect 15784 -13690 15836 -13659
rect 15784 -13724 15794 -13690
rect 15828 -13724 15836 -13690
rect 15784 -13769 15836 -13724
rect 15982 -13690 16034 -13659
rect 15982 -13724 15990 -13690
rect 16024 -13724 16034 -13690
rect 15982 -13769 16034 -13724
rect 16612 -13690 16664 -13659
rect 16612 -13724 16622 -13690
rect 16656 -13724 16664 -13690
rect 16612 -13769 16664 -13724
<< pdiff >>
rect -2970 -71 -2918 -59
rect -2970 -105 -2962 -71
rect -2928 -105 -2918 -71
rect -2970 -173 -2918 -105
rect -2970 -207 -2962 -173
rect -2928 -207 -2918 -173
rect -2970 -233 -2918 -207
rect -2340 -71 -2288 -59
rect -2340 -105 -2330 -71
rect -2296 -105 -2288 -71
rect -1406 -71 -1354 -59
rect -2340 -173 -2288 -105
rect -2340 -207 -2330 -173
rect -2296 -207 -2288 -173
rect -2340 -233 -2288 -207
rect -1406 -105 -1398 -71
rect -1364 -105 -1354 -71
rect -1406 -173 -1354 -105
rect -1406 -207 -1398 -173
rect -1364 -207 -1354 -173
rect -1406 -233 -1354 -207
rect -1144 -71 -1092 -59
rect -1144 -105 -1134 -71
rect -1100 -105 -1092 -71
rect -942 -71 -890 -59
rect -1144 -173 -1092 -105
rect -1144 -207 -1134 -173
rect -1100 -207 -1092 -173
rect -1144 -233 -1092 -207
rect -942 -105 -934 -71
rect -900 -105 -890 -71
rect -942 -139 -890 -105
rect -942 -173 -934 -139
rect -900 -173 -890 -139
rect -942 -207 -890 -173
rect -942 -241 -934 -207
rect -900 -241 -890 -207
rect -942 -259 -890 -241
rect -860 -71 -806 -59
rect -860 -105 -850 -71
rect -816 -105 -806 -71
rect -860 -139 -806 -105
rect -860 -173 -850 -139
rect -816 -173 -806 -139
rect -860 -207 -806 -173
rect -860 -241 -850 -207
rect -816 -241 -806 -207
rect -860 -259 -806 -241
rect -776 -71 -724 -59
rect -776 -105 -766 -71
rect -732 -105 -724 -71
rect -578 -71 -526 -59
rect -776 -139 -724 -105
rect -776 -173 -766 -139
rect -732 -173 -724 -139
rect -776 -207 -724 -173
rect -776 -241 -766 -207
rect -732 -241 -724 -207
rect -776 -259 -724 -241
rect -578 -105 -570 -71
rect -536 -105 -526 -71
rect -578 -173 -526 -105
rect -578 -207 -570 -173
rect -536 -207 -526 -173
rect -578 -233 -526 -207
rect -316 -71 -264 -59
rect -316 -105 -306 -71
rect -272 -105 -264 -71
rect -316 -173 -264 -105
rect -316 -207 -306 -173
rect -272 -207 -264 -173
rect -316 -233 -264 -207
rect -118 -78 -57 -59
rect -118 -112 -102 -78
rect -68 -112 -57 -78
rect -118 -146 -57 -112
rect -118 -180 -102 -146
rect -68 -180 -57 -146
rect -118 -259 -57 -180
rect -27 -85 29 -59
rect -27 -119 -16 -85
rect 18 -119 29 -85
rect -27 -173 29 -119
rect -27 -207 -16 -173
rect 18 -207 29 -173
rect -27 -259 29 -207
rect 59 -78 115 -59
rect 59 -112 70 -78
rect 104 -112 115 -78
rect 59 -146 115 -112
rect 59 -180 70 -146
rect 104 -180 115 -146
rect 59 -259 115 -180
rect 145 -85 201 -59
rect 145 -119 156 -85
rect 190 -119 201 -85
rect 145 -173 201 -119
rect 145 -207 156 -173
rect 190 -207 201 -173
rect 145 -259 201 -207
rect 231 -78 287 -59
rect 231 -112 242 -78
rect 276 -112 287 -78
rect 231 -146 287 -112
rect 231 -180 242 -146
rect 276 -180 287 -146
rect 231 -259 287 -180
rect 317 -85 373 -59
rect 317 -119 328 -85
rect 362 -119 373 -85
rect 317 -173 373 -119
rect 317 -207 328 -173
rect 362 -207 373 -173
rect 317 -259 373 -207
rect 403 -78 472 -59
rect 618 -71 670 -59
rect 403 -112 414 -78
rect 448 -112 472 -78
rect 403 -146 472 -112
rect 403 -180 414 -146
rect 448 -180 472 -146
rect 403 -259 472 -180
rect 618 -105 626 -71
rect 660 -105 670 -71
rect 618 -173 670 -105
rect 618 -207 626 -173
rect 660 -207 670 -173
rect 618 -233 670 -207
rect 880 -71 932 -59
rect 880 -105 890 -71
rect 924 -105 932 -71
rect 1078 -71 1130 -59
rect 880 -173 932 -105
rect 880 -207 890 -173
rect 924 -207 932 -173
rect 880 -233 932 -207
rect 1078 -105 1086 -71
rect 1120 -105 1130 -71
rect 1078 -173 1130 -105
rect 1078 -207 1086 -173
rect 1120 -207 1130 -173
rect 1078 -227 1130 -207
rect 1160 -71 1214 -59
rect 1160 -105 1170 -71
rect 1204 -105 1214 -71
rect 1160 -173 1214 -105
rect 1160 -207 1170 -173
rect 1204 -207 1214 -173
rect 1160 -227 1214 -207
rect 1244 -71 1300 -59
rect 1244 -105 1254 -71
rect 1288 -105 1300 -71
rect 1446 -71 1498 -59
rect 1244 -173 1300 -105
rect 1244 -207 1254 -173
rect 1288 -207 1300 -173
rect 1244 -227 1300 -207
rect 1446 -105 1454 -71
rect 1488 -105 1498 -71
rect 1446 -173 1498 -105
rect 1446 -207 1454 -173
rect 1488 -207 1498 -173
rect 1446 -233 1498 -207
rect 1708 -71 1760 -59
rect 1708 -105 1718 -71
rect 1752 -105 1760 -71
rect 1906 -71 1958 -59
rect 1708 -173 1760 -105
rect 1708 -207 1718 -173
rect 1752 -207 1760 -173
rect 1708 -233 1760 -207
rect 1906 -105 1914 -71
rect 1948 -105 1958 -71
rect 1906 -173 1958 -105
rect 1906 -207 1914 -173
rect 1948 -207 1958 -173
rect 1906 -233 1958 -207
rect 2168 -71 2220 -59
rect 2168 -105 2178 -71
rect 2212 -105 2220 -71
rect 2168 -173 2220 -105
rect 2168 -207 2178 -173
rect 2212 -207 2220 -173
rect 2168 -233 2220 -207
rect 2366 -78 2420 -59
rect 2366 -112 2375 -78
rect 2409 -112 2420 -78
rect 2366 -146 2420 -112
rect 2366 -180 2375 -146
rect 2409 -180 2420 -146
rect 2366 -259 2420 -180
rect 2450 -78 2522 -59
rect 2450 -112 2475 -78
rect 2509 -112 2522 -78
rect 2450 -146 2522 -112
rect 2450 -180 2475 -146
rect 2509 -180 2522 -146
rect 2450 -223 2522 -180
rect 2622 -78 2675 -59
rect 2622 -112 2633 -78
rect 2667 -112 2675 -78
rect 2622 -146 2675 -112
rect 2622 -180 2633 -146
rect 2667 -180 2675 -146
rect 2622 -223 2675 -180
rect 2729 -79 2782 -59
rect 2729 -113 2737 -79
rect 2771 -113 2782 -79
rect 2729 -147 2782 -113
rect 2729 -181 2737 -147
rect 2771 -181 2782 -147
rect 2729 -223 2782 -181
rect 2882 -78 2947 -59
rect 2882 -112 2893 -78
rect 2927 -112 2947 -78
rect 2882 -146 2947 -112
rect 2882 -180 2893 -146
rect 2927 -180 2947 -146
rect 2882 -223 2947 -180
rect 2450 -259 2500 -223
rect 2897 -259 2947 -223
rect 2977 -79 3048 -59
rect 3194 -71 3246 -59
rect 2977 -113 2991 -79
rect 3025 -113 3048 -79
rect 2977 -147 3048 -113
rect 2977 -181 2991 -147
rect 3025 -181 3048 -147
rect 2977 -259 3048 -181
rect 3194 -105 3202 -71
rect 3236 -105 3246 -71
rect 3194 -173 3246 -105
rect 3194 -207 3202 -173
rect 3236 -207 3246 -173
rect 3194 -233 3246 -207
rect 3456 -71 3508 -59
rect 3456 -105 3466 -71
rect 3500 -105 3508 -71
rect 4390 -71 4442 -59
rect 3456 -173 3508 -105
rect 3456 -207 3466 -173
rect 3500 -207 3508 -173
rect 3456 -233 3508 -207
rect 4390 -105 4398 -71
rect 4432 -105 4442 -71
rect 4390 -173 4442 -105
rect 4390 -207 4398 -173
rect 4432 -207 4442 -173
rect 4390 -233 4442 -207
rect 5388 -71 5440 -59
rect 5388 -105 5398 -71
rect 5432 -105 5440 -71
rect 6414 -71 6466 -59
rect 5388 -173 5440 -105
rect 5388 -207 5398 -173
rect 5432 -207 5440 -173
rect 5388 -233 5440 -207
rect 6414 -105 6422 -71
rect 6456 -105 6466 -71
rect 6414 -173 6466 -105
rect 6414 -207 6422 -173
rect 6456 -207 6466 -173
rect 6414 -233 6466 -207
rect 6676 -71 6728 -59
rect 6676 -105 6686 -71
rect 6720 -105 6728 -71
rect 6676 -173 6728 -105
rect 6676 -207 6686 -173
rect 6720 -207 6728 -173
rect 6676 -233 6728 -207
rect 6874 -78 6928 -59
rect 6874 -112 6883 -78
rect 6917 -112 6928 -78
rect 6874 -146 6928 -112
rect 6874 -180 6883 -146
rect 6917 -180 6928 -146
rect 6874 -259 6928 -180
rect 6958 -78 7030 -59
rect 6958 -112 6983 -78
rect 7017 -112 7030 -78
rect 6958 -146 7030 -112
rect 6958 -180 6983 -146
rect 7017 -180 7030 -146
rect 6958 -223 7030 -180
rect 7130 -78 7183 -59
rect 7130 -112 7141 -78
rect 7175 -112 7183 -78
rect 7130 -146 7183 -112
rect 7130 -180 7141 -146
rect 7175 -180 7183 -146
rect 7130 -223 7183 -180
rect 7237 -79 7290 -59
rect 7237 -113 7245 -79
rect 7279 -113 7290 -79
rect 7237 -147 7290 -113
rect 7237 -181 7245 -147
rect 7279 -181 7290 -147
rect 7237 -223 7290 -181
rect 7390 -78 7455 -59
rect 7390 -112 7401 -78
rect 7435 -112 7455 -78
rect 7390 -146 7455 -112
rect 7390 -180 7401 -146
rect 7435 -180 7455 -146
rect 7390 -223 7455 -180
rect 6958 -259 7008 -223
rect 7405 -259 7455 -223
rect 7485 -79 7556 -59
rect 7702 -71 7754 -59
rect 7485 -113 7499 -79
rect 7533 -113 7556 -79
rect 7485 -147 7556 -113
rect 7485 -181 7499 -147
rect 7533 -181 7556 -147
rect 7485 -259 7556 -181
rect 7702 -105 7710 -71
rect 7744 -105 7754 -71
rect 7702 -173 7754 -105
rect 7702 -207 7710 -173
rect 7744 -207 7754 -173
rect 7702 -233 7754 -207
rect 7964 -71 8016 -59
rect 7964 -105 7974 -71
rect 8008 -105 8016 -71
rect 7964 -173 8016 -105
rect 7964 -207 7974 -173
rect 8008 -207 8016 -173
rect 7964 -233 8016 -207
rect 8162 -78 8216 -59
rect 8162 -112 8171 -78
rect 8205 -112 8216 -78
rect 8162 -146 8216 -112
rect 8162 -180 8171 -146
rect 8205 -180 8216 -146
rect 8162 -259 8216 -180
rect 8246 -78 8318 -59
rect 8246 -112 8271 -78
rect 8305 -112 8318 -78
rect 8246 -146 8318 -112
rect 8246 -180 8271 -146
rect 8305 -180 8318 -146
rect 8246 -223 8318 -180
rect 8418 -78 8471 -59
rect 8418 -112 8429 -78
rect 8463 -112 8471 -78
rect 8418 -146 8471 -112
rect 8418 -180 8429 -146
rect 8463 -180 8471 -146
rect 8418 -223 8471 -180
rect 8525 -79 8578 -59
rect 8525 -113 8533 -79
rect 8567 -113 8578 -79
rect 8525 -147 8578 -113
rect 8525 -181 8533 -147
rect 8567 -181 8578 -147
rect 8525 -223 8578 -181
rect 8678 -78 8743 -59
rect 8678 -112 8689 -78
rect 8723 -112 8743 -78
rect 8678 -146 8743 -112
rect 8678 -180 8689 -146
rect 8723 -180 8743 -146
rect 8678 -223 8743 -180
rect 8246 -259 8296 -223
rect 8693 -259 8743 -223
rect 8773 -79 8844 -59
rect 8990 -71 9042 -59
rect 8773 -113 8787 -79
rect 8821 -113 8844 -79
rect 8773 -147 8844 -113
rect 8773 -181 8787 -147
rect 8821 -181 8844 -147
rect 8773 -259 8844 -181
rect 8990 -105 8998 -71
rect 9032 -105 9042 -71
rect 8990 -173 9042 -105
rect 8990 -207 8998 -173
rect 9032 -207 9042 -173
rect 8990 -233 9042 -207
rect 9252 -71 9304 -59
rect 9252 -105 9262 -71
rect 9296 -105 9304 -71
rect 9252 -173 9304 -105
rect 9252 -207 9262 -173
rect 9296 -207 9304 -173
rect 9252 -233 9304 -207
rect 9450 -78 9504 -59
rect 9450 -112 9459 -78
rect 9493 -112 9504 -78
rect 9450 -146 9504 -112
rect 9450 -180 9459 -146
rect 9493 -180 9504 -146
rect 9450 -259 9504 -180
rect 9534 -78 9606 -59
rect 9534 -112 9559 -78
rect 9593 -112 9606 -78
rect 9534 -146 9606 -112
rect 9534 -180 9559 -146
rect 9593 -180 9606 -146
rect 9534 -223 9606 -180
rect 9706 -78 9759 -59
rect 9706 -112 9717 -78
rect 9751 -112 9759 -78
rect 9706 -146 9759 -112
rect 9706 -180 9717 -146
rect 9751 -180 9759 -146
rect 9706 -223 9759 -180
rect 9813 -79 9866 -59
rect 9813 -113 9821 -79
rect 9855 -113 9866 -79
rect 9813 -147 9866 -113
rect 9813 -181 9821 -147
rect 9855 -181 9866 -147
rect 9813 -223 9866 -181
rect 9966 -78 10031 -59
rect 9966 -112 9977 -78
rect 10011 -112 10031 -78
rect 9966 -146 10031 -112
rect 9966 -180 9977 -146
rect 10011 -180 10031 -146
rect 9966 -223 10031 -180
rect 9534 -259 9584 -223
rect 9981 -259 10031 -223
rect 10061 -79 10132 -59
rect 10278 -71 10330 -59
rect 10061 -113 10075 -79
rect 10109 -113 10132 -79
rect 10061 -147 10132 -113
rect 10061 -181 10075 -147
rect 10109 -181 10132 -147
rect 10061 -259 10132 -181
rect 10278 -105 10286 -71
rect 10320 -105 10330 -71
rect 10278 -173 10330 -105
rect 10278 -207 10286 -173
rect 10320 -207 10330 -173
rect 10278 -233 10330 -207
rect 10540 -71 10592 -59
rect 10540 -105 10550 -71
rect 10584 -105 10592 -71
rect 10738 -71 10790 -59
rect 10540 -173 10592 -105
rect 10540 -207 10550 -173
rect 10584 -207 10592 -173
rect 10540 -233 10592 -207
rect 10738 -105 10746 -71
rect 10780 -105 10790 -71
rect 10738 -139 10790 -105
rect 10738 -173 10746 -139
rect 10780 -173 10790 -139
rect 10738 -207 10790 -173
rect 10738 -241 10746 -207
rect 10780 -241 10790 -207
rect 10738 -259 10790 -241
rect 10820 -71 10874 -59
rect 10820 -105 10830 -71
rect 10864 -105 10874 -71
rect 10820 -139 10874 -105
rect 10820 -173 10830 -139
rect 10864 -173 10874 -139
rect 10820 -207 10874 -173
rect 10820 -241 10830 -207
rect 10864 -241 10874 -207
rect 10820 -259 10874 -241
rect 10904 -71 10958 -59
rect 10904 -105 10914 -71
rect 10948 -105 10958 -71
rect 10904 -139 10958 -105
rect 10904 -173 10914 -139
rect 10948 -173 10958 -139
rect 10904 -259 10958 -173
rect 10988 -71 11042 -59
rect 10988 -105 10998 -71
rect 11032 -105 11042 -71
rect 10988 -139 11042 -105
rect 10988 -173 10998 -139
rect 11032 -173 11042 -139
rect 10988 -207 11042 -173
rect 10988 -241 10998 -207
rect 11032 -241 11042 -207
rect 10988 -259 11042 -241
rect 11072 -71 11126 -59
rect 11072 -105 11082 -71
rect 11116 -105 11126 -71
rect 11072 -139 11126 -105
rect 11072 -173 11082 -139
rect 11116 -173 11126 -139
rect 11072 -259 11126 -173
rect 11156 -71 11210 -59
rect 11156 -105 11166 -71
rect 11200 -105 11210 -71
rect 11156 -139 11210 -105
rect 11156 -173 11166 -139
rect 11200 -173 11210 -139
rect 11156 -207 11210 -173
rect 11156 -241 11166 -207
rect 11200 -241 11210 -207
rect 11156 -259 11210 -241
rect 11240 -71 11294 -59
rect 11240 -105 11250 -71
rect 11284 -105 11294 -71
rect 11240 -139 11294 -105
rect 11240 -173 11250 -139
rect 11284 -173 11294 -139
rect 11240 -259 11294 -173
rect 11324 -71 11378 -59
rect 11324 -105 11334 -71
rect 11368 -105 11378 -71
rect 11324 -139 11378 -105
rect 11324 -173 11334 -139
rect 11368 -173 11378 -139
rect 11324 -207 11378 -173
rect 11324 -241 11334 -207
rect 11368 -241 11378 -207
rect 11324 -259 11378 -241
rect 11408 -71 11460 -59
rect 11408 -105 11418 -71
rect 11452 -105 11460 -71
rect 11658 -71 11710 -59
rect 11408 -139 11460 -105
rect 11408 -173 11418 -139
rect 11452 -173 11460 -139
rect 11408 -259 11460 -173
rect 11658 -105 11666 -71
rect 11700 -105 11710 -71
rect 11658 -173 11710 -105
rect 11658 -207 11666 -173
rect 11700 -207 11710 -173
rect 11658 -233 11710 -207
rect 11920 -71 11972 -59
rect 11920 -105 11930 -71
rect 11964 -105 11972 -71
rect 13590 -71 13642 -59
rect 11920 -173 11972 -105
rect 11920 -207 11930 -173
rect 11964 -207 11972 -173
rect 11920 -233 11972 -207
rect 13590 -105 13598 -71
rect 13632 -105 13642 -71
rect 13590 -173 13642 -105
rect 13590 -207 13598 -173
rect 13632 -207 13642 -173
rect 13590 -233 13642 -207
rect 14588 -71 14640 -59
rect 14588 -105 14598 -71
rect 14632 -105 14640 -71
rect 14786 -71 14838 -59
rect 14588 -173 14640 -105
rect 14588 -207 14598 -173
rect 14632 -207 14640 -173
rect 14588 -233 14640 -207
rect 14786 -105 14794 -71
rect 14828 -105 14838 -71
rect 14786 -173 14838 -105
rect 14786 -207 14794 -173
rect 14828 -207 14838 -173
rect 14786 -233 14838 -207
rect 15784 -71 15836 -59
rect 15784 -105 15794 -71
rect 15828 -105 15836 -71
rect 15982 -71 16034 -59
rect 15784 -173 15836 -105
rect 15784 -207 15794 -173
rect 15828 -207 15836 -173
rect 15784 -233 15836 -207
rect 15982 -105 15990 -71
rect 16024 -105 16034 -71
rect 15982 -173 16034 -105
rect 15982 -207 15990 -173
rect 16024 -207 16034 -173
rect 15982 -233 16034 -207
rect 16612 -71 16664 -59
rect 16612 -105 16622 -71
rect 16656 -105 16664 -71
rect 16612 -173 16664 -105
rect 16612 -207 16622 -173
rect 16656 -207 16664 -173
rect 16612 -233 16664 -207
rect -2970 -905 -2918 -879
rect -2970 -939 -2962 -905
rect -2928 -939 -2918 -905
rect -2970 -1007 -2918 -939
rect -2970 -1041 -2962 -1007
rect -2928 -1041 -2918 -1007
rect -2970 -1053 -2918 -1041
rect -2340 -905 -2288 -879
rect -2340 -939 -2330 -905
rect -2296 -939 -2288 -905
rect -2340 -1007 -2288 -939
rect -2340 -1041 -2330 -1007
rect -2296 -1041 -2288 -1007
rect -1590 -905 -1538 -879
rect -1590 -939 -1582 -905
rect -1548 -939 -1538 -905
rect -1590 -1007 -1538 -939
rect -2340 -1053 -2288 -1041
rect -1590 -1041 -1582 -1007
rect -1548 -1041 -1538 -1007
rect -1590 -1053 -1538 -1041
rect -960 -905 -908 -879
rect -960 -939 -950 -905
rect -916 -939 -908 -905
rect -960 -1007 -908 -939
rect -960 -1041 -950 -1007
rect -916 -1041 -908 -1007
rect -960 -1053 -908 -1041
rect -854 -905 -802 -879
rect -854 -939 -846 -905
rect -812 -939 -802 -905
rect -854 -1007 -802 -939
rect -854 -1041 -846 -1007
rect -812 -1041 -802 -1007
rect -854 -1053 -802 -1041
rect -224 -905 -172 -879
rect -224 -939 -214 -905
rect -180 -939 -172 -905
rect -224 -1007 -172 -939
rect -224 -1041 -214 -1007
rect -180 -1041 -172 -1007
rect -26 -905 26 -879
rect -26 -939 -18 -905
rect 16 -939 26 -905
rect -26 -1007 26 -939
rect -224 -1053 -172 -1041
rect -26 -1041 -18 -1007
rect 16 -1041 26 -1007
rect -26 -1053 26 -1041
rect 236 -905 288 -879
rect 236 -939 246 -905
rect 280 -939 288 -905
rect 236 -1007 288 -939
rect 236 -1041 246 -1007
rect 280 -1041 288 -1007
rect 434 -931 505 -853
rect 434 -965 457 -931
rect 491 -965 505 -931
rect 434 -999 505 -965
rect 434 -1033 457 -999
rect 491 -1033 505 -999
rect 236 -1053 288 -1041
rect 434 -1053 505 -1033
rect 535 -889 585 -853
rect 982 -889 1032 -853
rect 535 -932 600 -889
rect 535 -966 555 -932
rect 589 -966 600 -932
rect 535 -1000 600 -966
rect 535 -1034 555 -1000
rect 589 -1034 600 -1000
rect 535 -1053 600 -1034
rect 700 -931 753 -889
rect 700 -965 711 -931
rect 745 -965 753 -931
rect 700 -999 753 -965
rect 700 -1033 711 -999
rect 745 -1033 753 -999
rect 700 -1053 753 -1033
rect 807 -932 860 -889
rect 807 -966 815 -932
rect 849 -966 860 -932
rect 807 -1000 860 -966
rect 807 -1034 815 -1000
rect 849 -1034 860 -1000
rect 807 -1053 860 -1034
rect 960 -932 1032 -889
rect 960 -966 973 -932
rect 1007 -966 1032 -932
rect 960 -1000 1032 -966
rect 960 -1034 973 -1000
rect 1007 -1034 1032 -1000
rect 960 -1053 1032 -1034
rect 1062 -932 1116 -853
rect 1062 -966 1073 -932
rect 1107 -966 1116 -932
rect 1062 -1000 1116 -966
rect 1062 -1034 1073 -1000
rect 1107 -1034 1116 -1000
rect 1062 -1053 1116 -1034
rect 1262 -905 1314 -879
rect 1262 -939 1270 -905
rect 1304 -939 1314 -905
rect 1262 -1007 1314 -939
rect 1262 -1041 1270 -1007
rect 1304 -1041 1314 -1007
rect 1262 -1053 1314 -1041
rect 1524 -905 1576 -879
rect 1524 -939 1534 -905
rect 1568 -939 1576 -905
rect 1524 -1007 1576 -939
rect 1524 -1041 1534 -1007
rect 1568 -1041 1576 -1007
rect 1722 -905 1774 -879
rect 1722 -939 1730 -905
rect 1764 -939 1774 -905
rect 1722 -1007 1774 -939
rect 1524 -1053 1576 -1041
rect 1722 -1041 1730 -1007
rect 1764 -1041 1774 -1007
rect 1722 -1053 1774 -1041
rect 2352 -905 2404 -879
rect 2352 -939 2362 -905
rect 2396 -939 2404 -905
rect 2352 -1007 2404 -939
rect 2352 -1041 2362 -1007
rect 2396 -1041 2404 -1007
rect 2550 -905 2602 -879
rect 2550 -939 2558 -905
rect 2592 -939 2602 -905
rect 2550 -1007 2602 -939
rect 2352 -1053 2404 -1041
rect 2550 -1041 2558 -1007
rect 2592 -1041 2602 -1007
rect 2550 -1053 2602 -1041
rect 2812 -905 2864 -879
rect 2812 -939 2822 -905
rect 2856 -939 2864 -905
rect 2812 -1007 2864 -939
rect 2812 -1041 2822 -1007
rect 2856 -1041 2864 -1007
rect 3010 -931 3081 -853
rect 3010 -965 3033 -931
rect 3067 -965 3081 -931
rect 3010 -999 3081 -965
rect 3010 -1033 3033 -999
rect 3067 -1033 3081 -999
rect 2812 -1053 2864 -1041
rect 3010 -1053 3081 -1033
rect 3111 -889 3161 -853
rect 3558 -889 3608 -853
rect 3111 -932 3176 -889
rect 3111 -966 3131 -932
rect 3165 -966 3176 -932
rect 3111 -1000 3176 -966
rect 3111 -1034 3131 -1000
rect 3165 -1034 3176 -1000
rect 3111 -1053 3176 -1034
rect 3276 -931 3329 -889
rect 3276 -965 3287 -931
rect 3321 -965 3329 -931
rect 3276 -999 3329 -965
rect 3276 -1033 3287 -999
rect 3321 -1033 3329 -999
rect 3276 -1053 3329 -1033
rect 3383 -932 3436 -889
rect 3383 -966 3391 -932
rect 3425 -966 3436 -932
rect 3383 -1000 3436 -966
rect 3383 -1034 3391 -1000
rect 3425 -1034 3436 -1000
rect 3383 -1053 3436 -1034
rect 3536 -932 3608 -889
rect 3536 -966 3549 -932
rect 3583 -966 3608 -932
rect 3536 -1000 3608 -966
rect 3536 -1034 3549 -1000
rect 3583 -1034 3608 -1000
rect 3536 -1053 3608 -1034
rect 3638 -932 3692 -853
rect 3638 -966 3649 -932
rect 3683 -966 3692 -932
rect 3638 -1000 3692 -966
rect 3638 -1034 3649 -1000
rect 3683 -1034 3692 -1000
rect 3638 -1053 3692 -1034
rect 3838 -905 3890 -879
rect 3838 -939 3846 -905
rect 3880 -939 3890 -905
rect 3838 -1007 3890 -939
rect 3838 -1041 3846 -1007
rect 3880 -1041 3890 -1007
rect 3838 -1053 3890 -1041
rect 4100 -905 4152 -879
rect 4100 -939 4110 -905
rect 4144 -939 4152 -905
rect 4100 -1007 4152 -939
rect 4100 -1041 4110 -1007
rect 4144 -1041 4152 -1007
rect 4298 -905 4350 -879
rect 4298 -939 4306 -905
rect 4340 -939 4350 -905
rect 4298 -1007 4350 -939
rect 4100 -1053 4152 -1041
rect 4298 -1041 4306 -1007
rect 4340 -1041 4350 -1007
rect 4298 -1053 4350 -1041
rect 4928 -905 4980 -879
rect 4928 -939 4938 -905
rect 4972 -939 4980 -905
rect 4928 -1007 4980 -939
rect 4928 -1041 4938 -1007
rect 4972 -1041 4980 -1007
rect 5126 -905 5178 -879
rect 5126 -939 5134 -905
rect 5168 -939 5178 -905
rect 5126 -1007 5178 -939
rect 4928 -1053 4980 -1041
rect 5126 -1041 5134 -1007
rect 5168 -1041 5178 -1007
rect 5126 -1053 5178 -1041
rect 5388 -905 5440 -879
rect 5388 -939 5398 -905
rect 5432 -939 5440 -905
rect 5388 -1007 5440 -939
rect 5388 -1041 5398 -1007
rect 5432 -1041 5440 -1007
rect 5586 -931 5657 -853
rect 5586 -965 5609 -931
rect 5643 -965 5657 -931
rect 5586 -999 5657 -965
rect 5586 -1033 5609 -999
rect 5643 -1033 5657 -999
rect 5388 -1053 5440 -1041
rect 5586 -1053 5657 -1033
rect 5687 -889 5737 -853
rect 6134 -889 6184 -853
rect 5687 -932 5752 -889
rect 5687 -966 5707 -932
rect 5741 -966 5752 -932
rect 5687 -1000 5752 -966
rect 5687 -1034 5707 -1000
rect 5741 -1034 5752 -1000
rect 5687 -1053 5752 -1034
rect 5852 -931 5905 -889
rect 5852 -965 5863 -931
rect 5897 -965 5905 -931
rect 5852 -999 5905 -965
rect 5852 -1033 5863 -999
rect 5897 -1033 5905 -999
rect 5852 -1053 5905 -1033
rect 5959 -932 6012 -889
rect 5959 -966 5967 -932
rect 6001 -966 6012 -932
rect 5959 -1000 6012 -966
rect 5959 -1034 5967 -1000
rect 6001 -1034 6012 -1000
rect 5959 -1053 6012 -1034
rect 6112 -932 6184 -889
rect 6112 -966 6125 -932
rect 6159 -966 6184 -932
rect 6112 -1000 6184 -966
rect 6112 -1034 6125 -1000
rect 6159 -1034 6184 -1000
rect 6112 -1053 6184 -1034
rect 6214 -932 6268 -853
rect 6214 -966 6225 -932
rect 6259 -966 6268 -932
rect 6214 -1000 6268 -966
rect 6214 -1034 6225 -1000
rect 6259 -1034 6268 -1000
rect 6214 -1053 6268 -1034
rect 6414 -905 6466 -879
rect 6414 -939 6422 -905
rect 6456 -939 6466 -905
rect 6414 -1007 6466 -939
rect 6414 -1041 6422 -1007
rect 6456 -1041 6466 -1007
rect 6414 -1053 6466 -1041
rect 6676 -905 6728 -879
rect 6676 -939 6686 -905
rect 6720 -939 6728 -905
rect 6676 -1007 6728 -939
rect 6676 -1041 6686 -1007
rect 6720 -1041 6728 -1007
rect 6874 -905 6926 -879
rect 6874 -939 6882 -905
rect 6916 -939 6926 -905
rect 6874 -1007 6926 -939
rect 6676 -1053 6728 -1041
rect 6874 -1041 6882 -1007
rect 6916 -1041 6926 -1007
rect 6874 -1053 6926 -1041
rect 7504 -905 7556 -879
rect 7504 -939 7514 -905
rect 7548 -939 7556 -905
rect 7504 -1007 7556 -939
rect 7504 -1041 7514 -1007
rect 7548 -1041 7556 -1007
rect 7702 -905 7754 -879
rect 7702 -939 7710 -905
rect 7744 -939 7754 -905
rect 7702 -1007 7754 -939
rect 7504 -1053 7556 -1041
rect 7702 -1041 7710 -1007
rect 7744 -1041 7754 -1007
rect 7702 -1053 7754 -1041
rect 7964 -905 8016 -879
rect 7964 -939 7974 -905
rect 8008 -939 8016 -905
rect 7964 -1007 8016 -939
rect 7964 -1041 7974 -1007
rect 8008 -1041 8016 -1007
rect 8162 -931 8233 -853
rect 8162 -965 8185 -931
rect 8219 -965 8233 -931
rect 8162 -999 8233 -965
rect 8162 -1033 8185 -999
rect 8219 -1033 8233 -999
rect 7964 -1053 8016 -1041
rect 8162 -1053 8233 -1033
rect 8263 -889 8313 -853
rect 8710 -889 8760 -853
rect 8263 -932 8328 -889
rect 8263 -966 8283 -932
rect 8317 -966 8328 -932
rect 8263 -1000 8328 -966
rect 8263 -1034 8283 -1000
rect 8317 -1034 8328 -1000
rect 8263 -1053 8328 -1034
rect 8428 -931 8481 -889
rect 8428 -965 8439 -931
rect 8473 -965 8481 -931
rect 8428 -999 8481 -965
rect 8428 -1033 8439 -999
rect 8473 -1033 8481 -999
rect 8428 -1053 8481 -1033
rect 8535 -932 8588 -889
rect 8535 -966 8543 -932
rect 8577 -966 8588 -932
rect 8535 -1000 8588 -966
rect 8535 -1034 8543 -1000
rect 8577 -1034 8588 -1000
rect 8535 -1053 8588 -1034
rect 8688 -932 8760 -889
rect 8688 -966 8701 -932
rect 8735 -966 8760 -932
rect 8688 -1000 8760 -966
rect 8688 -1034 8701 -1000
rect 8735 -1034 8760 -1000
rect 8688 -1053 8760 -1034
rect 8790 -932 8844 -853
rect 8790 -966 8801 -932
rect 8835 -966 8844 -932
rect 8790 -1000 8844 -966
rect 8790 -1034 8801 -1000
rect 8835 -1034 8844 -1000
rect 8790 -1053 8844 -1034
rect 8990 -905 9042 -879
rect 8990 -939 8998 -905
rect 9032 -939 9042 -905
rect 8990 -1007 9042 -939
rect 8990 -1041 8998 -1007
rect 9032 -1041 9042 -1007
rect 8990 -1053 9042 -1041
rect 9252 -905 9304 -879
rect 9252 -939 9262 -905
rect 9296 -939 9304 -905
rect 9252 -1007 9304 -939
rect 9252 -1041 9262 -1007
rect 9296 -1041 9304 -1007
rect 9450 -905 9502 -879
rect 9450 -939 9458 -905
rect 9492 -939 9502 -905
rect 9450 -1007 9502 -939
rect 9252 -1053 9304 -1041
rect 9450 -1041 9458 -1007
rect 9492 -1041 9502 -1007
rect 9450 -1053 9502 -1041
rect 10080 -905 10132 -879
rect 10080 -939 10090 -905
rect 10124 -939 10132 -905
rect 10080 -1007 10132 -939
rect 10080 -1041 10090 -1007
rect 10124 -1041 10132 -1007
rect 10370 -905 10422 -879
rect 10370 -939 10378 -905
rect 10412 -939 10422 -905
rect 10370 -1007 10422 -939
rect 10080 -1053 10132 -1041
rect 10370 -1041 10378 -1007
rect 10412 -1041 10422 -1007
rect 10370 -1053 10422 -1041
rect 10632 -905 10684 -879
rect 10632 -939 10642 -905
rect 10676 -939 10684 -905
rect 10632 -1007 10684 -939
rect 10632 -1041 10642 -1007
rect 10676 -1041 10684 -1007
rect 10632 -1053 10684 -1041
rect 10738 -931 10809 -853
rect 10738 -965 10761 -931
rect 10795 -965 10809 -931
rect 10738 -999 10809 -965
rect 10738 -1033 10761 -999
rect 10795 -1033 10809 -999
rect 10738 -1053 10809 -1033
rect 10839 -889 10889 -853
rect 11286 -889 11336 -853
rect 10839 -932 10904 -889
rect 10839 -966 10859 -932
rect 10893 -966 10904 -932
rect 10839 -1000 10904 -966
rect 10839 -1034 10859 -1000
rect 10893 -1034 10904 -1000
rect 10839 -1053 10904 -1034
rect 11004 -931 11057 -889
rect 11004 -965 11015 -931
rect 11049 -965 11057 -931
rect 11004 -999 11057 -965
rect 11004 -1033 11015 -999
rect 11049 -1033 11057 -999
rect 11004 -1053 11057 -1033
rect 11111 -932 11164 -889
rect 11111 -966 11119 -932
rect 11153 -966 11164 -932
rect 11111 -1000 11164 -966
rect 11111 -1034 11119 -1000
rect 11153 -1034 11164 -1000
rect 11111 -1053 11164 -1034
rect 11264 -932 11336 -889
rect 11264 -966 11277 -932
rect 11311 -966 11336 -932
rect 11264 -1000 11336 -966
rect 11264 -1034 11277 -1000
rect 11311 -1034 11336 -1000
rect 11264 -1053 11336 -1034
rect 11366 -932 11420 -853
rect 11366 -966 11377 -932
rect 11411 -966 11420 -932
rect 11366 -1000 11420 -966
rect 11366 -1034 11377 -1000
rect 11411 -1034 11420 -1000
rect 11366 -1053 11420 -1034
rect 11658 -905 11710 -879
rect 11658 -939 11666 -905
rect 11700 -939 11710 -905
rect 11658 -1007 11710 -939
rect 11658 -1041 11666 -1007
rect 11700 -1041 11710 -1007
rect 11658 -1053 11710 -1041
rect 11920 -905 11972 -879
rect 11920 -939 11930 -905
rect 11964 -939 11972 -905
rect 11920 -1007 11972 -939
rect 11920 -1041 11930 -1007
rect 11964 -1041 11972 -1007
rect 13682 -939 13735 -853
rect 13682 -973 13690 -939
rect 13724 -973 13735 -939
rect 13682 -1007 13735 -973
rect 11920 -1053 11972 -1041
rect 13682 -1041 13690 -1007
rect 13724 -1041 13735 -1007
rect 13682 -1053 13735 -1041
rect 13765 -931 13821 -853
rect 13765 -965 13776 -931
rect 13810 -965 13821 -931
rect 13765 -999 13821 -965
rect 13765 -1033 13776 -999
rect 13810 -1033 13821 -999
rect 13765 -1053 13821 -1033
rect 13851 -939 13907 -853
rect 13851 -973 13862 -939
rect 13896 -973 13907 -939
rect 13851 -1007 13907 -973
rect 13851 -1041 13862 -1007
rect 13896 -1041 13907 -1007
rect 13851 -1053 13907 -1041
rect 13937 -923 13993 -853
rect 13937 -957 13948 -923
rect 13982 -957 13993 -923
rect 13937 -991 13993 -957
rect 13937 -1025 13948 -991
rect 13982 -1025 13993 -991
rect 13937 -1053 13993 -1025
rect 14023 -939 14079 -853
rect 14023 -973 14034 -939
rect 14068 -973 14079 -939
rect 14023 -1007 14079 -973
rect 14023 -1041 14034 -1007
rect 14068 -1041 14079 -1007
rect 14023 -1053 14079 -1041
rect 14109 -877 14165 -853
rect 14109 -911 14120 -877
rect 14154 -911 14165 -877
rect 14109 -963 14165 -911
rect 14109 -997 14120 -963
rect 14154 -997 14165 -963
rect 14109 -1053 14165 -997
rect 14195 -983 14251 -853
rect 14195 -1017 14206 -983
rect 14240 -1017 14251 -983
rect 14195 -1053 14251 -1017
rect 14281 -877 14337 -853
rect 14281 -911 14292 -877
rect 14326 -911 14337 -877
rect 14281 -963 14337 -911
rect 14281 -997 14292 -963
rect 14326 -997 14337 -963
rect 14281 -1053 14337 -997
rect 14367 -983 14423 -853
rect 14367 -1017 14378 -983
rect 14412 -1017 14423 -983
rect 14367 -1053 14423 -1017
rect 14453 -877 14509 -853
rect 14453 -911 14464 -877
rect 14498 -911 14509 -877
rect 14453 -963 14509 -911
rect 14453 -997 14464 -963
rect 14498 -997 14509 -963
rect 14453 -1053 14509 -997
rect 14539 -983 14595 -853
rect 14539 -1017 14550 -983
rect 14584 -1017 14595 -983
rect 14539 -1053 14595 -1017
rect 14625 -877 14681 -853
rect 14625 -911 14636 -877
rect 14670 -911 14681 -877
rect 14625 -963 14681 -911
rect 14625 -997 14636 -963
rect 14670 -997 14681 -963
rect 14625 -1053 14681 -997
rect 14711 -983 14766 -853
rect 14711 -1017 14722 -983
rect 14756 -1017 14766 -983
rect 14711 -1053 14766 -1017
rect 14796 -877 14852 -853
rect 14796 -911 14807 -877
rect 14841 -911 14852 -877
rect 14796 -963 14852 -911
rect 14796 -997 14807 -963
rect 14841 -997 14852 -963
rect 14796 -1053 14852 -997
rect 14882 -983 14938 -853
rect 14882 -1017 14893 -983
rect 14927 -1017 14938 -983
rect 14882 -1053 14938 -1017
rect 14968 -877 15024 -853
rect 14968 -911 14979 -877
rect 15013 -911 15024 -877
rect 14968 -963 15024 -911
rect 14968 -997 14979 -963
rect 15013 -997 15024 -963
rect 14968 -1053 15024 -997
rect 15054 -983 15110 -853
rect 15054 -1017 15065 -983
rect 15099 -1017 15110 -983
rect 15054 -1053 15110 -1017
rect 15140 -877 15196 -853
rect 15140 -911 15151 -877
rect 15185 -911 15196 -877
rect 15140 -963 15196 -911
rect 15140 -997 15151 -963
rect 15185 -997 15196 -963
rect 15140 -1053 15196 -997
rect 15226 -983 15282 -853
rect 15226 -1017 15237 -983
rect 15271 -1017 15282 -983
rect 15226 -1053 15282 -1017
rect 15312 -877 15368 -853
rect 15312 -911 15323 -877
rect 15357 -911 15368 -877
rect 15312 -963 15368 -911
rect 15312 -997 15323 -963
rect 15357 -997 15368 -963
rect 15312 -1053 15368 -997
rect 15398 -983 15451 -853
rect 15398 -1017 15409 -983
rect 15443 -1017 15451 -983
rect 15398 -1053 15451 -1017
rect 15614 -905 15666 -879
rect 15614 -939 15622 -905
rect 15656 -939 15666 -905
rect 15614 -1007 15666 -939
rect 15614 -1041 15622 -1007
rect 15656 -1041 15666 -1007
rect 15614 -1053 15666 -1041
rect 16612 -905 16664 -879
rect 16612 -939 16622 -905
rect 16656 -939 16664 -905
rect 16612 -1007 16664 -939
rect 16612 -1041 16622 -1007
rect 16656 -1041 16664 -1007
rect 16612 -1053 16664 -1041
rect -2970 -1159 -2918 -1147
rect -2970 -1193 -2962 -1159
rect -2928 -1193 -2918 -1159
rect -2970 -1261 -2918 -1193
rect -2970 -1295 -2962 -1261
rect -2928 -1295 -2918 -1261
rect -2970 -1321 -2918 -1295
rect -2340 -1159 -2288 -1147
rect -2340 -1193 -2330 -1159
rect -2296 -1193 -2288 -1159
rect -1590 -1159 -1538 -1147
rect -2340 -1261 -2288 -1193
rect -2340 -1295 -2330 -1261
rect -2296 -1295 -2288 -1261
rect -2340 -1321 -2288 -1295
rect -1590 -1193 -1582 -1159
rect -1548 -1193 -1538 -1159
rect -1590 -1261 -1538 -1193
rect -1590 -1295 -1582 -1261
rect -1548 -1295 -1538 -1261
rect -1590 -1321 -1538 -1295
rect -960 -1159 -908 -1147
rect -960 -1193 -950 -1159
rect -916 -1193 -908 -1159
rect -960 -1261 -908 -1193
rect -960 -1295 -950 -1261
rect -916 -1295 -908 -1261
rect -960 -1321 -908 -1295
rect -854 -1159 -802 -1147
rect -854 -1193 -846 -1159
rect -812 -1193 -802 -1159
rect -854 -1261 -802 -1193
rect -854 -1295 -846 -1261
rect -812 -1295 -802 -1261
rect -854 -1321 -802 -1295
rect -224 -1159 -172 -1147
rect -224 -1193 -214 -1159
rect -180 -1193 -172 -1159
rect -26 -1159 26 -1147
rect -224 -1261 -172 -1193
rect -224 -1295 -214 -1261
rect -180 -1295 -172 -1261
rect -224 -1321 -172 -1295
rect -26 -1193 -18 -1159
rect 16 -1193 26 -1159
rect -26 -1261 26 -1193
rect -26 -1295 -18 -1261
rect 16 -1295 26 -1261
rect -26 -1321 26 -1295
rect 236 -1159 288 -1147
rect 236 -1193 246 -1159
rect 280 -1193 288 -1159
rect 236 -1261 288 -1193
rect 236 -1295 246 -1261
rect 280 -1295 288 -1261
rect 236 -1321 288 -1295
rect 434 -1166 488 -1147
rect 434 -1200 443 -1166
rect 477 -1200 488 -1166
rect 434 -1234 488 -1200
rect 434 -1268 443 -1234
rect 477 -1268 488 -1234
rect 434 -1347 488 -1268
rect 518 -1166 590 -1147
rect 518 -1200 543 -1166
rect 577 -1200 590 -1166
rect 518 -1234 590 -1200
rect 518 -1268 543 -1234
rect 577 -1268 590 -1234
rect 518 -1311 590 -1268
rect 690 -1166 743 -1147
rect 690 -1200 701 -1166
rect 735 -1200 743 -1166
rect 690 -1234 743 -1200
rect 690 -1268 701 -1234
rect 735 -1268 743 -1234
rect 690 -1311 743 -1268
rect 797 -1167 850 -1147
rect 797 -1201 805 -1167
rect 839 -1201 850 -1167
rect 797 -1235 850 -1201
rect 797 -1269 805 -1235
rect 839 -1269 850 -1235
rect 797 -1311 850 -1269
rect 950 -1166 1015 -1147
rect 950 -1200 961 -1166
rect 995 -1200 1015 -1166
rect 950 -1234 1015 -1200
rect 950 -1268 961 -1234
rect 995 -1268 1015 -1234
rect 950 -1311 1015 -1268
rect 518 -1347 568 -1311
rect 965 -1347 1015 -1311
rect 1045 -1167 1116 -1147
rect 1262 -1159 1314 -1147
rect 1045 -1201 1059 -1167
rect 1093 -1201 1116 -1167
rect 1045 -1235 1116 -1201
rect 1045 -1269 1059 -1235
rect 1093 -1269 1116 -1235
rect 1045 -1347 1116 -1269
rect 1262 -1193 1270 -1159
rect 1304 -1193 1314 -1159
rect 1262 -1261 1314 -1193
rect 1262 -1295 1270 -1261
rect 1304 -1295 1314 -1261
rect 1262 -1321 1314 -1295
rect 1524 -1159 1576 -1147
rect 1524 -1193 1534 -1159
rect 1568 -1193 1576 -1159
rect 1722 -1159 1774 -1147
rect 1524 -1261 1576 -1193
rect 1524 -1295 1534 -1261
rect 1568 -1295 1576 -1261
rect 1524 -1321 1576 -1295
rect 1722 -1193 1730 -1159
rect 1764 -1193 1774 -1159
rect 1722 -1261 1774 -1193
rect 1722 -1295 1730 -1261
rect 1764 -1295 1774 -1261
rect 1722 -1321 1774 -1295
rect 2352 -1159 2404 -1147
rect 2352 -1193 2362 -1159
rect 2396 -1193 2404 -1159
rect 2550 -1159 2602 -1147
rect 2352 -1261 2404 -1193
rect 2352 -1295 2362 -1261
rect 2396 -1295 2404 -1261
rect 2352 -1321 2404 -1295
rect 2550 -1193 2558 -1159
rect 2592 -1193 2602 -1159
rect 2550 -1261 2602 -1193
rect 2550 -1295 2558 -1261
rect 2592 -1295 2602 -1261
rect 2550 -1321 2602 -1295
rect 2812 -1159 2864 -1147
rect 2812 -1193 2822 -1159
rect 2856 -1193 2864 -1159
rect 2812 -1261 2864 -1193
rect 2812 -1295 2822 -1261
rect 2856 -1295 2864 -1261
rect 2812 -1321 2864 -1295
rect 3010 -1166 3064 -1147
rect 3010 -1200 3019 -1166
rect 3053 -1200 3064 -1166
rect 3010 -1234 3064 -1200
rect 3010 -1268 3019 -1234
rect 3053 -1268 3064 -1234
rect 3010 -1347 3064 -1268
rect 3094 -1166 3166 -1147
rect 3094 -1200 3119 -1166
rect 3153 -1200 3166 -1166
rect 3094 -1234 3166 -1200
rect 3094 -1268 3119 -1234
rect 3153 -1268 3166 -1234
rect 3094 -1311 3166 -1268
rect 3266 -1166 3319 -1147
rect 3266 -1200 3277 -1166
rect 3311 -1200 3319 -1166
rect 3266 -1234 3319 -1200
rect 3266 -1268 3277 -1234
rect 3311 -1268 3319 -1234
rect 3266 -1311 3319 -1268
rect 3373 -1167 3426 -1147
rect 3373 -1201 3381 -1167
rect 3415 -1201 3426 -1167
rect 3373 -1235 3426 -1201
rect 3373 -1269 3381 -1235
rect 3415 -1269 3426 -1235
rect 3373 -1311 3426 -1269
rect 3526 -1166 3591 -1147
rect 3526 -1200 3537 -1166
rect 3571 -1200 3591 -1166
rect 3526 -1234 3591 -1200
rect 3526 -1268 3537 -1234
rect 3571 -1268 3591 -1234
rect 3526 -1311 3591 -1268
rect 3094 -1347 3144 -1311
rect 3541 -1347 3591 -1311
rect 3621 -1167 3692 -1147
rect 3838 -1159 3890 -1147
rect 3621 -1201 3635 -1167
rect 3669 -1201 3692 -1167
rect 3621 -1235 3692 -1201
rect 3621 -1269 3635 -1235
rect 3669 -1269 3692 -1235
rect 3621 -1347 3692 -1269
rect 3838 -1193 3846 -1159
rect 3880 -1193 3890 -1159
rect 3838 -1261 3890 -1193
rect 3838 -1295 3846 -1261
rect 3880 -1295 3890 -1261
rect 3838 -1321 3890 -1295
rect 4100 -1159 4152 -1147
rect 4100 -1193 4110 -1159
rect 4144 -1193 4152 -1159
rect 4298 -1159 4350 -1147
rect 4100 -1261 4152 -1193
rect 4100 -1295 4110 -1261
rect 4144 -1295 4152 -1261
rect 4100 -1321 4152 -1295
rect 4298 -1193 4306 -1159
rect 4340 -1193 4350 -1159
rect 4298 -1261 4350 -1193
rect 4298 -1295 4306 -1261
rect 4340 -1295 4350 -1261
rect 4298 -1321 4350 -1295
rect 4928 -1159 4980 -1147
rect 4928 -1193 4938 -1159
rect 4972 -1193 4980 -1159
rect 5126 -1159 5178 -1147
rect 4928 -1261 4980 -1193
rect 4928 -1295 4938 -1261
rect 4972 -1295 4980 -1261
rect 4928 -1321 4980 -1295
rect 5126 -1193 5134 -1159
rect 5168 -1193 5178 -1159
rect 5126 -1261 5178 -1193
rect 5126 -1295 5134 -1261
rect 5168 -1295 5178 -1261
rect 5126 -1321 5178 -1295
rect 5388 -1159 5440 -1147
rect 5388 -1193 5398 -1159
rect 5432 -1193 5440 -1159
rect 5388 -1261 5440 -1193
rect 5388 -1295 5398 -1261
rect 5432 -1295 5440 -1261
rect 5388 -1321 5440 -1295
rect 5586 -1166 5640 -1147
rect 5586 -1200 5595 -1166
rect 5629 -1200 5640 -1166
rect 5586 -1234 5640 -1200
rect 5586 -1268 5595 -1234
rect 5629 -1268 5640 -1234
rect 5586 -1347 5640 -1268
rect 5670 -1166 5742 -1147
rect 5670 -1200 5695 -1166
rect 5729 -1200 5742 -1166
rect 5670 -1234 5742 -1200
rect 5670 -1268 5695 -1234
rect 5729 -1268 5742 -1234
rect 5670 -1311 5742 -1268
rect 5842 -1166 5895 -1147
rect 5842 -1200 5853 -1166
rect 5887 -1200 5895 -1166
rect 5842 -1234 5895 -1200
rect 5842 -1268 5853 -1234
rect 5887 -1268 5895 -1234
rect 5842 -1311 5895 -1268
rect 5949 -1167 6002 -1147
rect 5949 -1201 5957 -1167
rect 5991 -1201 6002 -1167
rect 5949 -1235 6002 -1201
rect 5949 -1269 5957 -1235
rect 5991 -1269 6002 -1235
rect 5949 -1311 6002 -1269
rect 6102 -1166 6167 -1147
rect 6102 -1200 6113 -1166
rect 6147 -1200 6167 -1166
rect 6102 -1234 6167 -1200
rect 6102 -1268 6113 -1234
rect 6147 -1268 6167 -1234
rect 6102 -1311 6167 -1268
rect 5670 -1347 5720 -1311
rect 6117 -1347 6167 -1311
rect 6197 -1167 6268 -1147
rect 6414 -1159 6466 -1147
rect 6197 -1201 6211 -1167
rect 6245 -1201 6268 -1167
rect 6197 -1235 6268 -1201
rect 6197 -1269 6211 -1235
rect 6245 -1269 6268 -1235
rect 6197 -1347 6268 -1269
rect 6414 -1193 6422 -1159
rect 6456 -1193 6466 -1159
rect 6414 -1261 6466 -1193
rect 6414 -1295 6422 -1261
rect 6456 -1295 6466 -1261
rect 6414 -1321 6466 -1295
rect 6676 -1159 6728 -1147
rect 6676 -1193 6686 -1159
rect 6720 -1193 6728 -1159
rect 6874 -1159 6926 -1147
rect 6676 -1261 6728 -1193
rect 6676 -1295 6686 -1261
rect 6720 -1295 6728 -1261
rect 6676 -1321 6728 -1295
rect 6874 -1193 6882 -1159
rect 6916 -1193 6926 -1159
rect 6874 -1261 6926 -1193
rect 6874 -1295 6882 -1261
rect 6916 -1295 6926 -1261
rect 6874 -1321 6926 -1295
rect 7504 -1159 7556 -1147
rect 7504 -1193 7514 -1159
rect 7548 -1193 7556 -1159
rect 7702 -1159 7754 -1147
rect 7504 -1261 7556 -1193
rect 7504 -1295 7514 -1261
rect 7548 -1295 7556 -1261
rect 7504 -1321 7556 -1295
rect 7702 -1193 7710 -1159
rect 7744 -1193 7754 -1159
rect 7702 -1261 7754 -1193
rect 7702 -1295 7710 -1261
rect 7744 -1295 7754 -1261
rect 7702 -1321 7754 -1295
rect 7964 -1159 8016 -1147
rect 7964 -1193 7974 -1159
rect 8008 -1193 8016 -1159
rect 7964 -1261 8016 -1193
rect 7964 -1295 7974 -1261
rect 8008 -1295 8016 -1261
rect 7964 -1321 8016 -1295
rect 8162 -1166 8216 -1147
rect 8162 -1200 8171 -1166
rect 8205 -1200 8216 -1166
rect 8162 -1234 8216 -1200
rect 8162 -1268 8171 -1234
rect 8205 -1268 8216 -1234
rect 8162 -1347 8216 -1268
rect 8246 -1166 8318 -1147
rect 8246 -1200 8271 -1166
rect 8305 -1200 8318 -1166
rect 8246 -1234 8318 -1200
rect 8246 -1268 8271 -1234
rect 8305 -1268 8318 -1234
rect 8246 -1311 8318 -1268
rect 8418 -1166 8471 -1147
rect 8418 -1200 8429 -1166
rect 8463 -1200 8471 -1166
rect 8418 -1234 8471 -1200
rect 8418 -1268 8429 -1234
rect 8463 -1268 8471 -1234
rect 8418 -1311 8471 -1268
rect 8525 -1167 8578 -1147
rect 8525 -1201 8533 -1167
rect 8567 -1201 8578 -1167
rect 8525 -1235 8578 -1201
rect 8525 -1269 8533 -1235
rect 8567 -1269 8578 -1235
rect 8525 -1311 8578 -1269
rect 8678 -1166 8743 -1147
rect 8678 -1200 8689 -1166
rect 8723 -1200 8743 -1166
rect 8678 -1234 8743 -1200
rect 8678 -1268 8689 -1234
rect 8723 -1268 8743 -1234
rect 8678 -1311 8743 -1268
rect 8246 -1347 8296 -1311
rect 8693 -1347 8743 -1311
rect 8773 -1167 8844 -1147
rect 8990 -1159 9042 -1147
rect 8773 -1201 8787 -1167
rect 8821 -1201 8844 -1167
rect 8773 -1235 8844 -1201
rect 8773 -1269 8787 -1235
rect 8821 -1269 8844 -1235
rect 8773 -1347 8844 -1269
rect 8990 -1193 8998 -1159
rect 9032 -1193 9042 -1159
rect 8990 -1261 9042 -1193
rect 8990 -1295 8998 -1261
rect 9032 -1295 9042 -1261
rect 8990 -1321 9042 -1295
rect 9252 -1159 9304 -1147
rect 9252 -1193 9262 -1159
rect 9296 -1193 9304 -1159
rect 9450 -1159 9502 -1147
rect 9252 -1261 9304 -1193
rect 9252 -1295 9262 -1261
rect 9296 -1295 9304 -1261
rect 9252 -1321 9304 -1295
rect 9450 -1193 9458 -1159
rect 9492 -1193 9502 -1159
rect 9450 -1261 9502 -1193
rect 9450 -1295 9458 -1261
rect 9492 -1295 9502 -1261
rect 9450 -1321 9502 -1295
rect 10080 -1159 10132 -1147
rect 10080 -1193 10090 -1159
rect 10124 -1193 10132 -1159
rect 10370 -1159 10422 -1147
rect 10080 -1261 10132 -1193
rect 10080 -1295 10090 -1261
rect 10124 -1295 10132 -1261
rect 10080 -1321 10132 -1295
rect 10370 -1193 10378 -1159
rect 10412 -1193 10422 -1159
rect 10370 -1261 10422 -1193
rect 10370 -1295 10378 -1261
rect 10412 -1295 10422 -1261
rect 10370 -1321 10422 -1295
rect 10632 -1159 10684 -1147
rect 10632 -1193 10642 -1159
rect 10676 -1193 10684 -1159
rect 10632 -1261 10684 -1193
rect 10632 -1295 10642 -1261
rect 10676 -1295 10684 -1261
rect 10632 -1321 10684 -1295
rect 10738 -1166 10792 -1147
rect 10738 -1200 10747 -1166
rect 10781 -1200 10792 -1166
rect 10738 -1234 10792 -1200
rect 10738 -1268 10747 -1234
rect 10781 -1268 10792 -1234
rect 10738 -1347 10792 -1268
rect 10822 -1166 10894 -1147
rect 10822 -1200 10847 -1166
rect 10881 -1200 10894 -1166
rect 10822 -1234 10894 -1200
rect 10822 -1268 10847 -1234
rect 10881 -1268 10894 -1234
rect 10822 -1311 10894 -1268
rect 10994 -1166 11047 -1147
rect 10994 -1200 11005 -1166
rect 11039 -1200 11047 -1166
rect 10994 -1234 11047 -1200
rect 10994 -1268 11005 -1234
rect 11039 -1268 11047 -1234
rect 10994 -1311 11047 -1268
rect 11101 -1167 11154 -1147
rect 11101 -1201 11109 -1167
rect 11143 -1201 11154 -1167
rect 11101 -1235 11154 -1201
rect 11101 -1269 11109 -1235
rect 11143 -1269 11154 -1235
rect 11101 -1311 11154 -1269
rect 11254 -1166 11319 -1147
rect 11254 -1200 11265 -1166
rect 11299 -1200 11319 -1166
rect 11254 -1234 11319 -1200
rect 11254 -1268 11265 -1234
rect 11299 -1268 11319 -1234
rect 11254 -1311 11319 -1268
rect 10822 -1347 10872 -1311
rect 11269 -1347 11319 -1311
rect 11349 -1167 11420 -1147
rect 11658 -1159 11710 -1147
rect 11349 -1201 11363 -1167
rect 11397 -1201 11420 -1167
rect 11349 -1235 11420 -1201
rect 11349 -1269 11363 -1235
rect 11397 -1269 11420 -1235
rect 11349 -1347 11420 -1269
rect 11658 -1193 11666 -1159
rect 11700 -1193 11710 -1159
rect 11658 -1261 11710 -1193
rect 11658 -1295 11666 -1261
rect 11700 -1295 11710 -1261
rect 11658 -1321 11710 -1295
rect 11920 -1159 11972 -1147
rect 11920 -1193 11930 -1159
rect 11964 -1193 11972 -1159
rect 11920 -1261 11972 -1193
rect 11920 -1295 11930 -1261
rect 11964 -1295 11972 -1261
rect 11920 -1321 11972 -1295
rect 12486 -1166 12547 -1147
rect 12486 -1200 12502 -1166
rect 12536 -1200 12547 -1166
rect 12486 -1234 12547 -1200
rect 12486 -1268 12502 -1234
rect 12536 -1268 12547 -1234
rect 12486 -1347 12547 -1268
rect 12577 -1173 12633 -1147
rect 12577 -1207 12588 -1173
rect 12622 -1207 12633 -1173
rect 12577 -1261 12633 -1207
rect 12577 -1295 12588 -1261
rect 12622 -1295 12633 -1261
rect 12577 -1347 12633 -1295
rect 12663 -1166 12719 -1147
rect 12663 -1200 12674 -1166
rect 12708 -1200 12719 -1166
rect 12663 -1234 12719 -1200
rect 12663 -1268 12674 -1234
rect 12708 -1268 12719 -1234
rect 12663 -1347 12719 -1268
rect 12749 -1173 12805 -1147
rect 12749 -1207 12760 -1173
rect 12794 -1207 12805 -1173
rect 12749 -1261 12805 -1207
rect 12749 -1295 12760 -1261
rect 12794 -1295 12805 -1261
rect 12749 -1347 12805 -1295
rect 12835 -1166 12891 -1147
rect 12835 -1200 12846 -1166
rect 12880 -1200 12891 -1166
rect 12835 -1234 12891 -1200
rect 12835 -1268 12846 -1234
rect 12880 -1268 12891 -1234
rect 12835 -1347 12891 -1268
rect 12921 -1173 12977 -1147
rect 12921 -1207 12932 -1173
rect 12966 -1207 12977 -1173
rect 12921 -1261 12977 -1207
rect 12921 -1295 12932 -1261
rect 12966 -1295 12977 -1261
rect 12921 -1347 12977 -1295
rect 13007 -1166 13076 -1147
rect 13222 -1159 13274 -1147
rect 13007 -1200 13018 -1166
rect 13052 -1200 13076 -1166
rect 13007 -1234 13076 -1200
rect 13007 -1268 13018 -1234
rect 13052 -1268 13076 -1234
rect 13007 -1347 13076 -1268
rect 13222 -1193 13230 -1159
rect 13264 -1193 13274 -1159
rect 13222 -1261 13274 -1193
rect 13222 -1295 13230 -1261
rect 13264 -1295 13274 -1261
rect 13222 -1321 13274 -1295
rect 13484 -1159 13536 -1147
rect 13484 -1193 13494 -1159
rect 13528 -1193 13536 -1159
rect 13682 -1159 13735 -1147
rect 13484 -1261 13536 -1193
rect 13484 -1295 13494 -1261
rect 13528 -1295 13536 -1261
rect 13484 -1321 13536 -1295
rect 13682 -1193 13690 -1159
rect 13724 -1193 13735 -1159
rect 13682 -1227 13735 -1193
rect 13682 -1261 13690 -1227
rect 13724 -1261 13735 -1227
rect 13682 -1347 13735 -1261
rect 13765 -1167 13821 -1147
rect 13765 -1201 13776 -1167
rect 13810 -1201 13821 -1167
rect 13765 -1235 13821 -1201
rect 13765 -1269 13776 -1235
rect 13810 -1269 13821 -1235
rect 13765 -1347 13821 -1269
rect 13851 -1159 13907 -1147
rect 13851 -1193 13862 -1159
rect 13896 -1193 13907 -1159
rect 13851 -1227 13907 -1193
rect 13851 -1261 13862 -1227
rect 13896 -1261 13907 -1227
rect 13851 -1347 13907 -1261
rect 13937 -1175 13993 -1147
rect 13937 -1209 13948 -1175
rect 13982 -1209 13993 -1175
rect 13937 -1243 13993 -1209
rect 13937 -1277 13948 -1243
rect 13982 -1277 13993 -1243
rect 13937 -1347 13993 -1277
rect 14023 -1159 14079 -1147
rect 14023 -1193 14034 -1159
rect 14068 -1193 14079 -1159
rect 14023 -1227 14079 -1193
rect 14023 -1261 14034 -1227
rect 14068 -1261 14079 -1227
rect 14023 -1347 14079 -1261
rect 14109 -1203 14165 -1147
rect 14109 -1237 14120 -1203
rect 14154 -1237 14165 -1203
rect 14109 -1289 14165 -1237
rect 14109 -1323 14120 -1289
rect 14154 -1323 14165 -1289
rect 14109 -1347 14165 -1323
rect 14195 -1183 14251 -1147
rect 14195 -1217 14206 -1183
rect 14240 -1217 14251 -1183
rect 14195 -1347 14251 -1217
rect 14281 -1203 14337 -1147
rect 14281 -1237 14292 -1203
rect 14326 -1237 14337 -1203
rect 14281 -1289 14337 -1237
rect 14281 -1323 14292 -1289
rect 14326 -1323 14337 -1289
rect 14281 -1347 14337 -1323
rect 14367 -1183 14423 -1147
rect 14367 -1217 14378 -1183
rect 14412 -1217 14423 -1183
rect 14367 -1347 14423 -1217
rect 14453 -1203 14509 -1147
rect 14453 -1237 14464 -1203
rect 14498 -1237 14509 -1203
rect 14453 -1289 14509 -1237
rect 14453 -1323 14464 -1289
rect 14498 -1323 14509 -1289
rect 14453 -1347 14509 -1323
rect 14539 -1183 14595 -1147
rect 14539 -1217 14550 -1183
rect 14584 -1217 14595 -1183
rect 14539 -1347 14595 -1217
rect 14625 -1203 14681 -1147
rect 14625 -1237 14636 -1203
rect 14670 -1237 14681 -1203
rect 14625 -1289 14681 -1237
rect 14625 -1323 14636 -1289
rect 14670 -1323 14681 -1289
rect 14625 -1347 14681 -1323
rect 14711 -1183 14766 -1147
rect 14711 -1217 14722 -1183
rect 14756 -1217 14766 -1183
rect 14711 -1347 14766 -1217
rect 14796 -1203 14852 -1147
rect 14796 -1237 14807 -1203
rect 14841 -1237 14852 -1203
rect 14796 -1289 14852 -1237
rect 14796 -1323 14807 -1289
rect 14841 -1323 14852 -1289
rect 14796 -1347 14852 -1323
rect 14882 -1183 14938 -1147
rect 14882 -1217 14893 -1183
rect 14927 -1217 14938 -1183
rect 14882 -1347 14938 -1217
rect 14968 -1203 15024 -1147
rect 14968 -1237 14979 -1203
rect 15013 -1237 15024 -1203
rect 14968 -1289 15024 -1237
rect 14968 -1323 14979 -1289
rect 15013 -1323 15024 -1289
rect 14968 -1347 15024 -1323
rect 15054 -1183 15110 -1147
rect 15054 -1217 15065 -1183
rect 15099 -1217 15110 -1183
rect 15054 -1347 15110 -1217
rect 15140 -1203 15196 -1147
rect 15140 -1237 15151 -1203
rect 15185 -1237 15196 -1203
rect 15140 -1289 15196 -1237
rect 15140 -1323 15151 -1289
rect 15185 -1323 15196 -1289
rect 15140 -1347 15196 -1323
rect 15226 -1183 15282 -1147
rect 15226 -1217 15237 -1183
rect 15271 -1217 15282 -1183
rect 15226 -1347 15282 -1217
rect 15312 -1203 15368 -1147
rect 15312 -1237 15323 -1203
rect 15357 -1237 15368 -1203
rect 15312 -1289 15368 -1237
rect 15312 -1323 15323 -1289
rect 15357 -1323 15368 -1289
rect 15312 -1347 15368 -1323
rect 15398 -1183 15451 -1147
rect 15614 -1159 15666 -1147
rect 15398 -1217 15409 -1183
rect 15443 -1217 15451 -1183
rect 15398 -1347 15451 -1217
rect 15614 -1193 15622 -1159
rect 15656 -1193 15666 -1159
rect 15614 -1261 15666 -1193
rect 15614 -1295 15622 -1261
rect 15656 -1295 15666 -1261
rect 15614 -1321 15666 -1295
rect 16612 -1159 16664 -1147
rect 16612 -1193 16622 -1159
rect 16656 -1193 16664 -1159
rect 16612 -1261 16664 -1193
rect 16612 -1295 16622 -1261
rect 16656 -1295 16664 -1261
rect 16612 -1321 16664 -1295
rect -2970 -1993 -2918 -1967
rect -2970 -2027 -2962 -1993
rect -2928 -2027 -2918 -1993
rect -2970 -2095 -2918 -2027
rect -2970 -2129 -2962 -2095
rect -2928 -2129 -2918 -2095
rect -2970 -2141 -2918 -2129
rect -2340 -1993 -2288 -1967
rect -2340 -2027 -2330 -1993
rect -2296 -2027 -2288 -1993
rect -2340 -2095 -2288 -2027
rect -2340 -2129 -2330 -2095
rect -2296 -2129 -2288 -2095
rect -1590 -1993 -1538 -1967
rect -1590 -2027 -1582 -1993
rect -1548 -2027 -1538 -1993
rect -1590 -2095 -1538 -2027
rect -2340 -2141 -2288 -2129
rect -1590 -2129 -1582 -2095
rect -1548 -2129 -1538 -2095
rect -1590 -2141 -1538 -2129
rect -960 -1993 -908 -1967
rect -960 -2027 -950 -1993
rect -916 -2027 -908 -1993
rect -960 -2095 -908 -2027
rect -960 -2129 -950 -2095
rect -916 -2129 -908 -2095
rect -960 -2141 -908 -2129
rect -854 -2019 -783 -1941
rect -854 -2053 -831 -2019
rect -797 -2053 -783 -2019
rect -854 -2087 -783 -2053
rect -854 -2121 -831 -2087
rect -797 -2121 -783 -2087
rect -854 -2141 -783 -2121
rect -753 -1977 -703 -1941
rect -306 -1977 -256 -1941
rect -753 -2020 -688 -1977
rect -753 -2054 -733 -2020
rect -699 -2054 -688 -2020
rect -753 -2088 -688 -2054
rect -753 -2122 -733 -2088
rect -699 -2122 -688 -2088
rect -753 -2141 -688 -2122
rect -588 -2019 -535 -1977
rect -588 -2053 -577 -2019
rect -543 -2053 -535 -2019
rect -588 -2087 -535 -2053
rect -588 -2121 -577 -2087
rect -543 -2121 -535 -2087
rect -588 -2141 -535 -2121
rect -481 -2020 -428 -1977
rect -481 -2054 -473 -2020
rect -439 -2054 -428 -2020
rect -481 -2088 -428 -2054
rect -481 -2122 -473 -2088
rect -439 -2122 -428 -2088
rect -481 -2141 -428 -2122
rect -328 -2020 -256 -1977
rect -328 -2054 -315 -2020
rect -281 -2054 -256 -2020
rect -328 -2088 -256 -2054
rect -328 -2122 -315 -2088
rect -281 -2122 -256 -2088
rect -328 -2141 -256 -2122
rect -226 -2020 -172 -1941
rect -226 -2054 -215 -2020
rect -181 -2054 -172 -2020
rect -226 -2088 -172 -2054
rect -226 -2122 -215 -2088
rect -181 -2122 -172 -2088
rect -226 -2141 -172 -2122
rect -26 -1993 26 -1967
rect -26 -2027 -18 -1993
rect 16 -2027 26 -1993
rect -26 -2095 26 -2027
rect -26 -2129 -18 -2095
rect 16 -2129 26 -2095
rect -26 -2141 26 -2129
rect 236 -1993 288 -1967
rect 236 -2027 246 -1993
rect 280 -2027 288 -1993
rect 236 -2095 288 -2027
rect 236 -2129 246 -2095
rect 280 -2129 288 -2095
rect 434 -2019 505 -1941
rect 434 -2053 457 -2019
rect 491 -2053 505 -2019
rect 434 -2087 505 -2053
rect 434 -2121 457 -2087
rect 491 -2121 505 -2087
rect 236 -2141 288 -2129
rect 434 -2141 505 -2121
rect 535 -1977 585 -1941
rect 982 -1977 1032 -1941
rect 535 -2020 600 -1977
rect 535 -2054 555 -2020
rect 589 -2054 600 -2020
rect 535 -2088 600 -2054
rect 535 -2122 555 -2088
rect 589 -2122 600 -2088
rect 535 -2141 600 -2122
rect 700 -2019 753 -1977
rect 700 -2053 711 -2019
rect 745 -2053 753 -2019
rect 700 -2087 753 -2053
rect 700 -2121 711 -2087
rect 745 -2121 753 -2087
rect 700 -2141 753 -2121
rect 807 -2020 860 -1977
rect 807 -2054 815 -2020
rect 849 -2054 860 -2020
rect 807 -2088 860 -2054
rect 807 -2122 815 -2088
rect 849 -2122 860 -2088
rect 807 -2141 860 -2122
rect 960 -2020 1032 -1977
rect 960 -2054 973 -2020
rect 1007 -2054 1032 -2020
rect 960 -2088 1032 -2054
rect 960 -2122 973 -2088
rect 1007 -2122 1032 -2088
rect 960 -2141 1032 -2122
rect 1062 -2020 1116 -1941
rect 1062 -2054 1073 -2020
rect 1107 -2054 1116 -2020
rect 1062 -2088 1116 -2054
rect 1062 -2122 1073 -2088
rect 1107 -2122 1116 -2088
rect 1062 -2141 1116 -2122
rect 1262 -1993 1314 -1967
rect 1262 -2027 1270 -1993
rect 1304 -2027 1314 -1993
rect 1262 -2095 1314 -2027
rect 1262 -2129 1270 -2095
rect 1304 -2129 1314 -2095
rect 1262 -2141 1314 -2129
rect 1524 -1993 1576 -1967
rect 1524 -2027 1534 -1993
rect 1568 -2027 1576 -1993
rect 1524 -2095 1576 -2027
rect 1524 -2129 1534 -2095
rect 1568 -2129 1576 -2095
rect 1722 -1993 1774 -1967
rect 1722 -2027 1730 -1993
rect 1764 -2027 1774 -1993
rect 1722 -2095 1774 -2027
rect 1524 -2141 1576 -2129
rect 1722 -2129 1730 -2095
rect 1764 -2129 1774 -2095
rect 1722 -2141 1774 -2129
rect 2352 -1993 2404 -1967
rect 2352 -2027 2362 -1993
rect 2396 -2027 2404 -1993
rect 2352 -2095 2404 -2027
rect 2352 -2129 2362 -2095
rect 2396 -2129 2404 -2095
rect 2550 -1993 2602 -1967
rect 2550 -2027 2558 -1993
rect 2592 -2027 2602 -1993
rect 2550 -2095 2602 -2027
rect 2352 -2141 2404 -2129
rect 2550 -2129 2558 -2095
rect 2592 -2129 2602 -2095
rect 2550 -2141 2602 -2129
rect 2812 -1993 2864 -1967
rect 2812 -2027 2822 -1993
rect 2856 -2027 2864 -1993
rect 2812 -2095 2864 -2027
rect 2812 -2129 2822 -2095
rect 2856 -2129 2864 -2095
rect 3010 -2019 3081 -1941
rect 3010 -2053 3033 -2019
rect 3067 -2053 3081 -2019
rect 3010 -2087 3081 -2053
rect 3010 -2121 3033 -2087
rect 3067 -2121 3081 -2087
rect 2812 -2141 2864 -2129
rect 3010 -2141 3081 -2121
rect 3111 -1977 3161 -1941
rect 3558 -1977 3608 -1941
rect 3111 -2020 3176 -1977
rect 3111 -2054 3131 -2020
rect 3165 -2054 3176 -2020
rect 3111 -2088 3176 -2054
rect 3111 -2122 3131 -2088
rect 3165 -2122 3176 -2088
rect 3111 -2141 3176 -2122
rect 3276 -2019 3329 -1977
rect 3276 -2053 3287 -2019
rect 3321 -2053 3329 -2019
rect 3276 -2087 3329 -2053
rect 3276 -2121 3287 -2087
rect 3321 -2121 3329 -2087
rect 3276 -2141 3329 -2121
rect 3383 -2020 3436 -1977
rect 3383 -2054 3391 -2020
rect 3425 -2054 3436 -2020
rect 3383 -2088 3436 -2054
rect 3383 -2122 3391 -2088
rect 3425 -2122 3436 -2088
rect 3383 -2141 3436 -2122
rect 3536 -2020 3608 -1977
rect 3536 -2054 3549 -2020
rect 3583 -2054 3608 -2020
rect 3536 -2088 3608 -2054
rect 3536 -2122 3549 -2088
rect 3583 -2122 3608 -2088
rect 3536 -2141 3608 -2122
rect 3638 -2020 3692 -1941
rect 3638 -2054 3649 -2020
rect 3683 -2054 3692 -2020
rect 3638 -2088 3692 -2054
rect 3638 -2122 3649 -2088
rect 3683 -2122 3692 -2088
rect 3638 -2141 3692 -2122
rect 3838 -1993 3890 -1967
rect 3838 -2027 3846 -1993
rect 3880 -2027 3890 -1993
rect 3838 -2095 3890 -2027
rect 3838 -2129 3846 -2095
rect 3880 -2129 3890 -2095
rect 3838 -2141 3890 -2129
rect 4100 -1993 4152 -1967
rect 4100 -2027 4110 -1993
rect 4144 -2027 4152 -1993
rect 4100 -2095 4152 -2027
rect 4100 -2129 4110 -2095
rect 4144 -2129 4152 -2095
rect 4298 -1993 4350 -1967
rect 4298 -2027 4306 -1993
rect 4340 -2027 4350 -1993
rect 4298 -2095 4350 -2027
rect 4100 -2141 4152 -2129
rect 4298 -2129 4306 -2095
rect 4340 -2129 4350 -2095
rect 4298 -2141 4350 -2129
rect 4928 -1993 4980 -1967
rect 4928 -2027 4938 -1993
rect 4972 -2027 4980 -1993
rect 4928 -2095 4980 -2027
rect 4928 -2129 4938 -2095
rect 4972 -2129 4980 -2095
rect 5126 -1993 5178 -1967
rect 5126 -2027 5134 -1993
rect 5168 -2027 5178 -1993
rect 5126 -2095 5178 -2027
rect 4928 -2141 4980 -2129
rect 5126 -2129 5134 -2095
rect 5168 -2129 5178 -2095
rect 5126 -2141 5178 -2129
rect 5388 -1993 5440 -1967
rect 5388 -2027 5398 -1993
rect 5432 -2027 5440 -1993
rect 5388 -2095 5440 -2027
rect 5388 -2129 5398 -2095
rect 5432 -2129 5440 -2095
rect 5586 -2019 5657 -1941
rect 5586 -2053 5609 -2019
rect 5643 -2053 5657 -2019
rect 5586 -2087 5657 -2053
rect 5586 -2121 5609 -2087
rect 5643 -2121 5657 -2087
rect 5388 -2141 5440 -2129
rect 5586 -2141 5657 -2121
rect 5687 -1977 5737 -1941
rect 6134 -1977 6184 -1941
rect 5687 -2020 5752 -1977
rect 5687 -2054 5707 -2020
rect 5741 -2054 5752 -2020
rect 5687 -2088 5752 -2054
rect 5687 -2122 5707 -2088
rect 5741 -2122 5752 -2088
rect 5687 -2141 5752 -2122
rect 5852 -2019 5905 -1977
rect 5852 -2053 5863 -2019
rect 5897 -2053 5905 -2019
rect 5852 -2087 5905 -2053
rect 5852 -2121 5863 -2087
rect 5897 -2121 5905 -2087
rect 5852 -2141 5905 -2121
rect 5959 -2020 6012 -1977
rect 5959 -2054 5967 -2020
rect 6001 -2054 6012 -2020
rect 5959 -2088 6012 -2054
rect 5959 -2122 5967 -2088
rect 6001 -2122 6012 -2088
rect 5959 -2141 6012 -2122
rect 6112 -2020 6184 -1977
rect 6112 -2054 6125 -2020
rect 6159 -2054 6184 -2020
rect 6112 -2088 6184 -2054
rect 6112 -2122 6125 -2088
rect 6159 -2122 6184 -2088
rect 6112 -2141 6184 -2122
rect 6214 -2020 6268 -1941
rect 6214 -2054 6225 -2020
rect 6259 -2054 6268 -2020
rect 6214 -2088 6268 -2054
rect 6214 -2122 6225 -2088
rect 6259 -2122 6268 -2088
rect 6214 -2141 6268 -2122
rect 6414 -1993 6466 -1967
rect 6414 -2027 6422 -1993
rect 6456 -2027 6466 -1993
rect 6414 -2095 6466 -2027
rect 6414 -2129 6422 -2095
rect 6456 -2129 6466 -2095
rect 6414 -2141 6466 -2129
rect 6676 -1993 6728 -1967
rect 6676 -2027 6686 -1993
rect 6720 -2027 6728 -1993
rect 6676 -2095 6728 -2027
rect 6676 -2129 6686 -2095
rect 6720 -2129 6728 -2095
rect 6874 -1993 6926 -1967
rect 6874 -2027 6882 -1993
rect 6916 -2027 6926 -1993
rect 6874 -2095 6926 -2027
rect 6676 -2141 6728 -2129
rect 6874 -2129 6882 -2095
rect 6916 -2129 6926 -2095
rect 6874 -2141 6926 -2129
rect 7504 -1993 7556 -1967
rect 7504 -2027 7514 -1993
rect 7548 -2027 7556 -1993
rect 7504 -2095 7556 -2027
rect 7504 -2129 7514 -2095
rect 7548 -2129 7556 -2095
rect 7702 -1993 7754 -1967
rect 7702 -2027 7710 -1993
rect 7744 -2027 7754 -1993
rect 7702 -2095 7754 -2027
rect 7504 -2141 7556 -2129
rect 7702 -2129 7710 -2095
rect 7744 -2129 7754 -2095
rect 7702 -2141 7754 -2129
rect 7964 -1993 8016 -1967
rect 7964 -2027 7974 -1993
rect 8008 -2027 8016 -1993
rect 7964 -2095 8016 -2027
rect 7964 -2129 7974 -2095
rect 8008 -2129 8016 -2095
rect 8162 -2019 8233 -1941
rect 8162 -2053 8185 -2019
rect 8219 -2053 8233 -2019
rect 8162 -2087 8233 -2053
rect 8162 -2121 8185 -2087
rect 8219 -2121 8233 -2087
rect 7964 -2141 8016 -2129
rect 8162 -2141 8233 -2121
rect 8263 -1977 8313 -1941
rect 8710 -1977 8760 -1941
rect 8263 -2020 8328 -1977
rect 8263 -2054 8283 -2020
rect 8317 -2054 8328 -2020
rect 8263 -2088 8328 -2054
rect 8263 -2122 8283 -2088
rect 8317 -2122 8328 -2088
rect 8263 -2141 8328 -2122
rect 8428 -2019 8481 -1977
rect 8428 -2053 8439 -2019
rect 8473 -2053 8481 -2019
rect 8428 -2087 8481 -2053
rect 8428 -2121 8439 -2087
rect 8473 -2121 8481 -2087
rect 8428 -2141 8481 -2121
rect 8535 -2020 8588 -1977
rect 8535 -2054 8543 -2020
rect 8577 -2054 8588 -2020
rect 8535 -2088 8588 -2054
rect 8535 -2122 8543 -2088
rect 8577 -2122 8588 -2088
rect 8535 -2141 8588 -2122
rect 8688 -2020 8760 -1977
rect 8688 -2054 8701 -2020
rect 8735 -2054 8760 -2020
rect 8688 -2088 8760 -2054
rect 8688 -2122 8701 -2088
rect 8735 -2122 8760 -2088
rect 8688 -2141 8760 -2122
rect 8790 -2020 8844 -1941
rect 8790 -2054 8801 -2020
rect 8835 -2054 8844 -2020
rect 8790 -2088 8844 -2054
rect 8790 -2122 8801 -2088
rect 8835 -2122 8844 -2088
rect 8790 -2141 8844 -2122
rect 8990 -1993 9042 -1967
rect 8990 -2027 8998 -1993
rect 9032 -2027 9042 -1993
rect 8990 -2095 9042 -2027
rect 8990 -2129 8998 -2095
rect 9032 -2129 9042 -2095
rect 8990 -2141 9042 -2129
rect 9252 -1993 9304 -1967
rect 9252 -2027 9262 -1993
rect 9296 -2027 9304 -1993
rect 9252 -2095 9304 -2027
rect 9252 -2129 9262 -2095
rect 9296 -2129 9304 -2095
rect 9450 -1993 9502 -1967
rect 9450 -2027 9458 -1993
rect 9492 -2027 9502 -1993
rect 9450 -2095 9502 -2027
rect 9252 -2141 9304 -2129
rect 9450 -2129 9458 -2095
rect 9492 -2129 9502 -2095
rect 9450 -2141 9502 -2129
rect 10080 -1993 10132 -1967
rect 10080 -2027 10090 -1993
rect 10124 -2027 10132 -1993
rect 10080 -2095 10132 -2027
rect 10080 -2129 10090 -2095
rect 10124 -2129 10132 -2095
rect 10370 -1993 10422 -1967
rect 10370 -2027 10378 -1993
rect 10412 -2027 10422 -1993
rect 10370 -2095 10422 -2027
rect 10080 -2141 10132 -2129
rect 10370 -2129 10378 -2095
rect 10412 -2129 10422 -2095
rect 10370 -2141 10422 -2129
rect 10632 -1993 10684 -1967
rect 10632 -2027 10642 -1993
rect 10676 -2027 10684 -1993
rect 10632 -2095 10684 -2027
rect 10632 -2129 10642 -2095
rect 10676 -2129 10684 -2095
rect 10632 -2141 10684 -2129
rect 10738 -2019 10809 -1941
rect 10738 -2053 10761 -2019
rect 10795 -2053 10809 -2019
rect 10738 -2087 10809 -2053
rect 10738 -2121 10761 -2087
rect 10795 -2121 10809 -2087
rect 10738 -2141 10809 -2121
rect 10839 -1977 10889 -1941
rect 11286 -1977 11336 -1941
rect 10839 -2020 10904 -1977
rect 10839 -2054 10859 -2020
rect 10893 -2054 10904 -2020
rect 10839 -2088 10904 -2054
rect 10839 -2122 10859 -2088
rect 10893 -2122 10904 -2088
rect 10839 -2141 10904 -2122
rect 11004 -2019 11057 -1977
rect 11004 -2053 11015 -2019
rect 11049 -2053 11057 -2019
rect 11004 -2087 11057 -2053
rect 11004 -2121 11015 -2087
rect 11049 -2121 11057 -2087
rect 11004 -2141 11057 -2121
rect 11111 -2020 11164 -1977
rect 11111 -2054 11119 -2020
rect 11153 -2054 11164 -2020
rect 11111 -2088 11164 -2054
rect 11111 -2122 11119 -2088
rect 11153 -2122 11164 -2088
rect 11111 -2141 11164 -2122
rect 11264 -2020 11336 -1977
rect 11264 -2054 11277 -2020
rect 11311 -2054 11336 -2020
rect 11264 -2088 11336 -2054
rect 11264 -2122 11277 -2088
rect 11311 -2122 11336 -2088
rect 11264 -2141 11336 -2122
rect 11366 -2020 11420 -1941
rect 11366 -2054 11377 -2020
rect 11411 -2054 11420 -2020
rect 11366 -2088 11420 -2054
rect 11366 -2122 11377 -2088
rect 11411 -2122 11420 -2088
rect 11366 -2141 11420 -2122
rect 11658 -1993 11710 -1967
rect 11658 -2027 11666 -1993
rect 11700 -2027 11710 -1993
rect 11658 -2095 11710 -2027
rect 11658 -2129 11666 -2095
rect 11700 -2129 11710 -2095
rect 11658 -2141 11710 -2129
rect 11920 -1993 11972 -1967
rect 11920 -2027 11930 -1993
rect 11964 -2027 11972 -1993
rect 11920 -2095 11972 -2027
rect 11920 -2129 11930 -2095
rect 11964 -2129 11972 -2095
rect 13682 -2027 13735 -1941
rect 13682 -2061 13690 -2027
rect 13724 -2061 13735 -2027
rect 13682 -2095 13735 -2061
rect 11920 -2141 11972 -2129
rect 13682 -2129 13690 -2095
rect 13724 -2129 13735 -2095
rect 13682 -2141 13735 -2129
rect 13765 -2019 13821 -1941
rect 13765 -2053 13776 -2019
rect 13810 -2053 13821 -2019
rect 13765 -2087 13821 -2053
rect 13765 -2121 13776 -2087
rect 13810 -2121 13821 -2087
rect 13765 -2141 13821 -2121
rect 13851 -2027 13907 -1941
rect 13851 -2061 13862 -2027
rect 13896 -2061 13907 -2027
rect 13851 -2095 13907 -2061
rect 13851 -2129 13862 -2095
rect 13896 -2129 13907 -2095
rect 13851 -2141 13907 -2129
rect 13937 -2011 13993 -1941
rect 13937 -2045 13948 -2011
rect 13982 -2045 13993 -2011
rect 13937 -2079 13993 -2045
rect 13937 -2113 13948 -2079
rect 13982 -2113 13993 -2079
rect 13937 -2141 13993 -2113
rect 14023 -2027 14079 -1941
rect 14023 -2061 14034 -2027
rect 14068 -2061 14079 -2027
rect 14023 -2095 14079 -2061
rect 14023 -2129 14034 -2095
rect 14068 -2129 14079 -2095
rect 14023 -2141 14079 -2129
rect 14109 -1965 14165 -1941
rect 14109 -1999 14120 -1965
rect 14154 -1999 14165 -1965
rect 14109 -2051 14165 -1999
rect 14109 -2085 14120 -2051
rect 14154 -2085 14165 -2051
rect 14109 -2141 14165 -2085
rect 14195 -2071 14251 -1941
rect 14195 -2105 14206 -2071
rect 14240 -2105 14251 -2071
rect 14195 -2141 14251 -2105
rect 14281 -1965 14337 -1941
rect 14281 -1999 14292 -1965
rect 14326 -1999 14337 -1965
rect 14281 -2051 14337 -1999
rect 14281 -2085 14292 -2051
rect 14326 -2085 14337 -2051
rect 14281 -2141 14337 -2085
rect 14367 -2071 14423 -1941
rect 14367 -2105 14378 -2071
rect 14412 -2105 14423 -2071
rect 14367 -2141 14423 -2105
rect 14453 -1965 14509 -1941
rect 14453 -1999 14464 -1965
rect 14498 -1999 14509 -1965
rect 14453 -2051 14509 -1999
rect 14453 -2085 14464 -2051
rect 14498 -2085 14509 -2051
rect 14453 -2141 14509 -2085
rect 14539 -2071 14595 -1941
rect 14539 -2105 14550 -2071
rect 14584 -2105 14595 -2071
rect 14539 -2141 14595 -2105
rect 14625 -1965 14681 -1941
rect 14625 -1999 14636 -1965
rect 14670 -1999 14681 -1965
rect 14625 -2051 14681 -1999
rect 14625 -2085 14636 -2051
rect 14670 -2085 14681 -2051
rect 14625 -2141 14681 -2085
rect 14711 -2071 14766 -1941
rect 14711 -2105 14722 -2071
rect 14756 -2105 14766 -2071
rect 14711 -2141 14766 -2105
rect 14796 -1965 14852 -1941
rect 14796 -1999 14807 -1965
rect 14841 -1999 14852 -1965
rect 14796 -2051 14852 -1999
rect 14796 -2085 14807 -2051
rect 14841 -2085 14852 -2051
rect 14796 -2141 14852 -2085
rect 14882 -2071 14938 -1941
rect 14882 -2105 14893 -2071
rect 14927 -2105 14938 -2071
rect 14882 -2141 14938 -2105
rect 14968 -1965 15024 -1941
rect 14968 -1999 14979 -1965
rect 15013 -1999 15024 -1965
rect 14968 -2051 15024 -1999
rect 14968 -2085 14979 -2051
rect 15013 -2085 15024 -2051
rect 14968 -2141 15024 -2085
rect 15054 -2071 15110 -1941
rect 15054 -2105 15065 -2071
rect 15099 -2105 15110 -2071
rect 15054 -2141 15110 -2105
rect 15140 -1965 15196 -1941
rect 15140 -1999 15151 -1965
rect 15185 -1999 15196 -1965
rect 15140 -2051 15196 -1999
rect 15140 -2085 15151 -2051
rect 15185 -2085 15196 -2051
rect 15140 -2141 15196 -2085
rect 15226 -2071 15282 -1941
rect 15226 -2105 15237 -2071
rect 15271 -2105 15282 -2071
rect 15226 -2141 15282 -2105
rect 15312 -1965 15368 -1941
rect 15312 -1999 15323 -1965
rect 15357 -1999 15368 -1965
rect 15312 -2051 15368 -1999
rect 15312 -2085 15323 -2051
rect 15357 -2085 15368 -2051
rect 15312 -2141 15368 -2085
rect 15398 -2071 15451 -1941
rect 15398 -2105 15409 -2071
rect 15443 -2105 15451 -2071
rect 15398 -2141 15451 -2105
rect 15614 -1993 15666 -1967
rect 15614 -2027 15622 -1993
rect 15656 -2027 15666 -1993
rect 15614 -2095 15666 -2027
rect 15614 -2129 15622 -2095
rect 15656 -2129 15666 -2095
rect 15614 -2141 15666 -2129
rect 16612 -1993 16664 -1967
rect 16612 -2027 16622 -1993
rect 16656 -2027 16664 -1993
rect 16612 -2095 16664 -2027
rect 16612 -2129 16622 -2095
rect 16656 -2129 16664 -2095
rect 16612 -2141 16664 -2129
rect -2970 -2247 -2918 -2235
rect -2970 -2281 -2962 -2247
rect -2928 -2281 -2918 -2247
rect -2970 -2349 -2918 -2281
rect -2970 -2383 -2962 -2349
rect -2928 -2383 -2918 -2349
rect -2970 -2409 -2918 -2383
rect -2340 -2247 -2288 -2235
rect -2340 -2281 -2330 -2247
rect -2296 -2281 -2288 -2247
rect -1590 -2247 -1538 -2235
rect -2340 -2349 -2288 -2281
rect -2340 -2383 -2330 -2349
rect -2296 -2383 -2288 -2349
rect -2340 -2409 -2288 -2383
rect -1590 -2281 -1582 -2247
rect -1548 -2281 -1538 -2247
rect -1590 -2349 -1538 -2281
rect -1590 -2383 -1582 -2349
rect -1548 -2383 -1538 -2349
rect -1590 -2409 -1538 -2383
rect -960 -2247 -908 -2235
rect -960 -2281 -950 -2247
rect -916 -2281 -908 -2247
rect -960 -2349 -908 -2281
rect -960 -2383 -950 -2349
rect -916 -2383 -908 -2349
rect -960 -2409 -908 -2383
rect -854 -2247 -802 -2235
rect -854 -2281 -846 -2247
rect -812 -2281 -802 -2247
rect -854 -2349 -802 -2281
rect -854 -2383 -846 -2349
rect -812 -2383 -802 -2349
rect -854 -2409 -802 -2383
rect -224 -2247 -172 -2235
rect -224 -2281 -214 -2247
rect -180 -2281 -172 -2247
rect -26 -2247 26 -2235
rect -224 -2349 -172 -2281
rect -224 -2383 -214 -2349
rect -180 -2383 -172 -2349
rect -224 -2409 -172 -2383
rect -26 -2281 -18 -2247
rect 16 -2281 26 -2247
rect -26 -2349 26 -2281
rect -26 -2383 -18 -2349
rect 16 -2383 26 -2349
rect -26 -2409 26 -2383
rect 236 -2247 288 -2235
rect 236 -2281 246 -2247
rect 280 -2281 288 -2247
rect 236 -2349 288 -2281
rect 236 -2383 246 -2349
rect 280 -2383 288 -2349
rect 236 -2409 288 -2383
rect 434 -2254 488 -2235
rect 434 -2288 443 -2254
rect 477 -2288 488 -2254
rect 434 -2322 488 -2288
rect 434 -2356 443 -2322
rect 477 -2356 488 -2322
rect 434 -2435 488 -2356
rect 518 -2254 590 -2235
rect 518 -2288 543 -2254
rect 577 -2288 590 -2254
rect 518 -2322 590 -2288
rect 518 -2356 543 -2322
rect 577 -2356 590 -2322
rect 518 -2399 590 -2356
rect 690 -2254 743 -2235
rect 690 -2288 701 -2254
rect 735 -2288 743 -2254
rect 690 -2322 743 -2288
rect 690 -2356 701 -2322
rect 735 -2356 743 -2322
rect 690 -2399 743 -2356
rect 797 -2255 850 -2235
rect 797 -2289 805 -2255
rect 839 -2289 850 -2255
rect 797 -2323 850 -2289
rect 797 -2357 805 -2323
rect 839 -2357 850 -2323
rect 797 -2399 850 -2357
rect 950 -2254 1015 -2235
rect 950 -2288 961 -2254
rect 995 -2288 1015 -2254
rect 950 -2322 1015 -2288
rect 950 -2356 961 -2322
rect 995 -2356 1015 -2322
rect 950 -2399 1015 -2356
rect 518 -2435 568 -2399
rect 965 -2435 1015 -2399
rect 1045 -2255 1116 -2235
rect 1262 -2247 1314 -2235
rect 1045 -2289 1059 -2255
rect 1093 -2289 1116 -2255
rect 1045 -2323 1116 -2289
rect 1045 -2357 1059 -2323
rect 1093 -2357 1116 -2323
rect 1045 -2435 1116 -2357
rect 1262 -2281 1270 -2247
rect 1304 -2281 1314 -2247
rect 1262 -2349 1314 -2281
rect 1262 -2383 1270 -2349
rect 1304 -2383 1314 -2349
rect 1262 -2409 1314 -2383
rect 1524 -2247 1576 -2235
rect 1524 -2281 1534 -2247
rect 1568 -2281 1576 -2247
rect 1722 -2247 1774 -2235
rect 1524 -2349 1576 -2281
rect 1524 -2383 1534 -2349
rect 1568 -2383 1576 -2349
rect 1524 -2409 1576 -2383
rect 1722 -2281 1730 -2247
rect 1764 -2281 1774 -2247
rect 1722 -2349 1774 -2281
rect 1722 -2383 1730 -2349
rect 1764 -2383 1774 -2349
rect 1722 -2409 1774 -2383
rect 2352 -2247 2404 -2235
rect 2352 -2281 2362 -2247
rect 2396 -2281 2404 -2247
rect 2550 -2247 2602 -2235
rect 2352 -2349 2404 -2281
rect 2352 -2383 2362 -2349
rect 2396 -2383 2404 -2349
rect 2352 -2409 2404 -2383
rect 2550 -2281 2558 -2247
rect 2592 -2281 2602 -2247
rect 2550 -2349 2602 -2281
rect 2550 -2383 2558 -2349
rect 2592 -2383 2602 -2349
rect 2550 -2409 2602 -2383
rect 2812 -2247 2864 -2235
rect 2812 -2281 2822 -2247
rect 2856 -2281 2864 -2247
rect 2812 -2349 2864 -2281
rect 2812 -2383 2822 -2349
rect 2856 -2383 2864 -2349
rect 2812 -2409 2864 -2383
rect 3010 -2254 3064 -2235
rect 3010 -2288 3019 -2254
rect 3053 -2288 3064 -2254
rect 3010 -2322 3064 -2288
rect 3010 -2356 3019 -2322
rect 3053 -2356 3064 -2322
rect 3010 -2435 3064 -2356
rect 3094 -2254 3166 -2235
rect 3094 -2288 3119 -2254
rect 3153 -2288 3166 -2254
rect 3094 -2322 3166 -2288
rect 3094 -2356 3119 -2322
rect 3153 -2356 3166 -2322
rect 3094 -2399 3166 -2356
rect 3266 -2254 3319 -2235
rect 3266 -2288 3277 -2254
rect 3311 -2288 3319 -2254
rect 3266 -2322 3319 -2288
rect 3266 -2356 3277 -2322
rect 3311 -2356 3319 -2322
rect 3266 -2399 3319 -2356
rect 3373 -2255 3426 -2235
rect 3373 -2289 3381 -2255
rect 3415 -2289 3426 -2255
rect 3373 -2323 3426 -2289
rect 3373 -2357 3381 -2323
rect 3415 -2357 3426 -2323
rect 3373 -2399 3426 -2357
rect 3526 -2254 3591 -2235
rect 3526 -2288 3537 -2254
rect 3571 -2288 3591 -2254
rect 3526 -2322 3591 -2288
rect 3526 -2356 3537 -2322
rect 3571 -2356 3591 -2322
rect 3526 -2399 3591 -2356
rect 3094 -2435 3144 -2399
rect 3541 -2435 3591 -2399
rect 3621 -2255 3692 -2235
rect 3838 -2247 3890 -2235
rect 3621 -2289 3635 -2255
rect 3669 -2289 3692 -2255
rect 3621 -2323 3692 -2289
rect 3621 -2357 3635 -2323
rect 3669 -2357 3692 -2323
rect 3621 -2435 3692 -2357
rect 3838 -2281 3846 -2247
rect 3880 -2281 3890 -2247
rect 3838 -2349 3890 -2281
rect 3838 -2383 3846 -2349
rect 3880 -2383 3890 -2349
rect 3838 -2409 3890 -2383
rect 4100 -2247 4152 -2235
rect 4100 -2281 4110 -2247
rect 4144 -2281 4152 -2247
rect 4298 -2247 4350 -2235
rect 4100 -2349 4152 -2281
rect 4100 -2383 4110 -2349
rect 4144 -2383 4152 -2349
rect 4100 -2409 4152 -2383
rect 4298 -2281 4306 -2247
rect 4340 -2281 4350 -2247
rect 4298 -2349 4350 -2281
rect 4298 -2383 4306 -2349
rect 4340 -2383 4350 -2349
rect 4298 -2409 4350 -2383
rect 4928 -2247 4980 -2235
rect 4928 -2281 4938 -2247
rect 4972 -2281 4980 -2247
rect 5126 -2247 5178 -2235
rect 4928 -2349 4980 -2281
rect 4928 -2383 4938 -2349
rect 4972 -2383 4980 -2349
rect 4928 -2409 4980 -2383
rect 5126 -2281 5134 -2247
rect 5168 -2281 5178 -2247
rect 5126 -2349 5178 -2281
rect 5126 -2383 5134 -2349
rect 5168 -2383 5178 -2349
rect 5126 -2409 5178 -2383
rect 5388 -2247 5440 -2235
rect 5388 -2281 5398 -2247
rect 5432 -2281 5440 -2247
rect 5388 -2349 5440 -2281
rect 5388 -2383 5398 -2349
rect 5432 -2383 5440 -2349
rect 5388 -2409 5440 -2383
rect 5586 -2254 5640 -2235
rect 5586 -2288 5595 -2254
rect 5629 -2288 5640 -2254
rect 5586 -2322 5640 -2288
rect 5586 -2356 5595 -2322
rect 5629 -2356 5640 -2322
rect 5586 -2435 5640 -2356
rect 5670 -2254 5742 -2235
rect 5670 -2288 5695 -2254
rect 5729 -2288 5742 -2254
rect 5670 -2322 5742 -2288
rect 5670 -2356 5695 -2322
rect 5729 -2356 5742 -2322
rect 5670 -2399 5742 -2356
rect 5842 -2254 5895 -2235
rect 5842 -2288 5853 -2254
rect 5887 -2288 5895 -2254
rect 5842 -2322 5895 -2288
rect 5842 -2356 5853 -2322
rect 5887 -2356 5895 -2322
rect 5842 -2399 5895 -2356
rect 5949 -2255 6002 -2235
rect 5949 -2289 5957 -2255
rect 5991 -2289 6002 -2255
rect 5949 -2323 6002 -2289
rect 5949 -2357 5957 -2323
rect 5991 -2357 6002 -2323
rect 5949 -2399 6002 -2357
rect 6102 -2254 6167 -2235
rect 6102 -2288 6113 -2254
rect 6147 -2288 6167 -2254
rect 6102 -2322 6167 -2288
rect 6102 -2356 6113 -2322
rect 6147 -2356 6167 -2322
rect 6102 -2399 6167 -2356
rect 5670 -2435 5720 -2399
rect 6117 -2435 6167 -2399
rect 6197 -2255 6268 -2235
rect 6414 -2247 6466 -2235
rect 6197 -2289 6211 -2255
rect 6245 -2289 6268 -2255
rect 6197 -2323 6268 -2289
rect 6197 -2357 6211 -2323
rect 6245 -2357 6268 -2323
rect 6197 -2435 6268 -2357
rect 6414 -2281 6422 -2247
rect 6456 -2281 6466 -2247
rect 6414 -2349 6466 -2281
rect 6414 -2383 6422 -2349
rect 6456 -2383 6466 -2349
rect 6414 -2409 6466 -2383
rect 6676 -2247 6728 -2235
rect 6676 -2281 6686 -2247
rect 6720 -2281 6728 -2247
rect 6874 -2247 6926 -2235
rect 6676 -2349 6728 -2281
rect 6676 -2383 6686 -2349
rect 6720 -2383 6728 -2349
rect 6676 -2409 6728 -2383
rect 6874 -2281 6882 -2247
rect 6916 -2281 6926 -2247
rect 6874 -2349 6926 -2281
rect 6874 -2383 6882 -2349
rect 6916 -2383 6926 -2349
rect 6874 -2409 6926 -2383
rect 7504 -2247 7556 -2235
rect 7504 -2281 7514 -2247
rect 7548 -2281 7556 -2247
rect 7702 -2247 7754 -2235
rect 7504 -2349 7556 -2281
rect 7504 -2383 7514 -2349
rect 7548 -2383 7556 -2349
rect 7504 -2409 7556 -2383
rect 7702 -2281 7710 -2247
rect 7744 -2281 7754 -2247
rect 7702 -2349 7754 -2281
rect 7702 -2383 7710 -2349
rect 7744 -2383 7754 -2349
rect 7702 -2409 7754 -2383
rect 7964 -2247 8016 -2235
rect 7964 -2281 7974 -2247
rect 8008 -2281 8016 -2247
rect 7964 -2349 8016 -2281
rect 7964 -2383 7974 -2349
rect 8008 -2383 8016 -2349
rect 7964 -2409 8016 -2383
rect 8162 -2254 8216 -2235
rect 8162 -2288 8171 -2254
rect 8205 -2288 8216 -2254
rect 8162 -2322 8216 -2288
rect 8162 -2356 8171 -2322
rect 8205 -2356 8216 -2322
rect 8162 -2435 8216 -2356
rect 8246 -2254 8318 -2235
rect 8246 -2288 8271 -2254
rect 8305 -2288 8318 -2254
rect 8246 -2322 8318 -2288
rect 8246 -2356 8271 -2322
rect 8305 -2356 8318 -2322
rect 8246 -2399 8318 -2356
rect 8418 -2254 8471 -2235
rect 8418 -2288 8429 -2254
rect 8463 -2288 8471 -2254
rect 8418 -2322 8471 -2288
rect 8418 -2356 8429 -2322
rect 8463 -2356 8471 -2322
rect 8418 -2399 8471 -2356
rect 8525 -2255 8578 -2235
rect 8525 -2289 8533 -2255
rect 8567 -2289 8578 -2255
rect 8525 -2323 8578 -2289
rect 8525 -2357 8533 -2323
rect 8567 -2357 8578 -2323
rect 8525 -2399 8578 -2357
rect 8678 -2254 8743 -2235
rect 8678 -2288 8689 -2254
rect 8723 -2288 8743 -2254
rect 8678 -2322 8743 -2288
rect 8678 -2356 8689 -2322
rect 8723 -2356 8743 -2322
rect 8678 -2399 8743 -2356
rect 8246 -2435 8296 -2399
rect 8693 -2435 8743 -2399
rect 8773 -2255 8844 -2235
rect 8990 -2247 9042 -2235
rect 8773 -2289 8787 -2255
rect 8821 -2289 8844 -2255
rect 8773 -2323 8844 -2289
rect 8773 -2357 8787 -2323
rect 8821 -2357 8844 -2323
rect 8773 -2435 8844 -2357
rect 8990 -2281 8998 -2247
rect 9032 -2281 9042 -2247
rect 8990 -2349 9042 -2281
rect 8990 -2383 8998 -2349
rect 9032 -2383 9042 -2349
rect 8990 -2409 9042 -2383
rect 9252 -2247 9304 -2235
rect 9252 -2281 9262 -2247
rect 9296 -2281 9304 -2247
rect 9450 -2247 9502 -2235
rect 9252 -2349 9304 -2281
rect 9252 -2383 9262 -2349
rect 9296 -2383 9304 -2349
rect 9252 -2409 9304 -2383
rect 9450 -2281 9458 -2247
rect 9492 -2281 9502 -2247
rect 9450 -2349 9502 -2281
rect 9450 -2383 9458 -2349
rect 9492 -2383 9502 -2349
rect 9450 -2409 9502 -2383
rect 10080 -2247 10132 -2235
rect 10080 -2281 10090 -2247
rect 10124 -2281 10132 -2247
rect 10370 -2247 10422 -2235
rect 10080 -2349 10132 -2281
rect 10080 -2383 10090 -2349
rect 10124 -2383 10132 -2349
rect 10080 -2409 10132 -2383
rect 10370 -2281 10378 -2247
rect 10412 -2281 10422 -2247
rect 10370 -2349 10422 -2281
rect 10370 -2383 10378 -2349
rect 10412 -2383 10422 -2349
rect 10370 -2409 10422 -2383
rect 10632 -2247 10684 -2235
rect 10632 -2281 10642 -2247
rect 10676 -2281 10684 -2247
rect 10632 -2349 10684 -2281
rect 10632 -2383 10642 -2349
rect 10676 -2383 10684 -2349
rect 10632 -2409 10684 -2383
rect 10738 -2254 10792 -2235
rect 10738 -2288 10747 -2254
rect 10781 -2288 10792 -2254
rect 10738 -2322 10792 -2288
rect 10738 -2356 10747 -2322
rect 10781 -2356 10792 -2322
rect 10738 -2435 10792 -2356
rect 10822 -2254 10894 -2235
rect 10822 -2288 10847 -2254
rect 10881 -2288 10894 -2254
rect 10822 -2322 10894 -2288
rect 10822 -2356 10847 -2322
rect 10881 -2356 10894 -2322
rect 10822 -2399 10894 -2356
rect 10994 -2254 11047 -2235
rect 10994 -2288 11005 -2254
rect 11039 -2288 11047 -2254
rect 10994 -2322 11047 -2288
rect 10994 -2356 11005 -2322
rect 11039 -2356 11047 -2322
rect 10994 -2399 11047 -2356
rect 11101 -2255 11154 -2235
rect 11101 -2289 11109 -2255
rect 11143 -2289 11154 -2255
rect 11101 -2323 11154 -2289
rect 11101 -2357 11109 -2323
rect 11143 -2357 11154 -2323
rect 11101 -2399 11154 -2357
rect 11254 -2254 11319 -2235
rect 11254 -2288 11265 -2254
rect 11299 -2288 11319 -2254
rect 11254 -2322 11319 -2288
rect 11254 -2356 11265 -2322
rect 11299 -2356 11319 -2322
rect 11254 -2399 11319 -2356
rect 10822 -2435 10872 -2399
rect 11269 -2435 11319 -2399
rect 11349 -2255 11420 -2235
rect 11658 -2247 11710 -2235
rect 11349 -2289 11363 -2255
rect 11397 -2289 11420 -2255
rect 11349 -2323 11420 -2289
rect 11349 -2357 11363 -2323
rect 11397 -2357 11420 -2323
rect 11349 -2435 11420 -2357
rect 11658 -2281 11666 -2247
rect 11700 -2281 11710 -2247
rect 11658 -2349 11710 -2281
rect 11658 -2383 11666 -2349
rect 11700 -2383 11710 -2349
rect 11658 -2409 11710 -2383
rect 11920 -2247 11972 -2235
rect 11920 -2281 11930 -2247
rect 11964 -2281 11972 -2247
rect 11920 -2349 11972 -2281
rect 11920 -2383 11930 -2349
rect 11964 -2383 11972 -2349
rect 11920 -2409 11972 -2383
rect 12486 -2254 12547 -2235
rect 12486 -2288 12502 -2254
rect 12536 -2288 12547 -2254
rect 12486 -2322 12547 -2288
rect 12486 -2356 12502 -2322
rect 12536 -2356 12547 -2322
rect 12486 -2435 12547 -2356
rect 12577 -2261 12633 -2235
rect 12577 -2295 12588 -2261
rect 12622 -2295 12633 -2261
rect 12577 -2349 12633 -2295
rect 12577 -2383 12588 -2349
rect 12622 -2383 12633 -2349
rect 12577 -2435 12633 -2383
rect 12663 -2254 12719 -2235
rect 12663 -2288 12674 -2254
rect 12708 -2288 12719 -2254
rect 12663 -2322 12719 -2288
rect 12663 -2356 12674 -2322
rect 12708 -2356 12719 -2322
rect 12663 -2435 12719 -2356
rect 12749 -2261 12805 -2235
rect 12749 -2295 12760 -2261
rect 12794 -2295 12805 -2261
rect 12749 -2349 12805 -2295
rect 12749 -2383 12760 -2349
rect 12794 -2383 12805 -2349
rect 12749 -2435 12805 -2383
rect 12835 -2254 12891 -2235
rect 12835 -2288 12846 -2254
rect 12880 -2288 12891 -2254
rect 12835 -2322 12891 -2288
rect 12835 -2356 12846 -2322
rect 12880 -2356 12891 -2322
rect 12835 -2435 12891 -2356
rect 12921 -2261 12977 -2235
rect 12921 -2295 12932 -2261
rect 12966 -2295 12977 -2261
rect 12921 -2349 12977 -2295
rect 12921 -2383 12932 -2349
rect 12966 -2383 12977 -2349
rect 12921 -2435 12977 -2383
rect 13007 -2254 13076 -2235
rect 13222 -2247 13274 -2235
rect 13007 -2288 13018 -2254
rect 13052 -2288 13076 -2254
rect 13007 -2322 13076 -2288
rect 13007 -2356 13018 -2322
rect 13052 -2356 13076 -2322
rect 13007 -2435 13076 -2356
rect 13222 -2281 13230 -2247
rect 13264 -2281 13274 -2247
rect 13222 -2349 13274 -2281
rect 13222 -2383 13230 -2349
rect 13264 -2383 13274 -2349
rect 13222 -2409 13274 -2383
rect 13484 -2247 13536 -2235
rect 13484 -2281 13494 -2247
rect 13528 -2281 13536 -2247
rect 13682 -2247 13735 -2235
rect 13484 -2349 13536 -2281
rect 13484 -2383 13494 -2349
rect 13528 -2383 13536 -2349
rect 13484 -2409 13536 -2383
rect 13682 -2281 13690 -2247
rect 13724 -2281 13735 -2247
rect 13682 -2315 13735 -2281
rect 13682 -2349 13690 -2315
rect 13724 -2349 13735 -2315
rect 13682 -2435 13735 -2349
rect 13765 -2255 13821 -2235
rect 13765 -2289 13776 -2255
rect 13810 -2289 13821 -2255
rect 13765 -2323 13821 -2289
rect 13765 -2357 13776 -2323
rect 13810 -2357 13821 -2323
rect 13765 -2435 13821 -2357
rect 13851 -2247 13907 -2235
rect 13851 -2281 13862 -2247
rect 13896 -2281 13907 -2247
rect 13851 -2315 13907 -2281
rect 13851 -2349 13862 -2315
rect 13896 -2349 13907 -2315
rect 13851 -2435 13907 -2349
rect 13937 -2263 13993 -2235
rect 13937 -2297 13948 -2263
rect 13982 -2297 13993 -2263
rect 13937 -2331 13993 -2297
rect 13937 -2365 13948 -2331
rect 13982 -2365 13993 -2331
rect 13937 -2435 13993 -2365
rect 14023 -2247 14079 -2235
rect 14023 -2281 14034 -2247
rect 14068 -2281 14079 -2247
rect 14023 -2315 14079 -2281
rect 14023 -2349 14034 -2315
rect 14068 -2349 14079 -2315
rect 14023 -2435 14079 -2349
rect 14109 -2291 14165 -2235
rect 14109 -2325 14120 -2291
rect 14154 -2325 14165 -2291
rect 14109 -2377 14165 -2325
rect 14109 -2411 14120 -2377
rect 14154 -2411 14165 -2377
rect 14109 -2435 14165 -2411
rect 14195 -2271 14251 -2235
rect 14195 -2305 14206 -2271
rect 14240 -2305 14251 -2271
rect 14195 -2435 14251 -2305
rect 14281 -2291 14337 -2235
rect 14281 -2325 14292 -2291
rect 14326 -2325 14337 -2291
rect 14281 -2377 14337 -2325
rect 14281 -2411 14292 -2377
rect 14326 -2411 14337 -2377
rect 14281 -2435 14337 -2411
rect 14367 -2271 14423 -2235
rect 14367 -2305 14378 -2271
rect 14412 -2305 14423 -2271
rect 14367 -2435 14423 -2305
rect 14453 -2291 14509 -2235
rect 14453 -2325 14464 -2291
rect 14498 -2325 14509 -2291
rect 14453 -2377 14509 -2325
rect 14453 -2411 14464 -2377
rect 14498 -2411 14509 -2377
rect 14453 -2435 14509 -2411
rect 14539 -2271 14595 -2235
rect 14539 -2305 14550 -2271
rect 14584 -2305 14595 -2271
rect 14539 -2435 14595 -2305
rect 14625 -2291 14681 -2235
rect 14625 -2325 14636 -2291
rect 14670 -2325 14681 -2291
rect 14625 -2377 14681 -2325
rect 14625 -2411 14636 -2377
rect 14670 -2411 14681 -2377
rect 14625 -2435 14681 -2411
rect 14711 -2271 14766 -2235
rect 14711 -2305 14722 -2271
rect 14756 -2305 14766 -2271
rect 14711 -2435 14766 -2305
rect 14796 -2291 14852 -2235
rect 14796 -2325 14807 -2291
rect 14841 -2325 14852 -2291
rect 14796 -2377 14852 -2325
rect 14796 -2411 14807 -2377
rect 14841 -2411 14852 -2377
rect 14796 -2435 14852 -2411
rect 14882 -2271 14938 -2235
rect 14882 -2305 14893 -2271
rect 14927 -2305 14938 -2271
rect 14882 -2435 14938 -2305
rect 14968 -2291 15024 -2235
rect 14968 -2325 14979 -2291
rect 15013 -2325 15024 -2291
rect 14968 -2377 15024 -2325
rect 14968 -2411 14979 -2377
rect 15013 -2411 15024 -2377
rect 14968 -2435 15024 -2411
rect 15054 -2271 15110 -2235
rect 15054 -2305 15065 -2271
rect 15099 -2305 15110 -2271
rect 15054 -2435 15110 -2305
rect 15140 -2291 15196 -2235
rect 15140 -2325 15151 -2291
rect 15185 -2325 15196 -2291
rect 15140 -2377 15196 -2325
rect 15140 -2411 15151 -2377
rect 15185 -2411 15196 -2377
rect 15140 -2435 15196 -2411
rect 15226 -2271 15282 -2235
rect 15226 -2305 15237 -2271
rect 15271 -2305 15282 -2271
rect 15226 -2435 15282 -2305
rect 15312 -2291 15368 -2235
rect 15312 -2325 15323 -2291
rect 15357 -2325 15368 -2291
rect 15312 -2377 15368 -2325
rect 15312 -2411 15323 -2377
rect 15357 -2411 15368 -2377
rect 15312 -2435 15368 -2411
rect 15398 -2271 15451 -2235
rect 15614 -2247 15666 -2235
rect 15398 -2305 15409 -2271
rect 15443 -2305 15451 -2271
rect 15398 -2435 15451 -2305
rect 15614 -2281 15622 -2247
rect 15656 -2281 15666 -2247
rect 15614 -2349 15666 -2281
rect 15614 -2383 15622 -2349
rect 15656 -2383 15666 -2349
rect 15614 -2409 15666 -2383
rect 16612 -2247 16664 -2235
rect 16612 -2281 16622 -2247
rect 16656 -2281 16664 -2247
rect 16612 -2349 16664 -2281
rect 16612 -2383 16622 -2349
rect 16656 -2383 16664 -2349
rect 16612 -2409 16664 -2383
rect -2970 -3081 -2918 -3055
rect -2970 -3115 -2962 -3081
rect -2928 -3115 -2918 -3081
rect -2970 -3183 -2918 -3115
rect -2970 -3217 -2962 -3183
rect -2928 -3217 -2918 -3183
rect -2970 -3229 -2918 -3217
rect -2340 -3081 -2288 -3055
rect -2340 -3115 -2330 -3081
rect -2296 -3115 -2288 -3081
rect -2340 -3183 -2288 -3115
rect -2340 -3217 -2330 -3183
rect -2296 -3217 -2288 -3183
rect -1958 -3081 -1906 -3061
rect -1958 -3115 -1950 -3081
rect -1916 -3115 -1906 -3081
rect -1958 -3183 -1906 -3115
rect -2340 -3229 -2288 -3217
rect -1958 -3217 -1950 -3183
rect -1916 -3217 -1906 -3183
rect -1958 -3229 -1906 -3217
rect -1876 -3081 -1822 -3061
rect -1876 -3115 -1866 -3081
rect -1832 -3115 -1822 -3081
rect -1876 -3183 -1822 -3115
rect -1876 -3217 -1866 -3183
rect -1832 -3217 -1822 -3183
rect -1876 -3229 -1822 -3217
rect -1792 -3081 -1736 -3061
rect -1792 -3115 -1782 -3081
rect -1748 -3115 -1736 -3081
rect -1792 -3183 -1736 -3115
rect -1792 -3217 -1782 -3183
rect -1748 -3217 -1736 -3183
rect -1590 -3081 -1538 -3055
rect -1590 -3115 -1582 -3081
rect -1548 -3115 -1538 -3081
rect -1590 -3183 -1538 -3115
rect -1792 -3229 -1736 -3217
rect -1590 -3217 -1582 -3183
rect -1548 -3217 -1538 -3183
rect -1590 -3229 -1538 -3217
rect -960 -3081 -908 -3055
rect -960 -3115 -950 -3081
rect -916 -3115 -908 -3081
rect -960 -3183 -908 -3115
rect -960 -3217 -950 -3183
rect -916 -3217 -908 -3183
rect -960 -3229 -908 -3217
rect -854 -3081 -802 -3055
rect -854 -3115 -846 -3081
rect -812 -3115 -802 -3081
rect -854 -3183 -802 -3115
rect -854 -3217 -846 -3183
rect -812 -3217 -802 -3183
rect -854 -3229 -802 -3217
rect -224 -3081 -172 -3055
rect -224 -3115 -214 -3081
rect -180 -3115 -172 -3081
rect -224 -3183 -172 -3115
rect -224 -3217 -214 -3183
rect -180 -3217 -172 -3183
rect -26 -3081 26 -3055
rect -26 -3115 -18 -3081
rect 16 -3115 26 -3081
rect -26 -3183 26 -3115
rect -224 -3229 -172 -3217
rect -26 -3217 -18 -3183
rect 16 -3217 26 -3183
rect -26 -3229 26 -3217
rect 236 -3081 288 -3055
rect 236 -3115 246 -3081
rect 280 -3115 288 -3081
rect 236 -3183 288 -3115
rect 236 -3217 246 -3183
rect 280 -3217 288 -3183
rect 434 -3107 505 -3029
rect 434 -3141 457 -3107
rect 491 -3141 505 -3107
rect 434 -3175 505 -3141
rect 434 -3209 457 -3175
rect 491 -3209 505 -3175
rect 236 -3229 288 -3217
rect 434 -3229 505 -3209
rect 535 -3065 585 -3029
rect 982 -3065 1032 -3029
rect 535 -3108 600 -3065
rect 535 -3142 555 -3108
rect 589 -3142 600 -3108
rect 535 -3176 600 -3142
rect 535 -3210 555 -3176
rect 589 -3210 600 -3176
rect 535 -3229 600 -3210
rect 700 -3107 753 -3065
rect 700 -3141 711 -3107
rect 745 -3141 753 -3107
rect 700 -3175 753 -3141
rect 700 -3209 711 -3175
rect 745 -3209 753 -3175
rect 700 -3229 753 -3209
rect 807 -3108 860 -3065
rect 807 -3142 815 -3108
rect 849 -3142 860 -3108
rect 807 -3176 860 -3142
rect 807 -3210 815 -3176
rect 849 -3210 860 -3176
rect 807 -3229 860 -3210
rect 960 -3108 1032 -3065
rect 960 -3142 973 -3108
rect 1007 -3142 1032 -3108
rect 960 -3176 1032 -3142
rect 960 -3210 973 -3176
rect 1007 -3210 1032 -3176
rect 960 -3229 1032 -3210
rect 1062 -3108 1116 -3029
rect 1062 -3142 1073 -3108
rect 1107 -3142 1116 -3108
rect 1062 -3176 1116 -3142
rect 1062 -3210 1073 -3176
rect 1107 -3210 1116 -3176
rect 1062 -3229 1116 -3210
rect 1262 -3081 1314 -3055
rect 1262 -3115 1270 -3081
rect 1304 -3115 1314 -3081
rect 1262 -3183 1314 -3115
rect 1262 -3217 1270 -3183
rect 1304 -3217 1314 -3183
rect 1262 -3229 1314 -3217
rect 1524 -3081 1576 -3055
rect 1524 -3115 1534 -3081
rect 1568 -3115 1576 -3081
rect 1524 -3183 1576 -3115
rect 1524 -3217 1534 -3183
rect 1568 -3217 1576 -3183
rect 1722 -3081 1774 -3055
rect 1722 -3115 1730 -3081
rect 1764 -3115 1774 -3081
rect 1722 -3183 1774 -3115
rect 1524 -3229 1576 -3217
rect 1722 -3217 1730 -3183
rect 1764 -3217 1774 -3183
rect 1722 -3229 1774 -3217
rect 2352 -3081 2404 -3055
rect 2352 -3115 2362 -3081
rect 2396 -3115 2404 -3081
rect 2352 -3183 2404 -3115
rect 2352 -3217 2362 -3183
rect 2396 -3217 2404 -3183
rect 2550 -3081 2602 -3055
rect 2550 -3115 2558 -3081
rect 2592 -3115 2602 -3081
rect 2550 -3183 2602 -3115
rect 2352 -3229 2404 -3217
rect 2550 -3217 2558 -3183
rect 2592 -3217 2602 -3183
rect 2550 -3229 2602 -3217
rect 2812 -3081 2864 -3055
rect 2812 -3115 2822 -3081
rect 2856 -3115 2864 -3081
rect 2812 -3183 2864 -3115
rect 2812 -3217 2822 -3183
rect 2856 -3217 2864 -3183
rect 3010 -3107 3081 -3029
rect 3010 -3141 3033 -3107
rect 3067 -3141 3081 -3107
rect 3010 -3175 3081 -3141
rect 3010 -3209 3033 -3175
rect 3067 -3209 3081 -3175
rect 2812 -3229 2864 -3217
rect 3010 -3229 3081 -3209
rect 3111 -3065 3161 -3029
rect 3558 -3065 3608 -3029
rect 3111 -3108 3176 -3065
rect 3111 -3142 3131 -3108
rect 3165 -3142 3176 -3108
rect 3111 -3176 3176 -3142
rect 3111 -3210 3131 -3176
rect 3165 -3210 3176 -3176
rect 3111 -3229 3176 -3210
rect 3276 -3107 3329 -3065
rect 3276 -3141 3287 -3107
rect 3321 -3141 3329 -3107
rect 3276 -3175 3329 -3141
rect 3276 -3209 3287 -3175
rect 3321 -3209 3329 -3175
rect 3276 -3229 3329 -3209
rect 3383 -3108 3436 -3065
rect 3383 -3142 3391 -3108
rect 3425 -3142 3436 -3108
rect 3383 -3176 3436 -3142
rect 3383 -3210 3391 -3176
rect 3425 -3210 3436 -3176
rect 3383 -3229 3436 -3210
rect 3536 -3108 3608 -3065
rect 3536 -3142 3549 -3108
rect 3583 -3142 3608 -3108
rect 3536 -3176 3608 -3142
rect 3536 -3210 3549 -3176
rect 3583 -3210 3608 -3176
rect 3536 -3229 3608 -3210
rect 3638 -3108 3692 -3029
rect 3638 -3142 3649 -3108
rect 3683 -3142 3692 -3108
rect 3638 -3176 3692 -3142
rect 3638 -3210 3649 -3176
rect 3683 -3210 3692 -3176
rect 3638 -3229 3692 -3210
rect 3838 -3081 3890 -3055
rect 3838 -3115 3846 -3081
rect 3880 -3115 3890 -3081
rect 3838 -3183 3890 -3115
rect 3838 -3217 3846 -3183
rect 3880 -3217 3890 -3183
rect 3838 -3229 3890 -3217
rect 4100 -3081 4152 -3055
rect 4100 -3115 4110 -3081
rect 4144 -3115 4152 -3081
rect 4100 -3183 4152 -3115
rect 4100 -3217 4110 -3183
rect 4144 -3217 4152 -3183
rect 4298 -3081 4350 -3055
rect 4298 -3115 4306 -3081
rect 4340 -3115 4350 -3081
rect 4298 -3183 4350 -3115
rect 4100 -3229 4152 -3217
rect 4298 -3217 4306 -3183
rect 4340 -3217 4350 -3183
rect 4298 -3229 4350 -3217
rect 4928 -3081 4980 -3055
rect 4928 -3115 4938 -3081
rect 4972 -3115 4980 -3081
rect 4928 -3183 4980 -3115
rect 4928 -3217 4938 -3183
rect 4972 -3217 4980 -3183
rect 5126 -3081 5178 -3055
rect 5126 -3115 5134 -3081
rect 5168 -3115 5178 -3081
rect 5126 -3183 5178 -3115
rect 4928 -3229 4980 -3217
rect 5126 -3217 5134 -3183
rect 5168 -3217 5178 -3183
rect 5126 -3229 5178 -3217
rect 5388 -3081 5440 -3055
rect 5388 -3115 5398 -3081
rect 5432 -3115 5440 -3081
rect 5388 -3183 5440 -3115
rect 5388 -3217 5398 -3183
rect 5432 -3217 5440 -3183
rect 5586 -3107 5657 -3029
rect 5586 -3141 5609 -3107
rect 5643 -3141 5657 -3107
rect 5586 -3175 5657 -3141
rect 5586 -3209 5609 -3175
rect 5643 -3209 5657 -3175
rect 5388 -3229 5440 -3217
rect 5586 -3229 5657 -3209
rect 5687 -3065 5737 -3029
rect 6134 -3065 6184 -3029
rect 5687 -3108 5752 -3065
rect 5687 -3142 5707 -3108
rect 5741 -3142 5752 -3108
rect 5687 -3176 5752 -3142
rect 5687 -3210 5707 -3176
rect 5741 -3210 5752 -3176
rect 5687 -3229 5752 -3210
rect 5852 -3107 5905 -3065
rect 5852 -3141 5863 -3107
rect 5897 -3141 5905 -3107
rect 5852 -3175 5905 -3141
rect 5852 -3209 5863 -3175
rect 5897 -3209 5905 -3175
rect 5852 -3229 5905 -3209
rect 5959 -3108 6012 -3065
rect 5959 -3142 5967 -3108
rect 6001 -3142 6012 -3108
rect 5959 -3176 6012 -3142
rect 5959 -3210 5967 -3176
rect 6001 -3210 6012 -3176
rect 5959 -3229 6012 -3210
rect 6112 -3108 6184 -3065
rect 6112 -3142 6125 -3108
rect 6159 -3142 6184 -3108
rect 6112 -3176 6184 -3142
rect 6112 -3210 6125 -3176
rect 6159 -3210 6184 -3176
rect 6112 -3229 6184 -3210
rect 6214 -3108 6268 -3029
rect 6214 -3142 6225 -3108
rect 6259 -3142 6268 -3108
rect 6214 -3176 6268 -3142
rect 6214 -3210 6225 -3176
rect 6259 -3210 6268 -3176
rect 6214 -3229 6268 -3210
rect 6414 -3081 6466 -3055
rect 6414 -3115 6422 -3081
rect 6456 -3115 6466 -3081
rect 6414 -3183 6466 -3115
rect 6414 -3217 6422 -3183
rect 6456 -3217 6466 -3183
rect 6414 -3229 6466 -3217
rect 6676 -3081 6728 -3055
rect 6676 -3115 6686 -3081
rect 6720 -3115 6728 -3081
rect 6676 -3183 6728 -3115
rect 6676 -3217 6686 -3183
rect 6720 -3217 6728 -3183
rect 6874 -3081 6926 -3055
rect 6874 -3115 6882 -3081
rect 6916 -3115 6926 -3081
rect 6874 -3183 6926 -3115
rect 6676 -3229 6728 -3217
rect 6874 -3217 6882 -3183
rect 6916 -3217 6926 -3183
rect 6874 -3229 6926 -3217
rect 7504 -3081 7556 -3055
rect 7504 -3115 7514 -3081
rect 7548 -3115 7556 -3081
rect 7504 -3183 7556 -3115
rect 7504 -3217 7514 -3183
rect 7548 -3217 7556 -3183
rect 7702 -3081 7754 -3055
rect 7702 -3115 7710 -3081
rect 7744 -3115 7754 -3081
rect 7702 -3183 7754 -3115
rect 7504 -3229 7556 -3217
rect 7702 -3217 7710 -3183
rect 7744 -3217 7754 -3183
rect 7702 -3229 7754 -3217
rect 7964 -3081 8016 -3055
rect 7964 -3115 7974 -3081
rect 8008 -3115 8016 -3081
rect 7964 -3183 8016 -3115
rect 7964 -3217 7974 -3183
rect 8008 -3217 8016 -3183
rect 8162 -3107 8233 -3029
rect 8162 -3141 8185 -3107
rect 8219 -3141 8233 -3107
rect 8162 -3175 8233 -3141
rect 8162 -3209 8185 -3175
rect 8219 -3209 8233 -3175
rect 7964 -3229 8016 -3217
rect 8162 -3229 8233 -3209
rect 8263 -3065 8313 -3029
rect 8710 -3065 8760 -3029
rect 8263 -3108 8328 -3065
rect 8263 -3142 8283 -3108
rect 8317 -3142 8328 -3108
rect 8263 -3176 8328 -3142
rect 8263 -3210 8283 -3176
rect 8317 -3210 8328 -3176
rect 8263 -3229 8328 -3210
rect 8428 -3107 8481 -3065
rect 8428 -3141 8439 -3107
rect 8473 -3141 8481 -3107
rect 8428 -3175 8481 -3141
rect 8428 -3209 8439 -3175
rect 8473 -3209 8481 -3175
rect 8428 -3229 8481 -3209
rect 8535 -3108 8588 -3065
rect 8535 -3142 8543 -3108
rect 8577 -3142 8588 -3108
rect 8535 -3176 8588 -3142
rect 8535 -3210 8543 -3176
rect 8577 -3210 8588 -3176
rect 8535 -3229 8588 -3210
rect 8688 -3108 8760 -3065
rect 8688 -3142 8701 -3108
rect 8735 -3142 8760 -3108
rect 8688 -3176 8760 -3142
rect 8688 -3210 8701 -3176
rect 8735 -3210 8760 -3176
rect 8688 -3229 8760 -3210
rect 8790 -3108 8844 -3029
rect 8790 -3142 8801 -3108
rect 8835 -3142 8844 -3108
rect 8790 -3176 8844 -3142
rect 8790 -3210 8801 -3176
rect 8835 -3210 8844 -3176
rect 8790 -3229 8844 -3210
rect 8990 -3081 9042 -3055
rect 8990 -3115 8998 -3081
rect 9032 -3115 9042 -3081
rect 8990 -3183 9042 -3115
rect 8990 -3217 8998 -3183
rect 9032 -3217 9042 -3183
rect 8990 -3229 9042 -3217
rect 9252 -3081 9304 -3055
rect 9252 -3115 9262 -3081
rect 9296 -3115 9304 -3081
rect 9252 -3183 9304 -3115
rect 9252 -3217 9262 -3183
rect 9296 -3217 9304 -3183
rect 9450 -3081 9502 -3055
rect 9450 -3115 9458 -3081
rect 9492 -3115 9502 -3081
rect 9450 -3183 9502 -3115
rect 9252 -3229 9304 -3217
rect 9450 -3217 9458 -3183
rect 9492 -3217 9502 -3183
rect 9450 -3229 9502 -3217
rect 10080 -3081 10132 -3055
rect 10080 -3115 10090 -3081
rect 10124 -3115 10132 -3081
rect 10080 -3183 10132 -3115
rect 10080 -3217 10090 -3183
rect 10124 -3217 10132 -3183
rect 10370 -3081 10422 -3055
rect 10370 -3115 10378 -3081
rect 10412 -3115 10422 -3081
rect 10370 -3183 10422 -3115
rect 10080 -3229 10132 -3217
rect 10370 -3217 10378 -3183
rect 10412 -3217 10422 -3183
rect 10370 -3229 10422 -3217
rect 10632 -3081 10684 -3055
rect 10632 -3115 10642 -3081
rect 10676 -3115 10684 -3081
rect 10632 -3183 10684 -3115
rect 10632 -3217 10642 -3183
rect 10676 -3217 10684 -3183
rect 10632 -3229 10684 -3217
rect 10738 -3107 10809 -3029
rect 10738 -3141 10761 -3107
rect 10795 -3141 10809 -3107
rect 10738 -3175 10809 -3141
rect 10738 -3209 10761 -3175
rect 10795 -3209 10809 -3175
rect 10738 -3229 10809 -3209
rect 10839 -3065 10889 -3029
rect 11286 -3065 11336 -3029
rect 10839 -3108 10904 -3065
rect 10839 -3142 10859 -3108
rect 10893 -3142 10904 -3108
rect 10839 -3176 10904 -3142
rect 10839 -3210 10859 -3176
rect 10893 -3210 10904 -3176
rect 10839 -3229 10904 -3210
rect 11004 -3107 11057 -3065
rect 11004 -3141 11015 -3107
rect 11049 -3141 11057 -3107
rect 11004 -3175 11057 -3141
rect 11004 -3209 11015 -3175
rect 11049 -3209 11057 -3175
rect 11004 -3229 11057 -3209
rect 11111 -3108 11164 -3065
rect 11111 -3142 11119 -3108
rect 11153 -3142 11164 -3108
rect 11111 -3176 11164 -3142
rect 11111 -3210 11119 -3176
rect 11153 -3210 11164 -3176
rect 11111 -3229 11164 -3210
rect 11264 -3108 11336 -3065
rect 11264 -3142 11277 -3108
rect 11311 -3142 11336 -3108
rect 11264 -3176 11336 -3142
rect 11264 -3210 11277 -3176
rect 11311 -3210 11336 -3176
rect 11264 -3229 11336 -3210
rect 11366 -3108 11420 -3029
rect 11366 -3142 11377 -3108
rect 11411 -3142 11420 -3108
rect 11366 -3176 11420 -3142
rect 11366 -3210 11377 -3176
rect 11411 -3210 11420 -3176
rect 11366 -3229 11420 -3210
rect 11658 -3081 11710 -3055
rect 11658 -3115 11666 -3081
rect 11700 -3115 11710 -3081
rect 11658 -3183 11710 -3115
rect 11658 -3217 11666 -3183
rect 11700 -3217 11710 -3183
rect 11658 -3229 11710 -3217
rect 11920 -3081 11972 -3055
rect 11920 -3115 11930 -3081
rect 11964 -3115 11972 -3081
rect 11920 -3183 11972 -3115
rect 11920 -3217 11930 -3183
rect 11964 -3217 11972 -3183
rect 13590 -3081 13642 -3055
rect 13590 -3115 13598 -3081
rect 13632 -3115 13642 -3081
rect 13590 -3183 13642 -3115
rect 11920 -3229 11972 -3217
rect 13590 -3217 13598 -3183
rect 13632 -3217 13642 -3183
rect 13590 -3229 13642 -3217
rect 14588 -3081 14640 -3055
rect 14588 -3115 14598 -3081
rect 14632 -3115 14640 -3081
rect 14588 -3183 14640 -3115
rect 14588 -3217 14598 -3183
rect 14632 -3217 14640 -3183
rect 14786 -3081 14838 -3055
rect 14786 -3115 14794 -3081
rect 14828 -3115 14838 -3081
rect 14786 -3183 14838 -3115
rect 14588 -3229 14640 -3217
rect 14786 -3217 14794 -3183
rect 14828 -3217 14838 -3183
rect 14786 -3229 14838 -3217
rect 15784 -3081 15836 -3055
rect 15784 -3115 15794 -3081
rect 15828 -3115 15836 -3081
rect 15784 -3183 15836 -3115
rect 15784 -3217 15794 -3183
rect 15828 -3217 15836 -3183
rect 15982 -3081 16034 -3055
rect 15982 -3115 15990 -3081
rect 16024 -3115 16034 -3081
rect 15982 -3183 16034 -3115
rect 15784 -3229 15836 -3217
rect 15982 -3217 15990 -3183
rect 16024 -3217 16034 -3183
rect 15982 -3229 16034 -3217
rect 16612 -3081 16664 -3055
rect 16612 -3115 16622 -3081
rect 16656 -3115 16664 -3081
rect 16612 -3183 16664 -3115
rect 16612 -3217 16622 -3183
rect 16656 -3217 16664 -3183
rect 16612 -3229 16664 -3217
rect -2970 -3335 -2918 -3323
rect -2970 -3369 -2962 -3335
rect -2928 -3369 -2918 -3335
rect -2970 -3437 -2918 -3369
rect -2970 -3471 -2962 -3437
rect -2928 -3471 -2918 -3437
rect -2970 -3497 -2918 -3471
rect -2340 -3335 -2288 -3323
rect -2340 -3369 -2330 -3335
rect -2296 -3369 -2288 -3335
rect -1590 -3335 -1538 -3323
rect -2340 -3437 -2288 -3369
rect -2340 -3471 -2330 -3437
rect -2296 -3471 -2288 -3437
rect -2340 -3497 -2288 -3471
rect -1590 -3369 -1582 -3335
rect -1548 -3369 -1538 -3335
rect -1590 -3437 -1538 -3369
rect -1590 -3471 -1582 -3437
rect -1548 -3471 -1538 -3437
rect -1590 -3497 -1538 -3471
rect -960 -3335 -908 -3323
rect -960 -3369 -950 -3335
rect -916 -3369 -908 -3335
rect -960 -3437 -908 -3369
rect -960 -3471 -950 -3437
rect -916 -3471 -908 -3437
rect -960 -3497 -908 -3471
rect -854 -3335 -802 -3323
rect -854 -3369 -846 -3335
rect -812 -3369 -802 -3335
rect -854 -3437 -802 -3369
rect -854 -3471 -846 -3437
rect -812 -3471 -802 -3437
rect -854 -3497 -802 -3471
rect -224 -3335 -172 -3323
rect -224 -3369 -214 -3335
rect -180 -3369 -172 -3335
rect -26 -3335 26 -3323
rect -224 -3437 -172 -3369
rect -224 -3471 -214 -3437
rect -180 -3471 -172 -3437
rect -224 -3497 -172 -3471
rect -26 -3369 -18 -3335
rect 16 -3369 26 -3335
rect -26 -3437 26 -3369
rect -26 -3471 -18 -3437
rect 16 -3471 26 -3437
rect -26 -3497 26 -3471
rect 236 -3335 288 -3323
rect 236 -3369 246 -3335
rect 280 -3369 288 -3335
rect 236 -3437 288 -3369
rect 236 -3471 246 -3437
rect 280 -3471 288 -3437
rect 236 -3497 288 -3471
rect 434 -3343 505 -3323
rect 434 -3377 457 -3343
rect 491 -3377 505 -3343
rect 434 -3411 505 -3377
rect 434 -3445 457 -3411
rect 491 -3445 505 -3411
rect 434 -3523 505 -3445
rect 535 -3342 600 -3323
rect 535 -3376 555 -3342
rect 589 -3376 600 -3342
rect 535 -3410 600 -3376
rect 535 -3444 555 -3410
rect 589 -3444 600 -3410
rect 535 -3487 600 -3444
rect 700 -3343 753 -3323
rect 700 -3377 711 -3343
rect 745 -3377 753 -3343
rect 700 -3411 753 -3377
rect 700 -3445 711 -3411
rect 745 -3445 753 -3411
rect 700 -3487 753 -3445
rect 807 -3342 860 -3323
rect 807 -3376 815 -3342
rect 849 -3376 860 -3342
rect 807 -3410 860 -3376
rect 807 -3444 815 -3410
rect 849 -3444 860 -3410
rect 807 -3487 860 -3444
rect 960 -3342 1032 -3323
rect 960 -3376 973 -3342
rect 1007 -3376 1032 -3342
rect 960 -3410 1032 -3376
rect 960 -3444 973 -3410
rect 1007 -3444 1032 -3410
rect 960 -3487 1032 -3444
rect 535 -3523 585 -3487
rect 982 -3523 1032 -3487
rect 1062 -3342 1116 -3323
rect 1262 -3335 1314 -3323
rect 1062 -3376 1073 -3342
rect 1107 -3376 1116 -3342
rect 1062 -3410 1116 -3376
rect 1062 -3444 1073 -3410
rect 1107 -3444 1116 -3410
rect 1062 -3523 1116 -3444
rect 1262 -3369 1270 -3335
rect 1304 -3369 1314 -3335
rect 1262 -3437 1314 -3369
rect 1262 -3471 1270 -3437
rect 1304 -3471 1314 -3437
rect 1262 -3497 1314 -3471
rect 1524 -3335 1576 -3323
rect 1524 -3369 1534 -3335
rect 1568 -3369 1576 -3335
rect 1722 -3335 1774 -3323
rect 1524 -3437 1576 -3369
rect 1524 -3471 1534 -3437
rect 1568 -3471 1576 -3437
rect 1524 -3497 1576 -3471
rect 1722 -3369 1730 -3335
rect 1764 -3369 1774 -3335
rect 1722 -3437 1774 -3369
rect 1722 -3471 1730 -3437
rect 1764 -3471 1774 -3437
rect 1722 -3497 1774 -3471
rect 2352 -3335 2404 -3323
rect 2352 -3369 2362 -3335
rect 2396 -3369 2404 -3335
rect 2550 -3335 2602 -3323
rect 2352 -3437 2404 -3369
rect 2352 -3471 2362 -3437
rect 2396 -3471 2404 -3437
rect 2352 -3497 2404 -3471
rect 2550 -3369 2558 -3335
rect 2592 -3369 2602 -3335
rect 2550 -3437 2602 -3369
rect 2550 -3471 2558 -3437
rect 2592 -3471 2602 -3437
rect 2550 -3497 2602 -3471
rect 2812 -3335 2864 -3323
rect 2812 -3369 2822 -3335
rect 2856 -3369 2864 -3335
rect 2812 -3437 2864 -3369
rect 2812 -3471 2822 -3437
rect 2856 -3471 2864 -3437
rect 2812 -3497 2864 -3471
rect 3010 -3343 3081 -3323
rect 3010 -3377 3033 -3343
rect 3067 -3377 3081 -3343
rect 3010 -3411 3081 -3377
rect 3010 -3445 3033 -3411
rect 3067 -3445 3081 -3411
rect 3010 -3523 3081 -3445
rect 3111 -3342 3176 -3323
rect 3111 -3376 3131 -3342
rect 3165 -3376 3176 -3342
rect 3111 -3410 3176 -3376
rect 3111 -3444 3131 -3410
rect 3165 -3444 3176 -3410
rect 3111 -3487 3176 -3444
rect 3276 -3343 3329 -3323
rect 3276 -3377 3287 -3343
rect 3321 -3377 3329 -3343
rect 3276 -3411 3329 -3377
rect 3276 -3445 3287 -3411
rect 3321 -3445 3329 -3411
rect 3276 -3487 3329 -3445
rect 3383 -3342 3436 -3323
rect 3383 -3376 3391 -3342
rect 3425 -3376 3436 -3342
rect 3383 -3410 3436 -3376
rect 3383 -3444 3391 -3410
rect 3425 -3444 3436 -3410
rect 3383 -3487 3436 -3444
rect 3536 -3342 3608 -3323
rect 3536 -3376 3549 -3342
rect 3583 -3376 3608 -3342
rect 3536 -3410 3608 -3376
rect 3536 -3444 3549 -3410
rect 3583 -3444 3608 -3410
rect 3536 -3487 3608 -3444
rect 3111 -3523 3161 -3487
rect 3558 -3523 3608 -3487
rect 3638 -3342 3692 -3323
rect 3838 -3335 3890 -3323
rect 3638 -3376 3649 -3342
rect 3683 -3376 3692 -3342
rect 3638 -3410 3692 -3376
rect 3638 -3444 3649 -3410
rect 3683 -3444 3692 -3410
rect 3638 -3523 3692 -3444
rect 3838 -3369 3846 -3335
rect 3880 -3369 3890 -3335
rect 3838 -3437 3890 -3369
rect 3838 -3471 3846 -3437
rect 3880 -3471 3890 -3437
rect 3838 -3497 3890 -3471
rect 4100 -3335 4152 -3323
rect 4100 -3369 4110 -3335
rect 4144 -3369 4152 -3335
rect 4298 -3335 4350 -3323
rect 4100 -3437 4152 -3369
rect 4100 -3471 4110 -3437
rect 4144 -3471 4152 -3437
rect 4100 -3497 4152 -3471
rect 4298 -3369 4306 -3335
rect 4340 -3369 4350 -3335
rect 4298 -3437 4350 -3369
rect 4298 -3471 4306 -3437
rect 4340 -3471 4350 -3437
rect 4298 -3497 4350 -3471
rect 4928 -3335 4980 -3323
rect 4928 -3369 4938 -3335
rect 4972 -3369 4980 -3335
rect 5126 -3335 5178 -3323
rect 4928 -3437 4980 -3369
rect 4928 -3471 4938 -3437
rect 4972 -3471 4980 -3437
rect 4928 -3497 4980 -3471
rect 5126 -3369 5134 -3335
rect 5168 -3369 5178 -3335
rect 5126 -3437 5178 -3369
rect 5126 -3471 5134 -3437
rect 5168 -3471 5178 -3437
rect 5126 -3497 5178 -3471
rect 5388 -3335 5440 -3323
rect 5388 -3369 5398 -3335
rect 5432 -3369 5440 -3335
rect 5388 -3437 5440 -3369
rect 5388 -3471 5398 -3437
rect 5432 -3471 5440 -3437
rect 5388 -3497 5440 -3471
rect 5586 -3343 5657 -3323
rect 5586 -3377 5609 -3343
rect 5643 -3377 5657 -3343
rect 5586 -3411 5657 -3377
rect 5586 -3445 5609 -3411
rect 5643 -3445 5657 -3411
rect 5586 -3523 5657 -3445
rect 5687 -3342 5752 -3323
rect 5687 -3376 5707 -3342
rect 5741 -3376 5752 -3342
rect 5687 -3410 5752 -3376
rect 5687 -3444 5707 -3410
rect 5741 -3444 5752 -3410
rect 5687 -3487 5752 -3444
rect 5852 -3343 5905 -3323
rect 5852 -3377 5863 -3343
rect 5897 -3377 5905 -3343
rect 5852 -3411 5905 -3377
rect 5852 -3445 5863 -3411
rect 5897 -3445 5905 -3411
rect 5852 -3487 5905 -3445
rect 5959 -3342 6012 -3323
rect 5959 -3376 5967 -3342
rect 6001 -3376 6012 -3342
rect 5959 -3410 6012 -3376
rect 5959 -3444 5967 -3410
rect 6001 -3444 6012 -3410
rect 5959 -3487 6012 -3444
rect 6112 -3342 6184 -3323
rect 6112 -3376 6125 -3342
rect 6159 -3376 6184 -3342
rect 6112 -3410 6184 -3376
rect 6112 -3444 6125 -3410
rect 6159 -3444 6184 -3410
rect 6112 -3487 6184 -3444
rect 5687 -3523 5737 -3487
rect 6134 -3523 6184 -3487
rect 6214 -3342 6268 -3323
rect 6414 -3335 6466 -3323
rect 6214 -3376 6225 -3342
rect 6259 -3376 6268 -3342
rect 6214 -3410 6268 -3376
rect 6214 -3444 6225 -3410
rect 6259 -3444 6268 -3410
rect 6214 -3523 6268 -3444
rect 6414 -3369 6422 -3335
rect 6456 -3369 6466 -3335
rect 6414 -3437 6466 -3369
rect 6414 -3471 6422 -3437
rect 6456 -3471 6466 -3437
rect 6414 -3497 6466 -3471
rect 6676 -3335 6728 -3323
rect 6676 -3369 6686 -3335
rect 6720 -3369 6728 -3335
rect 6874 -3335 6926 -3323
rect 6676 -3437 6728 -3369
rect 6676 -3471 6686 -3437
rect 6720 -3471 6728 -3437
rect 6676 -3497 6728 -3471
rect 6874 -3369 6882 -3335
rect 6916 -3369 6926 -3335
rect 6874 -3437 6926 -3369
rect 6874 -3471 6882 -3437
rect 6916 -3471 6926 -3437
rect 6874 -3497 6926 -3471
rect 7504 -3335 7556 -3323
rect 7504 -3369 7514 -3335
rect 7548 -3369 7556 -3335
rect 7702 -3335 7754 -3323
rect 7504 -3437 7556 -3369
rect 7504 -3471 7514 -3437
rect 7548 -3471 7556 -3437
rect 7504 -3497 7556 -3471
rect 7702 -3369 7710 -3335
rect 7744 -3369 7754 -3335
rect 7702 -3437 7754 -3369
rect 7702 -3471 7710 -3437
rect 7744 -3471 7754 -3437
rect 7702 -3497 7754 -3471
rect 7964 -3335 8016 -3323
rect 7964 -3369 7974 -3335
rect 8008 -3369 8016 -3335
rect 7964 -3437 8016 -3369
rect 7964 -3471 7974 -3437
rect 8008 -3471 8016 -3437
rect 7964 -3497 8016 -3471
rect 8162 -3343 8233 -3323
rect 8162 -3377 8185 -3343
rect 8219 -3377 8233 -3343
rect 8162 -3411 8233 -3377
rect 8162 -3445 8185 -3411
rect 8219 -3445 8233 -3411
rect 8162 -3523 8233 -3445
rect 8263 -3342 8328 -3323
rect 8263 -3376 8283 -3342
rect 8317 -3376 8328 -3342
rect 8263 -3410 8328 -3376
rect 8263 -3444 8283 -3410
rect 8317 -3444 8328 -3410
rect 8263 -3487 8328 -3444
rect 8428 -3343 8481 -3323
rect 8428 -3377 8439 -3343
rect 8473 -3377 8481 -3343
rect 8428 -3411 8481 -3377
rect 8428 -3445 8439 -3411
rect 8473 -3445 8481 -3411
rect 8428 -3487 8481 -3445
rect 8535 -3342 8588 -3323
rect 8535 -3376 8543 -3342
rect 8577 -3376 8588 -3342
rect 8535 -3410 8588 -3376
rect 8535 -3444 8543 -3410
rect 8577 -3444 8588 -3410
rect 8535 -3487 8588 -3444
rect 8688 -3342 8760 -3323
rect 8688 -3376 8701 -3342
rect 8735 -3376 8760 -3342
rect 8688 -3410 8760 -3376
rect 8688 -3444 8701 -3410
rect 8735 -3444 8760 -3410
rect 8688 -3487 8760 -3444
rect 8263 -3523 8313 -3487
rect 8710 -3523 8760 -3487
rect 8790 -3342 8844 -3323
rect 8990 -3335 9042 -3323
rect 8790 -3376 8801 -3342
rect 8835 -3376 8844 -3342
rect 8790 -3410 8844 -3376
rect 8790 -3444 8801 -3410
rect 8835 -3444 8844 -3410
rect 8790 -3523 8844 -3444
rect 8990 -3369 8998 -3335
rect 9032 -3369 9042 -3335
rect 8990 -3437 9042 -3369
rect 8990 -3471 8998 -3437
rect 9032 -3471 9042 -3437
rect 8990 -3497 9042 -3471
rect 9252 -3335 9304 -3323
rect 9252 -3369 9262 -3335
rect 9296 -3369 9304 -3335
rect 9450 -3335 9502 -3323
rect 9252 -3437 9304 -3369
rect 9252 -3471 9262 -3437
rect 9296 -3471 9304 -3437
rect 9252 -3497 9304 -3471
rect 9450 -3369 9458 -3335
rect 9492 -3369 9502 -3335
rect 9450 -3437 9502 -3369
rect 9450 -3471 9458 -3437
rect 9492 -3471 9502 -3437
rect 9450 -3497 9502 -3471
rect 10080 -3335 10132 -3323
rect 10080 -3369 10090 -3335
rect 10124 -3369 10132 -3335
rect 10370 -3335 10422 -3323
rect 10080 -3437 10132 -3369
rect 10080 -3471 10090 -3437
rect 10124 -3471 10132 -3437
rect 10080 -3497 10132 -3471
rect 10370 -3369 10378 -3335
rect 10412 -3369 10422 -3335
rect 10370 -3437 10422 -3369
rect 10370 -3471 10378 -3437
rect 10412 -3471 10422 -3437
rect 10370 -3497 10422 -3471
rect 10632 -3335 10684 -3323
rect 10632 -3369 10642 -3335
rect 10676 -3369 10684 -3335
rect 10632 -3437 10684 -3369
rect 10632 -3471 10642 -3437
rect 10676 -3471 10684 -3437
rect 10632 -3497 10684 -3471
rect 10738 -3343 10809 -3323
rect 10738 -3377 10761 -3343
rect 10795 -3377 10809 -3343
rect 10738 -3411 10809 -3377
rect 10738 -3445 10761 -3411
rect 10795 -3445 10809 -3411
rect 10738 -3523 10809 -3445
rect 10839 -3342 10904 -3323
rect 10839 -3376 10859 -3342
rect 10893 -3376 10904 -3342
rect 10839 -3410 10904 -3376
rect 10839 -3444 10859 -3410
rect 10893 -3444 10904 -3410
rect 10839 -3487 10904 -3444
rect 11004 -3343 11057 -3323
rect 11004 -3377 11015 -3343
rect 11049 -3377 11057 -3343
rect 11004 -3411 11057 -3377
rect 11004 -3445 11015 -3411
rect 11049 -3445 11057 -3411
rect 11004 -3487 11057 -3445
rect 11111 -3342 11164 -3323
rect 11111 -3376 11119 -3342
rect 11153 -3376 11164 -3342
rect 11111 -3410 11164 -3376
rect 11111 -3444 11119 -3410
rect 11153 -3444 11164 -3410
rect 11111 -3487 11164 -3444
rect 11264 -3342 11336 -3323
rect 11264 -3376 11277 -3342
rect 11311 -3376 11336 -3342
rect 11264 -3410 11336 -3376
rect 11264 -3444 11277 -3410
rect 11311 -3444 11336 -3410
rect 11264 -3487 11336 -3444
rect 10839 -3523 10889 -3487
rect 11286 -3523 11336 -3487
rect 11366 -3342 11420 -3323
rect 11658 -3335 11710 -3323
rect 11366 -3376 11377 -3342
rect 11411 -3376 11420 -3342
rect 11366 -3410 11420 -3376
rect 11366 -3444 11377 -3410
rect 11411 -3444 11420 -3410
rect 11366 -3523 11420 -3444
rect 11658 -3369 11666 -3335
rect 11700 -3369 11710 -3335
rect 11658 -3437 11710 -3369
rect 11658 -3471 11666 -3437
rect 11700 -3471 11710 -3437
rect 11658 -3497 11710 -3471
rect 11920 -3335 11972 -3323
rect 11920 -3369 11930 -3335
rect 11964 -3369 11972 -3335
rect 13590 -3335 13642 -3323
rect 11920 -3437 11972 -3369
rect 11920 -3471 11930 -3437
rect 11964 -3471 11972 -3437
rect 11920 -3497 11972 -3471
rect 13590 -3369 13598 -3335
rect 13632 -3369 13642 -3335
rect 13590 -3437 13642 -3369
rect 13590 -3471 13598 -3437
rect 13632 -3471 13642 -3437
rect 13590 -3497 13642 -3471
rect 14588 -3335 14640 -3323
rect 14588 -3369 14598 -3335
rect 14632 -3369 14640 -3335
rect 14786 -3335 14838 -3323
rect 14588 -3437 14640 -3369
rect 14588 -3471 14598 -3437
rect 14632 -3471 14640 -3437
rect 14588 -3497 14640 -3471
rect 14786 -3369 14794 -3335
rect 14828 -3369 14838 -3335
rect 14786 -3437 14838 -3369
rect 14786 -3471 14794 -3437
rect 14828 -3471 14838 -3437
rect 14786 -3497 14838 -3471
rect 15784 -3335 15836 -3323
rect 15784 -3369 15794 -3335
rect 15828 -3369 15836 -3335
rect 15982 -3335 16034 -3323
rect 15784 -3437 15836 -3369
rect 15784 -3471 15794 -3437
rect 15828 -3471 15836 -3437
rect 15784 -3497 15836 -3471
rect 15982 -3369 15990 -3335
rect 16024 -3369 16034 -3335
rect 15982 -3437 16034 -3369
rect 15982 -3471 15990 -3437
rect 16024 -3471 16034 -3437
rect 15982 -3497 16034 -3471
rect 16612 -3335 16664 -3323
rect 16612 -3369 16622 -3335
rect 16656 -3369 16664 -3335
rect 16612 -3437 16664 -3369
rect 16612 -3471 16622 -3437
rect 16656 -3471 16664 -3437
rect 16612 -3497 16664 -3471
rect -2970 -4169 -2918 -4143
rect -2970 -4203 -2962 -4169
rect -2928 -4203 -2918 -4169
rect -2970 -4271 -2918 -4203
rect -2970 -4305 -2962 -4271
rect -2928 -4305 -2918 -4271
rect -2970 -4317 -2918 -4305
rect -2340 -4169 -2288 -4143
rect -2340 -4203 -2330 -4169
rect -2296 -4203 -2288 -4169
rect -2340 -4271 -2288 -4203
rect -2340 -4305 -2330 -4271
rect -2296 -4305 -2288 -4271
rect -1590 -4169 -1538 -4143
rect -1590 -4203 -1582 -4169
rect -1548 -4203 -1538 -4169
rect -1590 -4271 -1538 -4203
rect -2340 -4317 -2288 -4305
rect -1590 -4305 -1582 -4271
rect -1548 -4305 -1538 -4271
rect -1590 -4317 -1538 -4305
rect -960 -4169 -908 -4143
rect -960 -4203 -950 -4169
rect -916 -4203 -908 -4169
rect -960 -4271 -908 -4203
rect -960 -4305 -950 -4271
rect -916 -4305 -908 -4271
rect -960 -4317 -908 -4305
rect -854 -4169 -802 -4143
rect -854 -4203 -846 -4169
rect -812 -4203 -802 -4169
rect -854 -4271 -802 -4203
rect -854 -4305 -846 -4271
rect -812 -4305 -802 -4271
rect -854 -4317 -802 -4305
rect -224 -4169 -172 -4143
rect -224 -4203 -214 -4169
rect -180 -4203 -172 -4169
rect -224 -4271 -172 -4203
rect -224 -4305 -214 -4271
rect -180 -4305 -172 -4271
rect -26 -4169 26 -4143
rect -26 -4203 -18 -4169
rect 16 -4203 26 -4169
rect -26 -4271 26 -4203
rect -224 -4317 -172 -4305
rect -26 -4305 -18 -4271
rect 16 -4305 26 -4271
rect -26 -4317 26 -4305
rect 236 -4169 288 -4143
rect 236 -4203 246 -4169
rect 280 -4203 288 -4169
rect 236 -4271 288 -4203
rect 236 -4305 246 -4271
rect 280 -4305 288 -4271
rect 434 -4196 488 -4117
rect 434 -4230 443 -4196
rect 477 -4230 488 -4196
rect 434 -4264 488 -4230
rect 434 -4298 443 -4264
rect 477 -4298 488 -4264
rect 236 -4317 288 -4305
rect 434 -4317 488 -4298
rect 518 -4153 568 -4117
rect 965 -4153 1015 -4117
rect 518 -4196 590 -4153
rect 518 -4230 543 -4196
rect 577 -4230 590 -4196
rect 518 -4264 590 -4230
rect 518 -4298 543 -4264
rect 577 -4298 590 -4264
rect 518 -4317 590 -4298
rect 690 -4196 743 -4153
rect 690 -4230 701 -4196
rect 735 -4230 743 -4196
rect 690 -4264 743 -4230
rect 690 -4298 701 -4264
rect 735 -4298 743 -4264
rect 690 -4317 743 -4298
rect 797 -4195 850 -4153
rect 797 -4229 805 -4195
rect 839 -4229 850 -4195
rect 797 -4263 850 -4229
rect 797 -4297 805 -4263
rect 839 -4297 850 -4263
rect 797 -4317 850 -4297
rect 950 -4196 1015 -4153
rect 950 -4230 961 -4196
rect 995 -4230 1015 -4196
rect 950 -4264 1015 -4230
rect 950 -4298 961 -4264
rect 995 -4298 1015 -4264
rect 950 -4317 1015 -4298
rect 1045 -4195 1116 -4117
rect 1045 -4229 1059 -4195
rect 1093 -4229 1116 -4195
rect 1045 -4263 1116 -4229
rect 1045 -4297 1059 -4263
rect 1093 -4297 1116 -4263
rect 1045 -4317 1116 -4297
rect 1262 -4169 1314 -4143
rect 1262 -4203 1270 -4169
rect 1304 -4203 1314 -4169
rect 1262 -4271 1314 -4203
rect 1262 -4305 1270 -4271
rect 1304 -4305 1314 -4271
rect 1262 -4317 1314 -4305
rect 1524 -4169 1576 -4143
rect 1524 -4203 1534 -4169
rect 1568 -4203 1576 -4169
rect 1524 -4271 1576 -4203
rect 1524 -4305 1534 -4271
rect 1568 -4305 1576 -4271
rect 1722 -4169 1774 -4143
rect 1722 -4203 1730 -4169
rect 1764 -4203 1774 -4169
rect 1722 -4271 1774 -4203
rect 1524 -4317 1576 -4305
rect 1722 -4305 1730 -4271
rect 1764 -4305 1774 -4271
rect 1722 -4317 1774 -4305
rect 2352 -4169 2404 -4143
rect 2352 -4203 2362 -4169
rect 2396 -4203 2404 -4169
rect 2352 -4271 2404 -4203
rect 2352 -4305 2362 -4271
rect 2396 -4305 2404 -4271
rect 2550 -4169 2602 -4143
rect 2550 -4203 2558 -4169
rect 2592 -4203 2602 -4169
rect 2550 -4271 2602 -4203
rect 2352 -4317 2404 -4305
rect 2550 -4305 2558 -4271
rect 2592 -4305 2602 -4271
rect 2550 -4317 2602 -4305
rect 2812 -4169 2864 -4143
rect 2812 -4203 2822 -4169
rect 2856 -4203 2864 -4169
rect 2812 -4271 2864 -4203
rect 2812 -4305 2822 -4271
rect 2856 -4305 2864 -4271
rect 3010 -4196 3064 -4117
rect 3010 -4230 3019 -4196
rect 3053 -4230 3064 -4196
rect 3010 -4264 3064 -4230
rect 3010 -4298 3019 -4264
rect 3053 -4298 3064 -4264
rect 2812 -4317 2864 -4305
rect 3010 -4317 3064 -4298
rect 3094 -4153 3144 -4117
rect 3541 -4153 3591 -4117
rect 3094 -4196 3166 -4153
rect 3094 -4230 3119 -4196
rect 3153 -4230 3166 -4196
rect 3094 -4264 3166 -4230
rect 3094 -4298 3119 -4264
rect 3153 -4298 3166 -4264
rect 3094 -4317 3166 -4298
rect 3266 -4196 3319 -4153
rect 3266 -4230 3277 -4196
rect 3311 -4230 3319 -4196
rect 3266 -4264 3319 -4230
rect 3266 -4298 3277 -4264
rect 3311 -4298 3319 -4264
rect 3266 -4317 3319 -4298
rect 3373 -4195 3426 -4153
rect 3373 -4229 3381 -4195
rect 3415 -4229 3426 -4195
rect 3373 -4263 3426 -4229
rect 3373 -4297 3381 -4263
rect 3415 -4297 3426 -4263
rect 3373 -4317 3426 -4297
rect 3526 -4196 3591 -4153
rect 3526 -4230 3537 -4196
rect 3571 -4230 3591 -4196
rect 3526 -4264 3591 -4230
rect 3526 -4298 3537 -4264
rect 3571 -4298 3591 -4264
rect 3526 -4317 3591 -4298
rect 3621 -4195 3692 -4117
rect 3621 -4229 3635 -4195
rect 3669 -4229 3692 -4195
rect 3621 -4263 3692 -4229
rect 3621 -4297 3635 -4263
rect 3669 -4297 3692 -4263
rect 3621 -4317 3692 -4297
rect 3838 -4169 3890 -4143
rect 3838 -4203 3846 -4169
rect 3880 -4203 3890 -4169
rect 3838 -4271 3890 -4203
rect 3838 -4305 3846 -4271
rect 3880 -4305 3890 -4271
rect 3838 -4317 3890 -4305
rect 4100 -4169 4152 -4143
rect 4100 -4203 4110 -4169
rect 4144 -4203 4152 -4169
rect 4100 -4271 4152 -4203
rect 4100 -4305 4110 -4271
rect 4144 -4305 4152 -4271
rect 4298 -4169 4350 -4143
rect 4298 -4203 4306 -4169
rect 4340 -4203 4350 -4169
rect 4298 -4271 4350 -4203
rect 4100 -4317 4152 -4305
rect 4298 -4305 4306 -4271
rect 4340 -4305 4350 -4271
rect 4298 -4317 4350 -4305
rect 4928 -4169 4980 -4143
rect 4928 -4203 4938 -4169
rect 4972 -4203 4980 -4169
rect 4928 -4271 4980 -4203
rect 4928 -4305 4938 -4271
rect 4972 -4305 4980 -4271
rect 5126 -4169 5178 -4143
rect 5126 -4203 5134 -4169
rect 5168 -4203 5178 -4169
rect 5126 -4271 5178 -4203
rect 4928 -4317 4980 -4305
rect 5126 -4305 5134 -4271
rect 5168 -4305 5178 -4271
rect 5126 -4317 5178 -4305
rect 5388 -4169 5440 -4143
rect 5388 -4203 5398 -4169
rect 5432 -4203 5440 -4169
rect 5388 -4271 5440 -4203
rect 5388 -4305 5398 -4271
rect 5432 -4305 5440 -4271
rect 5586 -4196 5640 -4117
rect 5586 -4230 5595 -4196
rect 5629 -4230 5640 -4196
rect 5586 -4264 5640 -4230
rect 5586 -4298 5595 -4264
rect 5629 -4298 5640 -4264
rect 5388 -4317 5440 -4305
rect 5586 -4317 5640 -4298
rect 5670 -4153 5720 -4117
rect 6117 -4153 6167 -4117
rect 5670 -4196 5742 -4153
rect 5670 -4230 5695 -4196
rect 5729 -4230 5742 -4196
rect 5670 -4264 5742 -4230
rect 5670 -4298 5695 -4264
rect 5729 -4298 5742 -4264
rect 5670 -4317 5742 -4298
rect 5842 -4196 5895 -4153
rect 5842 -4230 5853 -4196
rect 5887 -4230 5895 -4196
rect 5842 -4264 5895 -4230
rect 5842 -4298 5853 -4264
rect 5887 -4298 5895 -4264
rect 5842 -4317 5895 -4298
rect 5949 -4195 6002 -4153
rect 5949 -4229 5957 -4195
rect 5991 -4229 6002 -4195
rect 5949 -4263 6002 -4229
rect 5949 -4297 5957 -4263
rect 5991 -4297 6002 -4263
rect 5949 -4317 6002 -4297
rect 6102 -4196 6167 -4153
rect 6102 -4230 6113 -4196
rect 6147 -4230 6167 -4196
rect 6102 -4264 6167 -4230
rect 6102 -4298 6113 -4264
rect 6147 -4298 6167 -4264
rect 6102 -4317 6167 -4298
rect 6197 -4195 6268 -4117
rect 6197 -4229 6211 -4195
rect 6245 -4229 6268 -4195
rect 6197 -4263 6268 -4229
rect 6197 -4297 6211 -4263
rect 6245 -4297 6268 -4263
rect 6197 -4317 6268 -4297
rect 6414 -4169 6466 -4143
rect 6414 -4203 6422 -4169
rect 6456 -4203 6466 -4169
rect 6414 -4271 6466 -4203
rect 6414 -4305 6422 -4271
rect 6456 -4305 6466 -4271
rect 6414 -4317 6466 -4305
rect 6676 -4169 6728 -4143
rect 6676 -4203 6686 -4169
rect 6720 -4203 6728 -4169
rect 6676 -4271 6728 -4203
rect 6676 -4305 6686 -4271
rect 6720 -4305 6728 -4271
rect 6874 -4169 6926 -4143
rect 6874 -4203 6882 -4169
rect 6916 -4203 6926 -4169
rect 6874 -4271 6926 -4203
rect 6676 -4317 6728 -4305
rect 6874 -4305 6882 -4271
rect 6916 -4305 6926 -4271
rect 6874 -4317 6926 -4305
rect 7504 -4169 7556 -4143
rect 7504 -4203 7514 -4169
rect 7548 -4203 7556 -4169
rect 7504 -4271 7556 -4203
rect 7504 -4305 7514 -4271
rect 7548 -4305 7556 -4271
rect 7702 -4169 7754 -4143
rect 7702 -4203 7710 -4169
rect 7744 -4203 7754 -4169
rect 7702 -4271 7754 -4203
rect 7504 -4317 7556 -4305
rect 7702 -4305 7710 -4271
rect 7744 -4305 7754 -4271
rect 7702 -4317 7754 -4305
rect 7964 -4169 8016 -4143
rect 7964 -4203 7974 -4169
rect 8008 -4203 8016 -4169
rect 7964 -4271 8016 -4203
rect 7964 -4305 7974 -4271
rect 8008 -4305 8016 -4271
rect 8162 -4196 8216 -4117
rect 8162 -4230 8171 -4196
rect 8205 -4230 8216 -4196
rect 8162 -4264 8216 -4230
rect 8162 -4298 8171 -4264
rect 8205 -4298 8216 -4264
rect 7964 -4317 8016 -4305
rect 8162 -4317 8216 -4298
rect 8246 -4153 8296 -4117
rect 8693 -4153 8743 -4117
rect 8246 -4196 8318 -4153
rect 8246 -4230 8271 -4196
rect 8305 -4230 8318 -4196
rect 8246 -4264 8318 -4230
rect 8246 -4298 8271 -4264
rect 8305 -4298 8318 -4264
rect 8246 -4317 8318 -4298
rect 8418 -4196 8471 -4153
rect 8418 -4230 8429 -4196
rect 8463 -4230 8471 -4196
rect 8418 -4264 8471 -4230
rect 8418 -4298 8429 -4264
rect 8463 -4298 8471 -4264
rect 8418 -4317 8471 -4298
rect 8525 -4195 8578 -4153
rect 8525 -4229 8533 -4195
rect 8567 -4229 8578 -4195
rect 8525 -4263 8578 -4229
rect 8525 -4297 8533 -4263
rect 8567 -4297 8578 -4263
rect 8525 -4317 8578 -4297
rect 8678 -4196 8743 -4153
rect 8678 -4230 8689 -4196
rect 8723 -4230 8743 -4196
rect 8678 -4264 8743 -4230
rect 8678 -4298 8689 -4264
rect 8723 -4298 8743 -4264
rect 8678 -4317 8743 -4298
rect 8773 -4195 8844 -4117
rect 8773 -4229 8787 -4195
rect 8821 -4229 8844 -4195
rect 8773 -4263 8844 -4229
rect 8773 -4297 8787 -4263
rect 8821 -4297 8844 -4263
rect 8773 -4317 8844 -4297
rect 8990 -4169 9042 -4143
rect 8990 -4203 8998 -4169
rect 9032 -4203 9042 -4169
rect 8990 -4271 9042 -4203
rect 8990 -4305 8998 -4271
rect 9032 -4305 9042 -4271
rect 8990 -4317 9042 -4305
rect 9252 -4169 9304 -4143
rect 9252 -4203 9262 -4169
rect 9296 -4203 9304 -4169
rect 9252 -4271 9304 -4203
rect 9252 -4305 9262 -4271
rect 9296 -4305 9304 -4271
rect 9450 -4169 9502 -4143
rect 9450 -4203 9458 -4169
rect 9492 -4203 9502 -4169
rect 9450 -4271 9502 -4203
rect 9252 -4317 9304 -4305
rect 9450 -4305 9458 -4271
rect 9492 -4305 9502 -4271
rect 9450 -4317 9502 -4305
rect 10080 -4169 10132 -4143
rect 10080 -4203 10090 -4169
rect 10124 -4203 10132 -4169
rect 10080 -4271 10132 -4203
rect 10080 -4305 10090 -4271
rect 10124 -4305 10132 -4271
rect 10370 -4169 10422 -4143
rect 10370 -4203 10378 -4169
rect 10412 -4203 10422 -4169
rect 10370 -4271 10422 -4203
rect 10080 -4317 10132 -4305
rect 10370 -4305 10378 -4271
rect 10412 -4305 10422 -4271
rect 10370 -4317 10422 -4305
rect 10632 -4169 10684 -4143
rect 10632 -4203 10642 -4169
rect 10676 -4203 10684 -4169
rect 10632 -4271 10684 -4203
rect 10632 -4305 10642 -4271
rect 10676 -4305 10684 -4271
rect 10632 -4317 10684 -4305
rect 10738 -4196 10792 -4117
rect 10738 -4230 10747 -4196
rect 10781 -4230 10792 -4196
rect 10738 -4264 10792 -4230
rect 10738 -4298 10747 -4264
rect 10781 -4298 10792 -4264
rect 10738 -4317 10792 -4298
rect 10822 -4153 10872 -4117
rect 11269 -4153 11319 -4117
rect 10822 -4196 10894 -4153
rect 10822 -4230 10847 -4196
rect 10881 -4230 10894 -4196
rect 10822 -4264 10894 -4230
rect 10822 -4298 10847 -4264
rect 10881 -4298 10894 -4264
rect 10822 -4317 10894 -4298
rect 10994 -4196 11047 -4153
rect 10994 -4230 11005 -4196
rect 11039 -4230 11047 -4196
rect 10994 -4264 11047 -4230
rect 10994 -4298 11005 -4264
rect 11039 -4298 11047 -4264
rect 10994 -4317 11047 -4298
rect 11101 -4195 11154 -4153
rect 11101 -4229 11109 -4195
rect 11143 -4229 11154 -4195
rect 11101 -4263 11154 -4229
rect 11101 -4297 11109 -4263
rect 11143 -4297 11154 -4263
rect 11101 -4317 11154 -4297
rect 11254 -4196 11319 -4153
rect 11254 -4230 11265 -4196
rect 11299 -4230 11319 -4196
rect 11254 -4264 11319 -4230
rect 11254 -4298 11265 -4264
rect 11299 -4298 11319 -4264
rect 11254 -4317 11319 -4298
rect 11349 -4195 11420 -4117
rect 11349 -4229 11363 -4195
rect 11397 -4229 11420 -4195
rect 11349 -4263 11420 -4229
rect 11349 -4297 11363 -4263
rect 11397 -4297 11420 -4263
rect 11349 -4317 11420 -4297
rect 11658 -4169 11710 -4143
rect 11658 -4203 11666 -4169
rect 11700 -4203 11710 -4169
rect 11658 -4271 11710 -4203
rect 11658 -4305 11666 -4271
rect 11700 -4305 11710 -4271
rect 11658 -4317 11710 -4305
rect 11920 -4169 11972 -4143
rect 11920 -4203 11930 -4169
rect 11964 -4203 11972 -4169
rect 11920 -4271 11972 -4203
rect 11920 -4305 11930 -4271
rect 11964 -4305 11972 -4271
rect 12486 -4196 12547 -4117
rect 12486 -4230 12502 -4196
rect 12536 -4230 12547 -4196
rect 12486 -4264 12547 -4230
rect 12486 -4298 12502 -4264
rect 12536 -4298 12547 -4264
rect 11920 -4317 11972 -4305
rect 12486 -4317 12547 -4298
rect 12577 -4169 12633 -4117
rect 12577 -4203 12588 -4169
rect 12622 -4203 12633 -4169
rect 12577 -4257 12633 -4203
rect 12577 -4291 12588 -4257
rect 12622 -4291 12633 -4257
rect 12577 -4317 12633 -4291
rect 12663 -4196 12719 -4117
rect 12663 -4230 12674 -4196
rect 12708 -4230 12719 -4196
rect 12663 -4264 12719 -4230
rect 12663 -4298 12674 -4264
rect 12708 -4298 12719 -4264
rect 12663 -4317 12719 -4298
rect 12749 -4169 12805 -4117
rect 12749 -4203 12760 -4169
rect 12794 -4203 12805 -4169
rect 12749 -4257 12805 -4203
rect 12749 -4291 12760 -4257
rect 12794 -4291 12805 -4257
rect 12749 -4317 12805 -4291
rect 12835 -4196 12891 -4117
rect 12835 -4230 12846 -4196
rect 12880 -4230 12891 -4196
rect 12835 -4264 12891 -4230
rect 12835 -4298 12846 -4264
rect 12880 -4298 12891 -4264
rect 12835 -4317 12891 -4298
rect 12921 -4169 12977 -4117
rect 12921 -4203 12932 -4169
rect 12966 -4203 12977 -4169
rect 12921 -4257 12977 -4203
rect 12921 -4291 12932 -4257
rect 12966 -4291 12977 -4257
rect 12921 -4317 12977 -4291
rect 13007 -4196 13076 -4117
rect 13007 -4230 13018 -4196
rect 13052 -4230 13076 -4196
rect 13007 -4264 13076 -4230
rect 13007 -4298 13018 -4264
rect 13052 -4298 13076 -4264
rect 13007 -4317 13076 -4298
rect 13222 -4169 13274 -4143
rect 13222 -4203 13230 -4169
rect 13264 -4203 13274 -4169
rect 13222 -4271 13274 -4203
rect 13222 -4305 13230 -4271
rect 13264 -4305 13274 -4271
rect 13222 -4317 13274 -4305
rect 13484 -4169 13536 -4143
rect 13484 -4203 13494 -4169
rect 13528 -4203 13536 -4169
rect 13484 -4271 13536 -4203
rect 13484 -4305 13494 -4271
rect 13528 -4305 13536 -4271
rect 13682 -4203 13735 -4117
rect 13682 -4237 13690 -4203
rect 13724 -4237 13735 -4203
rect 13682 -4271 13735 -4237
rect 13484 -4317 13536 -4305
rect 13682 -4305 13690 -4271
rect 13724 -4305 13735 -4271
rect 13682 -4317 13735 -4305
rect 13765 -4195 13821 -4117
rect 13765 -4229 13776 -4195
rect 13810 -4229 13821 -4195
rect 13765 -4263 13821 -4229
rect 13765 -4297 13776 -4263
rect 13810 -4297 13821 -4263
rect 13765 -4317 13821 -4297
rect 13851 -4203 13907 -4117
rect 13851 -4237 13862 -4203
rect 13896 -4237 13907 -4203
rect 13851 -4271 13907 -4237
rect 13851 -4305 13862 -4271
rect 13896 -4305 13907 -4271
rect 13851 -4317 13907 -4305
rect 13937 -4187 13993 -4117
rect 13937 -4221 13948 -4187
rect 13982 -4221 13993 -4187
rect 13937 -4255 13993 -4221
rect 13937 -4289 13948 -4255
rect 13982 -4289 13993 -4255
rect 13937 -4317 13993 -4289
rect 14023 -4203 14079 -4117
rect 14023 -4237 14034 -4203
rect 14068 -4237 14079 -4203
rect 14023 -4271 14079 -4237
rect 14023 -4305 14034 -4271
rect 14068 -4305 14079 -4271
rect 14023 -4317 14079 -4305
rect 14109 -4141 14165 -4117
rect 14109 -4175 14120 -4141
rect 14154 -4175 14165 -4141
rect 14109 -4227 14165 -4175
rect 14109 -4261 14120 -4227
rect 14154 -4261 14165 -4227
rect 14109 -4317 14165 -4261
rect 14195 -4247 14251 -4117
rect 14195 -4281 14206 -4247
rect 14240 -4281 14251 -4247
rect 14195 -4317 14251 -4281
rect 14281 -4141 14337 -4117
rect 14281 -4175 14292 -4141
rect 14326 -4175 14337 -4141
rect 14281 -4227 14337 -4175
rect 14281 -4261 14292 -4227
rect 14326 -4261 14337 -4227
rect 14281 -4317 14337 -4261
rect 14367 -4247 14423 -4117
rect 14367 -4281 14378 -4247
rect 14412 -4281 14423 -4247
rect 14367 -4317 14423 -4281
rect 14453 -4141 14509 -4117
rect 14453 -4175 14464 -4141
rect 14498 -4175 14509 -4141
rect 14453 -4227 14509 -4175
rect 14453 -4261 14464 -4227
rect 14498 -4261 14509 -4227
rect 14453 -4317 14509 -4261
rect 14539 -4247 14595 -4117
rect 14539 -4281 14550 -4247
rect 14584 -4281 14595 -4247
rect 14539 -4317 14595 -4281
rect 14625 -4141 14681 -4117
rect 14625 -4175 14636 -4141
rect 14670 -4175 14681 -4141
rect 14625 -4227 14681 -4175
rect 14625 -4261 14636 -4227
rect 14670 -4261 14681 -4227
rect 14625 -4317 14681 -4261
rect 14711 -4247 14766 -4117
rect 14711 -4281 14722 -4247
rect 14756 -4281 14766 -4247
rect 14711 -4317 14766 -4281
rect 14796 -4141 14852 -4117
rect 14796 -4175 14807 -4141
rect 14841 -4175 14852 -4141
rect 14796 -4227 14852 -4175
rect 14796 -4261 14807 -4227
rect 14841 -4261 14852 -4227
rect 14796 -4317 14852 -4261
rect 14882 -4247 14938 -4117
rect 14882 -4281 14893 -4247
rect 14927 -4281 14938 -4247
rect 14882 -4317 14938 -4281
rect 14968 -4141 15024 -4117
rect 14968 -4175 14979 -4141
rect 15013 -4175 15024 -4141
rect 14968 -4227 15024 -4175
rect 14968 -4261 14979 -4227
rect 15013 -4261 15024 -4227
rect 14968 -4317 15024 -4261
rect 15054 -4247 15110 -4117
rect 15054 -4281 15065 -4247
rect 15099 -4281 15110 -4247
rect 15054 -4317 15110 -4281
rect 15140 -4141 15196 -4117
rect 15140 -4175 15151 -4141
rect 15185 -4175 15196 -4141
rect 15140 -4227 15196 -4175
rect 15140 -4261 15151 -4227
rect 15185 -4261 15196 -4227
rect 15140 -4317 15196 -4261
rect 15226 -4247 15282 -4117
rect 15226 -4281 15237 -4247
rect 15271 -4281 15282 -4247
rect 15226 -4317 15282 -4281
rect 15312 -4141 15368 -4117
rect 15312 -4175 15323 -4141
rect 15357 -4175 15368 -4141
rect 15312 -4227 15368 -4175
rect 15312 -4261 15323 -4227
rect 15357 -4261 15368 -4227
rect 15312 -4317 15368 -4261
rect 15398 -4247 15451 -4117
rect 15398 -4281 15409 -4247
rect 15443 -4281 15451 -4247
rect 15398 -4317 15451 -4281
rect 15614 -4169 15666 -4143
rect 15614 -4203 15622 -4169
rect 15656 -4203 15666 -4169
rect 15614 -4271 15666 -4203
rect 15614 -4305 15622 -4271
rect 15656 -4305 15666 -4271
rect 15614 -4317 15666 -4305
rect 16612 -4169 16664 -4143
rect 16612 -4203 16622 -4169
rect 16656 -4203 16664 -4169
rect 16612 -4271 16664 -4203
rect 16612 -4305 16622 -4271
rect 16656 -4305 16664 -4271
rect 16612 -4317 16664 -4305
rect -2970 -4423 -2918 -4411
rect -2970 -4457 -2962 -4423
rect -2928 -4457 -2918 -4423
rect -2970 -4525 -2918 -4457
rect -2970 -4559 -2962 -4525
rect -2928 -4559 -2918 -4525
rect -2970 -4585 -2918 -4559
rect -2340 -4423 -2288 -4411
rect -2340 -4457 -2330 -4423
rect -2296 -4457 -2288 -4423
rect -1590 -4423 -1538 -4411
rect -2340 -4525 -2288 -4457
rect -2340 -4559 -2330 -4525
rect -2296 -4559 -2288 -4525
rect -2340 -4585 -2288 -4559
rect -1590 -4457 -1582 -4423
rect -1548 -4457 -1538 -4423
rect -1590 -4525 -1538 -4457
rect -1590 -4559 -1582 -4525
rect -1548 -4559 -1538 -4525
rect -1590 -4585 -1538 -4559
rect -960 -4423 -908 -4411
rect -960 -4457 -950 -4423
rect -916 -4457 -908 -4423
rect -960 -4525 -908 -4457
rect -960 -4559 -950 -4525
rect -916 -4559 -908 -4525
rect -960 -4585 -908 -4559
rect -854 -4431 -783 -4411
rect -854 -4465 -831 -4431
rect -797 -4465 -783 -4431
rect -854 -4499 -783 -4465
rect -854 -4533 -831 -4499
rect -797 -4533 -783 -4499
rect -854 -4611 -783 -4533
rect -753 -4430 -688 -4411
rect -753 -4464 -733 -4430
rect -699 -4464 -688 -4430
rect -753 -4498 -688 -4464
rect -753 -4532 -733 -4498
rect -699 -4532 -688 -4498
rect -753 -4575 -688 -4532
rect -588 -4431 -535 -4411
rect -588 -4465 -577 -4431
rect -543 -4465 -535 -4431
rect -588 -4499 -535 -4465
rect -588 -4533 -577 -4499
rect -543 -4533 -535 -4499
rect -588 -4575 -535 -4533
rect -481 -4430 -428 -4411
rect -481 -4464 -473 -4430
rect -439 -4464 -428 -4430
rect -481 -4498 -428 -4464
rect -481 -4532 -473 -4498
rect -439 -4532 -428 -4498
rect -481 -4575 -428 -4532
rect -328 -4430 -256 -4411
rect -328 -4464 -315 -4430
rect -281 -4464 -256 -4430
rect -328 -4498 -256 -4464
rect -328 -4532 -315 -4498
rect -281 -4532 -256 -4498
rect -328 -4575 -256 -4532
rect -753 -4611 -703 -4575
rect -306 -4611 -256 -4575
rect -226 -4430 -172 -4411
rect -26 -4423 26 -4411
rect -226 -4464 -215 -4430
rect -181 -4464 -172 -4430
rect -226 -4498 -172 -4464
rect -226 -4532 -215 -4498
rect -181 -4532 -172 -4498
rect -226 -4611 -172 -4532
rect -26 -4457 -18 -4423
rect 16 -4457 26 -4423
rect -26 -4525 26 -4457
rect -26 -4559 -18 -4525
rect 16 -4559 26 -4525
rect -26 -4585 26 -4559
rect 236 -4423 288 -4411
rect 236 -4457 246 -4423
rect 280 -4457 288 -4423
rect 236 -4525 288 -4457
rect 236 -4559 246 -4525
rect 280 -4559 288 -4525
rect 236 -4585 288 -4559
rect 434 -4431 505 -4411
rect 434 -4465 457 -4431
rect 491 -4465 505 -4431
rect 434 -4499 505 -4465
rect 434 -4533 457 -4499
rect 491 -4533 505 -4499
rect 434 -4611 505 -4533
rect 535 -4430 600 -4411
rect 535 -4464 555 -4430
rect 589 -4464 600 -4430
rect 535 -4498 600 -4464
rect 535 -4532 555 -4498
rect 589 -4532 600 -4498
rect 535 -4575 600 -4532
rect 700 -4431 753 -4411
rect 700 -4465 711 -4431
rect 745 -4465 753 -4431
rect 700 -4499 753 -4465
rect 700 -4533 711 -4499
rect 745 -4533 753 -4499
rect 700 -4575 753 -4533
rect 807 -4430 860 -4411
rect 807 -4464 815 -4430
rect 849 -4464 860 -4430
rect 807 -4498 860 -4464
rect 807 -4532 815 -4498
rect 849 -4532 860 -4498
rect 807 -4575 860 -4532
rect 960 -4430 1032 -4411
rect 960 -4464 973 -4430
rect 1007 -4464 1032 -4430
rect 960 -4498 1032 -4464
rect 960 -4532 973 -4498
rect 1007 -4532 1032 -4498
rect 960 -4575 1032 -4532
rect 535 -4611 585 -4575
rect 982 -4611 1032 -4575
rect 1062 -4430 1116 -4411
rect 1262 -4423 1314 -4411
rect 1062 -4464 1073 -4430
rect 1107 -4464 1116 -4430
rect 1062 -4498 1116 -4464
rect 1062 -4532 1073 -4498
rect 1107 -4532 1116 -4498
rect 1062 -4611 1116 -4532
rect 1262 -4457 1270 -4423
rect 1304 -4457 1314 -4423
rect 1262 -4525 1314 -4457
rect 1262 -4559 1270 -4525
rect 1304 -4559 1314 -4525
rect 1262 -4585 1314 -4559
rect 1524 -4423 1576 -4411
rect 1524 -4457 1534 -4423
rect 1568 -4457 1576 -4423
rect 1722 -4423 1774 -4411
rect 1524 -4525 1576 -4457
rect 1524 -4559 1534 -4525
rect 1568 -4559 1576 -4525
rect 1524 -4585 1576 -4559
rect 1722 -4457 1730 -4423
rect 1764 -4457 1774 -4423
rect 1722 -4525 1774 -4457
rect 1722 -4559 1730 -4525
rect 1764 -4559 1774 -4525
rect 1722 -4585 1774 -4559
rect 2352 -4423 2404 -4411
rect 2352 -4457 2362 -4423
rect 2396 -4457 2404 -4423
rect 2550 -4423 2602 -4411
rect 2352 -4525 2404 -4457
rect 2352 -4559 2362 -4525
rect 2396 -4559 2404 -4525
rect 2352 -4585 2404 -4559
rect 2550 -4457 2558 -4423
rect 2592 -4457 2602 -4423
rect 2550 -4525 2602 -4457
rect 2550 -4559 2558 -4525
rect 2592 -4559 2602 -4525
rect 2550 -4585 2602 -4559
rect 2812 -4423 2864 -4411
rect 2812 -4457 2822 -4423
rect 2856 -4457 2864 -4423
rect 2812 -4525 2864 -4457
rect 2812 -4559 2822 -4525
rect 2856 -4559 2864 -4525
rect 2812 -4585 2864 -4559
rect 3010 -4431 3081 -4411
rect 3010 -4465 3033 -4431
rect 3067 -4465 3081 -4431
rect 3010 -4499 3081 -4465
rect 3010 -4533 3033 -4499
rect 3067 -4533 3081 -4499
rect 3010 -4611 3081 -4533
rect 3111 -4430 3176 -4411
rect 3111 -4464 3131 -4430
rect 3165 -4464 3176 -4430
rect 3111 -4498 3176 -4464
rect 3111 -4532 3131 -4498
rect 3165 -4532 3176 -4498
rect 3111 -4575 3176 -4532
rect 3276 -4431 3329 -4411
rect 3276 -4465 3287 -4431
rect 3321 -4465 3329 -4431
rect 3276 -4499 3329 -4465
rect 3276 -4533 3287 -4499
rect 3321 -4533 3329 -4499
rect 3276 -4575 3329 -4533
rect 3383 -4430 3436 -4411
rect 3383 -4464 3391 -4430
rect 3425 -4464 3436 -4430
rect 3383 -4498 3436 -4464
rect 3383 -4532 3391 -4498
rect 3425 -4532 3436 -4498
rect 3383 -4575 3436 -4532
rect 3536 -4430 3608 -4411
rect 3536 -4464 3549 -4430
rect 3583 -4464 3608 -4430
rect 3536 -4498 3608 -4464
rect 3536 -4532 3549 -4498
rect 3583 -4532 3608 -4498
rect 3536 -4575 3608 -4532
rect 3111 -4611 3161 -4575
rect 3558 -4611 3608 -4575
rect 3638 -4430 3692 -4411
rect 3838 -4423 3890 -4411
rect 3638 -4464 3649 -4430
rect 3683 -4464 3692 -4430
rect 3638 -4498 3692 -4464
rect 3638 -4532 3649 -4498
rect 3683 -4532 3692 -4498
rect 3638 -4611 3692 -4532
rect 3838 -4457 3846 -4423
rect 3880 -4457 3890 -4423
rect 3838 -4525 3890 -4457
rect 3838 -4559 3846 -4525
rect 3880 -4559 3890 -4525
rect 3838 -4585 3890 -4559
rect 4100 -4423 4152 -4411
rect 4100 -4457 4110 -4423
rect 4144 -4457 4152 -4423
rect 4298 -4423 4350 -4411
rect 4100 -4525 4152 -4457
rect 4100 -4559 4110 -4525
rect 4144 -4559 4152 -4525
rect 4100 -4585 4152 -4559
rect 4298 -4457 4306 -4423
rect 4340 -4457 4350 -4423
rect 4298 -4525 4350 -4457
rect 4298 -4559 4306 -4525
rect 4340 -4559 4350 -4525
rect 4298 -4585 4350 -4559
rect 4928 -4423 4980 -4411
rect 4928 -4457 4938 -4423
rect 4972 -4457 4980 -4423
rect 5126 -4423 5178 -4411
rect 4928 -4525 4980 -4457
rect 4928 -4559 4938 -4525
rect 4972 -4559 4980 -4525
rect 4928 -4585 4980 -4559
rect 5126 -4457 5134 -4423
rect 5168 -4457 5178 -4423
rect 5126 -4525 5178 -4457
rect 5126 -4559 5134 -4525
rect 5168 -4559 5178 -4525
rect 5126 -4585 5178 -4559
rect 5388 -4423 5440 -4411
rect 5388 -4457 5398 -4423
rect 5432 -4457 5440 -4423
rect 5388 -4525 5440 -4457
rect 5388 -4559 5398 -4525
rect 5432 -4559 5440 -4525
rect 5388 -4585 5440 -4559
rect 5586 -4431 5657 -4411
rect 5586 -4465 5609 -4431
rect 5643 -4465 5657 -4431
rect 5586 -4499 5657 -4465
rect 5586 -4533 5609 -4499
rect 5643 -4533 5657 -4499
rect 5586 -4611 5657 -4533
rect 5687 -4430 5752 -4411
rect 5687 -4464 5707 -4430
rect 5741 -4464 5752 -4430
rect 5687 -4498 5752 -4464
rect 5687 -4532 5707 -4498
rect 5741 -4532 5752 -4498
rect 5687 -4575 5752 -4532
rect 5852 -4431 5905 -4411
rect 5852 -4465 5863 -4431
rect 5897 -4465 5905 -4431
rect 5852 -4499 5905 -4465
rect 5852 -4533 5863 -4499
rect 5897 -4533 5905 -4499
rect 5852 -4575 5905 -4533
rect 5959 -4430 6012 -4411
rect 5959 -4464 5967 -4430
rect 6001 -4464 6012 -4430
rect 5959 -4498 6012 -4464
rect 5959 -4532 5967 -4498
rect 6001 -4532 6012 -4498
rect 5959 -4575 6012 -4532
rect 6112 -4430 6184 -4411
rect 6112 -4464 6125 -4430
rect 6159 -4464 6184 -4430
rect 6112 -4498 6184 -4464
rect 6112 -4532 6125 -4498
rect 6159 -4532 6184 -4498
rect 6112 -4575 6184 -4532
rect 5687 -4611 5737 -4575
rect 6134 -4611 6184 -4575
rect 6214 -4430 6268 -4411
rect 6414 -4423 6466 -4411
rect 6214 -4464 6225 -4430
rect 6259 -4464 6268 -4430
rect 6214 -4498 6268 -4464
rect 6214 -4532 6225 -4498
rect 6259 -4532 6268 -4498
rect 6214 -4611 6268 -4532
rect 6414 -4457 6422 -4423
rect 6456 -4457 6466 -4423
rect 6414 -4525 6466 -4457
rect 6414 -4559 6422 -4525
rect 6456 -4559 6466 -4525
rect 6414 -4585 6466 -4559
rect 6676 -4423 6728 -4411
rect 6676 -4457 6686 -4423
rect 6720 -4457 6728 -4423
rect 6874 -4423 6926 -4411
rect 6676 -4525 6728 -4457
rect 6676 -4559 6686 -4525
rect 6720 -4559 6728 -4525
rect 6676 -4585 6728 -4559
rect 6874 -4457 6882 -4423
rect 6916 -4457 6926 -4423
rect 6874 -4525 6926 -4457
rect 6874 -4559 6882 -4525
rect 6916 -4559 6926 -4525
rect 6874 -4585 6926 -4559
rect 7504 -4423 7556 -4411
rect 7504 -4457 7514 -4423
rect 7548 -4457 7556 -4423
rect 7702 -4423 7754 -4411
rect 7504 -4525 7556 -4457
rect 7504 -4559 7514 -4525
rect 7548 -4559 7556 -4525
rect 7504 -4585 7556 -4559
rect 7702 -4457 7710 -4423
rect 7744 -4457 7754 -4423
rect 7702 -4525 7754 -4457
rect 7702 -4559 7710 -4525
rect 7744 -4559 7754 -4525
rect 7702 -4585 7754 -4559
rect 7964 -4423 8016 -4411
rect 7964 -4457 7974 -4423
rect 8008 -4457 8016 -4423
rect 7964 -4525 8016 -4457
rect 7964 -4559 7974 -4525
rect 8008 -4559 8016 -4525
rect 7964 -4585 8016 -4559
rect 8162 -4431 8233 -4411
rect 8162 -4465 8185 -4431
rect 8219 -4465 8233 -4431
rect 8162 -4499 8233 -4465
rect 8162 -4533 8185 -4499
rect 8219 -4533 8233 -4499
rect 8162 -4611 8233 -4533
rect 8263 -4430 8328 -4411
rect 8263 -4464 8283 -4430
rect 8317 -4464 8328 -4430
rect 8263 -4498 8328 -4464
rect 8263 -4532 8283 -4498
rect 8317 -4532 8328 -4498
rect 8263 -4575 8328 -4532
rect 8428 -4431 8481 -4411
rect 8428 -4465 8439 -4431
rect 8473 -4465 8481 -4431
rect 8428 -4499 8481 -4465
rect 8428 -4533 8439 -4499
rect 8473 -4533 8481 -4499
rect 8428 -4575 8481 -4533
rect 8535 -4430 8588 -4411
rect 8535 -4464 8543 -4430
rect 8577 -4464 8588 -4430
rect 8535 -4498 8588 -4464
rect 8535 -4532 8543 -4498
rect 8577 -4532 8588 -4498
rect 8535 -4575 8588 -4532
rect 8688 -4430 8760 -4411
rect 8688 -4464 8701 -4430
rect 8735 -4464 8760 -4430
rect 8688 -4498 8760 -4464
rect 8688 -4532 8701 -4498
rect 8735 -4532 8760 -4498
rect 8688 -4575 8760 -4532
rect 8263 -4611 8313 -4575
rect 8710 -4611 8760 -4575
rect 8790 -4430 8844 -4411
rect 8990 -4423 9042 -4411
rect 8790 -4464 8801 -4430
rect 8835 -4464 8844 -4430
rect 8790 -4498 8844 -4464
rect 8790 -4532 8801 -4498
rect 8835 -4532 8844 -4498
rect 8790 -4611 8844 -4532
rect 8990 -4457 8998 -4423
rect 9032 -4457 9042 -4423
rect 8990 -4525 9042 -4457
rect 8990 -4559 8998 -4525
rect 9032 -4559 9042 -4525
rect 8990 -4585 9042 -4559
rect 9252 -4423 9304 -4411
rect 9252 -4457 9262 -4423
rect 9296 -4457 9304 -4423
rect 9450 -4423 9502 -4411
rect 9252 -4525 9304 -4457
rect 9252 -4559 9262 -4525
rect 9296 -4559 9304 -4525
rect 9252 -4585 9304 -4559
rect 9450 -4457 9458 -4423
rect 9492 -4457 9502 -4423
rect 9450 -4525 9502 -4457
rect 9450 -4559 9458 -4525
rect 9492 -4559 9502 -4525
rect 9450 -4585 9502 -4559
rect 10080 -4423 10132 -4411
rect 10080 -4457 10090 -4423
rect 10124 -4457 10132 -4423
rect 10370 -4423 10422 -4411
rect 10080 -4525 10132 -4457
rect 10080 -4559 10090 -4525
rect 10124 -4559 10132 -4525
rect 10080 -4585 10132 -4559
rect 10370 -4457 10378 -4423
rect 10412 -4457 10422 -4423
rect 10370 -4525 10422 -4457
rect 10370 -4559 10378 -4525
rect 10412 -4559 10422 -4525
rect 10370 -4585 10422 -4559
rect 10632 -4423 10684 -4411
rect 10632 -4457 10642 -4423
rect 10676 -4457 10684 -4423
rect 10632 -4525 10684 -4457
rect 10632 -4559 10642 -4525
rect 10676 -4559 10684 -4525
rect 10632 -4585 10684 -4559
rect 10738 -4431 10809 -4411
rect 10738 -4465 10761 -4431
rect 10795 -4465 10809 -4431
rect 10738 -4499 10809 -4465
rect 10738 -4533 10761 -4499
rect 10795 -4533 10809 -4499
rect 10738 -4611 10809 -4533
rect 10839 -4430 10904 -4411
rect 10839 -4464 10859 -4430
rect 10893 -4464 10904 -4430
rect 10839 -4498 10904 -4464
rect 10839 -4532 10859 -4498
rect 10893 -4532 10904 -4498
rect 10839 -4575 10904 -4532
rect 11004 -4431 11057 -4411
rect 11004 -4465 11015 -4431
rect 11049 -4465 11057 -4431
rect 11004 -4499 11057 -4465
rect 11004 -4533 11015 -4499
rect 11049 -4533 11057 -4499
rect 11004 -4575 11057 -4533
rect 11111 -4430 11164 -4411
rect 11111 -4464 11119 -4430
rect 11153 -4464 11164 -4430
rect 11111 -4498 11164 -4464
rect 11111 -4532 11119 -4498
rect 11153 -4532 11164 -4498
rect 11111 -4575 11164 -4532
rect 11264 -4430 11336 -4411
rect 11264 -4464 11277 -4430
rect 11311 -4464 11336 -4430
rect 11264 -4498 11336 -4464
rect 11264 -4532 11277 -4498
rect 11311 -4532 11336 -4498
rect 11264 -4575 11336 -4532
rect 10839 -4611 10889 -4575
rect 11286 -4611 11336 -4575
rect 11366 -4430 11420 -4411
rect 11658 -4423 11710 -4411
rect 11366 -4464 11377 -4430
rect 11411 -4464 11420 -4430
rect 11366 -4498 11420 -4464
rect 11366 -4532 11377 -4498
rect 11411 -4532 11420 -4498
rect 11366 -4611 11420 -4532
rect 11658 -4457 11666 -4423
rect 11700 -4457 11710 -4423
rect 11658 -4525 11710 -4457
rect 11658 -4559 11666 -4525
rect 11700 -4559 11710 -4525
rect 11658 -4585 11710 -4559
rect 11920 -4423 11972 -4411
rect 11920 -4457 11930 -4423
rect 11964 -4457 11972 -4423
rect 13682 -4423 13735 -4411
rect 11920 -4525 11972 -4457
rect 11920 -4559 11930 -4525
rect 11964 -4559 11972 -4525
rect 11920 -4585 11972 -4559
rect 13682 -4457 13690 -4423
rect 13724 -4457 13735 -4423
rect 13682 -4491 13735 -4457
rect 13682 -4525 13690 -4491
rect 13724 -4525 13735 -4491
rect 13682 -4611 13735 -4525
rect 13765 -4431 13821 -4411
rect 13765 -4465 13776 -4431
rect 13810 -4465 13821 -4431
rect 13765 -4499 13821 -4465
rect 13765 -4533 13776 -4499
rect 13810 -4533 13821 -4499
rect 13765 -4611 13821 -4533
rect 13851 -4423 13907 -4411
rect 13851 -4457 13862 -4423
rect 13896 -4457 13907 -4423
rect 13851 -4491 13907 -4457
rect 13851 -4525 13862 -4491
rect 13896 -4525 13907 -4491
rect 13851 -4611 13907 -4525
rect 13937 -4439 13993 -4411
rect 13937 -4473 13948 -4439
rect 13982 -4473 13993 -4439
rect 13937 -4507 13993 -4473
rect 13937 -4541 13948 -4507
rect 13982 -4541 13993 -4507
rect 13937 -4611 13993 -4541
rect 14023 -4423 14079 -4411
rect 14023 -4457 14034 -4423
rect 14068 -4457 14079 -4423
rect 14023 -4491 14079 -4457
rect 14023 -4525 14034 -4491
rect 14068 -4525 14079 -4491
rect 14023 -4611 14079 -4525
rect 14109 -4467 14165 -4411
rect 14109 -4501 14120 -4467
rect 14154 -4501 14165 -4467
rect 14109 -4553 14165 -4501
rect 14109 -4587 14120 -4553
rect 14154 -4587 14165 -4553
rect 14109 -4611 14165 -4587
rect 14195 -4447 14251 -4411
rect 14195 -4481 14206 -4447
rect 14240 -4481 14251 -4447
rect 14195 -4611 14251 -4481
rect 14281 -4467 14337 -4411
rect 14281 -4501 14292 -4467
rect 14326 -4501 14337 -4467
rect 14281 -4553 14337 -4501
rect 14281 -4587 14292 -4553
rect 14326 -4587 14337 -4553
rect 14281 -4611 14337 -4587
rect 14367 -4447 14423 -4411
rect 14367 -4481 14378 -4447
rect 14412 -4481 14423 -4447
rect 14367 -4611 14423 -4481
rect 14453 -4467 14509 -4411
rect 14453 -4501 14464 -4467
rect 14498 -4501 14509 -4467
rect 14453 -4553 14509 -4501
rect 14453 -4587 14464 -4553
rect 14498 -4587 14509 -4553
rect 14453 -4611 14509 -4587
rect 14539 -4447 14595 -4411
rect 14539 -4481 14550 -4447
rect 14584 -4481 14595 -4447
rect 14539 -4611 14595 -4481
rect 14625 -4467 14681 -4411
rect 14625 -4501 14636 -4467
rect 14670 -4501 14681 -4467
rect 14625 -4553 14681 -4501
rect 14625 -4587 14636 -4553
rect 14670 -4587 14681 -4553
rect 14625 -4611 14681 -4587
rect 14711 -4447 14766 -4411
rect 14711 -4481 14722 -4447
rect 14756 -4481 14766 -4447
rect 14711 -4611 14766 -4481
rect 14796 -4467 14852 -4411
rect 14796 -4501 14807 -4467
rect 14841 -4501 14852 -4467
rect 14796 -4553 14852 -4501
rect 14796 -4587 14807 -4553
rect 14841 -4587 14852 -4553
rect 14796 -4611 14852 -4587
rect 14882 -4447 14938 -4411
rect 14882 -4481 14893 -4447
rect 14927 -4481 14938 -4447
rect 14882 -4611 14938 -4481
rect 14968 -4467 15024 -4411
rect 14968 -4501 14979 -4467
rect 15013 -4501 15024 -4467
rect 14968 -4553 15024 -4501
rect 14968 -4587 14979 -4553
rect 15013 -4587 15024 -4553
rect 14968 -4611 15024 -4587
rect 15054 -4447 15110 -4411
rect 15054 -4481 15065 -4447
rect 15099 -4481 15110 -4447
rect 15054 -4611 15110 -4481
rect 15140 -4467 15196 -4411
rect 15140 -4501 15151 -4467
rect 15185 -4501 15196 -4467
rect 15140 -4553 15196 -4501
rect 15140 -4587 15151 -4553
rect 15185 -4587 15196 -4553
rect 15140 -4611 15196 -4587
rect 15226 -4447 15282 -4411
rect 15226 -4481 15237 -4447
rect 15271 -4481 15282 -4447
rect 15226 -4611 15282 -4481
rect 15312 -4467 15368 -4411
rect 15312 -4501 15323 -4467
rect 15357 -4501 15368 -4467
rect 15312 -4553 15368 -4501
rect 15312 -4587 15323 -4553
rect 15357 -4587 15368 -4553
rect 15312 -4611 15368 -4587
rect 15398 -4447 15451 -4411
rect 15614 -4423 15666 -4411
rect 15398 -4481 15409 -4447
rect 15443 -4481 15451 -4447
rect 15398 -4611 15451 -4481
rect 15614 -4457 15622 -4423
rect 15656 -4457 15666 -4423
rect 15614 -4525 15666 -4457
rect 15614 -4559 15622 -4525
rect 15656 -4559 15666 -4525
rect 15614 -4585 15666 -4559
rect 16612 -4423 16664 -4411
rect 16612 -4457 16622 -4423
rect 16656 -4457 16664 -4423
rect 16612 -4525 16664 -4457
rect 16612 -4559 16622 -4525
rect 16656 -4559 16664 -4525
rect 16612 -4585 16664 -4559
rect -2970 -5257 -2918 -5231
rect -2970 -5291 -2962 -5257
rect -2928 -5291 -2918 -5257
rect -2970 -5359 -2918 -5291
rect -2970 -5393 -2962 -5359
rect -2928 -5393 -2918 -5359
rect -2970 -5405 -2918 -5393
rect -2340 -5257 -2288 -5231
rect -2340 -5291 -2330 -5257
rect -2296 -5291 -2288 -5257
rect -2340 -5359 -2288 -5291
rect -2340 -5393 -2330 -5359
rect -2296 -5393 -2288 -5359
rect -1590 -5257 -1538 -5231
rect -1590 -5291 -1582 -5257
rect -1548 -5291 -1538 -5257
rect -1590 -5359 -1538 -5291
rect -2340 -5405 -2288 -5393
rect -1590 -5393 -1582 -5359
rect -1548 -5393 -1538 -5359
rect -1590 -5405 -1538 -5393
rect -960 -5257 -908 -5231
rect -960 -5291 -950 -5257
rect -916 -5291 -908 -5257
rect -960 -5359 -908 -5291
rect -960 -5393 -950 -5359
rect -916 -5393 -908 -5359
rect -960 -5405 -908 -5393
rect -854 -5257 -802 -5231
rect -854 -5291 -846 -5257
rect -812 -5291 -802 -5257
rect -854 -5359 -802 -5291
rect -854 -5393 -846 -5359
rect -812 -5393 -802 -5359
rect -854 -5405 -802 -5393
rect -224 -5257 -172 -5231
rect -224 -5291 -214 -5257
rect -180 -5291 -172 -5257
rect -224 -5359 -172 -5291
rect -224 -5393 -214 -5359
rect -180 -5393 -172 -5359
rect -26 -5257 26 -5231
rect -26 -5291 -18 -5257
rect 16 -5291 26 -5257
rect -26 -5359 26 -5291
rect -224 -5405 -172 -5393
rect -26 -5393 -18 -5359
rect 16 -5393 26 -5359
rect -26 -5405 26 -5393
rect 236 -5257 288 -5231
rect 236 -5291 246 -5257
rect 280 -5291 288 -5257
rect 236 -5359 288 -5291
rect 236 -5393 246 -5359
rect 280 -5393 288 -5359
rect 434 -5284 488 -5205
rect 434 -5318 443 -5284
rect 477 -5318 488 -5284
rect 434 -5352 488 -5318
rect 434 -5386 443 -5352
rect 477 -5386 488 -5352
rect 236 -5405 288 -5393
rect 434 -5405 488 -5386
rect 518 -5241 568 -5205
rect 965 -5241 1015 -5205
rect 518 -5284 590 -5241
rect 518 -5318 543 -5284
rect 577 -5318 590 -5284
rect 518 -5352 590 -5318
rect 518 -5386 543 -5352
rect 577 -5386 590 -5352
rect 518 -5405 590 -5386
rect 690 -5284 743 -5241
rect 690 -5318 701 -5284
rect 735 -5318 743 -5284
rect 690 -5352 743 -5318
rect 690 -5386 701 -5352
rect 735 -5386 743 -5352
rect 690 -5405 743 -5386
rect 797 -5283 850 -5241
rect 797 -5317 805 -5283
rect 839 -5317 850 -5283
rect 797 -5351 850 -5317
rect 797 -5385 805 -5351
rect 839 -5385 850 -5351
rect 797 -5405 850 -5385
rect 950 -5284 1015 -5241
rect 950 -5318 961 -5284
rect 995 -5318 1015 -5284
rect 950 -5352 1015 -5318
rect 950 -5386 961 -5352
rect 995 -5386 1015 -5352
rect 950 -5405 1015 -5386
rect 1045 -5283 1116 -5205
rect 1045 -5317 1059 -5283
rect 1093 -5317 1116 -5283
rect 1045 -5351 1116 -5317
rect 1045 -5385 1059 -5351
rect 1093 -5385 1116 -5351
rect 1045 -5405 1116 -5385
rect 1262 -5257 1314 -5231
rect 1262 -5291 1270 -5257
rect 1304 -5291 1314 -5257
rect 1262 -5359 1314 -5291
rect 1262 -5393 1270 -5359
rect 1304 -5393 1314 -5359
rect 1262 -5405 1314 -5393
rect 1524 -5257 1576 -5231
rect 1524 -5291 1534 -5257
rect 1568 -5291 1576 -5257
rect 1524 -5359 1576 -5291
rect 1524 -5393 1534 -5359
rect 1568 -5393 1576 -5359
rect 1722 -5257 1774 -5231
rect 1722 -5291 1730 -5257
rect 1764 -5291 1774 -5257
rect 1722 -5359 1774 -5291
rect 1524 -5405 1576 -5393
rect 1722 -5393 1730 -5359
rect 1764 -5393 1774 -5359
rect 1722 -5405 1774 -5393
rect 2352 -5257 2404 -5231
rect 2352 -5291 2362 -5257
rect 2396 -5291 2404 -5257
rect 2352 -5359 2404 -5291
rect 2352 -5393 2362 -5359
rect 2396 -5393 2404 -5359
rect 2550 -5257 2602 -5231
rect 2550 -5291 2558 -5257
rect 2592 -5291 2602 -5257
rect 2550 -5359 2602 -5291
rect 2352 -5405 2404 -5393
rect 2550 -5393 2558 -5359
rect 2592 -5393 2602 -5359
rect 2550 -5405 2602 -5393
rect 2812 -5257 2864 -5231
rect 2812 -5291 2822 -5257
rect 2856 -5291 2864 -5257
rect 2812 -5359 2864 -5291
rect 2812 -5393 2822 -5359
rect 2856 -5393 2864 -5359
rect 3010 -5284 3064 -5205
rect 3010 -5318 3019 -5284
rect 3053 -5318 3064 -5284
rect 3010 -5352 3064 -5318
rect 3010 -5386 3019 -5352
rect 3053 -5386 3064 -5352
rect 2812 -5405 2864 -5393
rect 3010 -5405 3064 -5386
rect 3094 -5241 3144 -5205
rect 3541 -5241 3591 -5205
rect 3094 -5284 3166 -5241
rect 3094 -5318 3119 -5284
rect 3153 -5318 3166 -5284
rect 3094 -5352 3166 -5318
rect 3094 -5386 3119 -5352
rect 3153 -5386 3166 -5352
rect 3094 -5405 3166 -5386
rect 3266 -5284 3319 -5241
rect 3266 -5318 3277 -5284
rect 3311 -5318 3319 -5284
rect 3266 -5352 3319 -5318
rect 3266 -5386 3277 -5352
rect 3311 -5386 3319 -5352
rect 3266 -5405 3319 -5386
rect 3373 -5283 3426 -5241
rect 3373 -5317 3381 -5283
rect 3415 -5317 3426 -5283
rect 3373 -5351 3426 -5317
rect 3373 -5385 3381 -5351
rect 3415 -5385 3426 -5351
rect 3373 -5405 3426 -5385
rect 3526 -5284 3591 -5241
rect 3526 -5318 3537 -5284
rect 3571 -5318 3591 -5284
rect 3526 -5352 3591 -5318
rect 3526 -5386 3537 -5352
rect 3571 -5386 3591 -5352
rect 3526 -5405 3591 -5386
rect 3621 -5283 3692 -5205
rect 3621 -5317 3635 -5283
rect 3669 -5317 3692 -5283
rect 3621 -5351 3692 -5317
rect 3621 -5385 3635 -5351
rect 3669 -5385 3692 -5351
rect 3621 -5405 3692 -5385
rect 3838 -5257 3890 -5231
rect 3838 -5291 3846 -5257
rect 3880 -5291 3890 -5257
rect 3838 -5359 3890 -5291
rect 3838 -5393 3846 -5359
rect 3880 -5393 3890 -5359
rect 3838 -5405 3890 -5393
rect 4100 -5257 4152 -5231
rect 4100 -5291 4110 -5257
rect 4144 -5291 4152 -5257
rect 4100 -5359 4152 -5291
rect 4100 -5393 4110 -5359
rect 4144 -5393 4152 -5359
rect 4298 -5257 4350 -5231
rect 4298 -5291 4306 -5257
rect 4340 -5291 4350 -5257
rect 4298 -5359 4350 -5291
rect 4100 -5405 4152 -5393
rect 4298 -5393 4306 -5359
rect 4340 -5393 4350 -5359
rect 4298 -5405 4350 -5393
rect 4928 -5257 4980 -5231
rect 4928 -5291 4938 -5257
rect 4972 -5291 4980 -5257
rect 4928 -5359 4980 -5291
rect 4928 -5393 4938 -5359
rect 4972 -5393 4980 -5359
rect 5126 -5257 5178 -5231
rect 5126 -5291 5134 -5257
rect 5168 -5291 5178 -5257
rect 5126 -5359 5178 -5291
rect 4928 -5405 4980 -5393
rect 5126 -5393 5134 -5359
rect 5168 -5393 5178 -5359
rect 5126 -5405 5178 -5393
rect 5388 -5257 5440 -5231
rect 5388 -5291 5398 -5257
rect 5432 -5291 5440 -5257
rect 5388 -5359 5440 -5291
rect 5388 -5393 5398 -5359
rect 5432 -5393 5440 -5359
rect 5586 -5284 5640 -5205
rect 5586 -5318 5595 -5284
rect 5629 -5318 5640 -5284
rect 5586 -5352 5640 -5318
rect 5586 -5386 5595 -5352
rect 5629 -5386 5640 -5352
rect 5388 -5405 5440 -5393
rect 5586 -5405 5640 -5386
rect 5670 -5241 5720 -5205
rect 6117 -5241 6167 -5205
rect 5670 -5284 5742 -5241
rect 5670 -5318 5695 -5284
rect 5729 -5318 5742 -5284
rect 5670 -5352 5742 -5318
rect 5670 -5386 5695 -5352
rect 5729 -5386 5742 -5352
rect 5670 -5405 5742 -5386
rect 5842 -5284 5895 -5241
rect 5842 -5318 5853 -5284
rect 5887 -5318 5895 -5284
rect 5842 -5352 5895 -5318
rect 5842 -5386 5853 -5352
rect 5887 -5386 5895 -5352
rect 5842 -5405 5895 -5386
rect 5949 -5283 6002 -5241
rect 5949 -5317 5957 -5283
rect 5991 -5317 6002 -5283
rect 5949 -5351 6002 -5317
rect 5949 -5385 5957 -5351
rect 5991 -5385 6002 -5351
rect 5949 -5405 6002 -5385
rect 6102 -5284 6167 -5241
rect 6102 -5318 6113 -5284
rect 6147 -5318 6167 -5284
rect 6102 -5352 6167 -5318
rect 6102 -5386 6113 -5352
rect 6147 -5386 6167 -5352
rect 6102 -5405 6167 -5386
rect 6197 -5283 6268 -5205
rect 6197 -5317 6211 -5283
rect 6245 -5317 6268 -5283
rect 6197 -5351 6268 -5317
rect 6197 -5385 6211 -5351
rect 6245 -5385 6268 -5351
rect 6197 -5405 6268 -5385
rect 6414 -5257 6466 -5231
rect 6414 -5291 6422 -5257
rect 6456 -5291 6466 -5257
rect 6414 -5359 6466 -5291
rect 6414 -5393 6422 -5359
rect 6456 -5393 6466 -5359
rect 6414 -5405 6466 -5393
rect 6676 -5257 6728 -5231
rect 6676 -5291 6686 -5257
rect 6720 -5291 6728 -5257
rect 6676 -5359 6728 -5291
rect 6676 -5393 6686 -5359
rect 6720 -5393 6728 -5359
rect 6874 -5257 6926 -5231
rect 6874 -5291 6882 -5257
rect 6916 -5291 6926 -5257
rect 6874 -5359 6926 -5291
rect 6676 -5405 6728 -5393
rect 6874 -5393 6882 -5359
rect 6916 -5393 6926 -5359
rect 6874 -5405 6926 -5393
rect 7504 -5257 7556 -5231
rect 7504 -5291 7514 -5257
rect 7548 -5291 7556 -5257
rect 7504 -5359 7556 -5291
rect 7504 -5393 7514 -5359
rect 7548 -5393 7556 -5359
rect 7702 -5257 7754 -5231
rect 7702 -5291 7710 -5257
rect 7744 -5291 7754 -5257
rect 7702 -5359 7754 -5291
rect 7504 -5405 7556 -5393
rect 7702 -5393 7710 -5359
rect 7744 -5393 7754 -5359
rect 7702 -5405 7754 -5393
rect 7964 -5257 8016 -5231
rect 7964 -5291 7974 -5257
rect 8008 -5291 8016 -5257
rect 7964 -5359 8016 -5291
rect 7964 -5393 7974 -5359
rect 8008 -5393 8016 -5359
rect 8162 -5284 8216 -5205
rect 8162 -5318 8171 -5284
rect 8205 -5318 8216 -5284
rect 8162 -5352 8216 -5318
rect 8162 -5386 8171 -5352
rect 8205 -5386 8216 -5352
rect 7964 -5405 8016 -5393
rect 8162 -5405 8216 -5386
rect 8246 -5241 8296 -5205
rect 8693 -5241 8743 -5205
rect 8246 -5284 8318 -5241
rect 8246 -5318 8271 -5284
rect 8305 -5318 8318 -5284
rect 8246 -5352 8318 -5318
rect 8246 -5386 8271 -5352
rect 8305 -5386 8318 -5352
rect 8246 -5405 8318 -5386
rect 8418 -5284 8471 -5241
rect 8418 -5318 8429 -5284
rect 8463 -5318 8471 -5284
rect 8418 -5352 8471 -5318
rect 8418 -5386 8429 -5352
rect 8463 -5386 8471 -5352
rect 8418 -5405 8471 -5386
rect 8525 -5283 8578 -5241
rect 8525 -5317 8533 -5283
rect 8567 -5317 8578 -5283
rect 8525 -5351 8578 -5317
rect 8525 -5385 8533 -5351
rect 8567 -5385 8578 -5351
rect 8525 -5405 8578 -5385
rect 8678 -5284 8743 -5241
rect 8678 -5318 8689 -5284
rect 8723 -5318 8743 -5284
rect 8678 -5352 8743 -5318
rect 8678 -5386 8689 -5352
rect 8723 -5386 8743 -5352
rect 8678 -5405 8743 -5386
rect 8773 -5283 8844 -5205
rect 8773 -5317 8787 -5283
rect 8821 -5317 8844 -5283
rect 8773 -5351 8844 -5317
rect 8773 -5385 8787 -5351
rect 8821 -5385 8844 -5351
rect 8773 -5405 8844 -5385
rect 8990 -5257 9042 -5231
rect 8990 -5291 8998 -5257
rect 9032 -5291 9042 -5257
rect 8990 -5359 9042 -5291
rect 8990 -5393 8998 -5359
rect 9032 -5393 9042 -5359
rect 8990 -5405 9042 -5393
rect 9252 -5257 9304 -5231
rect 9252 -5291 9262 -5257
rect 9296 -5291 9304 -5257
rect 9252 -5359 9304 -5291
rect 9252 -5393 9262 -5359
rect 9296 -5393 9304 -5359
rect 9450 -5257 9502 -5231
rect 9450 -5291 9458 -5257
rect 9492 -5291 9502 -5257
rect 9450 -5359 9502 -5291
rect 9252 -5405 9304 -5393
rect 9450 -5393 9458 -5359
rect 9492 -5393 9502 -5359
rect 9450 -5405 9502 -5393
rect 10080 -5257 10132 -5231
rect 10080 -5291 10090 -5257
rect 10124 -5291 10132 -5257
rect 10080 -5359 10132 -5291
rect 10080 -5393 10090 -5359
rect 10124 -5393 10132 -5359
rect 10370 -5257 10422 -5231
rect 10370 -5291 10378 -5257
rect 10412 -5291 10422 -5257
rect 10370 -5359 10422 -5291
rect 10080 -5405 10132 -5393
rect 10370 -5393 10378 -5359
rect 10412 -5393 10422 -5359
rect 10370 -5405 10422 -5393
rect 10632 -5257 10684 -5231
rect 10632 -5291 10642 -5257
rect 10676 -5291 10684 -5257
rect 10632 -5359 10684 -5291
rect 10632 -5393 10642 -5359
rect 10676 -5393 10684 -5359
rect 10632 -5405 10684 -5393
rect 10738 -5284 10792 -5205
rect 10738 -5318 10747 -5284
rect 10781 -5318 10792 -5284
rect 10738 -5352 10792 -5318
rect 10738 -5386 10747 -5352
rect 10781 -5386 10792 -5352
rect 10738 -5405 10792 -5386
rect 10822 -5241 10872 -5205
rect 11269 -5241 11319 -5205
rect 10822 -5284 10894 -5241
rect 10822 -5318 10847 -5284
rect 10881 -5318 10894 -5284
rect 10822 -5352 10894 -5318
rect 10822 -5386 10847 -5352
rect 10881 -5386 10894 -5352
rect 10822 -5405 10894 -5386
rect 10994 -5284 11047 -5241
rect 10994 -5318 11005 -5284
rect 11039 -5318 11047 -5284
rect 10994 -5352 11047 -5318
rect 10994 -5386 11005 -5352
rect 11039 -5386 11047 -5352
rect 10994 -5405 11047 -5386
rect 11101 -5283 11154 -5241
rect 11101 -5317 11109 -5283
rect 11143 -5317 11154 -5283
rect 11101 -5351 11154 -5317
rect 11101 -5385 11109 -5351
rect 11143 -5385 11154 -5351
rect 11101 -5405 11154 -5385
rect 11254 -5284 11319 -5241
rect 11254 -5318 11265 -5284
rect 11299 -5318 11319 -5284
rect 11254 -5352 11319 -5318
rect 11254 -5386 11265 -5352
rect 11299 -5386 11319 -5352
rect 11254 -5405 11319 -5386
rect 11349 -5283 11420 -5205
rect 11349 -5317 11363 -5283
rect 11397 -5317 11420 -5283
rect 11349 -5351 11420 -5317
rect 11349 -5385 11363 -5351
rect 11397 -5385 11420 -5351
rect 11349 -5405 11420 -5385
rect 11658 -5257 11710 -5231
rect 11658 -5291 11666 -5257
rect 11700 -5291 11710 -5257
rect 11658 -5359 11710 -5291
rect 11658 -5393 11666 -5359
rect 11700 -5393 11710 -5359
rect 11658 -5405 11710 -5393
rect 11920 -5257 11972 -5231
rect 11920 -5291 11930 -5257
rect 11964 -5291 11972 -5257
rect 11920 -5359 11972 -5291
rect 11920 -5393 11930 -5359
rect 11964 -5393 11972 -5359
rect 12486 -5284 12547 -5205
rect 12486 -5318 12502 -5284
rect 12536 -5318 12547 -5284
rect 12486 -5352 12547 -5318
rect 12486 -5386 12502 -5352
rect 12536 -5386 12547 -5352
rect 11920 -5405 11972 -5393
rect 12486 -5405 12547 -5386
rect 12577 -5257 12633 -5205
rect 12577 -5291 12588 -5257
rect 12622 -5291 12633 -5257
rect 12577 -5345 12633 -5291
rect 12577 -5379 12588 -5345
rect 12622 -5379 12633 -5345
rect 12577 -5405 12633 -5379
rect 12663 -5284 12719 -5205
rect 12663 -5318 12674 -5284
rect 12708 -5318 12719 -5284
rect 12663 -5352 12719 -5318
rect 12663 -5386 12674 -5352
rect 12708 -5386 12719 -5352
rect 12663 -5405 12719 -5386
rect 12749 -5257 12805 -5205
rect 12749 -5291 12760 -5257
rect 12794 -5291 12805 -5257
rect 12749 -5345 12805 -5291
rect 12749 -5379 12760 -5345
rect 12794 -5379 12805 -5345
rect 12749 -5405 12805 -5379
rect 12835 -5284 12891 -5205
rect 12835 -5318 12846 -5284
rect 12880 -5318 12891 -5284
rect 12835 -5352 12891 -5318
rect 12835 -5386 12846 -5352
rect 12880 -5386 12891 -5352
rect 12835 -5405 12891 -5386
rect 12921 -5257 12977 -5205
rect 12921 -5291 12932 -5257
rect 12966 -5291 12977 -5257
rect 12921 -5345 12977 -5291
rect 12921 -5379 12932 -5345
rect 12966 -5379 12977 -5345
rect 12921 -5405 12977 -5379
rect 13007 -5284 13076 -5205
rect 13007 -5318 13018 -5284
rect 13052 -5318 13076 -5284
rect 13007 -5352 13076 -5318
rect 13007 -5386 13018 -5352
rect 13052 -5386 13076 -5352
rect 13007 -5405 13076 -5386
rect 13222 -5257 13274 -5231
rect 13222 -5291 13230 -5257
rect 13264 -5291 13274 -5257
rect 13222 -5359 13274 -5291
rect 13222 -5393 13230 -5359
rect 13264 -5393 13274 -5359
rect 13222 -5405 13274 -5393
rect 13484 -5257 13536 -5231
rect 13484 -5291 13494 -5257
rect 13528 -5291 13536 -5257
rect 13484 -5359 13536 -5291
rect 13484 -5393 13494 -5359
rect 13528 -5393 13536 -5359
rect 13682 -5291 13735 -5205
rect 13682 -5325 13690 -5291
rect 13724 -5325 13735 -5291
rect 13682 -5359 13735 -5325
rect 13484 -5405 13536 -5393
rect 13682 -5393 13690 -5359
rect 13724 -5393 13735 -5359
rect 13682 -5405 13735 -5393
rect 13765 -5283 13821 -5205
rect 13765 -5317 13776 -5283
rect 13810 -5317 13821 -5283
rect 13765 -5351 13821 -5317
rect 13765 -5385 13776 -5351
rect 13810 -5385 13821 -5351
rect 13765 -5405 13821 -5385
rect 13851 -5291 13907 -5205
rect 13851 -5325 13862 -5291
rect 13896 -5325 13907 -5291
rect 13851 -5359 13907 -5325
rect 13851 -5393 13862 -5359
rect 13896 -5393 13907 -5359
rect 13851 -5405 13907 -5393
rect 13937 -5275 13993 -5205
rect 13937 -5309 13948 -5275
rect 13982 -5309 13993 -5275
rect 13937 -5343 13993 -5309
rect 13937 -5377 13948 -5343
rect 13982 -5377 13993 -5343
rect 13937 -5405 13993 -5377
rect 14023 -5291 14079 -5205
rect 14023 -5325 14034 -5291
rect 14068 -5325 14079 -5291
rect 14023 -5359 14079 -5325
rect 14023 -5393 14034 -5359
rect 14068 -5393 14079 -5359
rect 14023 -5405 14079 -5393
rect 14109 -5229 14165 -5205
rect 14109 -5263 14120 -5229
rect 14154 -5263 14165 -5229
rect 14109 -5315 14165 -5263
rect 14109 -5349 14120 -5315
rect 14154 -5349 14165 -5315
rect 14109 -5405 14165 -5349
rect 14195 -5335 14251 -5205
rect 14195 -5369 14206 -5335
rect 14240 -5369 14251 -5335
rect 14195 -5405 14251 -5369
rect 14281 -5229 14337 -5205
rect 14281 -5263 14292 -5229
rect 14326 -5263 14337 -5229
rect 14281 -5315 14337 -5263
rect 14281 -5349 14292 -5315
rect 14326 -5349 14337 -5315
rect 14281 -5405 14337 -5349
rect 14367 -5335 14423 -5205
rect 14367 -5369 14378 -5335
rect 14412 -5369 14423 -5335
rect 14367 -5405 14423 -5369
rect 14453 -5229 14509 -5205
rect 14453 -5263 14464 -5229
rect 14498 -5263 14509 -5229
rect 14453 -5315 14509 -5263
rect 14453 -5349 14464 -5315
rect 14498 -5349 14509 -5315
rect 14453 -5405 14509 -5349
rect 14539 -5335 14595 -5205
rect 14539 -5369 14550 -5335
rect 14584 -5369 14595 -5335
rect 14539 -5405 14595 -5369
rect 14625 -5229 14681 -5205
rect 14625 -5263 14636 -5229
rect 14670 -5263 14681 -5229
rect 14625 -5315 14681 -5263
rect 14625 -5349 14636 -5315
rect 14670 -5349 14681 -5315
rect 14625 -5405 14681 -5349
rect 14711 -5335 14766 -5205
rect 14711 -5369 14722 -5335
rect 14756 -5369 14766 -5335
rect 14711 -5405 14766 -5369
rect 14796 -5229 14852 -5205
rect 14796 -5263 14807 -5229
rect 14841 -5263 14852 -5229
rect 14796 -5315 14852 -5263
rect 14796 -5349 14807 -5315
rect 14841 -5349 14852 -5315
rect 14796 -5405 14852 -5349
rect 14882 -5335 14938 -5205
rect 14882 -5369 14893 -5335
rect 14927 -5369 14938 -5335
rect 14882 -5405 14938 -5369
rect 14968 -5229 15024 -5205
rect 14968 -5263 14979 -5229
rect 15013 -5263 15024 -5229
rect 14968 -5315 15024 -5263
rect 14968 -5349 14979 -5315
rect 15013 -5349 15024 -5315
rect 14968 -5405 15024 -5349
rect 15054 -5335 15110 -5205
rect 15054 -5369 15065 -5335
rect 15099 -5369 15110 -5335
rect 15054 -5405 15110 -5369
rect 15140 -5229 15196 -5205
rect 15140 -5263 15151 -5229
rect 15185 -5263 15196 -5229
rect 15140 -5315 15196 -5263
rect 15140 -5349 15151 -5315
rect 15185 -5349 15196 -5315
rect 15140 -5405 15196 -5349
rect 15226 -5335 15282 -5205
rect 15226 -5369 15237 -5335
rect 15271 -5369 15282 -5335
rect 15226 -5405 15282 -5369
rect 15312 -5229 15368 -5205
rect 15312 -5263 15323 -5229
rect 15357 -5263 15368 -5229
rect 15312 -5315 15368 -5263
rect 15312 -5349 15323 -5315
rect 15357 -5349 15368 -5315
rect 15312 -5405 15368 -5349
rect 15398 -5335 15451 -5205
rect 15398 -5369 15409 -5335
rect 15443 -5369 15451 -5335
rect 15398 -5405 15451 -5369
rect 15614 -5257 15666 -5231
rect 15614 -5291 15622 -5257
rect 15656 -5291 15666 -5257
rect 15614 -5359 15666 -5291
rect 15614 -5393 15622 -5359
rect 15656 -5393 15666 -5359
rect 15614 -5405 15666 -5393
rect 16612 -5257 16664 -5231
rect 16612 -5291 16622 -5257
rect 16656 -5291 16664 -5257
rect 16612 -5359 16664 -5291
rect 16612 -5393 16622 -5359
rect 16656 -5393 16664 -5359
rect 16612 -5405 16664 -5393
rect -2970 -5511 -2918 -5499
rect -2970 -5545 -2962 -5511
rect -2928 -5545 -2918 -5511
rect -2970 -5613 -2918 -5545
rect -2970 -5647 -2962 -5613
rect -2928 -5647 -2918 -5613
rect -2970 -5673 -2918 -5647
rect -2340 -5511 -2288 -5499
rect -2340 -5545 -2330 -5511
rect -2296 -5545 -2288 -5511
rect -1590 -5511 -1538 -5499
rect -2340 -5613 -2288 -5545
rect -2340 -5647 -2330 -5613
rect -2296 -5647 -2288 -5613
rect -2340 -5673 -2288 -5647
rect -1590 -5545 -1582 -5511
rect -1548 -5545 -1538 -5511
rect -1590 -5613 -1538 -5545
rect -1590 -5647 -1582 -5613
rect -1548 -5647 -1538 -5613
rect -1590 -5673 -1538 -5647
rect -960 -5511 -908 -5499
rect -960 -5545 -950 -5511
rect -916 -5545 -908 -5511
rect -960 -5613 -908 -5545
rect -960 -5647 -950 -5613
rect -916 -5647 -908 -5613
rect -960 -5673 -908 -5647
rect -854 -5511 -802 -5499
rect -854 -5545 -846 -5511
rect -812 -5545 -802 -5511
rect -854 -5613 -802 -5545
rect -854 -5647 -846 -5613
rect -812 -5647 -802 -5613
rect -854 -5673 -802 -5647
rect -224 -5511 -172 -5499
rect -224 -5545 -214 -5511
rect -180 -5545 -172 -5511
rect -26 -5511 26 -5499
rect -224 -5613 -172 -5545
rect -224 -5647 -214 -5613
rect -180 -5647 -172 -5613
rect -224 -5673 -172 -5647
rect -26 -5545 -18 -5511
rect 16 -5545 26 -5511
rect -26 -5613 26 -5545
rect -26 -5647 -18 -5613
rect 16 -5647 26 -5613
rect -26 -5673 26 -5647
rect 236 -5511 288 -5499
rect 236 -5545 246 -5511
rect 280 -5545 288 -5511
rect 236 -5613 288 -5545
rect 236 -5647 246 -5613
rect 280 -5647 288 -5613
rect 236 -5673 288 -5647
rect 434 -5519 505 -5499
rect 434 -5553 457 -5519
rect 491 -5553 505 -5519
rect 434 -5587 505 -5553
rect 434 -5621 457 -5587
rect 491 -5621 505 -5587
rect 434 -5699 505 -5621
rect 535 -5518 600 -5499
rect 535 -5552 555 -5518
rect 589 -5552 600 -5518
rect 535 -5586 600 -5552
rect 535 -5620 555 -5586
rect 589 -5620 600 -5586
rect 535 -5663 600 -5620
rect 700 -5519 753 -5499
rect 700 -5553 711 -5519
rect 745 -5553 753 -5519
rect 700 -5587 753 -5553
rect 700 -5621 711 -5587
rect 745 -5621 753 -5587
rect 700 -5663 753 -5621
rect 807 -5518 860 -5499
rect 807 -5552 815 -5518
rect 849 -5552 860 -5518
rect 807 -5586 860 -5552
rect 807 -5620 815 -5586
rect 849 -5620 860 -5586
rect 807 -5663 860 -5620
rect 960 -5518 1032 -5499
rect 960 -5552 973 -5518
rect 1007 -5552 1032 -5518
rect 960 -5586 1032 -5552
rect 960 -5620 973 -5586
rect 1007 -5620 1032 -5586
rect 960 -5663 1032 -5620
rect 535 -5699 585 -5663
rect 982 -5699 1032 -5663
rect 1062 -5518 1116 -5499
rect 1262 -5511 1314 -5499
rect 1062 -5552 1073 -5518
rect 1107 -5552 1116 -5518
rect 1062 -5586 1116 -5552
rect 1062 -5620 1073 -5586
rect 1107 -5620 1116 -5586
rect 1062 -5699 1116 -5620
rect 1262 -5545 1270 -5511
rect 1304 -5545 1314 -5511
rect 1262 -5613 1314 -5545
rect 1262 -5647 1270 -5613
rect 1304 -5647 1314 -5613
rect 1262 -5673 1314 -5647
rect 1524 -5511 1576 -5499
rect 1524 -5545 1534 -5511
rect 1568 -5545 1576 -5511
rect 1722 -5511 1774 -5499
rect 1524 -5613 1576 -5545
rect 1524 -5647 1534 -5613
rect 1568 -5647 1576 -5613
rect 1524 -5673 1576 -5647
rect 1722 -5545 1730 -5511
rect 1764 -5545 1774 -5511
rect 1722 -5613 1774 -5545
rect 1722 -5647 1730 -5613
rect 1764 -5647 1774 -5613
rect 1722 -5673 1774 -5647
rect 2352 -5511 2404 -5499
rect 2352 -5545 2362 -5511
rect 2396 -5545 2404 -5511
rect 2550 -5511 2602 -5499
rect 2352 -5613 2404 -5545
rect 2352 -5647 2362 -5613
rect 2396 -5647 2404 -5613
rect 2352 -5673 2404 -5647
rect 2550 -5545 2558 -5511
rect 2592 -5545 2602 -5511
rect 2550 -5613 2602 -5545
rect 2550 -5647 2558 -5613
rect 2592 -5647 2602 -5613
rect 2550 -5673 2602 -5647
rect 2812 -5511 2864 -5499
rect 2812 -5545 2822 -5511
rect 2856 -5545 2864 -5511
rect 2812 -5613 2864 -5545
rect 2812 -5647 2822 -5613
rect 2856 -5647 2864 -5613
rect 2812 -5673 2864 -5647
rect 3010 -5519 3081 -5499
rect 3010 -5553 3033 -5519
rect 3067 -5553 3081 -5519
rect 3010 -5587 3081 -5553
rect 3010 -5621 3033 -5587
rect 3067 -5621 3081 -5587
rect 3010 -5699 3081 -5621
rect 3111 -5518 3176 -5499
rect 3111 -5552 3131 -5518
rect 3165 -5552 3176 -5518
rect 3111 -5586 3176 -5552
rect 3111 -5620 3131 -5586
rect 3165 -5620 3176 -5586
rect 3111 -5663 3176 -5620
rect 3276 -5519 3329 -5499
rect 3276 -5553 3287 -5519
rect 3321 -5553 3329 -5519
rect 3276 -5587 3329 -5553
rect 3276 -5621 3287 -5587
rect 3321 -5621 3329 -5587
rect 3276 -5663 3329 -5621
rect 3383 -5518 3436 -5499
rect 3383 -5552 3391 -5518
rect 3425 -5552 3436 -5518
rect 3383 -5586 3436 -5552
rect 3383 -5620 3391 -5586
rect 3425 -5620 3436 -5586
rect 3383 -5663 3436 -5620
rect 3536 -5518 3608 -5499
rect 3536 -5552 3549 -5518
rect 3583 -5552 3608 -5518
rect 3536 -5586 3608 -5552
rect 3536 -5620 3549 -5586
rect 3583 -5620 3608 -5586
rect 3536 -5663 3608 -5620
rect 3111 -5699 3161 -5663
rect 3558 -5699 3608 -5663
rect 3638 -5518 3692 -5499
rect 3838 -5511 3890 -5499
rect 3638 -5552 3649 -5518
rect 3683 -5552 3692 -5518
rect 3638 -5586 3692 -5552
rect 3638 -5620 3649 -5586
rect 3683 -5620 3692 -5586
rect 3638 -5699 3692 -5620
rect 3838 -5545 3846 -5511
rect 3880 -5545 3890 -5511
rect 3838 -5613 3890 -5545
rect 3838 -5647 3846 -5613
rect 3880 -5647 3890 -5613
rect 3838 -5673 3890 -5647
rect 4100 -5511 4152 -5499
rect 4100 -5545 4110 -5511
rect 4144 -5545 4152 -5511
rect 4298 -5511 4350 -5499
rect 4100 -5613 4152 -5545
rect 4100 -5647 4110 -5613
rect 4144 -5647 4152 -5613
rect 4100 -5673 4152 -5647
rect 4298 -5545 4306 -5511
rect 4340 -5545 4350 -5511
rect 4298 -5613 4350 -5545
rect 4298 -5647 4306 -5613
rect 4340 -5647 4350 -5613
rect 4298 -5673 4350 -5647
rect 4928 -5511 4980 -5499
rect 4928 -5545 4938 -5511
rect 4972 -5545 4980 -5511
rect 5126 -5511 5178 -5499
rect 4928 -5613 4980 -5545
rect 4928 -5647 4938 -5613
rect 4972 -5647 4980 -5613
rect 4928 -5673 4980 -5647
rect 5126 -5545 5134 -5511
rect 5168 -5545 5178 -5511
rect 5126 -5613 5178 -5545
rect 5126 -5647 5134 -5613
rect 5168 -5647 5178 -5613
rect 5126 -5673 5178 -5647
rect 5388 -5511 5440 -5499
rect 5388 -5545 5398 -5511
rect 5432 -5545 5440 -5511
rect 5388 -5613 5440 -5545
rect 5388 -5647 5398 -5613
rect 5432 -5647 5440 -5613
rect 5388 -5673 5440 -5647
rect 5586 -5519 5657 -5499
rect 5586 -5553 5609 -5519
rect 5643 -5553 5657 -5519
rect 5586 -5587 5657 -5553
rect 5586 -5621 5609 -5587
rect 5643 -5621 5657 -5587
rect 5586 -5699 5657 -5621
rect 5687 -5518 5752 -5499
rect 5687 -5552 5707 -5518
rect 5741 -5552 5752 -5518
rect 5687 -5586 5752 -5552
rect 5687 -5620 5707 -5586
rect 5741 -5620 5752 -5586
rect 5687 -5663 5752 -5620
rect 5852 -5519 5905 -5499
rect 5852 -5553 5863 -5519
rect 5897 -5553 5905 -5519
rect 5852 -5587 5905 -5553
rect 5852 -5621 5863 -5587
rect 5897 -5621 5905 -5587
rect 5852 -5663 5905 -5621
rect 5959 -5518 6012 -5499
rect 5959 -5552 5967 -5518
rect 6001 -5552 6012 -5518
rect 5959 -5586 6012 -5552
rect 5959 -5620 5967 -5586
rect 6001 -5620 6012 -5586
rect 5959 -5663 6012 -5620
rect 6112 -5518 6184 -5499
rect 6112 -5552 6125 -5518
rect 6159 -5552 6184 -5518
rect 6112 -5586 6184 -5552
rect 6112 -5620 6125 -5586
rect 6159 -5620 6184 -5586
rect 6112 -5663 6184 -5620
rect 5687 -5699 5737 -5663
rect 6134 -5699 6184 -5663
rect 6214 -5518 6268 -5499
rect 6414 -5511 6466 -5499
rect 6214 -5552 6225 -5518
rect 6259 -5552 6268 -5518
rect 6214 -5586 6268 -5552
rect 6214 -5620 6225 -5586
rect 6259 -5620 6268 -5586
rect 6214 -5699 6268 -5620
rect 6414 -5545 6422 -5511
rect 6456 -5545 6466 -5511
rect 6414 -5613 6466 -5545
rect 6414 -5647 6422 -5613
rect 6456 -5647 6466 -5613
rect 6414 -5673 6466 -5647
rect 6676 -5511 6728 -5499
rect 6676 -5545 6686 -5511
rect 6720 -5545 6728 -5511
rect 6874 -5511 6926 -5499
rect 6676 -5613 6728 -5545
rect 6676 -5647 6686 -5613
rect 6720 -5647 6728 -5613
rect 6676 -5673 6728 -5647
rect 6874 -5545 6882 -5511
rect 6916 -5545 6926 -5511
rect 6874 -5613 6926 -5545
rect 6874 -5647 6882 -5613
rect 6916 -5647 6926 -5613
rect 6874 -5673 6926 -5647
rect 7504 -5511 7556 -5499
rect 7504 -5545 7514 -5511
rect 7548 -5545 7556 -5511
rect 7702 -5511 7754 -5499
rect 7504 -5613 7556 -5545
rect 7504 -5647 7514 -5613
rect 7548 -5647 7556 -5613
rect 7504 -5673 7556 -5647
rect 7702 -5545 7710 -5511
rect 7744 -5545 7754 -5511
rect 7702 -5613 7754 -5545
rect 7702 -5647 7710 -5613
rect 7744 -5647 7754 -5613
rect 7702 -5673 7754 -5647
rect 7964 -5511 8016 -5499
rect 7964 -5545 7974 -5511
rect 8008 -5545 8016 -5511
rect 7964 -5613 8016 -5545
rect 7964 -5647 7974 -5613
rect 8008 -5647 8016 -5613
rect 7964 -5673 8016 -5647
rect 8162 -5519 8233 -5499
rect 8162 -5553 8185 -5519
rect 8219 -5553 8233 -5519
rect 8162 -5587 8233 -5553
rect 8162 -5621 8185 -5587
rect 8219 -5621 8233 -5587
rect 8162 -5699 8233 -5621
rect 8263 -5518 8328 -5499
rect 8263 -5552 8283 -5518
rect 8317 -5552 8328 -5518
rect 8263 -5586 8328 -5552
rect 8263 -5620 8283 -5586
rect 8317 -5620 8328 -5586
rect 8263 -5663 8328 -5620
rect 8428 -5519 8481 -5499
rect 8428 -5553 8439 -5519
rect 8473 -5553 8481 -5519
rect 8428 -5587 8481 -5553
rect 8428 -5621 8439 -5587
rect 8473 -5621 8481 -5587
rect 8428 -5663 8481 -5621
rect 8535 -5518 8588 -5499
rect 8535 -5552 8543 -5518
rect 8577 -5552 8588 -5518
rect 8535 -5586 8588 -5552
rect 8535 -5620 8543 -5586
rect 8577 -5620 8588 -5586
rect 8535 -5663 8588 -5620
rect 8688 -5518 8760 -5499
rect 8688 -5552 8701 -5518
rect 8735 -5552 8760 -5518
rect 8688 -5586 8760 -5552
rect 8688 -5620 8701 -5586
rect 8735 -5620 8760 -5586
rect 8688 -5663 8760 -5620
rect 8263 -5699 8313 -5663
rect 8710 -5699 8760 -5663
rect 8790 -5518 8844 -5499
rect 8990 -5511 9042 -5499
rect 8790 -5552 8801 -5518
rect 8835 -5552 8844 -5518
rect 8790 -5586 8844 -5552
rect 8790 -5620 8801 -5586
rect 8835 -5620 8844 -5586
rect 8790 -5699 8844 -5620
rect 8990 -5545 8998 -5511
rect 9032 -5545 9042 -5511
rect 8990 -5613 9042 -5545
rect 8990 -5647 8998 -5613
rect 9032 -5647 9042 -5613
rect 8990 -5673 9042 -5647
rect 9252 -5511 9304 -5499
rect 9252 -5545 9262 -5511
rect 9296 -5545 9304 -5511
rect 9450 -5511 9502 -5499
rect 9252 -5613 9304 -5545
rect 9252 -5647 9262 -5613
rect 9296 -5647 9304 -5613
rect 9252 -5673 9304 -5647
rect 9450 -5545 9458 -5511
rect 9492 -5545 9502 -5511
rect 9450 -5613 9502 -5545
rect 9450 -5647 9458 -5613
rect 9492 -5647 9502 -5613
rect 9450 -5673 9502 -5647
rect 10080 -5511 10132 -5499
rect 10080 -5545 10090 -5511
rect 10124 -5545 10132 -5511
rect 10370 -5511 10422 -5499
rect 10080 -5613 10132 -5545
rect 10080 -5647 10090 -5613
rect 10124 -5647 10132 -5613
rect 10080 -5673 10132 -5647
rect 10370 -5545 10378 -5511
rect 10412 -5545 10422 -5511
rect 10370 -5613 10422 -5545
rect 10370 -5647 10378 -5613
rect 10412 -5647 10422 -5613
rect 10370 -5673 10422 -5647
rect 10632 -5511 10684 -5499
rect 10632 -5545 10642 -5511
rect 10676 -5545 10684 -5511
rect 10632 -5613 10684 -5545
rect 10632 -5647 10642 -5613
rect 10676 -5647 10684 -5613
rect 10632 -5673 10684 -5647
rect 10738 -5519 10809 -5499
rect 10738 -5553 10761 -5519
rect 10795 -5553 10809 -5519
rect 10738 -5587 10809 -5553
rect 10738 -5621 10761 -5587
rect 10795 -5621 10809 -5587
rect 10738 -5699 10809 -5621
rect 10839 -5518 10904 -5499
rect 10839 -5552 10859 -5518
rect 10893 -5552 10904 -5518
rect 10839 -5586 10904 -5552
rect 10839 -5620 10859 -5586
rect 10893 -5620 10904 -5586
rect 10839 -5663 10904 -5620
rect 11004 -5519 11057 -5499
rect 11004 -5553 11015 -5519
rect 11049 -5553 11057 -5519
rect 11004 -5587 11057 -5553
rect 11004 -5621 11015 -5587
rect 11049 -5621 11057 -5587
rect 11004 -5663 11057 -5621
rect 11111 -5518 11164 -5499
rect 11111 -5552 11119 -5518
rect 11153 -5552 11164 -5518
rect 11111 -5586 11164 -5552
rect 11111 -5620 11119 -5586
rect 11153 -5620 11164 -5586
rect 11111 -5663 11164 -5620
rect 11264 -5518 11336 -5499
rect 11264 -5552 11277 -5518
rect 11311 -5552 11336 -5518
rect 11264 -5586 11336 -5552
rect 11264 -5620 11277 -5586
rect 11311 -5620 11336 -5586
rect 11264 -5663 11336 -5620
rect 10839 -5699 10889 -5663
rect 11286 -5699 11336 -5663
rect 11366 -5518 11420 -5499
rect 11658 -5511 11710 -5499
rect 11366 -5552 11377 -5518
rect 11411 -5552 11420 -5518
rect 11366 -5586 11420 -5552
rect 11366 -5620 11377 -5586
rect 11411 -5620 11420 -5586
rect 11366 -5699 11420 -5620
rect 11658 -5545 11666 -5511
rect 11700 -5545 11710 -5511
rect 11658 -5613 11710 -5545
rect 11658 -5647 11666 -5613
rect 11700 -5647 11710 -5613
rect 11658 -5673 11710 -5647
rect 11920 -5511 11972 -5499
rect 11920 -5545 11930 -5511
rect 11964 -5545 11972 -5511
rect 13682 -5511 13735 -5499
rect 11920 -5613 11972 -5545
rect 11920 -5647 11930 -5613
rect 11964 -5647 11972 -5613
rect 11920 -5673 11972 -5647
rect 13682 -5545 13690 -5511
rect 13724 -5545 13735 -5511
rect 13682 -5579 13735 -5545
rect 13682 -5613 13690 -5579
rect 13724 -5613 13735 -5579
rect 13682 -5699 13735 -5613
rect 13765 -5519 13821 -5499
rect 13765 -5553 13776 -5519
rect 13810 -5553 13821 -5519
rect 13765 -5587 13821 -5553
rect 13765 -5621 13776 -5587
rect 13810 -5621 13821 -5587
rect 13765 -5699 13821 -5621
rect 13851 -5511 13907 -5499
rect 13851 -5545 13862 -5511
rect 13896 -5545 13907 -5511
rect 13851 -5579 13907 -5545
rect 13851 -5613 13862 -5579
rect 13896 -5613 13907 -5579
rect 13851 -5699 13907 -5613
rect 13937 -5527 13993 -5499
rect 13937 -5561 13948 -5527
rect 13982 -5561 13993 -5527
rect 13937 -5595 13993 -5561
rect 13937 -5629 13948 -5595
rect 13982 -5629 13993 -5595
rect 13937 -5699 13993 -5629
rect 14023 -5511 14079 -5499
rect 14023 -5545 14034 -5511
rect 14068 -5545 14079 -5511
rect 14023 -5579 14079 -5545
rect 14023 -5613 14034 -5579
rect 14068 -5613 14079 -5579
rect 14023 -5699 14079 -5613
rect 14109 -5555 14165 -5499
rect 14109 -5589 14120 -5555
rect 14154 -5589 14165 -5555
rect 14109 -5641 14165 -5589
rect 14109 -5675 14120 -5641
rect 14154 -5675 14165 -5641
rect 14109 -5699 14165 -5675
rect 14195 -5535 14251 -5499
rect 14195 -5569 14206 -5535
rect 14240 -5569 14251 -5535
rect 14195 -5699 14251 -5569
rect 14281 -5555 14337 -5499
rect 14281 -5589 14292 -5555
rect 14326 -5589 14337 -5555
rect 14281 -5641 14337 -5589
rect 14281 -5675 14292 -5641
rect 14326 -5675 14337 -5641
rect 14281 -5699 14337 -5675
rect 14367 -5535 14423 -5499
rect 14367 -5569 14378 -5535
rect 14412 -5569 14423 -5535
rect 14367 -5699 14423 -5569
rect 14453 -5555 14509 -5499
rect 14453 -5589 14464 -5555
rect 14498 -5589 14509 -5555
rect 14453 -5641 14509 -5589
rect 14453 -5675 14464 -5641
rect 14498 -5675 14509 -5641
rect 14453 -5699 14509 -5675
rect 14539 -5535 14595 -5499
rect 14539 -5569 14550 -5535
rect 14584 -5569 14595 -5535
rect 14539 -5699 14595 -5569
rect 14625 -5555 14681 -5499
rect 14625 -5589 14636 -5555
rect 14670 -5589 14681 -5555
rect 14625 -5641 14681 -5589
rect 14625 -5675 14636 -5641
rect 14670 -5675 14681 -5641
rect 14625 -5699 14681 -5675
rect 14711 -5535 14766 -5499
rect 14711 -5569 14722 -5535
rect 14756 -5569 14766 -5535
rect 14711 -5699 14766 -5569
rect 14796 -5555 14852 -5499
rect 14796 -5589 14807 -5555
rect 14841 -5589 14852 -5555
rect 14796 -5641 14852 -5589
rect 14796 -5675 14807 -5641
rect 14841 -5675 14852 -5641
rect 14796 -5699 14852 -5675
rect 14882 -5535 14938 -5499
rect 14882 -5569 14893 -5535
rect 14927 -5569 14938 -5535
rect 14882 -5699 14938 -5569
rect 14968 -5555 15024 -5499
rect 14968 -5589 14979 -5555
rect 15013 -5589 15024 -5555
rect 14968 -5641 15024 -5589
rect 14968 -5675 14979 -5641
rect 15013 -5675 15024 -5641
rect 14968 -5699 15024 -5675
rect 15054 -5535 15110 -5499
rect 15054 -5569 15065 -5535
rect 15099 -5569 15110 -5535
rect 15054 -5699 15110 -5569
rect 15140 -5555 15196 -5499
rect 15140 -5589 15151 -5555
rect 15185 -5589 15196 -5555
rect 15140 -5641 15196 -5589
rect 15140 -5675 15151 -5641
rect 15185 -5675 15196 -5641
rect 15140 -5699 15196 -5675
rect 15226 -5535 15282 -5499
rect 15226 -5569 15237 -5535
rect 15271 -5569 15282 -5535
rect 15226 -5699 15282 -5569
rect 15312 -5555 15368 -5499
rect 15312 -5589 15323 -5555
rect 15357 -5589 15368 -5555
rect 15312 -5641 15368 -5589
rect 15312 -5675 15323 -5641
rect 15357 -5675 15368 -5641
rect 15312 -5699 15368 -5675
rect 15398 -5535 15451 -5499
rect 15614 -5511 15666 -5499
rect 15398 -5569 15409 -5535
rect 15443 -5569 15451 -5535
rect 15398 -5699 15451 -5569
rect 15614 -5545 15622 -5511
rect 15656 -5545 15666 -5511
rect 15614 -5613 15666 -5545
rect 15614 -5647 15622 -5613
rect 15656 -5647 15666 -5613
rect 15614 -5673 15666 -5647
rect 16612 -5511 16664 -5499
rect 16612 -5545 16622 -5511
rect 16656 -5545 16664 -5511
rect 16612 -5613 16664 -5545
rect 16612 -5647 16622 -5613
rect 16656 -5647 16664 -5613
rect 16612 -5673 16664 -5647
rect -2970 -6345 -2918 -6319
rect -2970 -6379 -2962 -6345
rect -2928 -6379 -2918 -6345
rect -2970 -6447 -2918 -6379
rect -2970 -6481 -2962 -6447
rect -2928 -6481 -2918 -6447
rect -2970 -6493 -2918 -6481
rect -2340 -6345 -2288 -6319
rect -2340 -6379 -2330 -6345
rect -2296 -6379 -2288 -6345
rect -2340 -6447 -2288 -6379
rect -2340 -6481 -2330 -6447
rect -2296 -6481 -2288 -6447
rect -1406 -6345 -1354 -6319
rect -1406 -6379 -1398 -6345
rect -1364 -6379 -1354 -6345
rect -1406 -6447 -1354 -6379
rect -2340 -6493 -2288 -6481
rect -1406 -6481 -1398 -6447
rect -1364 -6481 -1354 -6447
rect -1406 -6493 -1354 -6481
rect -1144 -6345 -1092 -6319
rect -1144 -6379 -1134 -6345
rect -1100 -6379 -1092 -6345
rect -1144 -6447 -1092 -6379
rect -1144 -6481 -1134 -6447
rect -1100 -6481 -1092 -6447
rect -942 -6311 -890 -6293
rect -942 -6345 -934 -6311
rect -900 -6345 -890 -6311
rect -942 -6379 -890 -6345
rect -942 -6413 -934 -6379
rect -900 -6413 -890 -6379
rect -942 -6447 -890 -6413
rect -1144 -6493 -1092 -6481
rect -942 -6481 -934 -6447
rect -900 -6481 -890 -6447
rect -942 -6493 -890 -6481
rect -860 -6311 -806 -6293
rect -860 -6345 -850 -6311
rect -816 -6345 -806 -6311
rect -860 -6379 -806 -6345
rect -860 -6413 -850 -6379
rect -816 -6413 -806 -6379
rect -860 -6447 -806 -6413
rect -860 -6481 -850 -6447
rect -816 -6481 -806 -6447
rect -860 -6493 -806 -6481
rect -776 -6311 -724 -6293
rect -776 -6345 -766 -6311
rect -732 -6345 -724 -6311
rect -776 -6379 -724 -6345
rect -776 -6413 -766 -6379
rect -732 -6413 -724 -6379
rect -776 -6447 -724 -6413
rect -776 -6481 -766 -6447
rect -732 -6481 -724 -6447
rect -578 -6345 -526 -6319
rect -578 -6379 -570 -6345
rect -536 -6379 -526 -6345
rect -578 -6447 -526 -6379
rect -776 -6493 -724 -6481
rect -578 -6481 -570 -6447
rect -536 -6481 -526 -6447
rect -578 -6493 -526 -6481
rect -316 -6345 -264 -6319
rect -316 -6379 -306 -6345
rect -272 -6379 -264 -6345
rect -316 -6447 -264 -6379
rect -316 -6481 -306 -6447
rect -272 -6481 -264 -6447
rect -118 -6372 -57 -6293
rect -118 -6406 -102 -6372
rect -68 -6406 -57 -6372
rect -118 -6440 -57 -6406
rect -118 -6474 -102 -6440
rect -68 -6474 -57 -6440
rect -316 -6493 -264 -6481
rect -118 -6493 -57 -6474
rect -27 -6345 29 -6293
rect -27 -6379 -16 -6345
rect 18 -6379 29 -6345
rect -27 -6433 29 -6379
rect -27 -6467 -16 -6433
rect 18 -6467 29 -6433
rect -27 -6493 29 -6467
rect 59 -6372 115 -6293
rect 59 -6406 70 -6372
rect 104 -6406 115 -6372
rect 59 -6440 115 -6406
rect 59 -6474 70 -6440
rect 104 -6474 115 -6440
rect 59 -6493 115 -6474
rect 145 -6345 201 -6293
rect 145 -6379 156 -6345
rect 190 -6379 201 -6345
rect 145 -6433 201 -6379
rect 145 -6467 156 -6433
rect 190 -6467 201 -6433
rect 145 -6493 201 -6467
rect 231 -6372 287 -6293
rect 231 -6406 242 -6372
rect 276 -6406 287 -6372
rect 231 -6440 287 -6406
rect 231 -6474 242 -6440
rect 276 -6474 287 -6440
rect 231 -6493 287 -6474
rect 317 -6345 373 -6293
rect 317 -6379 328 -6345
rect 362 -6379 373 -6345
rect 317 -6433 373 -6379
rect 317 -6467 328 -6433
rect 362 -6467 373 -6433
rect 317 -6493 373 -6467
rect 403 -6372 472 -6293
rect 403 -6406 414 -6372
rect 448 -6406 472 -6372
rect 403 -6440 472 -6406
rect 403 -6474 414 -6440
rect 448 -6474 472 -6440
rect 403 -6493 472 -6474
rect 618 -6345 670 -6319
rect 618 -6379 626 -6345
rect 660 -6379 670 -6345
rect 618 -6447 670 -6379
rect 618 -6481 626 -6447
rect 660 -6481 670 -6447
rect 618 -6493 670 -6481
rect 880 -6345 932 -6319
rect 880 -6379 890 -6345
rect 924 -6379 932 -6345
rect 880 -6447 932 -6379
rect 880 -6481 890 -6447
rect 924 -6481 932 -6447
rect 1078 -6345 1130 -6325
rect 1078 -6379 1086 -6345
rect 1120 -6379 1130 -6345
rect 1078 -6447 1130 -6379
rect 880 -6493 932 -6481
rect 1078 -6481 1086 -6447
rect 1120 -6481 1130 -6447
rect 1078 -6493 1130 -6481
rect 1160 -6345 1214 -6325
rect 1160 -6379 1170 -6345
rect 1204 -6379 1214 -6345
rect 1160 -6447 1214 -6379
rect 1160 -6481 1170 -6447
rect 1204 -6481 1214 -6447
rect 1160 -6493 1214 -6481
rect 1244 -6345 1300 -6325
rect 1244 -6379 1254 -6345
rect 1288 -6379 1300 -6345
rect 1244 -6447 1300 -6379
rect 1244 -6481 1254 -6447
rect 1288 -6481 1300 -6447
rect 1446 -6345 1498 -6319
rect 1446 -6379 1454 -6345
rect 1488 -6379 1498 -6345
rect 1446 -6447 1498 -6379
rect 1244 -6493 1300 -6481
rect 1446 -6481 1454 -6447
rect 1488 -6481 1498 -6447
rect 1446 -6493 1498 -6481
rect 1708 -6345 1760 -6319
rect 1708 -6379 1718 -6345
rect 1752 -6379 1760 -6345
rect 1708 -6447 1760 -6379
rect 1708 -6481 1718 -6447
rect 1752 -6481 1760 -6447
rect 1906 -6345 1958 -6319
rect 1906 -6379 1914 -6345
rect 1948 -6379 1958 -6345
rect 1906 -6447 1958 -6379
rect 1708 -6493 1760 -6481
rect 1906 -6481 1914 -6447
rect 1948 -6481 1958 -6447
rect 1906 -6493 1958 -6481
rect 2168 -6345 2220 -6319
rect 2168 -6379 2178 -6345
rect 2212 -6379 2220 -6345
rect 2168 -6447 2220 -6379
rect 2168 -6481 2178 -6447
rect 2212 -6481 2220 -6447
rect 2366 -6372 2420 -6293
rect 2366 -6406 2375 -6372
rect 2409 -6406 2420 -6372
rect 2366 -6440 2420 -6406
rect 2366 -6474 2375 -6440
rect 2409 -6474 2420 -6440
rect 2168 -6493 2220 -6481
rect 2366 -6493 2420 -6474
rect 2450 -6329 2500 -6293
rect 2897 -6329 2947 -6293
rect 2450 -6372 2522 -6329
rect 2450 -6406 2475 -6372
rect 2509 -6406 2522 -6372
rect 2450 -6440 2522 -6406
rect 2450 -6474 2475 -6440
rect 2509 -6474 2522 -6440
rect 2450 -6493 2522 -6474
rect 2622 -6372 2675 -6329
rect 2622 -6406 2633 -6372
rect 2667 -6406 2675 -6372
rect 2622 -6440 2675 -6406
rect 2622 -6474 2633 -6440
rect 2667 -6474 2675 -6440
rect 2622 -6493 2675 -6474
rect 2729 -6371 2782 -6329
rect 2729 -6405 2737 -6371
rect 2771 -6405 2782 -6371
rect 2729 -6439 2782 -6405
rect 2729 -6473 2737 -6439
rect 2771 -6473 2782 -6439
rect 2729 -6493 2782 -6473
rect 2882 -6372 2947 -6329
rect 2882 -6406 2893 -6372
rect 2927 -6406 2947 -6372
rect 2882 -6440 2947 -6406
rect 2882 -6474 2893 -6440
rect 2927 -6474 2947 -6440
rect 2882 -6493 2947 -6474
rect 2977 -6371 3048 -6293
rect 2977 -6405 2991 -6371
rect 3025 -6405 3048 -6371
rect 2977 -6439 3048 -6405
rect 2977 -6473 2991 -6439
rect 3025 -6473 3048 -6439
rect 2977 -6493 3048 -6473
rect 3194 -6345 3246 -6319
rect 3194 -6379 3202 -6345
rect 3236 -6379 3246 -6345
rect 3194 -6447 3246 -6379
rect 3194 -6481 3202 -6447
rect 3236 -6481 3246 -6447
rect 3194 -6493 3246 -6481
rect 3456 -6345 3508 -6319
rect 3456 -6379 3466 -6345
rect 3500 -6379 3508 -6345
rect 3456 -6447 3508 -6379
rect 3456 -6481 3466 -6447
rect 3500 -6481 3508 -6447
rect 4390 -6345 4442 -6319
rect 4390 -6379 4398 -6345
rect 4432 -6379 4442 -6345
rect 4390 -6447 4442 -6379
rect 3456 -6493 3508 -6481
rect 4390 -6481 4398 -6447
rect 4432 -6481 4442 -6447
rect 4390 -6493 4442 -6481
rect 5388 -6345 5440 -6319
rect 5388 -6379 5398 -6345
rect 5432 -6379 5440 -6345
rect 5388 -6447 5440 -6379
rect 5388 -6481 5398 -6447
rect 5432 -6481 5440 -6447
rect 6414 -6345 6466 -6319
rect 6414 -6379 6422 -6345
rect 6456 -6379 6466 -6345
rect 6414 -6447 6466 -6379
rect 5388 -6493 5440 -6481
rect 6414 -6481 6422 -6447
rect 6456 -6481 6466 -6447
rect 6414 -6493 6466 -6481
rect 6676 -6345 6728 -6319
rect 6676 -6379 6686 -6345
rect 6720 -6379 6728 -6345
rect 6676 -6447 6728 -6379
rect 6676 -6481 6686 -6447
rect 6720 -6481 6728 -6447
rect 6874 -6372 6928 -6293
rect 6874 -6406 6883 -6372
rect 6917 -6406 6928 -6372
rect 6874 -6440 6928 -6406
rect 6874 -6474 6883 -6440
rect 6917 -6474 6928 -6440
rect 6676 -6493 6728 -6481
rect 6874 -6493 6928 -6474
rect 6958 -6329 7008 -6293
rect 7405 -6329 7455 -6293
rect 6958 -6372 7030 -6329
rect 6958 -6406 6983 -6372
rect 7017 -6406 7030 -6372
rect 6958 -6440 7030 -6406
rect 6958 -6474 6983 -6440
rect 7017 -6474 7030 -6440
rect 6958 -6493 7030 -6474
rect 7130 -6372 7183 -6329
rect 7130 -6406 7141 -6372
rect 7175 -6406 7183 -6372
rect 7130 -6440 7183 -6406
rect 7130 -6474 7141 -6440
rect 7175 -6474 7183 -6440
rect 7130 -6493 7183 -6474
rect 7237 -6371 7290 -6329
rect 7237 -6405 7245 -6371
rect 7279 -6405 7290 -6371
rect 7237 -6439 7290 -6405
rect 7237 -6473 7245 -6439
rect 7279 -6473 7290 -6439
rect 7237 -6493 7290 -6473
rect 7390 -6372 7455 -6329
rect 7390 -6406 7401 -6372
rect 7435 -6406 7455 -6372
rect 7390 -6440 7455 -6406
rect 7390 -6474 7401 -6440
rect 7435 -6474 7455 -6440
rect 7390 -6493 7455 -6474
rect 7485 -6371 7556 -6293
rect 7485 -6405 7499 -6371
rect 7533 -6405 7556 -6371
rect 7485 -6439 7556 -6405
rect 7485 -6473 7499 -6439
rect 7533 -6473 7556 -6439
rect 7485 -6493 7556 -6473
rect 7702 -6345 7754 -6319
rect 7702 -6379 7710 -6345
rect 7744 -6379 7754 -6345
rect 7702 -6447 7754 -6379
rect 7702 -6481 7710 -6447
rect 7744 -6481 7754 -6447
rect 7702 -6493 7754 -6481
rect 7964 -6345 8016 -6319
rect 7964 -6379 7974 -6345
rect 8008 -6379 8016 -6345
rect 7964 -6447 8016 -6379
rect 7964 -6481 7974 -6447
rect 8008 -6481 8016 -6447
rect 8162 -6372 8216 -6293
rect 8162 -6406 8171 -6372
rect 8205 -6406 8216 -6372
rect 8162 -6440 8216 -6406
rect 8162 -6474 8171 -6440
rect 8205 -6474 8216 -6440
rect 7964 -6493 8016 -6481
rect 8162 -6493 8216 -6474
rect 8246 -6329 8296 -6293
rect 8693 -6329 8743 -6293
rect 8246 -6372 8318 -6329
rect 8246 -6406 8271 -6372
rect 8305 -6406 8318 -6372
rect 8246 -6440 8318 -6406
rect 8246 -6474 8271 -6440
rect 8305 -6474 8318 -6440
rect 8246 -6493 8318 -6474
rect 8418 -6372 8471 -6329
rect 8418 -6406 8429 -6372
rect 8463 -6406 8471 -6372
rect 8418 -6440 8471 -6406
rect 8418 -6474 8429 -6440
rect 8463 -6474 8471 -6440
rect 8418 -6493 8471 -6474
rect 8525 -6371 8578 -6329
rect 8525 -6405 8533 -6371
rect 8567 -6405 8578 -6371
rect 8525 -6439 8578 -6405
rect 8525 -6473 8533 -6439
rect 8567 -6473 8578 -6439
rect 8525 -6493 8578 -6473
rect 8678 -6372 8743 -6329
rect 8678 -6406 8689 -6372
rect 8723 -6406 8743 -6372
rect 8678 -6440 8743 -6406
rect 8678 -6474 8689 -6440
rect 8723 -6474 8743 -6440
rect 8678 -6493 8743 -6474
rect 8773 -6371 8844 -6293
rect 8773 -6405 8787 -6371
rect 8821 -6405 8844 -6371
rect 8773 -6439 8844 -6405
rect 8773 -6473 8787 -6439
rect 8821 -6473 8844 -6439
rect 8773 -6493 8844 -6473
rect 8990 -6345 9042 -6319
rect 8990 -6379 8998 -6345
rect 9032 -6379 9042 -6345
rect 8990 -6447 9042 -6379
rect 8990 -6481 8998 -6447
rect 9032 -6481 9042 -6447
rect 8990 -6493 9042 -6481
rect 9252 -6345 9304 -6319
rect 9252 -6379 9262 -6345
rect 9296 -6379 9304 -6345
rect 9252 -6447 9304 -6379
rect 9252 -6481 9262 -6447
rect 9296 -6481 9304 -6447
rect 9450 -6372 9504 -6293
rect 9450 -6406 9459 -6372
rect 9493 -6406 9504 -6372
rect 9450 -6440 9504 -6406
rect 9450 -6474 9459 -6440
rect 9493 -6474 9504 -6440
rect 9252 -6493 9304 -6481
rect 9450 -6493 9504 -6474
rect 9534 -6329 9584 -6293
rect 9981 -6329 10031 -6293
rect 9534 -6372 9606 -6329
rect 9534 -6406 9559 -6372
rect 9593 -6406 9606 -6372
rect 9534 -6440 9606 -6406
rect 9534 -6474 9559 -6440
rect 9593 -6474 9606 -6440
rect 9534 -6493 9606 -6474
rect 9706 -6372 9759 -6329
rect 9706 -6406 9717 -6372
rect 9751 -6406 9759 -6372
rect 9706 -6440 9759 -6406
rect 9706 -6474 9717 -6440
rect 9751 -6474 9759 -6440
rect 9706 -6493 9759 -6474
rect 9813 -6371 9866 -6329
rect 9813 -6405 9821 -6371
rect 9855 -6405 9866 -6371
rect 9813 -6439 9866 -6405
rect 9813 -6473 9821 -6439
rect 9855 -6473 9866 -6439
rect 9813 -6493 9866 -6473
rect 9966 -6372 10031 -6329
rect 9966 -6406 9977 -6372
rect 10011 -6406 10031 -6372
rect 9966 -6440 10031 -6406
rect 9966 -6474 9977 -6440
rect 10011 -6474 10031 -6440
rect 9966 -6493 10031 -6474
rect 10061 -6371 10132 -6293
rect 10061 -6405 10075 -6371
rect 10109 -6405 10132 -6371
rect 10061 -6439 10132 -6405
rect 10061 -6473 10075 -6439
rect 10109 -6473 10132 -6439
rect 10061 -6493 10132 -6473
rect 10278 -6345 10330 -6319
rect 10278 -6379 10286 -6345
rect 10320 -6379 10330 -6345
rect 10278 -6447 10330 -6379
rect 10278 -6481 10286 -6447
rect 10320 -6481 10330 -6447
rect 10278 -6493 10330 -6481
rect 10540 -6345 10592 -6319
rect 10540 -6379 10550 -6345
rect 10584 -6379 10592 -6345
rect 10540 -6447 10592 -6379
rect 10540 -6481 10550 -6447
rect 10584 -6481 10592 -6447
rect 10738 -6311 10790 -6293
rect 10738 -6345 10746 -6311
rect 10780 -6345 10790 -6311
rect 10738 -6379 10790 -6345
rect 10738 -6413 10746 -6379
rect 10780 -6413 10790 -6379
rect 10738 -6447 10790 -6413
rect 10540 -6493 10592 -6481
rect 10738 -6481 10746 -6447
rect 10780 -6481 10790 -6447
rect 10738 -6493 10790 -6481
rect 10820 -6311 10874 -6293
rect 10820 -6345 10830 -6311
rect 10864 -6345 10874 -6311
rect 10820 -6379 10874 -6345
rect 10820 -6413 10830 -6379
rect 10864 -6413 10874 -6379
rect 10820 -6447 10874 -6413
rect 10820 -6481 10830 -6447
rect 10864 -6481 10874 -6447
rect 10820 -6493 10874 -6481
rect 10904 -6379 10958 -6293
rect 10904 -6413 10914 -6379
rect 10948 -6413 10958 -6379
rect 10904 -6447 10958 -6413
rect 10904 -6481 10914 -6447
rect 10948 -6481 10958 -6447
rect 10904 -6493 10958 -6481
rect 10988 -6311 11042 -6293
rect 10988 -6345 10998 -6311
rect 11032 -6345 11042 -6311
rect 10988 -6379 11042 -6345
rect 10988 -6413 10998 -6379
rect 11032 -6413 11042 -6379
rect 10988 -6447 11042 -6413
rect 10988 -6481 10998 -6447
rect 11032 -6481 11042 -6447
rect 10988 -6493 11042 -6481
rect 11072 -6379 11126 -6293
rect 11072 -6413 11082 -6379
rect 11116 -6413 11126 -6379
rect 11072 -6447 11126 -6413
rect 11072 -6481 11082 -6447
rect 11116 -6481 11126 -6447
rect 11072 -6493 11126 -6481
rect 11156 -6311 11210 -6293
rect 11156 -6345 11166 -6311
rect 11200 -6345 11210 -6311
rect 11156 -6379 11210 -6345
rect 11156 -6413 11166 -6379
rect 11200 -6413 11210 -6379
rect 11156 -6447 11210 -6413
rect 11156 -6481 11166 -6447
rect 11200 -6481 11210 -6447
rect 11156 -6493 11210 -6481
rect 11240 -6379 11294 -6293
rect 11240 -6413 11250 -6379
rect 11284 -6413 11294 -6379
rect 11240 -6447 11294 -6413
rect 11240 -6481 11250 -6447
rect 11284 -6481 11294 -6447
rect 11240 -6493 11294 -6481
rect 11324 -6311 11378 -6293
rect 11324 -6345 11334 -6311
rect 11368 -6345 11378 -6311
rect 11324 -6379 11378 -6345
rect 11324 -6413 11334 -6379
rect 11368 -6413 11378 -6379
rect 11324 -6447 11378 -6413
rect 11324 -6481 11334 -6447
rect 11368 -6481 11378 -6447
rect 11324 -6493 11378 -6481
rect 11408 -6379 11460 -6293
rect 11408 -6413 11418 -6379
rect 11452 -6413 11460 -6379
rect 11408 -6447 11460 -6413
rect 11408 -6481 11418 -6447
rect 11452 -6481 11460 -6447
rect 11658 -6345 11710 -6319
rect 11658 -6379 11666 -6345
rect 11700 -6379 11710 -6345
rect 11658 -6447 11710 -6379
rect 11408 -6493 11460 -6481
rect 11658 -6481 11666 -6447
rect 11700 -6481 11710 -6447
rect 11658 -6493 11710 -6481
rect 11920 -6345 11972 -6319
rect 11920 -6379 11930 -6345
rect 11964 -6379 11972 -6345
rect 11920 -6447 11972 -6379
rect 11920 -6481 11930 -6447
rect 11964 -6481 11972 -6447
rect 13590 -6345 13642 -6319
rect 13590 -6379 13598 -6345
rect 13632 -6379 13642 -6345
rect 13590 -6447 13642 -6379
rect 11920 -6493 11972 -6481
rect 13590 -6481 13598 -6447
rect 13632 -6481 13642 -6447
rect 13590 -6493 13642 -6481
rect 14588 -6345 14640 -6319
rect 14588 -6379 14598 -6345
rect 14632 -6379 14640 -6345
rect 14588 -6447 14640 -6379
rect 14588 -6481 14598 -6447
rect 14632 -6481 14640 -6447
rect 14786 -6345 14838 -6319
rect 14786 -6379 14794 -6345
rect 14828 -6379 14838 -6345
rect 14786 -6447 14838 -6379
rect 14588 -6493 14640 -6481
rect 14786 -6481 14794 -6447
rect 14828 -6481 14838 -6447
rect 14786 -6493 14838 -6481
rect 15784 -6345 15836 -6319
rect 15784 -6379 15794 -6345
rect 15828 -6379 15836 -6345
rect 15784 -6447 15836 -6379
rect 15784 -6481 15794 -6447
rect 15828 -6481 15836 -6447
rect 15982 -6345 16034 -6319
rect 15982 -6379 15990 -6345
rect 16024 -6379 16034 -6345
rect 15982 -6447 16034 -6379
rect 15784 -6493 15836 -6481
rect 15982 -6481 15990 -6447
rect 16024 -6481 16034 -6447
rect 15982 -6493 16034 -6481
rect 16612 -6345 16664 -6319
rect 16612 -6379 16622 -6345
rect 16656 -6379 16664 -6345
rect 16612 -6447 16664 -6379
rect 16612 -6481 16622 -6447
rect 16656 -6481 16664 -6447
rect 16612 -6493 16664 -6481
rect -2970 -6599 -2918 -6587
rect -2970 -6633 -2962 -6599
rect -2928 -6633 -2918 -6599
rect -2970 -6694 -2918 -6633
rect -2970 -6728 -2962 -6694
rect -2928 -6728 -2918 -6694
rect -2970 -6761 -2918 -6728
rect -2800 -6599 -2748 -6587
rect -2800 -6633 -2790 -6599
rect -2756 -6633 -2748 -6599
rect -2800 -6694 -2748 -6633
rect -2800 -6728 -2790 -6694
rect -2756 -6728 -2748 -6694
rect -2800 -6761 -2748 -6728
rect -2602 -6607 -2550 -6593
rect -2602 -6641 -2594 -6607
rect -2560 -6641 -2550 -6607
rect -2602 -6675 -2550 -6641
rect -2602 -6709 -2594 -6675
rect -2560 -6709 -2550 -6675
rect -2602 -6721 -2550 -6709
rect -2520 -6623 -2466 -6593
rect -2520 -6657 -2510 -6623
rect -2476 -6657 -2466 -6623
rect -2520 -6721 -2466 -6657
rect -2436 -6607 -2384 -6593
rect -2436 -6641 -2426 -6607
rect -2392 -6641 -2384 -6607
rect -2436 -6675 -2384 -6641
rect -2330 -6599 -2278 -6587
rect -2330 -6633 -2322 -6599
rect -2288 -6633 -2278 -6599
rect -2330 -6671 -2278 -6633
rect -2248 -6607 -2193 -6587
rect -2248 -6641 -2238 -6607
rect -2204 -6641 -2193 -6607
rect -2248 -6671 -2193 -6641
rect -2163 -6612 -2098 -6587
rect -2163 -6646 -2146 -6612
rect -2112 -6646 -2098 -6612
rect -2163 -6671 -2098 -6646
rect -2068 -6671 -1995 -6587
rect -1965 -6599 -1863 -6587
rect -1965 -6633 -1907 -6599
rect -1873 -6633 -1863 -6599
rect -1965 -6667 -1863 -6633
rect -1965 -6671 -1907 -6667
rect -2436 -6709 -2426 -6675
rect -2392 -6709 -2384 -6675
rect -2436 -6721 -2384 -6709
rect -1950 -6701 -1907 -6671
rect -1873 -6701 -1863 -6667
rect -1950 -6737 -1863 -6701
rect -1833 -6607 -1768 -6587
rect -1833 -6641 -1823 -6607
rect -1789 -6641 -1768 -6607
rect -1833 -6671 -1768 -6641
rect -1738 -6617 -1684 -6587
rect -1738 -6651 -1728 -6617
rect -1694 -6651 -1684 -6617
rect -1738 -6671 -1684 -6651
rect -1654 -6671 -1570 -6587
rect -1540 -6607 -1487 -6587
rect -1540 -6641 -1529 -6607
rect -1495 -6641 -1487 -6607
rect -1540 -6671 -1487 -6641
rect -1413 -6599 -1359 -6587
rect -1413 -6633 -1405 -6599
rect -1371 -6633 -1359 -6599
rect -1413 -6670 -1359 -6633
rect -1833 -6737 -1783 -6671
rect -1413 -6704 -1405 -6670
rect -1371 -6704 -1359 -6670
rect -1413 -6741 -1359 -6704
rect -1413 -6775 -1405 -6741
rect -1371 -6775 -1359 -6741
rect -1413 -6787 -1359 -6775
rect -1329 -6629 -1275 -6587
rect -1329 -6663 -1319 -6629
rect -1285 -6663 -1275 -6629
rect -1329 -6709 -1275 -6663
rect -1329 -6743 -1319 -6709
rect -1285 -6743 -1275 -6709
rect -1329 -6787 -1275 -6743
rect -1245 -6605 -1193 -6587
rect -1245 -6639 -1235 -6605
rect -1201 -6639 -1193 -6605
rect -1245 -6673 -1193 -6639
rect -1245 -6707 -1235 -6673
rect -1201 -6707 -1193 -6673
rect -1245 -6741 -1193 -6707
rect -1139 -6599 -1087 -6587
rect -1139 -6633 -1131 -6599
rect -1097 -6633 -1087 -6599
rect -1139 -6667 -1087 -6633
rect -1139 -6701 -1131 -6667
rect -1097 -6701 -1087 -6667
rect -1139 -6715 -1087 -6701
rect -1057 -6599 -990 -6587
rect -1057 -6633 -1034 -6599
rect -1000 -6633 -990 -6599
rect -1057 -6667 -990 -6633
rect -1057 -6701 -1034 -6667
rect -1000 -6701 -990 -6667
rect -1057 -6715 -990 -6701
rect -1245 -6775 -1235 -6741
rect -1201 -6775 -1193 -6741
rect -1245 -6787 -1193 -6775
rect -1042 -6735 -990 -6715
rect -1042 -6769 -1034 -6735
rect -1000 -6769 -990 -6735
rect -1042 -6787 -990 -6769
rect -960 -6599 -908 -6587
rect -960 -6633 -950 -6599
rect -916 -6633 -908 -6599
rect -960 -6670 -908 -6633
rect -960 -6704 -950 -6670
rect -916 -6704 -908 -6670
rect -960 -6741 -908 -6704
rect -960 -6775 -950 -6741
rect -916 -6775 -908 -6741
rect -854 -6599 -802 -6587
rect -854 -6633 -846 -6599
rect -812 -6633 -802 -6599
rect -854 -6701 -802 -6633
rect -854 -6735 -846 -6701
rect -812 -6735 -802 -6701
rect -854 -6761 -802 -6735
rect -224 -6599 -172 -6587
rect -224 -6633 -214 -6599
rect -180 -6633 -172 -6599
rect -26 -6599 26 -6587
rect -224 -6701 -172 -6633
rect -224 -6735 -214 -6701
rect -180 -6735 -172 -6701
rect -224 -6761 -172 -6735
rect -960 -6787 -908 -6775
rect -26 -6633 -18 -6599
rect 16 -6633 26 -6599
rect -26 -6701 26 -6633
rect -26 -6735 -18 -6701
rect 16 -6735 26 -6701
rect -26 -6761 26 -6735
rect 604 -6599 656 -6587
rect 604 -6633 614 -6599
rect 648 -6633 656 -6599
rect 604 -6701 656 -6633
rect 604 -6735 614 -6701
rect 648 -6735 656 -6701
rect 604 -6761 656 -6735
rect 710 -6599 762 -6587
rect 710 -6633 718 -6599
rect 752 -6633 762 -6599
rect 710 -6701 762 -6633
rect 710 -6735 718 -6701
rect 752 -6735 762 -6701
rect 710 -6761 762 -6735
rect 1340 -6599 1392 -6587
rect 1340 -6633 1350 -6599
rect 1384 -6633 1392 -6599
rect 1538 -6599 1590 -6587
rect 1340 -6701 1392 -6633
rect 1340 -6735 1350 -6701
rect 1384 -6735 1392 -6701
rect 1340 -6761 1392 -6735
rect 1538 -6633 1546 -6599
rect 1580 -6633 1590 -6599
rect 1538 -6701 1590 -6633
rect 1538 -6735 1546 -6701
rect 1580 -6735 1590 -6701
rect 1538 -6761 1590 -6735
rect 2168 -6599 2220 -6587
rect 2168 -6633 2178 -6599
rect 2212 -6633 2220 -6599
rect 2168 -6701 2220 -6633
rect 2168 -6735 2178 -6701
rect 2212 -6735 2220 -6701
rect 2168 -6761 2220 -6735
rect 2274 -6599 2326 -6587
rect 2274 -6633 2282 -6599
rect 2316 -6633 2326 -6599
rect 2274 -6701 2326 -6633
rect 2274 -6735 2282 -6701
rect 2316 -6735 2326 -6701
rect 2274 -6761 2326 -6735
rect 2904 -6599 2956 -6587
rect 2904 -6633 2914 -6599
rect 2948 -6633 2956 -6599
rect 3102 -6599 3154 -6587
rect 2904 -6701 2956 -6633
rect 2904 -6735 2914 -6701
rect 2948 -6735 2956 -6701
rect 2904 -6761 2956 -6735
rect 3102 -6633 3110 -6599
rect 3144 -6633 3154 -6599
rect 3102 -6701 3154 -6633
rect 3102 -6735 3110 -6701
rect 3144 -6735 3154 -6701
rect 3102 -6761 3154 -6735
rect 3732 -6599 3784 -6587
rect 3732 -6633 3742 -6599
rect 3776 -6633 3784 -6599
rect 3732 -6701 3784 -6633
rect 3732 -6735 3742 -6701
rect 3776 -6735 3784 -6701
rect 3732 -6761 3784 -6735
rect 3838 -6599 3890 -6587
rect 3838 -6633 3846 -6599
rect 3880 -6633 3890 -6599
rect 3838 -6701 3890 -6633
rect 3838 -6735 3846 -6701
rect 3880 -6735 3890 -6701
rect 3838 -6761 3890 -6735
rect 4468 -6599 4520 -6587
rect 4468 -6633 4478 -6599
rect 4512 -6633 4520 -6599
rect 4666 -6599 4718 -6587
rect 4468 -6701 4520 -6633
rect 4468 -6735 4478 -6701
rect 4512 -6735 4520 -6701
rect 4468 -6761 4520 -6735
rect 4666 -6633 4674 -6599
rect 4708 -6633 4718 -6599
rect 4666 -6701 4718 -6633
rect 4666 -6735 4674 -6701
rect 4708 -6735 4718 -6701
rect 4666 -6761 4718 -6735
rect 5296 -6599 5348 -6587
rect 5296 -6633 5306 -6599
rect 5340 -6633 5348 -6599
rect 5296 -6701 5348 -6633
rect 5296 -6735 5306 -6701
rect 5340 -6735 5348 -6701
rect 5296 -6761 5348 -6735
rect 5402 -6599 5454 -6587
rect 5402 -6633 5410 -6599
rect 5444 -6633 5454 -6599
rect 5402 -6701 5454 -6633
rect 5402 -6735 5410 -6701
rect 5444 -6735 5454 -6701
rect 5402 -6761 5454 -6735
rect 6032 -6599 6084 -6587
rect 6032 -6633 6042 -6599
rect 6076 -6633 6084 -6599
rect 6230 -6599 6282 -6587
rect 6032 -6701 6084 -6633
rect 6032 -6735 6042 -6701
rect 6076 -6735 6084 -6701
rect 6032 -6761 6084 -6735
rect 6230 -6633 6238 -6599
rect 6272 -6633 6282 -6599
rect 6230 -6701 6282 -6633
rect 6230 -6735 6238 -6701
rect 6272 -6735 6282 -6701
rect 6230 -6761 6282 -6735
rect 6860 -6599 6912 -6587
rect 6860 -6633 6870 -6599
rect 6904 -6633 6912 -6599
rect 6860 -6701 6912 -6633
rect 6860 -6735 6870 -6701
rect 6904 -6735 6912 -6701
rect 6860 -6761 6912 -6735
rect 6966 -6599 7018 -6587
rect 6966 -6633 6974 -6599
rect 7008 -6633 7018 -6599
rect 6966 -6701 7018 -6633
rect 6966 -6735 6974 -6701
rect 7008 -6735 7018 -6701
rect 6966 -6761 7018 -6735
rect 7596 -6599 7648 -6587
rect 7596 -6633 7606 -6599
rect 7640 -6633 7648 -6599
rect 7794 -6599 7846 -6587
rect 7596 -6701 7648 -6633
rect 7596 -6735 7606 -6701
rect 7640 -6735 7648 -6701
rect 7596 -6761 7648 -6735
rect 7794 -6633 7802 -6599
rect 7836 -6633 7846 -6599
rect 7794 -6701 7846 -6633
rect 7794 -6735 7802 -6701
rect 7836 -6735 7846 -6701
rect 7794 -6761 7846 -6735
rect 8424 -6599 8476 -6587
rect 8424 -6633 8434 -6599
rect 8468 -6633 8476 -6599
rect 8424 -6701 8476 -6633
rect 8424 -6735 8434 -6701
rect 8468 -6735 8476 -6701
rect 8424 -6761 8476 -6735
rect 8530 -6599 8582 -6587
rect 8530 -6633 8538 -6599
rect 8572 -6633 8582 -6599
rect 8530 -6701 8582 -6633
rect 8530 -6735 8538 -6701
rect 8572 -6735 8582 -6701
rect 8530 -6761 8582 -6735
rect 9160 -6599 9212 -6587
rect 9160 -6633 9170 -6599
rect 9204 -6633 9212 -6599
rect 15982 -6599 16034 -6587
rect 9160 -6701 9212 -6633
rect 9160 -6735 9170 -6701
rect 9204 -6735 9212 -6701
rect 9160 -6761 9212 -6735
rect 15982 -6633 15990 -6599
rect 16024 -6633 16034 -6599
rect 15982 -6701 16034 -6633
rect 15982 -6735 15990 -6701
rect 16024 -6735 16034 -6701
rect 15982 -6761 16034 -6735
rect 16612 -6599 16664 -6587
rect 16612 -6633 16622 -6599
rect 16656 -6633 16664 -6599
rect 16612 -6701 16664 -6633
rect 16612 -6735 16622 -6701
rect 16656 -6735 16664 -6701
rect 16612 -6761 16664 -6735
rect -2970 -7433 -2918 -7407
rect -2970 -7467 -2962 -7433
rect -2928 -7467 -2918 -7433
rect -2970 -7535 -2918 -7467
rect -2970 -7569 -2962 -7535
rect -2928 -7569 -2918 -7535
rect -2970 -7581 -2918 -7569
rect -2340 -7433 -2288 -7407
rect -2340 -7467 -2330 -7433
rect -2296 -7467 -2288 -7433
rect -2340 -7535 -2288 -7467
rect -2340 -7569 -2330 -7535
rect -2296 -7569 -2288 -7535
rect -1590 -7433 -1538 -7407
rect -1590 -7467 -1582 -7433
rect -1548 -7467 -1538 -7433
rect -1590 -7535 -1538 -7467
rect -2340 -7581 -2288 -7569
rect -1590 -7569 -1582 -7535
rect -1548 -7569 -1538 -7535
rect -1590 -7581 -1538 -7569
rect -960 -7433 -908 -7407
rect -960 -7467 -950 -7433
rect -916 -7467 -908 -7433
rect -960 -7535 -908 -7467
rect -960 -7569 -950 -7535
rect -916 -7569 -908 -7535
rect -960 -7581 -908 -7569
rect -854 -7433 -802 -7407
rect -854 -7467 -846 -7433
rect -812 -7467 -802 -7433
rect -854 -7535 -802 -7467
rect -854 -7569 -846 -7535
rect -812 -7569 -802 -7535
rect -854 -7581 -802 -7569
rect -224 -7433 -172 -7407
rect -224 -7467 -214 -7433
rect -180 -7467 -172 -7433
rect -224 -7535 -172 -7467
rect -224 -7569 -214 -7535
rect -180 -7569 -172 -7535
rect -26 -7433 26 -7407
rect -26 -7467 -18 -7433
rect 16 -7467 26 -7433
rect -26 -7535 26 -7467
rect -224 -7581 -172 -7569
rect -26 -7569 -18 -7535
rect 16 -7569 26 -7535
rect -26 -7581 26 -7569
rect 604 -7433 656 -7407
rect 604 -7467 614 -7433
rect 648 -7467 656 -7433
rect 604 -7535 656 -7467
rect 604 -7569 614 -7535
rect 648 -7569 656 -7535
rect 604 -7581 656 -7569
rect 710 -7433 762 -7407
rect 710 -7467 718 -7433
rect 752 -7467 762 -7433
rect 710 -7535 762 -7467
rect 710 -7569 718 -7535
rect 752 -7569 762 -7535
rect 710 -7581 762 -7569
rect 1340 -7433 1392 -7407
rect 1340 -7467 1350 -7433
rect 1384 -7467 1392 -7433
rect 1340 -7535 1392 -7467
rect 1340 -7569 1350 -7535
rect 1384 -7569 1392 -7535
rect 1538 -7433 1590 -7407
rect 1538 -7467 1546 -7433
rect 1580 -7467 1590 -7433
rect 1538 -7535 1590 -7467
rect 1340 -7581 1392 -7569
rect 1538 -7569 1546 -7535
rect 1580 -7569 1590 -7535
rect 1538 -7581 1590 -7569
rect 2168 -7433 2220 -7407
rect 2168 -7467 2178 -7433
rect 2212 -7467 2220 -7433
rect 2168 -7535 2220 -7467
rect 2168 -7569 2178 -7535
rect 2212 -7569 2220 -7535
rect 2168 -7581 2220 -7569
rect 2274 -7433 2326 -7407
rect 2274 -7467 2282 -7433
rect 2316 -7467 2326 -7433
rect 2274 -7535 2326 -7467
rect 2274 -7569 2282 -7535
rect 2316 -7569 2326 -7535
rect 2274 -7581 2326 -7569
rect 2536 -7433 2588 -7407
rect 2536 -7467 2546 -7433
rect 2580 -7467 2588 -7433
rect 2536 -7535 2588 -7467
rect 2536 -7569 2546 -7535
rect 2580 -7569 2588 -7535
rect 2918 -7433 2974 -7413
rect 2918 -7467 2930 -7433
rect 2964 -7467 2974 -7433
rect 2918 -7535 2974 -7467
rect 2536 -7581 2588 -7569
rect 2918 -7569 2930 -7535
rect 2964 -7569 2974 -7535
rect 2918 -7581 2974 -7569
rect 3004 -7433 3058 -7413
rect 3004 -7467 3014 -7433
rect 3048 -7467 3058 -7433
rect 3004 -7535 3058 -7467
rect 3004 -7569 3014 -7535
rect 3048 -7569 3058 -7535
rect 3004 -7581 3058 -7569
rect 3088 -7433 3140 -7413
rect 3088 -7467 3098 -7433
rect 3132 -7467 3140 -7433
rect 3088 -7535 3140 -7467
rect 3088 -7569 3098 -7535
rect 3132 -7569 3140 -7535
rect 3286 -7433 3338 -7407
rect 3286 -7467 3294 -7433
rect 3328 -7467 3338 -7433
rect 3286 -7535 3338 -7467
rect 3088 -7581 3140 -7569
rect 3286 -7569 3294 -7535
rect 3328 -7569 3338 -7535
rect 3286 -7581 3338 -7569
rect 3548 -7433 3600 -7407
rect 3548 -7467 3558 -7433
rect 3592 -7467 3600 -7433
rect 3548 -7535 3600 -7467
rect 3548 -7569 3558 -7535
rect 3592 -7569 3600 -7535
rect 3750 -7399 3802 -7381
rect 3750 -7433 3758 -7399
rect 3792 -7433 3802 -7399
rect 3750 -7467 3802 -7433
rect 3750 -7501 3758 -7467
rect 3792 -7501 3802 -7467
rect 3750 -7535 3802 -7501
rect 3548 -7581 3600 -7569
rect 3750 -7569 3758 -7535
rect 3792 -7569 3802 -7535
rect 3750 -7581 3802 -7569
rect 3832 -7399 3886 -7381
rect 3832 -7433 3842 -7399
rect 3876 -7433 3886 -7399
rect 3832 -7467 3886 -7433
rect 3832 -7501 3842 -7467
rect 3876 -7501 3886 -7467
rect 3832 -7535 3886 -7501
rect 3832 -7569 3842 -7535
rect 3876 -7569 3886 -7535
rect 3832 -7581 3886 -7569
rect 3916 -7399 3968 -7381
rect 3916 -7433 3926 -7399
rect 3960 -7433 3968 -7399
rect 3916 -7467 3968 -7433
rect 3916 -7501 3926 -7467
rect 3960 -7501 3968 -7467
rect 3916 -7535 3968 -7501
rect 3916 -7569 3926 -7535
rect 3960 -7569 3968 -7535
rect 4114 -7433 4166 -7407
rect 4114 -7467 4122 -7433
rect 4156 -7467 4166 -7433
rect 4114 -7535 4166 -7467
rect 3916 -7581 3968 -7569
rect 4114 -7569 4122 -7535
rect 4156 -7569 4166 -7535
rect 4114 -7581 4166 -7569
rect 4376 -7433 4428 -7407
rect 4376 -7467 4386 -7433
rect 4420 -7467 4428 -7433
rect 4376 -7535 4428 -7467
rect 4376 -7569 4386 -7535
rect 4420 -7569 4428 -7535
rect 4574 -7399 4626 -7381
rect 4574 -7433 4582 -7399
rect 4616 -7433 4626 -7399
rect 4574 -7467 4626 -7433
rect 4574 -7501 4582 -7467
rect 4616 -7501 4626 -7467
rect 4574 -7535 4626 -7501
rect 4376 -7581 4428 -7569
rect 4574 -7569 4582 -7535
rect 4616 -7569 4626 -7535
rect 4574 -7581 4626 -7569
rect 4656 -7399 4708 -7381
rect 4656 -7433 4666 -7399
rect 4700 -7433 4708 -7399
rect 4656 -7458 4708 -7433
rect 4656 -7467 4735 -7458
rect 4656 -7501 4666 -7467
rect 4700 -7501 4735 -7467
rect 4656 -7535 4735 -7501
rect 4656 -7569 4666 -7535
rect 4700 -7542 4735 -7535
rect 4765 -7542 4838 -7458
rect 4868 -7475 5052 -7458
rect 4868 -7509 4902 -7475
rect 4936 -7509 4977 -7475
rect 5011 -7509 5052 -7475
rect 4868 -7542 5052 -7509
rect 5082 -7542 5124 -7458
rect 5154 -7475 5220 -7458
rect 5154 -7509 5174 -7475
rect 5208 -7509 5220 -7475
rect 5154 -7542 5220 -7509
rect 5250 -7475 5306 -7458
rect 5250 -7509 5260 -7475
rect 5294 -7509 5306 -7475
rect 5250 -7542 5306 -7509
rect 4700 -7569 4708 -7542
rect 5494 -7433 5546 -7407
rect 5494 -7467 5502 -7433
rect 5536 -7467 5546 -7433
rect 5494 -7535 5546 -7467
rect 4656 -7581 4708 -7569
rect 5494 -7569 5502 -7535
rect 5536 -7569 5546 -7535
rect 5494 -7581 5546 -7569
rect 5756 -7433 5808 -7407
rect 5756 -7467 5766 -7433
rect 5800 -7467 5808 -7433
rect 5756 -7535 5808 -7467
rect 5756 -7569 5766 -7535
rect 5800 -7569 5808 -7535
rect 5954 -7393 6006 -7381
rect 5954 -7427 5962 -7393
rect 5996 -7427 6006 -7393
rect 5954 -7464 6006 -7427
rect 5954 -7498 5962 -7464
rect 5996 -7498 6006 -7464
rect 5954 -7535 6006 -7498
rect 5756 -7581 5808 -7569
rect 5954 -7569 5962 -7535
rect 5996 -7569 6006 -7535
rect 5954 -7581 6006 -7569
rect 6036 -7399 6088 -7381
rect 6036 -7433 6046 -7399
rect 6080 -7433 6088 -7399
rect 6036 -7453 6088 -7433
rect 6239 -7393 6291 -7381
rect 6239 -7427 6247 -7393
rect 6281 -7427 6291 -7393
rect 6036 -7467 6103 -7453
rect 6036 -7501 6046 -7467
rect 6080 -7501 6103 -7467
rect 6036 -7535 6103 -7501
rect 6036 -7569 6046 -7535
rect 6080 -7569 6103 -7535
rect 6036 -7581 6103 -7569
rect 6133 -7467 6185 -7453
rect 6133 -7501 6143 -7467
rect 6177 -7501 6185 -7467
rect 6133 -7535 6185 -7501
rect 6133 -7569 6143 -7535
rect 6177 -7569 6185 -7535
rect 6133 -7581 6185 -7569
rect 6239 -7461 6291 -7427
rect 6239 -7495 6247 -7461
rect 6281 -7495 6291 -7461
rect 6239 -7529 6291 -7495
rect 6239 -7563 6247 -7529
rect 6281 -7563 6291 -7529
rect 6239 -7581 6291 -7563
rect 6321 -7425 6375 -7381
rect 6321 -7459 6331 -7425
rect 6365 -7459 6375 -7425
rect 6321 -7505 6375 -7459
rect 6321 -7539 6331 -7505
rect 6365 -7539 6375 -7505
rect 6321 -7581 6375 -7539
rect 6405 -7393 6459 -7381
rect 6405 -7427 6417 -7393
rect 6451 -7427 6459 -7393
rect 6405 -7464 6459 -7427
rect 6405 -7498 6417 -7464
rect 6451 -7498 6459 -7464
rect 6829 -7497 6879 -7431
rect 6405 -7535 6459 -7498
rect 6405 -7569 6417 -7535
rect 6451 -7569 6459 -7535
rect 6405 -7581 6459 -7569
rect 6533 -7527 6586 -7497
rect 6533 -7561 6541 -7527
rect 6575 -7561 6586 -7527
rect 6533 -7581 6586 -7561
rect 6616 -7581 6700 -7497
rect 6730 -7517 6784 -7497
rect 6730 -7551 6740 -7517
rect 6774 -7551 6784 -7517
rect 6730 -7581 6784 -7551
rect 6814 -7527 6879 -7497
rect 6814 -7561 6835 -7527
rect 6869 -7561 6879 -7527
rect 6814 -7581 6879 -7561
rect 6909 -7467 6996 -7431
rect 6909 -7501 6919 -7467
rect 6953 -7497 6996 -7467
rect 7430 -7459 7482 -7447
rect 7430 -7493 7438 -7459
rect 7472 -7493 7482 -7459
rect 6953 -7501 7011 -7497
rect 6909 -7535 7011 -7501
rect 6909 -7569 6919 -7535
rect 6953 -7569 7011 -7535
rect 6909 -7581 7011 -7569
rect 7041 -7581 7114 -7497
rect 7144 -7522 7209 -7497
rect 7144 -7556 7158 -7522
rect 7192 -7556 7209 -7522
rect 7144 -7581 7209 -7556
rect 7239 -7527 7294 -7497
rect 7239 -7561 7250 -7527
rect 7284 -7561 7294 -7527
rect 7239 -7581 7294 -7561
rect 7324 -7535 7376 -7497
rect 7324 -7569 7334 -7535
rect 7368 -7569 7376 -7535
rect 7324 -7581 7376 -7569
rect 7430 -7527 7482 -7493
rect 7430 -7561 7438 -7527
rect 7472 -7561 7482 -7527
rect 7430 -7575 7482 -7561
rect 7512 -7511 7566 -7447
rect 7512 -7545 7522 -7511
rect 7556 -7545 7566 -7511
rect 7512 -7575 7566 -7545
rect 7596 -7459 7648 -7447
rect 7596 -7493 7606 -7459
rect 7640 -7493 7648 -7459
rect 7596 -7527 7648 -7493
rect 7596 -7561 7606 -7527
rect 7640 -7561 7648 -7527
rect 7596 -7575 7648 -7561
rect 7794 -7433 7846 -7407
rect 7794 -7467 7802 -7433
rect 7836 -7467 7846 -7433
rect 7794 -7535 7846 -7467
rect 7794 -7569 7802 -7535
rect 7836 -7569 7846 -7535
rect 7794 -7581 7846 -7569
rect 8424 -7433 8476 -7407
rect 8424 -7467 8434 -7433
rect 8468 -7467 8476 -7433
rect 8424 -7535 8476 -7467
rect 8424 -7569 8434 -7535
rect 8468 -7569 8476 -7535
rect 8424 -7581 8476 -7569
rect 8530 -7433 8582 -7407
rect 8530 -7467 8538 -7433
rect 8572 -7467 8582 -7433
rect 8530 -7535 8582 -7467
rect 8530 -7569 8538 -7535
rect 8572 -7569 8582 -7535
rect 8530 -7581 8582 -7569
rect 9160 -7433 9212 -7407
rect 9160 -7467 9170 -7433
rect 9204 -7467 9212 -7433
rect 9160 -7535 9212 -7467
rect 9160 -7569 9170 -7535
rect 9204 -7569 9212 -7535
rect 15982 -7433 16034 -7407
rect 15982 -7467 15990 -7433
rect 16024 -7467 16034 -7433
rect 15982 -7535 16034 -7467
rect 9160 -7581 9212 -7569
rect 15982 -7569 15990 -7535
rect 16024 -7569 16034 -7535
rect 15982 -7581 16034 -7569
rect 16612 -7433 16664 -7407
rect 16612 -7467 16622 -7433
rect 16656 -7467 16664 -7433
rect 16612 -7535 16664 -7467
rect 16612 -7569 16622 -7535
rect 16656 -7569 16664 -7535
rect 16612 -7581 16664 -7569
rect -2970 -7687 -2918 -7675
rect -2970 -7721 -2962 -7687
rect -2928 -7721 -2918 -7687
rect -2970 -7789 -2918 -7721
rect -2970 -7823 -2962 -7789
rect -2928 -7823 -2918 -7789
rect -2970 -7849 -2918 -7823
rect -2340 -7687 -2288 -7675
rect -2340 -7721 -2330 -7687
rect -2296 -7721 -2288 -7687
rect -1406 -7687 -1354 -7675
rect -2340 -7789 -2288 -7721
rect -2340 -7823 -2330 -7789
rect -2296 -7823 -2288 -7789
rect -2340 -7849 -2288 -7823
rect -1406 -7721 -1398 -7687
rect -1364 -7721 -1354 -7687
rect -1406 -7789 -1354 -7721
rect -1406 -7823 -1398 -7789
rect -1364 -7823 -1354 -7789
rect -1406 -7849 -1354 -7823
rect -1144 -7687 -1092 -7675
rect -1144 -7721 -1134 -7687
rect -1100 -7721 -1092 -7687
rect -942 -7687 -890 -7675
rect -1144 -7789 -1092 -7721
rect -1144 -7823 -1134 -7789
rect -1100 -7823 -1092 -7789
rect -1144 -7849 -1092 -7823
rect -942 -7721 -934 -7687
rect -900 -7721 -890 -7687
rect -942 -7755 -890 -7721
rect -942 -7789 -934 -7755
rect -900 -7789 -890 -7755
rect -942 -7823 -890 -7789
rect -942 -7857 -934 -7823
rect -900 -7857 -890 -7823
rect -942 -7875 -890 -7857
rect -860 -7687 -806 -7675
rect -860 -7721 -850 -7687
rect -816 -7721 -806 -7687
rect -860 -7755 -806 -7721
rect -860 -7789 -850 -7755
rect -816 -7789 -806 -7755
rect -860 -7823 -806 -7789
rect -860 -7857 -850 -7823
rect -816 -7857 -806 -7823
rect -860 -7875 -806 -7857
rect -776 -7687 -724 -7675
rect -776 -7721 -766 -7687
rect -732 -7721 -724 -7687
rect -578 -7687 -526 -7675
rect -776 -7755 -724 -7721
rect -776 -7789 -766 -7755
rect -732 -7789 -724 -7755
rect -776 -7823 -724 -7789
rect -776 -7857 -766 -7823
rect -732 -7857 -724 -7823
rect -776 -7875 -724 -7857
rect -578 -7721 -570 -7687
rect -536 -7721 -526 -7687
rect -578 -7789 -526 -7721
rect -578 -7823 -570 -7789
rect -536 -7823 -526 -7789
rect -578 -7849 -526 -7823
rect -316 -7687 -264 -7675
rect -316 -7721 -306 -7687
rect -272 -7721 -264 -7687
rect -316 -7789 -264 -7721
rect -316 -7823 -306 -7789
rect -272 -7823 -264 -7789
rect -316 -7849 -264 -7823
rect -118 -7694 -57 -7675
rect -118 -7728 -102 -7694
rect -68 -7728 -57 -7694
rect -118 -7762 -57 -7728
rect -118 -7796 -102 -7762
rect -68 -7796 -57 -7762
rect -118 -7875 -57 -7796
rect -27 -7701 29 -7675
rect -27 -7735 -16 -7701
rect 18 -7735 29 -7701
rect -27 -7789 29 -7735
rect -27 -7823 -16 -7789
rect 18 -7823 29 -7789
rect -27 -7875 29 -7823
rect 59 -7694 115 -7675
rect 59 -7728 70 -7694
rect 104 -7728 115 -7694
rect 59 -7762 115 -7728
rect 59 -7796 70 -7762
rect 104 -7796 115 -7762
rect 59 -7875 115 -7796
rect 145 -7701 201 -7675
rect 145 -7735 156 -7701
rect 190 -7735 201 -7701
rect 145 -7789 201 -7735
rect 145 -7823 156 -7789
rect 190 -7823 201 -7789
rect 145 -7875 201 -7823
rect 231 -7694 287 -7675
rect 231 -7728 242 -7694
rect 276 -7728 287 -7694
rect 231 -7762 287 -7728
rect 231 -7796 242 -7762
rect 276 -7796 287 -7762
rect 231 -7875 287 -7796
rect 317 -7701 373 -7675
rect 317 -7735 328 -7701
rect 362 -7735 373 -7701
rect 317 -7789 373 -7735
rect 317 -7823 328 -7789
rect 362 -7823 373 -7789
rect 317 -7875 373 -7823
rect 403 -7694 472 -7675
rect 618 -7687 670 -7675
rect 403 -7728 414 -7694
rect 448 -7728 472 -7694
rect 403 -7762 472 -7728
rect 403 -7796 414 -7762
rect 448 -7796 472 -7762
rect 403 -7875 472 -7796
rect 618 -7721 626 -7687
rect 660 -7721 670 -7687
rect 618 -7789 670 -7721
rect 618 -7823 626 -7789
rect 660 -7823 670 -7789
rect 618 -7849 670 -7823
rect 880 -7687 932 -7675
rect 880 -7721 890 -7687
rect 924 -7721 932 -7687
rect 1078 -7687 1130 -7675
rect 880 -7789 932 -7721
rect 880 -7823 890 -7789
rect 924 -7823 932 -7789
rect 880 -7849 932 -7823
rect 1078 -7721 1086 -7687
rect 1120 -7721 1130 -7687
rect 1078 -7789 1130 -7721
rect 1078 -7823 1086 -7789
rect 1120 -7823 1130 -7789
rect 1078 -7843 1130 -7823
rect 1160 -7687 1214 -7675
rect 1160 -7721 1170 -7687
rect 1204 -7721 1214 -7687
rect 1160 -7789 1214 -7721
rect 1160 -7823 1170 -7789
rect 1204 -7823 1214 -7789
rect 1160 -7843 1214 -7823
rect 1244 -7687 1300 -7675
rect 1244 -7721 1254 -7687
rect 1288 -7721 1300 -7687
rect 1446 -7687 1498 -7675
rect 1244 -7789 1300 -7721
rect 1244 -7823 1254 -7789
rect 1288 -7823 1300 -7789
rect 1244 -7843 1300 -7823
rect 1446 -7721 1454 -7687
rect 1488 -7721 1498 -7687
rect 1446 -7789 1498 -7721
rect 1446 -7823 1454 -7789
rect 1488 -7823 1498 -7789
rect 1446 -7849 1498 -7823
rect 1708 -7687 1760 -7675
rect 1708 -7721 1718 -7687
rect 1752 -7721 1760 -7687
rect 1906 -7687 1958 -7675
rect 1708 -7789 1760 -7721
rect 1708 -7823 1718 -7789
rect 1752 -7823 1760 -7789
rect 1708 -7849 1760 -7823
rect 1906 -7721 1914 -7687
rect 1948 -7721 1958 -7687
rect 1906 -7789 1958 -7721
rect 1906 -7823 1914 -7789
rect 1948 -7823 1958 -7789
rect 1906 -7849 1958 -7823
rect 2168 -7687 2220 -7675
rect 2168 -7721 2178 -7687
rect 2212 -7721 2220 -7687
rect 2168 -7789 2220 -7721
rect 2168 -7823 2178 -7789
rect 2212 -7823 2220 -7789
rect 2168 -7849 2220 -7823
rect 2366 -7694 2420 -7675
rect 2366 -7728 2375 -7694
rect 2409 -7728 2420 -7694
rect 2366 -7762 2420 -7728
rect 2366 -7796 2375 -7762
rect 2409 -7796 2420 -7762
rect 2366 -7875 2420 -7796
rect 2450 -7694 2522 -7675
rect 2450 -7728 2475 -7694
rect 2509 -7728 2522 -7694
rect 2450 -7762 2522 -7728
rect 2450 -7796 2475 -7762
rect 2509 -7796 2522 -7762
rect 2450 -7839 2522 -7796
rect 2622 -7694 2675 -7675
rect 2622 -7728 2633 -7694
rect 2667 -7728 2675 -7694
rect 2622 -7762 2675 -7728
rect 2622 -7796 2633 -7762
rect 2667 -7796 2675 -7762
rect 2622 -7839 2675 -7796
rect 2729 -7695 2782 -7675
rect 2729 -7729 2737 -7695
rect 2771 -7729 2782 -7695
rect 2729 -7763 2782 -7729
rect 2729 -7797 2737 -7763
rect 2771 -7797 2782 -7763
rect 2729 -7839 2782 -7797
rect 2882 -7694 2947 -7675
rect 2882 -7728 2893 -7694
rect 2927 -7728 2947 -7694
rect 2882 -7762 2947 -7728
rect 2882 -7796 2893 -7762
rect 2927 -7796 2947 -7762
rect 2882 -7839 2947 -7796
rect 2450 -7875 2500 -7839
rect 2897 -7875 2947 -7839
rect 2977 -7695 3048 -7675
rect 3194 -7687 3246 -7675
rect 2977 -7729 2991 -7695
rect 3025 -7729 3048 -7695
rect 2977 -7763 3048 -7729
rect 2977 -7797 2991 -7763
rect 3025 -7797 3048 -7763
rect 2977 -7875 3048 -7797
rect 3194 -7721 3202 -7687
rect 3236 -7721 3246 -7687
rect 3194 -7789 3246 -7721
rect 3194 -7823 3202 -7789
rect 3236 -7823 3246 -7789
rect 3194 -7849 3246 -7823
rect 3456 -7687 3508 -7675
rect 3456 -7721 3466 -7687
rect 3500 -7721 3508 -7687
rect 4390 -7687 4442 -7675
rect 3456 -7789 3508 -7721
rect 3456 -7823 3466 -7789
rect 3500 -7823 3508 -7789
rect 3456 -7849 3508 -7823
rect 4390 -7721 4398 -7687
rect 4432 -7721 4442 -7687
rect 4390 -7789 4442 -7721
rect 4390 -7823 4398 -7789
rect 4432 -7823 4442 -7789
rect 4390 -7849 4442 -7823
rect 5388 -7687 5440 -7675
rect 5388 -7721 5398 -7687
rect 5432 -7721 5440 -7687
rect 6414 -7687 6466 -7675
rect 5388 -7789 5440 -7721
rect 5388 -7823 5398 -7789
rect 5432 -7823 5440 -7789
rect 5388 -7849 5440 -7823
rect 6414 -7721 6422 -7687
rect 6456 -7721 6466 -7687
rect 6414 -7789 6466 -7721
rect 6414 -7823 6422 -7789
rect 6456 -7823 6466 -7789
rect 6414 -7849 6466 -7823
rect 6676 -7687 6728 -7675
rect 6676 -7721 6686 -7687
rect 6720 -7721 6728 -7687
rect 6676 -7789 6728 -7721
rect 6676 -7823 6686 -7789
rect 6720 -7823 6728 -7789
rect 6676 -7849 6728 -7823
rect 6874 -7694 6928 -7675
rect 6874 -7728 6883 -7694
rect 6917 -7728 6928 -7694
rect 6874 -7762 6928 -7728
rect 6874 -7796 6883 -7762
rect 6917 -7796 6928 -7762
rect 6874 -7875 6928 -7796
rect 6958 -7694 7030 -7675
rect 6958 -7728 6983 -7694
rect 7017 -7728 7030 -7694
rect 6958 -7762 7030 -7728
rect 6958 -7796 6983 -7762
rect 7017 -7796 7030 -7762
rect 6958 -7839 7030 -7796
rect 7130 -7694 7183 -7675
rect 7130 -7728 7141 -7694
rect 7175 -7728 7183 -7694
rect 7130 -7762 7183 -7728
rect 7130 -7796 7141 -7762
rect 7175 -7796 7183 -7762
rect 7130 -7839 7183 -7796
rect 7237 -7695 7290 -7675
rect 7237 -7729 7245 -7695
rect 7279 -7729 7290 -7695
rect 7237 -7763 7290 -7729
rect 7237 -7797 7245 -7763
rect 7279 -7797 7290 -7763
rect 7237 -7839 7290 -7797
rect 7390 -7694 7455 -7675
rect 7390 -7728 7401 -7694
rect 7435 -7728 7455 -7694
rect 7390 -7762 7455 -7728
rect 7390 -7796 7401 -7762
rect 7435 -7796 7455 -7762
rect 7390 -7839 7455 -7796
rect 6958 -7875 7008 -7839
rect 7405 -7875 7455 -7839
rect 7485 -7695 7556 -7675
rect 7702 -7687 7754 -7675
rect 7485 -7729 7499 -7695
rect 7533 -7729 7556 -7695
rect 7485 -7763 7556 -7729
rect 7485 -7797 7499 -7763
rect 7533 -7797 7556 -7763
rect 7485 -7875 7556 -7797
rect 7702 -7721 7710 -7687
rect 7744 -7721 7754 -7687
rect 7702 -7789 7754 -7721
rect 7702 -7823 7710 -7789
rect 7744 -7823 7754 -7789
rect 7702 -7849 7754 -7823
rect 7964 -7687 8016 -7675
rect 7964 -7721 7974 -7687
rect 8008 -7721 8016 -7687
rect 7964 -7789 8016 -7721
rect 7964 -7823 7974 -7789
rect 8008 -7823 8016 -7789
rect 7964 -7849 8016 -7823
rect 8162 -7694 8216 -7675
rect 8162 -7728 8171 -7694
rect 8205 -7728 8216 -7694
rect 8162 -7762 8216 -7728
rect 8162 -7796 8171 -7762
rect 8205 -7796 8216 -7762
rect 8162 -7875 8216 -7796
rect 8246 -7694 8318 -7675
rect 8246 -7728 8271 -7694
rect 8305 -7728 8318 -7694
rect 8246 -7762 8318 -7728
rect 8246 -7796 8271 -7762
rect 8305 -7796 8318 -7762
rect 8246 -7839 8318 -7796
rect 8418 -7694 8471 -7675
rect 8418 -7728 8429 -7694
rect 8463 -7728 8471 -7694
rect 8418 -7762 8471 -7728
rect 8418 -7796 8429 -7762
rect 8463 -7796 8471 -7762
rect 8418 -7839 8471 -7796
rect 8525 -7695 8578 -7675
rect 8525 -7729 8533 -7695
rect 8567 -7729 8578 -7695
rect 8525 -7763 8578 -7729
rect 8525 -7797 8533 -7763
rect 8567 -7797 8578 -7763
rect 8525 -7839 8578 -7797
rect 8678 -7694 8743 -7675
rect 8678 -7728 8689 -7694
rect 8723 -7728 8743 -7694
rect 8678 -7762 8743 -7728
rect 8678 -7796 8689 -7762
rect 8723 -7796 8743 -7762
rect 8678 -7839 8743 -7796
rect 8246 -7875 8296 -7839
rect 8693 -7875 8743 -7839
rect 8773 -7695 8844 -7675
rect 8990 -7687 9042 -7675
rect 8773 -7729 8787 -7695
rect 8821 -7729 8844 -7695
rect 8773 -7763 8844 -7729
rect 8773 -7797 8787 -7763
rect 8821 -7797 8844 -7763
rect 8773 -7875 8844 -7797
rect 8990 -7721 8998 -7687
rect 9032 -7721 9042 -7687
rect 8990 -7789 9042 -7721
rect 8990 -7823 8998 -7789
rect 9032 -7823 9042 -7789
rect 8990 -7849 9042 -7823
rect 9252 -7687 9304 -7675
rect 9252 -7721 9262 -7687
rect 9296 -7721 9304 -7687
rect 9252 -7789 9304 -7721
rect 9252 -7823 9262 -7789
rect 9296 -7823 9304 -7789
rect 9252 -7849 9304 -7823
rect 9450 -7694 9504 -7675
rect 9450 -7728 9459 -7694
rect 9493 -7728 9504 -7694
rect 9450 -7762 9504 -7728
rect 9450 -7796 9459 -7762
rect 9493 -7796 9504 -7762
rect 9450 -7875 9504 -7796
rect 9534 -7694 9606 -7675
rect 9534 -7728 9559 -7694
rect 9593 -7728 9606 -7694
rect 9534 -7762 9606 -7728
rect 9534 -7796 9559 -7762
rect 9593 -7796 9606 -7762
rect 9534 -7839 9606 -7796
rect 9706 -7694 9759 -7675
rect 9706 -7728 9717 -7694
rect 9751 -7728 9759 -7694
rect 9706 -7762 9759 -7728
rect 9706 -7796 9717 -7762
rect 9751 -7796 9759 -7762
rect 9706 -7839 9759 -7796
rect 9813 -7695 9866 -7675
rect 9813 -7729 9821 -7695
rect 9855 -7729 9866 -7695
rect 9813 -7763 9866 -7729
rect 9813 -7797 9821 -7763
rect 9855 -7797 9866 -7763
rect 9813 -7839 9866 -7797
rect 9966 -7694 10031 -7675
rect 9966 -7728 9977 -7694
rect 10011 -7728 10031 -7694
rect 9966 -7762 10031 -7728
rect 9966 -7796 9977 -7762
rect 10011 -7796 10031 -7762
rect 9966 -7839 10031 -7796
rect 9534 -7875 9584 -7839
rect 9981 -7875 10031 -7839
rect 10061 -7695 10132 -7675
rect 10278 -7687 10330 -7675
rect 10061 -7729 10075 -7695
rect 10109 -7729 10132 -7695
rect 10061 -7763 10132 -7729
rect 10061 -7797 10075 -7763
rect 10109 -7797 10132 -7763
rect 10061 -7875 10132 -7797
rect 10278 -7721 10286 -7687
rect 10320 -7721 10330 -7687
rect 10278 -7789 10330 -7721
rect 10278 -7823 10286 -7789
rect 10320 -7823 10330 -7789
rect 10278 -7849 10330 -7823
rect 10540 -7687 10592 -7675
rect 10540 -7721 10550 -7687
rect 10584 -7721 10592 -7687
rect 10738 -7687 10790 -7675
rect 10540 -7789 10592 -7721
rect 10540 -7823 10550 -7789
rect 10584 -7823 10592 -7789
rect 10540 -7849 10592 -7823
rect 10738 -7721 10746 -7687
rect 10780 -7721 10790 -7687
rect 10738 -7755 10790 -7721
rect 10738 -7789 10746 -7755
rect 10780 -7789 10790 -7755
rect 10738 -7823 10790 -7789
rect 10738 -7857 10746 -7823
rect 10780 -7857 10790 -7823
rect 10738 -7875 10790 -7857
rect 10820 -7687 10874 -7675
rect 10820 -7721 10830 -7687
rect 10864 -7721 10874 -7687
rect 10820 -7755 10874 -7721
rect 10820 -7789 10830 -7755
rect 10864 -7789 10874 -7755
rect 10820 -7823 10874 -7789
rect 10820 -7857 10830 -7823
rect 10864 -7857 10874 -7823
rect 10820 -7875 10874 -7857
rect 10904 -7687 10958 -7675
rect 10904 -7721 10914 -7687
rect 10948 -7721 10958 -7687
rect 10904 -7755 10958 -7721
rect 10904 -7789 10914 -7755
rect 10948 -7789 10958 -7755
rect 10904 -7875 10958 -7789
rect 10988 -7687 11042 -7675
rect 10988 -7721 10998 -7687
rect 11032 -7721 11042 -7687
rect 10988 -7755 11042 -7721
rect 10988 -7789 10998 -7755
rect 11032 -7789 11042 -7755
rect 10988 -7823 11042 -7789
rect 10988 -7857 10998 -7823
rect 11032 -7857 11042 -7823
rect 10988 -7875 11042 -7857
rect 11072 -7687 11126 -7675
rect 11072 -7721 11082 -7687
rect 11116 -7721 11126 -7687
rect 11072 -7755 11126 -7721
rect 11072 -7789 11082 -7755
rect 11116 -7789 11126 -7755
rect 11072 -7875 11126 -7789
rect 11156 -7687 11210 -7675
rect 11156 -7721 11166 -7687
rect 11200 -7721 11210 -7687
rect 11156 -7755 11210 -7721
rect 11156 -7789 11166 -7755
rect 11200 -7789 11210 -7755
rect 11156 -7823 11210 -7789
rect 11156 -7857 11166 -7823
rect 11200 -7857 11210 -7823
rect 11156 -7875 11210 -7857
rect 11240 -7687 11294 -7675
rect 11240 -7721 11250 -7687
rect 11284 -7721 11294 -7687
rect 11240 -7755 11294 -7721
rect 11240 -7789 11250 -7755
rect 11284 -7789 11294 -7755
rect 11240 -7875 11294 -7789
rect 11324 -7687 11378 -7675
rect 11324 -7721 11334 -7687
rect 11368 -7721 11378 -7687
rect 11324 -7755 11378 -7721
rect 11324 -7789 11334 -7755
rect 11368 -7789 11378 -7755
rect 11324 -7823 11378 -7789
rect 11324 -7857 11334 -7823
rect 11368 -7857 11378 -7823
rect 11324 -7875 11378 -7857
rect 11408 -7687 11460 -7675
rect 11408 -7721 11418 -7687
rect 11452 -7721 11460 -7687
rect 11658 -7687 11710 -7675
rect 11408 -7755 11460 -7721
rect 11408 -7789 11418 -7755
rect 11452 -7789 11460 -7755
rect 11408 -7875 11460 -7789
rect 11658 -7721 11666 -7687
rect 11700 -7721 11710 -7687
rect 11658 -7789 11710 -7721
rect 11658 -7823 11666 -7789
rect 11700 -7823 11710 -7789
rect 11658 -7849 11710 -7823
rect 11920 -7687 11972 -7675
rect 11920 -7721 11930 -7687
rect 11964 -7721 11972 -7687
rect 13590 -7687 13642 -7675
rect 11920 -7789 11972 -7721
rect 11920 -7823 11930 -7789
rect 11964 -7823 11972 -7789
rect 11920 -7849 11972 -7823
rect 13590 -7721 13598 -7687
rect 13632 -7721 13642 -7687
rect 13590 -7789 13642 -7721
rect 13590 -7823 13598 -7789
rect 13632 -7823 13642 -7789
rect 13590 -7849 13642 -7823
rect 14588 -7687 14640 -7675
rect 14588 -7721 14598 -7687
rect 14632 -7721 14640 -7687
rect 14786 -7687 14838 -7675
rect 14588 -7789 14640 -7721
rect 14588 -7823 14598 -7789
rect 14632 -7823 14640 -7789
rect 14588 -7849 14640 -7823
rect 14786 -7721 14794 -7687
rect 14828 -7721 14838 -7687
rect 14786 -7789 14838 -7721
rect 14786 -7823 14794 -7789
rect 14828 -7823 14838 -7789
rect 14786 -7849 14838 -7823
rect 15784 -7687 15836 -7675
rect 15784 -7721 15794 -7687
rect 15828 -7721 15836 -7687
rect 15982 -7687 16034 -7675
rect 15784 -7789 15836 -7721
rect 15784 -7823 15794 -7789
rect 15828 -7823 15836 -7789
rect 15784 -7849 15836 -7823
rect 15982 -7721 15990 -7687
rect 16024 -7721 16034 -7687
rect 15982 -7789 16034 -7721
rect 15982 -7823 15990 -7789
rect 16024 -7823 16034 -7789
rect 15982 -7849 16034 -7823
rect 16612 -7687 16664 -7675
rect 16612 -7721 16622 -7687
rect 16656 -7721 16664 -7687
rect 16612 -7789 16664 -7721
rect 16612 -7823 16622 -7789
rect 16656 -7823 16664 -7789
rect 16612 -7849 16664 -7823
rect -2970 -8521 -2918 -8495
rect -2970 -8555 -2962 -8521
rect -2928 -8555 -2918 -8521
rect -2970 -8623 -2918 -8555
rect -2970 -8657 -2962 -8623
rect -2928 -8657 -2918 -8623
rect -2970 -8669 -2918 -8657
rect -2340 -8521 -2288 -8495
rect -2340 -8555 -2330 -8521
rect -2296 -8555 -2288 -8521
rect -2340 -8623 -2288 -8555
rect -2340 -8657 -2330 -8623
rect -2296 -8657 -2288 -8623
rect -1590 -8521 -1538 -8495
rect -1590 -8555 -1582 -8521
rect -1548 -8555 -1538 -8521
rect -1590 -8623 -1538 -8555
rect -2340 -8669 -2288 -8657
rect -1590 -8657 -1582 -8623
rect -1548 -8657 -1538 -8623
rect -1590 -8669 -1538 -8657
rect -960 -8521 -908 -8495
rect -960 -8555 -950 -8521
rect -916 -8555 -908 -8521
rect -960 -8623 -908 -8555
rect -960 -8657 -950 -8623
rect -916 -8657 -908 -8623
rect -960 -8669 -908 -8657
rect -854 -8521 -802 -8495
rect -854 -8555 -846 -8521
rect -812 -8555 -802 -8521
rect -854 -8623 -802 -8555
rect -854 -8657 -846 -8623
rect -812 -8657 -802 -8623
rect -854 -8669 -802 -8657
rect -224 -8521 -172 -8495
rect -224 -8555 -214 -8521
rect -180 -8555 -172 -8521
rect -224 -8623 -172 -8555
rect -224 -8657 -214 -8623
rect -180 -8657 -172 -8623
rect -26 -8521 26 -8495
rect -26 -8555 -18 -8521
rect 16 -8555 26 -8521
rect -26 -8623 26 -8555
rect -224 -8669 -172 -8657
rect -26 -8657 -18 -8623
rect 16 -8657 26 -8623
rect -26 -8669 26 -8657
rect 236 -8521 288 -8495
rect 236 -8555 246 -8521
rect 280 -8555 288 -8521
rect 236 -8623 288 -8555
rect 236 -8657 246 -8623
rect 280 -8657 288 -8623
rect 434 -8547 505 -8469
rect 434 -8581 457 -8547
rect 491 -8581 505 -8547
rect 434 -8615 505 -8581
rect 434 -8649 457 -8615
rect 491 -8649 505 -8615
rect 236 -8669 288 -8657
rect 434 -8669 505 -8649
rect 535 -8505 585 -8469
rect 982 -8505 1032 -8469
rect 535 -8548 600 -8505
rect 535 -8582 555 -8548
rect 589 -8582 600 -8548
rect 535 -8616 600 -8582
rect 535 -8650 555 -8616
rect 589 -8650 600 -8616
rect 535 -8669 600 -8650
rect 700 -8547 753 -8505
rect 700 -8581 711 -8547
rect 745 -8581 753 -8547
rect 700 -8615 753 -8581
rect 700 -8649 711 -8615
rect 745 -8649 753 -8615
rect 700 -8669 753 -8649
rect 807 -8548 860 -8505
rect 807 -8582 815 -8548
rect 849 -8582 860 -8548
rect 807 -8616 860 -8582
rect 807 -8650 815 -8616
rect 849 -8650 860 -8616
rect 807 -8669 860 -8650
rect 960 -8548 1032 -8505
rect 960 -8582 973 -8548
rect 1007 -8582 1032 -8548
rect 960 -8616 1032 -8582
rect 960 -8650 973 -8616
rect 1007 -8650 1032 -8616
rect 960 -8669 1032 -8650
rect 1062 -8548 1116 -8469
rect 1062 -8582 1073 -8548
rect 1107 -8582 1116 -8548
rect 1062 -8616 1116 -8582
rect 1062 -8650 1073 -8616
rect 1107 -8650 1116 -8616
rect 1062 -8669 1116 -8650
rect 1262 -8521 1314 -8495
rect 1262 -8555 1270 -8521
rect 1304 -8555 1314 -8521
rect 1262 -8623 1314 -8555
rect 1262 -8657 1270 -8623
rect 1304 -8657 1314 -8623
rect 1262 -8669 1314 -8657
rect 1524 -8521 1576 -8495
rect 1524 -8555 1534 -8521
rect 1568 -8555 1576 -8521
rect 1524 -8623 1576 -8555
rect 1524 -8657 1534 -8623
rect 1568 -8657 1576 -8623
rect 1722 -8521 1774 -8495
rect 1722 -8555 1730 -8521
rect 1764 -8555 1774 -8521
rect 1722 -8623 1774 -8555
rect 1524 -8669 1576 -8657
rect 1722 -8657 1730 -8623
rect 1764 -8657 1774 -8623
rect 1722 -8669 1774 -8657
rect 2352 -8521 2404 -8495
rect 2352 -8555 2362 -8521
rect 2396 -8555 2404 -8521
rect 2352 -8623 2404 -8555
rect 2352 -8657 2362 -8623
rect 2396 -8657 2404 -8623
rect 2550 -8521 2602 -8495
rect 2550 -8555 2558 -8521
rect 2592 -8555 2602 -8521
rect 2550 -8623 2602 -8555
rect 2352 -8669 2404 -8657
rect 2550 -8657 2558 -8623
rect 2592 -8657 2602 -8623
rect 2550 -8669 2602 -8657
rect 2812 -8521 2864 -8495
rect 2812 -8555 2822 -8521
rect 2856 -8555 2864 -8521
rect 2812 -8623 2864 -8555
rect 2812 -8657 2822 -8623
rect 2856 -8657 2864 -8623
rect 3010 -8547 3081 -8469
rect 3010 -8581 3033 -8547
rect 3067 -8581 3081 -8547
rect 3010 -8615 3081 -8581
rect 3010 -8649 3033 -8615
rect 3067 -8649 3081 -8615
rect 2812 -8669 2864 -8657
rect 3010 -8669 3081 -8649
rect 3111 -8505 3161 -8469
rect 3558 -8505 3608 -8469
rect 3111 -8548 3176 -8505
rect 3111 -8582 3131 -8548
rect 3165 -8582 3176 -8548
rect 3111 -8616 3176 -8582
rect 3111 -8650 3131 -8616
rect 3165 -8650 3176 -8616
rect 3111 -8669 3176 -8650
rect 3276 -8547 3329 -8505
rect 3276 -8581 3287 -8547
rect 3321 -8581 3329 -8547
rect 3276 -8615 3329 -8581
rect 3276 -8649 3287 -8615
rect 3321 -8649 3329 -8615
rect 3276 -8669 3329 -8649
rect 3383 -8548 3436 -8505
rect 3383 -8582 3391 -8548
rect 3425 -8582 3436 -8548
rect 3383 -8616 3436 -8582
rect 3383 -8650 3391 -8616
rect 3425 -8650 3436 -8616
rect 3383 -8669 3436 -8650
rect 3536 -8548 3608 -8505
rect 3536 -8582 3549 -8548
rect 3583 -8582 3608 -8548
rect 3536 -8616 3608 -8582
rect 3536 -8650 3549 -8616
rect 3583 -8650 3608 -8616
rect 3536 -8669 3608 -8650
rect 3638 -8548 3692 -8469
rect 3638 -8582 3649 -8548
rect 3683 -8582 3692 -8548
rect 3638 -8616 3692 -8582
rect 3638 -8650 3649 -8616
rect 3683 -8650 3692 -8616
rect 3638 -8669 3692 -8650
rect 3838 -8521 3890 -8495
rect 3838 -8555 3846 -8521
rect 3880 -8555 3890 -8521
rect 3838 -8623 3890 -8555
rect 3838 -8657 3846 -8623
rect 3880 -8657 3890 -8623
rect 3838 -8669 3890 -8657
rect 4100 -8521 4152 -8495
rect 4100 -8555 4110 -8521
rect 4144 -8555 4152 -8521
rect 4100 -8623 4152 -8555
rect 4100 -8657 4110 -8623
rect 4144 -8657 4152 -8623
rect 4298 -8521 4350 -8495
rect 4298 -8555 4306 -8521
rect 4340 -8555 4350 -8521
rect 4298 -8623 4350 -8555
rect 4100 -8669 4152 -8657
rect 4298 -8657 4306 -8623
rect 4340 -8657 4350 -8623
rect 4298 -8669 4350 -8657
rect 4928 -8521 4980 -8495
rect 4928 -8555 4938 -8521
rect 4972 -8555 4980 -8521
rect 4928 -8623 4980 -8555
rect 4928 -8657 4938 -8623
rect 4972 -8657 4980 -8623
rect 5126 -8521 5178 -8495
rect 5126 -8555 5134 -8521
rect 5168 -8555 5178 -8521
rect 5126 -8623 5178 -8555
rect 4928 -8669 4980 -8657
rect 5126 -8657 5134 -8623
rect 5168 -8657 5178 -8623
rect 5126 -8669 5178 -8657
rect 5388 -8521 5440 -8495
rect 5388 -8555 5398 -8521
rect 5432 -8555 5440 -8521
rect 5388 -8623 5440 -8555
rect 5388 -8657 5398 -8623
rect 5432 -8657 5440 -8623
rect 5586 -8547 5657 -8469
rect 5586 -8581 5609 -8547
rect 5643 -8581 5657 -8547
rect 5586 -8615 5657 -8581
rect 5586 -8649 5609 -8615
rect 5643 -8649 5657 -8615
rect 5388 -8669 5440 -8657
rect 5586 -8669 5657 -8649
rect 5687 -8505 5737 -8469
rect 6134 -8505 6184 -8469
rect 5687 -8548 5752 -8505
rect 5687 -8582 5707 -8548
rect 5741 -8582 5752 -8548
rect 5687 -8616 5752 -8582
rect 5687 -8650 5707 -8616
rect 5741 -8650 5752 -8616
rect 5687 -8669 5752 -8650
rect 5852 -8547 5905 -8505
rect 5852 -8581 5863 -8547
rect 5897 -8581 5905 -8547
rect 5852 -8615 5905 -8581
rect 5852 -8649 5863 -8615
rect 5897 -8649 5905 -8615
rect 5852 -8669 5905 -8649
rect 5959 -8548 6012 -8505
rect 5959 -8582 5967 -8548
rect 6001 -8582 6012 -8548
rect 5959 -8616 6012 -8582
rect 5959 -8650 5967 -8616
rect 6001 -8650 6012 -8616
rect 5959 -8669 6012 -8650
rect 6112 -8548 6184 -8505
rect 6112 -8582 6125 -8548
rect 6159 -8582 6184 -8548
rect 6112 -8616 6184 -8582
rect 6112 -8650 6125 -8616
rect 6159 -8650 6184 -8616
rect 6112 -8669 6184 -8650
rect 6214 -8548 6268 -8469
rect 6214 -8582 6225 -8548
rect 6259 -8582 6268 -8548
rect 6214 -8616 6268 -8582
rect 6214 -8650 6225 -8616
rect 6259 -8650 6268 -8616
rect 6214 -8669 6268 -8650
rect 6414 -8521 6466 -8495
rect 6414 -8555 6422 -8521
rect 6456 -8555 6466 -8521
rect 6414 -8623 6466 -8555
rect 6414 -8657 6422 -8623
rect 6456 -8657 6466 -8623
rect 6414 -8669 6466 -8657
rect 6676 -8521 6728 -8495
rect 6676 -8555 6686 -8521
rect 6720 -8555 6728 -8521
rect 6676 -8623 6728 -8555
rect 6676 -8657 6686 -8623
rect 6720 -8657 6728 -8623
rect 6874 -8521 6926 -8495
rect 6874 -8555 6882 -8521
rect 6916 -8555 6926 -8521
rect 6874 -8623 6926 -8555
rect 6676 -8669 6728 -8657
rect 6874 -8657 6882 -8623
rect 6916 -8657 6926 -8623
rect 6874 -8669 6926 -8657
rect 7504 -8521 7556 -8495
rect 7504 -8555 7514 -8521
rect 7548 -8555 7556 -8521
rect 7504 -8623 7556 -8555
rect 7504 -8657 7514 -8623
rect 7548 -8657 7556 -8623
rect 7702 -8521 7754 -8495
rect 7702 -8555 7710 -8521
rect 7744 -8555 7754 -8521
rect 7702 -8623 7754 -8555
rect 7504 -8669 7556 -8657
rect 7702 -8657 7710 -8623
rect 7744 -8657 7754 -8623
rect 7702 -8669 7754 -8657
rect 7964 -8521 8016 -8495
rect 7964 -8555 7974 -8521
rect 8008 -8555 8016 -8521
rect 7964 -8623 8016 -8555
rect 7964 -8657 7974 -8623
rect 8008 -8657 8016 -8623
rect 8162 -8547 8233 -8469
rect 8162 -8581 8185 -8547
rect 8219 -8581 8233 -8547
rect 8162 -8615 8233 -8581
rect 8162 -8649 8185 -8615
rect 8219 -8649 8233 -8615
rect 7964 -8669 8016 -8657
rect 8162 -8669 8233 -8649
rect 8263 -8505 8313 -8469
rect 8710 -8505 8760 -8469
rect 8263 -8548 8328 -8505
rect 8263 -8582 8283 -8548
rect 8317 -8582 8328 -8548
rect 8263 -8616 8328 -8582
rect 8263 -8650 8283 -8616
rect 8317 -8650 8328 -8616
rect 8263 -8669 8328 -8650
rect 8428 -8547 8481 -8505
rect 8428 -8581 8439 -8547
rect 8473 -8581 8481 -8547
rect 8428 -8615 8481 -8581
rect 8428 -8649 8439 -8615
rect 8473 -8649 8481 -8615
rect 8428 -8669 8481 -8649
rect 8535 -8548 8588 -8505
rect 8535 -8582 8543 -8548
rect 8577 -8582 8588 -8548
rect 8535 -8616 8588 -8582
rect 8535 -8650 8543 -8616
rect 8577 -8650 8588 -8616
rect 8535 -8669 8588 -8650
rect 8688 -8548 8760 -8505
rect 8688 -8582 8701 -8548
rect 8735 -8582 8760 -8548
rect 8688 -8616 8760 -8582
rect 8688 -8650 8701 -8616
rect 8735 -8650 8760 -8616
rect 8688 -8669 8760 -8650
rect 8790 -8548 8844 -8469
rect 8790 -8582 8801 -8548
rect 8835 -8582 8844 -8548
rect 8790 -8616 8844 -8582
rect 8790 -8650 8801 -8616
rect 8835 -8650 8844 -8616
rect 8790 -8669 8844 -8650
rect 8990 -8521 9042 -8495
rect 8990 -8555 8998 -8521
rect 9032 -8555 9042 -8521
rect 8990 -8623 9042 -8555
rect 8990 -8657 8998 -8623
rect 9032 -8657 9042 -8623
rect 8990 -8669 9042 -8657
rect 9252 -8521 9304 -8495
rect 9252 -8555 9262 -8521
rect 9296 -8555 9304 -8521
rect 9252 -8623 9304 -8555
rect 9252 -8657 9262 -8623
rect 9296 -8657 9304 -8623
rect 9450 -8521 9502 -8495
rect 9450 -8555 9458 -8521
rect 9492 -8555 9502 -8521
rect 9450 -8623 9502 -8555
rect 9252 -8669 9304 -8657
rect 9450 -8657 9458 -8623
rect 9492 -8657 9502 -8623
rect 9450 -8669 9502 -8657
rect 10080 -8521 10132 -8495
rect 10080 -8555 10090 -8521
rect 10124 -8555 10132 -8521
rect 10080 -8623 10132 -8555
rect 10080 -8657 10090 -8623
rect 10124 -8657 10132 -8623
rect 10370 -8521 10422 -8495
rect 10370 -8555 10378 -8521
rect 10412 -8555 10422 -8521
rect 10370 -8623 10422 -8555
rect 10080 -8669 10132 -8657
rect 10370 -8657 10378 -8623
rect 10412 -8657 10422 -8623
rect 10370 -8669 10422 -8657
rect 10632 -8521 10684 -8495
rect 10632 -8555 10642 -8521
rect 10676 -8555 10684 -8521
rect 10632 -8623 10684 -8555
rect 10632 -8657 10642 -8623
rect 10676 -8657 10684 -8623
rect 10632 -8669 10684 -8657
rect 10738 -8547 10809 -8469
rect 10738 -8581 10761 -8547
rect 10795 -8581 10809 -8547
rect 10738 -8615 10809 -8581
rect 10738 -8649 10761 -8615
rect 10795 -8649 10809 -8615
rect 10738 -8669 10809 -8649
rect 10839 -8505 10889 -8469
rect 11286 -8505 11336 -8469
rect 10839 -8548 10904 -8505
rect 10839 -8582 10859 -8548
rect 10893 -8582 10904 -8548
rect 10839 -8616 10904 -8582
rect 10839 -8650 10859 -8616
rect 10893 -8650 10904 -8616
rect 10839 -8669 10904 -8650
rect 11004 -8547 11057 -8505
rect 11004 -8581 11015 -8547
rect 11049 -8581 11057 -8547
rect 11004 -8615 11057 -8581
rect 11004 -8649 11015 -8615
rect 11049 -8649 11057 -8615
rect 11004 -8669 11057 -8649
rect 11111 -8548 11164 -8505
rect 11111 -8582 11119 -8548
rect 11153 -8582 11164 -8548
rect 11111 -8616 11164 -8582
rect 11111 -8650 11119 -8616
rect 11153 -8650 11164 -8616
rect 11111 -8669 11164 -8650
rect 11264 -8548 11336 -8505
rect 11264 -8582 11277 -8548
rect 11311 -8582 11336 -8548
rect 11264 -8616 11336 -8582
rect 11264 -8650 11277 -8616
rect 11311 -8650 11336 -8616
rect 11264 -8669 11336 -8650
rect 11366 -8548 11420 -8469
rect 11366 -8582 11377 -8548
rect 11411 -8582 11420 -8548
rect 11366 -8616 11420 -8582
rect 11366 -8650 11377 -8616
rect 11411 -8650 11420 -8616
rect 11366 -8669 11420 -8650
rect 11658 -8521 11710 -8495
rect 11658 -8555 11666 -8521
rect 11700 -8555 11710 -8521
rect 11658 -8623 11710 -8555
rect 11658 -8657 11666 -8623
rect 11700 -8657 11710 -8623
rect 11658 -8669 11710 -8657
rect 11920 -8521 11972 -8495
rect 11920 -8555 11930 -8521
rect 11964 -8555 11972 -8521
rect 11920 -8623 11972 -8555
rect 11920 -8657 11930 -8623
rect 11964 -8657 11972 -8623
rect 13682 -8555 13735 -8469
rect 13682 -8589 13690 -8555
rect 13724 -8589 13735 -8555
rect 13682 -8623 13735 -8589
rect 11920 -8669 11972 -8657
rect 13682 -8657 13690 -8623
rect 13724 -8657 13735 -8623
rect 13682 -8669 13735 -8657
rect 13765 -8547 13821 -8469
rect 13765 -8581 13776 -8547
rect 13810 -8581 13821 -8547
rect 13765 -8615 13821 -8581
rect 13765 -8649 13776 -8615
rect 13810 -8649 13821 -8615
rect 13765 -8669 13821 -8649
rect 13851 -8555 13907 -8469
rect 13851 -8589 13862 -8555
rect 13896 -8589 13907 -8555
rect 13851 -8623 13907 -8589
rect 13851 -8657 13862 -8623
rect 13896 -8657 13907 -8623
rect 13851 -8669 13907 -8657
rect 13937 -8539 13993 -8469
rect 13937 -8573 13948 -8539
rect 13982 -8573 13993 -8539
rect 13937 -8607 13993 -8573
rect 13937 -8641 13948 -8607
rect 13982 -8641 13993 -8607
rect 13937 -8669 13993 -8641
rect 14023 -8555 14079 -8469
rect 14023 -8589 14034 -8555
rect 14068 -8589 14079 -8555
rect 14023 -8623 14079 -8589
rect 14023 -8657 14034 -8623
rect 14068 -8657 14079 -8623
rect 14023 -8669 14079 -8657
rect 14109 -8493 14165 -8469
rect 14109 -8527 14120 -8493
rect 14154 -8527 14165 -8493
rect 14109 -8579 14165 -8527
rect 14109 -8613 14120 -8579
rect 14154 -8613 14165 -8579
rect 14109 -8669 14165 -8613
rect 14195 -8599 14251 -8469
rect 14195 -8633 14206 -8599
rect 14240 -8633 14251 -8599
rect 14195 -8669 14251 -8633
rect 14281 -8493 14337 -8469
rect 14281 -8527 14292 -8493
rect 14326 -8527 14337 -8493
rect 14281 -8579 14337 -8527
rect 14281 -8613 14292 -8579
rect 14326 -8613 14337 -8579
rect 14281 -8669 14337 -8613
rect 14367 -8599 14423 -8469
rect 14367 -8633 14378 -8599
rect 14412 -8633 14423 -8599
rect 14367 -8669 14423 -8633
rect 14453 -8493 14509 -8469
rect 14453 -8527 14464 -8493
rect 14498 -8527 14509 -8493
rect 14453 -8579 14509 -8527
rect 14453 -8613 14464 -8579
rect 14498 -8613 14509 -8579
rect 14453 -8669 14509 -8613
rect 14539 -8599 14595 -8469
rect 14539 -8633 14550 -8599
rect 14584 -8633 14595 -8599
rect 14539 -8669 14595 -8633
rect 14625 -8493 14681 -8469
rect 14625 -8527 14636 -8493
rect 14670 -8527 14681 -8493
rect 14625 -8579 14681 -8527
rect 14625 -8613 14636 -8579
rect 14670 -8613 14681 -8579
rect 14625 -8669 14681 -8613
rect 14711 -8599 14766 -8469
rect 14711 -8633 14722 -8599
rect 14756 -8633 14766 -8599
rect 14711 -8669 14766 -8633
rect 14796 -8493 14852 -8469
rect 14796 -8527 14807 -8493
rect 14841 -8527 14852 -8493
rect 14796 -8579 14852 -8527
rect 14796 -8613 14807 -8579
rect 14841 -8613 14852 -8579
rect 14796 -8669 14852 -8613
rect 14882 -8599 14938 -8469
rect 14882 -8633 14893 -8599
rect 14927 -8633 14938 -8599
rect 14882 -8669 14938 -8633
rect 14968 -8493 15024 -8469
rect 14968 -8527 14979 -8493
rect 15013 -8527 15024 -8493
rect 14968 -8579 15024 -8527
rect 14968 -8613 14979 -8579
rect 15013 -8613 15024 -8579
rect 14968 -8669 15024 -8613
rect 15054 -8599 15110 -8469
rect 15054 -8633 15065 -8599
rect 15099 -8633 15110 -8599
rect 15054 -8669 15110 -8633
rect 15140 -8493 15196 -8469
rect 15140 -8527 15151 -8493
rect 15185 -8527 15196 -8493
rect 15140 -8579 15196 -8527
rect 15140 -8613 15151 -8579
rect 15185 -8613 15196 -8579
rect 15140 -8669 15196 -8613
rect 15226 -8599 15282 -8469
rect 15226 -8633 15237 -8599
rect 15271 -8633 15282 -8599
rect 15226 -8669 15282 -8633
rect 15312 -8493 15368 -8469
rect 15312 -8527 15323 -8493
rect 15357 -8527 15368 -8493
rect 15312 -8579 15368 -8527
rect 15312 -8613 15323 -8579
rect 15357 -8613 15368 -8579
rect 15312 -8669 15368 -8613
rect 15398 -8599 15451 -8469
rect 15398 -8633 15409 -8599
rect 15443 -8633 15451 -8599
rect 15398 -8669 15451 -8633
rect 15614 -8521 15666 -8495
rect 15614 -8555 15622 -8521
rect 15656 -8555 15666 -8521
rect 15614 -8623 15666 -8555
rect 15614 -8657 15622 -8623
rect 15656 -8657 15666 -8623
rect 15614 -8669 15666 -8657
rect 16612 -8521 16664 -8495
rect 16612 -8555 16622 -8521
rect 16656 -8555 16664 -8521
rect 16612 -8623 16664 -8555
rect 16612 -8657 16622 -8623
rect 16656 -8657 16664 -8623
rect 16612 -8669 16664 -8657
rect -2970 -8775 -2918 -8763
rect -2970 -8809 -2962 -8775
rect -2928 -8809 -2918 -8775
rect -2970 -8877 -2918 -8809
rect -2970 -8911 -2962 -8877
rect -2928 -8911 -2918 -8877
rect -2970 -8937 -2918 -8911
rect -2340 -8775 -2288 -8763
rect -2340 -8809 -2330 -8775
rect -2296 -8809 -2288 -8775
rect -1590 -8775 -1538 -8763
rect -2340 -8877 -2288 -8809
rect -2340 -8911 -2330 -8877
rect -2296 -8911 -2288 -8877
rect -2340 -8937 -2288 -8911
rect -1590 -8809 -1582 -8775
rect -1548 -8809 -1538 -8775
rect -1590 -8877 -1538 -8809
rect -1590 -8911 -1582 -8877
rect -1548 -8911 -1538 -8877
rect -1590 -8937 -1538 -8911
rect -960 -8775 -908 -8763
rect -960 -8809 -950 -8775
rect -916 -8809 -908 -8775
rect -960 -8877 -908 -8809
rect -960 -8911 -950 -8877
rect -916 -8911 -908 -8877
rect -960 -8937 -908 -8911
rect -854 -8775 -802 -8763
rect -854 -8809 -846 -8775
rect -812 -8809 -802 -8775
rect -854 -8877 -802 -8809
rect -854 -8911 -846 -8877
rect -812 -8911 -802 -8877
rect -854 -8937 -802 -8911
rect -224 -8775 -172 -8763
rect -224 -8809 -214 -8775
rect -180 -8809 -172 -8775
rect -26 -8775 26 -8763
rect -224 -8877 -172 -8809
rect -224 -8911 -214 -8877
rect -180 -8911 -172 -8877
rect -224 -8937 -172 -8911
rect -26 -8809 -18 -8775
rect 16 -8809 26 -8775
rect -26 -8877 26 -8809
rect -26 -8911 -18 -8877
rect 16 -8911 26 -8877
rect -26 -8937 26 -8911
rect 236 -8775 288 -8763
rect 236 -8809 246 -8775
rect 280 -8809 288 -8775
rect 236 -8877 288 -8809
rect 236 -8911 246 -8877
rect 280 -8911 288 -8877
rect 236 -8937 288 -8911
rect 434 -8782 488 -8763
rect 434 -8816 443 -8782
rect 477 -8816 488 -8782
rect 434 -8850 488 -8816
rect 434 -8884 443 -8850
rect 477 -8884 488 -8850
rect 434 -8963 488 -8884
rect 518 -8782 590 -8763
rect 518 -8816 543 -8782
rect 577 -8816 590 -8782
rect 518 -8850 590 -8816
rect 518 -8884 543 -8850
rect 577 -8884 590 -8850
rect 518 -8927 590 -8884
rect 690 -8782 743 -8763
rect 690 -8816 701 -8782
rect 735 -8816 743 -8782
rect 690 -8850 743 -8816
rect 690 -8884 701 -8850
rect 735 -8884 743 -8850
rect 690 -8927 743 -8884
rect 797 -8783 850 -8763
rect 797 -8817 805 -8783
rect 839 -8817 850 -8783
rect 797 -8851 850 -8817
rect 797 -8885 805 -8851
rect 839 -8885 850 -8851
rect 797 -8927 850 -8885
rect 950 -8782 1015 -8763
rect 950 -8816 961 -8782
rect 995 -8816 1015 -8782
rect 950 -8850 1015 -8816
rect 950 -8884 961 -8850
rect 995 -8884 1015 -8850
rect 950 -8927 1015 -8884
rect 518 -8963 568 -8927
rect 965 -8963 1015 -8927
rect 1045 -8783 1116 -8763
rect 1262 -8775 1314 -8763
rect 1045 -8817 1059 -8783
rect 1093 -8817 1116 -8783
rect 1045 -8851 1116 -8817
rect 1045 -8885 1059 -8851
rect 1093 -8885 1116 -8851
rect 1045 -8963 1116 -8885
rect 1262 -8809 1270 -8775
rect 1304 -8809 1314 -8775
rect 1262 -8877 1314 -8809
rect 1262 -8911 1270 -8877
rect 1304 -8911 1314 -8877
rect 1262 -8937 1314 -8911
rect 1524 -8775 1576 -8763
rect 1524 -8809 1534 -8775
rect 1568 -8809 1576 -8775
rect 1722 -8775 1774 -8763
rect 1524 -8877 1576 -8809
rect 1524 -8911 1534 -8877
rect 1568 -8911 1576 -8877
rect 1524 -8937 1576 -8911
rect 1722 -8809 1730 -8775
rect 1764 -8809 1774 -8775
rect 1722 -8877 1774 -8809
rect 1722 -8911 1730 -8877
rect 1764 -8911 1774 -8877
rect 1722 -8937 1774 -8911
rect 2352 -8775 2404 -8763
rect 2352 -8809 2362 -8775
rect 2396 -8809 2404 -8775
rect 2550 -8775 2602 -8763
rect 2352 -8877 2404 -8809
rect 2352 -8911 2362 -8877
rect 2396 -8911 2404 -8877
rect 2352 -8937 2404 -8911
rect 2550 -8809 2558 -8775
rect 2592 -8809 2602 -8775
rect 2550 -8877 2602 -8809
rect 2550 -8911 2558 -8877
rect 2592 -8911 2602 -8877
rect 2550 -8937 2602 -8911
rect 2812 -8775 2864 -8763
rect 2812 -8809 2822 -8775
rect 2856 -8809 2864 -8775
rect 2812 -8877 2864 -8809
rect 2812 -8911 2822 -8877
rect 2856 -8911 2864 -8877
rect 2812 -8937 2864 -8911
rect 3010 -8782 3064 -8763
rect 3010 -8816 3019 -8782
rect 3053 -8816 3064 -8782
rect 3010 -8850 3064 -8816
rect 3010 -8884 3019 -8850
rect 3053 -8884 3064 -8850
rect 3010 -8963 3064 -8884
rect 3094 -8782 3166 -8763
rect 3094 -8816 3119 -8782
rect 3153 -8816 3166 -8782
rect 3094 -8850 3166 -8816
rect 3094 -8884 3119 -8850
rect 3153 -8884 3166 -8850
rect 3094 -8927 3166 -8884
rect 3266 -8782 3319 -8763
rect 3266 -8816 3277 -8782
rect 3311 -8816 3319 -8782
rect 3266 -8850 3319 -8816
rect 3266 -8884 3277 -8850
rect 3311 -8884 3319 -8850
rect 3266 -8927 3319 -8884
rect 3373 -8783 3426 -8763
rect 3373 -8817 3381 -8783
rect 3415 -8817 3426 -8783
rect 3373 -8851 3426 -8817
rect 3373 -8885 3381 -8851
rect 3415 -8885 3426 -8851
rect 3373 -8927 3426 -8885
rect 3526 -8782 3591 -8763
rect 3526 -8816 3537 -8782
rect 3571 -8816 3591 -8782
rect 3526 -8850 3591 -8816
rect 3526 -8884 3537 -8850
rect 3571 -8884 3591 -8850
rect 3526 -8927 3591 -8884
rect 3094 -8963 3144 -8927
rect 3541 -8963 3591 -8927
rect 3621 -8783 3692 -8763
rect 3838 -8775 3890 -8763
rect 3621 -8817 3635 -8783
rect 3669 -8817 3692 -8783
rect 3621 -8851 3692 -8817
rect 3621 -8885 3635 -8851
rect 3669 -8885 3692 -8851
rect 3621 -8963 3692 -8885
rect 3838 -8809 3846 -8775
rect 3880 -8809 3890 -8775
rect 3838 -8877 3890 -8809
rect 3838 -8911 3846 -8877
rect 3880 -8911 3890 -8877
rect 3838 -8937 3890 -8911
rect 4100 -8775 4152 -8763
rect 4100 -8809 4110 -8775
rect 4144 -8809 4152 -8775
rect 4298 -8775 4350 -8763
rect 4100 -8877 4152 -8809
rect 4100 -8911 4110 -8877
rect 4144 -8911 4152 -8877
rect 4100 -8937 4152 -8911
rect 4298 -8809 4306 -8775
rect 4340 -8809 4350 -8775
rect 4298 -8877 4350 -8809
rect 4298 -8911 4306 -8877
rect 4340 -8911 4350 -8877
rect 4298 -8937 4350 -8911
rect 4928 -8775 4980 -8763
rect 4928 -8809 4938 -8775
rect 4972 -8809 4980 -8775
rect 5126 -8775 5178 -8763
rect 4928 -8877 4980 -8809
rect 4928 -8911 4938 -8877
rect 4972 -8911 4980 -8877
rect 4928 -8937 4980 -8911
rect 5126 -8809 5134 -8775
rect 5168 -8809 5178 -8775
rect 5126 -8877 5178 -8809
rect 5126 -8911 5134 -8877
rect 5168 -8911 5178 -8877
rect 5126 -8937 5178 -8911
rect 5388 -8775 5440 -8763
rect 5388 -8809 5398 -8775
rect 5432 -8809 5440 -8775
rect 5388 -8877 5440 -8809
rect 5388 -8911 5398 -8877
rect 5432 -8911 5440 -8877
rect 5388 -8937 5440 -8911
rect 5586 -8782 5640 -8763
rect 5586 -8816 5595 -8782
rect 5629 -8816 5640 -8782
rect 5586 -8850 5640 -8816
rect 5586 -8884 5595 -8850
rect 5629 -8884 5640 -8850
rect 5586 -8963 5640 -8884
rect 5670 -8782 5742 -8763
rect 5670 -8816 5695 -8782
rect 5729 -8816 5742 -8782
rect 5670 -8850 5742 -8816
rect 5670 -8884 5695 -8850
rect 5729 -8884 5742 -8850
rect 5670 -8927 5742 -8884
rect 5842 -8782 5895 -8763
rect 5842 -8816 5853 -8782
rect 5887 -8816 5895 -8782
rect 5842 -8850 5895 -8816
rect 5842 -8884 5853 -8850
rect 5887 -8884 5895 -8850
rect 5842 -8927 5895 -8884
rect 5949 -8783 6002 -8763
rect 5949 -8817 5957 -8783
rect 5991 -8817 6002 -8783
rect 5949 -8851 6002 -8817
rect 5949 -8885 5957 -8851
rect 5991 -8885 6002 -8851
rect 5949 -8927 6002 -8885
rect 6102 -8782 6167 -8763
rect 6102 -8816 6113 -8782
rect 6147 -8816 6167 -8782
rect 6102 -8850 6167 -8816
rect 6102 -8884 6113 -8850
rect 6147 -8884 6167 -8850
rect 6102 -8927 6167 -8884
rect 5670 -8963 5720 -8927
rect 6117 -8963 6167 -8927
rect 6197 -8783 6268 -8763
rect 6414 -8775 6466 -8763
rect 6197 -8817 6211 -8783
rect 6245 -8817 6268 -8783
rect 6197 -8851 6268 -8817
rect 6197 -8885 6211 -8851
rect 6245 -8885 6268 -8851
rect 6197 -8963 6268 -8885
rect 6414 -8809 6422 -8775
rect 6456 -8809 6466 -8775
rect 6414 -8877 6466 -8809
rect 6414 -8911 6422 -8877
rect 6456 -8911 6466 -8877
rect 6414 -8937 6466 -8911
rect 6676 -8775 6728 -8763
rect 6676 -8809 6686 -8775
rect 6720 -8809 6728 -8775
rect 6874 -8775 6926 -8763
rect 6676 -8877 6728 -8809
rect 6676 -8911 6686 -8877
rect 6720 -8911 6728 -8877
rect 6676 -8937 6728 -8911
rect 6874 -8809 6882 -8775
rect 6916 -8809 6926 -8775
rect 6874 -8877 6926 -8809
rect 6874 -8911 6882 -8877
rect 6916 -8911 6926 -8877
rect 6874 -8937 6926 -8911
rect 7504 -8775 7556 -8763
rect 7504 -8809 7514 -8775
rect 7548 -8809 7556 -8775
rect 7702 -8775 7754 -8763
rect 7504 -8877 7556 -8809
rect 7504 -8911 7514 -8877
rect 7548 -8911 7556 -8877
rect 7504 -8937 7556 -8911
rect 7702 -8809 7710 -8775
rect 7744 -8809 7754 -8775
rect 7702 -8877 7754 -8809
rect 7702 -8911 7710 -8877
rect 7744 -8911 7754 -8877
rect 7702 -8937 7754 -8911
rect 7964 -8775 8016 -8763
rect 7964 -8809 7974 -8775
rect 8008 -8809 8016 -8775
rect 7964 -8877 8016 -8809
rect 7964 -8911 7974 -8877
rect 8008 -8911 8016 -8877
rect 7964 -8937 8016 -8911
rect 8162 -8782 8216 -8763
rect 8162 -8816 8171 -8782
rect 8205 -8816 8216 -8782
rect 8162 -8850 8216 -8816
rect 8162 -8884 8171 -8850
rect 8205 -8884 8216 -8850
rect 8162 -8963 8216 -8884
rect 8246 -8782 8318 -8763
rect 8246 -8816 8271 -8782
rect 8305 -8816 8318 -8782
rect 8246 -8850 8318 -8816
rect 8246 -8884 8271 -8850
rect 8305 -8884 8318 -8850
rect 8246 -8927 8318 -8884
rect 8418 -8782 8471 -8763
rect 8418 -8816 8429 -8782
rect 8463 -8816 8471 -8782
rect 8418 -8850 8471 -8816
rect 8418 -8884 8429 -8850
rect 8463 -8884 8471 -8850
rect 8418 -8927 8471 -8884
rect 8525 -8783 8578 -8763
rect 8525 -8817 8533 -8783
rect 8567 -8817 8578 -8783
rect 8525 -8851 8578 -8817
rect 8525 -8885 8533 -8851
rect 8567 -8885 8578 -8851
rect 8525 -8927 8578 -8885
rect 8678 -8782 8743 -8763
rect 8678 -8816 8689 -8782
rect 8723 -8816 8743 -8782
rect 8678 -8850 8743 -8816
rect 8678 -8884 8689 -8850
rect 8723 -8884 8743 -8850
rect 8678 -8927 8743 -8884
rect 8246 -8963 8296 -8927
rect 8693 -8963 8743 -8927
rect 8773 -8783 8844 -8763
rect 8990 -8775 9042 -8763
rect 8773 -8817 8787 -8783
rect 8821 -8817 8844 -8783
rect 8773 -8851 8844 -8817
rect 8773 -8885 8787 -8851
rect 8821 -8885 8844 -8851
rect 8773 -8963 8844 -8885
rect 8990 -8809 8998 -8775
rect 9032 -8809 9042 -8775
rect 8990 -8877 9042 -8809
rect 8990 -8911 8998 -8877
rect 9032 -8911 9042 -8877
rect 8990 -8937 9042 -8911
rect 9252 -8775 9304 -8763
rect 9252 -8809 9262 -8775
rect 9296 -8809 9304 -8775
rect 9450 -8775 9502 -8763
rect 9252 -8877 9304 -8809
rect 9252 -8911 9262 -8877
rect 9296 -8911 9304 -8877
rect 9252 -8937 9304 -8911
rect 9450 -8809 9458 -8775
rect 9492 -8809 9502 -8775
rect 9450 -8877 9502 -8809
rect 9450 -8911 9458 -8877
rect 9492 -8911 9502 -8877
rect 9450 -8937 9502 -8911
rect 10080 -8775 10132 -8763
rect 10080 -8809 10090 -8775
rect 10124 -8809 10132 -8775
rect 10370 -8775 10422 -8763
rect 10080 -8877 10132 -8809
rect 10080 -8911 10090 -8877
rect 10124 -8911 10132 -8877
rect 10080 -8937 10132 -8911
rect 10370 -8809 10378 -8775
rect 10412 -8809 10422 -8775
rect 10370 -8877 10422 -8809
rect 10370 -8911 10378 -8877
rect 10412 -8911 10422 -8877
rect 10370 -8937 10422 -8911
rect 10632 -8775 10684 -8763
rect 10632 -8809 10642 -8775
rect 10676 -8809 10684 -8775
rect 10632 -8877 10684 -8809
rect 10632 -8911 10642 -8877
rect 10676 -8911 10684 -8877
rect 10632 -8937 10684 -8911
rect 10738 -8782 10792 -8763
rect 10738 -8816 10747 -8782
rect 10781 -8816 10792 -8782
rect 10738 -8850 10792 -8816
rect 10738 -8884 10747 -8850
rect 10781 -8884 10792 -8850
rect 10738 -8963 10792 -8884
rect 10822 -8782 10894 -8763
rect 10822 -8816 10847 -8782
rect 10881 -8816 10894 -8782
rect 10822 -8850 10894 -8816
rect 10822 -8884 10847 -8850
rect 10881 -8884 10894 -8850
rect 10822 -8927 10894 -8884
rect 10994 -8782 11047 -8763
rect 10994 -8816 11005 -8782
rect 11039 -8816 11047 -8782
rect 10994 -8850 11047 -8816
rect 10994 -8884 11005 -8850
rect 11039 -8884 11047 -8850
rect 10994 -8927 11047 -8884
rect 11101 -8783 11154 -8763
rect 11101 -8817 11109 -8783
rect 11143 -8817 11154 -8783
rect 11101 -8851 11154 -8817
rect 11101 -8885 11109 -8851
rect 11143 -8885 11154 -8851
rect 11101 -8927 11154 -8885
rect 11254 -8782 11319 -8763
rect 11254 -8816 11265 -8782
rect 11299 -8816 11319 -8782
rect 11254 -8850 11319 -8816
rect 11254 -8884 11265 -8850
rect 11299 -8884 11319 -8850
rect 11254 -8927 11319 -8884
rect 10822 -8963 10872 -8927
rect 11269 -8963 11319 -8927
rect 11349 -8783 11420 -8763
rect 11658 -8775 11710 -8763
rect 11349 -8817 11363 -8783
rect 11397 -8817 11420 -8783
rect 11349 -8851 11420 -8817
rect 11349 -8885 11363 -8851
rect 11397 -8885 11420 -8851
rect 11349 -8963 11420 -8885
rect 11658 -8809 11666 -8775
rect 11700 -8809 11710 -8775
rect 11658 -8877 11710 -8809
rect 11658 -8911 11666 -8877
rect 11700 -8911 11710 -8877
rect 11658 -8937 11710 -8911
rect 11920 -8775 11972 -8763
rect 11920 -8809 11930 -8775
rect 11964 -8809 11972 -8775
rect 11920 -8877 11972 -8809
rect 11920 -8911 11930 -8877
rect 11964 -8911 11972 -8877
rect 11920 -8937 11972 -8911
rect 12486 -8782 12547 -8763
rect 12486 -8816 12502 -8782
rect 12536 -8816 12547 -8782
rect 12486 -8850 12547 -8816
rect 12486 -8884 12502 -8850
rect 12536 -8884 12547 -8850
rect 12486 -8963 12547 -8884
rect 12577 -8789 12633 -8763
rect 12577 -8823 12588 -8789
rect 12622 -8823 12633 -8789
rect 12577 -8877 12633 -8823
rect 12577 -8911 12588 -8877
rect 12622 -8911 12633 -8877
rect 12577 -8963 12633 -8911
rect 12663 -8782 12719 -8763
rect 12663 -8816 12674 -8782
rect 12708 -8816 12719 -8782
rect 12663 -8850 12719 -8816
rect 12663 -8884 12674 -8850
rect 12708 -8884 12719 -8850
rect 12663 -8963 12719 -8884
rect 12749 -8789 12805 -8763
rect 12749 -8823 12760 -8789
rect 12794 -8823 12805 -8789
rect 12749 -8877 12805 -8823
rect 12749 -8911 12760 -8877
rect 12794 -8911 12805 -8877
rect 12749 -8963 12805 -8911
rect 12835 -8782 12891 -8763
rect 12835 -8816 12846 -8782
rect 12880 -8816 12891 -8782
rect 12835 -8850 12891 -8816
rect 12835 -8884 12846 -8850
rect 12880 -8884 12891 -8850
rect 12835 -8963 12891 -8884
rect 12921 -8789 12977 -8763
rect 12921 -8823 12932 -8789
rect 12966 -8823 12977 -8789
rect 12921 -8877 12977 -8823
rect 12921 -8911 12932 -8877
rect 12966 -8911 12977 -8877
rect 12921 -8963 12977 -8911
rect 13007 -8782 13076 -8763
rect 13222 -8775 13274 -8763
rect 13007 -8816 13018 -8782
rect 13052 -8816 13076 -8782
rect 13007 -8850 13076 -8816
rect 13007 -8884 13018 -8850
rect 13052 -8884 13076 -8850
rect 13007 -8963 13076 -8884
rect 13222 -8809 13230 -8775
rect 13264 -8809 13274 -8775
rect 13222 -8877 13274 -8809
rect 13222 -8911 13230 -8877
rect 13264 -8911 13274 -8877
rect 13222 -8937 13274 -8911
rect 13484 -8775 13536 -8763
rect 13484 -8809 13494 -8775
rect 13528 -8809 13536 -8775
rect 13682 -8775 13735 -8763
rect 13484 -8877 13536 -8809
rect 13484 -8911 13494 -8877
rect 13528 -8911 13536 -8877
rect 13484 -8937 13536 -8911
rect 13682 -8809 13690 -8775
rect 13724 -8809 13735 -8775
rect 13682 -8843 13735 -8809
rect 13682 -8877 13690 -8843
rect 13724 -8877 13735 -8843
rect 13682 -8963 13735 -8877
rect 13765 -8783 13821 -8763
rect 13765 -8817 13776 -8783
rect 13810 -8817 13821 -8783
rect 13765 -8851 13821 -8817
rect 13765 -8885 13776 -8851
rect 13810 -8885 13821 -8851
rect 13765 -8963 13821 -8885
rect 13851 -8775 13907 -8763
rect 13851 -8809 13862 -8775
rect 13896 -8809 13907 -8775
rect 13851 -8843 13907 -8809
rect 13851 -8877 13862 -8843
rect 13896 -8877 13907 -8843
rect 13851 -8963 13907 -8877
rect 13937 -8791 13993 -8763
rect 13937 -8825 13948 -8791
rect 13982 -8825 13993 -8791
rect 13937 -8859 13993 -8825
rect 13937 -8893 13948 -8859
rect 13982 -8893 13993 -8859
rect 13937 -8963 13993 -8893
rect 14023 -8775 14079 -8763
rect 14023 -8809 14034 -8775
rect 14068 -8809 14079 -8775
rect 14023 -8843 14079 -8809
rect 14023 -8877 14034 -8843
rect 14068 -8877 14079 -8843
rect 14023 -8963 14079 -8877
rect 14109 -8819 14165 -8763
rect 14109 -8853 14120 -8819
rect 14154 -8853 14165 -8819
rect 14109 -8905 14165 -8853
rect 14109 -8939 14120 -8905
rect 14154 -8939 14165 -8905
rect 14109 -8963 14165 -8939
rect 14195 -8799 14251 -8763
rect 14195 -8833 14206 -8799
rect 14240 -8833 14251 -8799
rect 14195 -8963 14251 -8833
rect 14281 -8819 14337 -8763
rect 14281 -8853 14292 -8819
rect 14326 -8853 14337 -8819
rect 14281 -8905 14337 -8853
rect 14281 -8939 14292 -8905
rect 14326 -8939 14337 -8905
rect 14281 -8963 14337 -8939
rect 14367 -8799 14423 -8763
rect 14367 -8833 14378 -8799
rect 14412 -8833 14423 -8799
rect 14367 -8963 14423 -8833
rect 14453 -8819 14509 -8763
rect 14453 -8853 14464 -8819
rect 14498 -8853 14509 -8819
rect 14453 -8905 14509 -8853
rect 14453 -8939 14464 -8905
rect 14498 -8939 14509 -8905
rect 14453 -8963 14509 -8939
rect 14539 -8799 14595 -8763
rect 14539 -8833 14550 -8799
rect 14584 -8833 14595 -8799
rect 14539 -8963 14595 -8833
rect 14625 -8819 14681 -8763
rect 14625 -8853 14636 -8819
rect 14670 -8853 14681 -8819
rect 14625 -8905 14681 -8853
rect 14625 -8939 14636 -8905
rect 14670 -8939 14681 -8905
rect 14625 -8963 14681 -8939
rect 14711 -8799 14766 -8763
rect 14711 -8833 14722 -8799
rect 14756 -8833 14766 -8799
rect 14711 -8963 14766 -8833
rect 14796 -8819 14852 -8763
rect 14796 -8853 14807 -8819
rect 14841 -8853 14852 -8819
rect 14796 -8905 14852 -8853
rect 14796 -8939 14807 -8905
rect 14841 -8939 14852 -8905
rect 14796 -8963 14852 -8939
rect 14882 -8799 14938 -8763
rect 14882 -8833 14893 -8799
rect 14927 -8833 14938 -8799
rect 14882 -8963 14938 -8833
rect 14968 -8819 15024 -8763
rect 14968 -8853 14979 -8819
rect 15013 -8853 15024 -8819
rect 14968 -8905 15024 -8853
rect 14968 -8939 14979 -8905
rect 15013 -8939 15024 -8905
rect 14968 -8963 15024 -8939
rect 15054 -8799 15110 -8763
rect 15054 -8833 15065 -8799
rect 15099 -8833 15110 -8799
rect 15054 -8963 15110 -8833
rect 15140 -8819 15196 -8763
rect 15140 -8853 15151 -8819
rect 15185 -8853 15196 -8819
rect 15140 -8905 15196 -8853
rect 15140 -8939 15151 -8905
rect 15185 -8939 15196 -8905
rect 15140 -8963 15196 -8939
rect 15226 -8799 15282 -8763
rect 15226 -8833 15237 -8799
rect 15271 -8833 15282 -8799
rect 15226 -8963 15282 -8833
rect 15312 -8819 15368 -8763
rect 15312 -8853 15323 -8819
rect 15357 -8853 15368 -8819
rect 15312 -8905 15368 -8853
rect 15312 -8939 15323 -8905
rect 15357 -8939 15368 -8905
rect 15312 -8963 15368 -8939
rect 15398 -8799 15451 -8763
rect 15614 -8775 15666 -8763
rect 15398 -8833 15409 -8799
rect 15443 -8833 15451 -8799
rect 15398 -8963 15451 -8833
rect 15614 -8809 15622 -8775
rect 15656 -8809 15666 -8775
rect 15614 -8877 15666 -8809
rect 15614 -8911 15622 -8877
rect 15656 -8911 15666 -8877
rect 15614 -8937 15666 -8911
rect 16612 -8775 16664 -8763
rect 16612 -8809 16622 -8775
rect 16656 -8809 16664 -8775
rect 16612 -8877 16664 -8809
rect 16612 -8911 16622 -8877
rect 16656 -8911 16664 -8877
rect 16612 -8937 16664 -8911
rect -2970 -9609 -2918 -9583
rect -2970 -9643 -2962 -9609
rect -2928 -9643 -2918 -9609
rect -2970 -9711 -2918 -9643
rect -2970 -9745 -2962 -9711
rect -2928 -9745 -2918 -9711
rect -2970 -9757 -2918 -9745
rect -2340 -9609 -2288 -9583
rect -2340 -9643 -2330 -9609
rect -2296 -9643 -2288 -9609
rect -2340 -9711 -2288 -9643
rect -2340 -9745 -2330 -9711
rect -2296 -9745 -2288 -9711
rect -1590 -9609 -1538 -9583
rect -1590 -9643 -1582 -9609
rect -1548 -9643 -1538 -9609
rect -1590 -9711 -1538 -9643
rect -2340 -9757 -2288 -9745
rect -1590 -9745 -1582 -9711
rect -1548 -9745 -1538 -9711
rect -1590 -9757 -1538 -9745
rect -960 -9609 -908 -9583
rect -960 -9643 -950 -9609
rect -916 -9643 -908 -9609
rect -960 -9711 -908 -9643
rect -960 -9745 -950 -9711
rect -916 -9745 -908 -9711
rect -960 -9757 -908 -9745
rect -854 -9635 -783 -9557
rect -854 -9669 -831 -9635
rect -797 -9669 -783 -9635
rect -854 -9703 -783 -9669
rect -854 -9737 -831 -9703
rect -797 -9737 -783 -9703
rect -854 -9757 -783 -9737
rect -753 -9593 -703 -9557
rect -306 -9593 -256 -9557
rect -753 -9636 -688 -9593
rect -753 -9670 -733 -9636
rect -699 -9670 -688 -9636
rect -753 -9704 -688 -9670
rect -753 -9738 -733 -9704
rect -699 -9738 -688 -9704
rect -753 -9757 -688 -9738
rect -588 -9635 -535 -9593
rect -588 -9669 -577 -9635
rect -543 -9669 -535 -9635
rect -588 -9703 -535 -9669
rect -588 -9737 -577 -9703
rect -543 -9737 -535 -9703
rect -588 -9757 -535 -9737
rect -481 -9636 -428 -9593
rect -481 -9670 -473 -9636
rect -439 -9670 -428 -9636
rect -481 -9704 -428 -9670
rect -481 -9738 -473 -9704
rect -439 -9738 -428 -9704
rect -481 -9757 -428 -9738
rect -328 -9636 -256 -9593
rect -328 -9670 -315 -9636
rect -281 -9670 -256 -9636
rect -328 -9704 -256 -9670
rect -328 -9738 -315 -9704
rect -281 -9738 -256 -9704
rect -328 -9757 -256 -9738
rect -226 -9636 -172 -9557
rect -226 -9670 -215 -9636
rect -181 -9670 -172 -9636
rect -226 -9704 -172 -9670
rect -226 -9738 -215 -9704
rect -181 -9738 -172 -9704
rect -226 -9757 -172 -9738
rect -26 -9609 26 -9583
rect -26 -9643 -18 -9609
rect 16 -9643 26 -9609
rect -26 -9711 26 -9643
rect -26 -9745 -18 -9711
rect 16 -9745 26 -9711
rect -26 -9757 26 -9745
rect 236 -9609 288 -9583
rect 236 -9643 246 -9609
rect 280 -9643 288 -9609
rect 236 -9711 288 -9643
rect 236 -9745 246 -9711
rect 280 -9745 288 -9711
rect 434 -9635 505 -9557
rect 434 -9669 457 -9635
rect 491 -9669 505 -9635
rect 434 -9703 505 -9669
rect 434 -9737 457 -9703
rect 491 -9737 505 -9703
rect 236 -9757 288 -9745
rect 434 -9757 505 -9737
rect 535 -9593 585 -9557
rect 982 -9593 1032 -9557
rect 535 -9636 600 -9593
rect 535 -9670 555 -9636
rect 589 -9670 600 -9636
rect 535 -9704 600 -9670
rect 535 -9738 555 -9704
rect 589 -9738 600 -9704
rect 535 -9757 600 -9738
rect 700 -9635 753 -9593
rect 700 -9669 711 -9635
rect 745 -9669 753 -9635
rect 700 -9703 753 -9669
rect 700 -9737 711 -9703
rect 745 -9737 753 -9703
rect 700 -9757 753 -9737
rect 807 -9636 860 -9593
rect 807 -9670 815 -9636
rect 849 -9670 860 -9636
rect 807 -9704 860 -9670
rect 807 -9738 815 -9704
rect 849 -9738 860 -9704
rect 807 -9757 860 -9738
rect 960 -9636 1032 -9593
rect 960 -9670 973 -9636
rect 1007 -9670 1032 -9636
rect 960 -9704 1032 -9670
rect 960 -9738 973 -9704
rect 1007 -9738 1032 -9704
rect 960 -9757 1032 -9738
rect 1062 -9636 1116 -9557
rect 1062 -9670 1073 -9636
rect 1107 -9670 1116 -9636
rect 1062 -9704 1116 -9670
rect 1062 -9738 1073 -9704
rect 1107 -9738 1116 -9704
rect 1062 -9757 1116 -9738
rect 1262 -9609 1314 -9583
rect 1262 -9643 1270 -9609
rect 1304 -9643 1314 -9609
rect 1262 -9711 1314 -9643
rect 1262 -9745 1270 -9711
rect 1304 -9745 1314 -9711
rect 1262 -9757 1314 -9745
rect 1524 -9609 1576 -9583
rect 1524 -9643 1534 -9609
rect 1568 -9643 1576 -9609
rect 1524 -9711 1576 -9643
rect 1524 -9745 1534 -9711
rect 1568 -9745 1576 -9711
rect 1722 -9609 1774 -9583
rect 1722 -9643 1730 -9609
rect 1764 -9643 1774 -9609
rect 1722 -9711 1774 -9643
rect 1524 -9757 1576 -9745
rect 1722 -9745 1730 -9711
rect 1764 -9745 1774 -9711
rect 1722 -9757 1774 -9745
rect 2352 -9609 2404 -9583
rect 2352 -9643 2362 -9609
rect 2396 -9643 2404 -9609
rect 2352 -9711 2404 -9643
rect 2352 -9745 2362 -9711
rect 2396 -9745 2404 -9711
rect 2550 -9609 2602 -9583
rect 2550 -9643 2558 -9609
rect 2592 -9643 2602 -9609
rect 2550 -9711 2602 -9643
rect 2352 -9757 2404 -9745
rect 2550 -9745 2558 -9711
rect 2592 -9745 2602 -9711
rect 2550 -9757 2602 -9745
rect 2812 -9609 2864 -9583
rect 2812 -9643 2822 -9609
rect 2856 -9643 2864 -9609
rect 2812 -9711 2864 -9643
rect 2812 -9745 2822 -9711
rect 2856 -9745 2864 -9711
rect 3010 -9635 3081 -9557
rect 3010 -9669 3033 -9635
rect 3067 -9669 3081 -9635
rect 3010 -9703 3081 -9669
rect 3010 -9737 3033 -9703
rect 3067 -9737 3081 -9703
rect 2812 -9757 2864 -9745
rect 3010 -9757 3081 -9737
rect 3111 -9593 3161 -9557
rect 3558 -9593 3608 -9557
rect 3111 -9636 3176 -9593
rect 3111 -9670 3131 -9636
rect 3165 -9670 3176 -9636
rect 3111 -9704 3176 -9670
rect 3111 -9738 3131 -9704
rect 3165 -9738 3176 -9704
rect 3111 -9757 3176 -9738
rect 3276 -9635 3329 -9593
rect 3276 -9669 3287 -9635
rect 3321 -9669 3329 -9635
rect 3276 -9703 3329 -9669
rect 3276 -9737 3287 -9703
rect 3321 -9737 3329 -9703
rect 3276 -9757 3329 -9737
rect 3383 -9636 3436 -9593
rect 3383 -9670 3391 -9636
rect 3425 -9670 3436 -9636
rect 3383 -9704 3436 -9670
rect 3383 -9738 3391 -9704
rect 3425 -9738 3436 -9704
rect 3383 -9757 3436 -9738
rect 3536 -9636 3608 -9593
rect 3536 -9670 3549 -9636
rect 3583 -9670 3608 -9636
rect 3536 -9704 3608 -9670
rect 3536 -9738 3549 -9704
rect 3583 -9738 3608 -9704
rect 3536 -9757 3608 -9738
rect 3638 -9636 3692 -9557
rect 3638 -9670 3649 -9636
rect 3683 -9670 3692 -9636
rect 3638 -9704 3692 -9670
rect 3638 -9738 3649 -9704
rect 3683 -9738 3692 -9704
rect 3638 -9757 3692 -9738
rect 3838 -9609 3890 -9583
rect 3838 -9643 3846 -9609
rect 3880 -9643 3890 -9609
rect 3838 -9711 3890 -9643
rect 3838 -9745 3846 -9711
rect 3880 -9745 3890 -9711
rect 3838 -9757 3890 -9745
rect 4100 -9609 4152 -9583
rect 4100 -9643 4110 -9609
rect 4144 -9643 4152 -9609
rect 4100 -9711 4152 -9643
rect 4100 -9745 4110 -9711
rect 4144 -9745 4152 -9711
rect 4298 -9609 4350 -9583
rect 4298 -9643 4306 -9609
rect 4340 -9643 4350 -9609
rect 4298 -9711 4350 -9643
rect 4100 -9757 4152 -9745
rect 4298 -9745 4306 -9711
rect 4340 -9745 4350 -9711
rect 4298 -9757 4350 -9745
rect 4928 -9609 4980 -9583
rect 4928 -9643 4938 -9609
rect 4972 -9643 4980 -9609
rect 4928 -9711 4980 -9643
rect 4928 -9745 4938 -9711
rect 4972 -9745 4980 -9711
rect 5126 -9609 5178 -9583
rect 5126 -9643 5134 -9609
rect 5168 -9643 5178 -9609
rect 5126 -9711 5178 -9643
rect 4928 -9757 4980 -9745
rect 5126 -9745 5134 -9711
rect 5168 -9745 5178 -9711
rect 5126 -9757 5178 -9745
rect 5388 -9609 5440 -9583
rect 5388 -9643 5398 -9609
rect 5432 -9643 5440 -9609
rect 5388 -9711 5440 -9643
rect 5388 -9745 5398 -9711
rect 5432 -9745 5440 -9711
rect 5586 -9635 5657 -9557
rect 5586 -9669 5609 -9635
rect 5643 -9669 5657 -9635
rect 5586 -9703 5657 -9669
rect 5586 -9737 5609 -9703
rect 5643 -9737 5657 -9703
rect 5388 -9757 5440 -9745
rect 5586 -9757 5657 -9737
rect 5687 -9593 5737 -9557
rect 6134 -9593 6184 -9557
rect 5687 -9636 5752 -9593
rect 5687 -9670 5707 -9636
rect 5741 -9670 5752 -9636
rect 5687 -9704 5752 -9670
rect 5687 -9738 5707 -9704
rect 5741 -9738 5752 -9704
rect 5687 -9757 5752 -9738
rect 5852 -9635 5905 -9593
rect 5852 -9669 5863 -9635
rect 5897 -9669 5905 -9635
rect 5852 -9703 5905 -9669
rect 5852 -9737 5863 -9703
rect 5897 -9737 5905 -9703
rect 5852 -9757 5905 -9737
rect 5959 -9636 6012 -9593
rect 5959 -9670 5967 -9636
rect 6001 -9670 6012 -9636
rect 5959 -9704 6012 -9670
rect 5959 -9738 5967 -9704
rect 6001 -9738 6012 -9704
rect 5959 -9757 6012 -9738
rect 6112 -9636 6184 -9593
rect 6112 -9670 6125 -9636
rect 6159 -9670 6184 -9636
rect 6112 -9704 6184 -9670
rect 6112 -9738 6125 -9704
rect 6159 -9738 6184 -9704
rect 6112 -9757 6184 -9738
rect 6214 -9636 6268 -9557
rect 6214 -9670 6225 -9636
rect 6259 -9670 6268 -9636
rect 6214 -9704 6268 -9670
rect 6214 -9738 6225 -9704
rect 6259 -9738 6268 -9704
rect 6214 -9757 6268 -9738
rect 6414 -9609 6466 -9583
rect 6414 -9643 6422 -9609
rect 6456 -9643 6466 -9609
rect 6414 -9711 6466 -9643
rect 6414 -9745 6422 -9711
rect 6456 -9745 6466 -9711
rect 6414 -9757 6466 -9745
rect 6676 -9609 6728 -9583
rect 6676 -9643 6686 -9609
rect 6720 -9643 6728 -9609
rect 6676 -9711 6728 -9643
rect 6676 -9745 6686 -9711
rect 6720 -9745 6728 -9711
rect 6874 -9609 6926 -9583
rect 6874 -9643 6882 -9609
rect 6916 -9643 6926 -9609
rect 6874 -9711 6926 -9643
rect 6676 -9757 6728 -9745
rect 6874 -9745 6882 -9711
rect 6916 -9745 6926 -9711
rect 6874 -9757 6926 -9745
rect 7504 -9609 7556 -9583
rect 7504 -9643 7514 -9609
rect 7548 -9643 7556 -9609
rect 7504 -9711 7556 -9643
rect 7504 -9745 7514 -9711
rect 7548 -9745 7556 -9711
rect 7702 -9609 7754 -9583
rect 7702 -9643 7710 -9609
rect 7744 -9643 7754 -9609
rect 7702 -9711 7754 -9643
rect 7504 -9757 7556 -9745
rect 7702 -9745 7710 -9711
rect 7744 -9745 7754 -9711
rect 7702 -9757 7754 -9745
rect 7964 -9609 8016 -9583
rect 7964 -9643 7974 -9609
rect 8008 -9643 8016 -9609
rect 7964 -9711 8016 -9643
rect 7964 -9745 7974 -9711
rect 8008 -9745 8016 -9711
rect 8162 -9635 8233 -9557
rect 8162 -9669 8185 -9635
rect 8219 -9669 8233 -9635
rect 8162 -9703 8233 -9669
rect 8162 -9737 8185 -9703
rect 8219 -9737 8233 -9703
rect 7964 -9757 8016 -9745
rect 8162 -9757 8233 -9737
rect 8263 -9593 8313 -9557
rect 8710 -9593 8760 -9557
rect 8263 -9636 8328 -9593
rect 8263 -9670 8283 -9636
rect 8317 -9670 8328 -9636
rect 8263 -9704 8328 -9670
rect 8263 -9738 8283 -9704
rect 8317 -9738 8328 -9704
rect 8263 -9757 8328 -9738
rect 8428 -9635 8481 -9593
rect 8428 -9669 8439 -9635
rect 8473 -9669 8481 -9635
rect 8428 -9703 8481 -9669
rect 8428 -9737 8439 -9703
rect 8473 -9737 8481 -9703
rect 8428 -9757 8481 -9737
rect 8535 -9636 8588 -9593
rect 8535 -9670 8543 -9636
rect 8577 -9670 8588 -9636
rect 8535 -9704 8588 -9670
rect 8535 -9738 8543 -9704
rect 8577 -9738 8588 -9704
rect 8535 -9757 8588 -9738
rect 8688 -9636 8760 -9593
rect 8688 -9670 8701 -9636
rect 8735 -9670 8760 -9636
rect 8688 -9704 8760 -9670
rect 8688 -9738 8701 -9704
rect 8735 -9738 8760 -9704
rect 8688 -9757 8760 -9738
rect 8790 -9636 8844 -9557
rect 8790 -9670 8801 -9636
rect 8835 -9670 8844 -9636
rect 8790 -9704 8844 -9670
rect 8790 -9738 8801 -9704
rect 8835 -9738 8844 -9704
rect 8790 -9757 8844 -9738
rect 8990 -9609 9042 -9583
rect 8990 -9643 8998 -9609
rect 9032 -9643 9042 -9609
rect 8990 -9711 9042 -9643
rect 8990 -9745 8998 -9711
rect 9032 -9745 9042 -9711
rect 8990 -9757 9042 -9745
rect 9252 -9609 9304 -9583
rect 9252 -9643 9262 -9609
rect 9296 -9643 9304 -9609
rect 9252 -9711 9304 -9643
rect 9252 -9745 9262 -9711
rect 9296 -9745 9304 -9711
rect 9450 -9609 9502 -9583
rect 9450 -9643 9458 -9609
rect 9492 -9643 9502 -9609
rect 9450 -9711 9502 -9643
rect 9252 -9757 9304 -9745
rect 9450 -9745 9458 -9711
rect 9492 -9745 9502 -9711
rect 9450 -9757 9502 -9745
rect 10080 -9609 10132 -9583
rect 10080 -9643 10090 -9609
rect 10124 -9643 10132 -9609
rect 10080 -9711 10132 -9643
rect 10080 -9745 10090 -9711
rect 10124 -9745 10132 -9711
rect 10370 -9609 10422 -9583
rect 10370 -9643 10378 -9609
rect 10412 -9643 10422 -9609
rect 10370 -9711 10422 -9643
rect 10080 -9757 10132 -9745
rect 10370 -9745 10378 -9711
rect 10412 -9745 10422 -9711
rect 10370 -9757 10422 -9745
rect 10632 -9609 10684 -9583
rect 10632 -9643 10642 -9609
rect 10676 -9643 10684 -9609
rect 10632 -9711 10684 -9643
rect 10632 -9745 10642 -9711
rect 10676 -9745 10684 -9711
rect 10632 -9757 10684 -9745
rect 10738 -9635 10809 -9557
rect 10738 -9669 10761 -9635
rect 10795 -9669 10809 -9635
rect 10738 -9703 10809 -9669
rect 10738 -9737 10761 -9703
rect 10795 -9737 10809 -9703
rect 10738 -9757 10809 -9737
rect 10839 -9593 10889 -9557
rect 11286 -9593 11336 -9557
rect 10839 -9636 10904 -9593
rect 10839 -9670 10859 -9636
rect 10893 -9670 10904 -9636
rect 10839 -9704 10904 -9670
rect 10839 -9738 10859 -9704
rect 10893 -9738 10904 -9704
rect 10839 -9757 10904 -9738
rect 11004 -9635 11057 -9593
rect 11004 -9669 11015 -9635
rect 11049 -9669 11057 -9635
rect 11004 -9703 11057 -9669
rect 11004 -9737 11015 -9703
rect 11049 -9737 11057 -9703
rect 11004 -9757 11057 -9737
rect 11111 -9636 11164 -9593
rect 11111 -9670 11119 -9636
rect 11153 -9670 11164 -9636
rect 11111 -9704 11164 -9670
rect 11111 -9738 11119 -9704
rect 11153 -9738 11164 -9704
rect 11111 -9757 11164 -9738
rect 11264 -9636 11336 -9593
rect 11264 -9670 11277 -9636
rect 11311 -9670 11336 -9636
rect 11264 -9704 11336 -9670
rect 11264 -9738 11277 -9704
rect 11311 -9738 11336 -9704
rect 11264 -9757 11336 -9738
rect 11366 -9636 11420 -9557
rect 11366 -9670 11377 -9636
rect 11411 -9670 11420 -9636
rect 11366 -9704 11420 -9670
rect 11366 -9738 11377 -9704
rect 11411 -9738 11420 -9704
rect 11366 -9757 11420 -9738
rect 11658 -9609 11710 -9583
rect 11658 -9643 11666 -9609
rect 11700 -9643 11710 -9609
rect 11658 -9711 11710 -9643
rect 11658 -9745 11666 -9711
rect 11700 -9745 11710 -9711
rect 11658 -9757 11710 -9745
rect 11920 -9609 11972 -9583
rect 11920 -9643 11930 -9609
rect 11964 -9643 11972 -9609
rect 11920 -9711 11972 -9643
rect 11920 -9745 11930 -9711
rect 11964 -9745 11972 -9711
rect 13682 -9643 13735 -9557
rect 13682 -9677 13690 -9643
rect 13724 -9677 13735 -9643
rect 13682 -9711 13735 -9677
rect 11920 -9757 11972 -9745
rect 13682 -9745 13690 -9711
rect 13724 -9745 13735 -9711
rect 13682 -9757 13735 -9745
rect 13765 -9635 13821 -9557
rect 13765 -9669 13776 -9635
rect 13810 -9669 13821 -9635
rect 13765 -9703 13821 -9669
rect 13765 -9737 13776 -9703
rect 13810 -9737 13821 -9703
rect 13765 -9757 13821 -9737
rect 13851 -9643 13907 -9557
rect 13851 -9677 13862 -9643
rect 13896 -9677 13907 -9643
rect 13851 -9711 13907 -9677
rect 13851 -9745 13862 -9711
rect 13896 -9745 13907 -9711
rect 13851 -9757 13907 -9745
rect 13937 -9627 13993 -9557
rect 13937 -9661 13948 -9627
rect 13982 -9661 13993 -9627
rect 13937 -9695 13993 -9661
rect 13937 -9729 13948 -9695
rect 13982 -9729 13993 -9695
rect 13937 -9757 13993 -9729
rect 14023 -9643 14079 -9557
rect 14023 -9677 14034 -9643
rect 14068 -9677 14079 -9643
rect 14023 -9711 14079 -9677
rect 14023 -9745 14034 -9711
rect 14068 -9745 14079 -9711
rect 14023 -9757 14079 -9745
rect 14109 -9581 14165 -9557
rect 14109 -9615 14120 -9581
rect 14154 -9615 14165 -9581
rect 14109 -9667 14165 -9615
rect 14109 -9701 14120 -9667
rect 14154 -9701 14165 -9667
rect 14109 -9757 14165 -9701
rect 14195 -9687 14251 -9557
rect 14195 -9721 14206 -9687
rect 14240 -9721 14251 -9687
rect 14195 -9757 14251 -9721
rect 14281 -9581 14337 -9557
rect 14281 -9615 14292 -9581
rect 14326 -9615 14337 -9581
rect 14281 -9667 14337 -9615
rect 14281 -9701 14292 -9667
rect 14326 -9701 14337 -9667
rect 14281 -9757 14337 -9701
rect 14367 -9687 14423 -9557
rect 14367 -9721 14378 -9687
rect 14412 -9721 14423 -9687
rect 14367 -9757 14423 -9721
rect 14453 -9581 14509 -9557
rect 14453 -9615 14464 -9581
rect 14498 -9615 14509 -9581
rect 14453 -9667 14509 -9615
rect 14453 -9701 14464 -9667
rect 14498 -9701 14509 -9667
rect 14453 -9757 14509 -9701
rect 14539 -9687 14595 -9557
rect 14539 -9721 14550 -9687
rect 14584 -9721 14595 -9687
rect 14539 -9757 14595 -9721
rect 14625 -9581 14681 -9557
rect 14625 -9615 14636 -9581
rect 14670 -9615 14681 -9581
rect 14625 -9667 14681 -9615
rect 14625 -9701 14636 -9667
rect 14670 -9701 14681 -9667
rect 14625 -9757 14681 -9701
rect 14711 -9687 14766 -9557
rect 14711 -9721 14722 -9687
rect 14756 -9721 14766 -9687
rect 14711 -9757 14766 -9721
rect 14796 -9581 14852 -9557
rect 14796 -9615 14807 -9581
rect 14841 -9615 14852 -9581
rect 14796 -9667 14852 -9615
rect 14796 -9701 14807 -9667
rect 14841 -9701 14852 -9667
rect 14796 -9757 14852 -9701
rect 14882 -9687 14938 -9557
rect 14882 -9721 14893 -9687
rect 14927 -9721 14938 -9687
rect 14882 -9757 14938 -9721
rect 14968 -9581 15024 -9557
rect 14968 -9615 14979 -9581
rect 15013 -9615 15024 -9581
rect 14968 -9667 15024 -9615
rect 14968 -9701 14979 -9667
rect 15013 -9701 15024 -9667
rect 14968 -9757 15024 -9701
rect 15054 -9687 15110 -9557
rect 15054 -9721 15065 -9687
rect 15099 -9721 15110 -9687
rect 15054 -9757 15110 -9721
rect 15140 -9581 15196 -9557
rect 15140 -9615 15151 -9581
rect 15185 -9615 15196 -9581
rect 15140 -9667 15196 -9615
rect 15140 -9701 15151 -9667
rect 15185 -9701 15196 -9667
rect 15140 -9757 15196 -9701
rect 15226 -9687 15282 -9557
rect 15226 -9721 15237 -9687
rect 15271 -9721 15282 -9687
rect 15226 -9757 15282 -9721
rect 15312 -9581 15368 -9557
rect 15312 -9615 15323 -9581
rect 15357 -9615 15368 -9581
rect 15312 -9667 15368 -9615
rect 15312 -9701 15323 -9667
rect 15357 -9701 15368 -9667
rect 15312 -9757 15368 -9701
rect 15398 -9687 15451 -9557
rect 15398 -9721 15409 -9687
rect 15443 -9721 15451 -9687
rect 15398 -9757 15451 -9721
rect 15614 -9609 15666 -9583
rect 15614 -9643 15622 -9609
rect 15656 -9643 15666 -9609
rect 15614 -9711 15666 -9643
rect 15614 -9745 15622 -9711
rect 15656 -9745 15666 -9711
rect 15614 -9757 15666 -9745
rect 16612 -9609 16664 -9583
rect 16612 -9643 16622 -9609
rect 16656 -9643 16664 -9609
rect 16612 -9711 16664 -9643
rect 16612 -9745 16622 -9711
rect 16656 -9745 16664 -9711
rect 16612 -9757 16664 -9745
rect -2970 -9863 -2918 -9851
rect -2970 -9897 -2962 -9863
rect -2928 -9897 -2918 -9863
rect -2970 -9965 -2918 -9897
rect -2970 -9999 -2962 -9965
rect -2928 -9999 -2918 -9965
rect -2970 -10025 -2918 -9999
rect -2340 -9863 -2288 -9851
rect -2340 -9897 -2330 -9863
rect -2296 -9897 -2288 -9863
rect -1590 -9863 -1538 -9851
rect -2340 -9965 -2288 -9897
rect -2340 -9999 -2330 -9965
rect -2296 -9999 -2288 -9965
rect -2340 -10025 -2288 -9999
rect -1590 -9897 -1582 -9863
rect -1548 -9897 -1538 -9863
rect -1590 -9965 -1538 -9897
rect -1590 -9999 -1582 -9965
rect -1548 -9999 -1538 -9965
rect -1590 -10025 -1538 -9999
rect -960 -9863 -908 -9851
rect -960 -9897 -950 -9863
rect -916 -9897 -908 -9863
rect -960 -9965 -908 -9897
rect -960 -9999 -950 -9965
rect -916 -9999 -908 -9965
rect -960 -10025 -908 -9999
rect -854 -9863 -802 -9851
rect -854 -9897 -846 -9863
rect -812 -9897 -802 -9863
rect -854 -9965 -802 -9897
rect -854 -9999 -846 -9965
rect -812 -9999 -802 -9965
rect -854 -10025 -802 -9999
rect -224 -9863 -172 -9851
rect -224 -9897 -214 -9863
rect -180 -9897 -172 -9863
rect -26 -9863 26 -9851
rect -224 -9965 -172 -9897
rect -224 -9999 -214 -9965
rect -180 -9999 -172 -9965
rect -224 -10025 -172 -9999
rect -26 -9897 -18 -9863
rect 16 -9897 26 -9863
rect -26 -9965 26 -9897
rect -26 -9999 -18 -9965
rect 16 -9999 26 -9965
rect -26 -10025 26 -9999
rect 236 -9863 288 -9851
rect 236 -9897 246 -9863
rect 280 -9897 288 -9863
rect 236 -9965 288 -9897
rect 236 -9999 246 -9965
rect 280 -9999 288 -9965
rect 236 -10025 288 -9999
rect 434 -9870 488 -9851
rect 434 -9904 443 -9870
rect 477 -9904 488 -9870
rect 434 -9938 488 -9904
rect 434 -9972 443 -9938
rect 477 -9972 488 -9938
rect 434 -10051 488 -9972
rect 518 -9870 590 -9851
rect 518 -9904 543 -9870
rect 577 -9904 590 -9870
rect 518 -9938 590 -9904
rect 518 -9972 543 -9938
rect 577 -9972 590 -9938
rect 518 -10015 590 -9972
rect 690 -9870 743 -9851
rect 690 -9904 701 -9870
rect 735 -9904 743 -9870
rect 690 -9938 743 -9904
rect 690 -9972 701 -9938
rect 735 -9972 743 -9938
rect 690 -10015 743 -9972
rect 797 -9871 850 -9851
rect 797 -9905 805 -9871
rect 839 -9905 850 -9871
rect 797 -9939 850 -9905
rect 797 -9973 805 -9939
rect 839 -9973 850 -9939
rect 797 -10015 850 -9973
rect 950 -9870 1015 -9851
rect 950 -9904 961 -9870
rect 995 -9904 1015 -9870
rect 950 -9938 1015 -9904
rect 950 -9972 961 -9938
rect 995 -9972 1015 -9938
rect 950 -10015 1015 -9972
rect 518 -10051 568 -10015
rect 965 -10051 1015 -10015
rect 1045 -9871 1116 -9851
rect 1262 -9863 1314 -9851
rect 1045 -9905 1059 -9871
rect 1093 -9905 1116 -9871
rect 1045 -9939 1116 -9905
rect 1045 -9973 1059 -9939
rect 1093 -9973 1116 -9939
rect 1045 -10051 1116 -9973
rect 1262 -9897 1270 -9863
rect 1304 -9897 1314 -9863
rect 1262 -9965 1314 -9897
rect 1262 -9999 1270 -9965
rect 1304 -9999 1314 -9965
rect 1262 -10025 1314 -9999
rect 1524 -9863 1576 -9851
rect 1524 -9897 1534 -9863
rect 1568 -9897 1576 -9863
rect 1722 -9863 1774 -9851
rect 1524 -9965 1576 -9897
rect 1524 -9999 1534 -9965
rect 1568 -9999 1576 -9965
rect 1524 -10025 1576 -9999
rect 1722 -9897 1730 -9863
rect 1764 -9897 1774 -9863
rect 1722 -9965 1774 -9897
rect 1722 -9999 1730 -9965
rect 1764 -9999 1774 -9965
rect 1722 -10025 1774 -9999
rect 2352 -9863 2404 -9851
rect 2352 -9897 2362 -9863
rect 2396 -9897 2404 -9863
rect 2550 -9863 2602 -9851
rect 2352 -9965 2404 -9897
rect 2352 -9999 2362 -9965
rect 2396 -9999 2404 -9965
rect 2352 -10025 2404 -9999
rect 2550 -9897 2558 -9863
rect 2592 -9897 2602 -9863
rect 2550 -9965 2602 -9897
rect 2550 -9999 2558 -9965
rect 2592 -9999 2602 -9965
rect 2550 -10025 2602 -9999
rect 2812 -9863 2864 -9851
rect 2812 -9897 2822 -9863
rect 2856 -9897 2864 -9863
rect 2812 -9965 2864 -9897
rect 2812 -9999 2822 -9965
rect 2856 -9999 2864 -9965
rect 2812 -10025 2864 -9999
rect 3010 -9870 3064 -9851
rect 3010 -9904 3019 -9870
rect 3053 -9904 3064 -9870
rect 3010 -9938 3064 -9904
rect 3010 -9972 3019 -9938
rect 3053 -9972 3064 -9938
rect 3010 -10051 3064 -9972
rect 3094 -9870 3166 -9851
rect 3094 -9904 3119 -9870
rect 3153 -9904 3166 -9870
rect 3094 -9938 3166 -9904
rect 3094 -9972 3119 -9938
rect 3153 -9972 3166 -9938
rect 3094 -10015 3166 -9972
rect 3266 -9870 3319 -9851
rect 3266 -9904 3277 -9870
rect 3311 -9904 3319 -9870
rect 3266 -9938 3319 -9904
rect 3266 -9972 3277 -9938
rect 3311 -9972 3319 -9938
rect 3266 -10015 3319 -9972
rect 3373 -9871 3426 -9851
rect 3373 -9905 3381 -9871
rect 3415 -9905 3426 -9871
rect 3373 -9939 3426 -9905
rect 3373 -9973 3381 -9939
rect 3415 -9973 3426 -9939
rect 3373 -10015 3426 -9973
rect 3526 -9870 3591 -9851
rect 3526 -9904 3537 -9870
rect 3571 -9904 3591 -9870
rect 3526 -9938 3591 -9904
rect 3526 -9972 3537 -9938
rect 3571 -9972 3591 -9938
rect 3526 -10015 3591 -9972
rect 3094 -10051 3144 -10015
rect 3541 -10051 3591 -10015
rect 3621 -9871 3692 -9851
rect 3838 -9863 3890 -9851
rect 3621 -9905 3635 -9871
rect 3669 -9905 3692 -9871
rect 3621 -9939 3692 -9905
rect 3621 -9973 3635 -9939
rect 3669 -9973 3692 -9939
rect 3621 -10051 3692 -9973
rect 3838 -9897 3846 -9863
rect 3880 -9897 3890 -9863
rect 3838 -9965 3890 -9897
rect 3838 -9999 3846 -9965
rect 3880 -9999 3890 -9965
rect 3838 -10025 3890 -9999
rect 4100 -9863 4152 -9851
rect 4100 -9897 4110 -9863
rect 4144 -9897 4152 -9863
rect 4298 -9863 4350 -9851
rect 4100 -9965 4152 -9897
rect 4100 -9999 4110 -9965
rect 4144 -9999 4152 -9965
rect 4100 -10025 4152 -9999
rect 4298 -9897 4306 -9863
rect 4340 -9897 4350 -9863
rect 4298 -9965 4350 -9897
rect 4298 -9999 4306 -9965
rect 4340 -9999 4350 -9965
rect 4298 -10025 4350 -9999
rect 4928 -9863 4980 -9851
rect 4928 -9897 4938 -9863
rect 4972 -9897 4980 -9863
rect 5126 -9863 5178 -9851
rect 4928 -9965 4980 -9897
rect 4928 -9999 4938 -9965
rect 4972 -9999 4980 -9965
rect 4928 -10025 4980 -9999
rect 5126 -9897 5134 -9863
rect 5168 -9897 5178 -9863
rect 5126 -9965 5178 -9897
rect 5126 -9999 5134 -9965
rect 5168 -9999 5178 -9965
rect 5126 -10025 5178 -9999
rect 5388 -9863 5440 -9851
rect 5388 -9897 5398 -9863
rect 5432 -9897 5440 -9863
rect 5388 -9965 5440 -9897
rect 5388 -9999 5398 -9965
rect 5432 -9999 5440 -9965
rect 5388 -10025 5440 -9999
rect 5586 -9870 5640 -9851
rect 5586 -9904 5595 -9870
rect 5629 -9904 5640 -9870
rect 5586 -9938 5640 -9904
rect 5586 -9972 5595 -9938
rect 5629 -9972 5640 -9938
rect 5586 -10051 5640 -9972
rect 5670 -9870 5742 -9851
rect 5670 -9904 5695 -9870
rect 5729 -9904 5742 -9870
rect 5670 -9938 5742 -9904
rect 5670 -9972 5695 -9938
rect 5729 -9972 5742 -9938
rect 5670 -10015 5742 -9972
rect 5842 -9870 5895 -9851
rect 5842 -9904 5853 -9870
rect 5887 -9904 5895 -9870
rect 5842 -9938 5895 -9904
rect 5842 -9972 5853 -9938
rect 5887 -9972 5895 -9938
rect 5842 -10015 5895 -9972
rect 5949 -9871 6002 -9851
rect 5949 -9905 5957 -9871
rect 5991 -9905 6002 -9871
rect 5949 -9939 6002 -9905
rect 5949 -9973 5957 -9939
rect 5991 -9973 6002 -9939
rect 5949 -10015 6002 -9973
rect 6102 -9870 6167 -9851
rect 6102 -9904 6113 -9870
rect 6147 -9904 6167 -9870
rect 6102 -9938 6167 -9904
rect 6102 -9972 6113 -9938
rect 6147 -9972 6167 -9938
rect 6102 -10015 6167 -9972
rect 5670 -10051 5720 -10015
rect 6117 -10051 6167 -10015
rect 6197 -9871 6268 -9851
rect 6414 -9863 6466 -9851
rect 6197 -9905 6211 -9871
rect 6245 -9905 6268 -9871
rect 6197 -9939 6268 -9905
rect 6197 -9973 6211 -9939
rect 6245 -9973 6268 -9939
rect 6197 -10051 6268 -9973
rect 6414 -9897 6422 -9863
rect 6456 -9897 6466 -9863
rect 6414 -9965 6466 -9897
rect 6414 -9999 6422 -9965
rect 6456 -9999 6466 -9965
rect 6414 -10025 6466 -9999
rect 6676 -9863 6728 -9851
rect 6676 -9897 6686 -9863
rect 6720 -9897 6728 -9863
rect 6874 -9863 6926 -9851
rect 6676 -9965 6728 -9897
rect 6676 -9999 6686 -9965
rect 6720 -9999 6728 -9965
rect 6676 -10025 6728 -9999
rect 6874 -9897 6882 -9863
rect 6916 -9897 6926 -9863
rect 6874 -9965 6926 -9897
rect 6874 -9999 6882 -9965
rect 6916 -9999 6926 -9965
rect 6874 -10025 6926 -9999
rect 7504 -9863 7556 -9851
rect 7504 -9897 7514 -9863
rect 7548 -9897 7556 -9863
rect 7702 -9863 7754 -9851
rect 7504 -9965 7556 -9897
rect 7504 -9999 7514 -9965
rect 7548 -9999 7556 -9965
rect 7504 -10025 7556 -9999
rect 7702 -9897 7710 -9863
rect 7744 -9897 7754 -9863
rect 7702 -9965 7754 -9897
rect 7702 -9999 7710 -9965
rect 7744 -9999 7754 -9965
rect 7702 -10025 7754 -9999
rect 7964 -9863 8016 -9851
rect 7964 -9897 7974 -9863
rect 8008 -9897 8016 -9863
rect 7964 -9965 8016 -9897
rect 7964 -9999 7974 -9965
rect 8008 -9999 8016 -9965
rect 7964 -10025 8016 -9999
rect 8162 -9870 8216 -9851
rect 8162 -9904 8171 -9870
rect 8205 -9904 8216 -9870
rect 8162 -9938 8216 -9904
rect 8162 -9972 8171 -9938
rect 8205 -9972 8216 -9938
rect 8162 -10051 8216 -9972
rect 8246 -9870 8318 -9851
rect 8246 -9904 8271 -9870
rect 8305 -9904 8318 -9870
rect 8246 -9938 8318 -9904
rect 8246 -9972 8271 -9938
rect 8305 -9972 8318 -9938
rect 8246 -10015 8318 -9972
rect 8418 -9870 8471 -9851
rect 8418 -9904 8429 -9870
rect 8463 -9904 8471 -9870
rect 8418 -9938 8471 -9904
rect 8418 -9972 8429 -9938
rect 8463 -9972 8471 -9938
rect 8418 -10015 8471 -9972
rect 8525 -9871 8578 -9851
rect 8525 -9905 8533 -9871
rect 8567 -9905 8578 -9871
rect 8525 -9939 8578 -9905
rect 8525 -9973 8533 -9939
rect 8567 -9973 8578 -9939
rect 8525 -10015 8578 -9973
rect 8678 -9870 8743 -9851
rect 8678 -9904 8689 -9870
rect 8723 -9904 8743 -9870
rect 8678 -9938 8743 -9904
rect 8678 -9972 8689 -9938
rect 8723 -9972 8743 -9938
rect 8678 -10015 8743 -9972
rect 8246 -10051 8296 -10015
rect 8693 -10051 8743 -10015
rect 8773 -9871 8844 -9851
rect 8990 -9863 9042 -9851
rect 8773 -9905 8787 -9871
rect 8821 -9905 8844 -9871
rect 8773 -9939 8844 -9905
rect 8773 -9973 8787 -9939
rect 8821 -9973 8844 -9939
rect 8773 -10051 8844 -9973
rect 8990 -9897 8998 -9863
rect 9032 -9897 9042 -9863
rect 8990 -9965 9042 -9897
rect 8990 -9999 8998 -9965
rect 9032 -9999 9042 -9965
rect 8990 -10025 9042 -9999
rect 9252 -9863 9304 -9851
rect 9252 -9897 9262 -9863
rect 9296 -9897 9304 -9863
rect 9450 -9863 9502 -9851
rect 9252 -9965 9304 -9897
rect 9252 -9999 9262 -9965
rect 9296 -9999 9304 -9965
rect 9252 -10025 9304 -9999
rect 9450 -9897 9458 -9863
rect 9492 -9897 9502 -9863
rect 9450 -9965 9502 -9897
rect 9450 -9999 9458 -9965
rect 9492 -9999 9502 -9965
rect 9450 -10025 9502 -9999
rect 10080 -9863 10132 -9851
rect 10080 -9897 10090 -9863
rect 10124 -9897 10132 -9863
rect 10370 -9863 10422 -9851
rect 10080 -9965 10132 -9897
rect 10080 -9999 10090 -9965
rect 10124 -9999 10132 -9965
rect 10080 -10025 10132 -9999
rect 10370 -9897 10378 -9863
rect 10412 -9897 10422 -9863
rect 10370 -9965 10422 -9897
rect 10370 -9999 10378 -9965
rect 10412 -9999 10422 -9965
rect 10370 -10025 10422 -9999
rect 10632 -9863 10684 -9851
rect 10632 -9897 10642 -9863
rect 10676 -9897 10684 -9863
rect 10632 -9965 10684 -9897
rect 10632 -9999 10642 -9965
rect 10676 -9999 10684 -9965
rect 10632 -10025 10684 -9999
rect 10738 -9870 10792 -9851
rect 10738 -9904 10747 -9870
rect 10781 -9904 10792 -9870
rect 10738 -9938 10792 -9904
rect 10738 -9972 10747 -9938
rect 10781 -9972 10792 -9938
rect 10738 -10051 10792 -9972
rect 10822 -9870 10894 -9851
rect 10822 -9904 10847 -9870
rect 10881 -9904 10894 -9870
rect 10822 -9938 10894 -9904
rect 10822 -9972 10847 -9938
rect 10881 -9972 10894 -9938
rect 10822 -10015 10894 -9972
rect 10994 -9870 11047 -9851
rect 10994 -9904 11005 -9870
rect 11039 -9904 11047 -9870
rect 10994 -9938 11047 -9904
rect 10994 -9972 11005 -9938
rect 11039 -9972 11047 -9938
rect 10994 -10015 11047 -9972
rect 11101 -9871 11154 -9851
rect 11101 -9905 11109 -9871
rect 11143 -9905 11154 -9871
rect 11101 -9939 11154 -9905
rect 11101 -9973 11109 -9939
rect 11143 -9973 11154 -9939
rect 11101 -10015 11154 -9973
rect 11254 -9870 11319 -9851
rect 11254 -9904 11265 -9870
rect 11299 -9904 11319 -9870
rect 11254 -9938 11319 -9904
rect 11254 -9972 11265 -9938
rect 11299 -9972 11319 -9938
rect 11254 -10015 11319 -9972
rect 10822 -10051 10872 -10015
rect 11269 -10051 11319 -10015
rect 11349 -9871 11420 -9851
rect 11658 -9863 11710 -9851
rect 11349 -9905 11363 -9871
rect 11397 -9905 11420 -9871
rect 11349 -9939 11420 -9905
rect 11349 -9973 11363 -9939
rect 11397 -9973 11420 -9939
rect 11349 -10051 11420 -9973
rect 11658 -9897 11666 -9863
rect 11700 -9897 11710 -9863
rect 11658 -9965 11710 -9897
rect 11658 -9999 11666 -9965
rect 11700 -9999 11710 -9965
rect 11658 -10025 11710 -9999
rect 11920 -9863 11972 -9851
rect 11920 -9897 11930 -9863
rect 11964 -9897 11972 -9863
rect 11920 -9965 11972 -9897
rect 11920 -9999 11930 -9965
rect 11964 -9999 11972 -9965
rect 11920 -10025 11972 -9999
rect 12486 -9870 12547 -9851
rect 12486 -9904 12502 -9870
rect 12536 -9904 12547 -9870
rect 12486 -9938 12547 -9904
rect 12486 -9972 12502 -9938
rect 12536 -9972 12547 -9938
rect 12486 -10051 12547 -9972
rect 12577 -9877 12633 -9851
rect 12577 -9911 12588 -9877
rect 12622 -9911 12633 -9877
rect 12577 -9965 12633 -9911
rect 12577 -9999 12588 -9965
rect 12622 -9999 12633 -9965
rect 12577 -10051 12633 -9999
rect 12663 -9870 12719 -9851
rect 12663 -9904 12674 -9870
rect 12708 -9904 12719 -9870
rect 12663 -9938 12719 -9904
rect 12663 -9972 12674 -9938
rect 12708 -9972 12719 -9938
rect 12663 -10051 12719 -9972
rect 12749 -9877 12805 -9851
rect 12749 -9911 12760 -9877
rect 12794 -9911 12805 -9877
rect 12749 -9965 12805 -9911
rect 12749 -9999 12760 -9965
rect 12794 -9999 12805 -9965
rect 12749 -10051 12805 -9999
rect 12835 -9870 12891 -9851
rect 12835 -9904 12846 -9870
rect 12880 -9904 12891 -9870
rect 12835 -9938 12891 -9904
rect 12835 -9972 12846 -9938
rect 12880 -9972 12891 -9938
rect 12835 -10051 12891 -9972
rect 12921 -9877 12977 -9851
rect 12921 -9911 12932 -9877
rect 12966 -9911 12977 -9877
rect 12921 -9965 12977 -9911
rect 12921 -9999 12932 -9965
rect 12966 -9999 12977 -9965
rect 12921 -10051 12977 -9999
rect 13007 -9870 13076 -9851
rect 13222 -9863 13274 -9851
rect 13007 -9904 13018 -9870
rect 13052 -9904 13076 -9870
rect 13007 -9938 13076 -9904
rect 13007 -9972 13018 -9938
rect 13052 -9972 13076 -9938
rect 13007 -10051 13076 -9972
rect 13222 -9897 13230 -9863
rect 13264 -9897 13274 -9863
rect 13222 -9965 13274 -9897
rect 13222 -9999 13230 -9965
rect 13264 -9999 13274 -9965
rect 13222 -10025 13274 -9999
rect 13484 -9863 13536 -9851
rect 13484 -9897 13494 -9863
rect 13528 -9897 13536 -9863
rect 13682 -9863 13735 -9851
rect 13484 -9965 13536 -9897
rect 13484 -9999 13494 -9965
rect 13528 -9999 13536 -9965
rect 13484 -10025 13536 -9999
rect 13682 -9897 13690 -9863
rect 13724 -9897 13735 -9863
rect 13682 -9931 13735 -9897
rect 13682 -9965 13690 -9931
rect 13724 -9965 13735 -9931
rect 13682 -10051 13735 -9965
rect 13765 -9871 13821 -9851
rect 13765 -9905 13776 -9871
rect 13810 -9905 13821 -9871
rect 13765 -9939 13821 -9905
rect 13765 -9973 13776 -9939
rect 13810 -9973 13821 -9939
rect 13765 -10051 13821 -9973
rect 13851 -9863 13907 -9851
rect 13851 -9897 13862 -9863
rect 13896 -9897 13907 -9863
rect 13851 -9931 13907 -9897
rect 13851 -9965 13862 -9931
rect 13896 -9965 13907 -9931
rect 13851 -10051 13907 -9965
rect 13937 -9879 13993 -9851
rect 13937 -9913 13948 -9879
rect 13982 -9913 13993 -9879
rect 13937 -9947 13993 -9913
rect 13937 -9981 13948 -9947
rect 13982 -9981 13993 -9947
rect 13937 -10051 13993 -9981
rect 14023 -9863 14079 -9851
rect 14023 -9897 14034 -9863
rect 14068 -9897 14079 -9863
rect 14023 -9931 14079 -9897
rect 14023 -9965 14034 -9931
rect 14068 -9965 14079 -9931
rect 14023 -10051 14079 -9965
rect 14109 -9907 14165 -9851
rect 14109 -9941 14120 -9907
rect 14154 -9941 14165 -9907
rect 14109 -9993 14165 -9941
rect 14109 -10027 14120 -9993
rect 14154 -10027 14165 -9993
rect 14109 -10051 14165 -10027
rect 14195 -9887 14251 -9851
rect 14195 -9921 14206 -9887
rect 14240 -9921 14251 -9887
rect 14195 -10051 14251 -9921
rect 14281 -9907 14337 -9851
rect 14281 -9941 14292 -9907
rect 14326 -9941 14337 -9907
rect 14281 -9993 14337 -9941
rect 14281 -10027 14292 -9993
rect 14326 -10027 14337 -9993
rect 14281 -10051 14337 -10027
rect 14367 -9887 14423 -9851
rect 14367 -9921 14378 -9887
rect 14412 -9921 14423 -9887
rect 14367 -10051 14423 -9921
rect 14453 -9907 14509 -9851
rect 14453 -9941 14464 -9907
rect 14498 -9941 14509 -9907
rect 14453 -9993 14509 -9941
rect 14453 -10027 14464 -9993
rect 14498 -10027 14509 -9993
rect 14453 -10051 14509 -10027
rect 14539 -9887 14595 -9851
rect 14539 -9921 14550 -9887
rect 14584 -9921 14595 -9887
rect 14539 -10051 14595 -9921
rect 14625 -9907 14681 -9851
rect 14625 -9941 14636 -9907
rect 14670 -9941 14681 -9907
rect 14625 -9993 14681 -9941
rect 14625 -10027 14636 -9993
rect 14670 -10027 14681 -9993
rect 14625 -10051 14681 -10027
rect 14711 -9887 14766 -9851
rect 14711 -9921 14722 -9887
rect 14756 -9921 14766 -9887
rect 14711 -10051 14766 -9921
rect 14796 -9907 14852 -9851
rect 14796 -9941 14807 -9907
rect 14841 -9941 14852 -9907
rect 14796 -9993 14852 -9941
rect 14796 -10027 14807 -9993
rect 14841 -10027 14852 -9993
rect 14796 -10051 14852 -10027
rect 14882 -9887 14938 -9851
rect 14882 -9921 14893 -9887
rect 14927 -9921 14938 -9887
rect 14882 -10051 14938 -9921
rect 14968 -9907 15024 -9851
rect 14968 -9941 14979 -9907
rect 15013 -9941 15024 -9907
rect 14968 -9993 15024 -9941
rect 14968 -10027 14979 -9993
rect 15013 -10027 15024 -9993
rect 14968 -10051 15024 -10027
rect 15054 -9887 15110 -9851
rect 15054 -9921 15065 -9887
rect 15099 -9921 15110 -9887
rect 15054 -10051 15110 -9921
rect 15140 -9907 15196 -9851
rect 15140 -9941 15151 -9907
rect 15185 -9941 15196 -9907
rect 15140 -9993 15196 -9941
rect 15140 -10027 15151 -9993
rect 15185 -10027 15196 -9993
rect 15140 -10051 15196 -10027
rect 15226 -9887 15282 -9851
rect 15226 -9921 15237 -9887
rect 15271 -9921 15282 -9887
rect 15226 -10051 15282 -9921
rect 15312 -9907 15368 -9851
rect 15312 -9941 15323 -9907
rect 15357 -9941 15368 -9907
rect 15312 -9993 15368 -9941
rect 15312 -10027 15323 -9993
rect 15357 -10027 15368 -9993
rect 15312 -10051 15368 -10027
rect 15398 -9887 15451 -9851
rect 15614 -9863 15666 -9851
rect 15398 -9921 15409 -9887
rect 15443 -9921 15451 -9887
rect 15398 -10051 15451 -9921
rect 15614 -9897 15622 -9863
rect 15656 -9897 15666 -9863
rect 15614 -9965 15666 -9897
rect 15614 -9999 15622 -9965
rect 15656 -9999 15666 -9965
rect 15614 -10025 15666 -9999
rect 16612 -9863 16664 -9851
rect 16612 -9897 16622 -9863
rect 16656 -9897 16664 -9863
rect 16612 -9965 16664 -9897
rect 16612 -9999 16622 -9965
rect 16656 -9999 16664 -9965
rect 16612 -10025 16664 -9999
rect -2970 -10697 -2918 -10671
rect -2970 -10731 -2962 -10697
rect -2928 -10731 -2918 -10697
rect -2970 -10799 -2918 -10731
rect -2970 -10833 -2962 -10799
rect -2928 -10833 -2918 -10799
rect -2970 -10845 -2918 -10833
rect -2340 -10697 -2288 -10671
rect -2340 -10731 -2330 -10697
rect -2296 -10731 -2288 -10697
rect -2340 -10799 -2288 -10731
rect -2340 -10833 -2330 -10799
rect -2296 -10833 -2288 -10799
rect -1958 -10697 -1906 -10677
rect -1958 -10731 -1950 -10697
rect -1916 -10731 -1906 -10697
rect -1958 -10799 -1906 -10731
rect -2340 -10845 -2288 -10833
rect -1958 -10833 -1950 -10799
rect -1916 -10833 -1906 -10799
rect -1958 -10845 -1906 -10833
rect -1876 -10697 -1822 -10677
rect -1876 -10731 -1866 -10697
rect -1832 -10731 -1822 -10697
rect -1876 -10799 -1822 -10731
rect -1876 -10833 -1866 -10799
rect -1832 -10833 -1822 -10799
rect -1876 -10845 -1822 -10833
rect -1792 -10697 -1736 -10677
rect -1792 -10731 -1782 -10697
rect -1748 -10731 -1736 -10697
rect -1792 -10799 -1736 -10731
rect -1792 -10833 -1782 -10799
rect -1748 -10833 -1736 -10799
rect -1590 -10697 -1538 -10671
rect -1590 -10731 -1582 -10697
rect -1548 -10731 -1538 -10697
rect -1590 -10799 -1538 -10731
rect -1792 -10845 -1736 -10833
rect -1590 -10833 -1582 -10799
rect -1548 -10833 -1538 -10799
rect -1590 -10845 -1538 -10833
rect -960 -10697 -908 -10671
rect -960 -10731 -950 -10697
rect -916 -10731 -908 -10697
rect -960 -10799 -908 -10731
rect -960 -10833 -950 -10799
rect -916 -10833 -908 -10799
rect -960 -10845 -908 -10833
rect -854 -10697 -802 -10671
rect -854 -10731 -846 -10697
rect -812 -10731 -802 -10697
rect -854 -10799 -802 -10731
rect -854 -10833 -846 -10799
rect -812 -10833 -802 -10799
rect -854 -10845 -802 -10833
rect -224 -10697 -172 -10671
rect -224 -10731 -214 -10697
rect -180 -10731 -172 -10697
rect -224 -10799 -172 -10731
rect -224 -10833 -214 -10799
rect -180 -10833 -172 -10799
rect -26 -10697 26 -10671
rect -26 -10731 -18 -10697
rect 16 -10731 26 -10697
rect -26 -10799 26 -10731
rect -224 -10845 -172 -10833
rect -26 -10833 -18 -10799
rect 16 -10833 26 -10799
rect -26 -10845 26 -10833
rect 236 -10697 288 -10671
rect 236 -10731 246 -10697
rect 280 -10731 288 -10697
rect 236 -10799 288 -10731
rect 236 -10833 246 -10799
rect 280 -10833 288 -10799
rect 434 -10723 505 -10645
rect 434 -10757 457 -10723
rect 491 -10757 505 -10723
rect 434 -10791 505 -10757
rect 434 -10825 457 -10791
rect 491 -10825 505 -10791
rect 236 -10845 288 -10833
rect 434 -10845 505 -10825
rect 535 -10681 585 -10645
rect 982 -10681 1032 -10645
rect 535 -10724 600 -10681
rect 535 -10758 555 -10724
rect 589 -10758 600 -10724
rect 535 -10792 600 -10758
rect 535 -10826 555 -10792
rect 589 -10826 600 -10792
rect 535 -10845 600 -10826
rect 700 -10723 753 -10681
rect 700 -10757 711 -10723
rect 745 -10757 753 -10723
rect 700 -10791 753 -10757
rect 700 -10825 711 -10791
rect 745 -10825 753 -10791
rect 700 -10845 753 -10825
rect 807 -10724 860 -10681
rect 807 -10758 815 -10724
rect 849 -10758 860 -10724
rect 807 -10792 860 -10758
rect 807 -10826 815 -10792
rect 849 -10826 860 -10792
rect 807 -10845 860 -10826
rect 960 -10724 1032 -10681
rect 960 -10758 973 -10724
rect 1007 -10758 1032 -10724
rect 960 -10792 1032 -10758
rect 960 -10826 973 -10792
rect 1007 -10826 1032 -10792
rect 960 -10845 1032 -10826
rect 1062 -10724 1116 -10645
rect 1062 -10758 1073 -10724
rect 1107 -10758 1116 -10724
rect 1062 -10792 1116 -10758
rect 1062 -10826 1073 -10792
rect 1107 -10826 1116 -10792
rect 1062 -10845 1116 -10826
rect 1262 -10697 1314 -10671
rect 1262 -10731 1270 -10697
rect 1304 -10731 1314 -10697
rect 1262 -10799 1314 -10731
rect 1262 -10833 1270 -10799
rect 1304 -10833 1314 -10799
rect 1262 -10845 1314 -10833
rect 1524 -10697 1576 -10671
rect 1524 -10731 1534 -10697
rect 1568 -10731 1576 -10697
rect 1524 -10799 1576 -10731
rect 1524 -10833 1534 -10799
rect 1568 -10833 1576 -10799
rect 1722 -10697 1774 -10671
rect 1722 -10731 1730 -10697
rect 1764 -10731 1774 -10697
rect 1722 -10799 1774 -10731
rect 1524 -10845 1576 -10833
rect 1722 -10833 1730 -10799
rect 1764 -10833 1774 -10799
rect 1722 -10845 1774 -10833
rect 2352 -10697 2404 -10671
rect 2352 -10731 2362 -10697
rect 2396 -10731 2404 -10697
rect 2352 -10799 2404 -10731
rect 2352 -10833 2362 -10799
rect 2396 -10833 2404 -10799
rect 2550 -10697 2602 -10671
rect 2550 -10731 2558 -10697
rect 2592 -10731 2602 -10697
rect 2550 -10799 2602 -10731
rect 2352 -10845 2404 -10833
rect 2550 -10833 2558 -10799
rect 2592 -10833 2602 -10799
rect 2550 -10845 2602 -10833
rect 2812 -10697 2864 -10671
rect 2812 -10731 2822 -10697
rect 2856 -10731 2864 -10697
rect 2812 -10799 2864 -10731
rect 2812 -10833 2822 -10799
rect 2856 -10833 2864 -10799
rect 3010 -10723 3081 -10645
rect 3010 -10757 3033 -10723
rect 3067 -10757 3081 -10723
rect 3010 -10791 3081 -10757
rect 3010 -10825 3033 -10791
rect 3067 -10825 3081 -10791
rect 2812 -10845 2864 -10833
rect 3010 -10845 3081 -10825
rect 3111 -10681 3161 -10645
rect 3558 -10681 3608 -10645
rect 3111 -10724 3176 -10681
rect 3111 -10758 3131 -10724
rect 3165 -10758 3176 -10724
rect 3111 -10792 3176 -10758
rect 3111 -10826 3131 -10792
rect 3165 -10826 3176 -10792
rect 3111 -10845 3176 -10826
rect 3276 -10723 3329 -10681
rect 3276 -10757 3287 -10723
rect 3321 -10757 3329 -10723
rect 3276 -10791 3329 -10757
rect 3276 -10825 3287 -10791
rect 3321 -10825 3329 -10791
rect 3276 -10845 3329 -10825
rect 3383 -10724 3436 -10681
rect 3383 -10758 3391 -10724
rect 3425 -10758 3436 -10724
rect 3383 -10792 3436 -10758
rect 3383 -10826 3391 -10792
rect 3425 -10826 3436 -10792
rect 3383 -10845 3436 -10826
rect 3536 -10724 3608 -10681
rect 3536 -10758 3549 -10724
rect 3583 -10758 3608 -10724
rect 3536 -10792 3608 -10758
rect 3536 -10826 3549 -10792
rect 3583 -10826 3608 -10792
rect 3536 -10845 3608 -10826
rect 3638 -10724 3692 -10645
rect 3638 -10758 3649 -10724
rect 3683 -10758 3692 -10724
rect 3638 -10792 3692 -10758
rect 3638 -10826 3649 -10792
rect 3683 -10826 3692 -10792
rect 3638 -10845 3692 -10826
rect 3838 -10697 3890 -10671
rect 3838 -10731 3846 -10697
rect 3880 -10731 3890 -10697
rect 3838 -10799 3890 -10731
rect 3838 -10833 3846 -10799
rect 3880 -10833 3890 -10799
rect 3838 -10845 3890 -10833
rect 4100 -10697 4152 -10671
rect 4100 -10731 4110 -10697
rect 4144 -10731 4152 -10697
rect 4100 -10799 4152 -10731
rect 4100 -10833 4110 -10799
rect 4144 -10833 4152 -10799
rect 4298 -10697 4350 -10671
rect 4298 -10731 4306 -10697
rect 4340 -10731 4350 -10697
rect 4298 -10799 4350 -10731
rect 4100 -10845 4152 -10833
rect 4298 -10833 4306 -10799
rect 4340 -10833 4350 -10799
rect 4298 -10845 4350 -10833
rect 4928 -10697 4980 -10671
rect 4928 -10731 4938 -10697
rect 4972 -10731 4980 -10697
rect 4928 -10799 4980 -10731
rect 4928 -10833 4938 -10799
rect 4972 -10833 4980 -10799
rect 5126 -10697 5178 -10671
rect 5126 -10731 5134 -10697
rect 5168 -10731 5178 -10697
rect 5126 -10799 5178 -10731
rect 4928 -10845 4980 -10833
rect 5126 -10833 5134 -10799
rect 5168 -10833 5178 -10799
rect 5126 -10845 5178 -10833
rect 5388 -10697 5440 -10671
rect 5388 -10731 5398 -10697
rect 5432 -10731 5440 -10697
rect 5388 -10799 5440 -10731
rect 5388 -10833 5398 -10799
rect 5432 -10833 5440 -10799
rect 5586 -10723 5657 -10645
rect 5586 -10757 5609 -10723
rect 5643 -10757 5657 -10723
rect 5586 -10791 5657 -10757
rect 5586 -10825 5609 -10791
rect 5643 -10825 5657 -10791
rect 5388 -10845 5440 -10833
rect 5586 -10845 5657 -10825
rect 5687 -10681 5737 -10645
rect 6134 -10681 6184 -10645
rect 5687 -10724 5752 -10681
rect 5687 -10758 5707 -10724
rect 5741 -10758 5752 -10724
rect 5687 -10792 5752 -10758
rect 5687 -10826 5707 -10792
rect 5741 -10826 5752 -10792
rect 5687 -10845 5752 -10826
rect 5852 -10723 5905 -10681
rect 5852 -10757 5863 -10723
rect 5897 -10757 5905 -10723
rect 5852 -10791 5905 -10757
rect 5852 -10825 5863 -10791
rect 5897 -10825 5905 -10791
rect 5852 -10845 5905 -10825
rect 5959 -10724 6012 -10681
rect 5959 -10758 5967 -10724
rect 6001 -10758 6012 -10724
rect 5959 -10792 6012 -10758
rect 5959 -10826 5967 -10792
rect 6001 -10826 6012 -10792
rect 5959 -10845 6012 -10826
rect 6112 -10724 6184 -10681
rect 6112 -10758 6125 -10724
rect 6159 -10758 6184 -10724
rect 6112 -10792 6184 -10758
rect 6112 -10826 6125 -10792
rect 6159 -10826 6184 -10792
rect 6112 -10845 6184 -10826
rect 6214 -10724 6268 -10645
rect 6214 -10758 6225 -10724
rect 6259 -10758 6268 -10724
rect 6214 -10792 6268 -10758
rect 6214 -10826 6225 -10792
rect 6259 -10826 6268 -10792
rect 6214 -10845 6268 -10826
rect 6414 -10697 6466 -10671
rect 6414 -10731 6422 -10697
rect 6456 -10731 6466 -10697
rect 6414 -10799 6466 -10731
rect 6414 -10833 6422 -10799
rect 6456 -10833 6466 -10799
rect 6414 -10845 6466 -10833
rect 6676 -10697 6728 -10671
rect 6676 -10731 6686 -10697
rect 6720 -10731 6728 -10697
rect 6676 -10799 6728 -10731
rect 6676 -10833 6686 -10799
rect 6720 -10833 6728 -10799
rect 6874 -10697 6926 -10671
rect 6874 -10731 6882 -10697
rect 6916 -10731 6926 -10697
rect 6874 -10799 6926 -10731
rect 6676 -10845 6728 -10833
rect 6874 -10833 6882 -10799
rect 6916 -10833 6926 -10799
rect 6874 -10845 6926 -10833
rect 7504 -10697 7556 -10671
rect 7504 -10731 7514 -10697
rect 7548 -10731 7556 -10697
rect 7504 -10799 7556 -10731
rect 7504 -10833 7514 -10799
rect 7548 -10833 7556 -10799
rect 7702 -10697 7754 -10671
rect 7702 -10731 7710 -10697
rect 7744 -10731 7754 -10697
rect 7702 -10799 7754 -10731
rect 7504 -10845 7556 -10833
rect 7702 -10833 7710 -10799
rect 7744 -10833 7754 -10799
rect 7702 -10845 7754 -10833
rect 7964 -10697 8016 -10671
rect 7964 -10731 7974 -10697
rect 8008 -10731 8016 -10697
rect 7964 -10799 8016 -10731
rect 7964 -10833 7974 -10799
rect 8008 -10833 8016 -10799
rect 8162 -10723 8233 -10645
rect 8162 -10757 8185 -10723
rect 8219 -10757 8233 -10723
rect 8162 -10791 8233 -10757
rect 8162 -10825 8185 -10791
rect 8219 -10825 8233 -10791
rect 7964 -10845 8016 -10833
rect 8162 -10845 8233 -10825
rect 8263 -10681 8313 -10645
rect 8710 -10681 8760 -10645
rect 8263 -10724 8328 -10681
rect 8263 -10758 8283 -10724
rect 8317 -10758 8328 -10724
rect 8263 -10792 8328 -10758
rect 8263 -10826 8283 -10792
rect 8317 -10826 8328 -10792
rect 8263 -10845 8328 -10826
rect 8428 -10723 8481 -10681
rect 8428 -10757 8439 -10723
rect 8473 -10757 8481 -10723
rect 8428 -10791 8481 -10757
rect 8428 -10825 8439 -10791
rect 8473 -10825 8481 -10791
rect 8428 -10845 8481 -10825
rect 8535 -10724 8588 -10681
rect 8535 -10758 8543 -10724
rect 8577 -10758 8588 -10724
rect 8535 -10792 8588 -10758
rect 8535 -10826 8543 -10792
rect 8577 -10826 8588 -10792
rect 8535 -10845 8588 -10826
rect 8688 -10724 8760 -10681
rect 8688 -10758 8701 -10724
rect 8735 -10758 8760 -10724
rect 8688 -10792 8760 -10758
rect 8688 -10826 8701 -10792
rect 8735 -10826 8760 -10792
rect 8688 -10845 8760 -10826
rect 8790 -10724 8844 -10645
rect 8790 -10758 8801 -10724
rect 8835 -10758 8844 -10724
rect 8790 -10792 8844 -10758
rect 8790 -10826 8801 -10792
rect 8835 -10826 8844 -10792
rect 8790 -10845 8844 -10826
rect 8990 -10697 9042 -10671
rect 8990 -10731 8998 -10697
rect 9032 -10731 9042 -10697
rect 8990 -10799 9042 -10731
rect 8990 -10833 8998 -10799
rect 9032 -10833 9042 -10799
rect 8990 -10845 9042 -10833
rect 9252 -10697 9304 -10671
rect 9252 -10731 9262 -10697
rect 9296 -10731 9304 -10697
rect 9252 -10799 9304 -10731
rect 9252 -10833 9262 -10799
rect 9296 -10833 9304 -10799
rect 9450 -10697 9502 -10671
rect 9450 -10731 9458 -10697
rect 9492 -10731 9502 -10697
rect 9450 -10799 9502 -10731
rect 9252 -10845 9304 -10833
rect 9450 -10833 9458 -10799
rect 9492 -10833 9502 -10799
rect 9450 -10845 9502 -10833
rect 10080 -10697 10132 -10671
rect 10080 -10731 10090 -10697
rect 10124 -10731 10132 -10697
rect 10080 -10799 10132 -10731
rect 10080 -10833 10090 -10799
rect 10124 -10833 10132 -10799
rect 10370 -10697 10422 -10671
rect 10370 -10731 10378 -10697
rect 10412 -10731 10422 -10697
rect 10370 -10799 10422 -10731
rect 10080 -10845 10132 -10833
rect 10370 -10833 10378 -10799
rect 10412 -10833 10422 -10799
rect 10370 -10845 10422 -10833
rect 10632 -10697 10684 -10671
rect 10632 -10731 10642 -10697
rect 10676 -10731 10684 -10697
rect 10632 -10799 10684 -10731
rect 10632 -10833 10642 -10799
rect 10676 -10833 10684 -10799
rect 10632 -10845 10684 -10833
rect 10738 -10723 10809 -10645
rect 10738 -10757 10761 -10723
rect 10795 -10757 10809 -10723
rect 10738 -10791 10809 -10757
rect 10738 -10825 10761 -10791
rect 10795 -10825 10809 -10791
rect 10738 -10845 10809 -10825
rect 10839 -10681 10889 -10645
rect 11286 -10681 11336 -10645
rect 10839 -10724 10904 -10681
rect 10839 -10758 10859 -10724
rect 10893 -10758 10904 -10724
rect 10839 -10792 10904 -10758
rect 10839 -10826 10859 -10792
rect 10893 -10826 10904 -10792
rect 10839 -10845 10904 -10826
rect 11004 -10723 11057 -10681
rect 11004 -10757 11015 -10723
rect 11049 -10757 11057 -10723
rect 11004 -10791 11057 -10757
rect 11004 -10825 11015 -10791
rect 11049 -10825 11057 -10791
rect 11004 -10845 11057 -10825
rect 11111 -10724 11164 -10681
rect 11111 -10758 11119 -10724
rect 11153 -10758 11164 -10724
rect 11111 -10792 11164 -10758
rect 11111 -10826 11119 -10792
rect 11153 -10826 11164 -10792
rect 11111 -10845 11164 -10826
rect 11264 -10724 11336 -10681
rect 11264 -10758 11277 -10724
rect 11311 -10758 11336 -10724
rect 11264 -10792 11336 -10758
rect 11264 -10826 11277 -10792
rect 11311 -10826 11336 -10792
rect 11264 -10845 11336 -10826
rect 11366 -10724 11420 -10645
rect 11366 -10758 11377 -10724
rect 11411 -10758 11420 -10724
rect 11366 -10792 11420 -10758
rect 11366 -10826 11377 -10792
rect 11411 -10826 11420 -10792
rect 11366 -10845 11420 -10826
rect 11658 -10697 11710 -10671
rect 11658 -10731 11666 -10697
rect 11700 -10731 11710 -10697
rect 11658 -10799 11710 -10731
rect 11658 -10833 11666 -10799
rect 11700 -10833 11710 -10799
rect 11658 -10845 11710 -10833
rect 11920 -10697 11972 -10671
rect 11920 -10731 11930 -10697
rect 11964 -10731 11972 -10697
rect 11920 -10799 11972 -10731
rect 11920 -10833 11930 -10799
rect 11964 -10833 11972 -10799
rect 13590 -10697 13642 -10671
rect 13590 -10731 13598 -10697
rect 13632 -10731 13642 -10697
rect 13590 -10799 13642 -10731
rect 11920 -10845 11972 -10833
rect 13590 -10833 13598 -10799
rect 13632 -10833 13642 -10799
rect 13590 -10845 13642 -10833
rect 14588 -10697 14640 -10671
rect 14588 -10731 14598 -10697
rect 14632 -10731 14640 -10697
rect 14588 -10799 14640 -10731
rect 14588 -10833 14598 -10799
rect 14632 -10833 14640 -10799
rect 14786 -10697 14838 -10671
rect 14786 -10731 14794 -10697
rect 14828 -10731 14838 -10697
rect 14786 -10799 14838 -10731
rect 14588 -10845 14640 -10833
rect 14786 -10833 14794 -10799
rect 14828 -10833 14838 -10799
rect 14786 -10845 14838 -10833
rect 15784 -10697 15836 -10671
rect 15784 -10731 15794 -10697
rect 15828 -10731 15836 -10697
rect 15784 -10799 15836 -10731
rect 15784 -10833 15794 -10799
rect 15828 -10833 15836 -10799
rect 15982 -10697 16034 -10671
rect 15982 -10731 15990 -10697
rect 16024 -10731 16034 -10697
rect 15982 -10799 16034 -10731
rect 15784 -10845 15836 -10833
rect 15982 -10833 15990 -10799
rect 16024 -10833 16034 -10799
rect 15982 -10845 16034 -10833
rect 16612 -10697 16664 -10671
rect 16612 -10731 16622 -10697
rect 16656 -10731 16664 -10697
rect 16612 -10799 16664 -10731
rect 16612 -10833 16622 -10799
rect 16656 -10833 16664 -10799
rect 16612 -10845 16664 -10833
rect -2970 -10951 -2918 -10939
rect -2970 -10985 -2962 -10951
rect -2928 -10985 -2918 -10951
rect -2970 -11053 -2918 -10985
rect -2970 -11087 -2962 -11053
rect -2928 -11087 -2918 -11053
rect -2970 -11113 -2918 -11087
rect -2340 -10951 -2288 -10939
rect -2340 -10985 -2330 -10951
rect -2296 -10985 -2288 -10951
rect -1590 -10951 -1538 -10939
rect -2340 -11053 -2288 -10985
rect -2340 -11087 -2330 -11053
rect -2296 -11087 -2288 -11053
rect -2340 -11113 -2288 -11087
rect -1590 -10985 -1582 -10951
rect -1548 -10985 -1538 -10951
rect -1590 -11053 -1538 -10985
rect -1590 -11087 -1582 -11053
rect -1548 -11087 -1538 -11053
rect -1590 -11113 -1538 -11087
rect -960 -10951 -908 -10939
rect -960 -10985 -950 -10951
rect -916 -10985 -908 -10951
rect -960 -11053 -908 -10985
rect -960 -11087 -950 -11053
rect -916 -11087 -908 -11053
rect -960 -11113 -908 -11087
rect -854 -10951 -802 -10939
rect -854 -10985 -846 -10951
rect -812 -10985 -802 -10951
rect -854 -11053 -802 -10985
rect -854 -11087 -846 -11053
rect -812 -11087 -802 -11053
rect -854 -11113 -802 -11087
rect -224 -10951 -172 -10939
rect -224 -10985 -214 -10951
rect -180 -10985 -172 -10951
rect -26 -10951 26 -10939
rect -224 -11053 -172 -10985
rect -224 -11087 -214 -11053
rect -180 -11087 -172 -11053
rect -224 -11113 -172 -11087
rect -26 -10985 -18 -10951
rect 16 -10985 26 -10951
rect -26 -11053 26 -10985
rect -26 -11087 -18 -11053
rect 16 -11087 26 -11053
rect -26 -11113 26 -11087
rect 236 -10951 288 -10939
rect 236 -10985 246 -10951
rect 280 -10985 288 -10951
rect 236 -11053 288 -10985
rect 236 -11087 246 -11053
rect 280 -11087 288 -11053
rect 236 -11113 288 -11087
rect 434 -10959 505 -10939
rect 434 -10993 457 -10959
rect 491 -10993 505 -10959
rect 434 -11027 505 -10993
rect 434 -11061 457 -11027
rect 491 -11061 505 -11027
rect 434 -11139 505 -11061
rect 535 -10958 600 -10939
rect 535 -10992 555 -10958
rect 589 -10992 600 -10958
rect 535 -11026 600 -10992
rect 535 -11060 555 -11026
rect 589 -11060 600 -11026
rect 535 -11103 600 -11060
rect 700 -10959 753 -10939
rect 700 -10993 711 -10959
rect 745 -10993 753 -10959
rect 700 -11027 753 -10993
rect 700 -11061 711 -11027
rect 745 -11061 753 -11027
rect 700 -11103 753 -11061
rect 807 -10958 860 -10939
rect 807 -10992 815 -10958
rect 849 -10992 860 -10958
rect 807 -11026 860 -10992
rect 807 -11060 815 -11026
rect 849 -11060 860 -11026
rect 807 -11103 860 -11060
rect 960 -10958 1032 -10939
rect 960 -10992 973 -10958
rect 1007 -10992 1032 -10958
rect 960 -11026 1032 -10992
rect 960 -11060 973 -11026
rect 1007 -11060 1032 -11026
rect 960 -11103 1032 -11060
rect 535 -11139 585 -11103
rect 982 -11139 1032 -11103
rect 1062 -10958 1116 -10939
rect 1262 -10951 1314 -10939
rect 1062 -10992 1073 -10958
rect 1107 -10992 1116 -10958
rect 1062 -11026 1116 -10992
rect 1062 -11060 1073 -11026
rect 1107 -11060 1116 -11026
rect 1062 -11139 1116 -11060
rect 1262 -10985 1270 -10951
rect 1304 -10985 1314 -10951
rect 1262 -11053 1314 -10985
rect 1262 -11087 1270 -11053
rect 1304 -11087 1314 -11053
rect 1262 -11113 1314 -11087
rect 1524 -10951 1576 -10939
rect 1524 -10985 1534 -10951
rect 1568 -10985 1576 -10951
rect 1722 -10951 1774 -10939
rect 1524 -11053 1576 -10985
rect 1524 -11087 1534 -11053
rect 1568 -11087 1576 -11053
rect 1524 -11113 1576 -11087
rect 1722 -10985 1730 -10951
rect 1764 -10985 1774 -10951
rect 1722 -11053 1774 -10985
rect 1722 -11087 1730 -11053
rect 1764 -11087 1774 -11053
rect 1722 -11113 1774 -11087
rect 2352 -10951 2404 -10939
rect 2352 -10985 2362 -10951
rect 2396 -10985 2404 -10951
rect 2550 -10951 2602 -10939
rect 2352 -11053 2404 -10985
rect 2352 -11087 2362 -11053
rect 2396 -11087 2404 -11053
rect 2352 -11113 2404 -11087
rect 2550 -10985 2558 -10951
rect 2592 -10985 2602 -10951
rect 2550 -11053 2602 -10985
rect 2550 -11087 2558 -11053
rect 2592 -11087 2602 -11053
rect 2550 -11113 2602 -11087
rect 2812 -10951 2864 -10939
rect 2812 -10985 2822 -10951
rect 2856 -10985 2864 -10951
rect 2812 -11053 2864 -10985
rect 2812 -11087 2822 -11053
rect 2856 -11087 2864 -11053
rect 2812 -11113 2864 -11087
rect 3010 -10959 3081 -10939
rect 3010 -10993 3033 -10959
rect 3067 -10993 3081 -10959
rect 3010 -11027 3081 -10993
rect 3010 -11061 3033 -11027
rect 3067 -11061 3081 -11027
rect 3010 -11139 3081 -11061
rect 3111 -10958 3176 -10939
rect 3111 -10992 3131 -10958
rect 3165 -10992 3176 -10958
rect 3111 -11026 3176 -10992
rect 3111 -11060 3131 -11026
rect 3165 -11060 3176 -11026
rect 3111 -11103 3176 -11060
rect 3276 -10959 3329 -10939
rect 3276 -10993 3287 -10959
rect 3321 -10993 3329 -10959
rect 3276 -11027 3329 -10993
rect 3276 -11061 3287 -11027
rect 3321 -11061 3329 -11027
rect 3276 -11103 3329 -11061
rect 3383 -10958 3436 -10939
rect 3383 -10992 3391 -10958
rect 3425 -10992 3436 -10958
rect 3383 -11026 3436 -10992
rect 3383 -11060 3391 -11026
rect 3425 -11060 3436 -11026
rect 3383 -11103 3436 -11060
rect 3536 -10958 3608 -10939
rect 3536 -10992 3549 -10958
rect 3583 -10992 3608 -10958
rect 3536 -11026 3608 -10992
rect 3536 -11060 3549 -11026
rect 3583 -11060 3608 -11026
rect 3536 -11103 3608 -11060
rect 3111 -11139 3161 -11103
rect 3558 -11139 3608 -11103
rect 3638 -10958 3692 -10939
rect 3838 -10951 3890 -10939
rect 3638 -10992 3649 -10958
rect 3683 -10992 3692 -10958
rect 3638 -11026 3692 -10992
rect 3638 -11060 3649 -11026
rect 3683 -11060 3692 -11026
rect 3638 -11139 3692 -11060
rect 3838 -10985 3846 -10951
rect 3880 -10985 3890 -10951
rect 3838 -11053 3890 -10985
rect 3838 -11087 3846 -11053
rect 3880 -11087 3890 -11053
rect 3838 -11113 3890 -11087
rect 4100 -10951 4152 -10939
rect 4100 -10985 4110 -10951
rect 4144 -10985 4152 -10951
rect 4298 -10951 4350 -10939
rect 4100 -11053 4152 -10985
rect 4100 -11087 4110 -11053
rect 4144 -11087 4152 -11053
rect 4100 -11113 4152 -11087
rect 4298 -10985 4306 -10951
rect 4340 -10985 4350 -10951
rect 4298 -11053 4350 -10985
rect 4298 -11087 4306 -11053
rect 4340 -11087 4350 -11053
rect 4298 -11113 4350 -11087
rect 4928 -10951 4980 -10939
rect 4928 -10985 4938 -10951
rect 4972 -10985 4980 -10951
rect 5126 -10951 5178 -10939
rect 4928 -11053 4980 -10985
rect 4928 -11087 4938 -11053
rect 4972 -11087 4980 -11053
rect 4928 -11113 4980 -11087
rect 5126 -10985 5134 -10951
rect 5168 -10985 5178 -10951
rect 5126 -11053 5178 -10985
rect 5126 -11087 5134 -11053
rect 5168 -11087 5178 -11053
rect 5126 -11113 5178 -11087
rect 5388 -10951 5440 -10939
rect 5388 -10985 5398 -10951
rect 5432 -10985 5440 -10951
rect 5388 -11053 5440 -10985
rect 5388 -11087 5398 -11053
rect 5432 -11087 5440 -11053
rect 5388 -11113 5440 -11087
rect 5586 -10959 5657 -10939
rect 5586 -10993 5609 -10959
rect 5643 -10993 5657 -10959
rect 5586 -11027 5657 -10993
rect 5586 -11061 5609 -11027
rect 5643 -11061 5657 -11027
rect 5586 -11139 5657 -11061
rect 5687 -10958 5752 -10939
rect 5687 -10992 5707 -10958
rect 5741 -10992 5752 -10958
rect 5687 -11026 5752 -10992
rect 5687 -11060 5707 -11026
rect 5741 -11060 5752 -11026
rect 5687 -11103 5752 -11060
rect 5852 -10959 5905 -10939
rect 5852 -10993 5863 -10959
rect 5897 -10993 5905 -10959
rect 5852 -11027 5905 -10993
rect 5852 -11061 5863 -11027
rect 5897 -11061 5905 -11027
rect 5852 -11103 5905 -11061
rect 5959 -10958 6012 -10939
rect 5959 -10992 5967 -10958
rect 6001 -10992 6012 -10958
rect 5959 -11026 6012 -10992
rect 5959 -11060 5967 -11026
rect 6001 -11060 6012 -11026
rect 5959 -11103 6012 -11060
rect 6112 -10958 6184 -10939
rect 6112 -10992 6125 -10958
rect 6159 -10992 6184 -10958
rect 6112 -11026 6184 -10992
rect 6112 -11060 6125 -11026
rect 6159 -11060 6184 -11026
rect 6112 -11103 6184 -11060
rect 5687 -11139 5737 -11103
rect 6134 -11139 6184 -11103
rect 6214 -10958 6268 -10939
rect 6414 -10951 6466 -10939
rect 6214 -10992 6225 -10958
rect 6259 -10992 6268 -10958
rect 6214 -11026 6268 -10992
rect 6214 -11060 6225 -11026
rect 6259 -11060 6268 -11026
rect 6214 -11139 6268 -11060
rect 6414 -10985 6422 -10951
rect 6456 -10985 6466 -10951
rect 6414 -11053 6466 -10985
rect 6414 -11087 6422 -11053
rect 6456 -11087 6466 -11053
rect 6414 -11113 6466 -11087
rect 6676 -10951 6728 -10939
rect 6676 -10985 6686 -10951
rect 6720 -10985 6728 -10951
rect 6874 -10951 6926 -10939
rect 6676 -11053 6728 -10985
rect 6676 -11087 6686 -11053
rect 6720 -11087 6728 -11053
rect 6676 -11113 6728 -11087
rect 6874 -10985 6882 -10951
rect 6916 -10985 6926 -10951
rect 6874 -11053 6926 -10985
rect 6874 -11087 6882 -11053
rect 6916 -11087 6926 -11053
rect 6874 -11113 6926 -11087
rect 7504 -10951 7556 -10939
rect 7504 -10985 7514 -10951
rect 7548 -10985 7556 -10951
rect 7702 -10951 7754 -10939
rect 7504 -11053 7556 -10985
rect 7504 -11087 7514 -11053
rect 7548 -11087 7556 -11053
rect 7504 -11113 7556 -11087
rect 7702 -10985 7710 -10951
rect 7744 -10985 7754 -10951
rect 7702 -11053 7754 -10985
rect 7702 -11087 7710 -11053
rect 7744 -11087 7754 -11053
rect 7702 -11113 7754 -11087
rect 7964 -10951 8016 -10939
rect 7964 -10985 7974 -10951
rect 8008 -10985 8016 -10951
rect 7964 -11053 8016 -10985
rect 7964 -11087 7974 -11053
rect 8008 -11087 8016 -11053
rect 7964 -11113 8016 -11087
rect 8162 -10959 8233 -10939
rect 8162 -10993 8185 -10959
rect 8219 -10993 8233 -10959
rect 8162 -11027 8233 -10993
rect 8162 -11061 8185 -11027
rect 8219 -11061 8233 -11027
rect 8162 -11139 8233 -11061
rect 8263 -10958 8328 -10939
rect 8263 -10992 8283 -10958
rect 8317 -10992 8328 -10958
rect 8263 -11026 8328 -10992
rect 8263 -11060 8283 -11026
rect 8317 -11060 8328 -11026
rect 8263 -11103 8328 -11060
rect 8428 -10959 8481 -10939
rect 8428 -10993 8439 -10959
rect 8473 -10993 8481 -10959
rect 8428 -11027 8481 -10993
rect 8428 -11061 8439 -11027
rect 8473 -11061 8481 -11027
rect 8428 -11103 8481 -11061
rect 8535 -10958 8588 -10939
rect 8535 -10992 8543 -10958
rect 8577 -10992 8588 -10958
rect 8535 -11026 8588 -10992
rect 8535 -11060 8543 -11026
rect 8577 -11060 8588 -11026
rect 8535 -11103 8588 -11060
rect 8688 -10958 8760 -10939
rect 8688 -10992 8701 -10958
rect 8735 -10992 8760 -10958
rect 8688 -11026 8760 -10992
rect 8688 -11060 8701 -11026
rect 8735 -11060 8760 -11026
rect 8688 -11103 8760 -11060
rect 8263 -11139 8313 -11103
rect 8710 -11139 8760 -11103
rect 8790 -10958 8844 -10939
rect 8990 -10951 9042 -10939
rect 8790 -10992 8801 -10958
rect 8835 -10992 8844 -10958
rect 8790 -11026 8844 -10992
rect 8790 -11060 8801 -11026
rect 8835 -11060 8844 -11026
rect 8790 -11139 8844 -11060
rect 8990 -10985 8998 -10951
rect 9032 -10985 9042 -10951
rect 8990 -11053 9042 -10985
rect 8990 -11087 8998 -11053
rect 9032 -11087 9042 -11053
rect 8990 -11113 9042 -11087
rect 9252 -10951 9304 -10939
rect 9252 -10985 9262 -10951
rect 9296 -10985 9304 -10951
rect 9450 -10951 9502 -10939
rect 9252 -11053 9304 -10985
rect 9252 -11087 9262 -11053
rect 9296 -11087 9304 -11053
rect 9252 -11113 9304 -11087
rect 9450 -10985 9458 -10951
rect 9492 -10985 9502 -10951
rect 9450 -11053 9502 -10985
rect 9450 -11087 9458 -11053
rect 9492 -11087 9502 -11053
rect 9450 -11113 9502 -11087
rect 10080 -10951 10132 -10939
rect 10080 -10985 10090 -10951
rect 10124 -10985 10132 -10951
rect 10370 -10951 10422 -10939
rect 10080 -11053 10132 -10985
rect 10080 -11087 10090 -11053
rect 10124 -11087 10132 -11053
rect 10080 -11113 10132 -11087
rect 10370 -10985 10378 -10951
rect 10412 -10985 10422 -10951
rect 10370 -11053 10422 -10985
rect 10370 -11087 10378 -11053
rect 10412 -11087 10422 -11053
rect 10370 -11113 10422 -11087
rect 10632 -10951 10684 -10939
rect 10632 -10985 10642 -10951
rect 10676 -10985 10684 -10951
rect 10632 -11053 10684 -10985
rect 10632 -11087 10642 -11053
rect 10676 -11087 10684 -11053
rect 10632 -11113 10684 -11087
rect 10738 -10959 10809 -10939
rect 10738 -10993 10761 -10959
rect 10795 -10993 10809 -10959
rect 10738 -11027 10809 -10993
rect 10738 -11061 10761 -11027
rect 10795 -11061 10809 -11027
rect 10738 -11139 10809 -11061
rect 10839 -10958 10904 -10939
rect 10839 -10992 10859 -10958
rect 10893 -10992 10904 -10958
rect 10839 -11026 10904 -10992
rect 10839 -11060 10859 -11026
rect 10893 -11060 10904 -11026
rect 10839 -11103 10904 -11060
rect 11004 -10959 11057 -10939
rect 11004 -10993 11015 -10959
rect 11049 -10993 11057 -10959
rect 11004 -11027 11057 -10993
rect 11004 -11061 11015 -11027
rect 11049 -11061 11057 -11027
rect 11004 -11103 11057 -11061
rect 11111 -10958 11164 -10939
rect 11111 -10992 11119 -10958
rect 11153 -10992 11164 -10958
rect 11111 -11026 11164 -10992
rect 11111 -11060 11119 -11026
rect 11153 -11060 11164 -11026
rect 11111 -11103 11164 -11060
rect 11264 -10958 11336 -10939
rect 11264 -10992 11277 -10958
rect 11311 -10992 11336 -10958
rect 11264 -11026 11336 -10992
rect 11264 -11060 11277 -11026
rect 11311 -11060 11336 -11026
rect 11264 -11103 11336 -11060
rect 10839 -11139 10889 -11103
rect 11286 -11139 11336 -11103
rect 11366 -10958 11420 -10939
rect 11658 -10951 11710 -10939
rect 11366 -10992 11377 -10958
rect 11411 -10992 11420 -10958
rect 11366 -11026 11420 -10992
rect 11366 -11060 11377 -11026
rect 11411 -11060 11420 -11026
rect 11366 -11139 11420 -11060
rect 11658 -10985 11666 -10951
rect 11700 -10985 11710 -10951
rect 11658 -11053 11710 -10985
rect 11658 -11087 11666 -11053
rect 11700 -11087 11710 -11053
rect 11658 -11113 11710 -11087
rect 11920 -10951 11972 -10939
rect 11920 -10985 11930 -10951
rect 11964 -10985 11972 -10951
rect 13590 -10951 13642 -10939
rect 11920 -11053 11972 -10985
rect 11920 -11087 11930 -11053
rect 11964 -11087 11972 -11053
rect 11920 -11113 11972 -11087
rect 13590 -10985 13598 -10951
rect 13632 -10985 13642 -10951
rect 13590 -11053 13642 -10985
rect 13590 -11087 13598 -11053
rect 13632 -11087 13642 -11053
rect 13590 -11113 13642 -11087
rect 14588 -10951 14640 -10939
rect 14588 -10985 14598 -10951
rect 14632 -10985 14640 -10951
rect 14786 -10951 14838 -10939
rect 14588 -11053 14640 -10985
rect 14588 -11087 14598 -11053
rect 14632 -11087 14640 -11053
rect 14588 -11113 14640 -11087
rect 14786 -10985 14794 -10951
rect 14828 -10985 14838 -10951
rect 14786 -11053 14838 -10985
rect 14786 -11087 14794 -11053
rect 14828 -11087 14838 -11053
rect 14786 -11113 14838 -11087
rect 15784 -10951 15836 -10939
rect 15784 -10985 15794 -10951
rect 15828 -10985 15836 -10951
rect 15982 -10951 16034 -10939
rect 15784 -11053 15836 -10985
rect 15784 -11087 15794 -11053
rect 15828 -11087 15836 -11053
rect 15784 -11113 15836 -11087
rect 15982 -10985 15990 -10951
rect 16024 -10985 16034 -10951
rect 15982 -11053 16034 -10985
rect 15982 -11087 15990 -11053
rect 16024 -11087 16034 -11053
rect 15982 -11113 16034 -11087
rect 16612 -10951 16664 -10939
rect 16612 -10985 16622 -10951
rect 16656 -10985 16664 -10951
rect 16612 -11053 16664 -10985
rect 16612 -11087 16622 -11053
rect 16656 -11087 16664 -11053
rect 16612 -11113 16664 -11087
rect -2970 -11785 -2918 -11759
rect -2970 -11819 -2962 -11785
rect -2928 -11819 -2918 -11785
rect -2970 -11887 -2918 -11819
rect -2970 -11921 -2962 -11887
rect -2928 -11921 -2918 -11887
rect -2970 -11933 -2918 -11921
rect -2340 -11785 -2288 -11759
rect -2340 -11819 -2330 -11785
rect -2296 -11819 -2288 -11785
rect -2340 -11887 -2288 -11819
rect -2340 -11921 -2330 -11887
rect -2296 -11921 -2288 -11887
rect -1590 -11785 -1538 -11759
rect -1590 -11819 -1582 -11785
rect -1548 -11819 -1538 -11785
rect -1590 -11887 -1538 -11819
rect -2340 -11933 -2288 -11921
rect -1590 -11921 -1582 -11887
rect -1548 -11921 -1538 -11887
rect -1590 -11933 -1538 -11921
rect -960 -11785 -908 -11759
rect -960 -11819 -950 -11785
rect -916 -11819 -908 -11785
rect -960 -11887 -908 -11819
rect -960 -11921 -950 -11887
rect -916 -11921 -908 -11887
rect -960 -11933 -908 -11921
rect -854 -11785 -802 -11759
rect -854 -11819 -846 -11785
rect -812 -11819 -802 -11785
rect -854 -11887 -802 -11819
rect -854 -11921 -846 -11887
rect -812 -11921 -802 -11887
rect -854 -11933 -802 -11921
rect -224 -11785 -172 -11759
rect -224 -11819 -214 -11785
rect -180 -11819 -172 -11785
rect -224 -11887 -172 -11819
rect -224 -11921 -214 -11887
rect -180 -11921 -172 -11887
rect -26 -11785 26 -11759
rect -26 -11819 -18 -11785
rect 16 -11819 26 -11785
rect -26 -11887 26 -11819
rect -224 -11933 -172 -11921
rect -26 -11921 -18 -11887
rect 16 -11921 26 -11887
rect -26 -11933 26 -11921
rect 236 -11785 288 -11759
rect 236 -11819 246 -11785
rect 280 -11819 288 -11785
rect 236 -11887 288 -11819
rect 236 -11921 246 -11887
rect 280 -11921 288 -11887
rect 434 -11812 488 -11733
rect 434 -11846 443 -11812
rect 477 -11846 488 -11812
rect 434 -11880 488 -11846
rect 434 -11914 443 -11880
rect 477 -11914 488 -11880
rect 236 -11933 288 -11921
rect 434 -11933 488 -11914
rect 518 -11769 568 -11733
rect 965 -11769 1015 -11733
rect 518 -11812 590 -11769
rect 518 -11846 543 -11812
rect 577 -11846 590 -11812
rect 518 -11880 590 -11846
rect 518 -11914 543 -11880
rect 577 -11914 590 -11880
rect 518 -11933 590 -11914
rect 690 -11812 743 -11769
rect 690 -11846 701 -11812
rect 735 -11846 743 -11812
rect 690 -11880 743 -11846
rect 690 -11914 701 -11880
rect 735 -11914 743 -11880
rect 690 -11933 743 -11914
rect 797 -11811 850 -11769
rect 797 -11845 805 -11811
rect 839 -11845 850 -11811
rect 797 -11879 850 -11845
rect 797 -11913 805 -11879
rect 839 -11913 850 -11879
rect 797 -11933 850 -11913
rect 950 -11812 1015 -11769
rect 950 -11846 961 -11812
rect 995 -11846 1015 -11812
rect 950 -11880 1015 -11846
rect 950 -11914 961 -11880
rect 995 -11914 1015 -11880
rect 950 -11933 1015 -11914
rect 1045 -11811 1116 -11733
rect 1045 -11845 1059 -11811
rect 1093 -11845 1116 -11811
rect 1045 -11879 1116 -11845
rect 1045 -11913 1059 -11879
rect 1093 -11913 1116 -11879
rect 1045 -11933 1116 -11913
rect 1262 -11785 1314 -11759
rect 1262 -11819 1270 -11785
rect 1304 -11819 1314 -11785
rect 1262 -11887 1314 -11819
rect 1262 -11921 1270 -11887
rect 1304 -11921 1314 -11887
rect 1262 -11933 1314 -11921
rect 1524 -11785 1576 -11759
rect 1524 -11819 1534 -11785
rect 1568 -11819 1576 -11785
rect 1524 -11887 1576 -11819
rect 1524 -11921 1534 -11887
rect 1568 -11921 1576 -11887
rect 1722 -11785 1774 -11759
rect 1722 -11819 1730 -11785
rect 1764 -11819 1774 -11785
rect 1722 -11887 1774 -11819
rect 1524 -11933 1576 -11921
rect 1722 -11921 1730 -11887
rect 1764 -11921 1774 -11887
rect 1722 -11933 1774 -11921
rect 2352 -11785 2404 -11759
rect 2352 -11819 2362 -11785
rect 2396 -11819 2404 -11785
rect 2352 -11887 2404 -11819
rect 2352 -11921 2362 -11887
rect 2396 -11921 2404 -11887
rect 2550 -11785 2602 -11759
rect 2550 -11819 2558 -11785
rect 2592 -11819 2602 -11785
rect 2550 -11887 2602 -11819
rect 2352 -11933 2404 -11921
rect 2550 -11921 2558 -11887
rect 2592 -11921 2602 -11887
rect 2550 -11933 2602 -11921
rect 2812 -11785 2864 -11759
rect 2812 -11819 2822 -11785
rect 2856 -11819 2864 -11785
rect 2812 -11887 2864 -11819
rect 2812 -11921 2822 -11887
rect 2856 -11921 2864 -11887
rect 3010 -11812 3064 -11733
rect 3010 -11846 3019 -11812
rect 3053 -11846 3064 -11812
rect 3010 -11880 3064 -11846
rect 3010 -11914 3019 -11880
rect 3053 -11914 3064 -11880
rect 2812 -11933 2864 -11921
rect 3010 -11933 3064 -11914
rect 3094 -11769 3144 -11733
rect 3541 -11769 3591 -11733
rect 3094 -11812 3166 -11769
rect 3094 -11846 3119 -11812
rect 3153 -11846 3166 -11812
rect 3094 -11880 3166 -11846
rect 3094 -11914 3119 -11880
rect 3153 -11914 3166 -11880
rect 3094 -11933 3166 -11914
rect 3266 -11812 3319 -11769
rect 3266 -11846 3277 -11812
rect 3311 -11846 3319 -11812
rect 3266 -11880 3319 -11846
rect 3266 -11914 3277 -11880
rect 3311 -11914 3319 -11880
rect 3266 -11933 3319 -11914
rect 3373 -11811 3426 -11769
rect 3373 -11845 3381 -11811
rect 3415 -11845 3426 -11811
rect 3373 -11879 3426 -11845
rect 3373 -11913 3381 -11879
rect 3415 -11913 3426 -11879
rect 3373 -11933 3426 -11913
rect 3526 -11812 3591 -11769
rect 3526 -11846 3537 -11812
rect 3571 -11846 3591 -11812
rect 3526 -11880 3591 -11846
rect 3526 -11914 3537 -11880
rect 3571 -11914 3591 -11880
rect 3526 -11933 3591 -11914
rect 3621 -11811 3692 -11733
rect 3621 -11845 3635 -11811
rect 3669 -11845 3692 -11811
rect 3621 -11879 3692 -11845
rect 3621 -11913 3635 -11879
rect 3669 -11913 3692 -11879
rect 3621 -11933 3692 -11913
rect 3838 -11785 3890 -11759
rect 3838 -11819 3846 -11785
rect 3880 -11819 3890 -11785
rect 3838 -11887 3890 -11819
rect 3838 -11921 3846 -11887
rect 3880 -11921 3890 -11887
rect 3838 -11933 3890 -11921
rect 4100 -11785 4152 -11759
rect 4100 -11819 4110 -11785
rect 4144 -11819 4152 -11785
rect 4100 -11887 4152 -11819
rect 4100 -11921 4110 -11887
rect 4144 -11921 4152 -11887
rect 4298 -11785 4350 -11759
rect 4298 -11819 4306 -11785
rect 4340 -11819 4350 -11785
rect 4298 -11887 4350 -11819
rect 4100 -11933 4152 -11921
rect 4298 -11921 4306 -11887
rect 4340 -11921 4350 -11887
rect 4298 -11933 4350 -11921
rect 4928 -11785 4980 -11759
rect 4928 -11819 4938 -11785
rect 4972 -11819 4980 -11785
rect 4928 -11887 4980 -11819
rect 4928 -11921 4938 -11887
rect 4972 -11921 4980 -11887
rect 5126 -11785 5178 -11759
rect 5126 -11819 5134 -11785
rect 5168 -11819 5178 -11785
rect 5126 -11887 5178 -11819
rect 4928 -11933 4980 -11921
rect 5126 -11921 5134 -11887
rect 5168 -11921 5178 -11887
rect 5126 -11933 5178 -11921
rect 5388 -11785 5440 -11759
rect 5388 -11819 5398 -11785
rect 5432 -11819 5440 -11785
rect 5388 -11887 5440 -11819
rect 5388 -11921 5398 -11887
rect 5432 -11921 5440 -11887
rect 5586 -11812 5640 -11733
rect 5586 -11846 5595 -11812
rect 5629 -11846 5640 -11812
rect 5586 -11880 5640 -11846
rect 5586 -11914 5595 -11880
rect 5629 -11914 5640 -11880
rect 5388 -11933 5440 -11921
rect 5586 -11933 5640 -11914
rect 5670 -11769 5720 -11733
rect 6117 -11769 6167 -11733
rect 5670 -11812 5742 -11769
rect 5670 -11846 5695 -11812
rect 5729 -11846 5742 -11812
rect 5670 -11880 5742 -11846
rect 5670 -11914 5695 -11880
rect 5729 -11914 5742 -11880
rect 5670 -11933 5742 -11914
rect 5842 -11812 5895 -11769
rect 5842 -11846 5853 -11812
rect 5887 -11846 5895 -11812
rect 5842 -11880 5895 -11846
rect 5842 -11914 5853 -11880
rect 5887 -11914 5895 -11880
rect 5842 -11933 5895 -11914
rect 5949 -11811 6002 -11769
rect 5949 -11845 5957 -11811
rect 5991 -11845 6002 -11811
rect 5949 -11879 6002 -11845
rect 5949 -11913 5957 -11879
rect 5991 -11913 6002 -11879
rect 5949 -11933 6002 -11913
rect 6102 -11812 6167 -11769
rect 6102 -11846 6113 -11812
rect 6147 -11846 6167 -11812
rect 6102 -11880 6167 -11846
rect 6102 -11914 6113 -11880
rect 6147 -11914 6167 -11880
rect 6102 -11933 6167 -11914
rect 6197 -11811 6268 -11733
rect 6197 -11845 6211 -11811
rect 6245 -11845 6268 -11811
rect 6197 -11879 6268 -11845
rect 6197 -11913 6211 -11879
rect 6245 -11913 6268 -11879
rect 6197 -11933 6268 -11913
rect 6414 -11785 6466 -11759
rect 6414 -11819 6422 -11785
rect 6456 -11819 6466 -11785
rect 6414 -11887 6466 -11819
rect 6414 -11921 6422 -11887
rect 6456 -11921 6466 -11887
rect 6414 -11933 6466 -11921
rect 6676 -11785 6728 -11759
rect 6676 -11819 6686 -11785
rect 6720 -11819 6728 -11785
rect 6676 -11887 6728 -11819
rect 6676 -11921 6686 -11887
rect 6720 -11921 6728 -11887
rect 6874 -11785 6926 -11759
rect 6874 -11819 6882 -11785
rect 6916 -11819 6926 -11785
rect 6874 -11887 6926 -11819
rect 6676 -11933 6728 -11921
rect 6874 -11921 6882 -11887
rect 6916 -11921 6926 -11887
rect 6874 -11933 6926 -11921
rect 7504 -11785 7556 -11759
rect 7504 -11819 7514 -11785
rect 7548 -11819 7556 -11785
rect 7504 -11887 7556 -11819
rect 7504 -11921 7514 -11887
rect 7548 -11921 7556 -11887
rect 7702 -11785 7754 -11759
rect 7702 -11819 7710 -11785
rect 7744 -11819 7754 -11785
rect 7702 -11887 7754 -11819
rect 7504 -11933 7556 -11921
rect 7702 -11921 7710 -11887
rect 7744 -11921 7754 -11887
rect 7702 -11933 7754 -11921
rect 7964 -11785 8016 -11759
rect 7964 -11819 7974 -11785
rect 8008 -11819 8016 -11785
rect 7964 -11887 8016 -11819
rect 7964 -11921 7974 -11887
rect 8008 -11921 8016 -11887
rect 8162 -11812 8216 -11733
rect 8162 -11846 8171 -11812
rect 8205 -11846 8216 -11812
rect 8162 -11880 8216 -11846
rect 8162 -11914 8171 -11880
rect 8205 -11914 8216 -11880
rect 7964 -11933 8016 -11921
rect 8162 -11933 8216 -11914
rect 8246 -11769 8296 -11733
rect 8693 -11769 8743 -11733
rect 8246 -11812 8318 -11769
rect 8246 -11846 8271 -11812
rect 8305 -11846 8318 -11812
rect 8246 -11880 8318 -11846
rect 8246 -11914 8271 -11880
rect 8305 -11914 8318 -11880
rect 8246 -11933 8318 -11914
rect 8418 -11812 8471 -11769
rect 8418 -11846 8429 -11812
rect 8463 -11846 8471 -11812
rect 8418 -11880 8471 -11846
rect 8418 -11914 8429 -11880
rect 8463 -11914 8471 -11880
rect 8418 -11933 8471 -11914
rect 8525 -11811 8578 -11769
rect 8525 -11845 8533 -11811
rect 8567 -11845 8578 -11811
rect 8525 -11879 8578 -11845
rect 8525 -11913 8533 -11879
rect 8567 -11913 8578 -11879
rect 8525 -11933 8578 -11913
rect 8678 -11812 8743 -11769
rect 8678 -11846 8689 -11812
rect 8723 -11846 8743 -11812
rect 8678 -11880 8743 -11846
rect 8678 -11914 8689 -11880
rect 8723 -11914 8743 -11880
rect 8678 -11933 8743 -11914
rect 8773 -11811 8844 -11733
rect 8773 -11845 8787 -11811
rect 8821 -11845 8844 -11811
rect 8773 -11879 8844 -11845
rect 8773 -11913 8787 -11879
rect 8821 -11913 8844 -11879
rect 8773 -11933 8844 -11913
rect 8990 -11785 9042 -11759
rect 8990 -11819 8998 -11785
rect 9032 -11819 9042 -11785
rect 8990 -11887 9042 -11819
rect 8990 -11921 8998 -11887
rect 9032 -11921 9042 -11887
rect 8990 -11933 9042 -11921
rect 9252 -11785 9304 -11759
rect 9252 -11819 9262 -11785
rect 9296 -11819 9304 -11785
rect 9252 -11887 9304 -11819
rect 9252 -11921 9262 -11887
rect 9296 -11921 9304 -11887
rect 9450 -11785 9502 -11759
rect 9450 -11819 9458 -11785
rect 9492 -11819 9502 -11785
rect 9450 -11887 9502 -11819
rect 9252 -11933 9304 -11921
rect 9450 -11921 9458 -11887
rect 9492 -11921 9502 -11887
rect 9450 -11933 9502 -11921
rect 10080 -11785 10132 -11759
rect 10080 -11819 10090 -11785
rect 10124 -11819 10132 -11785
rect 10080 -11887 10132 -11819
rect 10080 -11921 10090 -11887
rect 10124 -11921 10132 -11887
rect 10370 -11785 10422 -11759
rect 10370 -11819 10378 -11785
rect 10412 -11819 10422 -11785
rect 10370 -11887 10422 -11819
rect 10080 -11933 10132 -11921
rect 10370 -11921 10378 -11887
rect 10412 -11921 10422 -11887
rect 10370 -11933 10422 -11921
rect 10632 -11785 10684 -11759
rect 10632 -11819 10642 -11785
rect 10676 -11819 10684 -11785
rect 10632 -11887 10684 -11819
rect 10632 -11921 10642 -11887
rect 10676 -11921 10684 -11887
rect 10632 -11933 10684 -11921
rect 10738 -11812 10792 -11733
rect 10738 -11846 10747 -11812
rect 10781 -11846 10792 -11812
rect 10738 -11880 10792 -11846
rect 10738 -11914 10747 -11880
rect 10781 -11914 10792 -11880
rect 10738 -11933 10792 -11914
rect 10822 -11769 10872 -11733
rect 11269 -11769 11319 -11733
rect 10822 -11812 10894 -11769
rect 10822 -11846 10847 -11812
rect 10881 -11846 10894 -11812
rect 10822 -11880 10894 -11846
rect 10822 -11914 10847 -11880
rect 10881 -11914 10894 -11880
rect 10822 -11933 10894 -11914
rect 10994 -11812 11047 -11769
rect 10994 -11846 11005 -11812
rect 11039 -11846 11047 -11812
rect 10994 -11880 11047 -11846
rect 10994 -11914 11005 -11880
rect 11039 -11914 11047 -11880
rect 10994 -11933 11047 -11914
rect 11101 -11811 11154 -11769
rect 11101 -11845 11109 -11811
rect 11143 -11845 11154 -11811
rect 11101 -11879 11154 -11845
rect 11101 -11913 11109 -11879
rect 11143 -11913 11154 -11879
rect 11101 -11933 11154 -11913
rect 11254 -11812 11319 -11769
rect 11254 -11846 11265 -11812
rect 11299 -11846 11319 -11812
rect 11254 -11880 11319 -11846
rect 11254 -11914 11265 -11880
rect 11299 -11914 11319 -11880
rect 11254 -11933 11319 -11914
rect 11349 -11811 11420 -11733
rect 11349 -11845 11363 -11811
rect 11397 -11845 11420 -11811
rect 11349 -11879 11420 -11845
rect 11349 -11913 11363 -11879
rect 11397 -11913 11420 -11879
rect 11349 -11933 11420 -11913
rect 11658 -11785 11710 -11759
rect 11658 -11819 11666 -11785
rect 11700 -11819 11710 -11785
rect 11658 -11887 11710 -11819
rect 11658 -11921 11666 -11887
rect 11700 -11921 11710 -11887
rect 11658 -11933 11710 -11921
rect 11920 -11785 11972 -11759
rect 11920 -11819 11930 -11785
rect 11964 -11819 11972 -11785
rect 11920 -11887 11972 -11819
rect 11920 -11921 11930 -11887
rect 11964 -11921 11972 -11887
rect 12486 -11812 12547 -11733
rect 12486 -11846 12502 -11812
rect 12536 -11846 12547 -11812
rect 12486 -11880 12547 -11846
rect 12486 -11914 12502 -11880
rect 12536 -11914 12547 -11880
rect 11920 -11933 11972 -11921
rect 12486 -11933 12547 -11914
rect 12577 -11785 12633 -11733
rect 12577 -11819 12588 -11785
rect 12622 -11819 12633 -11785
rect 12577 -11873 12633 -11819
rect 12577 -11907 12588 -11873
rect 12622 -11907 12633 -11873
rect 12577 -11933 12633 -11907
rect 12663 -11812 12719 -11733
rect 12663 -11846 12674 -11812
rect 12708 -11846 12719 -11812
rect 12663 -11880 12719 -11846
rect 12663 -11914 12674 -11880
rect 12708 -11914 12719 -11880
rect 12663 -11933 12719 -11914
rect 12749 -11785 12805 -11733
rect 12749 -11819 12760 -11785
rect 12794 -11819 12805 -11785
rect 12749 -11873 12805 -11819
rect 12749 -11907 12760 -11873
rect 12794 -11907 12805 -11873
rect 12749 -11933 12805 -11907
rect 12835 -11812 12891 -11733
rect 12835 -11846 12846 -11812
rect 12880 -11846 12891 -11812
rect 12835 -11880 12891 -11846
rect 12835 -11914 12846 -11880
rect 12880 -11914 12891 -11880
rect 12835 -11933 12891 -11914
rect 12921 -11785 12977 -11733
rect 12921 -11819 12932 -11785
rect 12966 -11819 12977 -11785
rect 12921 -11873 12977 -11819
rect 12921 -11907 12932 -11873
rect 12966 -11907 12977 -11873
rect 12921 -11933 12977 -11907
rect 13007 -11812 13076 -11733
rect 13007 -11846 13018 -11812
rect 13052 -11846 13076 -11812
rect 13007 -11880 13076 -11846
rect 13007 -11914 13018 -11880
rect 13052 -11914 13076 -11880
rect 13007 -11933 13076 -11914
rect 13222 -11785 13274 -11759
rect 13222 -11819 13230 -11785
rect 13264 -11819 13274 -11785
rect 13222 -11887 13274 -11819
rect 13222 -11921 13230 -11887
rect 13264 -11921 13274 -11887
rect 13222 -11933 13274 -11921
rect 13484 -11785 13536 -11759
rect 13484 -11819 13494 -11785
rect 13528 -11819 13536 -11785
rect 13484 -11887 13536 -11819
rect 13484 -11921 13494 -11887
rect 13528 -11921 13536 -11887
rect 13682 -11819 13735 -11733
rect 13682 -11853 13690 -11819
rect 13724 -11853 13735 -11819
rect 13682 -11887 13735 -11853
rect 13484 -11933 13536 -11921
rect 13682 -11921 13690 -11887
rect 13724 -11921 13735 -11887
rect 13682 -11933 13735 -11921
rect 13765 -11811 13821 -11733
rect 13765 -11845 13776 -11811
rect 13810 -11845 13821 -11811
rect 13765 -11879 13821 -11845
rect 13765 -11913 13776 -11879
rect 13810 -11913 13821 -11879
rect 13765 -11933 13821 -11913
rect 13851 -11819 13907 -11733
rect 13851 -11853 13862 -11819
rect 13896 -11853 13907 -11819
rect 13851 -11887 13907 -11853
rect 13851 -11921 13862 -11887
rect 13896 -11921 13907 -11887
rect 13851 -11933 13907 -11921
rect 13937 -11803 13993 -11733
rect 13937 -11837 13948 -11803
rect 13982 -11837 13993 -11803
rect 13937 -11871 13993 -11837
rect 13937 -11905 13948 -11871
rect 13982 -11905 13993 -11871
rect 13937 -11933 13993 -11905
rect 14023 -11819 14079 -11733
rect 14023 -11853 14034 -11819
rect 14068 -11853 14079 -11819
rect 14023 -11887 14079 -11853
rect 14023 -11921 14034 -11887
rect 14068 -11921 14079 -11887
rect 14023 -11933 14079 -11921
rect 14109 -11757 14165 -11733
rect 14109 -11791 14120 -11757
rect 14154 -11791 14165 -11757
rect 14109 -11843 14165 -11791
rect 14109 -11877 14120 -11843
rect 14154 -11877 14165 -11843
rect 14109 -11933 14165 -11877
rect 14195 -11863 14251 -11733
rect 14195 -11897 14206 -11863
rect 14240 -11897 14251 -11863
rect 14195 -11933 14251 -11897
rect 14281 -11757 14337 -11733
rect 14281 -11791 14292 -11757
rect 14326 -11791 14337 -11757
rect 14281 -11843 14337 -11791
rect 14281 -11877 14292 -11843
rect 14326 -11877 14337 -11843
rect 14281 -11933 14337 -11877
rect 14367 -11863 14423 -11733
rect 14367 -11897 14378 -11863
rect 14412 -11897 14423 -11863
rect 14367 -11933 14423 -11897
rect 14453 -11757 14509 -11733
rect 14453 -11791 14464 -11757
rect 14498 -11791 14509 -11757
rect 14453 -11843 14509 -11791
rect 14453 -11877 14464 -11843
rect 14498 -11877 14509 -11843
rect 14453 -11933 14509 -11877
rect 14539 -11863 14595 -11733
rect 14539 -11897 14550 -11863
rect 14584 -11897 14595 -11863
rect 14539 -11933 14595 -11897
rect 14625 -11757 14681 -11733
rect 14625 -11791 14636 -11757
rect 14670 -11791 14681 -11757
rect 14625 -11843 14681 -11791
rect 14625 -11877 14636 -11843
rect 14670 -11877 14681 -11843
rect 14625 -11933 14681 -11877
rect 14711 -11863 14766 -11733
rect 14711 -11897 14722 -11863
rect 14756 -11897 14766 -11863
rect 14711 -11933 14766 -11897
rect 14796 -11757 14852 -11733
rect 14796 -11791 14807 -11757
rect 14841 -11791 14852 -11757
rect 14796 -11843 14852 -11791
rect 14796 -11877 14807 -11843
rect 14841 -11877 14852 -11843
rect 14796 -11933 14852 -11877
rect 14882 -11863 14938 -11733
rect 14882 -11897 14893 -11863
rect 14927 -11897 14938 -11863
rect 14882 -11933 14938 -11897
rect 14968 -11757 15024 -11733
rect 14968 -11791 14979 -11757
rect 15013 -11791 15024 -11757
rect 14968 -11843 15024 -11791
rect 14968 -11877 14979 -11843
rect 15013 -11877 15024 -11843
rect 14968 -11933 15024 -11877
rect 15054 -11863 15110 -11733
rect 15054 -11897 15065 -11863
rect 15099 -11897 15110 -11863
rect 15054 -11933 15110 -11897
rect 15140 -11757 15196 -11733
rect 15140 -11791 15151 -11757
rect 15185 -11791 15196 -11757
rect 15140 -11843 15196 -11791
rect 15140 -11877 15151 -11843
rect 15185 -11877 15196 -11843
rect 15140 -11933 15196 -11877
rect 15226 -11863 15282 -11733
rect 15226 -11897 15237 -11863
rect 15271 -11897 15282 -11863
rect 15226 -11933 15282 -11897
rect 15312 -11757 15368 -11733
rect 15312 -11791 15323 -11757
rect 15357 -11791 15368 -11757
rect 15312 -11843 15368 -11791
rect 15312 -11877 15323 -11843
rect 15357 -11877 15368 -11843
rect 15312 -11933 15368 -11877
rect 15398 -11863 15451 -11733
rect 15398 -11897 15409 -11863
rect 15443 -11897 15451 -11863
rect 15398 -11933 15451 -11897
rect 15614 -11785 15666 -11759
rect 15614 -11819 15622 -11785
rect 15656 -11819 15666 -11785
rect 15614 -11887 15666 -11819
rect 15614 -11921 15622 -11887
rect 15656 -11921 15666 -11887
rect 15614 -11933 15666 -11921
rect 16612 -11785 16664 -11759
rect 16612 -11819 16622 -11785
rect 16656 -11819 16664 -11785
rect 16612 -11887 16664 -11819
rect 16612 -11921 16622 -11887
rect 16656 -11921 16664 -11887
rect 16612 -11933 16664 -11921
rect -2970 -12039 -2918 -12027
rect -2970 -12073 -2962 -12039
rect -2928 -12073 -2918 -12039
rect -2970 -12141 -2918 -12073
rect -2970 -12175 -2962 -12141
rect -2928 -12175 -2918 -12141
rect -2970 -12201 -2918 -12175
rect -2340 -12039 -2288 -12027
rect -2340 -12073 -2330 -12039
rect -2296 -12073 -2288 -12039
rect -1590 -12039 -1538 -12027
rect -2340 -12141 -2288 -12073
rect -2340 -12175 -2330 -12141
rect -2296 -12175 -2288 -12141
rect -2340 -12201 -2288 -12175
rect -1590 -12073 -1582 -12039
rect -1548 -12073 -1538 -12039
rect -1590 -12141 -1538 -12073
rect -1590 -12175 -1582 -12141
rect -1548 -12175 -1538 -12141
rect -1590 -12201 -1538 -12175
rect -960 -12039 -908 -12027
rect -960 -12073 -950 -12039
rect -916 -12073 -908 -12039
rect -960 -12141 -908 -12073
rect -960 -12175 -950 -12141
rect -916 -12175 -908 -12141
rect -960 -12201 -908 -12175
rect -854 -12047 -783 -12027
rect -854 -12081 -831 -12047
rect -797 -12081 -783 -12047
rect -854 -12115 -783 -12081
rect -854 -12149 -831 -12115
rect -797 -12149 -783 -12115
rect -854 -12227 -783 -12149
rect -753 -12046 -688 -12027
rect -753 -12080 -733 -12046
rect -699 -12080 -688 -12046
rect -753 -12114 -688 -12080
rect -753 -12148 -733 -12114
rect -699 -12148 -688 -12114
rect -753 -12191 -688 -12148
rect -588 -12047 -535 -12027
rect -588 -12081 -577 -12047
rect -543 -12081 -535 -12047
rect -588 -12115 -535 -12081
rect -588 -12149 -577 -12115
rect -543 -12149 -535 -12115
rect -588 -12191 -535 -12149
rect -481 -12046 -428 -12027
rect -481 -12080 -473 -12046
rect -439 -12080 -428 -12046
rect -481 -12114 -428 -12080
rect -481 -12148 -473 -12114
rect -439 -12148 -428 -12114
rect -481 -12191 -428 -12148
rect -328 -12046 -256 -12027
rect -328 -12080 -315 -12046
rect -281 -12080 -256 -12046
rect -328 -12114 -256 -12080
rect -328 -12148 -315 -12114
rect -281 -12148 -256 -12114
rect -328 -12191 -256 -12148
rect -753 -12227 -703 -12191
rect -306 -12227 -256 -12191
rect -226 -12046 -172 -12027
rect -26 -12039 26 -12027
rect -226 -12080 -215 -12046
rect -181 -12080 -172 -12046
rect -226 -12114 -172 -12080
rect -226 -12148 -215 -12114
rect -181 -12148 -172 -12114
rect -226 -12227 -172 -12148
rect -26 -12073 -18 -12039
rect 16 -12073 26 -12039
rect -26 -12141 26 -12073
rect -26 -12175 -18 -12141
rect 16 -12175 26 -12141
rect -26 -12201 26 -12175
rect 236 -12039 288 -12027
rect 236 -12073 246 -12039
rect 280 -12073 288 -12039
rect 236 -12141 288 -12073
rect 236 -12175 246 -12141
rect 280 -12175 288 -12141
rect 236 -12201 288 -12175
rect 434 -12047 505 -12027
rect 434 -12081 457 -12047
rect 491 -12081 505 -12047
rect 434 -12115 505 -12081
rect 434 -12149 457 -12115
rect 491 -12149 505 -12115
rect 434 -12227 505 -12149
rect 535 -12046 600 -12027
rect 535 -12080 555 -12046
rect 589 -12080 600 -12046
rect 535 -12114 600 -12080
rect 535 -12148 555 -12114
rect 589 -12148 600 -12114
rect 535 -12191 600 -12148
rect 700 -12047 753 -12027
rect 700 -12081 711 -12047
rect 745 -12081 753 -12047
rect 700 -12115 753 -12081
rect 700 -12149 711 -12115
rect 745 -12149 753 -12115
rect 700 -12191 753 -12149
rect 807 -12046 860 -12027
rect 807 -12080 815 -12046
rect 849 -12080 860 -12046
rect 807 -12114 860 -12080
rect 807 -12148 815 -12114
rect 849 -12148 860 -12114
rect 807 -12191 860 -12148
rect 960 -12046 1032 -12027
rect 960 -12080 973 -12046
rect 1007 -12080 1032 -12046
rect 960 -12114 1032 -12080
rect 960 -12148 973 -12114
rect 1007 -12148 1032 -12114
rect 960 -12191 1032 -12148
rect 535 -12227 585 -12191
rect 982 -12227 1032 -12191
rect 1062 -12046 1116 -12027
rect 1262 -12039 1314 -12027
rect 1062 -12080 1073 -12046
rect 1107 -12080 1116 -12046
rect 1062 -12114 1116 -12080
rect 1062 -12148 1073 -12114
rect 1107 -12148 1116 -12114
rect 1062 -12227 1116 -12148
rect 1262 -12073 1270 -12039
rect 1304 -12073 1314 -12039
rect 1262 -12141 1314 -12073
rect 1262 -12175 1270 -12141
rect 1304 -12175 1314 -12141
rect 1262 -12201 1314 -12175
rect 1524 -12039 1576 -12027
rect 1524 -12073 1534 -12039
rect 1568 -12073 1576 -12039
rect 1722 -12039 1774 -12027
rect 1524 -12141 1576 -12073
rect 1524 -12175 1534 -12141
rect 1568 -12175 1576 -12141
rect 1524 -12201 1576 -12175
rect 1722 -12073 1730 -12039
rect 1764 -12073 1774 -12039
rect 1722 -12141 1774 -12073
rect 1722 -12175 1730 -12141
rect 1764 -12175 1774 -12141
rect 1722 -12201 1774 -12175
rect 2352 -12039 2404 -12027
rect 2352 -12073 2362 -12039
rect 2396 -12073 2404 -12039
rect 2550 -12039 2602 -12027
rect 2352 -12141 2404 -12073
rect 2352 -12175 2362 -12141
rect 2396 -12175 2404 -12141
rect 2352 -12201 2404 -12175
rect 2550 -12073 2558 -12039
rect 2592 -12073 2602 -12039
rect 2550 -12141 2602 -12073
rect 2550 -12175 2558 -12141
rect 2592 -12175 2602 -12141
rect 2550 -12201 2602 -12175
rect 2812 -12039 2864 -12027
rect 2812 -12073 2822 -12039
rect 2856 -12073 2864 -12039
rect 2812 -12141 2864 -12073
rect 2812 -12175 2822 -12141
rect 2856 -12175 2864 -12141
rect 2812 -12201 2864 -12175
rect 3010 -12047 3081 -12027
rect 3010 -12081 3033 -12047
rect 3067 -12081 3081 -12047
rect 3010 -12115 3081 -12081
rect 3010 -12149 3033 -12115
rect 3067 -12149 3081 -12115
rect 3010 -12227 3081 -12149
rect 3111 -12046 3176 -12027
rect 3111 -12080 3131 -12046
rect 3165 -12080 3176 -12046
rect 3111 -12114 3176 -12080
rect 3111 -12148 3131 -12114
rect 3165 -12148 3176 -12114
rect 3111 -12191 3176 -12148
rect 3276 -12047 3329 -12027
rect 3276 -12081 3287 -12047
rect 3321 -12081 3329 -12047
rect 3276 -12115 3329 -12081
rect 3276 -12149 3287 -12115
rect 3321 -12149 3329 -12115
rect 3276 -12191 3329 -12149
rect 3383 -12046 3436 -12027
rect 3383 -12080 3391 -12046
rect 3425 -12080 3436 -12046
rect 3383 -12114 3436 -12080
rect 3383 -12148 3391 -12114
rect 3425 -12148 3436 -12114
rect 3383 -12191 3436 -12148
rect 3536 -12046 3608 -12027
rect 3536 -12080 3549 -12046
rect 3583 -12080 3608 -12046
rect 3536 -12114 3608 -12080
rect 3536 -12148 3549 -12114
rect 3583 -12148 3608 -12114
rect 3536 -12191 3608 -12148
rect 3111 -12227 3161 -12191
rect 3558 -12227 3608 -12191
rect 3638 -12046 3692 -12027
rect 3838 -12039 3890 -12027
rect 3638 -12080 3649 -12046
rect 3683 -12080 3692 -12046
rect 3638 -12114 3692 -12080
rect 3638 -12148 3649 -12114
rect 3683 -12148 3692 -12114
rect 3638 -12227 3692 -12148
rect 3838 -12073 3846 -12039
rect 3880 -12073 3890 -12039
rect 3838 -12141 3890 -12073
rect 3838 -12175 3846 -12141
rect 3880 -12175 3890 -12141
rect 3838 -12201 3890 -12175
rect 4100 -12039 4152 -12027
rect 4100 -12073 4110 -12039
rect 4144 -12073 4152 -12039
rect 4298 -12039 4350 -12027
rect 4100 -12141 4152 -12073
rect 4100 -12175 4110 -12141
rect 4144 -12175 4152 -12141
rect 4100 -12201 4152 -12175
rect 4298 -12073 4306 -12039
rect 4340 -12073 4350 -12039
rect 4298 -12141 4350 -12073
rect 4298 -12175 4306 -12141
rect 4340 -12175 4350 -12141
rect 4298 -12201 4350 -12175
rect 4928 -12039 4980 -12027
rect 4928 -12073 4938 -12039
rect 4972 -12073 4980 -12039
rect 5126 -12039 5178 -12027
rect 4928 -12141 4980 -12073
rect 4928 -12175 4938 -12141
rect 4972 -12175 4980 -12141
rect 4928 -12201 4980 -12175
rect 5126 -12073 5134 -12039
rect 5168 -12073 5178 -12039
rect 5126 -12141 5178 -12073
rect 5126 -12175 5134 -12141
rect 5168 -12175 5178 -12141
rect 5126 -12201 5178 -12175
rect 5388 -12039 5440 -12027
rect 5388 -12073 5398 -12039
rect 5432 -12073 5440 -12039
rect 5388 -12141 5440 -12073
rect 5388 -12175 5398 -12141
rect 5432 -12175 5440 -12141
rect 5388 -12201 5440 -12175
rect 5586 -12047 5657 -12027
rect 5586 -12081 5609 -12047
rect 5643 -12081 5657 -12047
rect 5586 -12115 5657 -12081
rect 5586 -12149 5609 -12115
rect 5643 -12149 5657 -12115
rect 5586 -12227 5657 -12149
rect 5687 -12046 5752 -12027
rect 5687 -12080 5707 -12046
rect 5741 -12080 5752 -12046
rect 5687 -12114 5752 -12080
rect 5687 -12148 5707 -12114
rect 5741 -12148 5752 -12114
rect 5687 -12191 5752 -12148
rect 5852 -12047 5905 -12027
rect 5852 -12081 5863 -12047
rect 5897 -12081 5905 -12047
rect 5852 -12115 5905 -12081
rect 5852 -12149 5863 -12115
rect 5897 -12149 5905 -12115
rect 5852 -12191 5905 -12149
rect 5959 -12046 6012 -12027
rect 5959 -12080 5967 -12046
rect 6001 -12080 6012 -12046
rect 5959 -12114 6012 -12080
rect 5959 -12148 5967 -12114
rect 6001 -12148 6012 -12114
rect 5959 -12191 6012 -12148
rect 6112 -12046 6184 -12027
rect 6112 -12080 6125 -12046
rect 6159 -12080 6184 -12046
rect 6112 -12114 6184 -12080
rect 6112 -12148 6125 -12114
rect 6159 -12148 6184 -12114
rect 6112 -12191 6184 -12148
rect 5687 -12227 5737 -12191
rect 6134 -12227 6184 -12191
rect 6214 -12046 6268 -12027
rect 6414 -12039 6466 -12027
rect 6214 -12080 6225 -12046
rect 6259 -12080 6268 -12046
rect 6214 -12114 6268 -12080
rect 6214 -12148 6225 -12114
rect 6259 -12148 6268 -12114
rect 6214 -12227 6268 -12148
rect 6414 -12073 6422 -12039
rect 6456 -12073 6466 -12039
rect 6414 -12141 6466 -12073
rect 6414 -12175 6422 -12141
rect 6456 -12175 6466 -12141
rect 6414 -12201 6466 -12175
rect 6676 -12039 6728 -12027
rect 6676 -12073 6686 -12039
rect 6720 -12073 6728 -12039
rect 6874 -12039 6926 -12027
rect 6676 -12141 6728 -12073
rect 6676 -12175 6686 -12141
rect 6720 -12175 6728 -12141
rect 6676 -12201 6728 -12175
rect 6874 -12073 6882 -12039
rect 6916 -12073 6926 -12039
rect 6874 -12141 6926 -12073
rect 6874 -12175 6882 -12141
rect 6916 -12175 6926 -12141
rect 6874 -12201 6926 -12175
rect 7504 -12039 7556 -12027
rect 7504 -12073 7514 -12039
rect 7548 -12073 7556 -12039
rect 7702 -12039 7754 -12027
rect 7504 -12141 7556 -12073
rect 7504 -12175 7514 -12141
rect 7548 -12175 7556 -12141
rect 7504 -12201 7556 -12175
rect 7702 -12073 7710 -12039
rect 7744 -12073 7754 -12039
rect 7702 -12141 7754 -12073
rect 7702 -12175 7710 -12141
rect 7744 -12175 7754 -12141
rect 7702 -12201 7754 -12175
rect 7964 -12039 8016 -12027
rect 7964 -12073 7974 -12039
rect 8008 -12073 8016 -12039
rect 7964 -12141 8016 -12073
rect 7964 -12175 7974 -12141
rect 8008 -12175 8016 -12141
rect 7964 -12201 8016 -12175
rect 8162 -12047 8233 -12027
rect 8162 -12081 8185 -12047
rect 8219 -12081 8233 -12047
rect 8162 -12115 8233 -12081
rect 8162 -12149 8185 -12115
rect 8219 -12149 8233 -12115
rect 8162 -12227 8233 -12149
rect 8263 -12046 8328 -12027
rect 8263 -12080 8283 -12046
rect 8317 -12080 8328 -12046
rect 8263 -12114 8328 -12080
rect 8263 -12148 8283 -12114
rect 8317 -12148 8328 -12114
rect 8263 -12191 8328 -12148
rect 8428 -12047 8481 -12027
rect 8428 -12081 8439 -12047
rect 8473 -12081 8481 -12047
rect 8428 -12115 8481 -12081
rect 8428 -12149 8439 -12115
rect 8473 -12149 8481 -12115
rect 8428 -12191 8481 -12149
rect 8535 -12046 8588 -12027
rect 8535 -12080 8543 -12046
rect 8577 -12080 8588 -12046
rect 8535 -12114 8588 -12080
rect 8535 -12148 8543 -12114
rect 8577 -12148 8588 -12114
rect 8535 -12191 8588 -12148
rect 8688 -12046 8760 -12027
rect 8688 -12080 8701 -12046
rect 8735 -12080 8760 -12046
rect 8688 -12114 8760 -12080
rect 8688 -12148 8701 -12114
rect 8735 -12148 8760 -12114
rect 8688 -12191 8760 -12148
rect 8263 -12227 8313 -12191
rect 8710 -12227 8760 -12191
rect 8790 -12046 8844 -12027
rect 8990 -12039 9042 -12027
rect 8790 -12080 8801 -12046
rect 8835 -12080 8844 -12046
rect 8790 -12114 8844 -12080
rect 8790 -12148 8801 -12114
rect 8835 -12148 8844 -12114
rect 8790 -12227 8844 -12148
rect 8990 -12073 8998 -12039
rect 9032 -12073 9042 -12039
rect 8990 -12141 9042 -12073
rect 8990 -12175 8998 -12141
rect 9032 -12175 9042 -12141
rect 8990 -12201 9042 -12175
rect 9252 -12039 9304 -12027
rect 9252 -12073 9262 -12039
rect 9296 -12073 9304 -12039
rect 9450 -12039 9502 -12027
rect 9252 -12141 9304 -12073
rect 9252 -12175 9262 -12141
rect 9296 -12175 9304 -12141
rect 9252 -12201 9304 -12175
rect 9450 -12073 9458 -12039
rect 9492 -12073 9502 -12039
rect 9450 -12141 9502 -12073
rect 9450 -12175 9458 -12141
rect 9492 -12175 9502 -12141
rect 9450 -12201 9502 -12175
rect 10080 -12039 10132 -12027
rect 10080 -12073 10090 -12039
rect 10124 -12073 10132 -12039
rect 10370 -12039 10422 -12027
rect 10080 -12141 10132 -12073
rect 10080 -12175 10090 -12141
rect 10124 -12175 10132 -12141
rect 10080 -12201 10132 -12175
rect 10370 -12073 10378 -12039
rect 10412 -12073 10422 -12039
rect 10370 -12141 10422 -12073
rect 10370 -12175 10378 -12141
rect 10412 -12175 10422 -12141
rect 10370 -12201 10422 -12175
rect 10632 -12039 10684 -12027
rect 10632 -12073 10642 -12039
rect 10676 -12073 10684 -12039
rect 10632 -12141 10684 -12073
rect 10632 -12175 10642 -12141
rect 10676 -12175 10684 -12141
rect 10632 -12201 10684 -12175
rect 10738 -12047 10809 -12027
rect 10738 -12081 10761 -12047
rect 10795 -12081 10809 -12047
rect 10738 -12115 10809 -12081
rect 10738 -12149 10761 -12115
rect 10795 -12149 10809 -12115
rect 10738 -12227 10809 -12149
rect 10839 -12046 10904 -12027
rect 10839 -12080 10859 -12046
rect 10893 -12080 10904 -12046
rect 10839 -12114 10904 -12080
rect 10839 -12148 10859 -12114
rect 10893 -12148 10904 -12114
rect 10839 -12191 10904 -12148
rect 11004 -12047 11057 -12027
rect 11004 -12081 11015 -12047
rect 11049 -12081 11057 -12047
rect 11004 -12115 11057 -12081
rect 11004 -12149 11015 -12115
rect 11049 -12149 11057 -12115
rect 11004 -12191 11057 -12149
rect 11111 -12046 11164 -12027
rect 11111 -12080 11119 -12046
rect 11153 -12080 11164 -12046
rect 11111 -12114 11164 -12080
rect 11111 -12148 11119 -12114
rect 11153 -12148 11164 -12114
rect 11111 -12191 11164 -12148
rect 11264 -12046 11336 -12027
rect 11264 -12080 11277 -12046
rect 11311 -12080 11336 -12046
rect 11264 -12114 11336 -12080
rect 11264 -12148 11277 -12114
rect 11311 -12148 11336 -12114
rect 11264 -12191 11336 -12148
rect 10839 -12227 10889 -12191
rect 11286 -12227 11336 -12191
rect 11366 -12046 11420 -12027
rect 11658 -12039 11710 -12027
rect 11366 -12080 11377 -12046
rect 11411 -12080 11420 -12046
rect 11366 -12114 11420 -12080
rect 11366 -12148 11377 -12114
rect 11411 -12148 11420 -12114
rect 11366 -12227 11420 -12148
rect 11658 -12073 11666 -12039
rect 11700 -12073 11710 -12039
rect 11658 -12141 11710 -12073
rect 11658 -12175 11666 -12141
rect 11700 -12175 11710 -12141
rect 11658 -12201 11710 -12175
rect 11920 -12039 11972 -12027
rect 11920 -12073 11930 -12039
rect 11964 -12073 11972 -12039
rect 13682 -12039 13735 -12027
rect 11920 -12141 11972 -12073
rect 11920 -12175 11930 -12141
rect 11964 -12175 11972 -12141
rect 11920 -12201 11972 -12175
rect 13682 -12073 13690 -12039
rect 13724 -12073 13735 -12039
rect 13682 -12107 13735 -12073
rect 13682 -12141 13690 -12107
rect 13724 -12141 13735 -12107
rect 13682 -12227 13735 -12141
rect 13765 -12047 13821 -12027
rect 13765 -12081 13776 -12047
rect 13810 -12081 13821 -12047
rect 13765 -12115 13821 -12081
rect 13765 -12149 13776 -12115
rect 13810 -12149 13821 -12115
rect 13765 -12227 13821 -12149
rect 13851 -12039 13907 -12027
rect 13851 -12073 13862 -12039
rect 13896 -12073 13907 -12039
rect 13851 -12107 13907 -12073
rect 13851 -12141 13862 -12107
rect 13896 -12141 13907 -12107
rect 13851 -12227 13907 -12141
rect 13937 -12055 13993 -12027
rect 13937 -12089 13948 -12055
rect 13982 -12089 13993 -12055
rect 13937 -12123 13993 -12089
rect 13937 -12157 13948 -12123
rect 13982 -12157 13993 -12123
rect 13937 -12227 13993 -12157
rect 14023 -12039 14079 -12027
rect 14023 -12073 14034 -12039
rect 14068 -12073 14079 -12039
rect 14023 -12107 14079 -12073
rect 14023 -12141 14034 -12107
rect 14068 -12141 14079 -12107
rect 14023 -12227 14079 -12141
rect 14109 -12083 14165 -12027
rect 14109 -12117 14120 -12083
rect 14154 -12117 14165 -12083
rect 14109 -12169 14165 -12117
rect 14109 -12203 14120 -12169
rect 14154 -12203 14165 -12169
rect 14109 -12227 14165 -12203
rect 14195 -12063 14251 -12027
rect 14195 -12097 14206 -12063
rect 14240 -12097 14251 -12063
rect 14195 -12227 14251 -12097
rect 14281 -12083 14337 -12027
rect 14281 -12117 14292 -12083
rect 14326 -12117 14337 -12083
rect 14281 -12169 14337 -12117
rect 14281 -12203 14292 -12169
rect 14326 -12203 14337 -12169
rect 14281 -12227 14337 -12203
rect 14367 -12063 14423 -12027
rect 14367 -12097 14378 -12063
rect 14412 -12097 14423 -12063
rect 14367 -12227 14423 -12097
rect 14453 -12083 14509 -12027
rect 14453 -12117 14464 -12083
rect 14498 -12117 14509 -12083
rect 14453 -12169 14509 -12117
rect 14453 -12203 14464 -12169
rect 14498 -12203 14509 -12169
rect 14453 -12227 14509 -12203
rect 14539 -12063 14595 -12027
rect 14539 -12097 14550 -12063
rect 14584 -12097 14595 -12063
rect 14539 -12227 14595 -12097
rect 14625 -12083 14681 -12027
rect 14625 -12117 14636 -12083
rect 14670 -12117 14681 -12083
rect 14625 -12169 14681 -12117
rect 14625 -12203 14636 -12169
rect 14670 -12203 14681 -12169
rect 14625 -12227 14681 -12203
rect 14711 -12063 14766 -12027
rect 14711 -12097 14722 -12063
rect 14756 -12097 14766 -12063
rect 14711 -12227 14766 -12097
rect 14796 -12083 14852 -12027
rect 14796 -12117 14807 -12083
rect 14841 -12117 14852 -12083
rect 14796 -12169 14852 -12117
rect 14796 -12203 14807 -12169
rect 14841 -12203 14852 -12169
rect 14796 -12227 14852 -12203
rect 14882 -12063 14938 -12027
rect 14882 -12097 14893 -12063
rect 14927 -12097 14938 -12063
rect 14882 -12227 14938 -12097
rect 14968 -12083 15024 -12027
rect 14968 -12117 14979 -12083
rect 15013 -12117 15024 -12083
rect 14968 -12169 15024 -12117
rect 14968 -12203 14979 -12169
rect 15013 -12203 15024 -12169
rect 14968 -12227 15024 -12203
rect 15054 -12063 15110 -12027
rect 15054 -12097 15065 -12063
rect 15099 -12097 15110 -12063
rect 15054 -12227 15110 -12097
rect 15140 -12083 15196 -12027
rect 15140 -12117 15151 -12083
rect 15185 -12117 15196 -12083
rect 15140 -12169 15196 -12117
rect 15140 -12203 15151 -12169
rect 15185 -12203 15196 -12169
rect 15140 -12227 15196 -12203
rect 15226 -12063 15282 -12027
rect 15226 -12097 15237 -12063
rect 15271 -12097 15282 -12063
rect 15226 -12227 15282 -12097
rect 15312 -12083 15368 -12027
rect 15312 -12117 15323 -12083
rect 15357 -12117 15368 -12083
rect 15312 -12169 15368 -12117
rect 15312 -12203 15323 -12169
rect 15357 -12203 15368 -12169
rect 15312 -12227 15368 -12203
rect 15398 -12063 15451 -12027
rect 15614 -12039 15666 -12027
rect 15398 -12097 15409 -12063
rect 15443 -12097 15451 -12063
rect 15398 -12227 15451 -12097
rect 15614 -12073 15622 -12039
rect 15656 -12073 15666 -12039
rect 15614 -12141 15666 -12073
rect 15614 -12175 15622 -12141
rect 15656 -12175 15666 -12141
rect 15614 -12201 15666 -12175
rect 16612 -12039 16664 -12027
rect 16612 -12073 16622 -12039
rect 16656 -12073 16664 -12039
rect 16612 -12141 16664 -12073
rect 16612 -12175 16622 -12141
rect 16656 -12175 16664 -12141
rect 16612 -12201 16664 -12175
rect -2970 -12873 -2918 -12847
rect -2970 -12907 -2962 -12873
rect -2928 -12907 -2918 -12873
rect -2970 -12975 -2918 -12907
rect -2970 -13009 -2962 -12975
rect -2928 -13009 -2918 -12975
rect -2970 -13021 -2918 -13009
rect -2340 -12873 -2288 -12847
rect -2340 -12907 -2330 -12873
rect -2296 -12907 -2288 -12873
rect -2340 -12975 -2288 -12907
rect -2340 -13009 -2330 -12975
rect -2296 -13009 -2288 -12975
rect -1590 -12873 -1538 -12847
rect -1590 -12907 -1582 -12873
rect -1548 -12907 -1538 -12873
rect -1590 -12975 -1538 -12907
rect -2340 -13021 -2288 -13009
rect -1590 -13009 -1582 -12975
rect -1548 -13009 -1538 -12975
rect -1590 -13021 -1538 -13009
rect -960 -12873 -908 -12847
rect -960 -12907 -950 -12873
rect -916 -12907 -908 -12873
rect -960 -12975 -908 -12907
rect -960 -13009 -950 -12975
rect -916 -13009 -908 -12975
rect -960 -13021 -908 -13009
rect -854 -12873 -802 -12847
rect -854 -12907 -846 -12873
rect -812 -12907 -802 -12873
rect -854 -12975 -802 -12907
rect -854 -13009 -846 -12975
rect -812 -13009 -802 -12975
rect -854 -13021 -802 -13009
rect -224 -12873 -172 -12847
rect -224 -12907 -214 -12873
rect -180 -12907 -172 -12873
rect -224 -12975 -172 -12907
rect -224 -13009 -214 -12975
rect -180 -13009 -172 -12975
rect -26 -12873 26 -12847
rect -26 -12907 -18 -12873
rect 16 -12907 26 -12873
rect -26 -12975 26 -12907
rect -224 -13021 -172 -13009
rect -26 -13009 -18 -12975
rect 16 -13009 26 -12975
rect -26 -13021 26 -13009
rect 236 -12873 288 -12847
rect 236 -12907 246 -12873
rect 280 -12907 288 -12873
rect 236 -12975 288 -12907
rect 236 -13009 246 -12975
rect 280 -13009 288 -12975
rect 434 -12900 488 -12821
rect 434 -12934 443 -12900
rect 477 -12934 488 -12900
rect 434 -12968 488 -12934
rect 434 -13002 443 -12968
rect 477 -13002 488 -12968
rect 236 -13021 288 -13009
rect 434 -13021 488 -13002
rect 518 -12857 568 -12821
rect 965 -12857 1015 -12821
rect 518 -12900 590 -12857
rect 518 -12934 543 -12900
rect 577 -12934 590 -12900
rect 518 -12968 590 -12934
rect 518 -13002 543 -12968
rect 577 -13002 590 -12968
rect 518 -13021 590 -13002
rect 690 -12900 743 -12857
rect 690 -12934 701 -12900
rect 735 -12934 743 -12900
rect 690 -12968 743 -12934
rect 690 -13002 701 -12968
rect 735 -13002 743 -12968
rect 690 -13021 743 -13002
rect 797 -12899 850 -12857
rect 797 -12933 805 -12899
rect 839 -12933 850 -12899
rect 797 -12967 850 -12933
rect 797 -13001 805 -12967
rect 839 -13001 850 -12967
rect 797 -13021 850 -13001
rect 950 -12900 1015 -12857
rect 950 -12934 961 -12900
rect 995 -12934 1015 -12900
rect 950 -12968 1015 -12934
rect 950 -13002 961 -12968
rect 995 -13002 1015 -12968
rect 950 -13021 1015 -13002
rect 1045 -12899 1116 -12821
rect 1045 -12933 1059 -12899
rect 1093 -12933 1116 -12899
rect 1045 -12967 1116 -12933
rect 1045 -13001 1059 -12967
rect 1093 -13001 1116 -12967
rect 1045 -13021 1116 -13001
rect 1262 -12873 1314 -12847
rect 1262 -12907 1270 -12873
rect 1304 -12907 1314 -12873
rect 1262 -12975 1314 -12907
rect 1262 -13009 1270 -12975
rect 1304 -13009 1314 -12975
rect 1262 -13021 1314 -13009
rect 1524 -12873 1576 -12847
rect 1524 -12907 1534 -12873
rect 1568 -12907 1576 -12873
rect 1524 -12975 1576 -12907
rect 1524 -13009 1534 -12975
rect 1568 -13009 1576 -12975
rect 1722 -12873 1774 -12847
rect 1722 -12907 1730 -12873
rect 1764 -12907 1774 -12873
rect 1722 -12975 1774 -12907
rect 1524 -13021 1576 -13009
rect 1722 -13009 1730 -12975
rect 1764 -13009 1774 -12975
rect 1722 -13021 1774 -13009
rect 2352 -12873 2404 -12847
rect 2352 -12907 2362 -12873
rect 2396 -12907 2404 -12873
rect 2352 -12975 2404 -12907
rect 2352 -13009 2362 -12975
rect 2396 -13009 2404 -12975
rect 2550 -12873 2602 -12847
rect 2550 -12907 2558 -12873
rect 2592 -12907 2602 -12873
rect 2550 -12975 2602 -12907
rect 2352 -13021 2404 -13009
rect 2550 -13009 2558 -12975
rect 2592 -13009 2602 -12975
rect 2550 -13021 2602 -13009
rect 2812 -12873 2864 -12847
rect 2812 -12907 2822 -12873
rect 2856 -12907 2864 -12873
rect 2812 -12975 2864 -12907
rect 2812 -13009 2822 -12975
rect 2856 -13009 2864 -12975
rect 3010 -12900 3064 -12821
rect 3010 -12934 3019 -12900
rect 3053 -12934 3064 -12900
rect 3010 -12968 3064 -12934
rect 3010 -13002 3019 -12968
rect 3053 -13002 3064 -12968
rect 2812 -13021 2864 -13009
rect 3010 -13021 3064 -13002
rect 3094 -12857 3144 -12821
rect 3541 -12857 3591 -12821
rect 3094 -12900 3166 -12857
rect 3094 -12934 3119 -12900
rect 3153 -12934 3166 -12900
rect 3094 -12968 3166 -12934
rect 3094 -13002 3119 -12968
rect 3153 -13002 3166 -12968
rect 3094 -13021 3166 -13002
rect 3266 -12900 3319 -12857
rect 3266 -12934 3277 -12900
rect 3311 -12934 3319 -12900
rect 3266 -12968 3319 -12934
rect 3266 -13002 3277 -12968
rect 3311 -13002 3319 -12968
rect 3266 -13021 3319 -13002
rect 3373 -12899 3426 -12857
rect 3373 -12933 3381 -12899
rect 3415 -12933 3426 -12899
rect 3373 -12967 3426 -12933
rect 3373 -13001 3381 -12967
rect 3415 -13001 3426 -12967
rect 3373 -13021 3426 -13001
rect 3526 -12900 3591 -12857
rect 3526 -12934 3537 -12900
rect 3571 -12934 3591 -12900
rect 3526 -12968 3591 -12934
rect 3526 -13002 3537 -12968
rect 3571 -13002 3591 -12968
rect 3526 -13021 3591 -13002
rect 3621 -12899 3692 -12821
rect 3621 -12933 3635 -12899
rect 3669 -12933 3692 -12899
rect 3621 -12967 3692 -12933
rect 3621 -13001 3635 -12967
rect 3669 -13001 3692 -12967
rect 3621 -13021 3692 -13001
rect 3838 -12873 3890 -12847
rect 3838 -12907 3846 -12873
rect 3880 -12907 3890 -12873
rect 3838 -12975 3890 -12907
rect 3838 -13009 3846 -12975
rect 3880 -13009 3890 -12975
rect 3838 -13021 3890 -13009
rect 4100 -12873 4152 -12847
rect 4100 -12907 4110 -12873
rect 4144 -12907 4152 -12873
rect 4100 -12975 4152 -12907
rect 4100 -13009 4110 -12975
rect 4144 -13009 4152 -12975
rect 4298 -12873 4350 -12847
rect 4298 -12907 4306 -12873
rect 4340 -12907 4350 -12873
rect 4298 -12975 4350 -12907
rect 4100 -13021 4152 -13009
rect 4298 -13009 4306 -12975
rect 4340 -13009 4350 -12975
rect 4298 -13021 4350 -13009
rect 4928 -12873 4980 -12847
rect 4928 -12907 4938 -12873
rect 4972 -12907 4980 -12873
rect 4928 -12975 4980 -12907
rect 4928 -13009 4938 -12975
rect 4972 -13009 4980 -12975
rect 5126 -12873 5178 -12847
rect 5126 -12907 5134 -12873
rect 5168 -12907 5178 -12873
rect 5126 -12975 5178 -12907
rect 4928 -13021 4980 -13009
rect 5126 -13009 5134 -12975
rect 5168 -13009 5178 -12975
rect 5126 -13021 5178 -13009
rect 5388 -12873 5440 -12847
rect 5388 -12907 5398 -12873
rect 5432 -12907 5440 -12873
rect 5388 -12975 5440 -12907
rect 5388 -13009 5398 -12975
rect 5432 -13009 5440 -12975
rect 5586 -12900 5640 -12821
rect 5586 -12934 5595 -12900
rect 5629 -12934 5640 -12900
rect 5586 -12968 5640 -12934
rect 5586 -13002 5595 -12968
rect 5629 -13002 5640 -12968
rect 5388 -13021 5440 -13009
rect 5586 -13021 5640 -13002
rect 5670 -12857 5720 -12821
rect 6117 -12857 6167 -12821
rect 5670 -12900 5742 -12857
rect 5670 -12934 5695 -12900
rect 5729 -12934 5742 -12900
rect 5670 -12968 5742 -12934
rect 5670 -13002 5695 -12968
rect 5729 -13002 5742 -12968
rect 5670 -13021 5742 -13002
rect 5842 -12900 5895 -12857
rect 5842 -12934 5853 -12900
rect 5887 -12934 5895 -12900
rect 5842 -12968 5895 -12934
rect 5842 -13002 5853 -12968
rect 5887 -13002 5895 -12968
rect 5842 -13021 5895 -13002
rect 5949 -12899 6002 -12857
rect 5949 -12933 5957 -12899
rect 5991 -12933 6002 -12899
rect 5949 -12967 6002 -12933
rect 5949 -13001 5957 -12967
rect 5991 -13001 6002 -12967
rect 5949 -13021 6002 -13001
rect 6102 -12900 6167 -12857
rect 6102 -12934 6113 -12900
rect 6147 -12934 6167 -12900
rect 6102 -12968 6167 -12934
rect 6102 -13002 6113 -12968
rect 6147 -13002 6167 -12968
rect 6102 -13021 6167 -13002
rect 6197 -12899 6268 -12821
rect 6197 -12933 6211 -12899
rect 6245 -12933 6268 -12899
rect 6197 -12967 6268 -12933
rect 6197 -13001 6211 -12967
rect 6245 -13001 6268 -12967
rect 6197 -13021 6268 -13001
rect 6414 -12873 6466 -12847
rect 6414 -12907 6422 -12873
rect 6456 -12907 6466 -12873
rect 6414 -12975 6466 -12907
rect 6414 -13009 6422 -12975
rect 6456 -13009 6466 -12975
rect 6414 -13021 6466 -13009
rect 6676 -12873 6728 -12847
rect 6676 -12907 6686 -12873
rect 6720 -12907 6728 -12873
rect 6676 -12975 6728 -12907
rect 6676 -13009 6686 -12975
rect 6720 -13009 6728 -12975
rect 6874 -12873 6926 -12847
rect 6874 -12907 6882 -12873
rect 6916 -12907 6926 -12873
rect 6874 -12975 6926 -12907
rect 6676 -13021 6728 -13009
rect 6874 -13009 6882 -12975
rect 6916 -13009 6926 -12975
rect 6874 -13021 6926 -13009
rect 7504 -12873 7556 -12847
rect 7504 -12907 7514 -12873
rect 7548 -12907 7556 -12873
rect 7504 -12975 7556 -12907
rect 7504 -13009 7514 -12975
rect 7548 -13009 7556 -12975
rect 7702 -12873 7754 -12847
rect 7702 -12907 7710 -12873
rect 7744 -12907 7754 -12873
rect 7702 -12975 7754 -12907
rect 7504 -13021 7556 -13009
rect 7702 -13009 7710 -12975
rect 7744 -13009 7754 -12975
rect 7702 -13021 7754 -13009
rect 7964 -12873 8016 -12847
rect 7964 -12907 7974 -12873
rect 8008 -12907 8016 -12873
rect 7964 -12975 8016 -12907
rect 7964 -13009 7974 -12975
rect 8008 -13009 8016 -12975
rect 8162 -12900 8216 -12821
rect 8162 -12934 8171 -12900
rect 8205 -12934 8216 -12900
rect 8162 -12968 8216 -12934
rect 8162 -13002 8171 -12968
rect 8205 -13002 8216 -12968
rect 7964 -13021 8016 -13009
rect 8162 -13021 8216 -13002
rect 8246 -12857 8296 -12821
rect 8693 -12857 8743 -12821
rect 8246 -12900 8318 -12857
rect 8246 -12934 8271 -12900
rect 8305 -12934 8318 -12900
rect 8246 -12968 8318 -12934
rect 8246 -13002 8271 -12968
rect 8305 -13002 8318 -12968
rect 8246 -13021 8318 -13002
rect 8418 -12900 8471 -12857
rect 8418 -12934 8429 -12900
rect 8463 -12934 8471 -12900
rect 8418 -12968 8471 -12934
rect 8418 -13002 8429 -12968
rect 8463 -13002 8471 -12968
rect 8418 -13021 8471 -13002
rect 8525 -12899 8578 -12857
rect 8525 -12933 8533 -12899
rect 8567 -12933 8578 -12899
rect 8525 -12967 8578 -12933
rect 8525 -13001 8533 -12967
rect 8567 -13001 8578 -12967
rect 8525 -13021 8578 -13001
rect 8678 -12900 8743 -12857
rect 8678 -12934 8689 -12900
rect 8723 -12934 8743 -12900
rect 8678 -12968 8743 -12934
rect 8678 -13002 8689 -12968
rect 8723 -13002 8743 -12968
rect 8678 -13021 8743 -13002
rect 8773 -12899 8844 -12821
rect 8773 -12933 8787 -12899
rect 8821 -12933 8844 -12899
rect 8773 -12967 8844 -12933
rect 8773 -13001 8787 -12967
rect 8821 -13001 8844 -12967
rect 8773 -13021 8844 -13001
rect 8990 -12873 9042 -12847
rect 8990 -12907 8998 -12873
rect 9032 -12907 9042 -12873
rect 8990 -12975 9042 -12907
rect 8990 -13009 8998 -12975
rect 9032 -13009 9042 -12975
rect 8990 -13021 9042 -13009
rect 9252 -12873 9304 -12847
rect 9252 -12907 9262 -12873
rect 9296 -12907 9304 -12873
rect 9252 -12975 9304 -12907
rect 9252 -13009 9262 -12975
rect 9296 -13009 9304 -12975
rect 9450 -12873 9502 -12847
rect 9450 -12907 9458 -12873
rect 9492 -12907 9502 -12873
rect 9450 -12975 9502 -12907
rect 9252 -13021 9304 -13009
rect 9450 -13009 9458 -12975
rect 9492 -13009 9502 -12975
rect 9450 -13021 9502 -13009
rect 10080 -12873 10132 -12847
rect 10080 -12907 10090 -12873
rect 10124 -12907 10132 -12873
rect 10080 -12975 10132 -12907
rect 10080 -13009 10090 -12975
rect 10124 -13009 10132 -12975
rect 10370 -12873 10422 -12847
rect 10370 -12907 10378 -12873
rect 10412 -12907 10422 -12873
rect 10370 -12975 10422 -12907
rect 10080 -13021 10132 -13009
rect 10370 -13009 10378 -12975
rect 10412 -13009 10422 -12975
rect 10370 -13021 10422 -13009
rect 10632 -12873 10684 -12847
rect 10632 -12907 10642 -12873
rect 10676 -12907 10684 -12873
rect 10632 -12975 10684 -12907
rect 10632 -13009 10642 -12975
rect 10676 -13009 10684 -12975
rect 10632 -13021 10684 -13009
rect 10738 -12900 10792 -12821
rect 10738 -12934 10747 -12900
rect 10781 -12934 10792 -12900
rect 10738 -12968 10792 -12934
rect 10738 -13002 10747 -12968
rect 10781 -13002 10792 -12968
rect 10738 -13021 10792 -13002
rect 10822 -12857 10872 -12821
rect 11269 -12857 11319 -12821
rect 10822 -12900 10894 -12857
rect 10822 -12934 10847 -12900
rect 10881 -12934 10894 -12900
rect 10822 -12968 10894 -12934
rect 10822 -13002 10847 -12968
rect 10881 -13002 10894 -12968
rect 10822 -13021 10894 -13002
rect 10994 -12900 11047 -12857
rect 10994 -12934 11005 -12900
rect 11039 -12934 11047 -12900
rect 10994 -12968 11047 -12934
rect 10994 -13002 11005 -12968
rect 11039 -13002 11047 -12968
rect 10994 -13021 11047 -13002
rect 11101 -12899 11154 -12857
rect 11101 -12933 11109 -12899
rect 11143 -12933 11154 -12899
rect 11101 -12967 11154 -12933
rect 11101 -13001 11109 -12967
rect 11143 -13001 11154 -12967
rect 11101 -13021 11154 -13001
rect 11254 -12900 11319 -12857
rect 11254 -12934 11265 -12900
rect 11299 -12934 11319 -12900
rect 11254 -12968 11319 -12934
rect 11254 -13002 11265 -12968
rect 11299 -13002 11319 -12968
rect 11254 -13021 11319 -13002
rect 11349 -12899 11420 -12821
rect 11349 -12933 11363 -12899
rect 11397 -12933 11420 -12899
rect 11349 -12967 11420 -12933
rect 11349 -13001 11363 -12967
rect 11397 -13001 11420 -12967
rect 11349 -13021 11420 -13001
rect 11658 -12873 11710 -12847
rect 11658 -12907 11666 -12873
rect 11700 -12907 11710 -12873
rect 11658 -12975 11710 -12907
rect 11658 -13009 11666 -12975
rect 11700 -13009 11710 -12975
rect 11658 -13021 11710 -13009
rect 11920 -12873 11972 -12847
rect 11920 -12907 11930 -12873
rect 11964 -12907 11972 -12873
rect 11920 -12975 11972 -12907
rect 11920 -13009 11930 -12975
rect 11964 -13009 11972 -12975
rect 12486 -12900 12547 -12821
rect 12486 -12934 12502 -12900
rect 12536 -12934 12547 -12900
rect 12486 -12968 12547 -12934
rect 12486 -13002 12502 -12968
rect 12536 -13002 12547 -12968
rect 11920 -13021 11972 -13009
rect 12486 -13021 12547 -13002
rect 12577 -12873 12633 -12821
rect 12577 -12907 12588 -12873
rect 12622 -12907 12633 -12873
rect 12577 -12961 12633 -12907
rect 12577 -12995 12588 -12961
rect 12622 -12995 12633 -12961
rect 12577 -13021 12633 -12995
rect 12663 -12900 12719 -12821
rect 12663 -12934 12674 -12900
rect 12708 -12934 12719 -12900
rect 12663 -12968 12719 -12934
rect 12663 -13002 12674 -12968
rect 12708 -13002 12719 -12968
rect 12663 -13021 12719 -13002
rect 12749 -12873 12805 -12821
rect 12749 -12907 12760 -12873
rect 12794 -12907 12805 -12873
rect 12749 -12961 12805 -12907
rect 12749 -12995 12760 -12961
rect 12794 -12995 12805 -12961
rect 12749 -13021 12805 -12995
rect 12835 -12900 12891 -12821
rect 12835 -12934 12846 -12900
rect 12880 -12934 12891 -12900
rect 12835 -12968 12891 -12934
rect 12835 -13002 12846 -12968
rect 12880 -13002 12891 -12968
rect 12835 -13021 12891 -13002
rect 12921 -12873 12977 -12821
rect 12921 -12907 12932 -12873
rect 12966 -12907 12977 -12873
rect 12921 -12961 12977 -12907
rect 12921 -12995 12932 -12961
rect 12966 -12995 12977 -12961
rect 12921 -13021 12977 -12995
rect 13007 -12900 13076 -12821
rect 13007 -12934 13018 -12900
rect 13052 -12934 13076 -12900
rect 13007 -12968 13076 -12934
rect 13007 -13002 13018 -12968
rect 13052 -13002 13076 -12968
rect 13007 -13021 13076 -13002
rect 13222 -12873 13274 -12847
rect 13222 -12907 13230 -12873
rect 13264 -12907 13274 -12873
rect 13222 -12975 13274 -12907
rect 13222 -13009 13230 -12975
rect 13264 -13009 13274 -12975
rect 13222 -13021 13274 -13009
rect 13484 -12873 13536 -12847
rect 13484 -12907 13494 -12873
rect 13528 -12907 13536 -12873
rect 13484 -12975 13536 -12907
rect 13484 -13009 13494 -12975
rect 13528 -13009 13536 -12975
rect 13682 -12907 13735 -12821
rect 13682 -12941 13690 -12907
rect 13724 -12941 13735 -12907
rect 13682 -12975 13735 -12941
rect 13484 -13021 13536 -13009
rect 13682 -13009 13690 -12975
rect 13724 -13009 13735 -12975
rect 13682 -13021 13735 -13009
rect 13765 -12899 13821 -12821
rect 13765 -12933 13776 -12899
rect 13810 -12933 13821 -12899
rect 13765 -12967 13821 -12933
rect 13765 -13001 13776 -12967
rect 13810 -13001 13821 -12967
rect 13765 -13021 13821 -13001
rect 13851 -12907 13907 -12821
rect 13851 -12941 13862 -12907
rect 13896 -12941 13907 -12907
rect 13851 -12975 13907 -12941
rect 13851 -13009 13862 -12975
rect 13896 -13009 13907 -12975
rect 13851 -13021 13907 -13009
rect 13937 -12891 13993 -12821
rect 13937 -12925 13948 -12891
rect 13982 -12925 13993 -12891
rect 13937 -12959 13993 -12925
rect 13937 -12993 13948 -12959
rect 13982 -12993 13993 -12959
rect 13937 -13021 13993 -12993
rect 14023 -12907 14079 -12821
rect 14023 -12941 14034 -12907
rect 14068 -12941 14079 -12907
rect 14023 -12975 14079 -12941
rect 14023 -13009 14034 -12975
rect 14068 -13009 14079 -12975
rect 14023 -13021 14079 -13009
rect 14109 -12845 14165 -12821
rect 14109 -12879 14120 -12845
rect 14154 -12879 14165 -12845
rect 14109 -12931 14165 -12879
rect 14109 -12965 14120 -12931
rect 14154 -12965 14165 -12931
rect 14109 -13021 14165 -12965
rect 14195 -12951 14251 -12821
rect 14195 -12985 14206 -12951
rect 14240 -12985 14251 -12951
rect 14195 -13021 14251 -12985
rect 14281 -12845 14337 -12821
rect 14281 -12879 14292 -12845
rect 14326 -12879 14337 -12845
rect 14281 -12931 14337 -12879
rect 14281 -12965 14292 -12931
rect 14326 -12965 14337 -12931
rect 14281 -13021 14337 -12965
rect 14367 -12951 14423 -12821
rect 14367 -12985 14378 -12951
rect 14412 -12985 14423 -12951
rect 14367 -13021 14423 -12985
rect 14453 -12845 14509 -12821
rect 14453 -12879 14464 -12845
rect 14498 -12879 14509 -12845
rect 14453 -12931 14509 -12879
rect 14453 -12965 14464 -12931
rect 14498 -12965 14509 -12931
rect 14453 -13021 14509 -12965
rect 14539 -12951 14595 -12821
rect 14539 -12985 14550 -12951
rect 14584 -12985 14595 -12951
rect 14539 -13021 14595 -12985
rect 14625 -12845 14681 -12821
rect 14625 -12879 14636 -12845
rect 14670 -12879 14681 -12845
rect 14625 -12931 14681 -12879
rect 14625 -12965 14636 -12931
rect 14670 -12965 14681 -12931
rect 14625 -13021 14681 -12965
rect 14711 -12951 14766 -12821
rect 14711 -12985 14722 -12951
rect 14756 -12985 14766 -12951
rect 14711 -13021 14766 -12985
rect 14796 -12845 14852 -12821
rect 14796 -12879 14807 -12845
rect 14841 -12879 14852 -12845
rect 14796 -12931 14852 -12879
rect 14796 -12965 14807 -12931
rect 14841 -12965 14852 -12931
rect 14796 -13021 14852 -12965
rect 14882 -12951 14938 -12821
rect 14882 -12985 14893 -12951
rect 14927 -12985 14938 -12951
rect 14882 -13021 14938 -12985
rect 14968 -12845 15024 -12821
rect 14968 -12879 14979 -12845
rect 15013 -12879 15024 -12845
rect 14968 -12931 15024 -12879
rect 14968 -12965 14979 -12931
rect 15013 -12965 15024 -12931
rect 14968 -13021 15024 -12965
rect 15054 -12951 15110 -12821
rect 15054 -12985 15065 -12951
rect 15099 -12985 15110 -12951
rect 15054 -13021 15110 -12985
rect 15140 -12845 15196 -12821
rect 15140 -12879 15151 -12845
rect 15185 -12879 15196 -12845
rect 15140 -12931 15196 -12879
rect 15140 -12965 15151 -12931
rect 15185 -12965 15196 -12931
rect 15140 -13021 15196 -12965
rect 15226 -12951 15282 -12821
rect 15226 -12985 15237 -12951
rect 15271 -12985 15282 -12951
rect 15226 -13021 15282 -12985
rect 15312 -12845 15368 -12821
rect 15312 -12879 15323 -12845
rect 15357 -12879 15368 -12845
rect 15312 -12931 15368 -12879
rect 15312 -12965 15323 -12931
rect 15357 -12965 15368 -12931
rect 15312 -13021 15368 -12965
rect 15398 -12951 15451 -12821
rect 15398 -12985 15409 -12951
rect 15443 -12985 15451 -12951
rect 15398 -13021 15451 -12985
rect 15614 -12873 15666 -12847
rect 15614 -12907 15622 -12873
rect 15656 -12907 15666 -12873
rect 15614 -12975 15666 -12907
rect 15614 -13009 15622 -12975
rect 15656 -13009 15666 -12975
rect 15614 -13021 15666 -13009
rect 16612 -12873 16664 -12847
rect 16612 -12907 16622 -12873
rect 16656 -12907 16664 -12873
rect 16612 -12975 16664 -12907
rect 16612 -13009 16622 -12975
rect 16656 -13009 16664 -12975
rect 16612 -13021 16664 -13009
rect -2970 -13127 -2918 -13115
rect -2970 -13161 -2962 -13127
rect -2928 -13161 -2918 -13127
rect -2970 -13229 -2918 -13161
rect -2970 -13263 -2962 -13229
rect -2928 -13263 -2918 -13229
rect -2970 -13289 -2918 -13263
rect -2340 -13127 -2288 -13115
rect -2340 -13161 -2330 -13127
rect -2296 -13161 -2288 -13127
rect -1590 -13127 -1538 -13115
rect -2340 -13229 -2288 -13161
rect -2340 -13263 -2330 -13229
rect -2296 -13263 -2288 -13229
rect -2340 -13289 -2288 -13263
rect -1590 -13161 -1582 -13127
rect -1548 -13161 -1538 -13127
rect -1590 -13229 -1538 -13161
rect -1590 -13263 -1582 -13229
rect -1548 -13263 -1538 -13229
rect -1590 -13289 -1538 -13263
rect -960 -13127 -908 -13115
rect -960 -13161 -950 -13127
rect -916 -13161 -908 -13127
rect -960 -13229 -908 -13161
rect -960 -13263 -950 -13229
rect -916 -13263 -908 -13229
rect -960 -13289 -908 -13263
rect -854 -13127 -802 -13115
rect -854 -13161 -846 -13127
rect -812 -13161 -802 -13127
rect -854 -13229 -802 -13161
rect -854 -13263 -846 -13229
rect -812 -13263 -802 -13229
rect -854 -13289 -802 -13263
rect -224 -13127 -172 -13115
rect -224 -13161 -214 -13127
rect -180 -13161 -172 -13127
rect -26 -13127 26 -13115
rect -224 -13229 -172 -13161
rect -224 -13263 -214 -13229
rect -180 -13263 -172 -13229
rect -224 -13289 -172 -13263
rect -26 -13161 -18 -13127
rect 16 -13161 26 -13127
rect -26 -13229 26 -13161
rect -26 -13263 -18 -13229
rect 16 -13263 26 -13229
rect -26 -13289 26 -13263
rect 236 -13127 288 -13115
rect 236 -13161 246 -13127
rect 280 -13161 288 -13127
rect 236 -13229 288 -13161
rect 236 -13263 246 -13229
rect 280 -13263 288 -13229
rect 236 -13289 288 -13263
rect 434 -13135 505 -13115
rect 434 -13169 457 -13135
rect 491 -13169 505 -13135
rect 434 -13203 505 -13169
rect 434 -13237 457 -13203
rect 491 -13237 505 -13203
rect 434 -13315 505 -13237
rect 535 -13134 600 -13115
rect 535 -13168 555 -13134
rect 589 -13168 600 -13134
rect 535 -13202 600 -13168
rect 535 -13236 555 -13202
rect 589 -13236 600 -13202
rect 535 -13279 600 -13236
rect 700 -13135 753 -13115
rect 700 -13169 711 -13135
rect 745 -13169 753 -13135
rect 700 -13203 753 -13169
rect 700 -13237 711 -13203
rect 745 -13237 753 -13203
rect 700 -13279 753 -13237
rect 807 -13134 860 -13115
rect 807 -13168 815 -13134
rect 849 -13168 860 -13134
rect 807 -13202 860 -13168
rect 807 -13236 815 -13202
rect 849 -13236 860 -13202
rect 807 -13279 860 -13236
rect 960 -13134 1032 -13115
rect 960 -13168 973 -13134
rect 1007 -13168 1032 -13134
rect 960 -13202 1032 -13168
rect 960 -13236 973 -13202
rect 1007 -13236 1032 -13202
rect 960 -13279 1032 -13236
rect 535 -13315 585 -13279
rect 982 -13315 1032 -13279
rect 1062 -13134 1116 -13115
rect 1262 -13127 1314 -13115
rect 1062 -13168 1073 -13134
rect 1107 -13168 1116 -13134
rect 1062 -13202 1116 -13168
rect 1062 -13236 1073 -13202
rect 1107 -13236 1116 -13202
rect 1062 -13315 1116 -13236
rect 1262 -13161 1270 -13127
rect 1304 -13161 1314 -13127
rect 1262 -13229 1314 -13161
rect 1262 -13263 1270 -13229
rect 1304 -13263 1314 -13229
rect 1262 -13289 1314 -13263
rect 1524 -13127 1576 -13115
rect 1524 -13161 1534 -13127
rect 1568 -13161 1576 -13127
rect 1722 -13127 1774 -13115
rect 1524 -13229 1576 -13161
rect 1524 -13263 1534 -13229
rect 1568 -13263 1576 -13229
rect 1524 -13289 1576 -13263
rect 1722 -13161 1730 -13127
rect 1764 -13161 1774 -13127
rect 1722 -13229 1774 -13161
rect 1722 -13263 1730 -13229
rect 1764 -13263 1774 -13229
rect 1722 -13289 1774 -13263
rect 2352 -13127 2404 -13115
rect 2352 -13161 2362 -13127
rect 2396 -13161 2404 -13127
rect 2550 -13127 2602 -13115
rect 2352 -13229 2404 -13161
rect 2352 -13263 2362 -13229
rect 2396 -13263 2404 -13229
rect 2352 -13289 2404 -13263
rect 2550 -13161 2558 -13127
rect 2592 -13161 2602 -13127
rect 2550 -13229 2602 -13161
rect 2550 -13263 2558 -13229
rect 2592 -13263 2602 -13229
rect 2550 -13289 2602 -13263
rect 2812 -13127 2864 -13115
rect 2812 -13161 2822 -13127
rect 2856 -13161 2864 -13127
rect 2812 -13229 2864 -13161
rect 2812 -13263 2822 -13229
rect 2856 -13263 2864 -13229
rect 2812 -13289 2864 -13263
rect 3010 -13135 3081 -13115
rect 3010 -13169 3033 -13135
rect 3067 -13169 3081 -13135
rect 3010 -13203 3081 -13169
rect 3010 -13237 3033 -13203
rect 3067 -13237 3081 -13203
rect 3010 -13315 3081 -13237
rect 3111 -13134 3176 -13115
rect 3111 -13168 3131 -13134
rect 3165 -13168 3176 -13134
rect 3111 -13202 3176 -13168
rect 3111 -13236 3131 -13202
rect 3165 -13236 3176 -13202
rect 3111 -13279 3176 -13236
rect 3276 -13135 3329 -13115
rect 3276 -13169 3287 -13135
rect 3321 -13169 3329 -13135
rect 3276 -13203 3329 -13169
rect 3276 -13237 3287 -13203
rect 3321 -13237 3329 -13203
rect 3276 -13279 3329 -13237
rect 3383 -13134 3436 -13115
rect 3383 -13168 3391 -13134
rect 3425 -13168 3436 -13134
rect 3383 -13202 3436 -13168
rect 3383 -13236 3391 -13202
rect 3425 -13236 3436 -13202
rect 3383 -13279 3436 -13236
rect 3536 -13134 3608 -13115
rect 3536 -13168 3549 -13134
rect 3583 -13168 3608 -13134
rect 3536 -13202 3608 -13168
rect 3536 -13236 3549 -13202
rect 3583 -13236 3608 -13202
rect 3536 -13279 3608 -13236
rect 3111 -13315 3161 -13279
rect 3558 -13315 3608 -13279
rect 3638 -13134 3692 -13115
rect 3838 -13127 3890 -13115
rect 3638 -13168 3649 -13134
rect 3683 -13168 3692 -13134
rect 3638 -13202 3692 -13168
rect 3638 -13236 3649 -13202
rect 3683 -13236 3692 -13202
rect 3638 -13315 3692 -13236
rect 3838 -13161 3846 -13127
rect 3880 -13161 3890 -13127
rect 3838 -13229 3890 -13161
rect 3838 -13263 3846 -13229
rect 3880 -13263 3890 -13229
rect 3838 -13289 3890 -13263
rect 4100 -13127 4152 -13115
rect 4100 -13161 4110 -13127
rect 4144 -13161 4152 -13127
rect 4298 -13127 4350 -13115
rect 4100 -13229 4152 -13161
rect 4100 -13263 4110 -13229
rect 4144 -13263 4152 -13229
rect 4100 -13289 4152 -13263
rect 4298 -13161 4306 -13127
rect 4340 -13161 4350 -13127
rect 4298 -13229 4350 -13161
rect 4298 -13263 4306 -13229
rect 4340 -13263 4350 -13229
rect 4298 -13289 4350 -13263
rect 4928 -13127 4980 -13115
rect 4928 -13161 4938 -13127
rect 4972 -13161 4980 -13127
rect 5126 -13127 5178 -13115
rect 4928 -13229 4980 -13161
rect 4928 -13263 4938 -13229
rect 4972 -13263 4980 -13229
rect 4928 -13289 4980 -13263
rect 5126 -13161 5134 -13127
rect 5168 -13161 5178 -13127
rect 5126 -13229 5178 -13161
rect 5126 -13263 5134 -13229
rect 5168 -13263 5178 -13229
rect 5126 -13289 5178 -13263
rect 5388 -13127 5440 -13115
rect 5388 -13161 5398 -13127
rect 5432 -13161 5440 -13127
rect 5388 -13229 5440 -13161
rect 5388 -13263 5398 -13229
rect 5432 -13263 5440 -13229
rect 5388 -13289 5440 -13263
rect 5586 -13135 5657 -13115
rect 5586 -13169 5609 -13135
rect 5643 -13169 5657 -13135
rect 5586 -13203 5657 -13169
rect 5586 -13237 5609 -13203
rect 5643 -13237 5657 -13203
rect 5586 -13315 5657 -13237
rect 5687 -13134 5752 -13115
rect 5687 -13168 5707 -13134
rect 5741 -13168 5752 -13134
rect 5687 -13202 5752 -13168
rect 5687 -13236 5707 -13202
rect 5741 -13236 5752 -13202
rect 5687 -13279 5752 -13236
rect 5852 -13135 5905 -13115
rect 5852 -13169 5863 -13135
rect 5897 -13169 5905 -13135
rect 5852 -13203 5905 -13169
rect 5852 -13237 5863 -13203
rect 5897 -13237 5905 -13203
rect 5852 -13279 5905 -13237
rect 5959 -13134 6012 -13115
rect 5959 -13168 5967 -13134
rect 6001 -13168 6012 -13134
rect 5959 -13202 6012 -13168
rect 5959 -13236 5967 -13202
rect 6001 -13236 6012 -13202
rect 5959 -13279 6012 -13236
rect 6112 -13134 6184 -13115
rect 6112 -13168 6125 -13134
rect 6159 -13168 6184 -13134
rect 6112 -13202 6184 -13168
rect 6112 -13236 6125 -13202
rect 6159 -13236 6184 -13202
rect 6112 -13279 6184 -13236
rect 5687 -13315 5737 -13279
rect 6134 -13315 6184 -13279
rect 6214 -13134 6268 -13115
rect 6414 -13127 6466 -13115
rect 6214 -13168 6225 -13134
rect 6259 -13168 6268 -13134
rect 6214 -13202 6268 -13168
rect 6214 -13236 6225 -13202
rect 6259 -13236 6268 -13202
rect 6214 -13315 6268 -13236
rect 6414 -13161 6422 -13127
rect 6456 -13161 6466 -13127
rect 6414 -13229 6466 -13161
rect 6414 -13263 6422 -13229
rect 6456 -13263 6466 -13229
rect 6414 -13289 6466 -13263
rect 6676 -13127 6728 -13115
rect 6676 -13161 6686 -13127
rect 6720 -13161 6728 -13127
rect 6874 -13127 6926 -13115
rect 6676 -13229 6728 -13161
rect 6676 -13263 6686 -13229
rect 6720 -13263 6728 -13229
rect 6676 -13289 6728 -13263
rect 6874 -13161 6882 -13127
rect 6916 -13161 6926 -13127
rect 6874 -13229 6926 -13161
rect 6874 -13263 6882 -13229
rect 6916 -13263 6926 -13229
rect 6874 -13289 6926 -13263
rect 7504 -13127 7556 -13115
rect 7504 -13161 7514 -13127
rect 7548 -13161 7556 -13127
rect 7702 -13127 7754 -13115
rect 7504 -13229 7556 -13161
rect 7504 -13263 7514 -13229
rect 7548 -13263 7556 -13229
rect 7504 -13289 7556 -13263
rect 7702 -13161 7710 -13127
rect 7744 -13161 7754 -13127
rect 7702 -13229 7754 -13161
rect 7702 -13263 7710 -13229
rect 7744 -13263 7754 -13229
rect 7702 -13289 7754 -13263
rect 7964 -13127 8016 -13115
rect 7964 -13161 7974 -13127
rect 8008 -13161 8016 -13127
rect 7964 -13229 8016 -13161
rect 7964 -13263 7974 -13229
rect 8008 -13263 8016 -13229
rect 7964 -13289 8016 -13263
rect 8162 -13135 8233 -13115
rect 8162 -13169 8185 -13135
rect 8219 -13169 8233 -13135
rect 8162 -13203 8233 -13169
rect 8162 -13237 8185 -13203
rect 8219 -13237 8233 -13203
rect 8162 -13315 8233 -13237
rect 8263 -13134 8328 -13115
rect 8263 -13168 8283 -13134
rect 8317 -13168 8328 -13134
rect 8263 -13202 8328 -13168
rect 8263 -13236 8283 -13202
rect 8317 -13236 8328 -13202
rect 8263 -13279 8328 -13236
rect 8428 -13135 8481 -13115
rect 8428 -13169 8439 -13135
rect 8473 -13169 8481 -13135
rect 8428 -13203 8481 -13169
rect 8428 -13237 8439 -13203
rect 8473 -13237 8481 -13203
rect 8428 -13279 8481 -13237
rect 8535 -13134 8588 -13115
rect 8535 -13168 8543 -13134
rect 8577 -13168 8588 -13134
rect 8535 -13202 8588 -13168
rect 8535 -13236 8543 -13202
rect 8577 -13236 8588 -13202
rect 8535 -13279 8588 -13236
rect 8688 -13134 8760 -13115
rect 8688 -13168 8701 -13134
rect 8735 -13168 8760 -13134
rect 8688 -13202 8760 -13168
rect 8688 -13236 8701 -13202
rect 8735 -13236 8760 -13202
rect 8688 -13279 8760 -13236
rect 8263 -13315 8313 -13279
rect 8710 -13315 8760 -13279
rect 8790 -13134 8844 -13115
rect 8990 -13127 9042 -13115
rect 8790 -13168 8801 -13134
rect 8835 -13168 8844 -13134
rect 8790 -13202 8844 -13168
rect 8790 -13236 8801 -13202
rect 8835 -13236 8844 -13202
rect 8790 -13315 8844 -13236
rect 8990 -13161 8998 -13127
rect 9032 -13161 9042 -13127
rect 8990 -13229 9042 -13161
rect 8990 -13263 8998 -13229
rect 9032 -13263 9042 -13229
rect 8990 -13289 9042 -13263
rect 9252 -13127 9304 -13115
rect 9252 -13161 9262 -13127
rect 9296 -13161 9304 -13127
rect 9450 -13127 9502 -13115
rect 9252 -13229 9304 -13161
rect 9252 -13263 9262 -13229
rect 9296 -13263 9304 -13229
rect 9252 -13289 9304 -13263
rect 9450 -13161 9458 -13127
rect 9492 -13161 9502 -13127
rect 9450 -13229 9502 -13161
rect 9450 -13263 9458 -13229
rect 9492 -13263 9502 -13229
rect 9450 -13289 9502 -13263
rect 10080 -13127 10132 -13115
rect 10080 -13161 10090 -13127
rect 10124 -13161 10132 -13127
rect 10370 -13127 10422 -13115
rect 10080 -13229 10132 -13161
rect 10080 -13263 10090 -13229
rect 10124 -13263 10132 -13229
rect 10080 -13289 10132 -13263
rect 10370 -13161 10378 -13127
rect 10412 -13161 10422 -13127
rect 10370 -13229 10422 -13161
rect 10370 -13263 10378 -13229
rect 10412 -13263 10422 -13229
rect 10370 -13289 10422 -13263
rect 10632 -13127 10684 -13115
rect 10632 -13161 10642 -13127
rect 10676 -13161 10684 -13127
rect 10632 -13229 10684 -13161
rect 10632 -13263 10642 -13229
rect 10676 -13263 10684 -13229
rect 10632 -13289 10684 -13263
rect 10738 -13135 10809 -13115
rect 10738 -13169 10761 -13135
rect 10795 -13169 10809 -13135
rect 10738 -13203 10809 -13169
rect 10738 -13237 10761 -13203
rect 10795 -13237 10809 -13203
rect 10738 -13315 10809 -13237
rect 10839 -13134 10904 -13115
rect 10839 -13168 10859 -13134
rect 10893 -13168 10904 -13134
rect 10839 -13202 10904 -13168
rect 10839 -13236 10859 -13202
rect 10893 -13236 10904 -13202
rect 10839 -13279 10904 -13236
rect 11004 -13135 11057 -13115
rect 11004 -13169 11015 -13135
rect 11049 -13169 11057 -13135
rect 11004 -13203 11057 -13169
rect 11004 -13237 11015 -13203
rect 11049 -13237 11057 -13203
rect 11004 -13279 11057 -13237
rect 11111 -13134 11164 -13115
rect 11111 -13168 11119 -13134
rect 11153 -13168 11164 -13134
rect 11111 -13202 11164 -13168
rect 11111 -13236 11119 -13202
rect 11153 -13236 11164 -13202
rect 11111 -13279 11164 -13236
rect 11264 -13134 11336 -13115
rect 11264 -13168 11277 -13134
rect 11311 -13168 11336 -13134
rect 11264 -13202 11336 -13168
rect 11264 -13236 11277 -13202
rect 11311 -13236 11336 -13202
rect 11264 -13279 11336 -13236
rect 10839 -13315 10889 -13279
rect 11286 -13315 11336 -13279
rect 11366 -13134 11420 -13115
rect 11658 -13127 11710 -13115
rect 11366 -13168 11377 -13134
rect 11411 -13168 11420 -13134
rect 11366 -13202 11420 -13168
rect 11366 -13236 11377 -13202
rect 11411 -13236 11420 -13202
rect 11366 -13315 11420 -13236
rect 11658 -13161 11666 -13127
rect 11700 -13161 11710 -13127
rect 11658 -13229 11710 -13161
rect 11658 -13263 11666 -13229
rect 11700 -13263 11710 -13229
rect 11658 -13289 11710 -13263
rect 11920 -13127 11972 -13115
rect 11920 -13161 11930 -13127
rect 11964 -13161 11972 -13127
rect 13682 -13127 13735 -13115
rect 11920 -13229 11972 -13161
rect 11920 -13263 11930 -13229
rect 11964 -13263 11972 -13229
rect 11920 -13289 11972 -13263
rect 13682 -13161 13690 -13127
rect 13724 -13161 13735 -13127
rect 13682 -13195 13735 -13161
rect 13682 -13229 13690 -13195
rect 13724 -13229 13735 -13195
rect 13682 -13315 13735 -13229
rect 13765 -13135 13821 -13115
rect 13765 -13169 13776 -13135
rect 13810 -13169 13821 -13135
rect 13765 -13203 13821 -13169
rect 13765 -13237 13776 -13203
rect 13810 -13237 13821 -13203
rect 13765 -13315 13821 -13237
rect 13851 -13127 13907 -13115
rect 13851 -13161 13862 -13127
rect 13896 -13161 13907 -13127
rect 13851 -13195 13907 -13161
rect 13851 -13229 13862 -13195
rect 13896 -13229 13907 -13195
rect 13851 -13315 13907 -13229
rect 13937 -13143 13993 -13115
rect 13937 -13177 13948 -13143
rect 13982 -13177 13993 -13143
rect 13937 -13211 13993 -13177
rect 13937 -13245 13948 -13211
rect 13982 -13245 13993 -13211
rect 13937 -13315 13993 -13245
rect 14023 -13127 14079 -13115
rect 14023 -13161 14034 -13127
rect 14068 -13161 14079 -13127
rect 14023 -13195 14079 -13161
rect 14023 -13229 14034 -13195
rect 14068 -13229 14079 -13195
rect 14023 -13315 14079 -13229
rect 14109 -13171 14165 -13115
rect 14109 -13205 14120 -13171
rect 14154 -13205 14165 -13171
rect 14109 -13257 14165 -13205
rect 14109 -13291 14120 -13257
rect 14154 -13291 14165 -13257
rect 14109 -13315 14165 -13291
rect 14195 -13151 14251 -13115
rect 14195 -13185 14206 -13151
rect 14240 -13185 14251 -13151
rect 14195 -13315 14251 -13185
rect 14281 -13171 14337 -13115
rect 14281 -13205 14292 -13171
rect 14326 -13205 14337 -13171
rect 14281 -13257 14337 -13205
rect 14281 -13291 14292 -13257
rect 14326 -13291 14337 -13257
rect 14281 -13315 14337 -13291
rect 14367 -13151 14423 -13115
rect 14367 -13185 14378 -13151
rect 14412 -13185 14423 -13151
rect 14367 -13315 14423 -13185
rect 14453 -13171 14509 -13115
rect 14453 -13205 14464 -13171
rect 14498 -13205 14509 -13171
rect 14453 -13257 14509 -13205
rect 14453 -13291 14464 -13257
rect 14498 -13291 14509 -13257
rect 14453 -13315 14509 -13291
rect 14539 -13151 14595 -13115
rect 14539 -13185 14550 -13151
rect 14584 -13185 14595 -13151
rect 14539 -13315 14595 -13185
rect 14625 -13171 14681 -13115
rect 14625 -13205 14636 -13171
rect 14670 -13205 14681 -13171
rect 14625 -13257 14681 -13205
rect 14625 -13291 14636 -13257
rect 14670 -13291 14681 -13257
rect 14625 -13315 14681 -13291
rect 14711 -13151 14766 -13115
rect 14711 -13185 14722 -13151
rect 14756 -13185 14766 -13151
rect 14711 -13315 14766 -13185
rect 14796 -13171 14852 -13115
rect 14796 -13205 14807 -13171
rect 14841 -13205 14852 -13171
rect 14796 -13257 14852 -13205
rect 14796 -13291 14807 -13257
rect 14841 -13291 14852 -13257
rect 14796 -13315 14852 -13291
rect 14882 -13151 14938 -13115
rect 14882 -13185 14893 -13151
rect 14927 -13185 14938 -13151
rect 14882 -13315 14938 -13185
rect 14968 -13171 15024 -13115
rect 14968 -13205 14979 -13171
rect 15013 -13205 15024 -13171
rect 14968 -13257 15024 -13205
rect 14968 -13291 14979 -13257
rect 15013 -13291 15024 -13257
rect 14968 -13315 15024 -13291
rect 15054 -13151 15110 -13115
rect 15054 -13185 15065 -13151
rect 15099 -13185 15110 -13151
rect 15054 -13315 15110 -13185
rect 15140 -13171 15196 -13115
rect 15140 -13205 15151 -13171
rect 15185 -13205 15196 -13171
rect 15140 -13257 15196 -13205
rect 15140 -13291 15151 -13257
rect 15185 -13291 15196 -13257
rect 15140 -13315 15196 -13291
rect 15226 -13151 15282 -13115
rect 15226 -13185 15237 -13151
rect 15271 -13185 15282 -13151
rect 15226 -13315 15282 -13185
rect 15312 -13171 15368 -13115
rect 15312 -13205 15323 -13171
rect 15357 -13205 15368 -13171
rect 15312 -13257 15368 -13205
rect 15312 -13291 15323 -13257
rect 15357 -13291 15368 -13257
rect 15312 -13315 15368 -13291
rect 15398 -13151 15451 -13115
rect 15614 -13127 15666 -13115
rect 15398 -13185 15409 -13151
rect 15443 -13185 15451 -13151
rect 15398 -13315 15451 -13185
rect 15614 -13161 15622 -13127
rect 15656 -13161 15666 -13127
rect 15614 -13229 15666 -13161
rect 15614 -13263 15622 -13229
rect 15656 -13263 15666 -13229
rect 15614 -13289 15666 -13263
rect 16612 -13127 16664 -13115
rect 16612 -13161 16622 -13127
rect 16656 -13161 16664 -13127
rect 16612 -13229 16664 -13161
rect 16612 -13263 16622 -13229
rect 16656 -13263 16664 -13229
rect 16612 -13289 16664 -13263
rect -2970 -13961 -2918 -13935
rect -2970 -13995 -2962 -13961
rect -2928 -13995 -2918 -13961
rect -2970 -14063 -2918 -13995
rect -2970 -14097 -2962 -14063
rect -2928 -14097 -2918 -14063
rect -2970 -14109 -2918 -14097
rect -2340 -13961 -2288 -13935
rect -2340 -13995 -2330 -13961
rect -2296 -13995 -2288 -13961
rect -2340 -14063 -2288 -13995
rect -2340 -14097 -2330 -14063
rect -2296 -14097 -2288 -14063
rect -1406 -13961 -1354 -13935
rect -1406 -13995 -1398 -13961
rect -1364 -13995 -1354 -13961
rect -1406 -14063 -1354 -13995
rect -2340 -14109 -2288 -14097
rect -1406 -14097 -1398 -14063
rect -1364 -14097 -1354 -14063
rect -1406 -14109 -1354 -14097
rect -1144 -13961 -1092 -13935
rect -1144 -13995 -1134 -13961
rect -1100 -13995 -1092 -13961
rect -1144 -14063 -1092 -13995
rect -1144 -14097 -1134 -14063
rect -1100 -14097 -1092 -14063
rect -942 -13927 -890 -13909
rect -942 -13961 -934 -13927
rect -900 -13961 -890 -13927
rect -942 -13995 -890 -13961
rect -942 -14029 -934 -13995
rect -900 -14029 -890 -13995
rect -942 -14063 -890 -14029
rect -1144 -14109 -1092 -14097
rect -942 -14097 -934 -14063
rect -900 -14097 -890 -14063
rect -942 -14109 -890 -14097
rect -860 -13927 -806 -13909
rect -860 -13961 -850 -13927
rect -816 -13961 -806 -13927
rect -860 -13995 -806 -13961
rect -860 -14029 -850 -13995
rect -816 -14029 -806 -13995
rect -860 -14063 -806 -14029
rect -860 -14097 -850 -14063
rect -816 -14097 -806 -14063
rect -860 -14109 -806 -14097
rect -776 -13927 -724 -13909
rect -776 -13961 -766 -13927
rect -732 -13961 -724 -13927
rect -776 -13995 -724 -13961
rect -776 -14029 -766 -13995
rect -732 -14029 -724 -13995
rect -776 -14063 -724 -14029
rect -776 -14097 -766 -14063
rect -732 -14097 -724 -14063
rect -578 -13961 -526 -13935
rect -578 -13995 -570 -13961
rect -536 -13995 -526 -13961
rect -578 -14063 -526 -13995
rect -776 -14109 -724 -14097
rect -578 -14097 -570 -14063
rect -536 -14097 -526 -14063
rect -578 -14109 -526 -14097
rect -316 -13961 -264 -13935
rect -316 -13995 -306 -13961
rect -272 -13995 -264 -13961
rect -316 -14063 -264 -13995
rect -316 -14097 -306 -14063
rect -272 -14097 -264 -14063
rect -118 -13988 -57 -13909
rect -118 -14022 -102 -13988
rect -68 -14022 -57 -13988
rect -118 -14056 -57 -14022
rect -118 -14090 -102 -14056
rect -68 -14090 -57 -14056
rect -316 -14109 -264 -14097
rect -118 -14109 -57 -14090
rect -27 -13961 29 -13909
rect -27 -13995 -16 -13961
rect 18 -13995 29 -13961
rect -27 -14049 29 -13995
rect -27 -14083 -16 -14049
rect 18 -14083 29 -14049
rect -27 -14109 29 -14083
rect 59 -13988 115 -13909
rect 59 -14022 70 -13988
rect 104 -14022 115 -13988
rect 59 -14056 115 -14022
rect 59 -14090 70 -14056
rect 104 -14090 115 -14056
rect 59 -14109 115 -14090
rect 145 -13961 201 -13909
rect 145 -13995 156 -13961
rect 190 -13995 201 -13961
rect 145 -14049 201 -13995
rect 145 -14083 156 -14049
rect 190 -14083 201 -14049
rect 145 -14109 201 -14083
rect 231 -13988 287 -13909
rect 231 -14022 242 -13988
rect 276 -14022 287 -13988
rect 231 -14056 287 -14022
rect 231 -14090 242 -14056
rect 276 -14090 287 -14056
rect 231 -14109 287 -14090
rect 317 -13961 373 -13909
rect 317 -13995 328 -13961
rect 362 -13995 373 -13961
rect 317 -14049 373 -13995
rect 317 -14083 328 -14049
rect 362 -14083 373 -14049
rect 317 -14109 373 -14083
rect 403 -13988 472 -13909
rect 403 -14022 414 -13988
rect 448 -14022 472 -13988
rect 403 -14056 472 -14022
rect 403 -14090 414 -14056
rect 448 -14090 472 -14056
rect 403 -14109 472 -14090
rect 618 -13961 670 -13935
rect 618 -13995 626 -13961
rect 660 -13995 670 -13961
rect 618 -14063 670 -13995
rect 618 -14097 626 -14063
rect 660 -14097 670 -14063
rect 618 -14109 670 -14097
rect 880 -13961 932 -13935
rect 880 -13995 890 -13961
rect 924 -13995 932 -13961
rect 880 -14063 932 -13995
rect 880 -14097 890 -14063
rect 924 -14097 932 -14063
rect 1078 -13961 1130 -13941
rect 1078 -13995 1086 -13961
rect 1120 -13995 1130 -13961
rect 1078 -14063 1130 -13995
rect 880 -14109 932 -14097
rect 1078 -14097 1086 -14063
rect 1120 -14097 1130 -14063
rect 1078 -14109 1130 -14097
rect 1160 -13961 1214 -13941
rect 1160 -13995 1170 -13961
rect 1204 -13995 1214 -13961
rect 1160 -14063 1214 -13995
rect 1160 -14097 1170 -14063
rect 1204 -14097 1214 -14063
rect 1160 -14109 1214 -14097
rect 1244 -13961 1300 -13941
rect 1244 -13995 1254 -13961
rect 1288 -13995 1300 -13961
rect 1244 -14063 1300 -13995
rect 1244 -14097 1254 -14063
rect 1288 -14097 1300 -14063
rect 1446 -13961 1498 -13935
rect 1446 -13995 1454 -13961
rect 1488 -13995 1498 -13961
rect 1446 -14063 1498 -13995
rect 1244 -14109 1300 -14097
rect 1446 -14097 1454 -14063
rect 1488 -14097 1498 -14063
rect 1446 -14109 1498 -14097
rect 1708 -13961 1760 -13935
rect 1708 -13995 1718 -13961
rect 1752 -13995 1760 -13961
rect 1708 -14063 1760 -13995
rect 1708 -14097 1718 -14063
rect 1752 -14097 1760 -14063
rect 1906 -13961 1958 -13935
rect 1906 -13995 1914 -13961
rect 1948 -13995 1958 -13961
rect 1906 -14063 1958 -13995
rect 1708 -14109 1760 -14097
rect 1906 -14097 1914 -14063
rect 1948 -14097 1958 -14063
rect 1906 -14109 1958 -14097
rect 2168 -13961 2220 -13935
rect 2168 -13995 2178 -13961
rect 2212 -13995 2220 -13961
rect 2168 -14063 2220 -13995
rect 2168 -14097 2178 -14063
rect 2212 -14097 2220 -14063
rect 2366 -13988 2420 -13909
rect 2366 -14022 2375 -13988
rect 2409 -14022 2420 -13988
rect 2366 -14056 2420 -14022
rect 2366 -14090 2375 -14056
rect 2409 -14090 2420 -14056
rect 2168 -14109 2220 -14097
rect 2366 -14109 2420 -14090
rect 2450 -13945 2500 -13909
rect 2897 -13945 2947 -13909
rect 2450 -13988 2522 -13945
rect 2450 -14022 2475 -13988
rect 2509 -14022 2522 -13988
rect 2450 -14056 2522 -14022
rect 2450 -14090 2475 -14056
rect 2509 -14090 2522 -14056
rect 2450 -14109 2522 -14090
rect 2622 -13988 2675 -13945
rect 2622 -14022 2633 -13988
rect 2667 -14022 2675 -13988
rect 2622 -14056 2675 -14022
rect 2622 -14090 2633 -14056
rect 2667 -14090 2675 -14056
rect 2622 -14109 2675 -14090
rect 2729 -13987 2782 -13945
rect 2729 -14021 2737 -13987
rect 2771 -14021 2782 -13987
rect 2729 -14055 2782 -14021
rect 2729 -14089 2737 -14055
rect 2771 -14089 2782 -14055
rect 2729 -14109 2782 -14089
rect 2882 -13988 2947 -13945
rect 2882 -14022 2893 -13988
rect 2927 -14022 2947 -13988
rect 2882 -14056 2947 -14022
rect 2882 -14090 2893 -14056
rect 2927 -14090 2947 -14056
rect 2882 -14109 2947 -14090
rect 2977 -13987 3048 -13909
rect 2977 -14021 2991 -13987
rect 3025 -14021 3048 -13987
rect 2977 -14055 3048 -14021
rect 2977 -14089 2991 -14055
rect 3025 -14089 3048 -14055
rect 2977 -14109 3048 -14089
rect 3194 -13961 3246 -13935
rect 3194 -13995 3202 -13961
rect 3236 -13995 3246 -13961
rect 3194 -14063 3246 -13995
rect 3194 -14097 3202 -14063
rect 3236 -14097 3246 -14063
rect 3194 -14109 3246 -14097
rect 3456 -13961 3508 -13935
rect 3456 -13995 3466 -13961
rect 3500 -13995 3508 -13961
rect 3456 -14063 3508 -13995
rect 3456 -14097 3466 -14063
rect 3500 -14097 3508 -14063
rect 4390 -13961 4442 -13935
rect 4390 -13995 4398 -13961
rect 4432 -13995 4442 -13961
rect 4390 -14063 4442 -13995
rect 3456 -14109 3508 -14097
rect 4390 -14097 4398 -14063
rect 4432 -14097 4442 -14063
rect 4390 -14109 4442 -14097
rect 5388 -13961 5440 -13935
rect 5388 -13995 5398 -13961
rect 5432 -13995 5440 -13961
rect 5388 -14063 5440 -13995
rect 5388 -14097 5398 -14063
rect 5432 -14097 5440 -14063
rect 6414 -13961 6466 -13935
rect 6414 -13995 6422 -13961
rect 6456 -13995 6466 -13961
rect 6414 -14063 6466 -13995
rect 5388 -14109 5440 -14097
rect 6414 -14097 6422 -14063
rect 6456 -14097 6466 -14063
rect 6414 -14109 6466 -14097
rect 6676 -13961 6728 -13935
rect 6676 -13995 6686 -13961
rect 6720 -13995 6728 -13961
rect 6676 -14063 6728 -13995
rect 6676 -14097 6686 -14063
rect 6720 -14097 6728 -14063
rect 6874 -13988 6928 -13909
rect 6874 -14022 6883 -13988
rect 6917 -14022 6928 -13988
rect 6874 -14056 6928 -14022
rect 6874 -14090 6883 -14056
rect 6917 -14090 6928 -14056
rect 6676 -14109 6728 -14097
rect 6874 -14109 6928 -14090
rect 6958 -13945 7008 -13909
rect 7405 -13945 7455 -13909
rect 6958 -13988 7030 -13945
rect 6958 -14022 6983 -13988
rect 7017 -14022 7030 -13988
rect 6958 -14056 7030 -14022
rect 6958 -14090 6983 -14056
rect 7017 -14090 7030 -14056
rect 6958 -14109 7030 -14090
rect 7130 -13988 7183 -13945
rect 7130 -14022 7141 -13988
rect 7175 -14022 7183 -13988
rect 7130 -14056 7183 -14022
rect 7130 -14090 7141 -14056
rect 7175 -14090 7183 -14056
rect 7130 -14109 7183 -14090
rect 7237 -13987 7290 -13945
rect 7237 -14021 7245 -13987
rect 7279 -14021 7290 -13987
rect 7237 -14055 7290 -14021
rect 7237 -14089 7245 -14055
rect 7279 -14089 7290 -14055
rect 7237 -14109 7290 -14089
rect 7390 -13988 7455 -13945
rect 7390 -14022 7401 -13988
rect 7435 -14022 7455 -13988
rect 7390 -14056 7455 -14022
rect 7390 -14090 7401 -14056
rect 7435 -14090 7455 -14056
rect 7390 -14109 7455 -14090
rect 7485 -13987 7556 -13909
rect 7485 -14021 7499 -13987
rect 7533 -14021 7556 -13987
rect 7485 -14055 7556 -14021
rect 7485 -14089 7499 -14055
rect 7533 -14089 7556 -14055
rect 7485 -14109 7556 -14089
rect 7702 -13961 7754 -13935
rect 7702 -13995 7710 -13961
rect 7744 -13995 7754 -13961
rect 7702 -14063 7754 -13995
rect 7702 -14097 7710 -14063
rect 7744 -14097 7754 -14063
rect 7702 -14109 7754 -14097
rect 7964 -13961 8016 -13935
rect 7964 -13995 7974 -13961
rect 8008 -13995 8016 -13961
rect 7964 -14063 8016 -13995
rect 7964 -14097 7974 -14063
rect 8008 -14097 8016 -14063
rect 8162 -13988 8216 -13909
rect 8162 -14022 8171 -13988
rect 8205 -14022 8216 -13988
rect 8162 -14056 8216 -14022
rect 8162 -14090 8171 -14056
rect 8205 -14090 8216 -14056
rect 7964 -14109 8016 -14097
rect 8162 -14109 8216 -14090
rect 8246 -13945 8296 -13909
rect 8693 -13945 8743 -13909
rect 8246 -13988 8318 -13945
rect 8246 -14022 8271 -13988
rect 8305 -14022 8318 -13988
rect 8246 -14056 8318 -14022
rect 8246 -14090 8271 -14056
rect 8305 -14090 8318 -14056
rect 8246 -14109 8318 -14090
rect 8418 -13988 8471 -13945
rect 8418 -14022 8429 -13988
rect 8463 -14022 8471 -13988
rect 8418 -14056 8471 -14022
rect 8418 -14090 8429 -14056
rect 8463 -14090 8471 -14056
rect 8418 -14109 8471 -14090
rect 8525 -13987 8578 -13945
rect 8525 -14021 8533 -13987
rect 8567 -14021 8578 -13987
rect 8525 -14055 8578 -14021
rect 8525 -14089 8533 -14055
rect 8567 -14089 8578 -14055
rect 8525 -14109 8578 -14089
rect 8678 -13988 8743 -13945
rect 8678 -14022 8689 -13988
rect 8723 -14022 8743 -13988
rect 8678 -14056 8743 -14022
rect 8678 -14090 8689 -14056
rect 8723 -14090 8743 -14056
rect 8678 -14109 8743 -14090
rect 8773 -13987 8844 -13909
rect 8773 -14021 8787 -13987
rect 8821 -14021 8844 -13987
rect 8773 -14055 8844 -14021
rect 8773 -14089 8787 -14055
rect 8821 -14089 8844 -14055
rect 8773 -14109 8844 -14089
rect 8990 -13961 9042 -13935
rect 8990 -13995 8998 -13961
rect 9032 -13995 9042 -13961
rect 8990 -14063 9042 -13995
rect 8990 -14097 8998 -14063
rect 9032 -14097 9042 -14063
rect 8990 -14109 9042 -14097
rect 9252 -13961 9304 -13935
rect 9252 -13995 9262 -13961
rect 9296 -13995 9304 -13961
rect 9252 -14063 9304 -13995
rect 9252 -14097 9262 -14063
rect 9296 -14097 9304 -14063
rect 9450 -13988 9504 -13909
rect 9450 -14022 9459 -13988
rect 9493 -14022 9504 -13988
rect 9450 -14056 9504 -14022
rect 9450 -14090 9459 -14056
rect 9493 -14090 9504 -14056
rect 9252 -14109 9304 -14097
rect 9450 -14109 9504 -14090
rect 9534 -13945 9584 -13909
rect 9981 -13945 10031 -13909
rect 9534 -13988 9606 -13945
rect 9534 -14022 9559 -13988
rect 9593 -14022 9606 -13988
rect 9534 -14056 9606 -14022
rect 9534 -14090 9559 -14056
rect 9593 -14090 9606 -14056
rect 9534 -14109 9606 -14090
rect 9706 -13988 9759 -13945
rect 9706 -14022 9717 -13988
rect 9751 -14022 9759 -13988
rect 9706 -14056 9759 -14022
rect 9706 -14090 9717 -14056
rect 9751 -14090 9759 -14056
rect 9706 -14109 9759 -14090
rect 9813 -13987 9866 -13945
rect 9813 -14021 9821 -13987
rect 9855 -14021 9866 -13987
rect 9813 -14055 9866 -14021
rect 9813 -14089 9821 -14055
rect 9855 -14089 9866 -14055
rect 9813 -14109 9866 -14089
rect 9966 -13988 10031 -13945
rect 9966 -14022 9977 -13988
rect 10011 -14022 10031 -13988
rect 9966 -14056 10031 -14022
rect 9966 -14090 9977 -14056
rect 10011 -14090 10031 -14056
rect 9966 -14109 10031 -14090
rect 10061 -13987 10132 -13909
rect 10061 -14021 10075 -13987
rect 10109 -14021 10132 -13987
rect 10061 -14055 10132 -14021
rect 10061 -14089 10075 -14055
rect 10109 -14089 10132 -14055
rect 10061 -14109 10132 -14089
rect 10278 -13961 10330 -13935
rect 10278 -13995 10286 -13961
rect 10320 -13995 10330 -13961
rect 10278 -14063 10330 -13995
rect 10278 -14097 10286 -14063
rect 10320 -14097 10330 -14063
rect 10278 -14109 10330 -14097
rect 10540 -13961 10592 -13935
rect 10540 -13995 10550 -13961
rect 10584 -13995 10592 -13961
rect 10540 -14063 10592 -13995
rect 10540 -14097 10550 -14063
rect 10584 -14097 10592 -14063
rect 10738 -13927 10790 -13909
rect 10738 -13961 10746 -13927
rect 10780 -13961 10790 -13927
rect 10738 -13995 10790 -13961
rect 10738 -14029 10746 -13995
rect 10780 -14029 10790 -13995
rect 10738 -14063 10790 -14029
rect 10540 -14109 10592 -14097
rect 10738 -14097 10746 -14063
rect 10780 -14097 10790 -14063
rect 10738 -14109 10790 -14097
rect 10820 -13927 10874 -13909
rect 10820 -13961 10830 -13927
rect 10864 -13961 10874 -13927
rect 10820 -13995 10874 -13961
rect 10820 -14029 10830 -13995
rect 10864 -14029 10874 -13995
rect 10820 -14063 10874 -14029
rect 10820 -14097 10830 -14063
rect 10864 -14097 10874 -14063
rect 10820 -14109 10874 -14097
rect 10904 -13995 10958 -13909
rect 10904 -14029 10914 -13995
rect 10948 -14029 10958 -13995
rect 10904 -14063 10958 -14029
rect 10904 -14097 10914 -14063
rect 10948 -14097 10958 -14063
rect 10904 -14109 10958 -14097
rect 10988 -13927 11042 -13909
rect 10988 -13961 10998 -13927
rect 11032 -13961 11042 -13927
rect 10988 -13995 11042 -13961
rect 10988 -14029 10998 -13995
rect 11032 -14029 11042 -13995
rect 10988 -14063 11042 -14029
rect 10988 -14097 10998 -14063
rect 11032 -14097 11042 -14063
rect 10988 -14109 11042 -14097
rect 11072 -13995 11126 -13909
rect 11072 -14029 11082 -13995
rect 11116 -14029 11126 -13995
rect 11072 -14063 11126 -14029
rect 11072 -14097 11082 -14063
rect 11116 -14097 11126 -14063
rect 11072 -14109 11126 -14097
rect 11156 -13927 11210 -13909
rect 11156 -13961 11166 -13927
rect 11200 -13961 11210 -13927
rect 11156 -13995 11210 -13961
rect 11156 -14029 11166 -13995
rect 11200 -14029 11210 -13995
rect 11156 -14063 11210 -14029
rect 11156 -14097 11166 -14063
rect 11200 -14097 11210 -14063
rect 11156 -14109 11210 -14097
rect 11240 -13995 11294 -13909
rect 11240 -14029 11250 -13995
rect 11284 -14029 11294 -13995
rect 11240 -14063 11294 -14029
rect 11240 -14097 11250 -14063
rect 11284 -14097 11294 -14063
rect 11240 -14109 11294 -14097
rect 11324 -13927 11378 -13909
rect 11324 -13961 11334 -13927
rect 11368 -13961 11378 -13927
rect 11324 -13995 11378 -13961
rect 11324 -14029 11334 -13995
rect 11368 -14029 11378 -13995
rect 11324 -14063 11378 -14029
rect 11324 -14097 11334 -14063
rect 11368 -14097 11378 -14063
rect 11324 -14109 11378 -14097
rect 11408 -13995 11460 -13909
rect 11408 -14029 11418 -13995
rect 11452 -14029 11460 -13995
rect 11408 -14063 11460 -14029
rect 11408 -14097 11418 -14063
rect 11452 -14097 11460 -14063
rect 11658 -13961 11710 -13935
rect 11658 -13995 11666 -13961
rect 11700 -13995 11710 -13961
rect 11658 -14063 11710 -13995
rect 11408 -14109 11460 -14097
rect 11658 -14097 11666 -14063
rect 11700 -14097 11710 -14063
rect 11658 -14109 11710 -14097
rect 11920 -13961 11972 -13935
rect 11920 -13995 11930 -13961
rect 11964 -13995 11972 -13961
rect 11920 -14063 11972 -13995
rect 11920 -14097 11930 -14063
rect 11964 -14097 11972 -14063
rect 13590 -13961 13642 -13935
rect 13590 -13995 13598 -13961
rect 13632 -13995 13642 -13961
rect 13590 -14063 13642 -13995
rect 11920 -14109 11972 -14097
rect 13590 -14097 13598 -14063
rect 13632 -14097 13642 -14063
rect 13590 -14109 13642 -14097
rect 14588 -13961 14640 -13935
rect 14588 -13995 14598 -13961
rect 14632 -13995 14640 -13961
rect 14588 -14063 14640 -13995
rect 14588 -14097 14598 -14063
rect 14632 -14097 14640 -14063
rect 14786 -13961 14838 -13935
rect 14786 -13995 14794 -13961
rect 14828 -13995 14838 -13961
rect 14786 -14063 14838 -13995
rect 14588 -14109 14640 -14097
rect 14786 -14097 14794 -14063
rect 14828 -14097 14838 -14063
rect 14786 -14109 14838 -14097
rect 15784 -13961 15836 -13935
rect 15784 -13995 15794 -13961
rect 15828 -13995 15836 -13961
rect 15784 -14063 15836 -13995
rect 15784 -14097 15794 -14063
rect 15828 -14097 15836 -14063
rect 15982 -13961 16034 -13935
rect 15982 -13995 15990 -13961
rect 16024 -13995 16034 -13961
rect 15982 -14063 16034 -13995
rect 15784 -14109 15836 -14097
rect 15982 -14097 15990 -14063
rect 16024 -14097 16034 -14063
rect 15982 -14109 16034 -14097
rect 16612 -13961 16664 -13935
rect 16612 -13995 16622 -13961
rect 16656 -13995 16664 -13961
rect 16612 -14063 16664 -13995
rect 16612 -14097 16622 -14063
rect 16656 -14097 16664 -14063
rect 16612 -14109 16664 -14097
<< ndiffc >>
rect -2962 -478 -2928 -444
rect -2330 -478 -2296 -444
rect -1398 -471 -1364 -437
rect -1134 -471 -1100 -437
rect -934 -429 -900 -395
rect -934 -497 -900 -463
rect -766 -429 -732 -395
rect -766 -497 -732 -463
rect -570 -471 -536 -437
rect -306 -471 -272 -437
rect -16 -495 18 -461
rect 70 -484 104 -450
rect 156 -495 190 -461
rect 242 -484 276 -450
rect 328 -495 362 -461
rect 626 -471 660 -437
rect 890 -471 924 -437
rect 1169 -486 1203 -452
rect 1253 -488 1287 -454
rect 1454 -471 1488 -437
rect 1718 -471 1752 -437
rect 1914 -471 1948 -437
rect 2178 -471 2212 -437
rect 2375 -486 2409 -452
rect 2472 -486 2506 -452
rect 2632 -486 2666 -452
rect 2737 -486 2771 -452
rect 2893 -486 2927 -452
rect 2991 -486 3025 -452
rect 3202 -471 3236 -437
rect 3466 -471 3500 -437
rect 4398 -478 4432 -444
rect 5398 -478 5432 -444
rect 6422 -471 6456 -437
rect 6686 -471 6720 -437
rect 6883 -486 6917 -452
rect 6980 -486 7014 -452
rect 7140 -486 7174 -452
rect 7245 -486 7279 -452
rect 7401 -486 7435 -452
rect 7499 -486 7533 -452
rect 7710 -471 7744 -437
rect 7974 -471 8008 -437
rect 8171 -486 8205 -452
rect 8268 -486 8302 -452
rect 8428 -486 8462 -452
rect 8533 -486 8567 -452
rect 8689 -486 8723 -452
rect 8787 -486 8821 -452
rect 8998 -471 9032 -437
rect 9262 -471 9296 -437
rect 9459 -486 9493 -452
rect 9556 -486 9590 -452
rect 9716 -486 9750 -452
rect 9821 -486 9855 -452
rect 9977 -486 10011 -452
rect 10075 -486 10109 -452
rect 10286 -471 10320 -437
rect 10550 -471 10584 -437
rect 10746 -429 10780 -395
rect 10746 -497 10780 -463
rect 10830 -497 10864 -463
rect 10914 -429 10948 -395
rect 10914 -497 10948 -463
rect 10998 -497 11032 -463
rect 11082 -429 11116 -395
rect 11082 -497 11116 -463
rect 11166 -429 11200 -395
rect 11250 -497 11284 -463
rect 11334 -429 11368 -395
rect 11418 -429 11452 -395
rect 11418 -497 11452 -463
rect 11666 -471 11700 -437
rect 11930 -471 11964 -437
rect 13598 -478 13632 -444
rect 14598 -478 14632 -444
rect 14794 -478 14828 -444
rect 15794 -478 15828 -444
rect 15990 -478 16024 -444
rect 16622 -478 16656 -444
rect -2962 -668 -2928 -634
rect -2330 -668 -2296 -634
rect -1582 -668 -1548 -634
rect -950 -668 -916 -634
rect -846 -668 -812 -634
rect -214 -668 -180 -634
rect -18 -675 16 -641
rect 246 -675 280 -641
rect 457 -660 491 -626
rect 555 -660 589 -626
rect 711 -660 745 -626
rect 816 -660 850 -626
rect 976 -660 1010 -626
rect 1073 -660 1107 -626
rect 1270 -675 1304 -641
rect 1534 -675 1568 -641
rect 1730 -668 1764 -634
rect 2362 -668 2396 -634
rect 2558 -675 2592 -641
rect 2822 -675 2856 -641
rect 3033 -660 3067 -626
rect 3131 -660 3165 -626
rect 3287 -660 3321 -626
rect 3392 -660 3426 -626
rect 3552 -660 3586 -626
rect 3649 -660 3683 -626
rect 3846 -675 3880 -641
rect 4110 -675 4144 -641
rect 4306 -668 4340 -634
rect 4938 -668 4972 -634
rect 5134 -675 5168 -641
rect 5398 -675 5432 -641
rect 5609 -660 5643 -626
rect 5707 -660 5741 -626
rect 5863 -660 5897 -626
rect 5968 -660 6002 -626
rect 6128 -660 6162 -626
rect 6225 -660 6259 -626
rect 6422 -675 6456 -641
rect 6686 -675 6720 -641
rect 6882 -668 6916 -634
rect 7514 -668 7548 -634
rect 7710 -675 7744 -641
rect 7974 -675 8008 -641
rect 8185 -660 8219 -626
rect 8283 -660 8317 -626
rect 8439 -660 8473 -626
rect 8544 -660 8578 -626
rect 8704 -660 8738 -626
rect 8801 -660 8835 -626
rect 8998 -675 9032 -641
rect 9262 -675 9296 -641
rect 9458 -668 9492 -634
rect 10090 -668 10124 -634
rect 10378 -675 10412 -641
rect 10642 -675 10676 -641
rect 10761 -660 10795 -626
rect 10859 -660 10893 -626
rect 11015 -660 11049 -626
rect 11120 -660 11154 -626
rect 11280 -660 11314 -626
rect 11377 -660 11411 -626
rect 11666 -675 11700 -641
rect 11930 -675 11964 -641
rect 13690 -649 13724 -615
rect 13776 -662 13810 -628
rect 13862 -662 13896 -628
rect 13948 -662 13982 -628
rect 14034 -662 14068 -628
rect 14120 -662 14154 -628
rect 14206 -653 14240 -619
rect 14292 -662 14326 -628
rect 14378 -653 14412 -619
rect 14464 -662 14498 -628
rect 14550 -653 14584 -619
rect 14636 -662 14670 -628
rect 14722 -653 14756 -619
rect 14807 -662 14841 -628
rect 14893 -653 14927 -619
rect 14979 -662 15013 -628
rect 15065 -653 15099 -619
rect 15151 -662 15185 -628
rect 15237 -653 15271 -619
rect 15323 -662 15357 -628
rect 15409 -653 15443 -619
rect 15622 -668 15656 -634
rect 16622 -668 16656 -634
rect -2962 -1566 -2928 -1532
rect -2330 -1566 -2296 -1532
rect -1582 -1566 -1548 -1532
rect -950 -1566 -916 -1532
rect -846 -1566 -812 -1532
rect -214 -1566 -180 -1532
rect -18 -1559 16 -1525
rect 246 -1559 280 -1525
rect 443 -1574 477 -1540
rect 540 -1574 574 -1540
rect 700 -1574 734 -1540
rect 805 -1574 839 -1540
rect 961 -1574 995 -1540
rect 1059 -1574 1093 -1540
rect 1270 -1559 1304 -1525
rect 1534 -1559 1568 -1525
rect 1730 -1566 1764 -1532
rect 2362 -1566 2396 -1532
rect 2558 -1559 2592 -1525
rect 2822 -1559 2856 -1525
rect 3019 -1574 3053 -1540
rect 3116 -1574 3150 -1540
rect 3276 -1574 3310 -1540
rect 3381 -1574 3415 -1540
rect 3537 -1574 3571 -1540
rect 3635 -1574 3669 -1540
rect 3846 -1559 3880 -1525
rect 4110 -1559 4144 -1525
rect 4306 -1566 4340 -1532
rect 4938 -1566 4972 -1532
rect 5134 -1559 5168 -1525
rect 5398 -1559 5432 -1525
rect 5595 -1574 5629 -1540
rect 5692 -1574 5726 -1540
rect 5852 -1574 5886 -1540
rect 5957 -1574 5991 -1540
rect 6113 -1574 6147 -1540
rect 6211 -1574 6245 -1540
rect 6422 -1559 6456 -1525
rect 6686 -1559 6720 -1525
rect 6882 -1566 6916 -1532
rect 7514 -1566 7548 -1532
rect 7710 -1559 7744 -1525
rect 7974 -1559 8008 -1525
rect 8171 -1574 8205 -1540
rect 8268 -1574 8302 -1540
rect 8428 -1574 8462 -1540
rect 8533 -1574 8567 -1540
rect 8689 -1574 8723 -1540
rect 8787 -1574 8821 -1540
rect 8998 -1559 9032 -1525
rect 9262 -1559 9296 -1525
rect 9458 -1566 9492 -1532
rect 10090 -1566 10124 -1532
rect 10378 -1559 10412 -1525
rect 10642 -1559 10676 -1525
rect 10747 -1574 10781 -1540
rect 10844 -1574 10878 -1540
rect 11004 -1574 11038 -1540
rect 11109 -1574 11143 -1540
rect 11265 -1574 11299 -1540
rect 11363 -1574 11397 -1540
rect 11666 -1559 11700 -1525
rect 11930 -1559 11964 -1525
rect 12588 -1583 12622 -1549
rect 12674 -1572 12708 -1538
rect 12760 -1583 12794 -1549
rect 12846 -1572 12880 -1538
rect 12932 -1583 12966 -1549
rect 13230 -1559 13264 -1525
rect 13494 -1559 13528 -1525
rect 13690 -1585 13724 -1551
rect 13776 -1572 13810 -1538
rect 13862 -1572 13896 -1538
rect 13948 -1572 13982 -1538
rect 14034 -1572 14068 -1538
rect 14120 -1572 14154 -1538
rect 14206 -1581 14240 -1547
rect 14292 -1572 14326 -1538
rect 14378 -1581 14412 -1547
rect 14464 -1572 14498 -1538
rect 14550 -1581 14584 -1547
rect 14636 -1572 14670 -1538
rect 14722 -1581 14756 -1547
rect 14807 -1572 14841 -1538
rect 14893 -1581 14927 -1547
rect 14979 -1572 15013 -1538
rect 15065 -1581 15099 -1547
rect 15151 -1572 15185 -1538
rect 15237 -1581 15271 -1547
rect 15323 -1572 15357 -1538
rect 15409 -1581 15443 -1547
rect 15622 -1566 15656 -1532
rect 16622 -1566 16656 -1532
rect -2962 -1756 -2928 -1722
rect -2330 -1756 -2296 -1722
rect -1582 -1756 -1548 -1722
rect -950 -1756 -916 -1722
rect -831 -1748 -797 -1714
rect -733 -1748 -699 -1714
rect -577 -1748 -543 -1714
rect -472 -1748 -438 -1714
rect -312 -1748 -278 -1714
rect -215 -1748 -181 -1714
rect -18 -1763 16 -1729
rect 246 -1763 280 -1729
rect 457 -1748 491 -1714
rect 555 -1748 589 -1714
rect 711 -1748 745 -1714
rect 816 -1748 850 -1714
rect 976 -1748 1010 -1714
rect 1073 -1748 1107 -1714
rect 1270 -1763 1304 -1729
rect 1534 -1763 1568 -1729
rect 1730 -1756 1764 -1722
rect 2362 -1756 2396 -1722
rect 2558 -1763 2592 -1729
rect 2822 -1763 2856 -1729
rect 3033 -1748 3067 -1714
rect 3131 -1748 3165 -1714
rect 3287 -1748 3321 -1714
rect 3392 -1748 3426 -1714
rect 3552 -1748 3586 -1714
rect 3649 -1748 3683 -1714
rect 3846 -1763 3880 -1729
rect 4110 -1763 4144 -1729
rect 4306 -1756 4340 -1722
rect 4938 -1756 4972 -1722
rect 5134 -1763 5168 -1729
rect 5398 -1763 5432 -1729
rect 5609 -1748 5643 -1714
rect 5707 -1748 5741 -1714
rect 5863 -1748 5897 -1714
rect 5968 -1748 6002 -1714
rect 6128 -1748 6162 -1714
rect 6225 -1748 6259 -1714
rect 6422 -1763 6456 -1729
rect 6686 -1763 6720 -1729
rect 6882 -1756 6916 -1722
rect 7514 -1756 7548 -1722
rect 7710 -1763 7744 -1729
rect 7974 -1763 8008 -1729
rect 8185 -1748 8219 -1714
rect 8283 -1748 8317 -1714
rect 8439 -1748 8473 -1714
rect 8544 -1748 8578 -1714
rect 8704 -1748 8738 -1714
rect 8801 -1748 8835 -1714
rect 8998 -1763 9032 -1729
rect 9262 -1763 9296 -1729
rect 9458 -1756 9492 -1722
rect 10090 -1756 10124 -1722
rect 10378 -1763 10412 -1729
rect 10642 -1763 10676 -1729
rect 10761 -1748 10795 -1714
rect 10859 -1748 10893 -1714
rect 11015 -1748 11049 -1714
rect 11120 -1748 11154 -1714
rect 11280 -1748 11314 -1714
rect 11377 -1748 11411 -1714
rect 11666 -1763 11700 -1729
rect 11930 -1763 11964 -1729
rect 13690 -1737 13724 -1703
rect 13776 -1750 13810 -1716
rect 13862 -1750 13896 -1716
rect 13948 -1750 13982 -1716
rect 14034 -1750 14068 -1716
rect 14120 -1750 14154 -1716
rect 14206 -1741 14240 -1707
rect 14292 -1750 14326 -1716
rect 14378 -1741 14412 -1707
rect 14464 -1750 14498 -1716
rect 14550 -1741 14584 -1707
rect 14636 -1750 14670 -1716
rect 14722 -1741 14756 -1707
rect 14807 -1750 14841 -1716
rect 14893 -1741 14927 -1707
rect 14979 -1750 15013 -1716
rect 15065 -1741 15099 -1707
rect 15151 -1750 15185 -1716
rect 15237 -1741 15271 -1707
rect 15323 -1750 15357 -1716
rect 15409 -1741 15443 -1707
rect 15622 -1756 15656 -1722
rect 16622 -1756 16656 -1722
rect -2962 -2654 -2928 -2620
rect -2330 -2654 -2296 -2620
rect -1582 -2654 -1548 -2620
rect -950 -2654 -916 -2620
rect -846 -2654 -812 -2620
rect -214 -2654 -180 -2620
rect -18 -2647 16 -2613
rect 246 -2647 280 -2613
rect 443 -2662 477 -2628
rect 540 -2662 574 -2628
rect 700 -2662 734 -2628
rect 805 -2662 839 -2628
rect 961 -2662 995 -2628
rect 1059 -2662 1093 -2628
rect 1270 -2647 1304 -2613
rect 1534 -2647 1568 -2613
rect 1730 -2654 1764 -2620
rect 2362 -2654 2396 -2620
rect 2558 -2647 2592 -2613
rect 2822 -2647 2856 -2613
rect 3019 -2662 3053 -2628
rect 3116 -2662 3150 -2628
rect 3276 -2662 3310 -2628
rect 3381 -2662 3415 -2628
rect 3537 -2662 3571 -2628
rect 3635 -2662 3669 -2628
rect 3846 -2647 3880 -2613
rect 4110 -2647 4144 -2613
rect 4306 -2654 4340 -2620
rect 4938 -2654 4972 -2620
rect 5134 -2647 5168 -2613
rect 5398 -2647 5432 -2613
rect 5595 -2662 5629 -2628
rect 5692 -2662 5726 -2628
rect 5852 -2662 5886 -2628
rect 5957 -2662 5991 -2628
rect 6113 -2662 6147 -2628
rect 6211 -2662 6245 -2628
rect 6422 -2647 6456 -2613
rect 6686 -2647 6720 -2613
rect 6882 -2654 6916 -2620
rect 7514 -2654 7548 -2620
rect 7710 -2647 7744 -2613
rect 7974 -2647 8008 -2613
rect 8171 -2662 8205 -2628
rect 8268 -2662 8302 -2628
rect 8428 -2662 8462 -2628
rect 8533 -2662 8567 -2628
rect 8689 -2662 8723 -2628
rect 8787 -2662 8821 -2628
rect 8998 -2647 9032 -2613
rect 9262 -2647 9296 -2613
rect 9458 -2654 9492 -2620
rect 10090 -2654 10124 -2620
rect 10378 -2647 10412 -2613
rect 10642 -2647 10676 -2613
rect 10747 -2662 10781 -2628
rect 10844 -2662 10878 -2628
rect 11004 -2662 11038 -2628
rect 11109 -2662 11143 -2628
rect 11265 -2662 11299 -2628
rect 11363 -2662 11397 -2628
rect 11666 -2647 11700 -2613
rect 11930 -2647 11964 -2613
rect 12588 -2671 12622 -2637
rect 12674 -2660 12708 -2626
rect 12760 -2671 12794 -2637
rect 12846 -2660 12880 -2626
rect 12932 -2671 12966 -2637
rect 13230 -2647 13264 -2613
rect 13494 -2647 13528 -2613
rect 13690 -2673 13724 -2639
rect 13776 -2660 13810 -2626
rect 13862 -2660 13896 -2626
rect 13948 -2660 13982 -2626
rect 14034 -2660 14068 -2626
rect 14120 -2660 14154 -2626
rect 14206 -2669 14240 -2635
rect 14292 -2660 14326 -2626
rect 14378 -2669 14412 -2635
rect 14464 -2660 14498 -2626
rect 14550 -2669 14584 -2635
rect 14636 -2660 14670 -2626
rect 14722 -2669 14756 -2635
rect 14807 -2660 14841 -2626
rect 14893 -2669 14927 -2635
rect 14979 -2660 15013 -2626
rect 15065 -2669 15099 -2635
rect 15151 -2660 15185 -2626
rect 15237 -2669 15271 -2635
rect 15323 -2660 15357 -2626
rect 15409 -2669 15443 -2635
rect 15622 -2654 15656 -2620
rect 16622 -2654 16656 -2620
rect -2962 -2844 -2928 -2810
rect -2330 -2844 -2296 -2810
rect -1867 -2836 -1833 -2802
rect -1783 -2834 -1749 -2800
rect -1582 -2844 -1548 -2810
rect -950 -2844 -916 -2810
rect -846 -2844 -812 -2810
rect -214 -2844 -180 -2810
rect -18 -2851 16 -2817
rect 246 -2851 280 -2817
rect 457 -2836 491 -2802
rect 555 -2836 589 -2802
rect 711 -2836 745 -2802
rect 816 -2836 850 -2802
rect 976 -2836 1010 -2802
rect 1073 -2836 1107 -2802
rect 1270 -2851 1304 -2817
rect 1534 -2851 1568 -2817
rect 1730 -2844 1764 -2810
rect 2362 -2844 2396 -2810
rect 2558 -2851 2592 -2817
rect 2822 -2851 2856 -2817
rect 3033 -2836 3067 -2802
rect 3131 -2836 3165 -2802
rect 3287 -2836 3321 -2802
rect 3392 -2836 3426 -2802
rect 3552 -2836 3586 -2802
rect 3649 -2836 3683 -2802
rect 3846 -2851 3880 -2817
rect 4110 -2851 4144 -2817
rect 4306 -2844 4340 -2810
rect 4938 -2844 4972 -2810
rect 5134 -2851 5168 -2817
rect 5398 -2851 5432 -2817
rect 5609 -2836 5643 -2802
rect 5707 -2836 5741 -2802
rect 5863 -2836 5897 -2802
rect 5968 -2836 6002 -2802
rect 6128 -2836 6162 -2802
rect 6225 -2836 6259 -2802
rect 6422 -2851 6456 -2817
rect 6686 -2851 6720 -2817
rect 6882 -2844 6916 -2810
rect 7514 -2844 7548 -2810
rect 7710 -2851 7744 -2817
rect 7974 -2851 8008 -2817
rect 8185 -2836 8219 -2802
rect 8283 -2836 8317 -2802
rect 8439 -2836 8473 -2802
rect 8544 -2836 8578 -2802
rect 8704 -2836 8738 -2802
rect 8801 -2836 8835 -2802
rect 8998 -2851 9032 -2817
rect 9262 -2851 9296 -2817
rect 9458 -2844 9492 -2810
rect 10090 -2844 10124 -2810
rect 10378 -2851 10412 -2817
rect 10642 -2851 10676 -2817
rect 10761 -2836 10795 -2802
rect 10859 -2836 10893 -2802
rect 11015 -2836 11049 -2802
rect 11120 -2836 11154 -2802
rect 11280 -2836 11314 -2802
rect 11377 -2836 11411 -2802
rect 11666 -2851 11700 -2817
rect 11930 -2851 11964 -2817
rect 13598 -2844 13632 -2810
rect 14598 -2844 14632 -2810
rect 14794 -2844 14828 -2810
rect 15794 -2844 15828 -2810
rect 15990 -2844 16024 -2810
rect 16622 -2844 16656 -2810
rect -2962 -3742 -2928 -3708
rect -2330 -3742 -2296 -3708
rect -1582 -3742 -1548 -3708
rect -950 -3742 -916 -3708
rect -846 -3742 -812 -3708
rect -214 -3742 -180 -3708
rect -18 -3735 16 -3701
rect 246 -3735 280 -3701
rect 457 -3750 491 -3716
rect 555 -3750 589 -3716
rect 711 -3750 745 -3716
rect 816 -3750 850 -3716
rect 976 -3750 1010 -3716
rect 1073 -3750 1107 -3716
rect 1270 -3735 1304 -3701
rect 1534 -3735 1568 -3701
rect 1730 -3742 1764 -3708
rect 2362 -3742 2396 -3708
rect 2558 -3735 2592 -3701
rect 2822 -3735 2856 -3701
rect 3033 -3750 3067 -3716
rect 3131 -3750 3165 -3716
rect 3287 -3750 3321 -3716
rect 3392 -3750 3426 -3716
rect 3552 -3750 3586 -3716
rect 3649 -3750 3683 -3716
rect 3846 -3735 3880 -3701
rect 4110 -3735 4144 -3701
rect 4306 -3742 4340 -3708
rect 4938 -3742 4972 -3708
rect 5134 -3735 5168 -3701
rect 5398 -3735 5432 -3701
rect 5609 -3750 5643 -3716
rect 5707 -3750 5741 -3716
rect 5863 -3750 5897 -3716
rect 5968 -3750 6002 -3716
rect 6128 -3750 6162 -3716
rect 6225 -3750 6259 -3716
rect 6422 -3735 6456 -3701
rect 6686 -3735 6720 -3701
rect 6882 -3742 6916 -3708
rect 7514 -3742 7548 -3708
rect 7710 -3735 7744 -3701
rect 7974 -3735 8008 -3701
rect 8185 -3750 8219 -3716
rect 8283 -3750 8317 -3716
rect 8439 -3750 8473 -3716
rect 8544 -3750 8578 -3716
rect 8704 -3750 8738 -3716
rect 8801 -3750 8835 -3716
rect 8998 -3735 9032 -3701
rect 9262 -3735 9296 -3701
rect 9458 -3742 9492 -3708
rect 10090 -3742 10124 -3708
rect 10378 -3735 10412 -3701
rect 10642 -3735 10676 -3701
rect 10761 -3750 10795 -3716
rect 10859 -3750 10893 -3716
rect 11015 -3750 11049 -3716
rect 11120 -3750 11154 -3716
rect 11280 -3750 11314 -3716
rect 11377 -3750 11411 -3716
rect 11666 -3735 11700 -3701
rect 11930 -3735 11964 -3701
rect 13598 -3742 13632 -3708
rect 14598 -3742 14632 -3708
rect 14794 -3742 14828 -3708
rect 15794 -3742 15828 -3708
rect 15990 -3742 16024 -3708
rect 16622 -3742 16656 -3708
rect -2962 -3932 -2928 -3898
rect -2330 -3932 -2296 -3898
rect -1582 -3932 -1548 -3898
rect -950 -3932 -916 -3898
rect -846 -3932 -812 -3898
rect -214 -3932 -180 -3898
rect -18 -3939 16 -3905
rect 246 -3939 280 -3905
rect 443 -3924 477 -3890
rect 540 -3924 574 -3890
rect 700 -3924 734 -3890
rect 805 -3924 839 -3890
rect 961 -3924 995 -3890
rect 1059 -3924 1093 -3890
rect 1270 -3939 1304 -3905
rect 1534 -3939 1568 -3905
rect 1730 -3932 1764 -3898
rect 2362 -3932 2396 -3898
rect 2558 -3939 2592 -3905
rect 2822 -3939 2856 -3905
rect 3019 -3924 3053 -3890
rect 3116 -3924 3150 -3890
rect 3276 -3924 3310 -3890
rect 3381 -3924 3415 -3890
rect 3537 -3924 3571 -3890
rect 3635 -3924 3669 -3890
rect 3846 -3939 3880 -3905
rect 4110 -3939 4144 -3905
rect 4306 -3932 4340 -3898
rect 4938 -3932 4972 -3898
rect 5134 -3939 5168 -3905
rect 5398 -3939 5432 -3905
rect 5595 -3924 5629 -3890
rect 5692 -3924 5726 -3890
rect 5852 -3924 5886 -3890
rect 5957 -3924 5991 -3890
rect 6113 -3924 6147 -3890
rect 6211 -3924 6245 -3890
rect 6422 -3939 6456 -3905
rect 6686 -3939 6720 -3905
rect 6882 -3932 6916 -3898
rect 7514 -3932 7548 -3898
rect 7710 -3939 7744 -3905
rect 7974 -3939 8008 -3905
rect 8171 -3924 8205 -3890
rect 8268 -3924 8302 -3890
rect 8428 -3924 8462 -3890
rect 8533 -3924 8567 -3890
rect 8689 -3924 8723 -3890
rect 8787 -3924 8821 -3890
rect 8998 -3939 9032 -3905
rect 9262 -3939 9296 -3905
rect 9458 -3932 9492 -3898
rect 10090 -3932 10124 -3898
rect 10378 -3939 10412 -3905
rect 10642 -3939 10676 -3905
rect 10747 -3924 10781 -3890
rect 10844 -3924 10878 -3890
rect 11004 -3924 11038 -3890
rect 11109 -3924 11143 -3890
rect 11265 -3924 11299 -3890
rect 11363 -3924 11397 -3890
rect 11666 -3939 11700 -3905
rect 11930 -3939 11964 -3905
rect 12588 -3915 12622 -3881
rect 12674 -3926 12708 -3892
rect 12760 -3915 12794 -3881
rect 12846 -3926 12880 -3892
rect 12932 -3915 12966 -3881
rect 13230 -3939 13264 -3905
rect 13494 -3939 13528 -3905
rect 13690 -3913 13724 -3879
rect 13776 -3926 13810 -3892
rect 13862 -3926 13896 -3892
rect 13948 -3926 13982 -3892
rect 14034 -3926 14068 -3892
rect 14120 -3926 14154 -3892
rect 14206 -3917 14240 -3883
rect 14292 -3926 14326 -3892
rect 14378 -3917 14412 -3883
rect 14464 -3926 14498 -3892
rect 14550 -3917 14584 -3883
rect 14636 -3926 14670 -3892
rect 14722 -3917 14756 -3883
rect 14807 -3926 14841 -3892
rect 14893 -3917 14927 -3883
rect 14979 -3926 15013 -3892
rect 15065 -3917 15099 -3883
rect 15151 -3926 15185 -3892
rect 15237 -3917 15271 -3883
rect 15323 -3926 15357 -3892
rect 15409 -3917 15443 -3883
rect 15622 -3932 15656 -3898
rect 16622 -3932 16656 -3898
rect -2962 -4830 -2928 -4796
rect -2330 -4830 -2296 -4796
rect -1582 -4830 -1548 -4796
rect -950 -4830 -916 -4796
rect -831 -4838 -797 -4804
rect -733 -4838 -699 -4804
rect -577 -4838 -543 -4804
rect -472 -4838 -438 -4804
rect -312 -4838 -278 -4804
rect -215 -4838 -181 -4804
rect -18 -4823 16 -4789
rect 246 -4823 280 -4789
rect 457 -4838 491 -4804
rect 555 -4838 589 -4804
rect 711 -4838 745 -4804
rect 816 -4838 850 -4804
rect 976 -4838 1010 -4804
rect 1073 -4838 1107 -4804
rect 1270 -4823 1304 -4789
rect 1534 -4823 1568 -4789
rect 1730 -4830 1764 -4796
rect 2362 -4830 2396 -4796
rect 2558 -4823 2592 -4789
rect 2822 -4823 2856 -4789
rect 3033 -4838 3067 -4804
rect 3131 -4838 3165 -4804
rect 3287 -4838 3321 -4804
rect 3392 -4838 3426 -4804
rect 3552 -4838 3586 -4804
rect 3649 -4838 3683 -4804
rect 3846 -4823 3880 -4789
rect 4110 -4823 4144 -4789
rect 4306 -4830 4340 -4796
rect 4938 -4830 4972 -4796
rect 5134 -4823 5168 -4789
rect 5398 -4823 5432 -4789
rect 5609 -4838 5643 -4804
rect 5707 -4838 5741 -4804
rect 5863 -4838 5897 -4804
rect 5968 -4838 6002 -4804
rect 6128 -4838 6162 -4804
rect 6225 -4838 6259 -4804
rect 6422 -4823 6456 -4789
rect 6686 -4823 6720 -4789
rect 6882 -4830 6916 -4796
rect 7514 -4830 7548 -4796
rect 7710 -4823 7744 -4789
rect 7974 -4823 8008 -4789
rect 8185 -4838 8219 -4804
rect 8283 -4838 8317 -4804
rect 8439 -4838 8473 -4804
rect 8544 -4838 8578 -4804
rect 8704 -4838 8738 -4804
rect 8801 -4838 8835 -4804
rect 8998 -4823 9032 -4789
rect 9262 -4823 9296 -4789
rect 9458 -4830 9492 -4796
rect 10090 -4830 10124 -4796
rect 10378 -4823 10412 -4789
rect 10642 -4823 10676 -4789
rect 10761 -4838 10795 -4804
rect 10859 -4838 10893 -4804
rect 11015 -4838 11049 -4804
rect 11120 -4838 11154 -4804
rect 11280 -4838 11314 -4804
rect 11377 -4838 11411 -4804
rect 11666 -4823 11700 -4789
rect 11930 -4823 11964 -4789
rect 13690 -4849 13724 -4815
rect 13776 -4836 13810 -4802
rect 13862 -4836 13896 -4802
rect 13948 -4836 13982 -4802
rect 14034 -4836 14068 -4802
rect 14120 -4836 14154 -4802
rect 14206 -4845 14240 -4811
rect 14292 -4836 14326 -4802
rect 14378 -4845 14412 -4811
rect 14464 -4836 14498 -4802
rect 14550 -4845 14584 -4811
rect 14636 -4836 14670 -4802
rect 14722 -4845 14756 -4811
rect 14807 -4836 14841 -4802
rect 14893 -4845 14927 -4811
rect 14979 -4836 15013 -4802
rect 15065 -4845 15099 -4811
rect 15151 -4836 15185 -4802
rect 15237 -4845 15271 -4811
rect 15323 -4836 15357 -4802
rect 15409 -4845 15443 -4811
rect 15622 -4830 15656 -4796
rect 16622 -4830 16656 -4796
rect -2962 -5020 -2928 -4986
rect -2330 -5020 -2296 -4986
rect -1582 -5020 -1548 -4986
rect -950 -5020 -916 -4986
rect -846 -5020 -812 -4986
rect -214 -5020 -180 -4986
rect -18 -5027 16 -4993
rect 246 -5027 280 -4993
rect 443 -5012 477 -4978
rect 540 -5012 574 -4978
rect 700 -5012 734 -4978
rect 805 -5012 839 -4978
rect 961 -5012 995 -4978
rect 1059 -5012 1093 -4978
rect 1270 -5027 1304 -4993
rect 1534 -5027 1568 -4993
rect 1730 -5020 1764 -4986
rect 2362 -5020 2396 -4986
rect 2558 -5027 2592 -4993
rect 2822 -5027 2856 -4993
rect 3019 -5012 3053 -4978
rect 3116 -5012 3150 -4978
rect 3276 -5012 3310 -4978
rect 3381 -5012 3415 -4978
rect 3537 -5012 3571 -4978
rect 3635 -5012 3669 -4978
rect 3846 -5027 3880 -4993
rect 4110 -5027 4144 -4993
rect 4306 -5020 4340 -4986
rect 4938 -5020 4972 -4986
rect 5134 -5027 5168 -4993
rect 5398 -5027 5432 -4993
rect 5595 -5012 5629 -4978
rect 5692 -5012 5726 -4978
rect 5852 -5012 5886 -4978
rect 5957 -5012 5991 -4978
rect 6113 -5012 6147 -4978
rect 6211 -5012 6245 -4978
rect 6422 -5027 6456 -4993
rect 6686 -5027 6720 -4993
rect 6882 -5020 6916 -4986
rect 7514 -5020 7548 -4986
rect 7710 -5027 7744 -4993
rect 7974 -5027 8008 -4993
rect 8171 -5012 8205 -4978
rect 8268 -5012 8302 -4978
rect 8428 -5012 8462 -4978
rect 8533 -5012 8567 -4978
rect 8689 -5012 8723 -4978
rect 8787 -5012 8821 -4978
rect 8998 -5027 9032 -4993
rect 9262 -5027 9296 -4993
rect 9458 -5020 9492 -4986
rect 10090 -5020 10124 -4986
rect 10378 -5027 10412 -4993
rect 10642 -5027 10676 -4993
rect 10747 -5012 10781 -4978
rect 10844 -5012 10878 -4978
rect 11004 -5012 11038 -4978
rect 11109 -5012 11143 -4978
rect 11265 -5012 11299 -4978
rect 11363 -5012 11397 -4978
rect 11666 -5027 11700 -4993
rect 11930 -5027 11964 -4993
rect 12588 -5003 12622 -4969
rect 12674 -5014 12708 -4980
rect 12760 -5003 12794 -4969
rect 12846 -5014 12880 -4980
rect 12932 -5003 12966 -4969
rect 13230 -5027 13264 -4993
rect 13494 -5027 13528 -4993
rect 13690 -5001 13724 -4967
rect 13776 -5014 13810 -4980
rect 13862 -5014 13896 -4980
rect 13948 -5014 13982 -4980
rect 14034 -5014 14068 -4980
rect 14120 -5014 14154 -4980
rect 14206 -5005 14240 -4971
rect 14292 -5014 14326 -4980
rect 14378 -5005 14412 -4971
rect 14464 -5014 14498 -4980
rect 14550 -5005 14584 -4971
rect 14636 -5014 14670 -4980
rect 14722 -5005 14756 -4971
rect 14807 -5014 14841 -4980
rect 14893 -5005 14927 -4971
rect 14979 -5014 15013 -4980
rect 15065 -5005 15099 -4971
rect 15151 -5014 15185 -4980
rect 15237 -5005 15271 -4971
rect 15323 -5014 15357 -4980
rect 15409 -5005 15443 -4971
rect 15622 -5020 15656 -4986
rect 16622 -5020 16656 -4986
rect -2962 -5918 -2928 -5884
rect -2330 -5918 -2296 -5884
rect -1582 -5918 -1548 -5884
rect -950 -5918 -916 -5884
rect -846 -5918 -812 -5884
rect -214 -5918 -180 -5884
rect -18 -5911 16 -5877
rect 246 -5911 280 -5877
rect 457 -5926 491 -5892
rect 555 -5926 589 -5892
rect 711 -5926 745 -5892
rect 816 -5926 850 -5892
rect 976 -5926 1010 -5892
rect 1073 -5926 1107 -5892
rect 1270 -5911 1304 -5877
rect 1534 -5911 1568 -5877
rect 1730 -5918 1764 -5884
rect 2362 -5918 2396 -5884
rect 2558 -5911 2592 -5877
rect 2822 -5911 2856 -5877
rect 3033 -5926 3067 -5892
rect 3131 -5926 3165 -5892
rect 3287 -5926 3321 -5892
rect 3392 -5926 3426 -5892
rect 3552 -5926 3586 -5892
rect 3649 -5926 3683 -5892
rect 3846 -5911 3880 -5877
rect 4110 -5911 4144 -5877
rect 4306 -5918 4340 -5884
rect 4938 -5918 4972 -5884
rect 5134 -5911 5168 -5877
rect 5398 -5911 5432 -5877
rect 5609 -5926 5643 -5892
rect 5707 -5926 5741 -5892
rect 5863 -5926 5897 -5892
rect 5968 -5926 6002 -5892
rect 6128 -5926 6162 -5892
rect 6225 -5926 6259 -5892
rect 6422 -5911 6456 -5877
rect 6686 -5911 6720 -5877
rect 6882 -5918 6916 -5884
rect 7514 -5918 7548 -5884
rect 7710 -5911 7744 -5877
rect 7974 -5911 8008 -5877
rect 8185 -5926 8219 -5892
rect 8283 -5926 8317 -5892
rect 8439 -5926 8473 -5892
rect 8544 -5926 8578 -5892
rect 8704 -5926 8738 -5892
rect 8801 -5926 8835 -5892
rect 8998 -5911 9032 -5877
rect 9262 -5911 9296 -5877
rect 9458 -5918 9492 -5884
rect 10090 -5918 10124 -5884
rect 10378 -5911 10412 -5877
rect 10642 -5911 10676 -5877
rect 10761 -5926 10795 -5892
rect 10859 -5926 10893 -5892
rect 11015 -5926 11049 -5892
rect 11120 -5926 11154 -5892
rect 11280 -5926 11314 -5892
rect 11377 -5926 11411 -5892
rect 11666 -5911 11700 -5877
rect 11930 -5911 11964 -5877
rect 13690 -5937 13724 -5903
rect 13776 -5924 13810 -5890
rect 13862 -5924 13896 -5890
rect 13948 -5924 13982 -5890
rect 14034 -5924 14068 -5890
rect 14120 -5924 14154 -5890
rect 14206 -5933 14240 -5899
rect 14292 -5924 14326 -5890
rect 14378 -5933 14412 -5899
rect 14464 -5924 14498 -5890
rect 14550 -5933 14584 -5899
rect 14636 -5924 14670 -5890
rect 14722 -5933 14756 -5899
rect 14807 -5924 14841 -5890
rect 14893 -5933 14927 -5899
rect 14979 -5924 15013 -5890
rect 15065 -5933 15099 -5899
rect 15151 -5924 15185 -5890
rect 15237 -5933 15271 -5899
rect 15323 -5924 15357 -5890
rect 15409 -5933 15443 -5899
rect 15622 -5918 15656 -5884
rect 16622 -5918 16656 -5884
rect -2962 -6108 -2928 -6074
rect -2330 -6108 -2296 -6074
rect -1398 -6115 -1364 -6081
rect -1134 -6115 -1100 -6081
rect -934 -6089 -900 -6055
rect -934 -6157 -900 -6123
rect -766 -6089 -732 -6055
rect -766 -6157 -732 -6123
rect -570 -6115 -536 -6081
rect -306 -6115 -272 -6081
rect -16 -6091 18 -6057
rect 70 -6102 104 -6068
rect 156 -6091 190 -6057
rect 242 -6102 276 -6068
rect 328 -6091 362 -6057
rect 626 -6115 660 -6081
rect 890 -6115 924 -6081
rect 1169 -6100 1203 -6066
rect 1253 -6098 1287 -6064
rect 1454 -6115 1488 -6081
rect 1718 -6115 1752 -6081
rect 1914 -6115 1948 -6081
rect 2178 -6115 2212 -6081
rect 2375 -6100 2409 -6066
rect 2472 -6100 2506 -6066
rect 2632 -6100 2666 -6066
rect 2737 -6100 2771 -6066
rect 2893 -6100 2927 -6066
rect 2991 -6100 3025 -6066
rect 3202 -6115 3236 -6081
rect 3466 -6115 3500 -6081
rect 4398 -6108 4432 -6074
rect 5398 -6108 5432 -6074
rect 6422 -6115 6456 -6081
rect 6686 -6115 6720 -6081
rect 6883 -6100 6917 -6066
rect 6980 -6100 7014 -6066
rect 7140 -6100 7174 -6066
rect 7245 -6100 7279 -6066
rect 7401 -6100 7435 -6066
rect 7499 -6100 7533 -6066
rect 7710 -6115 7744 -6081
rect 7974 -6115 8008 -6081
rect 8171 -6100 8205 -6066
rect 8268 -6100 8302 -6066
rect 8428 -6100 8462 -6066
rect 8533 -6100 8567 -6066
rect 8689 -6100 8723 -6066
rect 8787 -6100 8821 -6066
rect 8998 -6115 9032 -6081
rect 9262 -6115 9296 -6081
rect 9459 -6100 9493 -6066
rect 9556 -6100 9590 -6066
rect 9716 -6100 9750 -6066
rect 9821 -6100 9855 -6066
rect 9977 -6100 10011 -6066
rect 10075 -6100 10109 -6066
rect 10286 -6115 10320 -6081
rect 10550 -6115 10584 -6081
rect 10746 -6089 10780 -6055
rect 10746 -6157 10780 -6123
rect 10830 -6089 10864 -6055
rect 10914 -6089 10948 -6055
rect 10914 -6157 10948 -6123
rect 10998 -6089 11032 -6055
rect 11082 -6089 11116 -6055
rect 11082 -6157 11116 -6123
rect 11166 -6157 11200 -6123
rect 11250 -6089 11284 -6055
rect 11334 -6157 11368 -6123
rect 11418 -6089 11452 -6055
rect 11418 -6157 11452 -6123
rect 11666 -6115 11700 -6081
rect 11930 -6115 11964 -6081
rect 13598 -6108 13632 -6074
rect 14598 -6108 14632 -6074
rect 14794 -6108 14828 -6074
rect 15794 -6108 15828 -6074
rect 15990 -6108 16024 -6074
rect 16622 -6108 16656 -6074
rect -2962 -7004 -2928 -6970
rect -2790 -7004 -2756 -6970
rect -2594 -6999 -2560 -6965
rect -2510 -7025 -2476 -6991
rect -2426 -6999 -2392 -6965
rect -2322 -7025 -2288 -6991
rect -2237 -7011 -2203 -6977
rect -2126 -7011 -2092 -6977
rect -1927 -7017 -1893 -6983
rect -1808 -7011 -1774 -6977
rect -1705 -7011 -1671 -6977
rect -1507 -7011 -1473 -6977
rect -1401 -6956 -1367 -6922
rect -1401 -7024 -1367 -6990
rect -1317 -6995 -1283 -6961
rect -1233 -6954 -1199 -6920
rect -1233 -7022 -1199 -6988
rect -1129 -6999 -1095 -6965
rect -1034 -7025 -1000 -6991
rect -950 -6987 -916 -6953
rect -846 -7006 -812 -6972
rect -214 -7006 -180 -6972
rect -18 -7006 16 -6972
rect 614 -7006 648 -6972
rect 718 -7006 752 -6972
rect 1350 -7006 1384 -6972
rect 1546 -7006 1580 -6972
rect 2178 -7006 2212 -6972
rect 2282 -7006 2316 -6972
rect 2914 -7006 2948 -6972
rect 3110 -7006 3144 -6972
rect 3742 -7006 3776 -6972
rect 3846 -7006 3880 -6972
rect 4478 -7006 4512 -6972
rect 4674 -7006 4708 -6972
rect 5306 -7006 5340 -6972
rect 5410 -7006 5444 -6972
rect 6042 -7006 6076 -6972
rect 6238 -7006 6272 -6972
rect 6870 -7006 6904 -6972
rect 6974 -7006 7008 -6972
rect 7606 -7006 7640 -6972
rect 7802 -7006 7836 -6972
rect 8434 -7006 8468 -6972
rect 8538 -7006 8572 -6972
rect 9170 -7006 9204 -6972
rect 15990 -7006 16024 -6972
rect 16622 -7006 16656 -6972
rect -2962 -7196 -2928 -7162
rect -2330 -7196 -2296 -7162
rect -1582 -7196 -1548 -7162
rect -950 -7196 -916 -7162
rect -846 -7196 -812 -7162
rect -214 -7196 -180 -7162
rect -18 -7196 16 -7162
rect 614 -7196 648 -7162
rect 718 -7196 752 -7162
rect 1350 -7196 1384 -7162
rect 1546 -7196 1580 -7162
rect 2178 -7196 2212 -7162
rect 2282 -7203 2316 -7169
rect 2546 -7203 2580 -7169
rect 2931 -7186 2965 -7152
rect 3015 -7188 3049 -7154
rect 3294 -7203 3328 -7169
rect 3558 -7203 3592 -7169
rect 3758 -7177 3792 -7143
rect 3758 -7245 3792 -7211
rect 3926 -7177 3960 -7143
rect 3926 -7245 3960 -7211
rect 4122 -7203 4156 -7169
rect 4386 -7203 4420 -7169
rect 4582 -7196 4616 -7162
rect 4666 -7177 4700 -7143
rect 4873 -7192 4907 -7158
rect 5108 -7192 5142 -7158
rect 5176 -7192 5210 -7158
rect 5260 -7192 5294 -7158
rect 5502 -7203 5536 -7169
rect 5766 -7203 5800 -7169
rect 5962 -7215 5996 -7181
rect 6046 -7177 6080 -7143
rect 6141 -7203 6175 -7169
rect 6245 -7180 6279 -7146
rect 6245 -7248 6279 -7214
rect 6329 -7207 6363 -7173
rect 6413 -7178 6447 -7144
rect 6413 -7246 6447 -7212
rect 6519 -7191 6553 -7157
rect 6717 -7191 6751 -7157
rect 6820 -7191 6854 -7157
rect 6939 -7185 6973 -7151
rect 7138 -7191 7172 -7157
rect 7249 -7191 7283 -7157
rect 7334 -7177 7368 -7143
rect 7438 -7203 7472 -7169
rect 7522 -7177 7556 -7143
rect 7606 -7203 7640 -7169
rect 7802 -7196 7836 -7162
rect 8434 -7196 8468 -7162
rect 8538 -7196 8572 -7162
rect 9170 -7196 9204 -7162
rect 15990 -7196 16024 -7162
rect 16622 -7196 16656 -7162
rect -2962 -8094 -2928 -8060
rect -2330 -8094 -2296 -8060
rect -1398 -8087 -1364 -8053
rect -1134 -8087 -1100 -8053
rect -934 -8045 -900 -8011
rect -934 -8113 -900 -8079
rect -766 -8045 -732 -8011
rect -766 -8113 -732 -8079
rect -570 -8087 -536 -8053
rect -306 -8087 -272 -8053
rect -16 -8111 18 -8077
rect 70 -8100 104 -8066
rect 156 -8111 190 -8077
rect 242 -8100 276 -8066
rect 328 -8111 362 -8077
rect 626 -8087 660 -8053
rect 890 -8087 924 -8053
rect 1169 -8102 1203 -8068
rect 1253 -8104 1287 -8070
rect 1454 -8087 1488 -8053
rect 1718 -8087 1752 -8053
rect 1914 -8087 1948 -8053
rect 2178 -8087 2212 -8053
rect 2375 -8102 2409 -8068
rect 2472 -8102 2506 -8068
rect 2632 -8102 2666 -8068
rect 2737 -8102 2771 -8068
rect 2893 -8102 2927 -8068
rect 2991 -8102 3025 -8068
rect 3202 -8087 3236 -8053
rect 3466 -8087 3500 -8053
rect 4398 -8094 4432 -8060
rect 5398 -8094 5432 -8060
rect 6422 -8087 6456 -8053
rect 6686 -8087 6720 -8053
rect 6883 -8102 6917 -8068
rect 6980 -8102 7014 -8068
rect 7140 -8102 7174 -8068
rect 7245 -8102 7279 -8068
rect 7401 -8102 7435 -8068
rect 7499 -8102 7533 -8068
rect 7710 -8087 7744 -8053
rect 7974 -8087 8008 -8053
rect 8171 -8102 8205 -8068
rect 8268 -8102 8302 -8068
rect 8428 -8102 8462 -8068
rect 8533 -8102 8567 -8068
rect 8689 -8102 8723 -8068
rect 8787 -8102 8821 -8068
rect 8998 -8087 9032 -8053
rect 9262 -8087 9296 -8053
rect 9459 -8102 9493 -8068
rect 9556 -8102 9590 -8068
rect 9716 -8102 9750 -8068
rect 9821 -8102 9855 -8068
rect 9977 -8102 10011 -8068
rect 10075 -8102 10109 -8068
rect 10286 -8087 10320 -8053
rect 10550 -8087 10584 -8053
rect 10746 -8045 10780 -8011
rect 10746 -8113 10780 -8079
rect 10830 -8113 10864 -8079
rect 10914 -8045 10948 -8011
rect 10914 -8113 10948 -8079
rect 10998 -8113 11032 -8079
rect 11082 -8045 11116 -8011
rect 11082 -8113 11116 -8079
rect 11166 -8045 11200 -8011
rect 11250 -8113 11284 -8079
rect 11334 -8045 11368 -8011
rect 11418 -8045 11452 -8011
rect 11418 -8113 11452 -8079
rect 11666 -8087 11700 -8053
rect 11930 -8087 11964 -8053
rect 13598 -8094 13632 -8060
rect 14598 -8094 14632 -8060
rect 14794 -8094 14828 -8060
rect 15794 -8094 15828 -8060
rect 15990 -8094 16024 -8060
rect 16622 -8094 16656 -8060
rect -2962 -8284 -2928 -8250
rect -2330 -8284 -2296 -8250
rect -1582 -8284 -1548 -8250
rect -950 -8284 -916 -8250
rect -846 -8284 -812 -8250
rect -214 -8284 -180 -8250
rect -18 -8291 16 -8257
rect 246 -8291 280 -8257
rect 457 -8276 491 -8242
rect 555 -8276 589 -8242
rect 711 -8276 745 -8242
rect 816 -8276 850 -8242
rect 976 -8276 1010 -8242
rect 1073 -8276 1107 -8242
rect 1270 -8291 1304 -8257
rect 1534 -8291 1568 -8257
rect 1730 -8284 1764 -8250
rect 2362 -8284 2396 -8250
rect 2558 -8291 2592 -8257
rect 2822 -8291 2856 -8257
rect 3033 -8276 3067 -8242
rect 3131 -8276 3165 -8242
rect 3287 -8276 3321 -8242
rect 3392 -8276 3426 -8242
rect 3552 -8276 3586 -8242
rect 3649 -8276 3683 -8242
rect 3846 -8291 3880 -8257
rect 4110 -8291 4144 -8257
rect 4306 -8284 4340 -8250
rect 4938 -8284 4972 -8250
rect 5134 -8291 5168 -8257
rect 5398 -8291 5432 -8257
rect 5609 -8276 5643 -8242
rect 5707 -8276 5741 -8242
rect 5863 -8276 5897 -8242
rect 5968 -8276 6002 -8242
rect 6128 -8276 6162 -8242
rect 6225 -8276 6259 -8242
rect 6422 -8291 6456 -8257
rect 6686 -8291 6720 -8257
rect 6882 -8284 6916 -8250
rect 7514 -8284 7548 -8250
rect 7710 -8291 7744 -8257
rect 7974 -8291 8008 -8257
rect 8185 -8276 8219 -8242
rect 8283 -8276 8317 -8242
rect 8439 -8276 8473 -8242
rect 8544 -8276 8578 -8242
rect 8704 -8276 8738 -8242
rect 8801 -8276 8835 -8242
rect 8998 -8291 9032 -8257
rect 9262 -8291 9296 -8257
rect 9458 -8284 9492 -8250
rect 10090 -8284 10124 -8250
rect 10378 -8291 10412 -8257
rect 10642 -8291 10676 -8257
rect 10761 -8276 10795 -8242
rect 10859 -8276 10893 -8242
rect 11015 -8276 11049 -8242
rect 11120 -8276 11154 -8242
rect 11280 -8276 11314 -8242
rect 11377 -8276 11411 -8242
rect 11666 -8291 11700 -8257
rect 11930 -8291 11964 -8257
rect 13690 -8265 13724 -8231
rect 13776 -8278 13810 -8244
rect 13862 -8278 13896 -8244
rect 13948 -8278 13982 -8244
rect 14034 -8278 14068 -8244
rect 14120 -8278 14154 -8244
rect 14206 -8269 14240 -8235
rect 14292 -8278 14326 -8244
rect 14378 -8269 14412 -8235
rect 14464 -8278 14498 -8244
rect 14550 -8269 14584 -8235
rect 14636 -8278 14670 -8244
rect 14722 -8269 14756 -8235
rect 14807 -8278 14841 -8244
rect 14893 -8269 14927 -8235
rect 14979 -8278 15013 -8244
rect 15065 -8269 15099 -8235
rect 15151 -8278 15185 -8244
rect 15237 -8269 15271 -8235
rect 15323 -8278 15357 -8244
rect 15409 -8269 15443 -8235
rect 15622 -8284 15656 -8250
rect 16622 -8284 16656 -8250
rect -2962 -9182 -2928 -9148
rect -2330 -9182 -2296 -9148
rect -1582 -9182 -1548 -9148
rect -950 -9182 -916 -9148
rect -846 -9182 -812 -9148
rect -214 -9182 -180 -9148
rect -18 -9175 16 -9141
rect 246 -9175 280 -9141
rect 443 -9190 477 -9156
rect 540 -9190 574 -9156
rect 700 -9190 734 -9156
rect 805 -9190 839 -9156
rect 961 -9190 995 -9156
rect 1059 -9190 1093 -9156
rect 1270 -9175 1304 -9141
rect 1534 -9175 1568 -9141
rect 1730 -9182 1764 -9148
rect 2362 -9182 2396 -9148
rect 2558 -9175 2592 -9141
rect 2822 -9175 2856 -9141
rect 3019 -9190 3053 -9156
rect 3116 -9190 3150 -9156
rect 3276 -9190 3310 -9156
rect 3381 -9190 3415 -9156
rect 3537 -9190 3571 -9156
rect 3635 -9190 3669 -9156
rect 3846 -9175 3880 -9141
rect 4110 -9175 4144 -9141
rect 4306 -9182 4340 -9148
rect 4938 -9182 4972 -9148
rect 5134 -9175 5168 -9141
rect 5398 -9175 5432 -9141
rect 5595 -9190 5629 -9156
rect 5692 -9190 5726 -9156
rect 5852 -9190 5886 -9156
rect 5957 -9190 5991 -9156
rect 6113 -9190 6147 -9156
rect 6211 -9190 6245 -9156
rect 6422 -9175 6456 -9141
rect 6686 -9175 6720 -9141
rect 6882 -9182 6916 -9148
rect 7514 -9182 7548 -9148
rect 7710 -9175 7744 -9141
rect 7974 -9175 8008 -9141
rect 8171 -9190 8205 -9156
rect 8268 -9190 8302 -9156
rect 8428 -9190 8462 -9156
rect 8533 -9190 8567 -9156
rect 8689 -9190 8723 -9156
rect 8787 -9190 8821 -9156
rect 8998 -9175 9032 -9141
rect 9262 -9175 9296 -9141
rect 9458 -9182 9492 -9148
rect 10090 -9182 10124 -9148
rect 10378 -9175 10412 -9141
rect 10642 -9175 10676 -9141
rect 10747 -9190 10781 -9156
rect 10844 -9190 10878 -9156
rect 11004 -9190 11038 -9156
rect 11109 -9190 11143 -9156
rect 11265 -9190 11299 -9156
rect 11363 -9190 11397 -9156
rect 11666 -9175 11700 -9141
rect 11930 -9175 11964 -9141
rect 12588 -9199 12622 -9165
rect 12674 -9188 12708 -9154
rect 12760 -9199 12794 -9165
rect 12846 -9188 12880 -9154
rect 12932 -9199 12966 -9165
rect 13230 -9175 13264 -9141
rect 13494 -9175 13528 -9141
rect 13690 -9201 13724 -9167
rect 13776 -9188 13810 -9154
rect 13862 -9188 13896 -9154
rect 13948 -9188 13982 -9154
rect 14034 -9188 14068 -9154
rect 14120 -9188 14154 -9154
rect 14206 -9197 14240 -9163
rect 14292 -9188 14326 -9154
rect 14378 -9197 14412 -9163
rect 14464 -9188 14498 -9154
rect 14550 -9197 14584 -9163
rect 14636 -9188 14670 -9154
rect 14722 -9197 14756 -9163
rect 14807 -9188 14841 -9154
rect 14893 -9197 14927 -9163
rect 14979 -9188 15013 -9154
rect 15065 -9197 15099 -9163
rect 15151 -9188 15185 -9154
rect 15237 -9197 15271 -9163
rect 15323 -9188 15357 -9154
rect 15409 -9197 15443 -9163
rect 15622 -9182 15656 -9148
rect 16622 -9182 16656 -9148
rect -2962 -9372 -2928 -9338
rect -2330 -9372 -2296 -9338
rect -1582 -9372 -1548 -9338
rect -950 -9372 -916 -9338
rect -831 -9364 -797 -9330
rect -733 -9364 -699 -9330
rect -577 -9364 -543 -9330
rect -472 -9364 -438 -9330
rect -312 -9364 -278 -9330
rect -215 -9364 -181 -9330
rect -18 -9379 16 -9345
rect 246 -9379 280 -9345
rect 457 -9364 491 -9330
rect 555 -9364 589 -9330
rect 711 -9364 745 -9330
rect 816 -9364 850 -9330
rect 976 -9364 1010 -9330
rect 1073 -9364 1107 -9330
rect 1270 -9379 1304 -9345
rect 1534 -9379 1568 -9345
rect 1730 -9372 1764 -9338
rect 2362 -9372 2396 -9338
rect 2558 -9379 2592 -9345
rect 2822 -9379 2856 -9345
rect 3033 -9364 3067 -9330
rect 3131 -9364 3165 -9330
rect 3287 -9364 3321 -9330
rect 3392 -9364 3426 -9330
rect 3552 -9364 3586 -9330
rect 3649 -9364 3683 -9330
rect 3846 -9379 3880 -9345
rect 4110 -9379 4144 -9345
rect 4306 -9372 4340 -9338
rect 4938 -9372 4972 -9338
rect 5134 -9379 5168 -9345
rect 5398 -9379 5432 -9345
rect 5609 -9364 5643 -9330
rect 5707 -9364 5741 -9330
rect 5863 -9364 5897 -9330
rect 5968 -9364 6002 -9330
rect 6128 -9364 6162 -9330
rect 6225 -9364 6259 -9330
rect 6422 -9379 6456 -9345
rect 6686 -9379 6720 -9345
rect 6882 -9372 6916 -9338
rect 7514 -9372 7548 -9338
rect 7710 -9379 7744 -9345
rect 7974 -9379 8008 -9345
rect 8185 -9364 8219 -9330
rect 8283 -9364 8317 -9330
rect 8439 -9364 8473 -9330
rect 8544 -9364 8578 -9330
rect 8704 -9364 8738 -9330
rect 8801 -9364 8835 -9330
rect 8998 -9379 9032 -9345
rect 9262 -9379 9296 -9345
rect 9458 -9372 9492 -9338
rect 10090 -9372 10124 -9338
rect 10378 -9379 10412 -9345
rect 10642 -9379 10676 -9345
rect 10761 -9364 10795 -9330
rect 10859 -9364 10893 -9330
rect 11015 -9364 11049 -9330
rect 11120 -9364 11154 -9330
rect 11280 -9364 11314 -9330
rect 11377 -9364 11411 -9330
rect 11666 -9379 11700 -9345
rect 11930 -9379 11964 -9345
rect 13690 -9353 13724 -9319
rect 13776 -9366 13810 -9332
rect 13862 -9366 13896 -9332
rect 13948 -9366 13982 -9332
rect 14034 -9366 14068 -9332
rect 14120 -9366 14154 -9332
rect 14206 -9357 14240 -9323
rect 14292 -9366 14326 -9332
rect 14378 -9357 14412 -9323
rect 14464 -9366 14498 -9332
rect 14550 -9357 14584 -9323
rect 14636 -9366 14670 -9332
rect 14722 -9357 14756 -9323
rect 14807 -9366 14841 -9332
rect 14893 -9357 14927 -9323
rect 14979 -9366 15013 -9332
rect 15065 -9357 15099 -9323
rect 15151 -9366 15185 -9332
rect 15237 -9357 15271 -9323
rect 15323 -9366 15357 -9332
rect 15409 -9357 15443 -9323
rect 15622 -9372 15656 -9338
rect 16622 -9372 16656 -9338
rect -2962 -10270 -2928 -10236
rect -2330 -10270 -2296 -10236
rect -1582 -10270 -1548 -10236
rect -950 -10270 -916 -10236
rect -846 -10270 -812 -10236
rect -214 -10270 -180 -10236
rect -18 -10263 16 -10229
rect 246 -10263 280 -10229
rect 443 -10278 477 -10244
rect 540 -10278 574 -10244
rect 700 -10278 734 -10244
rect 805 -10278 839 -10244
rect 961 -10278 995 -10244
rect 1059 -10278 1093 -10244
rect 1270 -10263 1304 -10229
rect 1534 -10263 1568 -10229
rect 1730 -10270 1764 -10236
rect 2362 -10270 2396 -10236
rect 2558 -10263 2592 -10229
rect 2822 -10263 2856 -10229
rect 3019 -10278 3053 -10244
rect 3116 -10278 3150 -10244
rect 3276 -10278 3310 -10244
rect 3381 -10278 3415 -10244
rect 3537 -10278 3571 -10244
rect 3635 -10278 3669 -10244
rect 3846 -10263 3880 -10229
rect 4110 -10263 4144 -10229
rect 4306 -10270 4340 -10236
rect 4938 -10270 4972 -10236
rect 5134 -10263 5168 -10229
rect 5398 -10263 5432 -10229
rect 5595 -10278 5629 -10244
rect 5692 -10278 5726 -10244
rect 5852 -10278 5886 -10244
rect 5957 -10278 5991 -10244
rect 6113 -10278 6147 -10244
rect 6211 -10278 6245 -10244
rect 6422 -10263 6456 -10229
rect 6686 -10263 6720 -10229
rect 6882 -10270 6916 -10236
rect 7514 -10270 7548 -10236
rect 7710 -10263 7744 -10229
rect 7974 -10263 8008 -10229
rect 8171 -10278 8205 -10244
rect 8268 -10278 8302 -10244
rect 8428 -10278 8462 -10244
rect 8533 -10278 8567 -10244
rect 8689 -10278 8723 -10244
rect 8787 -10278 8821 -10244
rect 8998 -10263 9032 -10229
rect 9262 -10263 9296 -10229
rect 9458 -10270 9492 -10236
rect 10090 -10270 10124 -10236
rect 10378 -10263 10412 -10229
rect 10642 -10263 10676 -10229
rect 10747 -10278 10781 -10244
rect 10844 -10278 10878 -10244
rect 11004 -10278 11038 -10244
rect 11109 -10278 11143 -10244
rect 11265 -10278 11299 -10244
rect 11363 -10278 11397 -10244
rect 11666 -10263 11700 -10229
rect 11930 -10263 11964 -10229
rect 12588 -10287 12622 -10253
rect 12674 -10276 12708 -10242
rect 12760 -10287 12794 -10253
rect 12846 -10276 12880 -10242
rect 12932 -10287 12966 -10253
rect 13230 -10263 13264 -10229
rect 13494 -10263 13528 -10229
rect 13690 -10289 13724 -10255
rect 13776 -10276 13810 -10242
rect 13862 -10276 13896 -10242
rect 13948 -10276 13982 -10242
rect 14034 -10276 14068 -10242
rect 14120 -10276 14154 -10242
rect 14206 -10285 14240 -10251
rect 14292 -10276 14326 -10242
rect 14378 -10285 14412 -10251
rect 14464 -10276 14498 -10242
rect 14550 -10285 14584 -10251
rect 14636 -10276 14670 -10242
rect 14722 -10285 14756 -10251
rect 14807 -10276 14841 -10242
rect 14893 -10285 14927 -10251
rect 14979 -10276 15013 -10242
rect 15065 -10285 15099 -10251
rect 15151 -10276 15185 -10242
rect 15237 -10285 15271 -10251
rect 15323 -10276 15357 -10242
rect 15409 -10285 15443 -10251
rect 15622 -10270 15656 -10236
rect 16622 -10270 16656 -10236
rect -2962 -10460 -2928 -10426
rect -2330 -10460 -2296 -10426
rect -1867 -10452 -1833 -10418
rect -1783 -10450 -1749 -10416
rect -1582 -10460 -1548 -10426
rect -950 -10460 -916 -10426
rect -846 -10460 -812 -10426
rect -214 -10460 -180 -10426
rect -18 -10467 16 -10433
rect 246 -10467 280 -10433
rect 457 -10452 491 -10418
rect 555 -10452 589 -10418
rect 711 -10452 745 -10418
rect 816 -10452 850 -10418
rect 976 -10452 1010 -10418
rect 1073 -10452 1107 -10418
rect 1270 -10467 1304 -10433
rect 1534 -10467 1568 -10433
rect 1730 -10460 1764 -10426
rect 2362 -10460 2396 -10426
rect 2558 -10467 2592 -10433
rect 2822 -10467 2856 -10433
rect 3033 -10452 3067 -10418
rect 3131 -10452 3165 -10418
rect 3287 -10452 3321 -10418
rect 3392 -10452 3426 -10418
rect 3552 -10452 3586 -10418
rect 3649 -10452 3683 -10418
rect 3846 -10467 3880 -10433
rect 4110 -10467 4144 -10433
rect 4306 -10460 4340 -10426
rect 4938 -10460 4972 -10426
rect 5134 -10467 5168 -10433
rect 5398 -10467 5432 -10433
rect 5609 -10452 5643 -10418
rect 5707 -10452 5741 -10418
rect 5863 -10452 5897 -10418
rect 5968 -10452 6002 -10418
rect 6128 -10452 6162 -10418
rect 6225 -10452 6259 -10418
rect 6422 -10467 6456 -10433
rect 6686 -10467 6720 -10433
rect 6882 -10460 6916 -10426
rect 7514 -10460 7548 -10426
rect 7710 -10467 7744 -10433
rect 7974 -10467 8008 -10433
rect 8185 -10452 8219 -10418
rect 8283 -10452 8317 -10418
rect 8439 -10452 8473 -10418
rect 8544 -10452 8578 -10418
rect 8704 -10452 8738 -10418
rect 8801 -10452 8835 -10418
rect 8998 -10467 9032 -10433
rect 9262 -10467 9296 -10433
rect 9458 -10460 9492 -10426
rect 10090 -10460 10124 -10426
rect 10378 -10467 10412 -10433
rect 10642 -10467 10676 -10433
rect 10761 -10452 10795 -10418
rect 10859 -10452 10893 -10418
rect 11015 -10452 11049 -10418
rect 11120 -10452 11154 -10418
rect 11280 -10452 11314 -10418
rect 11377 -10452 11411 -10418
rect 11666 -10467 11700 -10433
rect 11930 -10467 11964 -10433
rect 13598 -10460 13632 -10426
rect 14598 -10460 14632 -10426
rect 14794 -10460 14828 -10426
rect 15794 -10460 15828 -10426
rect 15990 -10460 16024 -10426
rect 16622 -10460 16656 -10426
rect -2962 -11358 -2928 -11324
rect -2330 -11358 -2296 -11324
rect -1582 -11358 -1548 -11324
rect -950 -11358 -916 -11324
rect -846 -11358 -812 -11324
rect -214 -11358 -180 -11324
rect -18 -11351 16 -11317
rect 246 -11351 280 -11317
rect 457 -11366 491 -11332
rect 555 -11366 589 -11332
rect 711 -11366 745 -11332
rect 816 -11366 850 -11332
rect 976 -11366 1010 -11332
rect 1073 -11366 1107 -11332
rect 1270 -11351 1304 -11317
rect 1534 -11351 1568 -11317
rect 1730 -11358 1764 -11324
rect 2362 -11358 2396 -11324
rect 2558 -11351 2592 -11317
rect 2822 -11351 2856 -11317
rect 3033 -11366 3067 -11332
rect 3131 -11366 3165 -11332
rect 3287 -11366 3321 -11332
rect 3392 -11366 3426 -11332
rect 3552 -11366 3586 -11332
rect 3649 -11366 3683 -11332
rect 3846 -11351 3880 -11317
rect 4110 -11351 4144 -11317
rect 4306 -11358 4340 -11324
rect 4938 -11358 4972 -11324
rect 5134 -11351 5168 -11317
rect 5398 -11351 5432 -11317
rect 5609 -11366 5643 -11332
rect 5707 -11366 5741 -11332
rect 5863 -11366 5897 -11332
rect 5968 -11366 6002 -11332
rect 6128 -11366 6162 -11332
rect 6225 -11366 6259 -11332
rect 6422 -11351 6456 -11317
rect 6686 -11351 6720 -11317
rect 6882 -11358 6916 -11324
rect 7514 -11358 7548 -11324
rect 7710 -11351 7744 -11317
rect 7974 -11351 8008 -11317
rect 8185 -11366 8219 -11332
rect 8283 -11366 8317 -11332
rect 8439 -11366 8473 -11332
rect 8544 -11366 8578 -11332
rect 8704 -11366 8738 -11332
rect 8801 -11366 8835 -11332
rect 8998 -11351 9032 -11317
rect 9262 -11351 9296 -11317
rect 9458 -11358 9492 -11324
rect 10090 -11358 10124 -11324
rect 10378 -11351 10412 -11317
rect 10642 -11351 10676 -11317
rect 10761 -11366 10795 -11332
rect 10859 -11366 10893 -11332
rect 11015 -11366 11049 -11332
rect 11120 -11366 11154 -11332
rect 11280 -11366 11314 -11332
rect 11377 -11366 11411 -11332
rect 11666 -11351 11700 -11317
rect 11930 -11351 11964 -11317
rect 13598 -11358 13632 -11324
rect 14598 -11358 14632 -11324
rect 14794 -11358 14828 -11324
rect 15794 -11358 15828 -11324
rect 15990 -11358 16024 -11324
rect 16622 -11358 16656 -11324
rect -2962 -11548 -2928 -11514
rect -2330 -11548 -2296 -11514
rect -1582 -11548 -1548 -11514
rect -950 -11548 -916 -11514
rect -846 -11548 -812 -11514
rect -214 -11548 -180 -11514
rect -18 -11555 16 -11521
rect 246 -11555 280 -11521
rect 443 -11540 477 -11506
rect 540 -11540 574 -11506
rect 700 -11540 734 -11506
rect 805 -11540 839 -11506
rect 961 -11540 995 -11506
rect 1059 -11540 1093 -11506
rect 1270 -11555 1304 -11521
rect 1534 -11555 1568 -11521
rect 1730 -11548 1764 -11514
rect 2362 -11548 2396 -11514
rect 2558 -11555 2592 -11521
rect 2822 -11555 2856 -11521
rect 3019 -11540 3053 -11506
rect 3116 -11540 3150 -11506
rect 3276 -11540 3310 -11506
rect 3381 -11540 3415 -11506
rect 3537 -11540 3571 -11506
rect 3635 -11540 3669 -11506
rect 3846 -11555 3880 -11521
rect 4110 -11555 4144 -11521
rect 4306 -11548 4340 -11514
rect 4938 -11548 4972 -11514
rect 5134 -11555 5168 -11521
rect 5398 -11555 5432 -11521
rect 5595 -11540 5629 -11506
rect 5692 -11540 5726 -11506
rect 5852 -11540 5886 -11506
rect 5957 -11540 5991 -11506
rect 6113 -11540 6147 -11506
rect 6211 -11540 6245 -11506
rect 6422 -11555 6456 -11521
rect 6686 -11555 6720 -11521
rect 6882 -11548 6916 -11514
rect 7514 -11548 7548 -11514
rect 7710 -11555 7744 -11521
rect 7974 -11555 8008 -11521
rect 8171 -11540 8205 -11506
rect 8268 -11540 8302 -11506
rect 8428 -11540 8462 -11506
rect 8533 -11540 8567 -11506
rect 8689 -11540 8723 -11506
rect 8787 -11540 8821 -11506
rect 8998 -11555 9032 -11521
rect 9262 -11555 9296 -11521
rect 9458 -11548 9492 -11514
rect 10090 -11548 10124 -11514
rect 10378 -11555 10412 -11521
rect 10642 -11555 10676 -11521
rect 10747 -11540 10781 -11506
rect 10844 -11540 10878 -11506
rect 11004 -11540 11038 -11506
rect 11109 -11540 11143 -11506
rect 11265 -11540 11299 -11506
rect 11363 -11540 11397 -11506
rect 11666 -11555 11700 -11521
rect 11930 -11555 11964 -11521
rect 12588 -11531 12622 -11497
rect 12674 -11542 12708 -11508
rect 12760 -11531 12794 -11497
rect 12846 -11542 12880 -11508
rect 12932 -11531 12966 -11497
rect 13230 -11555 13264 -11521
rect 13494 -11555 13528 -11521
rect 13690 -11529 13724 -11495
rect 13776 -11542 13810 -11508
rect 13862 -11542 13896 -11508
rect 13948 -11542 13982 -11508
rect 14034 -11542 14068 -11508
rect 14120 -11542 14154 -11508
rect 14206 -11533 14240 -11499
rect 14292 -11542 14326 -11508
rect 14378 -11533 14412 -11499
rect 14464 -11542 14498 -11508
rect 14550 -11533 14584 -11499
rect 14636 -11542 14670 -11508
rect 14722 -11533 14756 -11499
rect 14807 -11542 14841 -11508
rect 14893 -11533 14927 -11499
rect 14979 -11542 15013 -11508
rect 15065 -11533 15099 -11499
rect 15151 -11542 15185 -11508
rect 15237 -11533 15271 -11499
rect 15323 -11542 15357 -11508
rect 15409 -11533 15443 -11499
rect 15622 -11548 15656 -11514
rect 16622 -11548 16656 -11514
rect -2962 -12446 -2928 -12412
rect -2330 -12446 -2296 -12412
rect -1582 -12446 -1548 -12412
rect -950 -12446 -916 -12412
rect -831 -12454 -797 -12420
rect -733 -12454 -699 -12420
rect -577 -12454 -543 -12420
rect -472 -12454 -438 -12420
rect -312 -12454 -278 -12420
rect -215 -12454 -181 -12420
rect -18 -12439 16 -12405
rect 246 -12439 280 -12405
rect 457 -12454 491 -12420
rect 555 -12454 589 -12420
rect 711 -12454 745 -12420
rect 816 -12454 850 -12420
rect 976 -12454 1010 -12420
rect 1073 -12454 1107 -12420
rect 1270 -12439 1304 -12405
rect 1534 -12439 1568 -12405
rect 1730 -12446 1764 -12412
rect 2362 -12446 2396 -12412
rect 2558 -12439 2592 -12405
rect 2822 -12439 2856 -12405
rect 3033 -12454 3067 -12420
rect 3131 -12454 3165 -12420
rect 3287 -12454 3321 -12420
rect 3392 -12454 3426 -12420
rect 3552 -12454 3586 -12420
rect 3649 -12454 3683 -12420
rect 3846 -12439 3880 -12405
rect 4110 -12439 4144 -12405
rect 4306 -12446 4340 -12412
rect 4938 -12446 4972 -12412
rect 5134 -12439 5168 -12405
rect 5398 -12439 5432 -12405
rect 5609 -12454 5643 -12420
rect 5707 -12454 5741 -12420
rect 5863 -12454 5897 -12420
rect 5968 -12454 6002 -12420
rect 6128 -12454 6162 -12420
rect 6225 -12454 6259 -12420
rect 6422 -12439 6456 -12405
rect 6686 -12439 6720 -12405
rect 6882 -12446 6916 -12412
rect 7514 -12446 7548 -12412
rect 7710 -12439 7744 -12405
rect 7974 -12439 8008 -12405
rect 8185 -12454 8219 -12420
rect 8283 -12454 8317 -12420
rect 8439 -12454 8473 -12420
rect 8544 -12454 8578 -12420
rect 8704 -12454 8738 -12420
rect 8801 -12454 8835 -12420
rect 8998 -12439 9032 -12405
rect 9262 -12439 9296 -12405
rect 9458 -12446 9492 -12412
rect 10090 -12446 10124 -12412
rect 10378 -12439 10412 -12405
rect 10642 -12439 10676 -12405
rect 10761 -12454 10795 -12420
rect 10859 -12454 10893 -12420
rect 11015 -12454 11049 -12420
rect 11120 -12454 11154 -12420
rect 11280 -12454 11314 -12420
rect 11377 -12454 11411 -12420
rect 11666 -12439 11700 -12405
rect 11930 -12439 11964 -12405
rect 13690 -12465 13724 -12431
rect 13776 -12452 13810 -12418
rect 13862 -12452 13896 -12418
rect 13948 -12452 13982 -12418
rect 14034 -12452 14068 -12418
rect 14120 -12452 14154 -12418
rect 14206 -12461 14240 -12427
rect 14292 -12452 14326 -12418
rect 14378 -12461 14412 -12427
rect 14464 -12452 14498 -12418
rect 14550 -12461 14584 -12427
rect 14636 -12452 14670 -12418
rect 14722 -12461 14756 -12427
rect 14807 -12452 14841 -12418
rect 14893 -12461 14927 -12427
rect 14979 -12452 15013 -12418
rect 15065 -12461 15099 -12427
rect 15151 -12452 15185 -12418
rect 15237 -12461 15271 -12427
rect 15323 -12452 15357 -12418
rect 15409 -12461 15443 -12427
rect 15622 -12446 15656 -12412
rect 16622 -12446 16656 -12412
rect -2962 -12636 -2928 -12602
rect -2330 -12636 -2296 -12602
rect -1582 -12636 -1548 -12602
rect -950 -12636 -916 -12602
rect -846 -12636 -812 -12602
rect -214 -12636 -180 -12602
rect -18 -12643 16 -12609
rect 246 -12643 280 -12609
rect 443 -12628 477 -12594
rect 540 -12628 574 -12594
rect 700 -12628 734 -12594
rect 805 -12628 839 -12594
rect 961 -12628 995 -12594
rect 1059 -12628 1093 -12594
rect 1270 -12643 1304 -12609
rect 1534 -12643 1568 -12609
rect 1730 -12636 1764 -12602
rect 2362 -12636 2396 -12602
rect 2558 -12643 2592 -12609
rect 2822 -12643 2856 -12609
rect 3019 -12628 3053 -12594
rect 3116 -12628 3150 -12594
rect 3276 -12628 3310 -12594
rect 3381 -12628 3415 -12594
rect 3537 -12628 3571 -12594
rect 3635 -12628 3669 -12594
rect 3846 -12643 3880 -12609
rect 4110 -12643 4144 -12609
rect 4306 -12636 4340 -12602
rect 4938 -12636 4972 -12602
rect 5134 -12643 5168 -12609
rect 5398 -12643 5432 -12609
rect 5595 -12628 5629 -12594
rect 5692 -12628 5726 -12594
rect 5852 -12628 5886 -12594
rect 5957 -12628 5991 -12594
rect 6113 -12628 6147 -12594
rect 6211 -12628 6245 -12594
rect 6422 -12643 6456 -12609
rect 6686 -12643 6720 -12609
rect 6882 -12636 6916 -12602
rect 7514 -12636 7548 -12602
rect 7710 -12643 7744 -12609
rect 7974 -12643 8008 -12609
rect 8171 -12628 8205 -12594
rect 8268 -12628 8302 -12594
rect 8428 -12628 8462 -12594
rect 8533 -12628 8567 -12594
rect 8689 -12628 8723 -12594
rect 8787 -12628 8821 -12594
rect 8998 -12643 9032 -12609
rect 9262 -12643 9296 -12609
rect 9458 -12636 9492 -12602
rect 10090 -12636 10124 -12602
rect 10378 -12643 10412 -12609
rect 10642 -12643 10676 -12609
rect 10747 -12628 10781 -12594
rect 10844 -12628 10878 -12594
rect 11004 -12628 11038 -12594
rect 11109 -12628 11143 -12594
rect 11265 -12628 11299 -12594
rect 11363 -12628 11397 -12594
rect 11666 -12643 11700 -12609
rect 11930 -12643 11964 -12609
rect 12588 -12619 12622 -12585
rect 12674 -12630 12708 -12596
rect 12760 -12619 12794 -12585
rect 12846 -12630 12880 -12596
rect 12932 -12619 12966 -12585
rect 13230 -12643 13264 -12609
rect 13494 -12643 13528 -12609
rect 13690 -12617 13724 -12583
rect 13776 -12630 13810 -12596
rect 13862 -12630 13896 -12596
rect 13948 -12630 13982 -12596
rect 14034 -12630 14068 -12596
rect 14120 -12630 14154 -12596
rect 14206 -12621 14240 -12587
rect 14292 -12630 14326 -12596
rect 14378 -12621 14412 -12587
rect 14464 -12630 14498 -12596
rect 14550 -12621 14584 -12587
rect 14636 -12630 14670 -12596
rect 14722 -12621 14756 -12587
rect 14807 -12630 14841 -12596
rect 14893 -12621 14927 -12587
rect 14979 -12630 15013 -12596
rect 15065 -12621 15099 -12587
rect 15151 -12630 15185 -12596
rect 15237 -12621 15271 -12587
rect 15323 -12630 15357 -12596
rect 15409 -12621 15443 -12587
rect 15622 -12636 15656 -12602
rect 16622 -12636 16656 -12602
rect -2962 -13534 -2928 -13500
rect -2330 -13534 -2296 -13500
rect -1582 -13534 -1548 -13500
rect -950 -13534 -916 -13500
rect -846 -13534 -812 -13500
rect -214 -13534 -180 -13500
rect -18 -13527 16 -13493
rect 246 -13527 280 -13493
rect 457 -13542 491 -13508
rect 555 -13542 589 -13508
rect 711 -13542 745 -13508
rect 816 -13542 850 -13508
rect 976 -13542 1010 -13508
rect 1073 -13542 1107 -13508
rect 1270 -13527 1304 -13493
rect 1534 -13527 1568 -13493
rect 1730 -13534 1764 -13500
rect 2362 -13534 2396 -13500
rect 2558 -13527 2592 -13493
rect 2822 -13527 2856 -13493
rect 3033 -13542 3067 -13508
rect 3131 -13542 3165 -13508
rect 3287 -13542 3321 -13508
rect 3392 -13542 3426 -13508
rect 3552 -13542 3586 -13508
rect 3649 -13542 3683 -13508
rect 3846 -13527 3880 -13493
rect 4110 -13527 4144 -13493
rect 4306 -13534 4340 -13500
rect 4938 -13534 4972 -13500
rect 5134 -13527 5168 -13493
rect 5398 -13527 5432 -13493
rect 5609 -13542 5643 -13508
rect 5707 -13542 5741 -13508
rect 5863 -13542 5897 -13508
rect 5968 -13542 6002 -13508
rect 6128 -13542 6162 -13508
rect 6225 -13542 6259 -13508
rect 6422 -13527 6456 -13493
rect 6686 -13527 6720 -13493
rect 6882 -13534 6916 -13500
rect 7514 -13534 7548 -13500
rect 7710 -13527 7744 -13493
rect 7974 -13527 8008 -13493
rect 8185 -13542 8219 -13508
rect 8283 -13542 8317 -13508
rect 8439 -13542 8473 -13508
rect 8544 -13542 8578 -13508
rect 8704 -13542 8738 -13508
rect 8801 -13542 8835 -13508
rect 8998 -13527 9032 -13493
rect 9262 -13527 9296 -13493
rect 9458 -13534 9492 -13500
rect 10090 -13534 10124 -13500
rect 10378 -13527 10412 -13493
rect 10642 -13527 10676 -13493
rect 10761 -13542 10795 -13508
rect 10859 -13542 10893 -13508
rect 11015 -13542 11049 -13508
rect 11120 -13542 11154 -13508
rect 11280 -13542 11314 -13508
rect 11377 -13542 11411 -13508
rect 11666 -13527 11700 -13493
rect 11930 -13527 11964 -13493
rect 13690 -13553 13724 -13519
rect 13776 -13540 13810 -13506
rect 13862 -13540 13896 -13506
rect 13948 -13540 13982 -13506
rect 14034 -13540 14068 -13506
rect 14120 -13540 14154 -13506
rect 14206 -13549 14240 -13515
rect 14292 -13540 14326 -13506
rect 14378 -13549 14412 -13515
rect 14464 -13540 14498 -13506
rect 14550 -13549 14584 -13515
rect 14636 -13540 14670 -13506
rect 14722 -13549 14756 -13515
rect 14807 -13540 14841 -13506
rect 14893 -13549 14927 -13515
rect 14979 -13540 15013 -13506
rect 15065 -13549 15099 -13515
rect 15151 -13540 15185 -13506
rect 15237 -13549 15271 -13515
rect 15323 -13540 15357 -13506
rect 15409 -13549 15443 -13515
rect 15622 -13534 15656 -13500
rect 16622 -13534 16656 -13500
rect -2962 -13724 -2928 -13690
rect -2330 -13724 -2296 -13690
rect -1398 -13731 -1364 -13697
rect -1134 -13731 -1100 -13697
rect -934 -13705 -900 -13671
rect -934 -13773 -900 -13739
rect -766 -13705 -732 -13671
rect -766 -13773 -732 -13739
rect -570 -13731 -536 -13697
rect -306 -13731 -272 -13697
rect -16 -13707 18 -13673
rect 70 -13718 104 -13684
rect 156 -13707 190 -13673
rect 242 -13718 276 -13684
rect 328 -13707 362 -13673
rect 626 -13731 660 -13697
rect 890 -13731 924 -13697
rect 1169 -13716 1203 -13682
rect 1253 -13714 1287 -13680
rect 1454 -13731 1488 -13697
rect 1718 -13731 1752 -13697
rect 1914 -13731 1948 -13697
rect 2178 -13731 2212 -13697
rect 2375 -13716 2409 -13682
rect 2472 -13716 2506 -13682
rect 2632 -13716 2666 -13682
rect 2737 -13716 2771 -13682
rect 2893 -13716 2927 -13682
rect 2991 -13716 3025 -13682
rect 3202 -13731 3236 -13697
rect 3466 -13731 3500 -13697
rect 4398 -13724 4432 -13690
rect 5398 -13724 5432 -13690
rect 6422 -13731 6456 -13697
rect 6686 -13731 6720 -13697
rect 6883 -13716 6917 -13682
rect 6980 -13716 7014 -13682
rect 7140 -13716 7174 -13682
rect 7245 -13716 7279 -13682
rect 7401 -13716 7435 -13682
rect 7499 -13716 7533 -13682
rect 7710 -13731 7744 -13697
rect 7974 -13731 8008 -13697
rect 8171 -13716 8205 -13682
rect 8268 -13716 8302 -13682
rect 8428 -13716 8462 -13682
rect 8533 -13716 8567 -13682
rect 8689 -13716 8723 -13682
rect 8787 -13716 8821 -13682
rect 8998 -13731 9032 -13697
rect 9262 -13731 9296 -13697
rect 9459 -13716 9493 -13682
rect 9556 -13716 9590 -13682
rect 9716 -13716 9750 -13682
rect 9821 -13716 9855 -13682
rect 9977 -13716 10011 -13682
rect 10075 -13716 10109 -13682
rect 10286 -13731 10320 -13697
rect 10550 -13731 10584 -13697
rect 10746 -13705 10780 -13671
rect 10746 -13773 10780 -13739
rect 10830 -13705 10864 -13671
rect 10914 -13705 10948 -13671
rect 10914 -13773 10948 -13739
rect 10998 -13705 11032 -13671
rect 11082 -13705 11116 -13671
rect 11082 -13773 11116 -13739
rect 11166 -13773 11200 -13739
rect 11250 -13705 11284 -13671
rect 11334 -13773 11368 -13739
rect 11418 -13705 11452 -13671
rect 11418 -13773 11452 -13739
rect 11666 -13731 11700 -13697
rect 11930 -13731 11964 -13697
rect 13598 -13724 13632 -13690
rect 14598 -13724 14632 -13690
rect 14794 -13724 14828 -13690
rect 15794 -13724 15828 -13690
rect 15990 -13724 16024 -13690
rect 16622 -13724 16656 -13690
<< pdiffc >>
rect -2962 -105 -2928 -71
rect -2962 -207 -2928 -173
rect -2330 -105 -2296 -71
rect -2330 -207 -2296 -173
rect -1398 -105 -1364 -71
rect -1398 -207 -1364 -173
rect -1134 -105 -1100 -71
rect -1134 -207 -1100 -173
rect -934 -105 -900 -71
rect -934 -173 -900 -139
rect -934 -241 -900 -207
rect -850 -105 -816 -71
rect -850 -173 -816 -139
rect -850 -241 -816 -207
rect -766 -105 -732 -71
rect -766 -173 -732 -139
rect -766 -241 -732 -207
rect -570 -105 -536 -71
rect -570 -207 -536 -173
rect -306 -105 -272 -71
rect -306 -207 -272 -173
rect -102 -112 -68 -78
rect -102 -180 -68 -146
rect -16 -119 18 -85
rect -16 -207 18 -173
rect 70 -112 104 -78
rect 70 -180 104 -146
rect 156 -119 190 -85
rect 156 -207 190 -173
rect 242 -112 276 -78
rect 242 -180 276 -146
rect 328 -119 362 -85
rect 328 -207 362 -173
rect 414 -112 448 -78
rect 414 -180 448 -146
rect 626 -105 660 -71
rect 626 -207 660 -173
rect 890 -105 924 -71
rect 890 -207 924 -173
rect 1086 -105 1120 -71
rect 1086 -207 1120 -173
rect 1170 -105 1204 -71
rect 1170 -207 1204 -173
rect 1254 -105 1288 -71
rect 1254 -207 1288 -173
rect 1454 -105 1488 -71
rect 1454 -207 1488 -173
rect 1718 -105 1752 -71
rect 1718 -207 1752 -173
rect 1914 -105 1948 -71
rect 1914 -207 1948 -173
rect 2178 -105 2212 -71
rect 2178 -207 2212 -173
rect 2375 -112 2409 -78
rect 2375 -180 2409 -146
rect 2475 -112 2509 -78
rect 2475 -180 2509 -146
rect 2633 -112 2667 -78
rect 2633 -180 2667 -146
rect 2737 -113 2771 -79
rect 2737 -181 2771 -147
rect 2893 -112 2927 -78
rect 2893 -180 2927 -146
rect 2991 -113 3025 -79
rect 2991 -181 3025 -147
rect 3202 -105 3236 -71
rect 3202 -207 3236 -173
rect 3466 -105 3500 -71
rect 3466 -207 3500 -173
rect 4398 -105 4432 -71
rect 4398 -207 4432 -173
rect 5398 -105 5432 -71
rect 5398 -207 5432 -173
rect 6422 -105 6456 -71
rect 6422 -207 6456 -173
rect 6686 -105 6720 -71
rect 6686 -207 6720 -173
rect 6883 -112 6917 -78
rect 6883 -180 6917 -146
rect 6983 -112 7017 -78
rect 6983 -180 7017 -146
rect 7141 -112 7175 -78
rect 7141 -180 7175 -146
rect 7245 -113 7279 -79
rect 7245 -181 7279 -147
rect 7401 -112 7435 -78
rect 7401 -180 7435 -146
rect 7499 -113 7533 -79
rect 7499 -181 7533 -147
rect 7710 -105 7744 -71
rect 7710 -207 7744 -173
rect 7974 -105 8008 -71
rect 7974 -207 8008 -173
rect 8171 -112 8205 -78
rect 8171 -180 8205 -146
rect 8271 -112 8305 -78
rect 8271 -180 8305 -146
rect 8429 -112 8463 -78
rect 8429 -180 8463 -146
rect 8533 -113 8567 -79
rect 8533 -181 8567 -147
rect 8689 -112 8723 -78
rect 8689 -180 8723 -146
rect 8787 -113 8821 -79
rect 8787 -181 8821 -147
rect 8998 -105 9032 -71
rect 8998 -207 9032 -173
rect 9262 -105 9296 -71
rect 9262 -207 9296 -173
rect 9459 -112 9493 -78
rect 9459 -180 9493 -146
rect 9559 -112 9593 -78
rect 9559 -180 9593 -146
rect 9717 -112 9751 -78
rect 9717 -180 9751 -146
rect 9821 -113 9855 -79
rect 9821 -181 9855 -147
rect 9977 -112 10011 -78
rect 9977 -180 10011 -146
rect 10075 -113 10109 -79
rect 10075 -181 10109 -147
rect 10286 -105 10320 -71
rect 10286 -207 10320 -173
rect 10550 -105 10584 -71
rect 10550 -207 10584 -173
rect 10746 -105 10780 -71
rect 10746 -173 10780 -139
rect 10746 -241 10780 -207
rect 10830 -105 10864 -71
rect 10830 -173 10864 -139
rect 10830 -241 10864 -207
rect 10914 -105 10948 -71
rect 10914 -173 10948 -139
rect 10998 -105 11032 -71
rect 10998 -173 11032 -139
rect 10998 -241 11032 -207
rect 11082 -105 11116 -71
rect 11082 -173 11116 -139
rect 11166 -105 11200 -71
rect 11166 -173 11200 -139
rect 11166 -241 11200 -207
rect 11250 -105 11284 -71
rect 11250 -173 11284 -139
rect 11334 -105 11368 -71
rect 11334 -173 11368 -139
rect 11334 -241 11368 -207
rect 11418 -105 11452 -71
rect 11418 -173 11452 -139
rect 11666 -105 11700 -71
rect 11666 -207 11700 -173
rect 11930 -105 11964 -71
rect 11930 -207 11964 -173
rect 13598 -105 13632 -71
rect 13598 -207 13632 -173
rect 14598 -105 14632 -71
rect 14598 -207 14632 -173
rect 14794 -105 14828 -71
rect 14794 -207 14828 -173
rect 15794 -105 15828 -71
rect 15794 -207 15828 -173
rect 15990 -105 16024 -71
rect 15990 -207 16024 -173
rect 16622 -105 16656 -71
rect 16622 -207 16656 -173
rect -2962 -939 -2928 -905
rect -2962 -1041 -2928 -1007
rect -2330 -939 -2296 -905
rect -2330 -1041 -2296 -1007
rect -1582 -939 -1548 -905
rect -1582 -1041 -1548 -1007
rect -950 -939 -916 -905
rect -950 -1041 -916 -1007
rect -846 -939 -812 -905
rect -846 -1041 -812 -1007
rect -214 -939 -180 -905
rect -214 -1041 -180 -1007
rect -18 -939 16 -905
rect -18 -1041 16 -1007
rect 246 -939 280 -905
rect 246 -1041 280 -1007
rect 457 -965 491 -931
rect 457 -1033 491 -999
rect 555 -966 589 -932
rect 555 -1034 589 -1000
rect 711 -965 745 -931
rect 711 -1033 745 -999
rect 815 -966 849 -932
rect 815 -1034 849 -1000
rect 973 -966 1007 -932
rect 973 -1034 1007 -1000
rect 1073 -966 1107 -932
rect 1073 -1034 1107 -1000
rect 1270 -939 1304 -905
rect 1270 -1041 1304 -1007
rect 1534 -939 1568 -905
rect 1534 -1041 1568 -1007
rect 1730 -939 1764 -905
rect 1730 -1041 1764 -1007
rect 2362 -939 2396 -905
rect 2362 -1041 2396 -1007
rect 2558 -939 2592 -905
rect 2558 -1041 2592 -1007
rect 2822 -939 2856 -905
rect 2822 -1041 2856 -1007
rect 3033 -965 3067 -931
rect 3033 -1033 3067 -999
rect 3131 -966 3165 -932
rect 3131 -1034 3165 -1000
rect 3287 -965 3321 -931
rect 3287 -1033 3321 -999
rect 3391 -966 3425 -932
rect 3391 -1034 3425 -1000
rect 3549 -966 3583 -932
rect 3549 -1034 3583 -1000
rect 3649 -966 3683 -932
rect 3649 -1034 3683 -1000
rect 3846 -939 3880 -905
rect 3846 -1041 3880 -1007
rect 4110 -939 4144 -905
rect 4110 -1041 4144 -1007
rect 4306 -939 4340 -905
rect 4306 -1041 4340 -1007
rect 4938 -939 4972 -905
rect 4938 -1041 4972 -1007
rect 5134 -939 5168 -905
rect 5134 -1041 5168 -1007
rect 5398 -939 5432 -905
rect 5398 -1041 5432 -1007
rect 5609 -965 5643 -931
rect 5609 -1033 5643 -999
rect 5707 -966 5741 -932
rect 5707 -1034 5741 -1000
rect 5863 -965 5897 -931
rect 5863 -1033 5897 -999
rect 5967 -966 6001 -932
rect 5967 -1034 6001 -1000
rect 6125 -966 6159 -932
rect 6125 -1034 6159 -1000
rect 6225 -966 6259 -932
rect 6225 -1034 6259 -1000
rect 6422 -939 6456 -905
rect 6422 -1041 6456 -1007
rect 6686 -939 6720 -905
rect 6686 -1041 6720 -1007
rect 6882 -939 6916 -905
rect 6882 -1041 6916 -1007
rect 7514 -939 7548 -905
rect 7514 -1041 7548 -1007
rect 7710 -939 7744 -905
rect 7710 -1041 7744 -1007
rect 7974 -939 8008 -905
rect 7974 -1041 8008 -1007
rect 8185 -965 8219 -931
rect 8185 -1033 8219 -999
rect 8283 -966 8317 -932
rect 8283 -1034 8317 -1000
rect 8439 -965 8473 -931
rect 8439 -1033 8473 -999
rect 8543 -966 8577 -932
rect 8543 -1034 8577 -1000
rect 8701 -966 8735 -932
rect 8701 -1034 8735 -1000
rect 8801 -966 8835 -932
rect 8801 -1034 8835 -1000
rect 8998 -939 9032 -905
rect 8998 -1041 9032 -1007
rect 9262 -939 9296 -905
rect 9262 -1041 9296 -1007
rect 9458 -939 9492 -905
rect 9458 -1041 9492 -1007
rect 10090 -939 10124 -905
rect 10090 -1041 10124 -1007
rect 10378 -939 10412 -905
rect 10378 -1041 10412 -1007
rect 10642 -939 10676 -905
rect 10642 -1041 10676 -1007
rect 10761 -965 10795 -931
rect 10761 -1033 10795 -999
rect 10859 -966 10893 -932
rect 10859 -1034 10893 -1000
rect 11015 -965 11049 -931
rect 11015 -1033 11049 -999
rect 11119 -966 11153 -932
rect 11119 -1034 11153 -1000
rect 11277 -966 11311 -932
rect 11277 -1034 11311 -1000
rect 11377 -966 11411 -932
rect 11377 -1034 11411 -1000
rect 11666 -939 11700 -905
rect 11666 -1041 11700 -1007
rect 11930 -939 11964 -905
rect 11930 -1041 11964 -1007
rect 13690 -973 13724 -939
rect 13690 -1041 13724 -1007
rect 13776 -965 13810 -931
rect 13776 -1033 13810 -999
rect 13862 -973 13896 -939
rect 13862 -1041 13896 -1007
rect 13948 -957 13982 -923
rect 13948 -1025 13982 -991
rect 14034 -973 14068 -939
rect 14034 -1041 14068 -1007
rect 14120 -911 14154 -877
rect 14120 -997 14154 -963
rect 14206 -1017 14240 -983
rect 14292 -911 14326 -877
rect 14292 -997 14326 -963
rect 14378 -1017 14412 -983
rect 14464 -911 14498 -877
rect 14464 -997 14498 -963
rect 14550 -1017 14584 -983
rect 14636 -911 14670 -877
rect 14636 -997 14670 -963
rect 14722 -1017 14756 -983
rect 14807 -911 14841 -877
rect 14807 -997 14841 -963
rect 14893 -1017 14927 -983
rect 14979 -911 15013 -877
rect 14979 -997 15013 -963
rect 15065 -1017 15099 -983
rect 15151 -911 15185 -877
rect 15151 -997 15185 -963
rect 15237 -1017 15271 -983
rect 15323 -911 15357 -877
rect 15323 -997 15357 -963
rect 15409 -1017 15443 -983
rect 15622 -939 15656 -905
rect 15622 -1041 15656 -1007
rect 16622 -939 16656 -905
rect 16622 -1041 16656 -1007
rect -2962 -1193 -2928 -1159
rect -2962 -1295 -2928 -1261
rect -2330 -1193 -2296 -1159
rect -2330 -1295 -2296 -1261
rect -1582 -1193 -1548 -1159
rect -1582 -1295 -1548 -1261
rect -950 -1193 -916 -1159
rect -950 -1295 -916 -1261
rect -846 -1193 -812 -1159
rect -846 -1295 -812 -1261
rect -214 -1193 -180 -1159
rect -214 -1295 -180 -1261
rect -18 -1193 16 -1159
rect -18 -1295 16 -1261
rect 246 -1193 280 -1159
rect 246 -1295 280 -1261
rect 443 -1200 477 -1166
rect 443 -1268 477 -1234
rect 543 -1200 577 -1166
rect 543 -1268 577 -1234
rect 701 -1200 735 -1166
rect 701 -1268 735 -1234
rect 805 -1201 839 -1167
rect 805 -1269 839 -1235
rect 961 -1200 995 -1166
rect 961 -1268 995 -1234
rect 1059 -1201 1093 -1167
rect 1059 -1269 1093 -1235
rect 1270 -1193 1304 -1159
rect 1270 -1295 1304 -1261
rect 1534 -1193 1568 -1159
rect 1534 -1295 1568 -1261
rect 1730 -1193 1764 -1159
rect 1730 -1295 1764 -1261
rect 2362 -1193 2396 -1159
rect 2362 -1295 2396 -1261
rect 2558 -1193 2592 -1159
rect 2558 -1295 2592 -1261
rect 2822 -1193 2856 -1159
rect 2822 -1295 2856 -1261
rect 3019 -1200 3053 -1166
rect 3019 -1268 3053 -1234
rect 3119 -1200 3153 -1166
rect 3119 -1268 3153 -1234
rect 3277 -1200 3311 -1166
rect 3277 -1268 3311 -1234
rect 3381 -1201 3415 -1167
rect 3381 -1269 3415 -1235
rect 3537 -1200 3571 -1166
rect 3537 -1268 3571 -1234
rect 3635 -1201 3669 -1167
rect 3635 -1269 3669 -1235
rect 3846 -1193 3880 -1159
rect 3846 -1295 3880 -1261
rect 4110 -1193 4144 -1159
rect 4110 -1295 4144 -1261
rect 4306 -1193 4340 -1159
rect 4306 -1295 4340 -1261
rect 4938 -1193 4972 -1159
rect 4938 -1295 4972 -1261
rect 5134 -1193 5168 -1159
rect 5134 -1295 5168 -1261
rect 5398 -1193 5432 -1159
rect 5398 -1295 5432 -1261
rect 5595 -1200 5629 -1166
rect 5595 -1268 5629 -1234
rect 5695 -1200 5729 -1166
rect 5695 -1268 5729 -1234
rect 5853 -1200 5887 -1166
rect 5853 -1268 5887 -1234
rect 5957 -1201 5991 -1167
rect 5957 -1269 5991 -1235
rect 6113 -1200 6147 -1166
rect 6113 -1268 6147 -1234
rect 6211 -1201 6245 -1167
rect 6211 -1269 6245 -1235
rect 6422 -1193 6456 -1159
rect 6422 -1295 6456 -1261
rect 6686 -1193 6720 -1159
rect 6686 -1295 6720 -1261
rect 6882 -1193 6916 -1159
rect 6882 -1295 6916 -1261
rect 7514 -1193 7548 -1159
rect 7514 -1295 7548 -1261
rect 7710 -1193 7744 -1159
rect 7710 -1295 7744 -1261
rect 7974 -1193 8008 -1159
rect 7974 -1295 8008 -1261
rect 8171 -1200 8205 -1166
rect 8171 -1268 8205 -1234
rect 8271 -1200 8305 -1166
rect 8271 -1268 8305 -1234
rect 8429 -1200 8463 -1166
rect 8429 -1268 8463 -1234
rect 8533 -1201 8567 -1167
rect 8533 -1269 8567 -1235
rect 8689 -1200 8723 -1166
rect 8689 -1268 8723 -1234
rect 8787 -1201 8821 -1167
rect 8787 -1269 8821 -1235
rect 8998 -1193 9032 -1159
rect 8998 -1295 9032 -1261
rect 9262 -1193 9296 -1159
rect 9262 -1295 9296 -1261
rect 9458 -1193 9492 -1159
rect 9458 -1295 9492 -1261
rect 10090 -1193 10124 -1159
rect 10090 -1295 10124 -1261
rect 10378 -1193 10412 -1159
rect 10378 -1295 10412 -1261
rect 10642 -1193 10676 -1159
rect 10642 -1295 10676 -1261
rect 10747 -1200 10781 -1166
rect 10747 -1268 10781 -1234
rect 10847 -1200 10881 -1166
rect 10847 -1268 10881 -1234
rect 11005 -1200 11039 -1166
rect 11005 -1268 11039 -1234
rect 11109 -1201 11143 -1167
rect 11109 -1269 11143 -1235
rect 11265 -1200 11299 -1166
rect 11265 -1268 11299 -1234
rect 11363 -1201 11397 -1167
rect 11363 -1269 11397 -1235
rect 11666 -1193 11700 -1159
rect 11666 -1295 11700 -1261
rect 11930 -1193 11964 -1159
rect 11930 -1295 11964 -1261
rect 12502 -1200 12536 -1166
rect 12502 -1268 12536 -1234
rect 12588 -1207 12622 -1173
rect 12588 -1295 12622 -1261
rect 12674 -1200 12708 -1166
rect 12674 -1268 12708 -1234
rect 12760 -1207 12794 -1173
rect 12760 -1295 12794 -1261
rect 12846 -1200 12880 -1166
rect 12846 -1268 12880 -1234
rect 12932 -1207 12966 -1173
rect 12932 -1295 12966 -1261
rect 13018 -1200 13052 -1166
rect 13018 -1268 13052 -1234
rect 13230 -1193 13264 -1159
rect 13230 -1295 13264 -1261
rect 13494 -1193 13528 -1159
rect 13494 -1295 13528 -1261
rect 13690 -1193 13724 -1159
rect 13690 -1261 13724 -1227
rect 13776 -1201 13810 -1167
rect 13776 -1269 13810 -1235
rect 13862 -1193 13896 -1159
rect 13862 -1261 13896 -1227
rect 13948 -1209 13982 -1175
rect 13948 -1277 13982 -1243
rect 14034 -1193 14068 -1159
rect 14034 -1261 14068 -1227
rect 14120 -1237 14154 -1203
rect 14120 -1323 14154 -1289
rect 14206 -1217 14240 -1183
rect 14292 -1237 14326 -1203
rect 14292 -1323 14326 -1289
rect 14378 -1217 14412 -1183
rect 14464 -1237 14498 -1203
rect 14464 -1323 14498 -1289
rect 14550 -1217 14584 -1183
rect 14636 -1237 14670 -1203
rect 14636 -1323 14670 -1289
rect 14722 -1217 14756 -1183
rect 14807 -1237 14841 -1203
rect 14807 -1323 14841 -1289
rect 14893 -1217 14927 -1183
rect 14979 -1237 15013 -1203
rect 14979 -1323 15013 -1289
rect 15065 -1217 15099 -1183
rect 15151 -1237 15185 -1203
rect 15151 -1323 15185 -1289
rect 15237 -1217 15271 -1183
rect 15323 -1237 15357 -1203
rect 15323 -1323 15357 -1289
rect 15409 -1217 15443 -1183
rect 15622 -1193 15656 -1159
rect 15622 -1295 15656 -1261
rect 16622 -1193 16656 -1159
rect 16622 -1295 16656 -1261
rect -2962 -2027 -2928 -1993
rect -2962 -2129 -2928 -2095
rect -2330 -2027 -2296 -1993
rect -2330 -2129 -2296 -2095
rect -1582 -2027 -1548 -1993
rect -1582 -2129 -1548 -2095
rect -950 -2027 -916 -1993
rect -950 -2129 -916 -2095
rect -831 -2053 -797 -2019
rect -831 -2121 -797 -2087
rect -733 -2054 -699 -2020
rect -733 -2122 -699 -2088
rect -577 -2053 -543 -2019
rect -577 -2121 -543 -2087
rect -473 -2054 -439 -2020
rect -473 -2122 -439 -2088
rect -315 -2054 -281 -2020
rect -315 -2122 -281 -2088
rect -215 -2054 -181 -2020
rect -215 -2122 -181 -2088
rect -18 -2027 16 -1993
rect -18 -2129 16 -2095
rect 246 -2027 280 -1993
rect 246 -2129 280 -2095
rect 457 -2053 491 -2019
rect 457 -2121 491 -2087
rect 555 -2054 589 -2020
rect 555 -2122 589 -2088
rect 711 -2053 745 -2019
rect 711 -2121 745 -2087
rect 815 -2054 849 -2020
rect 815 -2122 849 -2088
rect 973 -2054 1007 -2020
rect 973 -2122 1007 -2088
rect 1073 -2054 1107 -2020
rect 1073 -2122 1107 -2088
rect 1270 -2027 1304 -1993
rect 1270 -2129 1304 -2095
rect 1534 -2027 1568 -1993
rect 1534 -2129 1568 -2095
rect 1730 -2027 1764 -1993
rect 1730 -2129 1764 -2095
rect 2362 -2027 2396 -1993
rect 2362 -2129 2396 -2095
rect 2558 -2027 2592 -1993
rect 2558 -2129 2592 -2095
rect 2822 -2027 2856 -1993
rect 2822 -2129 2856 -2095
rect 3033 -2053 3067 -2019
rect 3033 -2121 3067 -2087
rect 3131 -2054 3165 -2020
rect 3131 -2122 3165 -2088
rect 3287 -2053 3321 -2019
rect 3287 -2121 3321 -2087
rect 3391 -2054 3425 -2020
rect 3391 -2122 3425 -2088
rect 3549 -2054 3583 -2020
rect 3549 -2122 3583 -2088
rect 3649 -2054 3683 -2020
rect 3649 -2122 3683 -2088
rect 3846 -2027 3880 -1993
rect 3846 -2129 3880 -2095
rect 4110 -2027 4144 -1993
rect 4110 -2129 4144 -2095
rect 4306 -2027 4340 -1993
rect 4306 -2129 4340 -2095
rect 4938 -2027 4972 -1993
rect 4938 -2129 4972 -2095
rect 5134 -2027 5168 -1993
rect 5134 -2129 5168 -2095
rect 5398 -2027 5432 -1993
rect 5398 -2129 5432 -2095
rect 5609 -2053 5643 -2019
rect 5609 -2121 5643 -2087
rect 5707 -2054 5741 -2020
rect 5707 -2122 5741 -2088
rect 5863 -2053 5897 -2019
rect 5863 -2121 5897 -2087
rect 5967 -2054 6001 -2020
rect 5967 -2122 6001 -2088
rect 6125 -2054 6159 -2020
rect 6125 -2122 6159 -2088
rect 6225 -2054 6259 -2020
rect 6225 -2122 6259 -2088
rect 6422 -2027 6456 -1993
rect 6422 -2129 6456 -2095
rect 6686 -2027 6720 -1993
rect 6686 -2129 6720 -2095
rect 6882 -2027 6916 -1993
rect 6882 -2129 6916 -2095
rect 7514 -2027 7548 -1993
rect 7514 -2129 7548 -2095
rect 7710 -2027 7744 -1993
rect 7710 -2129 7744 -2095
rect 7974 -2027 8008 -1993
rect 7974 -2129 8008 -2095
rect 8185 -2053 8219 -2019
rect 8185 -2121 8219 -2087
rect 8283 -2054 8317 -2020
rect 8283 -2122 8317 -2088
rect 8439 -2053 8473 -2019
rect 8439 -2121 8473 -2087
rect 8543 -2054 8577 -2020
rect 8543 -2122 8577 -2088
rect 8701 -2054 8735 -2020
rect 8701 -2122 8735 -2088
rect 8801 -2054 8835 -2020
rect 8801 -2122 8835 -2088
rect 8998 -2027 9032 -1993
rect 8998 -2129 9032 -2095
rect 9262 -2027 9296 -1993
rect 9262 -2129 9296 -2095
rect 9458 -2027 9492 -1993
rect 9458 -2129 9492 -2095
rect 10090 -2027 10124 -1993
rect 10090 -2129 10124 -2095
rect 10378 -2027 10412 -1993
rect 10378 -2129 10412 -2095
rect 10642 -2027 10676 -1993
rect 10642 -2129 10676 -2095
rect 10761 -2053 10795 -2019
rect 10761 -2121 10795 -2087
rect 10859 -2054 10893 -2020
rect 10859 -2122 10893 -2088
rect 11015 -2053 11049 -2019
rect 11015 -2121 11049 -2087
rect 11119 -2054 11153 -2020
rect 11119 -2122 11153 -2088
rect 11277 -2054 11311 -2020
rect 11277 -2122 11311 -2088
rect 11377 -2054 11411 -2020
rect 11377 -2122 11411 -2088
rect 11666 -2027 11700 -1993
rect 11666 -2129 11700 -2095
rect 11930 -2027 11964 -1993
rect 11930 -2129 11964 -2095
rect 13690 -2061 13724 -2027
rect 13690 -2129 13724 -2095
rect 13776 -2053 13810 -2019
rect 13776 -2121 13810 -2087
rect 13862 -2061 13896 -2027
rect 13862 -2129 13896 -2095
rect 13948 -2045 13982 -2011
rect 13948 -2113 13982 -2079
rect 14034 -2061 14068 -2027
rect 14034 -2129 14068 -2095
rect 14120 -1999 14154 -1965
rect 14120 -2085 14154 -2051
rect 14206 -2105 14240 -2071
rect 14292 -1999 14326 -1965
rect 14292 -2085 14326 -2051
rect 14378 -2105 14412 -2071
rect 14464 -1999 14498 -1965
rect 14464 -2085 14498 -2051
rect 14550 -2105 14584 -2071
rect 14636 -1999 14670 -1965
rect 14636 -2085 14670 -2051
rect 14722 -2105 14756 -2071
rect 14807 -1999 14841 -1965
rect 14807 -2085 14841 -2051
rect 14893 -2105 14927 -2071
rect 14979 -1999 15013 -1965
rect 14979 -2085 15013 -2051
rect 15065 -2105 15099 -2071
rect 15151 -1999 15185 -1965
rect 15151 -2085 15185 -2051
rect 15237 -2105 15271 -2071
rect 15323 -1999 15357 -1965
rect 15323 -2085 15357 -2051
rect 15409 -2105 15443 -2071
rect 15622 -2027 15656 -1993
rect 15622 -2129 15656 -2095
rect 16622 -2027 16656 -1993
rect 16622 -2129 16656 -2095
rect -2962 -2281 -2928 -2247
rect -2962 -2383 -2928 -2349
rect -2330 -2281 -2296 -2247
rect -2330 -2383 -2296 -2349
rect -1582 -2281 -1548 -2247
rect -1582 -2383 -1548 -2349
rect -950 -2281 -916 -2247
rect -950 -2383 -916 -2349
rect -846 -2281 -812 -2247
rect -846 -2383 -812 -2349
rect -214 -2281 -180 -2247
rect -214 -2383 -180 -2349
rect -18 -2281 16 -2247
rect -18 -2383 16 -2349
rect 246 -2281 280 -2247
rect 246 -2383 280 -2349
rect 443 -2288 477 -2254
rect 443 -2356 477 -2322
rect 543 -2288 577 -2254
rect 543 -2356 577 -2322
rect 701 -2288 735 -2254
rect 701 -2356 735 -2322
rect 805 -2289 839 -2255
rect 805 -2357 839 -2323
rect 961 -2288 995 -2254
rect 961 -2356 995 -2322
rect 1059 -2289 1093 -2255
rect 1059 -2357 1093 -2323
rect 1270 -2281 1304 -2247
rect 1270 -2383 1304 -2349
rect 1534 -2281 1568 -2247
rect 1534 -2383 1568 -2349
rect 1730 -2281 1764 -2247
rect 1730 -2383 1764 -2349
rect 2362 -2281 2396 -2247
rect 2362 -2383 2396 -2349
rect 2558 -2281 2592 -2247
rect 2558 -2383 2592 -2349
rect 2822 -2281 2856 -2247
rect 2822 -2383 2856 -2349
rect 3019 -2288 3053 -2254
rect 3019 -2356 3053 -2322
rect 3119 -2288 3153 -2254
rect 3119 -2356 3153 -2322
rect 3277 -2288 3311 -2254
rect 3277 -2356 3311 -2322
rect 3381 -2289 3415 -2255
rect 3381 -2357 3415 -2323
rect 3537 -2288 3571 -2254
rect 3537 -2356 3571 -2322
rect 3635 -2289 3669 -2255
rect 3635 -2357 3669 -2323
rect 3846 -2281 3880 -2247
rect 3846 -2383 3880 -2349
rect 4110 -2281 4144 -2247
rect 4110 -2383 4144 -2349
rect 4306 -2281 4340 -2247
rect 4306 -2383 4340 -2349
rect 4938 -2281 4972 -2247
rect 4938 -2383 4972 -2349
rect 5134 -2281 5168 -2247
rect 5134 -2383 5168 -2349
rect 5398 -2281 5432 -2247
rect 5398 -2383 5432 -2349
rect 5595 -2288 5629 -2254
rect 5595 -2356 5629 -2322
rect 5695 -2288 5729 -2254
rect 5695 -2356 5729 -2322
rect 5853 -2288 5887 -2254
rect 5853 -2356 5887 -2322
rect 5957 -2289 5991 -2255
rect 5957 -2357 5991 -2323
rect 6113 -2288 6147 -2254
rect 6113 -2356 6147 -2322
rect 6211 -2289 6245 -2255
rect 6211 -2357 6245 -2323
rect 6422 -2281 6456 -2247
rect 6422 -2383 6456 -2349
rect 6686 -2281 6720 -2247
rect 6686 -2383 6720 -2349
rect 6882 -2281 6916 -2247
rect 6882 -2383 6916 -2349
rect 7514 -2281 7548 -2247
rect 7514 -2383 7548 -2349
rect 7710 -2281 7744 -2247
rect 7710 -2383 7744 -2349
rect 7974 -2281 8008 -2247
rect 7974 -2383 8008 -2349
rect 8171 -2288 8205 -2254
rect 8171 -2356 8205 -2322
rect 8271 -2288 8305 -2254
rect 8271 -2356 8305 -2322
rect 8429 -2288 8463 -2254
rect 8429 -2356 8463 -2322
rect 8533 -2289 8567 -2255
rect 8533 -2357 8567 -2323
rect 8689 -2288 8723 -2254
rect 8689 -2356 8723 -2322
rect 8787 -2289 8821 -2255
rect 8787 -2357 8821 -2323
rect 8998 -2281 9032 -2247
rect 8998 -2383 9032 -2349
rect 9262 -2281 9296 -2247
rect 9262 -2383 9296 -2349
rect 9458 -2281 9492 -2247
rect 9458 -2383 9492 -2349
rect 10090 -2281 10124 -2247
rect 10090 -2383 10124 -2349
rect 10378 -2281 10412 -2247
rect 10378 -2383 10412 -2349
rect 10642 -2281 10676 -2247
rect 10642 -2383 10676 -2349
rect 10747 -2288 10781 -2254
rect 10747 -2356 10781 -2322
rect 10847 -2288 10881 -2254
rect 10847 -2356 10881 -2322
rect 11005 -2288 11039 -2254
rect 11005 -2356 11039 -2322
rect 11109 -2289 11143 -2255
rect 11109 -2357 11143 -2323
rect 11265 -2288 11299 -2254
rect 11265 -2356 11299 -2322
rect 11363 -2289 11397 -2255
rect 11363 -2357 11397 -2323
rect 11666 -2281 11700 -2247
rect 11666 -2383 11700 -2349
rect 11930 -2281 11964 -2247
rect 11930 -2383 11964 -2349
rect 12502 -2288 12536 -2254
rect 12502 -2356 12536 -2322
rect 12588 -2295 12622 -2261
rect 12588 -2383 12622 -2349
rect 12674 -2288 12708 -2254
rect 12674 -2356 12708 -2322
rect 12760 -2295 12794 -2261
rect 12760 -2383 12794 -2349
rect 12846 -2288 12880 -2254
rect 12846 -2356 12880 -2322
rect 12932 -2295 12966 -2261
rect 12932 -2383 12966 -2349
rect 13018 -2288 13052 -2254
rect 13018 -2356 13052 -2322
rect 13230 -2281 13264 -2247
rect 13230 -2383 13264 -2349
rect 13494 -2281 13528 -2247
rect 13494 -2383 13528 -2349
rect 13690 -2281 13724 -2247
rect 13690 -2349 13724 -2315
rect 13776 -2289 13810 -2255
rect 13776 -2357 13810 -2323
rect 13862 -2281 13896 -2247
rect 13862 -2349 13896 -2315
rect 13948 -2297 13982 -2263
rect 13948 -2365 13982 -2331
rect 14034 -2281 14068 -2247
rect 14034 -2349 14068 -2315
rect 14120 -2325 14154 -2291
rect 14120 -2411 14154 -2377
rect 14206 -2305 14240 -2271
rect 14292 -2325 14326 -2291
rect 14292 -2411 14326 -2377
rect 14378 -2305 14412 -2271
rect 14464 -2325 14498 -2291
rect 14464 -2411 14498 -2377
rect 14550 -2305 14584 -2271
rect 14636 -2325 14670 -2291
rect 14636 -2411 14670 -2377
rect 14722 -2305 14756 -2271
rect 14807 -2325 14841 -2291
rect 14807 -2411 14841 -2377
rect 14893 -2305 14927 -2271
rect 14979 -2325 15013 -2291
rect 14979 -2411 15013 -2377
rect 15065 -2305 15099 -2271
rect 15151 -2325 15185 -2291
rect 15151 -2411 15185 -2377
rect 15237 -2305 15271 -2271
rect 15323 -2325 15357 -2291
rect 15323 -2411 15357 -2377
rect 15409 -2305 15443 -2271
rect 15622 -2281 15656 -2247
rect 15622 -2383 15656 -2349
rect 16622 -2281 16656 -2247
rect 16622 -2383 16656 -2349
rect -2962 -3115 -2928 -3081
rect -2962 -3217 -2928 -3183
rect -2330 -3115 -2296 -3081
rect -2330 -3217 -2296 -3183
rect -1950 -3115 -1916 -3081
rect -1950 -3217 -1916 -3183
rect -1866 -3115 -1832 -3081
rect -1866 -3217 -1832 -3183
rect -1782 -3115 -1748 -3081
rect -1782 -3217 -1748 -3183
rect -1582 -3115 -1548 -3081
rect -1582 -3217 -1548 -3183
rect -950 -3115 -916 -3081
rect -950 -3217 -916 -3183
rect -846 -3115 -812 -3081
rect -846 -3217 -812 -3183
rect -214 -3115 -180 -3081
rect -214 -3217 -180 -3183
rect -18 -3115 16 -3081
rect -18 -3217 16 -3183
rect 246 -3115 280 -3081
rect 246 -3217 280 -3183
rect 457 -3141 491 -3107
rect 457 -3209 491 -3175
rect 555 -3142 589 -3108
rect 555 -3210 589 -3176
rect 711 -3141 745 -3107
rect 711 -3209 745 -3175
rect 815 -3142 849 -3108
rect 815 -3210 849 -3176
rect 973 -3142 1007 -3108
rect 973 -3210 1007 -3176
rect 1073 -3142 1107 -3108
rect 1073 -3210 1107 -3176
rect 1270 -3115 1304 -3081
rect 1270 -3217 1304 -3183
rect 1534 -3115 1568 -3081
rect 1534 -3217 1568 -3183
rect 1730 -3115 1764 -3081
rect 1730 -3217 1764 -3183
rect 2362 -3115 2396 -3081
rect 2362 -3217 2396 -3183
rect 2558 -3115 2592 -3081
rect 2558 -3217 2592 -3183
rect 2822 -3115 2856 -3081
rect 2822 -3217 2856 -3183
rect 3033 -3141 3067 -3107
rect 3033 -3209 3067 -3175
rect 3131 -3142 3165 -3108
rect 3131 -3210 3165 -3176
rect 3287 -3141 3321 -3107
rect 3287 -3209 3321 -3175
rect 3391 -3142 3425 -3108
rect 3391 -3210 3425 -3176
rect 3549 -3142 3583 -3108
rect 3549 -3210 3583 -3176
rect 3649 -3142 3683 -3108
rect 3649 -3210 3683 -3176
rect 3846 -3115 3880 -3081
rect 3846 -3217 3880 -3183
rect 4110 -3115 4144 -3081
rect 4110 -3217 4144 -3183
rect 4306 -3115 4340 -3081
rect 4306 -3217 4340 -3183
rect 4938 -3115 4972 -3081
rect 4938 -3217 4972 -3183
rect 5134 -3115 5168 -3081
rect 5134 -3217 5168 -3183
rect 5398 -3115 5432 -3081
rect 5398 -3217 5432 -3183
rect 5609 -3141 5643 -3107
rect 5609 -3209 5643 -3175
rect 5707 -3142 5741 -3108
rect 5707 -3210 5741 -3176
rect 5863 -3141 5897 -3107
rect 5863 -3209 5897 -3175
rect 5967 -3142 6001 -3108
rect 5967 -3210 6001 -3176
rect 6125 -3142 6159 -3108
rect 6125 -3210 6159 -3176
rect 6225 -3142 6259 -3108
rect 6225 -3210 6259 -3176
rect 6422 -3115 6456 -3081
rect 6422 -3217 6456 -3183
rect 6686 -3115 6720 -3081
rect 6686 -3217 6720 -3183
rect 6882 -3115 6916 -3081
rect 6882 -3217 6916 -3183
rect 7514 -3115 7548 -3081
rect 7514 -3217 7548 -3183
rect 7710 -3115 7744 -3081
rect 7710 -3217 7744 -3183
rect 7974 -3115 8008 -3081
rect 7974 -3217 8008 -3183
rect 8185 -3141 8219 -3107
rect 8185 -3209 8219 -3175
rect 8283 -3142 8317 -3108
rect 8283 -3210 8317 -3176
rect 8439 -3141 8473 -3107
rect 8439 -3209 8473 -3175
rect 8543 -3142 8577 -3108
rect 8543 -3210 8577 -3176
rect 8701 -3142 8735 -3108
rect 8701 -3210 8735 -3176
rect 8801 -3142 8835 -3108
rect 8801 -3210 8835 -3176
rect 8998 -3115 9032 -3081
rect 8998 -3217 9032 -3183
rect 9262 -3115 9296 -3081
rect 9262 -3217 9296 -3183
rect 9458 -3115 9492 -3081
rect 9458 -3217 9492 -3183
rect 10090 -3115 10124 -3081
rect 10090 -3217 10124 -3183
rect 10378 -3115 10412 -3081
rect 10378 -3217 10412 -3183
rect 10642 -3115 10676 -3081
rect 10642 -3217 10676 -3183
rect 10761 -3141 10795 -3107
rect 10761 -3209 10795 -3175
rect 10859 -3142 10893 -3108
rect 10859 -3210 10893 -3176
rect 11015 -3141 11049 -3107
rect 11015 -3209 11049 -3175
rect 11119 -3142 11153 -3108
rect 11119 -3210 11153 -3176
rect 11277 -3142 11311 -3108
rect 11277 -3210 11311 -3176
rect 11377 -3142 11411 -3108
rect 11377 -3210 11411 -3176
rect 11666 -3115 11700 -3081
rect 11666 -3217 11700 -3183
rect 11930 -3115 11964 -3081
rect 11930 -3217 11964 -3183
rect 13598 -3115 13632 -3081
rect 13598 -3217 13632 -3183
rect 14598 -3115 14632 -3081
rect 14598 -3217 14632 -3183
rect 14794 -3115 14828 -3081
rect 14794 -3217 14828 -3183
rect 15794 -3115 15828 -3081
rect 15794 -3217 15828 -3183
rect 15990 -3115 16024 -3081
rect 15990 -3217 16024 -3183
rect 16622 -3115 16656 -3081
rect 16622 -3217 16656 -3183
rect -2962 -3369 -2928 -3335
rect -2962 -3471 -2928 -3437
rect -2330 -3369 -2296 -3335
rect -2330 -3471 -2296 -3437
rect -1582 -3369 -1548 -3335
rect -1582 -3471 -1548 -3437
rect -950 -3369 -916 -3335
rect -950 -3471 -916 -3437
rect -846 -3369 -812 -3335
rect -846 -3471 -812 -3437
rect -214 -3369 -180 -3335
rect -214 -3471 -180 -3437
rect -18 -3369 16 -3335
rect -18 -3471 16 -3437
rect 246 -3369 280 -3335
rect 246 -3471 280 -3437
rect 457 -3377 491 -3343
rect 457 -3445 491 -3411
rect 555 -3376 589 -3342
rect 555 -3444 589 -3410
rect 711 -3377 745 -3343
rect 711 -3445 745 -3411
rect 815 -3376 849 -3342
rect 815 -3444 849 -3410
rect 973 -3376 1007 -3342
rect 973 -3444 1007 -3410
rect 1073 -3376 1107 -3342
rect 1073 -3444 1107 -3410
rect 1270 -3369 1304 -3335
rect 1270 -3471 1304 -3437
rect 1534 -3369 1568 -3335
rect 1534 -3471 1568 -3437
rect 1730 -3369 1764 -3335
rect 1730 -3471 1764 -3437
rect 2362 -3369 2396 -3335
rect 2362 -3471 2396 -3437
rect 2558 -3369 2592 -3335
rect 2558 -3471 2592 -3437
rect 2822 -3369 2856 -3335
rect 2822 -3471 2856 -3437
rect 3033 -3377 3067 -3343
rect 3033 -3445 3067 -3411
rect 3131 -3376 3165 -3342
rect 3131 -3444 3165 -3410
rect 3287 -3377 3321 -3343
rect 3287 -3445 3321 -3411
rect 3391 -3376 3425 -3342
rect 3391 -3444 3425 -3410
rect 3549 -3376 3583 -3342
rect 3549 -3444 3583 -3410
rect 3649 -3376 3683 -3342
rect 3649 -3444 3683 -3410
rect 3846 -3369 3880 -3335
rect 3846 -3471 3880 -3437
rect 4110 -3369 4144 -3335
rect 4110 -3471 4144 -3437
rect 4306 -3369 4340 -3335
rect 4306 -3471 4340 -3437
rect 4938 -3369 4972 -3335
rect 4938 -3471 4972 -3437
rect 5134 -3369 5168 -3335
rect 5134 -3471 5168 -3437
rect 5398 -3369 5432 -3335
rect 5398 -3471 5432 -3437
rect 5609 -3377 5643 -3343
rect 5609 -3445 5643 -3411
rect 5707 -3376 5741 -3342
rect 5707 -3444 5741 -3410
rect 5863 -3377 5897 -3343
rect 5863 -3445 5897 -3411
rect 5967 -3376 6001 -3342
rect 5967 -3444 6001 -3410
rect 6125 -3376 6159 -3342
rect 6125 -3444 6159 -3410
rect 6225 -3376 6259 -3342
rect 6225 -3444 6259 -3410
rect 6422 -3369 6456 -3335
rect 6422 -3471 6456 -3437
rect 6686 -3369 6720 -3335
rect 6686 -3471 6720 -3437
rect 6882 -3369 6916 -3335
rect 6882 -3471 6916 -3437
rect 7514 -3369 7548 -3335
rect 7514 -3471 7548 -3437
rect 7710 -3369 7744 -3335
rect 7710 -3471 7744 -3437
rect 7974 -3369 8008 -3335
rect 7974 -3471 8008 -3437
rect 8185 -3377 8219 -3343
rect 8185 -3445 8219 -3411
rect 8283 -3376 8317 -3342
rect 8283 -3444 8317 -3410
rect 8439 -3377 8473 -3343
rect 8439 -3445 8473 -3411
rect 8543 -3376 8577 -3342
rect 8543 -3444 8577 -3410
rect 8701 -3376 8735 -3342
rect 8701 -3444 8735 -3410
rect 8801 -3376 8835 -3342
rect 8801 -3444 8835 -3410
rect 8998 -3369 9032 -3335
rect 8998 -3471 9032 -3437
rect 9262 -3369 9296 -3335
rect 9262 -3471 9296 -3437
rect 9458 -3369 9492 -3335
rect 9458 -3471 9492 -3437
rect 10090 -3369 10124 -3335
rect 10090 -3471 10124 -3437
rect 10378 -3369 10412 -3335
rect 10378 -3471 10412 -3437
rect 10642 -3369 10676 -3335
rect 10642 -3471 10676 -3437
rect 10761 -3377 10795 -3343
rect 10761 -3445 10795 -3411
rect 10859 -3376 10893 -3342
rect 10859 -3444 10893 -3410
rect 11015 -3377 11049 -3343
rect 11015 -3445 11049 -3411
rect 11119 -3376 11153 -3342
rect 11119 -3444 11153 -3410
rect 11277 -3376 11311 -3342
rect 11277 -3444 11311 -3410
rect 11377 -3376 11411 -3342
rect 11377 -3444 11411 -3410
rect 11666 -3369 11700 -3335
rect 11666 -3471 11700 -3437
rect 11930 -3369 11964 -3335
rect 11930 -3471 11964 -3437
rect 13598 -3369 13632 -3335
rect 13598 -3471 13632 -3437
rect 14598 -3369 14632 -3335
rect 14598 -3471 14632 -3437
rect 14794 -3369 14828 -3335
rect 14794 -3471 14828 -3437
rect 15794 -3369 15828 -3335
rect 15794 -3471 15828 -3437
rect 15990 -3369 16024 -3335
rect 15990 -3471 16024 -3437
rect 16622 -3369 16656 -3335
rect 16622 -3471 16656 -3437
rect -2962 -4203 -2928 -4169
rect -2962 -4305 -2928 -4271
rect -2330 -4203 -2296 -4169
rect -2330 -4305 -2296 -4271
rect -1582 -4203 -1548 -4169
rect -1582 -4305 -1548 -4271
rect -950 -4203 -916 -4169
rect -950 -4305 -916 -4271
rect -846 -4203 -812 -4169
rect -846 -4305 -812 -4271
rect -214 -4203 -180 -4169
rect -214 -4305 -180 -4271
rect -18 -4203 16 -4169
rect -18 -4305 16 -4271
rect 246 -4203 280 -4169
rect 246 -4305 280 -4271
rect 443 -4230 477 -4196
rect 443 -4298 477 -4264
rect 543 -4230 577 -4196
rect 543 -4298 577 -4264
rect 701 -4230 735 -4196
rect 701 -4298 735 -4264
rect 805 -4229 839 -4195
rect 805 -4297 839 -4263
rect 961 -4230 995 -4196
rect 961 -4298 995 -4264
rect 1059 -4229 1093 -4195
rect 1059 -4297 1093 -4263
rect 1270 -4203 1304 -4169
rect 1270 -4305 1304 -4271
rect 1534 -4203 1568 -4169
rect 1534 -4305 1568 -4271
rect 1730 -4203 1764 -4169
rect 1730 -4305 1764 -4271
rect 2362 -4203 2396 -4169
rect 2362 -4305 2396 -4271
rect 2558 -4203 2592 -4169
rect 2558 -4305 2592 -4271
rect 2822 -4203 2856 -4169
rect 2822 -4305 2856 -4271
rect 3019 -4230 3053 -4196
rect 3019 -4298 3053 -4264
rect 3119 -4230 3153 -4196
rect 3119 -4298 3153 -4264
rect 3277 -4230 3311 -4196
rect 3277 -4298 3311 -4264
rect 3381 -4229 3415 -4195
rect 3381 -4297 3415 -4263
rect 3537 -4230 3571 -4196
rect 3537 -4298 3571 -4264
rect 3635 -4229 3669 -4195
rect 3635 -4297 3669 -4263
rect 3846 -4203 3880 -4169
rect 3846 -4305 3880 -4271
rect 4110 -4203 4144 -4169
rect 4110 -4305 4144 -4271
rect 4306 -4203 4340 -4169
rect 4306 -4305 4340 -4271
rect 4938 -4203 4972 -4169
rect 4938 -4305 4972 -4271
rect 5134 -4203 5168 -4169
rect 5134 -4305 5168 -4271
rect 5398 -4203 5432 -4169
rect 5398 -4305 5432 -4271
rect 5595 -4230 5629 -4196
rect 5595 -4298 5629 -4264
rect 5695 -4230 5729 -4196
rect 5695 -4298 5729 -4264
rect 5853 -4230 5887 -4196
rect 5853 -4298 5887 -4264
rect 5957 -4229 5991 -4195
rect 5957 -4297 5991 -4263
rect 6113 -4230 6147 -4196
rect 6113 -4298 6147 -4264
rect 6211 -4229 6245 -4195
rect 6211 -4297 6245 -4263
rect 6422 -4203 6456 -4169
rect 6422 -4305 6456 -4271
rect 6686 -4203 6720 -4169
rect 6686 -4305 6720 -4271
rect 6882 -4203 6916 -4169
rect 6882 -4305 6916 -4271
rect 7514 -4203 7548 -4169
rect 7514 -4305 7548 -4271
rect 7710 -4203 7744 -4169
rect 7710 -4305 7744 -4271
rect 7974 -4203 8008 -4169
rect 7974 -4305 8008 -4271
rect 8171 -4230 8205 -4196
rect 8171 -4298 8205 -4264
rect 8271 -4230 8305 -4196
rect 8271 -4298 8305 -4264
rect 8429 -4230 8463 -4196
rect 8429 -4298 8463 -4264
rect 8533 -4229 8567 -4195
rect 8533 -4297 8567 -4263
rect 8689 -4230 8723 -4196
rect 8689 -4298 8723 -4264
rect 8787 -4229 8821 -4195
rect 8787 -4297 8821 -4263
rect 8998 -4203 9032 -4169
rect 8998 -4305 9032 -4271
rect 9262 -4203 9296 -4169
rect 9262 -4305 9296 -4271
rect 9458 -4203 9492 -4169
rect 9458 -4305 9492 -4271
rect 10090 -4203 10124 -4169
rect 10090 -4305 10124 -4271
rect 10378 -4203 10412 -4169
rect 10378 -4305 10412 -4271
rect 10642 -4203 10676 -4169
rect 10642 -4305 10676 -4271
rect 10747 -4230 10781 -4196
rect 10747 -4298 10781 -4264
rect 10847 -4230 10881 -4196
rect 10847 -4298 10881 -4264
rect 11005 -4230 11039 -4196
rect 11005 -4298 11039 -4264
rect 11109 -4229 11143 -4195
rect 11109 -4297 11143 -4263
rect 11265 -4230 11299 -4196
rect 11265 -4298 11299 -4264
rect 11363 -4229 11397 -4195
rect 11363 -4297 11397 -4263
rect 11666 -4203 11700 -4169
rect 11666 -4305 11700 -4271
rect 11930 -4203 11964 -4169
rect 11930 -4305 11964 -4271
rect 12502 -4230 12536 -4196
rect 12502 -4298 12536 -4264
rect 12588 -4203 12622 -4169
rect 12588 -4291 12622 -4257
rect 12674 -4230 12708 -4196
rect 12674 -4298 12708 -4264
rect 12760 -4203 12794 -4169
rect 12760 -4291 12794 -4257
rect 12846 -4230 12880 -4196
rect 12846 -4298 12880 -4264
rect 12932 -4203 12966 -4169
rect 12932 -4291 12966 -4257
rect 13018 -4230 13052 -4196
rect 13018 -4298 13052 -4264
rect 13230 -4203 13264 -4169
rect 13230 -4305 13264 -4271
rect 13494 -4203 13528 -4169
rect 13494 -4305 13528 -4271
rect 13690 -4237 13724 -4203
rect 13690 -4305 13724 -4271
rect 13776 -4229 13810 -4195
rect 13776 -4297 13810 -4263
rect 13862 -4237 13896 -4203
rect 13862 -4305 13896 -4271
rect 13948 -4221 13982 -4187
rect 13948 -4289 13982 -4255
rect 14034 -4237 14068 -4203
rect 14034 -4305 14068 -4271
rect 14120 -4175 14154 -4141
rect 14120 -4261 14154 -4227
rect 14206 -4281 14240 -4247
rect 14292 -4175 14326 -4141
rect 14292 -4261 14326 -4227
rect 14378 -4281 14412 -4247
rect 14464 -4175 14498 -4141
rect 14464 -4261 14498 -4227
rect 14550 -4281 14584 -4247
rect 14636 -4175 14670 -4141
rect 14636 -4261 14670 -4227
rect 14722 -4281 14756 -4247
rect 14807 -4175 14841 -4141
rect 14807 -4261 14841 -4227
rect 14893 -4281 14927 -4247
rect 14979 -4175 15013 -4141
rect 14979 -4261 15013 -4227
rect 15065 -4281 15099 -4247
rect 15151 -4175 15185 -4141
rect 15151 -4261 15185 -4227
rect 15237 -4281 15271 -4247
rect 15323 -4175 15357 -4141
rect 15323 -4261 15357 -4227
rect 15409 -4281 15443 -4247
rect 15622 -4203 15656 -4169
rect 15622 -4305 15656 -4271
rect 16622 -4203 16656 -4169
rect 16622 -4305 16656 -4271
rect -2962 -4457 -2928 -4423
rect -2962 -4559 -2928 -4525
rect -2330 -4457 -2296 -4423
rect -2330 -4559 -2296 -4525
rect -1582 -4457 -1548 -4423
rect -1582 -4559 -1548 -4525
rect -950 -4457 -916 -4423
rect -950 -4559 -916 -4525
rect -831 -4465 -797 -4431
rect -831 -4533 -797 -4499
rect -733 -4464 -699 -4430
rect -733 -4532 -699 -4498
rect -577 -4465 -543 -4431
rect -577 -4533 -543 -4499
rect -473 -4464 -439 -4430
rect -473 -4532 -439 -4498
rect -315 -4464 -281 -4430
rect -315 -4532 -281 -4498
rect -215 -4464 -181 -4430
rect -215 -4532 -181 -4498
rect -18 -4457 16 -4423
rect -18 -4559 16 -4525
rect 246 -4457 280 -4423
rect 246 -4559 280 -4525
rect 457 -4465 491 -4431
rect 457 -4533 491 -4499
rect 555 -4464 589 -4430
rect 555 -4532 589 -4498
rect 711 -4465 745 -4431
rect 711 -4533 745 -4499
rect 815 -4464 849 -4430
rect 815 -4532 849 -4498
rect 973 -4464 1007 -4430
rect 973 -4532 1007 -4498
rect 1073 -4464 1107 -4430
rect 1073 -4532 1107 -4498
rect 1270 -4457 1304 -4423
rect 1270 -4559 1304 -4525
rect 1534 -4457 1568 -4423
rect 1534 -4559 1568 -4525
rect 1730 -4457 1764 -4423
rect 1730 -4559 1764 -4525
rect 2362 -4457 2396 -4423
rect 2362 -4559 2396 -4525
rect 2558 -4457 2592 -4423
rect 2558 -4559 2592 -4525
rect 2822 -4457 2856 -4423
rect 2822 -4559 2856 -4525
rect 3033 -4465 3067 -4431
rect 3033 -4533 3067 -4499
rect 3131 -4464 3165 -4430
rect 3131 -4532 3165 -4498
rect 3287 -4465 3321 -4431
rect 3287 -4533 3321 -4499
rect 3391 -4464 3425 -4430
rect 3391 -4532 3425 -4498
rect 3549 -4464 3583 -4430
rect 3549 -4532 3583 -4498
rect 3649 -4464 3683 -4430
rect 3649 -4532 3683 -4498
rect 3846 -4457 3880 -4423
rect 3846 -4559 3880 -4525
rect 4110 -4457 4144 -4423
rect 4110 -4559 4144 -4525
rect 4306 -4457 4340 -4423
rect 4306 -4559 4340 -4525
rect 4938 -4457 4972 -4423
rect 4938 -4559 4972 -4525
rect 5134 -4457 5168 -4423
rect 5134 -4559 5168 -4525
rect 5398 -4457 5432 -4423
rect 5398 -4559 5432 -4525
rect 5609 -4465 5643 -4431
rect 5609 -4533 5643 -4499
rect 5707 -4464 5741 -4430
rect 5707 -4532 5741 -4498
rect 5863 -4465 5897 -4431
rect 5863 -4533 5897 -4499
rect 5967 -4464 6001 -4430
rect 5967 -4532 6001 -4498
rect 6125 -4464 6159 -4430
rect 6125 -4532 6159 -4498
rect 6225 -4464 6259 -4430
rect 6225 -4532 6259 -4498
rect 6422 -4457 6456 -4423
rect 6422 -4559 6456 -4525
rect 6686 -4457 6720 -4423
rect 6686 -4559 6720 -4525
rect 6882 -4457 6916 -4423
rect 6882 -4559 6916 -4525
rect 7514 -4457 7548 -4423
rect 7514 -4559 7548 -4525
rect 7710 -4457 7744 -4423
rect 7710 -4559 7744 -4525
rect 7974 -4457 8008 -4423
rect 7974 -4559 8008 -4525
rect 8185 -4465 8219 -4431
rect 8185 -4533 8219 -4499
rect 8283 -4464 8317 -4430
rect 8283 -4532 8317 -4498
rect 8439 -4465 8473 -4431
rect 8439 -4533 8473 -4499
rect 8543 -4464 8577 -4430
rect 8543 -4532 8577 -4498
rect 8701 -4464 8735 -4430
rect 8701 -4532 8735 -4498
rect 8801 -4464 8835 -4430
rect 8801 -4532 8835 -4498
rect 8998 -4457 9032 -4423
rect 8998 -4559 9032 -4525
rect 9262 -4457 9296 -4423
rect 9262 -4559 9296 -4525
rect 9458 -4457 9492 -4423
rect 9458 -4559 9492 -4525
rect 10090 -4457 10124 -4423
rect 10090 -4559 10124 -4525
rect 10378 -4457 10412 -4423
rect 10378 -4559 10412 -4525
rect 10642 -4457 10676 -4423
rect 10642 -4559 10676 -4525
rect 10761 -4465 10795 -4431
rect 10761 -4533 10795 -4499
rect 10859 -4464 10893 -4430
rect 10859 -4532 10893 -4498
rect 11015 -4465 11049 -4431
rect 11015 -4533 11049 -4499
rect 11119 -4464 11153 -4430
rect 11119 -4532 11153 -4498
rect 11277 -4464 11311 -4430
rect 11277 -4532 11311 -4498
rect 11377 -4464 11411 -4430
rect 11377 -4532 11411 -4498
rect 11666 -4457 11700 -4423
rect 11666 -4559 11700 -4525
rect 11930 -4457 11964 -4423
rect 11930 -4559 11964 -4525
rect 13690 -4457 13724 -4423
rect 13690 -4525 13724 -4491
rect 13776 -4465 13810 -4431
rect 13776 -4533 13810 -4499
rect 13862 -4457 13896 -4423
rect 13862 -4525 13896 -4491
rect 13948 -4473 13982 -4439
rect 13948 -4541 13982 -4507
rect 14034 -4457 14068 -4423
rect 14034 -4525 14068 -4491
rect 14120 -4501 14154 -4467
rect 14120 -4587 14154 -4553
rect 14206 -4481 14240 -4447
rect 14292 -4501 14326 -4467
rect 14292 -4587 14326 -4553
rect 14378 -4481 14412 -4447
rect 14464 -4501 14498 -4467
rect 14464 -4587 14498 -4553
rect 14550 -4481 14584 -4447
rect 14636 -4501 14670 -4467
rect 14636 -4587 14670 -4553
rect 14722 -4481 14756 -4447
rect 14807 -4501 14841 -4467
rect 14807 -4587 14841 -4553
rect 14893 -4481 14927 -4447
rect 14979 -4501 15013 -4467
rect 14979 -4587 15013 -4553
rect 15065 -4481 15099 -4447
rect 15151 -4501 15185 -4467
rect 15151 -4587 15185 -4553
rect 15237 -4481 15271 -4447
rect 15323 -4501 15357 -4467
rect 15323 -4587 15357 -4553
rect 15409 -4481 15443 -4447
rect 15622 -4457 15656 -4423
rect 15622 -4559 15656 -4525
rect 16622 -4457 16656 -4423
rect 16622 -4559 16656 -4525
rect -2962 -5291 -2928 -5257
rect -2962 -5393 -2928 -5359
rect -2330 -5291 -2296 -5257
rect -2330 -5393 -2296 -5359
rect -1582 -5291 -1548 -5257
rect -1582 -5393 -1548 -5359
rect -950 -5291 -916 -5257
rect -950 -5393 -916 -5359
rect -846 -5291 -812 -5257
rect -846 -5393 -812 -5359
rect -214 -5291 -180 -5257
rect -214 -5393 -180 -5359
rect -18 -5291 16 -5257
rect -18 -5393 16 -5359
rect 246 -5291 280 -5257
rect 246 -5393 280 -5359
rect 443 -5318 477 -5284
rect 443 -5386 477 -5352
rect 543 -5318 577 -5284
rect 543 -5386 577 -5352
rect 701 -5318 735 -5284
rect 701 -5386 735 -5352
rect 805 -5317 839 -5283
rect 805 -5385 839 -5351
rect 961 -5318 995 -5284
rect 961 -5386 995 -5352
rect 1059 -5317 1093 -5283
rect 1059 -5385 1093 -5351
rect 1270 -5291 1304 -5257
rect 1270 -5393 1304 -5359
rect 1534 -5291 1568 -5257
rect 1534 -5393 1568 -5359
rect 1730 -5291 1764 -5257
rect 1730 -5393 1764 -5359
rect 2362 -5291 2396 -5257
rect 2362 -5393 2396 -5359
rect 2558 -5291 2592 -5257
rect 2558 -5393 2592 -5359
rect 2822 -5291 2856 -5257
rect 2822 -5393 2856 -5359
rect 3019 -5318 3053 -5284
rect 3019 -5386 3053 -5352
rect 3119 -5318 3153 -5284
rect 3119 -5386 3153 -5352
rect 3277 -5318 3311 -5284
rect 3277 -5386 3311 -5352
rect 3381 -5317 3415 -5283
rect 3381 -5385 3415 -5351
rect 3537 -5318 3571 -5284
rect 3537 -5386 3571 -5352
rect 3635 -5317 3669 -5283
rect 3635 -5385 3669 -5351
rect 3846 -5291 3880 -5257
rect 3846 -5393 3880 -5359
rect 4110 -5291 4144 -5257
rect 4110 -5393 4144 -5359
rect 4306 -5291 4340 -5257
rect 4306 -5393 4340 -5359
rect 4938 -5291 4972 -5257
rect 4938 -5393 4972 -5359
rect 5134 -5291 5168 -5257
rect 5134 -5393 5168 -5359
rect 5398 -5291 5432 -5257
rect 5398 -5393 5432 -5359
rect 5595 -5318 5629 -5284
rect 5595 -5386 5629 -5352
rect 5695 -5318 5729 -5284
rect 5695 -5386 5729 -5352
rect 5853 -5318 5887 -5284
rect 5853 -5386 5887 -5352
rect 5957 -5317 5991 -5283
rect 5957 -5385 5991 -5351
rect 6113 -5318 6147 -5284
rect 6113 -5386 6147 -5352
rect 6211 -5317 6245 -5283
rect 6211 -5385 6245 -5351
rect 6422 -5291 6456 -5257
rect 6422 -5393 6456 -5359
rect 6686 -5291 6720 -5257
rect 6686 -5393 6720 -5359
rect 6882 -5291 6916 -5257
rect 6882 -5393 6916 -5359
rect 7514 -5291 7548 -5257
rect 7514 -5393 7548 -5359
rect 7710 -5291 7744 -5257
rect 7710 -5393 7744 -5359
rect 7974 -5291 8008 -5257
rect 7974 -5393 8008 -5359
rect 8171 -5318 8205 -5284
rect 8171 -5386 8205 -5352
rect 8271 -5318 8305 -5284
rect 8271 -5386 8305 -5352
rect 8429 -5318 8463 -5284
rect 8429 -5386 8463 -5352
rect 8533 -5317 8567 -5283
rect 8533 -5385 8567 -5351
rect 8689 -5318 8723 -5284
rect 8689 -5386 8723 -5352
rect 8787 -5317 8821 -5283
rect 8787 -5385 8821 -5351
rect 8998 -5291 9032 -5257
rect 8998 -5393 9032 -5359
rect 9262 -5291 9296 -5257
rect 9262 -5393 9296 -5359
rect 9458 -5291 9492 -5257
rect 9458 -5393 9492 -5359
rect 10090 -5291 10124 -5257
rect 10090 -5393 10124 -5359
rect 10378 -5291 10412 -5257
rect 10378 -5393 10412 -5359
rect 10642 -5291 10676 -5257
rect 10642 -5393 10676 -5359
rect 10747 -5318 10781 -5284
rect 10747 -5386 10781 -5352
rect 10847 -5318 10881 -5284
rect 10847 -5386 10881 -5352
rect 11005 -5318 11039 -5284
rect 11005 -5386 11039 -5352
rect 11109 -5317 11143 -5283
rect 11109 -5385 11143 -5351
rect 11265 -5318 11299 -5284
rect 11265 -5386 11299 -5352
rect 11363 -5317 11397 -5283
rect 11363 -5385 11397 -5351
rect 11666 -5291 11700 -5257
rect 11666 -5393 11700 -5359
rect 11930 -5291 11964 -5257
rect 11930 -5393 11964 -5359
rect 12502 -5318 12536 -5284
rect 12502 -5386 12536 -5352
rect 12588 -5291 12622 -5257
rect 12588 -5379 12622 -5345
rect 12674 -5318 12708 -5284
rect 12674 -5386 12708 -5352
rect 12760 -5291 12794 -5257
rect 12760 -5379 12794 -5345
rect 12846 -5318 12880 -5284
rect 12846 -5386 12880 -5352
rect 12932 -5291 12966 -5257
rect 12932 -5379 12966 -5345
rect 13018 -5318 13052 -5284
rect 13018 -5386 13052 -5352
rect 13230 -5291 13264 -5257
rect 13230 -5393 13264 -5359
rect 13494 -5291 13528 -5257
rect 13494 -5393 13528 -5359
rect 13690 -5325 13724 -5291
rect 13690 -5393 13724 -5359
rect 13776 -5317 13810 -5283
rect 13776 -5385 13810 -5351
rect 13862 -5325 13896 -5291
rect 13862 -5393 13896 -5359
rect 13948 -5309 13982 -5275
rect 13948 -5377 13982 -5343
rect 14034 -5325 14068 -5291
rect 14034 -5393 14068 -5359
rect 14120 -5263 14154 -5229
rect 14120 -5349 14154 -5315
rect 14206 -5369 14240 -5335
rect 14292 -5263 14326 -5229
rect 14292 -5349 14326 -5315
rect 14378 -5369 14412 -5335
rect 14464 -5263 14498 -5229
rect 14464 -5349 14498 -5315
rect 14550 -5369 14584 -5335
rect 14636 -5263 14670 -5229
rect 14636 -5349 14670 -5315
rect 14722 -5369 14756 -5335
rect 14807 -5263 14841 -5229
rect 14807 -5349 14841 -5315
rect 14893 -5369 14927 -5335
rect 14979 -5263 15013 -5229
rect 14979 -5349 15013 -5315
rect 15065 -5369 15099 -5335
rect 15151 -5263 15185 -5229
rect 15151 -5349 15185 -5315
rect 15237 -5369 15271 -5335
rect 15323 -5263 15357 -5229
rect 15323 -5349 15357 -5315
rect 15409 -5369 15443 -5335
rect 15622 -5291 15656 -5257
rect 15622 -5393 15656 -5359
rect 16622 -5291 16656 -5257
rect 16622 -5393 16656 -5359
rect -2962 -5545 -2928 -5511
rect -2962 -5647 -2928 -5613
rect -2330 -5545 -2296 -5511
rect -2330 -5647 -2296 -5613
rect -1582 -5545 -1548 -5511
rect -1582 -5647 -1548 -5613
rect -950 -5545 -916 -5511
rect -950 -5647 -916 -5613
rect -846 -5545 -812 -5511
rect -846 -5647 -812 -5613
rect -214 -5545 -180 -5511
rect -214 -5647 -180 -5613
rect -18 -5545 16 -5511
rect -18 -5647 16 -5613
rect 246 -5545 280 -5511
rect 246 -5647 280 -5613
rect 457 -5553 491 -5519
rect 457 -5621 491 -5587
rect 555 -5552 589 -5518
rect 555 -5620 589 -5586
rect 711 -5553 745 -5519
rect 711 -5621 745 -5587
rect 815 -5552 849 -5518
rect 815 -5620 849 -5586
rect 973 -5552 1007 -5518
rect 973 -5620 1007 -5586
rect 1073 -5552 1107 -5518
rect 1073 -5620 1107 -5586
rect 1270 -5545 1304 -5511
rect 1270 -5647 1304 -5613
rect 1534 -5545 1568 -5511
rect 1534 -5647 1568 -5613
rect 1730 -5545 1764 -5511
rect 1730 -5647 1764 -5613
rect 2362 -5545 2396 -5511
rect 2362 -5647 2396 -5613
rect 2558 -5545 2592 -5511
rect 2558 -5647 2592 -5613
rect 2822 -5545 2856 -5511
rect 2822 -5647 2856 -5613
rect 3033 -5553 3067 -5519
rect 3033 -5621 3067 -5587
rect 3131 -5552 3165 -5518
rect 3131 -5620 3165 -5586
rect 3287 -5553 3321 -5519
rect 3287 -5621 3321 -5587
rect 3391 -5552 3425 -5518
rect 3391 -5620 3425 -5586
rect 3549 -5552 3583 -5518
rect 3549 -5620 3583 -5586
rect 3649 -5552 3683 -5518
rect 3649 -5620 3683 -5586
rect 3846 -5545 3880 -5511
rect 3846 -5647 3880 -5613
rect 4110 -5545 4144 -5511
rect 4110 -5647 4144 -5613
rect 4306 -5545 4340 -5511
rect 4306 -5647 4340 -5613
rect 4938 -5545 4972 -5511
rect 4938 -5647 4972 -5613
rect 5134 -5545 5168 -5511
rect 5134 -5647 5168 -5613
rect 5398 -5545 5432 -5511
rect 5398 -5647 5432 -5613
rect 5609 -5553 5643 -5519
rect 5609 -5621 5643 -5587
rect 5707 -5552 5741 -5518
rect 5707 -5620 5741 -5586
rect 5863 -5553 5897 -5519
rect 5863 -5621 5897 -5587
rect 5967 -5552 6001 -5518
rect 5967 -5620 6001 -5586
rect 6125 -5552 6159 -5518
rect 6125 -5620 6159 -5586
rect 6225 -5552 6259 -5518
rect 6225 -5620 6259 -5586
rect 6422 -5545 6456 -5511
rect 6422 -5647 6456 -5613
rect 6686 -5545 6720 -5511
rect 6686 -5647 6720 -5613
rect 6882 -5545 6916 -5511
rect 6882 -5647 6916 -5613
rect 7514 -5545 7548 -5511
rect 7514 -5647 7548 -5613
rect 7710 -5545 7744 -5511
rect 7710 -5647 7744 -5613
rect 7974 -5545 8008 -5511
rect 7974 -5647 8008 -5613
rect 8185 -5553 8219 -5519
rect 8185 -5621 8219 -5587
rect 8283 -5552 8317 -5518
rect 8283 -5620 8317 -5586
rect 8439 -5553 8473 -5519
rect 8439 -5621 8473 -5587
rect 8543 -5552 8577 -5518
rect 8543 -5620 8577 -5586
rect 8701 -5552 8735 -5518
rect 8701 -5620 8735 -5586
rect 8801 -5552 8835 -5518
rect 8801 -5620 8835 -5586
rect 8998 -5545 9032 -5511
rect 8998 -5647 9032 -5613
rect 9262 -5545 9296 -5511
rect 9262 -5647 9296 -5613
rect 9458 -5545 9492 -5511
rect 9458 -5647 9492 -5613
rect 10090 -5545 10124 -5511
rect 10090 -5647 10124 -5613
rect 10378 -5545 10412 -5511
rect 10378 -5647 10412 -5613
rect 10642 -5545 10676 -5511
rect 10642 -5647 10676 -5613
rect 10761 -5553 10795 -5519
rect 10761 -5621 10795 -5587
rect 10859 -5552 10893 -5518
rect 10859 -5620 10893 -5586
rect 11015 -5553 11049 -5519
rect 11015 -5621 11049 -5587
rect 11119 -5552 11153 -5518
rect 11119 -5620 11153 -5586
rect 11277 -5552 11311 -5518
rect 11277 -5620 11311 -5586
rect 11377 -5552 11411 -5518
rect 11377 -5620 11411 -5586
rect 11666 -5545 11700 -5511
rect 11666 -5647 11700 -5613
rect 11930 -5545 11964 -5511
rect 11930 -5647 11964 -5613
rect 13690 -5545 13724 -5511
rect 13690 -5613 13724 -5579
rect 13776 -5553 13810 -5519
rect 13776 -5621 13810 -5587
rect 13862 -5545 13896 -5511
rect 13862 -5613 13896 -5579
rect 13948 -5561 13982 -5527
rect 13948 -5629 13982 -5595
rect 14034 -5545 14068 -5511
rect 14034 -5613 14068 -5579
rect 14120 -5589 14154 -5555
rect 14120 -5675 14154 -5641
rect 14206 -5569 14240 -5535
rect 14292 -5589 14326 -5555
rect 14292 -5675 14326 -5641
rect 14378 -5569 14412 -5535
rect 14464 -5589 14498 -5555
rect 14464 -5675 14498 -5641
rect 14550 -5569 14584 -5535
rect 14636 -5589 14670 -5555
rect 14636 -5675 14670 -5641
rect 14722 -5569 14756 -5535
rect 14807 -5589 14841 -5555
rect 14807 -5675 14841 -5641
rect 14893 -5569 14927 -5535
rect 14979 -5589 15013 -5555
rect 14979 -5675 15013 -5641
rect 15065 -5569 15099 -5535
rect 15151 -5589 15185 -5555
rect 15151 -5675 15185 -5641
rect 15237 -5569 15271 -5535
rect 15323 -5589 15357 -5555
rect 15323 -5675 15357 -5641
rect 15409 -5569 15443 -5535
rect 15622 -5545 15656 -5511
rect 15622 -5647 15656 -5613
rect 16622 -5545 16656 -5511
rect 16622 -5647 16656 -5613
rect -2962 -6379 -2928 -6345
rect -2962 -6481 -2928 -6447
rect -2330 -6379 -2296 -6345
rect -2330 -6481 -2296 -6447
rect -1398 -6379 -1364 -6345
rect -1398 -6481 -1364 -6447
rect -1134 -6379 -1100 -6345
rect -1134 -6481 -1100 -6447
rect -934 -6345 -900 -6311
rect -934 -6413 -900 -6379
rect -934 -6481 -900 -6447
rect -850 -6345 -816 -6311
rect -850 -6413 -816 -6379
rect -850 -6481 -816 -6447
rect -766 -6345 -732 -6311
rect -766 -6413 -732 -6379
rect -766 -6481 -732 -6447
rect -570 -6379 -536 -6345
rect -570 -6481 -536 -6447
rect -306 -6379 -272 -6345
rect -306 -6481 -272 -6447
rect -102 -6406 -68 -6372
rect -102 -6474 -68 -6440
rect -16 -6379 18 -6345
rect -16 -6467 18 -6433
rect 70 -6406 104 -6372
rect 70 -6474 104 -6440
rect 156 -6379 190 -6345
rect 156 -6467 190 -6433
rect 242 -6406 276 -6372
rect 242 -6474 276 -6440
rect 328 -6379 362 -6345
rect 328 -6467 362 -6433
rect 414 -6406 448 -6372
rect 414 -6474 448 -6440
rect 626 -6379 660 -6345
rect 626 -6481 660 -6447
rect 890 -6379 924 -6345
rect 890 -6481 924 -6447
rect 1086 -6379 1120 -6345
rect 1086 -6481 1120 -6447
rect 1170 -6379 1204 -6345
rect 1170 -6481 1204 -6447
rect 1254 -6379 1288 -6345
rect 1254 -6481 1288 -6447
rect 1454 -6379 1488 -6345
rect 1454 -6481 1488 -6447
rect 1718 -6379 1752 -6345
rect 1718 -6481 1752 -6447
rect 1914 -6379 1948 -6345
rect 1914 -6481 1948 -6447
rect 2178 -6379 2212 -6345
rect 2178 -6481 2212 -6447
rect 2375 -6406 2409 -6372
rect 2375 -6474 2409 -6440
rect 2475 -6406 2509 -6372
rect 2475 -6474 2509 -6440
rect 2633 -6406 2667 -6372
rect 2633 -6474 2667 -6440
rect 2737 -6405 2771 -6371
rect 2737 -6473 2771 -6439
rect 2893 -6406 2927 -6372
rect 2893 -6474 2927 -6440
rect 2991 -6405 3025 -6371
rect 2991 -6473 3025 -6439
rect 3202 -6379 3236 -6345
rect 3202 -6481 3236 -6447
rect 3466 -6379 3500 -6345
rect 3466 -6481 3500 -6447
rect 4398 -6379 4432 -6345
rect 4398 -6481 4432 -6447
rect 5398 -6379 5432 -6345
rect 5398 -6481 5432 -6447
rect 6422 -6379 6456 -6345
rect 6422 -6481 6456 -6447
rect 6686 -6379 6720 -6345
rect 6686 -6481 6720 -6447
rect 6883 -6406 6917 -6372
rect 6883 -6474 6917 -6440
rect 6983 -6406 7017 -6372
rect 6983 -6474 7017 -6440
rect 7141 -6406 7175 -6372
rect 7141 -6474 7175 -6440
rect 7245 -6405 7279 -6371
rect 7245 -6473 7279 -6439
rect 7401 -6406 7435 -6372
rect 7401 -6474 7435 -6440
rect 7499 -6405 7533 -6371
rect 7499 -6473 7533 -6439
rect 7710 -6379 7744 -6345
rect 7710 -6481 7744 -6447
rect 7974 -6379 8008 -6345
rect 7974 -6481 8008 -6447
rect 8171 -6406 8205 -6372
rect 8171 -6474 8205 -6440
rect 8271 -6406 8305 -6372
rect 8271 -6474 8305 -6440
rect 8429 -6406 8463 -6372
rect 8429 -6474 8463 -6440
rect 8533 -6405 8567 -6371
rect 8533 -6473 8567 -6439
rect 8689 -6406 8723 -6372
rect 8689 -6474 8723 -6440
rect 8787 -6405 8821 -6371
rect 8787 -6473 8821 -6439
rect 8998 -6379 9032 -6345
rect 8998 -6481 9032 -6447
rect 9262 -6379 9296 -6345
rect 9262 -6481 9296 -6447
rect 9459 -6406 9493 -6372
rect 9459 -6474 9493 -6440
rect 9559 -6406 9593 -6372
rect 9559 -6474 9593 -6440
rect 9717 -6406 9751 -6372
rect 9717 -6474 9751 -6440
rect 9821 -6405 9855 -6371
rect 9821 -6473 9855 -6439
rect 9977 -6406 10011 -6372
rect 9977 -6474 10011 -6440
rect 10075 -6405 10109 -6371
rect 10075 -6473 10109 -6439
rect 10286 -6379 10320 -6345
rect 10286 -6481 10320 -6447
rect 10550 -6379 10584 -6345
rect 10550 -6481 10584 -6447
rect 10746 -6345 10780 -6311
rect 10746 -6413 10780 -6379
rect 10746 -6481 10780 -6447
rect 10830 -6345 10864 -6311
rect 10830 -6413 10864 -6379
rect 10830 -6481 10864 -6447
rect 10914 -6413 10948 -6379
rect 10914 -6481 10948 -6447
rect 10998 -6345 11032 -6311
rect 10998 -6413 11032 -6379
rect 10998 -6481 11032 -6447
rect 11082 -6413 11116 -6379
rect 11082 -6481 11116 -6447
rect 11166 -6345 11200 -6311
rect 11166 -6413 11200 -6379
rect 11166 -6481 11200 -6447
rect 11250 -6413 11284 -6379
rect 11250 -6481 11284 -6447
rect 11334 -6345 11368 -6311
rect 11334 -6413 11368 -6379
rect 11334 -6481 11368 -6447
rect 11418 -6413 11452 -6379
rect 11418 -6481 11452 -6447
rect 11666 -6379 11700 -6345
rect 11666 -6481 11700 -6447
rect 11930 -6379 11964 -6345
rect 11930 -6481 11964 -6447
rect 13598 -6379 13632 -6345
rect 13598 -6481 13632 -6447
rect 14598 -6379 14632 -6345
rect 14598 -6481 14632 -6447
rect 14794 -6379 14828 -6345
rect 14794 -6481 14828 -6447
rect 15794 -6379 15828 -6345
rect 15794 -6481 15828 -6447
rect 15990 -6379 16024 -6345
rect 15990 -6481 16024 -6447
rect 16622 -6379 16656 -6345
rect 16622 -6481 16656 -6447
rect -2962 -6633 -2928 -6599
rect -2962 -6728 -2928 -6694
rect -2790 -6633 -2756 -6599
rect -2790 -6728 -2756 -6694
rect -2594 -6641 -2560 -6607
rect -2594 -6709 -2560 -6675
rect -2510 -6657 -2476 -6623
rect -2426 -6641 -2392 -6607
rect -2322 -6633 -2288 -6599
rect -2238 -6641 -2204 -6607
rect -2146 -6646 -2112 -6612
rect -1907 -6633 -1873 -6599
rect -2426 -6709 -2392 -6675
rect -1907 -6701 -1873 -6667
rect -1823 -6641 -1789 -6607
rect -1728 -6651 -1694 -6617
rect -1529 -6641 -1495 -6607
rect -1405 -6633 -1371 -6599
rect -1405 -6704 -1371 -6670
rect -1405 -6775 -1371 -6741
rect -1319 -6663 -1285 -6629
rect -1319 -6743 -1285 -6709
rect -1235 -6639 -1201 -6605
rect -1235 -6707 -1201 -6673
rect -1131 -6633 -1097 -6599
rect -1131 -6701 -1097 -6667
rect -1034 -6633 -1000 -6599
rect -1034 -6701 -1000 -6667
rect -1235 -6775 -1201 -6741
rect -1034 -6769 -1000 -6735
rect -950 -6633 -916 -6599
rect -950 -6704 -916 -6670
rect -950 -6775 -916 -6741
rect -846 -6633 -812 -6599
rect -846 -6735 -812 -6701
rect -214 -6633 -180 -6599
rect -214 -6735 -180 -6701
rect -18 -6633 16 -6599
rect -18 -6735 16 -6701
rect 614 -6633 648 -6599
rect 614 -6735 648 -6701
rect 718 -6633 752 -6599
rect 718 -6735 752 -6701
rect 1350 -6633 1384 -6599
rect 1350 -6735 1384 -6701
rect 1546 -6633 1580 -6599
rect 1546 -6735 1580 -6701
rect 2178 -6633 2212 -6599
rect 2178 -6735 2212 -6701
rect 2282 -6633 2316 -6599
rect 2282 -6735 2316 -6701
rect 2914 -6633 2948 -6599
rect 2914 -6735 2948 -6701
rect 3110 -6633 3144 -6599
rect 3110 -6735 3144 -6701
rect 3742 -6633 3776 -6599
rect 3742 -6735 3776 -6701
rect 3846 -6633 3880 -6599
rect 3846 -6735 3880 -6701
rect 4478 -6633 4512 -6599
rect 4478 -6735 4512 -6701
rect 4674 -6633 4708 -6599
rect 4674 -6735 4708 -6701
rect 5306 -6633 5340 -6599
rect 5306 -6735 5340 -6701
rect 5410 -6633 5444 -6599
rect 5410 -6735 5444 -6701
rect 6042 -6633 6076 -6599
rect 6042 -6735 6076 -6701
rect 6238 -6633 6272 -6599
rect 6238 -6735 6272 -6701
rect 6870 -6633 6904 -6599
rect 6870 -6735 6904 -6701
rect 6974 -6633 7008 -6599
rect 6974 -6735 7008 -6701
rect 7606 -6633 7640 -6599
rect 7606 -6735 7640 -6701
rect 7802 -6633 7836 -6599
rect 7802 -6735 7836 -6701
rect 8434 -6633 8468 -6599
rect 8434 -6735 8468 -6701
rect 8538 -6633 8572 -6599
rect 8538 -6735 8572 -6701
rect 9170 -6633 9204 -6599
rect 9170 -6735 9204 -6701
rect 15990 -6633 16024 -6599
rect 15990 -6735 16024 -6701
rect 16622 -6633 16656 -6599
rect 16622 -6735 16656 -6701
rect -2962 -7467 -2928 -7433
rect -2962 -7569 -2928 -7535
rect -2330 -7467 -2296 -7433
rect -2330 -7569 -2296 -7535
rect -1582 -7467 -1548 -7433
rect -1582 -7569 -1548 -7535
rect -950 -7467 -916 -7433
rect -950 -7569 -916 -7535
rect -846 -7467 -812 -7433
rect -846 -7569 -812 -7535
rect -214 -7467 -180 -7433
rect -214 -7569 -180 -7535
rect -18 -7467 16 -7433
rect -18 -7569 16 -7535
rect 614 -7467 648 -7433
rect 614 -7569 648 -7535
rect 718 -7467 752 -7433
rect 718 -7569 752 -7535
rect 1350 -7467 1384 -7433
rect 1350 -7569 1384 -7535
rect 1546 -7467 1580 -7433
rect 1546 -7569 1580 -7535
rect 2178 -7467 2212 -7433
rect 2178 -7569 2212 -7535
rect 2282 -7467 2316 -7433
rect 2282 -7569 2316 -7535
rect 2546 -7467 2580 -7433
rect 2546 -7569 2580 -7535
rect 2930 -7467 2964 -7433
rect 2930 -7569 2964 -7535
rect 3014 -7467 3048 -7433
rect 3014 -7569 3048 -7535
rect 3098 -7467 3132 -7433
rect 3098 -7569 3132 -7535
rect 3294 -7467 3328 -7433
rect 3294 -7569 3328 -7535
rect 3558 -7467 3592 -7433
rect 3558 -7569 3592 -7535
rect 3758 -7433 3792 -7399
rect 3758 -7501 3792 -7467
rect 3758 -7569 3792 -7535
rect 3842 -7433 3876 -7399
rect 3842 -7501 3876 -7467
rect 3842 -7569 3876 -7535
rect 3926 -7433 3960 -7399
rect 3926 -7501 3960 -7467
rect 3926 -7569 3960 -7535
rect 4122 -7467 4156 -7433
rect 4122 -7569 4156 -7535
rect 4386 -7467 4420 -7433
rect 4386 -7569 4420 -7535
rect 4582 -7433 4616 -7399
rect 4582 -7501 4616 -7467
rect 4582 -7569 4616 -7535
rect 4666 -7433 4700 -7399
rect 4666 -7501 4700 -7467
rect 4666 -7569 4700 -7535
rect 4902 -7509 4936 -7475
rect 4977 -7509 5011 -7475
rect 5174 -7509 5208 -7475
rect 5260 -7509 5294 -7475
rect 5502 -7467 5536 -7433
rect 5502 -7569 5536 -7535
rect 5766 -7467 5800 -7433
rect 5766 -7569 5800 -7535
rect 5962 -7427 5996 -7393
rect 5962 -7498 5996 -7464
rect 5962 -7569 5996 -7535
rect 6046 -7433 6080 -7399
rect 6247 -7427 6281 -7393
rect 6046 -7501 6080 -7467
rect 6046 -7569 6080 -7535
rect 6143 -7501 6177 -7467
rect 6143 -7569 6177 -7535
rect 6247 -7495 6281 -7461
rect 6247 -7563 6281 -7529
rect 6331 -7459 6365 -7425
rect 6331 -7539 6365 -7505
rect 6417 -7427 6451 -7393
rect 6417 -7498 6451 -7464
rect 6417 -7569 6451 -7535
rect 6541 -7561 6575 -7527
rect 6740 -7551 6774 -7517
rect 6835 -7561 6869 -7527
rect 6919 -7501 6953 -7467
rect 7438 -7493 7472 -7459
rect 6919 -7569 6953 -7535
rect 7158 -7556 7192 -7522
rect 7250 -7561 7284 -7527
rect 7334 -7569 7368 -7535
rect 7438 -7561 7472 -7527
rect 7522 -7545 7556 -7511
rect 7606 -7493 7640 -7459
rect 7606 -7561 7640 -7527
rect 7802 -7467 7836 -7433
rect 7802 -7569 7836 -7535
rect 8434 -7467 8468 -7433
rect 8434 -7569 8468 -7535
rect 8538 -7467 8572 -7433
rect 8538 -7569 8572 -7535
rect 9170 -7467 9204 -7433
rect 9170 -7569 9204 -7535
rect 15990 -7467 16024 -7433
rect 15990 -7569 16024 -7535
rect 16622 -7467 16656 -7433
rect 16622 -7569 16656 -7535
rect -2962 -7721 -2928 -7687
rect -2962 -7823 -2928 -7789
rect -2330 -7721 -2296 -7687
rect -2330 -7823 -2296 -7789
rect -1398 -7721 -1364 -7687
rect -1398 -7823 -1364 -7789
rect -1134 -7721 -1100 -7687
rect -1134 -7823 -1100 -7789
rect -934 -7721 -900 -7687
rect -934 -7789 -900 -7755
rect -934 -7857 -900 -7823
rect -850 -7721 -816 -7687
rect -850 -7789 -816 -7755
rect -850 -7857 -816 -7823
rect -766 -7721 -732 -7687
rect -766 -7789 -732 -7755
rect -766 -7857 -732 -7823
rect -570 -7721 -536 -7687
rect -570 -7823 -536 -7789
rect -306 -7721 -272 -7687
rect -306 -7823 -272 -7789
rect -102 -7728 -68 -7694
rect -102 -7796 -68 -7762
rect -16 -7735 18 -7701
rect -16 -7823 18 -7789
rect 70 -7728 104 -7694
rect 70 -7796 104 -7762
rect 156 -7735 190 -7701
rect 156 -7823 190 -7789
rect 242 -7728 276 -7694
rect 242 -7796 276 -7762
rect 328 -7735 362 -7701
rect 328 -7823 362 -7789
rect 414 -7728 448 -7694
rect 414 -7796 448 -7762
rect 626 -7721 660 -7687
rect 626 -7823 660 -7789
rect 890 -7721 924 -7687
rect 890 -7823 924 -7789
rect 1086 -7721 1120 -7687
rect 1086 -7823 1120 -7789
rect 1170 -7721 1204 -7687
rect 1170 -7823 1204 -7789
rect 1254 -7721 1288 -7687
rect 1254 -7823 1288 -7789
rect 1454 -7721 1488 -7687
rect 1454 -7823 1488 -7789
rect 1718 -7721 1752 -7687
rect 1718 -7823 1752 -7789
rect 1914 -7721 1948 -7687
rect 1914 -7823 1948 -7789
rect 2178 -7721 2212 -7687
rect 2178 -7823 2212 -7789
rect 2375 -7728 2409 -7694
rect 2375 -7796 2409 -7762
rect 2475 -7728 2509 -7694
rect 2475 -7796 2509 -7762
rect 2633 -7728 2667 -7694
rect 2633 -7796 2667 -7762
rect 2737 -7729 2771 -7695
rect 2737 -7797 2771 -7763
rect 2893 -7728 2927 -7694
rect 2893 -7796 2927 -7762
rect 2991 -7729 3025 -7695
rect 2991 -7797 3025 -7763
rect 3202 -7721 3236 -7687
rect 3202 -7823 3236 -7789
rect 3466 -7721 3500 -7687
rect 3466 -7823 3500 -7789
rect 4398 -7721 4432 -7687
rect 4398 -7823 4432 -7789
rect 5398 -7721 5432 -7687
rect 5398 -7823 5432 -7789
rect 6422 -7721 6456 -7687
rect 6422 -7823 6456 -7789
rect 6686 -7721 6720 -7687
rect 6686 -7823 6720 -7789
rect 6883 -7728 6917 -7694
rect 6883 -7796 6917 -7762
rect 6983 -7728 7017 -7694
rect 6983 -7796 7017 -7762
rect 7141 -7728 7175 -7694
rect 7141 -7796 7175 -7762
rect 7245 -7729 7279 -7695
rect 7245 -7797 7279 -7763
rect 7401 -7728 7435 -7694
rect 7401 -7796 7435 -7762
rect 7499 -7729 7533 -7695
rect 7499 -7797 7533 -7763
rect 7710 -7721 7744 -7687
rect 7710 -7823 7744 -7789
rect 7974 -7721 8008 -7687
rect 7974 -7823 8008 -7789
rect 8171 -7728 8205 -7694
rect 8171 -7796 8205 -7762
rect 8271 -7728 8305 -7694
rect 8271 -7796 8305 -7762
rect 8429 -7728 8463 -7694
rect 8429 -7796 8463 -7762
rect 8533 -7729 8567 -7695
rect 8533 -7797 8567 -7763
rect 8689 -7728 8723 -7694
rect 8689 -7796 8723 -7762
rect 8787 -7729 8821 -7695
rect 8787 -7797 8821 -7763
rect 8998 -7721 9032 -7687
rect 8998 -7823 9032 -7789
rect 9262 -7721 9296 -7687
rect 9262 -7823 9296 -7789
rect 9459 -7728 9493 -7694
rect 9459 -7796 9493 -7762
rect 9559 -7728 9593 -7694
rect 9559 -7796 9593 -7762
rect 9717 -7728 9751 -7694
rect 9717 -7796 9751 -7762
rect 9821 -7729 9855 -7695
rect 9821 -7797 9855 -7763
rect 9977 -7728 10011 -7694
rect 9977 -7796 10011 -7762
rect 10075 -7729 10109 -7695
rect 10075 -7797 10109 -7763
rect 10286 -7721 10320 -7687
rect 10286 -7823 10320 -7789
rect 10550 -7721 10584 -7687
rect 10550 -7823 10584 -7789
rect 10746 -7721 10780 -7687
rect 10746 -7789 10780 -7755
rect 10746 -7857 10780 -7823
rect 10830 -7721 10864 -7687
rect 10830 -7789 10864 -7755
rect 10830 -7857 10864 -7823
rect 10914 -7721 10948 -7687
rect 10914 -7789 10948 -7755
rect 10998 -7721 11032 -7687
rect 10998 -7789 11032 -7755
rect 10998 -7857 11032 -7823
rect 11082 -7721 11116 -7687
rect 11082 -7789 11116 -7755
rect 11166 -7721 11200 -7687
rect 11166 -7789 11200 -7755
rect 11166 -7857 11200 -7823
rect 11250 -7721 11284 -7687
rect 11250 -7789 11284 -7755
rect 11334 -7721 11368 -7687
rect 11334 -7789 11368 -7755
rect 11334 -7857 11368 -7823
rect 11418 -7721 11452 -7687
rect 11418 -7789 11452 -7755
rect 11666 -7721 11700 -7687
rect 11666 -7823 11700 -7789
rect 11930 -7721 11964 -7687
rect 11930 -7823 11964 -7789
rect 13598 -7721 13632 -7687
rect 13598 -7823 13632 -7789
rect 14598 -7721 14632 -7687
rect 14598 -7823 14632 -7789
rect 14794 -7721 14828 -7687
rect 14794 -7823 14828 -7789
rect 15794 -7721 15828 -7687
rect 15794 -7823 15828 -7789
rect 15990 -7721 16024 -7687
rect 15990 -7823 16024 -7789
rect 16622 -7721 16656 -7687
rect 16622 -7823 16656 -7789
rect -2962 -8555 -2928 -8521
rect -2962 -8657 -2928 -8623
rect -2330 -8555 -2296 -8521
rect -2330 -8657 -2296 -8623
rect -1582 -8555 -1548 -8521
rect -1582 -8657 -1548 -8623
rect -950 -8555 -916 -8521
rect -950 -8657 -916 -8623
rect -846 -8555 -812 -8521
rect -846 -8657 -812 -8623
rect -214 -8555 -180 -8521
rect -214 -8657 -180 -8623
rect -18 -8555 16 -8521
rect -18 -8657 16 -8623
rect 246 -8555 280 -8521
rect 246 -8657 280 -8623
rect 457 -8581 491 -8547
rect 457 -8649 491 -8615
rect 555 -8582 589 -8548
rect 555 -8650 589 -8616
rect 711 -8581 745 -8547
rect 711 -8649 745 -8615
rect 815 -8582 849 -8548
rect 815 -8650 849 -8616
rect 973 -8582 1007 -8548
rect 973 -8650 1007 -8616
rect 1073 -8582 1107 -8548
rect 1073 -8650 1107 -8616
rect 1270 -8555 1304 -8521
rect 1270 -8657 1304 -8623
rect 1534 -8555 1568 -8521
rect 1534 -8657 1568 -8623
rect 1730 -8555 1764 -8521
rect 1730 -8657 1764 -8623
rect 2362 -8555 2396 -8521
rect 2362 -8657 2396 -8623
rect 2558 -8555 2592 -8521
rect 2558 -8657 2592 -8623
rect 2822 -8555 2856 -8521
rect 2822 -8657 2856 -8623
rect 3033 -8581 3067 -8547
rect 3033 -8649 3067 -8615
rect 3131 -8582 3165 -8548
rect 3131 -8650 3165 -8616
rect 3287 -8581 3321 -8547
rect 3287 -8649 3321 -8615
rect 3391 -8582 3425 -8548
rect 3391 -8650 3425 -8616
rect 3549 -8582 3583 -8548
rect 3549 -8650 3583 -8616
rect 3649 -8582 3683 -8548
rect 3649 -8650 3683 -8616
rect 3846 -8555 3880 -8521
rect 3846 -8657 3880 -8623
rect 4110 -8555 4144 -8521
rect 4110 -8657 4144 -8623
rect 4306 -8555 4340 -8521
rect 4306 -8657 4340 -8623
rect 4938 -8555 4972 -8521
rect 4938 -8657 4972 -8623
rect 5134 -8555 5168 -8521
rect 5134 -8657 5168 -8623
rect 5398 -8555 5432 -8521
rect 5398 -8657 5432 -8623
rect 5609 -8581 5643 -8547
rect 5609 -8649 5643 -8615
rect 5707 -8582 5741 -8548
rect 5707 -8650 5741 -8616
rect 5863 -8581 5897 -8547
rect 5863 -8649 5897 -8615
rect 5967 -8582 6001 -8548
rect 5967 -8650 6001 -8616
rect 6125 -8582 6159 -8548
rect 6125 -8650 6159 -8616
rect 6225 -8582 6259 -8548
rect 6225 -8650 6259 -8616
rect 6422 -8555 6456 -8521
rect 6422 -8657 6456 -8623
rect 6686 -8555 6720 -8521
rect 6686 -8657 6720 -8623
rect 6882 -8555 6916 -8521
rect 6882 -8657 6916 -8623
rect 7514 -8555 7548 -8521
rect 7514 -8657 7548 -8623
rect 7710 -8555 7744 -8521
rect 7710 -8657 7744 -8623
rect 7974 -8555 8008 -8521
rect 7974 -8657 8008 -8623
rect 8185 -8581 8219 -8547
rect 8185 -8649 8219 -8615
rect 8283 -8582 8317 -8548
rect 8283 -8650 8317 -8616
rect 8439 -8581 8473 -8547
rect 8439 -8649 8473 -8615
rect 8543 -8582 8577 -8548
rect 8543 -8650 8577 -8616
rect 8701 -8582 8735 -8548
rect 8701 -8650 8735 -8616
rect 8801 -8582 8835 -8548
rect 8801 -8650 8835 -8616
rect 8998 -8555 9032 -8521
rect 8998 -8657 9032 -8623
rect 9262 -8555 9296 -8521
rect 9262 -8657 9296 -8623
rect 9458 -8555 9492 -8521
rect 9458 -8657 9492 -8623
rect 10090 -8555 10124 -8521
rect 10090 -8657 10124 -8623
rect 10378 -8555 10412 -8521
rect 10378 -8657 10412 -8623
rect 10642 -8555 10676 -8521
rect 10642 -8657 10676 -8623
rect 10761 -8581 10795 -8547
rect 10761 -8649 10795 -8615
rect 10859 -8582 10893 -8548
rect 10859 -8650 10893 -8616
rect 11015 -8581 11049 -8547
rect 11015 -8649 11049 -8615
rect 11119 -8582 11153 -8548
rect 11119 -8650 11153 -8616
rect 11277 -8582 11311 -8548
rect 11277 -8650 11311 -8616
rect 11377 -8582 11411 -8548
rect 11377 -8650 11411 -8616
rect 11666 -8555 11700 -8521
rect 11666 -8657 11700 -8623
rect 11930 -8555 11964 -8521
rect 11930 -8657 11964 -8623
rect 13690 -8589 13724 -8555
rect 13690 -8657 13724 -8623
rect 13776 -8581 13810 -8547
rect 13776 -8649 13810 -8615
rect 13862 -8589 13896 -8555
rect 13862 -8657 13896 -8623
rect 13948 -8573 13982 -8539
rect 13948 -8641 13982 -8607
rect 14034 -8589 14068 -8555
rect 14034 -8657 14068 -8623
rect 14120 -8527 14154 -8493
rect 14120 -8613 14154 -8579
rect 14206 -8633 14240 -8599
rect 14292 -8527 14326 -8493
rect 14292 -8613 14326 -8579
rect 14378 -8633 14412 -8599
rect 14464 -8527 14498 -8493
rect 14464 -8613 14498 -8579
rect 14550 -8633 14584 -8599
rect 14636 -8527 14670 -8493
rect 14636 -8613 14670 -8579
rect 14722 -8633 14756 -8599
rect 14807 -8527 14841 -8493
rect 14807 -8613 14841 -8579
rect 14893 -8633 14927 -8599
rect 14979 -8527 15013 -8493
rect 14979 -8613 15013 -8579
rect 15065 -8633 15099 -8599
rect 15151 -8527 15185 -8493
rect 15151 -8613 15185 -8579
rect 15237 -8633 15271 -8599
rect 15323 -8527 15357 -8493
rect 15323 -8613 15357 -8579
rect 15409 -8633 15443 -8599
rect 15622 -8555 15656 -8521
rect 15622 -8657 15656 -8623
rect 16622 -8555 16656 -8521
rect 16622 -8657 16656 -8623
rect -2962 -8809 -2928 -8775
rect -2962 -8911 -2928 -8877
rect -2330 -8809 -2296 -8775
rect -2330 -8911 -2296 -8877
rect -1582 -8809 -1548 -8775
rect -1582 -8911 -1548 -8877
rect -950 -8809 -916 -8775
rect -950 -8911 -916 -8877
rect -846 -8809 -812 -8775
rect -846 -8911 -812 -8877
rect -214 -8809 -180 -8775
rect -214 -8911 -180 -8877
rect -18 -8809 16 -8775
rect -18 -8911 16 -8877
rect 246 -8809 280 -8775
rect 246 -8911 280 -8877
rect 443 -8816 477 -8782
rect 443 -8884 477 -8850
rect 543 -8816 577 -8782
rect 543 -8884 577 -8850
rect 701 -8816 735 -8782
rect 701 -8884 735 -8850
rect 805 -8817 839 -8783
rect 805 -8885 839 -8851
rect 961 -8816 995 -8782
rect 961 -8884 995 -8850
rect 1059 -8817 1093 -8783
rect 1059 -8885 1093 -8851
rect 1270 -8809 1304 -8775
rect 1270 -8911 1304 -8877
rect 1534 -8809 1568 -8775
rect 1534 -8911 1568 -8877
rect 1730 -8809 1764 -8775
rect 1730 -8911 1764 -8877
rect 2362 -8809 2396 -8775
rect 2362 -8911 2396 -8877
rect 2558 -8809 2592 -8775
rect 2558 -8911 2592 -8877
rect 2822 -8809 2856 -8775
rect 2822 -8911 2856 -8877
rect 3019 -8816 3053 -8782
rect 3019 -8884 3053 -8850
rect 3119 -8816 3153 -8782
rect 3119 -8884 3153 -8850
rect 3277 -8816 3311 -8782
rect 3277 -8884 3311 -8850
rect 3381 -8817 3415 -8783
rect 3381 -8885 3415 -8851
rect 3537 -8816 3571 -8782
rect 3537 -8884 3571 -8850
rect 3635 -8817 3669 -8783
rect 3635 -8885 3669 -8851
rect 3846 -8809 3880 -8775
rect 3846 -8911 3880 -8877
rect 4110 -8809 4144 -8775
rect 4110 -8911 4144 -8877
rect 4306 -8809 4340 -8775
rect 4306 -8911 4340 -8877
rect 4938 -8809 4972 -8775
rect 4938 -8911 4972 -8877
rect 5134 -8809 5168 -8775
rect 5134 -8911 5168 -8877
rect 5398 -8809 5432 -8775
rect 5398 -8911 5432 -8877
rect 5595 -8816 5629 -8782
rect 5595 -8884 5629 -8850
rect 5695 -8816 5729 -8782
rect 5695 -8884 5729 -8850
rect 5853 -8816 5887 -8782
rect 5853 -8884 5887 -8850
rect 5957 -8817 5991 -8783
rect 5957 -8885 5991 -8851
rect 6113 -8816 6147 -8782
rect 6113 -8884 6147 -8850
rect 6211 -8817 6245 -8783
rect 6211 -8885 6245 -8851
rect 6422 -8809 6456 -8775
rect 6422 -8911 6456 -8877
rect 6686 -8809 6720 -8775
rect 6686 -8911 6720 -8877
rect 6882 -8809 6916 -8775
rect 6882 -8911 6916 -8877
rect 7514 -8809 7548 -8775
rect 7514 -8911 7548 -8877
rect 7710 -8809 7744 -8775
rect 7710 -8911 7744 -8877
rect 7974 -8809 8008 -8775
rect 7974 -8911 8008 -8877
rect 8171 -8816 8205 -8782
rect 8171 -8884 8205 -8850
rect 8271 -8816 8305 -8782
rect 8271 -8884 8305 -8850
rect 8429 -8816 8463 -8782
rect 8429 -8884 8463 -8850
rect 8533 -8817 8567 -8783
rect 8533 -8885 8567 -8851
rect 8689 -8816 8723 -8782
rect 8689 -8884 8723 -8850
rect 8787 -8817 8821 -8783
rect 8787 -8885 8821 -8851
rect 8998 -8809 9032 -8775
rect 8998 -8911 9032 -8877
rect 9262 -8809 9296 -8775
rect 9262 -8911 9296 -8877
rect 9458 -8809 9492 -8775
rect 9458 -8911 9492 -8877
rect 10090 -8809 10124 -8775
rect 10090 -8911 10124 -8877
rect 10378 -8809 10412 -8775
rect 10378 -8911 10412 -8877
rect 10642 -8809 10676 -8775
rect 10642 -8911 10676 -8877
rect 10747 -8816 10781 -8782
rect 10747 -8884 10781 -8850
rect 10847 -8816 10881 -8782
rect 10847 -8884 10881 -8850
rect 11005 -8816 11039 -8782
rect 11005 -8884 11039 -8850
rect 11109 -8817 11143 -8783
rect 11109 -8885 11143 -8851
rect 11265 -8816 11299 -8782
rect 11265 -8884 11299 -8850
rect 11363 -8817 11397 -8783
rect 11363 -8885 11397 -8851
rect 11666 -8809 11700 -8775
rect 11666 -8911 11700 -8877
rect 11930 -8809 11964 -8775
rect 11930 -8911 11964 -8877
rect 12502 -8816 12536 -8782
rect 12502 -8884 12536 -8850
rect 12588 -8823 12622 -8789
rect 12588 -8911 12622 -8877
rect 12674 -8816 12708 -8782
rect 12674 -8884 12708 -8850
rect 12760 -8823 12794 -8789
rect 12760 -8911 12794 -8877
rect 12846 -8816 12880 -8782
rect 12846 -8884 12880 -8850
rect 12932 -8823 12966 -8789
rect 12932 -8911 12966 -8877
rect 13018 -8816 13052 -8782
rect 13018 -8884 13052 -8850
rect 13230 -8809 13264 -8775
rect 13230 -8911 13264 -8877
rect 13494 -8809 13528 -8775
rect 13494 -8911 13528 -8877
rect 13690 -8809 13724 -8775
rect 13690 -8877 13724 -8843
rect 13776 -8817 13810 -8783
rect 13776 -8885 13810 -8851
rect 13862 -8809 13896 -8775
rect 13862 -8877 13896 -8843
rect 13948 -8825 13982 -8791
rect 13948 -8893 13982 -8859
rect 14034 -8809 14068 -8775
rect 14034 -8877 14068 -8843
rect 14120 -8853 14154 -8819
rect 14120 -8939 14154 -8905
rect 14206 -8833 14240 -8799
rect 14292 -8853 14326 -8819
rect 14292 -8939 14326 -8905
rect 14378 -8833 14412 -8799
rect 14464 -8853 14498 -8819
rect 14464 -8939 14498 -8905
rect 14550 -8833 14584 -8799
rect 14636 -8853 14670 -8819
rect 14636 -8939 14670 -8905
rect 14722 -8833 14756 -8799
rect 14807 -8853 14841 -8819
rect 14807 -8939 14841 -8905
rect 14893 -8833 14927 -8799
rect 14979 -8853 15013 -8819
rect 14979 -8939 15013 -8905
rect 15065 -8833 15099 -8799
rect 15151 -8853 15185 -8819
rect 15151 -8939 15185 -8905
rect 15237 -8833 15271 -8799
rect 15323 -8853 15357 -8819
rect 15323 -8939 15357 -8905
rect 15409 -8833 15443 -8799
rect 15622 -8809 15656 -8775
rect 15622 -8911 15656 -8877
rect 16622 -8809 16656 -8775
rect 16622 -8911 16656 -8877
rect -2962 -9643 -2928 -9609
rect -2962 -9745 -2928 -9711
rect -2330 -9643 -2296 -9609
rect -2330 -9745 -2296 -9711
rect -1582 -9643 -1548 -9609
rect -1582 -9745 -1548 -9711
rect -950 -9643 -916 -9609
rect -950 -9745 -916 -9711
rect -831 -9669 -797 -9635
rect -831 -9737 -797 -9703
rect -733 -9670 -699 -9636
rect -733 -9738 -699 -9704
rect -577 -9669 -543 -9635
rect -577 -9737 -543 -9703
rect -473 -9670 -439 -9636
rect -473 -9738 -439 -9704
rect -315 -9670 -281 -9636
rect -315 -9738 -281 -9704
rect -215 -9670 -181 -9636
rect -215 -9738 -181 -9704
rect -18 -9643 16 -9609
rect -18 -9745 16 -9711
rect 246 -9643 280 -9609
rect 246 -9745 280 -9711
rect 457 -9669 491 -9635
rect 457 -9737 491 -9703
rect 555 -9670 589 -9636
rect 555 -9738 589 -9704
rect 711 -9669 745 -9635
rect 711 -9737 745 -9703
rect 815 -9670 849 -9636
rect 815 -9738 849 -9704
rect 973 -9670 1007 -9636
rect 973 -9738 1007 -9704
rect 1073 -9670 1107 -9636
rect 1073 -9738 1107 -9704
rect 1270 -9643 1304 -9609
rect 1270 -9745 1304 -9711
rect 1534 -9643 1568 -9609
rect 1534 -9745 1568 -9711
rect 1730 -9643 1764 -9609
rect 1730 -9745 1764 -9711
rect 2362 -9643 2396 -9609
rect 2362 -9745 2396 -9711
rect 2558 -9643 2592 -9609
rect 2558 -9745 2592 -9711
rect 2822 -9643 2856 -9609
rect 2822 -9745 2856 -9711
rect 3033 -9669 3067 -9635
rect 3033 -9737 3067 -9703
rect 3131 -9670 3165 -9636
rect 3131 -9738 3165 -9704
rect 3287 -9669 3321 -9635
rect 3287 -9737 3321 -9703
rect 3391 -9670 3425 -9636
rect 3391 -9738 3425 -9704
rect 3549 -9670 3583 -9636
rect 3549 -9738 3583 -9704
rect 3649 -9670 3683 -9636
rect 3649 -9738 3683 -9704
rect 3846 -9643 3880 -9609
rect 3846 -9745 3880 -9711
rect 4110 -9643 4144 -9609
rect 4110 -9745 4144 -9711
rect 4306 -9643 4340 -9609
rect 4306 -9745 4340 -9711
rect 4938 -9643 4972 -9609
rect 4938 -9745 4972 -9711
rect 5134 -9643 5168 -9609
rect 5134 -9745 5168 -9711
rect 5398 -9643 5432 -9609
rect 5398 -9745 5432 -9711
rect 5609 -9669 5643 -9635
rect 5609 -9737 5643 -9703
rect 5707 -9670 5741 -9636
rect 5707 -9738 5741 -9704
rect 5863 -9669 5897 -9635
rect 5863 -9737 5897 -9703
rect 5967 -9670 6001 -9636
rect 5967 -9738 6001 -9704
rect 6125 -9670 6159 -9636
rect 6125 -9738 6159 -9704
rect 6225 -9670 6259 -9636
rect 6225 -9738 6259 -9704
rect 6422 -9643 6456 -9609
rect 6422 -9745 6456 -9711
rect 6686 -9643 6720 -9609
rect 6686 -9745 6720 -9711
rect 6882 -9643 6916 -9609
rect 6882 -9745 6916 -9711
rect 7514 -9643 7548 -9609
rect 7514 -9745 7548 -9711
rect 7710 -9643 7744 -9609
rect 7710 -9745 7744 -9711
rect 7974 -9643 8008 -9609
rect 7974 -9745 8008 -9711
rect 8185 -9669 8219 -9635
rect 8185 -9737 8219 -9703
rect 8283 -9670 8317 -9636
rect 8283 -9738 8317 -9704
rect 8439 -9669 8473 -9635
rect 8439 -9737 8473 -9703
rect 8543 -9670 8577 -9636
rect 8543 -9738 8577 -9704
rect 8701 -9670 8735 -9636
rect 8701 -9738 8735 -9704
rect 8801 -9670 8835 -9636
rect 8801 -9738 8835 -9704
rect 8998 -9643 9032 -9609
rect 8998 -9745 9032 -9711
rect 9262 -9643 9296 -9609
rect 9262 -9745 9296 -9711
rect 9458 -9643 9492 -9609
rect 9458 -9745 9492 -9711
rect 10090 -9643 10124 -9609
rect 10090 -9745 10124 -9711
rect 10378 -9643 10412 -9609
rect 10378 -9745 10412 -9711
rect 10642 -9643 10676 -9609
rect 10642 -9745 10676 -9711
rect 10761 -9669 10795 -9635
rect 10761 -9737 10795 -9703
rect 10859 -9670 10893 -9636
rect 10859 -9738 10893 -9704
rect 11015 -9669 11049 -9635
rect 11015 -9737 11049 -9703
rect 11119 -9670 11153 -9636
rect 11119 -9738 11153 -9704
rect 11277 -9670 11311 -9636
rect 11277 -9738 11311 -9704
rect 11377 -9670 11411 -9636
rect 11377 -9738 11411 -9704
rect 11666 -9643 11700 -9609
rect 11666 -9745 11700 -9711
rect 11930 -9643 11964 -9609
rect 11930 -9745 11964 -9711
rect 13690 -9677 13724 -9643
rect 13690 -9745 13724 -9711
rect 13776 -9669 13810 -9635
rect 13776 -9737 13810 -9703
rect 13862 -9677 13896 -9643
rect 13862 -9745 13896 -9711
rect 13948 -9661 13982 -9627
rect 13948 -9729 13982 -9695
rect 14034 -9677 14068 -9643
rect 14034 -9745 14068 -9711
rect 14120 -9615 14154 -9581
rect 14120 -9701 14154 -9667
rect 14206 -9721 14240 -9687
rect 14292 -9615 14326 -9581
rect 14292 -9701 14326 -9667
rect 14378 -9721 14412 -9687
rect 14464 -9615 14498 -9581
rect 14464 -9701 14498 -9667
rect 14550 -9721 14584 -9687
rect 14636 -9615 14670 -9581
rect 14636 -9701 14670 -9667
rect 14722 -9721 14756 -9687
rect 14807 -9615 14841 -9581
rect 14807 -9701 14841 -9667
rect 14893 -9721 14927 -9687
rect 14979 -9615 15013 -9581
rect 14979 -9701 15013 -9667
rect 15065 -9721 15099 -9687
rect 15151 -9615 15185 -9581
rect 15151 -9701 15185 -9667
rect 15237 -9721 15271 -9687
rect 15323 -9615 15357 -9581
rect 15323 -9701 15357 -9667
rect 15409 -9721 15443 -9687
rect 15622 -9643 15656 -9609
rect 15622 -9745 15656 -9711
rect 16622 -9643 16656 -9609
rect 16622 -9745 16656 -9711
rect -2962 -9897 -2928 -9863
rect -2962 -9999 -2928 -9965
rect -2330 -9897 -2296 -9863
rect -2330 -9999 -2296 -9965
rect -1582 -9897 -1548 -9863
rect -1582 -9999 -1548 -9965
rect -950 -9897 -916 -9863
rect -950 -9999 -916 -9965
rect -846 -9897 -812 -9863
rect -846 -9999 -812 -9965
rect -214 -9897 -180 -9863
rect -214 -9999 -180 -9965
rect -18 -9897 16 -9863
rect -18 -9999 16 -9965
rect 246 -9897 280 -9863
rect 246 -9999 280 -9965
rect 443 -9904 477 -9870
rect 443 -9972 477 -9938
rect 543 -9904 577 -9870
rect 543 -9972 577 -9938
rect 701 -9904 735 -9870
rect 701 -9972 735 -9938
rect 805 -9905 839 -9871
rect 805 -9973 839 -9939
rect 961 -9904 995 -9870
rect 961 -9972 995 -9938
rect 1059 -9905 1093 -9871
rect 1059 -9973 1093 -9939
rect 1270 -9897 1304 -9863
rect 1270 -9999 1304 -9965
rect 1534 -9897 1568 -9863
rect 1534 -9999 1568 -9965
rect 1730 -9897 1764 -9863
rect 1730 -9999 1764 -9965
rect 2362 -9897 2396 -9863
rect 2362 -9999 2396 -9965
rect 2558 -9897 2592 -9863
rect 2558 -9999 2592 -9965
rect 2822 -9897 2856 -9863
rect 2822 -9999 2856 -9965
rect 3019 -9904 3053 -9870
rect 3019 -9972 3053 -9938
rect 3119 -9904 3153 -9870
rect 3119 -9972 3153 -9938
rect 3277 -9904 3311 -9870
rect 3277 -9972 3311 -9938
rect 3381 -9905 3415 -9871
rect 3381 -9973 3415 -9939
rect 3537 -9904 3571 -9870
rect 3537 -9972 3571 -9938
rect 3635 -9905 3669 -9871
rect 3635 -9973 3669 -9939
rect 3846 -9897 3880 -9863
rect 3846 -9999 3880 -9965
rect 4110 -9897 4144 -9863
rect 4110 -9999 4144 -9965
rect 4306 -9897 4340 -9863
rect 4306 -9999 4340 -9965
rect 4938 -9897 4972 -9863
rect 4938 -9999 4972 -9965
rect 5134 -9897 5168 -9863
rect 5134 -9999 5168 -9965
rect 5398 -9897 5432 -9863
rect 5398 -9999 5432 -9965
rect 5595 -9904 5629 -9870
rect 5595 -9972 5629 -9938
rect 5695 -9904 5729 -9870
rect 5695 -9972 5729 -9938
rect 5853 -9904 5887 -9870
rect 5853 -9972 5887 -9938
rect 5957 -9905 5991 -9871
rect 5957 -9973 5991 -9939
rect 6113 -9904 6147 -9870
rect 6113 -9972 6147 -9938
rect 6211 -9905 6245 -9871
rect 6211 -9973 6245 -9939
rect 6422 -9897 6456 -9863
rect 6422 -9999 6456 -9965
rect 6686 -9897 6720 -9863
rect 6686 -9999 6720 -9965
rect 6882 -9897 6916 -9863
rect 6882 -9999 6916 -9965
rect 7514 -9897 7548 -9863
rect 7514 -9999 7548 -9965
rect 7710 -9897 7744 -9863
rect 7710 -9999 7744 -9965
rect 7974 -9897 8008 -9863
rect 7974 -9999 8008 -9965
rect 8171 -9904 8205 -9870
rect 8171 -9972 8205 -9938
rect 8271 -9904 8305 -9870
rect 8271 -9972 8305 -9938
rect 8429 -9904 8463 -9870
rect 8429 -9972 8463 -9938
rect 8533 -9905 8567 -9871
rect 8533 -9973 8567 -9939
rect 8689 -9904 8723 -9870
rect 8689 -9972 8723 -9938
rect 8787 -9905 8821 -9871
rect 8787 -9973 8821 -9939
rect 8998 -9897 9032 -9863
rect 8998 -9999 9032 -9965
rect 9262 -9897 9296 -9863
rect 9262 -9999 9296 -9965
rect 9458 -9897 9492 -9863
rect 9458 -9999 9492 -9965
rect 10090 -9897 10124 -9863
rect 10090 -9999 10124 -9965
rect 10378 -9897 10412 -9863
rect 10378 -9999 10412 -9965
rect 10642 -9897 10676 -9863
rect 10642 -9999 10676 -9965
rect 10747 -9904 10781 -9870
rect 10747 -9972 10781 -9938
rect 10847 -9904 10881 -9870
rect 10847 -9972 10881 -9938
rect 11005 -9904 11039 -9870
rect 11005 -9972 11039 -9938
rect 11109 -9905 11143 -9871
rect 11109 -9973 11143 -9939
rect 11265 -9904 11299 -9870
rect 11265 -9972 11299 -9938
rect 11363 -9905 11397 -9871
rect 11363 -9973 11397 -9939
rect 11666 -9897 11700 -9863
rect 11666 -9999 11700 -9965
rect 11930 -9897 11964 -9863
rect 11930 -9999 11964 -9965
rect 12502 -9904 12536 -9870
rect 12502 -9972 12536 -9938
rect 12588 -9911 12622 -9877
rect 12588 -9999 12622 -9965
rect 12674 -9904 12708 -9870
rect 12674 -9972 12708 -9938
rect 12760 -9911 12794 -9877
rect 12760 -9999 12794 -9965
rect 12846 -9904 12880 -9870
rect 12846 -9972 12880 -9938
rect 12932 -9911 12966 -9877
rect 12932 -9999 12966 -9965
rect 13018 -9904 13052 -9870
rect 13018 -9972 13052 -9938
rect 13230 -9897 13264 -9863
rect 13230 -9999 13264 -9965
rect 13494 -9897 13528 -9863
rect 13494 -9999 13528 -9965
rect 13690 -9897 13724 -9863
rect 13690 -9965 13724 -9931
rect 13776 -9905 13810 -9871
rect 13776 -9973 13810 -9939
rect 13862 -9897 13896 -9863
rect 13862 -9965 13896 -9931
rect 13948 -9913 13982 -9879
rect 13948 -9981 13982 -9947
rect 14034 -9897 14068 -9863
rect 14034 -9965 14068 -9931
rect 14120 -9941 14154 -9907
rect 14120 -10027 14154 -9993
rect 14206 -9921 14240 -9887
rect 14292 -9941 14326 -9907
rect 14292 -10027 14326 -9993
rect 14378 -9921 14412 -9887
rect 14464 -9941 14498 -9907
rect 14464 -10027 14498 -9993
rect 14550 -9921 14584 -9887
rect 14636 -9941 14670 -9907
rect 14636 -10027 14670 -9993
rect 14722 -9921 14756 -9887
rect 14807 -9941 14841 -9907
rect 14807 -10027 14841 -9993
rect 14893 -9921 14927 -9887
rect 14979 -9941 15013 -9907
rect 14979 -10027 15013 -9993
rect 15065 -9921 15099 -9887
rect 15151 -9941 15185 -9907
rect 15151 -10027 15185 -9993
rect 15237 -9921 15271 -9887
rect 15323 -9941 15357 -9907
rect 15323 -10027 15357 -9993
rect 15409 -9921 15443 -9887
rect 15622 -9897 15656 -9863
rect 15622 -9999 15656 -9965
rect 16622 -9897 16656 -9863
rect 16622 -9999 16656 -9965
rect -2962 -10731 -2928 -10697
rect -2962 -10833 -2928 -10799
rect -2330 -10731 -2296 -10697
rect -2330 -10833 -2296 -10799
rect -1950 -10731 -1916 -10697
rect -1950 -10833 -1916 -10799
rect -1866 -10731 -1832 -10697
rect -1866 -10833 -1832 -10799
rect -1782 -10731 -1748 -10697
rect -1782 -10833 -1748 -10799
rect -1582 -10731 -1548 -10697
rect -1582 -10833 -1548 -10799
rect -950 -10731 -916 -10697
rect -950 -10833 -916 -10799
rect -846 -10731 -812 -10697
rect -846 -10833 -812 -10799
rect -214 -10731 -180 -10697
rect -214 -10833 -180 -10799
rect -18 -10731 16 -10697
rect -18 -10833 16 -10799
rect 246 -10731 280 -10697
rect 246 -10833 280 -10799
rect 457 -10757 491 -10723
rect 457 -10825 491 -10791
rect 555 -10758 589 -10724
rect 555 -10826 589 -10792
rect 711 -10757 745 -10723
rect 711 -10825 745 -10791
rect 815 -10758 849 -10724
rect 815 -10826 849 -10792
rect 973 -10758 1007 -10724
rect 973 -10826 1007 -10792
rect 1073 -10758 1107 -10724
rect 1073 -10826 1107 -10792
rect 1270 -10731 1304 -10697
rect 1270 -10833 1304 -10799
rect 1534 -10731 1568 -10697
rect 1534 -10833 1568 -10799
rect 1730 -10731 1764 -10697
rect 1730 -10833 1764 -10799
rect 2362 -10731 2396 -10697
rect 2362 -10833 2396 -10799
rect 2558 -10731 2592 -10697
rect 2558 -10833 2592 -10799
rect 2822 -10731 2856 -10697
rect 2822 -10833 2856 -10799
rect 3033 -10757 3067 -10723
rect 3033 -10825 3067 -10791
rect 3131 -10758 3165 -10724
rect 3131 -10826 3165 -10792
rect 3287 -10757 3321 -10723
rect 3287 -10825 3321 -10791
rect 3391 -10758 3425 -10724
rect 3391 -10826 3425 -10792
rect 3549 -10758 3583 -10724
rect 3549 -10826 3583 -10792
rect 3649 -10758 3683 -10724
rect 3649 -10826 3683 -10792
rect 3846 -10731 3880 -10697
rect 3846 -10833 3880 -10799
rect 4110 -10731 4144 -10697
rect 4110 -10833 4144 -10799
rect 4306 -10731 4340 -10697
rect 4306 -10833 4340 -10799
rect 4938 -10731 4972 -10697
rect 4938 -10833 4972 -10799
rect 5134 -10731 5168 -10697
rect 5134 -10833 5168 -10799
rect 5398 -10731 5432 -10697
rect 5398 -10833 5432 -10799
rect 5609 -10757 5643 -10723
rect 5609 -10825 5643 -10791
rect 5707 -10758 5741 -10724
rect 5707 -10826 5741 -10792
rect 5863 -10757 5897 -10723
rect 5863 -10825 5897 -10791
rect 5967 -10758 6001 -10724
rect 5967 -10826 6001 -10792
rect 6125 -10758 6159 -10724
rect 6125 -10826 6159 -10792
rect 6225 -10758 6259 -10724
rect 6225 -10826 6259 -10792
rect 6422 -10731 6456 -10697
rect 6422 -10833 6456 -10799
rect 6686 -10731 6720 -10697
rect 6686 -10833 6720 -10799
rect 6882 -10731 6916 -10697
rect 6882 -10833 6916 -10799
rect 7514 -10731 7548 -10697
rect 7514 -10833 7548 -10799
rect 7710 -10731 7744 -10697
rect 7710 -10833 7744 -10799
rect 7974 -10731 8008 -10697
rect 7974 -10833 8008 -10799
rect 8185 -10757 8219 -10723
rect 8185 -10825 8219 -10791
rect 8283 -10758 8317 -10724
rect 8283 -10826 8317 -10792
rect 8439 -10757 8473 -10723
rect 8439 -10825 8473 -10791
rect 8543 -10758 8577 -10724
rect 8543 -10826 8577 -10792
rect 8701 -10758 8735 -10724
rect 8701 -10826 8735 -10792
rect 8801 -10758 8835 -10724
rect 8801 -10826 8835 -10792
rect 8998 -10731 9032 -10697
rect 8998 -10833 9032 -10799
rect 9262 -10731 9296 -10697
rect 9262 -10833 9296 -10799
rect 9458 -10731 9492 -10697
rect 9458 -10833 9492 -10799
rect 10090 -10731 10124 -10697
rect 10090 -10833 10124 -10799
rect 10378 -10731 10412 -10697
rect 10378 -10833 10412 -10799
rect 10642 -10731 10676 -10697
rect 10642 -10833 10676 -10799
rect 10761 -10757 10795 -10723
rect 10761 -10825 10795 -10791
rect 10859 -10758 10893 -10724
rect 10859 -10826 10893 -10792
rect 11015 -10757 11049 -10723
rect 11015 -10825 11049 -10791
rect 11119 -10758 11153 -10724
rect 11119 -10826 11153 -10792
rect 11277 -10758 11311 -10724
rect 11277 -10826 11311 -10792
rect 11377 -10758 11411 -10724
rect 11377 -10826 11411 -10792
rect 11666 -10731 11700 -10697
rect 11666 -10833 11700 -10799
rect 11930 -10731 11964 -10697
rect 11930 -10833 11964 -10799
rect 13598 -10731 13632 -10697
rect 13598 -10833 13632 -10799
rect 14598 -10731 14632 -10697
rect 14598 -10833 14632 -10799
rect 14794 -10731 14828 -10697
rect 14794 -10833 14828 -10799
rect 15794 -10731 15828 -10697
rect 15794 -10833 15828 -10799
rect 15990 -10731 16024 -10697
rect 15990 -10833 16024 -10799
rect 16622 -10731 16656 -10697
rect 16622 -10833 16656 -10799
rect -2962 -10985 -2928 -10951
rect -2962 -11087 -2928 -11053
rect -2330 -10985 -2296 -10951
rect -2330 -11087 -2296 -11053
rect -1582 -10985 -1548 -10951
rect -1582 -11087 -1548 -11053
rect -950 -10985 -916 -10951
rect -950 -11087 -916 -11053
rect -846 -10985 -812 -10951
rect -846 -11087 -812 -11053
rect -214 -10985 -180 -10951
rect -214 -11087 -180 -11053
rect -18 -10985 16 -10951
rect -18 -11087 16 -11053
rect 246 -10985 280 -10951
rect 246 -11087 280 -11053
rect 457 -10993 491 -10959
rect 457 -11061 491 -11027
rect 555 -10992 589 -10958
rect 555 -11060 589 -11026
rect 711 -10993 745 -10959
rect 711 -11061 745 -11027
rect 815 -10992 849 -10958
rect 815 -11060 849 -11026
rect 973 -10992 1007 -10958
rect 973 -11060 1007 -11026
rect 1073 -10992 1107 -10958
rect 1073 -11060 1107 -11026
rect 1270 -10985 1304 -10951
rect 1270 -11087 1304 -11053
rect 1534 -10985 1568 -10951
rect 1534 -11087 1568 -11053
rect 1730 -10985 1764 -10951
rect 1730 -11087 1764 -11053
rect 2362 -10985 2396 -10951
rect 2362 -11087 2396 -11053
rect 2558 -10985 2592 -10951
rect 2558 -11087 2592 -11053
rect 2822 -10985 2856 -10951
rect 2822 -11087 2856 -11053
rect 3033 -10993 3067 -10959
rect 3033 -11061 3067 -11027
rect 3131 -10992 3165 -10958
rect 3131 -11060 3165 -11026
rect 3287 -10993 3321 -10959
rect 3287 -11061 3321 -11027
rect 3391 -10992 3425 -10958
rect 3391 -11060 3425 -11026
rect 3549 -10992 3583 -10958
rect 3549 -11060 3583 -11026
rect 3649 -10992 3683 -10958
rect 3649 -11060 3683 -11026
rect 3846 -10985 3880 -10951
rect 3846 -11087 3880 -11053
rect 4110 -10985 4144 -10951
rect 4110 -11087 4144 -11053
rect 4306 -10985 4340 -10951
rect 4306 -11087 4340 -11053
rect 4938 -10985 4972 -10951
rect 4938 -11087 4972 -11053
rect 5134 -10985 5168 -10951
rect 5134 -11087 5168 -11053
rect 5398 -10985 5432 -10951
rect 5398 -11087 5432 -11053
rect 5609 -10993 5643 -10959
rect 5609 -11061 5643 -11027
rect 5707 -10992 5741 -10958
rect 5707 -11060 5741 -11026
rect 5863 -10993 5897 -10959
rect 5863 -11061 5897 -11027
rect 5967 -10992 6001 -10958
rect 5967 -11060 6001 -11026
rect 6125 -10992 6159 -10958
rect 6125 -11060 6159 -11026
rect 6225 -10992 6259 -10958
rect 6225 -11060 6259 -11026
rect 6422 -10985 6456 -10951
rect 6422 -11087 6456 -11053
rect 6686 -10985 6720 -10951
rect 6686 -11087 6720 -11053
rect 6882 -10985 6916 -10951
rect 6882 -11087 6916 -11053
rect 7514 -10985 7548 -10951
rect 7514 -11087 7548 -11053
rect 7710 -10985 7744 -10951
rect 7710 -11087 7744 -11053
rect 7974 -10985 8008 -10951
rect 7974 -11087 8008 -11053
rect 8185 -10993 8219 -10959
rect 8185 -11061 8219 -11027
rect 8283 -10992 8317 -10958
rect 8283 -11060 8317 -11026
rect 8439 -10993 8473 -10959
rect 8439 -11061 8473 -11027
rect 8543 -10992 8577 -10958
rect 8543 -11060 8577 -11026
rect 8701 -10992 8735 -10958
rect 8701 -11060 8735 -11026
rect 8801 -10992 8835 -10958
rect 8801 -11060 8835 -11026
rect 8998 -10985 9032 -10951
rect 8998 -11087 9032 -11053
rect 9262 -10985 9296 -10951
rect 9262 -11087 9296 -11053
rect 9458 -10985 9492 -10951
rect 9458 -11087 9492 -11053
rect 10090 -10985 10124 -10951
rect 10090 -11087 10124 -11053
rect 10378 -10985 10412 -10951
rect 10378 -11087 10412 -11053
rect 10642 -10985 10676 -10951
rect 10642 -11087 10676 -11053
rect 10761 -10993 10795 -10959
rect 10761 -11061 10795 -11027
rect 10859 -10992 10893 -10958
rect 10859 -11060 10893 -11026
rect 11015 -10993 11049 -10959
rect 11015 -11061 11049 -11027
rect 11119 -10992 11153 -10958
rect 11119 -11060 11153 -11026
rect 11277 -10992 11311 -10958
rect 11277 -11060 11311 -11026
rect 11377 -10992 11411 -10958
rect 11377 -11060 11411 -11026
rect 11666 -10985 11700 -10951
rect 11666 -11087 11700 -11053
rect 11930 -10985 11964 -10951
rect 11930 -11087 11964 -11053
rect 13598 -10985 13632 -10951
rect 13598 -11087 13632 -11053
rect 14598 -10985 14632 -10951
rect 14598 -11087 14632 -11053
rect 14794 -10985 14828 -10951
rect 14794 -11087 14828 -11053
rect 15794 -10985 15828 -10951
rect 15794 -11087 15828 -11053
rect 15990 -10985 16024 -10951
rect 15990 -11087 16024 -11053
rect 16622 -10985 16656 -10951
rect 16622 -11087 16656 -11053
rect -2962 -11819 -2928 -11785
rect -2962 -11921 -2928 -11887
rect -2330 -11819 -2296 -11785
rect -2330 -11921 -2296 -11887
rect -1582 -11819 -1548 -11785
rect -1582 -11921 -1548 -11887
rect -950 -11819 -916 -11785
rect -950 -11921 -916 -11887
rect -846 -11819 -812 -11785
rect -846 -11921 -812 -11887
rect -214 -11819 -180 -11785
rect -214 -11921 -180 -11887
rect -18 -11819 16 -11785
rect -18 -11921 16 -11887
rect 246 -11819 280 -11785
rect 246 -11921 280 -11887
rect 443 -11846 477 -11812
rect 443 -11914 477 -11880
rect 543 -11846 577 -11812
rect 543 -11914 577 -11880
rect 701 -11846 735 -11812
rect 701 -11914 735 -11880
rect 805 -11845 839 -11811
rect 805 -11913 839 -11879
rect 961 -11846 995 -11812
rect 961 -11914 995 -11880
rect 1059 -11845 1093 -11811
rect 1059 -11913 1093 -11879
rect 1270 -11819 1304 -11785
rect 1270 -11921 1304 -11887
rect 1534 -11819 1568 -11785
rect 1534 -11921 1568 -11887
rect 1730 -11819 1764 -11785
rect 1730 -11921 1764 -11887
rect 2362 -11819 2396 -11785
rect 2362 -11921 2396 -11887
rect 2558 -11819 2592 -11785
rect 2558 -11921 2592 -11887
rect 2822 -11819 2856 -11785
rect 2822 -11921 2856 -11887
rect 3019 -11846 3053 -11812
rect 3019 -11914 3053 -11880
rect 3119 -11846 3153 -11812
rect 3119 -11914 3153 -11880
rect 3277 -11846 3311 -11812
rect 3277 -11914 3311 -11880
rect 3381 -11845 3415 -11811
rect 3381 -11913 3415 -11879
rect 3537 -11846 3571 -11812
rect 3537 -11914 3571 -11880
rect 3635 -11845 3669 -11811
rect 3635 -11913 3669 -11879
rect 3846 -11819 3880 -11785
rect 3846 -11921 3880 -11887
rect 4110 -11819 4144 -11785
rect 4110 -11921 4144 -11887
rect 4306 -11819 4340 -11785
rect 4306 -11921 4340 -11887
rect 4938 -11819 4972 -11785
rect 4938 -11921 4972 -11887
rect 5134 -11819 5168 -11785
rect 5134 -11921 5168 -11887
rect 5398 -11819 5432 -11785
rect 5398 -11921 5432 -11887
rect 5595 -11846 5629 -11812
rect 5595 -11914 5629 -11880
rect 5695 -11846 5729 -11812
rect 5695 -11914 5729 -11880
rect 5853 -11846 5887 -11812
rect 5853 -11914 5887 -11880
rect 5957 -11845 5991 -11811
rect 5957 -11913 5991 -11879
rect 6113 -11846 6147 -11812
rect 6113 -11914 6147 -11880
rect 6211 -11845 6245 -11811
rect 6211 -11913 6245 -11879
rect 6422 -11819 6456 -11785
rect 6422 -11921 6456 -11887
rect 6686 -11819 6720 -11785
rect 6686 -11921 6720 -11887
rect 6882 -11819 6916 -11785
rect 6882 -11921 6916 -11887
rect 7514 -11819 7548 -11785
rect 7514 -11921 7548 -11887
rect 7710 -11819 7744 -11785
rect 7710 -11921 7744 -11887
rect 7974 -11819 8008 -11785
rect 7974 -11921 8008 -11887
rect 8171 -11846 8205 -11812
rect 8171 -11914 8205 -11880
rect 8271 -11846 8305 -11812
rect 8271 -11914 8305 -11880
rect 8429 -11846 8463 -11812
rect 8429 -11914 8463 -11880
rect 8533 -11845 8567 -11811
rect 8533 -11913 8567 -11879
rect 8689 -11846 8723 -11812
rect 8689 -11914 8723 -11880
rect 8787 -11845 8821 -11811
rect 8787 -11913 8821 -11879
rect 8998 -11819 9032 -11785
rect 8998 -11921 9032 -11887
rect 9262 -11819 9296 -11785
rect 9262 -11921 9296 -11887
rect 9458 -11819 9492 -11785
rect 9458 -11921 9492 -11887
rect 10090 -11819 10124 -11785
rect 10090 -11921 10124 -11887
rect 10378 -11819 10412 -11785
rect 10378 -11921 10412 -11887
rect 10642 -11819 10676 -11785
rect 10642 -11921 10676 -11887
rect 10747 -11846 10781 -11812
rect 10747 -11914 10781 -11880
rect 10847 -11846 10881 -11812
rect 10847 -11914 10881 -11880
rect 11005 -11846 11039 -11812
rect 11005 -11914 11039 -11880
rect 11109 -11845 11143 -11811
rect 11109 -11913 11143 -11879
rect 11265 -11846 11299 -11812
rect 11265 -11914 11299 -11880
rect 11363 -11845 11397 -11811
rect 11363 -11913 11397 -11879
rect 11666 -11819 11700 -11785
rect 11666 -11921 11700 -11887
rect 11930 -11819 11964 -11785
rect 11930 -11921 11964 -11887
rect 12502 -11846 12536 -11812
rect 12502 -11914 12536 -11880
rect 12588 -11819 12622 -11785
rect 12588 -11907 12622 -11873
rect 12674 -11846 12708 -11812
rect 12674 -11914 12708 -11880
rect 12760 -11819 12794 -11785
rect 12760 -11907 12794 -11873
rect 12846 -11846 12880 -11812
rect 12846 -11914 12880 -11880
rect 12932 -11819 12966 -11785
rect 12932 -11907 12966 -11873
rect 13018 -11846 13052 -11812
rect 13018 -11914 13052 -11880
rect 13230 -11819 13264 -11785
rect 13230 -11921 13264 -11887
rect 13494 -11819 13528 -11785
rect 13494 -11921 13528 -11887
rect 13690 -11853 13724 -11819
rect 13690 -11921 13724 -11887
rect 13776 -11845 13810 -11811
rect 13776 -11913 13810 -11879
rect 13862 -11853 13896 -11819
rect 13862 -11921 13896 -11887
rect 13948 -11837 13982 -11803
rect 13948 -11905 13982 -11871
rect 14034 -11853 14068 -11819
rect 14034 -11921 14068 -11887
rect 14120 -11791 14154 -11757
rect 14120 -11877 14154 -11843
rect 14206 -11897 14240 -11863
rect 14292 -11791 14326 -11757
rect 14292 -11877 14326 -11843
rect 14378 -11897 14412 -11863
rect 14464 -11791 14498 -11757
rect 14464 -11877 14498 -11843
rect 14550 -11897 14584 -11863
rect 14636 -11791 14670 -11757
rect 14636 -11877 14670 -11843
rect 14722 -11897 14756 -11863
rect 14807 -11791 14841 -11757
rect 14807 -11877 14841 -11843
rect 14893 -11897 14927 -11863
rect 14979 -11791 15013 -11757
rect 14979 -11877 15013 -11843
rect 15065 -11897 15099 -11863
rect 15151 -11791 15185 -11757
rect 15151 -11877 15185 -11843
rect 15237 -11897 15271 -11863
rect 15323 -11791 15357 -11757
rect 15323 -11877 15357 -11843
rect 15409 -11897 15443 -11863
rect 15622 -11819 15656 -11785
rect 15622 -11921 15656 -11887
rect 16622 -11819 16656 -11785
rect 16622 -11921 16656 -11887
rect -2962 -12073 -2928 -12039
rect -2962 -12175 -2928 -12141
rect -2330 -12073 -2296 -12039
rect -2330 -12175 -2296 -12141
rect -1582 -12073 -1548 -12039
rect -1582 -12175 -1548 -12141
rect -950 -12073 -916 -12039
rect -950 -12175 -916 -12141
rect -831 -12081 -797 -12047
rect -831 -12149 -797 -12115
rect -733 -12080 -699 -12046
rect -733 -12148 -699 -12114
rect -577 -12081 -543 -12047
rect -577 -12149 -543 -12115
rect -473 -12080 -439 -12046
rect -473 -12148 -439 -12114
rect -315 -12080 -281 -12046
rect -315 -12148 -281 -12114
rect -215 -12080 -181 -12046
rect -215 -12148 -181 -12114
rect -18 -12073 16 -12039
rect -18 -12175 16 -12141
rect 246 -12073 280 -12039
rect 246 -12175 280 -12141
rect 457 -12081 491 -12047
rect 457 -12149 491 -12115
rect 555 -12080 589 -12046
rect 555 -12148 589 -12114
rect 711 -12081 745 -12047
rect 711 -12149 745 -12115
rect 815 -12080 849 -12046
rect 815 -12148 849 -12114
rect 973 -12080 1007 -12046
rect 973 -12148 1007 -12114
rect 1073 -12080 1107 -12046
rect 1073 -12148 1107 -12114
rect 1270 -12073 1304 -12039
rect 1270 -12175 1304 -12141
rect 1534 -12073 1568 -12039
rect 1534 -12175 1568 -12141
rect 1730 -12073 1764 -12039
rect 1730 -12175 1764 -12141
rect 2362 -12073 2396 -12039
rect 2362 -12175 2396 -12141
rect 2558 -12073 2592 -12039
rect 2558 -12175 2592 -12141
rect 2822 -12073 2856 -12039
rect 2822 -12175 2856 -12141
rect 3033 -12081 3067 -12047
rect 3033 -12149 3067 -12115
rect 3131 -12080 3165 -12046
rect 3131 -12148 3165 -12114
rect 3287 -12081 3321 -12047
rect 3287 -12149 3321 -12115
rect 3391 -12080 3425 -12046
rect 3391 -12148 3425 -12114
rect 3549 -12080 3583 -12046
rect 3549 -12148 3583 -12114
rect 3649 -12080 3683 -12046
rect 3649 -12148 3683 -12114
rect 3846 -12073 3880 -12039
rect 3846 -12175 3880 -12141
rect 4110 -12073 4144 -12039
rect 4110 -12175 4144 -12141
rect 4306 -12073 4340 -12039
rect 4306 -12175 4340 -12141
rect 4938 -12073 4972 -12039
rect 4938 -12175 4972 -12141
rect 5134 -12073 5168 -12039
rect 5134 -12175 5168 -12141
rect 5398 -12073 5432 -12039
rect 5398 -12175 5432 -12141
rect 5609 -12081 5643 -12047
rect 5609 -12149 5643 -12115
rect 5707 -12080 5741 -12046
rect 5707 -12148 5741 -12114
rect 5863 -12081 5897 -12047
rect 5863 -12149 5897 -12115
rect 5967 -12080 6001 -12046
rect 5967 -12148 6001 -12114
rect 6125 -12080 6159 -12046
rect 6125 -12148 6159 -12114
rect 6225 -12080 6259 -12046
rect 6225 -12148 6259 -12114
rect 6422 -12073 6456 -12039
rect 6422 -12175 6456 -12141
rect 6686 -12073 6720 -12039
rect 6686 -12175 6720 -12141
rect 6882 -12073 6916 -12039
rect 6882 -12175 6916 -12141
rect 7514 -12073 7548 -12039
rect 7514 -12175 7548 -12141
rect 7710 -12073 7744 -12039
rect 7710 -12175 7744 -12141
rect 7974 -12073 8008 -12039
rect 7974 -12175 8008 -12141
rect 8185 -12081 8219 -12047
rect 8185 -12149 8219 -12115
rect 8283 -12080 8317 -12046
rect 8283 -12148 8317 -12114
rect 8439 -12081 8473 -12047
rect 8439 -12149 8473 -12115
rect 8543 -12080 8577 -12046
rect 8543 -12148 8577 -12114
rect 8701 -12080 8735 -12046
rect 8701 -12148 8735 -12114
rect 8801 -12080 8835 -12046
rect 8801 -12148 8835 -12114
rect 8998 -12073 9032 -12039
rect 8998 -12175 9032 -12141
rect 9262 -12073 9296 -12039
rect 9262 -12175 9296 -12141
rect 9458 -12073 9492 -12039
rect 9458 -12175 9492 -12141
rect 10090 -12073 10124 -12039
rect 10090 -12175 10124 -12141
rect 10378 -12073 10412 -12039
rect 10378 -12175 10412 -12141
rect 10642 -12073 10676 -12039
rect 10642 -12175 10676 -12141
rect 10761 -12081 10795 -12047
rect 10761 -12149 10795 -12115
rect 10859 -12080 10893 -12046
rect 10859 -12148 10893 -12114
rect 11015 -12081 11049 -12047
rect 11015 -12149 11049 -12115
rect 11119 -12080 11153 -12046
rect 11119 -12148 11153 -12114
rect 11277 -12080 11311 -12046
rect 11277 -12148 11311 -12114
rect 11377 -12080 11411 -12046
rect 11377 -12148 11411 -12114
rect 11666 -12073 11700 -12039
rect 11666 -12175 11700 -12141
rect 11930 -12073 11964 -12039
rect 11930 -12175 11964 -12141
rect 13690 -12073 13724 -12039
rect 13690 -12141 13724 -12107
rect 13776 -12081 13810 -12047
rect 13776 -12149 13810 -12115
rect 13862 -12073 13896 -12039
rect 13862 -12141 13896 -12107
rect 13948 -12089 13982 -12055
rect 13948 -12157 13982 -12123
rect 14034 -12073 14068 -12039
rect 14034 -12141 14068 -12107
rect 14120 -12117 14154 -12083
rect 14120 -12203 14154 -12169
rect 14206 -12097 14240 -12063
rect 14292 -12117 14326 -12083
rect 14292 -12203 14326 -12169
rect 14378 -12097 14412 -12063
rect 14464 -12117 14498 -12083
rect 14464 -12203 14498 -12169
rect 14550 -12097 14584 -12063
rect 14636 -12117 14670 -12083
rect 14636 -12203 14670 -12169
rect 14722 -12097 14756 -12063
rect 14807 -12117 14841 -12083
rect 14807 -12203 14841 -12169
rect 14893 -12097 14927 -12063
rect 14979 -12117 15013 -12083
rect 14979 -12203 15013 -12169
rect 15065 -12097 15099 -12063
rect 15151 -12117 15185 -12083
rect 15151 -12203 15185 -12169
rect 15237 -12097 15271 -12063
rect 15323 -12117 15357 -12083
rect 15323 -12203 15357 -12169
rect 15409 -12097 15443 -12063
rect 15622 -12073 15656 -12039
rect 15622 -12175 15656 -12141
rect 16622 -12073 16656 -12039
rect 16622 -12175 16656 -12141
rect -2962 -12907 -2928 -12873
rect -2962 -13009 -2928 -12975
rect -2330 -12907 -2296 -12873
rect -2330 -13009 -2296 -12975
rect -1582 -12907 -1548 -12873
rect -1582 -13009 -1548 -12975
rect -950 -12907 -916 -12873
rect -950 -13009 -916 -12975
rect -846 -12907 -812 -12873
rect -846 -13009 -812 -12975
rect -214 -12907 -180 -12873
rect -214 -13009 -180 -12975
rect -18 -12907 16 -12873
rect -18 -13009 16 -12975
rect 246 -12907 280 -12873
rect 246 -13009 280 -12975
rect 443 -12934 477 -12900
rect 443 -13002 477 -12968
rect 543 -12934 577 -12900
rect 543 -13002 577 -12968
rect 701 -12934 735 -12900
rect 701 -13002 735 -12968
rect 805 -12933 839 -12899
rect 805 -13001 839 -12967
rect 961 -12934 995 -12900
rect 961 -13002 995 -12968
rect 1059 -12933 1093 -12899
rect 1059 -13001 1093 -12967
rect 1270 -12907 1304 -12873
rect 1270 -13009 1304 -12975
rect 1534 -12907 1568 -12873
rect 1534 -13009 1568 -12975
rect 1730 -12907 1764 -12873
rect 1730 -13009 1764 -12975
rect 2362 -12907 2396 -12873
rect 2362 -13009 2396 -12975
rect 2558 -12907 2592 -12873
rect 2558 -13009 2592 -12975
rect 2822 -12907 2856 -12873
rect 2822 -13009 2856 -12975
rect 3019 -12934 3053 -12900
rect 3019 -13002 3053 -12968
rect 3119 -12934 3153 -12900
rect 3119 -13002 3153 -12968
rect 3277 -12934 3311 -12900
rect 3277 -13002 3311 -12968
rect 3381 -12933 3415 -12899
rect 3381 -13001 3415 -12967
rect 3537 -12934 3571 -12900
rect 3537 -13002 3571 -12968
rect 3635 -12933 3669 -12899
rect 3635 -13001 3669 -12967
rect 3846 -12907 3880 -12873
rect 3846 -13009 3880 -12975
rect 4110 -12907 4144 -12873
rect 4110 -13009 4144 -12975
rect 4306 -12907 4340 -12873
rect 4306 -13009 4340 -12975
rect 4938 -12907 4972 -12873
rect 4938 -13009 4972 -12975
rect 5134 -12907 5168 -12873
rect 5134 -13009 5168 -12975
rect 5398 -12907 5432 -12873
rect 5398 -13009 5432 -12975
rect 5595 -12934 5629 -12900
rect 5595 -13002 5629 -12968
rect 5695 -12934 5729 -12900
rect 5695 -13002 5729 -12968
rect 5853 -12934 5887 -12900
rect 5853 -13002 5887 -12968
rect 5957 -12933 5991 -12899
rect 5957 -13001 5991 -12967
rect 6113 -12934 6147 -12900
rect 6113 -13002 6147 -12968
rect 6211 -12933 6245 -12899
rect 6211 -13001 6245 -12967
rect 6422 -12907 6456 -12873
rect 6422 -13009 6456 -12975
rect 6686 -12907 6720 -12873
rect 6686 -13009 6720 -12975
rect 6882 -12907 6916 -12873
rect 6882 -13009 6916 -12975
rect 7514 -12907 7548 -12873
rect 7514 -13009 7548 -12975
rect 7710 -12907 7744 -12873
rect 7710 -13009 7744 -12975
rect 7974 -12907 8008 -12873
rect 7974 -13009 8008 -12975
rect 8171 -12934 8205 -12900
rect 8171 -13002 8205 -12968
rect 8271 -12934 8305 -12900
rect 8271 -13002 8305 -12968
rect 8429 -12934 8463 -12900
rect 8429 -13002 8463 -12968
rect 8533 -12933 8567 -12899
rect 8533 -13001 8567 -12967
rect 8689 -12934 8723 -12900
rect 8689 -13002 8723 -12968
rect 8787 -12933 8821 -12899
rect 8787 -13001 8821 -12967
rect 8998 -12907 9032 -12873
rect 8998 -13009 9032 -12975
rect 9262 -12907 9296 -12873
rect 9262 -13009 9296 -12975
rect 9458 -12907 9492 -12873
rect 9458 -13009 9492 -12975
rect 10090 -12907 10124 -12873
rect 10090 -13009 10124 -12975
rect 10378 -12907 10412 -12873
rect 10378 -13009 10412 -12975
rect 10642 -12907 10676 -12873
rect 10642 -13009 10676 -12975
rect 10747 -12934 10781 -12900
rect 10747 -13002 10781 -12968
rect 10847 -12934 10881 -12900
rect 10847 -13002 10881 -12968
rect 11005 -12934 11039 -12900
rect 11005 -13002 11039 -12968
rect 11109 -12933 11143 -12899
rect 11109 -13001 11143 -12967
rect 11265 -12934 11299 -12900
rect 11265 -13002 11299 -12968
rect 11363 -12933 11397 -12899
rect 11363 -13001 11397 -12967
rect 11666 -12907 11700 -12873
rect 11666 -13009 11700 -12975
rect 11930 -12907 11964 -12873
rect 11930 -13009 11964 -12975
rect 12502 -12934 12536 -12900
rect 12502 -13002 12536 -12968
rect 12588 -12907 12622 -12873
rect 12588 -12995 12622 -12961
rect 12674 -12934 12708 -12900
rect 12674 -13002 12708 -12968
rect 12760 -12907 12794 -12873
rect 12760 -12995 12794 -12961
rect 12846 -12934 12880 -12900
rect 12846 -13002 12880 -12968
rect 12932 -12907 12966 -12873
rect 12932 -12995 12966 -12961
rect 13018 -12934 13052 -12900
rect 13018 -13002 13052 -12968
rect 13230 -12907 13264 -12873
rect 13230 -13009 13264 -12975
rect 13494 -12907 13528 -12873
rect 13494 -13009 13528 -12975
rect 13690 -12941 13724 -12907
rect 13690 -13009 13724 -12975
rect 13776 -12933 13810 -12899
rect 13776 -13001 13810 -12967
rect 13862 -12941 13896 -12907
rect 13862 -13009 13896 -12975
rect 13948 -12925 13982 -12891
rect 13948 -12993 13982 -12959
rect 14034 -12941 14068 -12907
rect 14034 -13009 14068 -12975
rect 14120 -12879 14154 -12845
rect 14120 -12965 14154 -12931
rect 14206 -12985 14240 -12951
rect 14292 -12879 14326 -12845
rect 14292 -12965 14326 -12931
rect 14378 -12985 14412 -12951
rect 14464 -12879 14498 -12845
rect 14464 -12965 14498 -12931
rect 14550 -12985 14584 -12951
rect 14636 -12879 14670 -12845
rect 14636 -12965 14670 -12931
rect 14722 -12985 14756 -12951
rect 14807 -12879 14841 -12845
rect 14807 -12965 14841 -12931
rect 14893 -12985 14927 -12951
rect 14979 -12879 15013 -12845
rect 14979 -12965 15013 -12931
rect 15065 -12985 15099 -12951
rect 15151 -12879 15185 -12845
rect 15151 -12965 15185 -12931
rect 15237 -12985 15271 -12951
rect 15323 -12879 15357 -12845
rect 15323 -12965 15357 -12931
rect 15409 -12985 15443 -12951
rect 15622 -12907 15656 -12873
rect 15622 -13009 15656 -12975
rect 16622 -12907 16656 -12873
rect 16622 -13009 16656 -12975
rect -2962 -13161 -2928 -13127
rect -2962 -13263 -2928 -13229
rect -2330 -13161 -2296 -13127
rect -2330 -13263 -2296 -13229
rect -1582 -13161 -1548 -13127
rect -1582 -13263 -1548 -13229
rect -950 -13161 -916 -13127
rect -950 -13263 -916 -13229
rect -846 -13161 -812 -13127
rect -846 -13263 -812 -13229
rect -214 -13161 -180 -13127
rect -214 -13263 -180 -13229
rect -18 -13161 16 -13127
rect -18 -13263 16 -13229
rect 246 -13161 280 -13127
rect 246 -13263 280 -13229
rect 457 -13169 491 -13135
rect 457 -13237 491 -13203
rect 555 -13168 589 -13134
rect 555 -13236 589 -13202
rect 711 -13169 745 -13135
rect 711 -13237 745 -13203
rect 815 -13168 849 -13134
rect 815 -13236 849 -13202
rect 973 -13168 1007 -13134
rect 973 -13236 1007 -13202
rect 1073 -13168 1107 -13134
rect 1073 -13236 1107 -13202
rect 1270 -13161 1304 -13127
rect 1270 -13263 1304 -13229
rect 1534 -13161 1568 -13127
rect 1534 -13263 1568 -13229
rect 1730 -13161 1764 -13127
rect 1730 -13263 1764 -13229
rect 2362 -13161 2396 -13127
rect 2362 -13263 2396 -13229
rect 2558 -13161 2592 -13127
rect 2558 -13263 2592 -13229
rect 2822 -13161 2856 -13127
rect 2822 -13263 2856 -13229
rect 3033 -13169 3067 -13135
rect 3033 -13237 3067 -13203
rect 3131 -13168 3165 -13134
rect 3131 -13236 3165 -13202
rect 3287 -13169 3321 -13135
rect 3287 -13237 3321 -13203
rect 3391 -13168 3425 -13134
rect 3391 -13236 3425 -13202
rect 3549 -13168 3583 -13134
rect 3549 -13236 3583 -13202
rect 3649 -13168 3683 -13134
rect 3649 -13236 3683 -13202
rect 3846 -13161 3880 -13127
rect 3846 -13263 3880 -13229
rect 4110 -13161 4144 -13127
rect 4110 -13263 4144 -13229
rect 4306 -13161 4340 -13127
rect 4306 -13263 4340 -13229
rect 4938 -13161 4972 -13127
rect 4938 -13263 4972 -13229
rect 5134 -13161 5168 -13127
rect 5134 -13263 5168 -13229
rect 5398 -13161 5432 -13127
rect 5398 -13263 5432 -13229
rect 5609 -13169 5643 -13135
rect 5609 -13237 5643 -13203
rect 5707 -13168 5741 -13134
rect 5707 -13236 5741 -13202
rect 5863 -13169 5897 -13135
rect 5863 -13237 5897 -13203
rect 5967 -13168 6001 -13134
rect 5967 -13236 6001 -13202
rect 6125 -13168 6159 -13134
rect 6125 -13236 6159 -13202
rect 6225 -13168 6259 -13134
rect 6225 -13236 6259 -13202
rect 6422 -13161 6456 -13127
rect 6422 -13263 6456 -13229
rect 6686 -13161 6720 -13127
rect 6686 -13263 6720 -13229
rect 6882 -13161 6916 -13127
rect 6882 -13263 6916 -13229
rect 7514 -13161 7548 -13127
rect 7514 -13263 7548 -13229
rect 7710 -13161 7744 -13127
rect 7710 -13263 7744 -13229
rect 7974 -13161 8008 -13127
rect 7974 -13263 8008 -13229
rect 8185 -13169 8219 -13135
rect 8185 -13237 8219 -13203
rect 8283 -13168 8317 -13134
rect 8283 -13236 8317 -13202
rect 8439 -13169 8473 -13135
rect 8439 -13237 8473 -13203
rect 8543 -13168 8577 -13134
rect 8543 -13236 8577 -13202
rect 8701 -13168 8735 -13134
rect 8701 -13236 8735 -13202
rect 8801 -13168 8835 -13134
rect 8801 -13236 8835 -13202
rect 8998 -13161 9032 -13127
rect 8998 -13263 9032 -13229
rect 9262 -13161 9296 -13127
rect 9262 -13263 9296 -13229
rect 9458 -13161 9492 -13127
rect 9458 -13263 9492 -13229
rect 10090 -13161 10124 -13127
rect 10090 -13263 10124 -13229
rect 10378 -13161 10412 -13127
rect 10378 -13263 10412 -13229
rect 10642 -13161 10676 -13127
rect 10642 -13263 10676 -13229
rect 10761 -13169 10795 -13135
rect 10761 -13237 10795 -13203
rect 10859 -13168 10893 -13134
rect 10859 -13236 10893 -13202
rect 11015 -13169 11049 -13135
rect 11015 -13237 11049 -13203
rect 11119 -13168 11153 -13134
rect 11119 -13236 11153 -13202
rect 11277 -13168 11311 -13134
rect 11277 -13236 11311 -13202
rect 11377 -13168 11411 -13134
rect 11377 -13236 11411 -13202
rect 11666 -13161 11700 -13127
rect 11666 -13263 11700 -13229
rect 11930 -13161 11964 -13127
rect 11930 -13263 11964 -13229
rect 13690 -13161 13724 -13127
rect 13690 -13229 13724 -13195
rect 13776 -13169 13810 -13135
rect 13776 -13237 13810 -13203
rect 13862 -13161 13896 -13127
rect 13862 -13229 13896 -13195
rect 13948 -13177 13982 -13143
rect 13948 -13245 13982 -13211
rect 14034 -13161 14068 -13127
rect 14034 -13229 14068 -13195
rect 14120 -13205 14154 -13171
rect 14120 -13291 14154 -13257
rect 14206 -13185 14240 -13151
rect 14292 -13205 14326 -13171
rect 14292 -13291 14326 -13257
rect 14378 -13185 14412 -13151
rect 14464 -13205 14498 -13171
rect 14464 -13291 14498 -13257
rect 14550 -13185 14584 -13151
rect 14636 -13205 14670 -13171
rect 14636 -13291 14670 -13257
rect 14722 -13185 14756 -13151
rect 14807 -13205 14841 -13171
rect 14807 -13291 14841 -13257
rect 14893 -13185 14927 -13151
rect 14979 -13205 15013 -13171
rect 14979 -13291 15013 -13257
rect 15065 -13185 15099 -13151
rect 15151 -13205 15185 -13171
rect 15151 -13291 15185 -13257
rect 15237 -13185 15271 -13151
rect 15323 -13205 15357 -13171
rect 15323 -13291 15357 -13257
rect 15409 -13185 15443 -13151
rect 15622 -13161 15656 -13127
rect 15622 -13263 15656 -13229
rect 16622 -13161 16656 -13127
rect 16622 -13263 16656 -13229
rect -2962 -13995 -2928 -13961
rect -2962 -14097 -2928 -14063
rect -2330 -13995 -2296 -13961
rect -2330 -14097 -2296 -14063
rect -1398 -13995 -1364 -13961
rect -1398 -14097 -1364 -14063
rect -1134 -13995 -1100 -13961
rect -1134 -14097 -1100 -14063
rect -934 -13961 -900 -13927
rect -934 -14029 -900 -13995
rect -934 -14097 -900 -14063
rect -850 -13961 -816 -13927
rect -850 -14029 -816 -13995
rect -850 -14097 -816 -14063
rect -766 -13961 -732 -13927
rect -766 -14029 -732 -13995
rect -766 -14097 -732 -14063
rect -570 -13995 -536 -13961
rect -570 -14097 -536 -14063
rect -306 -13995 -272 -13961
rect -306 -14097 -272 -14063
rect -102 -14022 -68 -13988
rect -102 -14090 -68 -14056
rect -16 -13995 18 -13961
rect -16 -14083 18 -14049
rect 70 -14022 104 -13988
rect 70 -14090 104 -14056
rect 156 -13995 190 -13961
rect 156 -14083 190 -14049
rect 242 -14022 276 -13988
rect 242 -14090 276 -14056
rect 328 -13995 362 -13961
rect 328 -14083 362 -14049
rect 414 -14022 448 -13988
rect 414 -14090 448 -14056
rect 626 -13995 660 -13961
rect 626 -14097 660 -14063
rect 890 -13995 924 -13961
rect 890 -14097 924 -14063
rect 1086 -13995 1120 -13961
rect 1086 -14097 1120 -14063
rect 1170 -13995 1204 -13961
rect 1170 -14097 1204 -14063
rect 1254 -13995 1288 -13961
rect 1254 -14097 1288 -14063
rect 1454 -13995 1488 -13961
rect 1454 -14097 1488 -14063
rect 1718 -13995 1752 -13961
rect 1718 -14097 1752 -14063
rect 1914 -13995 1948 -13961
rect 1914 -14097 1948 -14063
rect 2178 -13995 2212 -13961
rect 2178 -14097 2212 -14063
rect 2375 -14022 2409 -13988
rect 2375 -14090 2409 -14056
rect 2475 -14022 2509 -13988
rect 2475 -14090 2509 -14056
rect 2633 -14022 2667 -13988
rect 2633 -14090 2667 -14056
rect 2737 -14021 2771 -13987
rect 2737 -14089 2771 -14055
rect 2893 -14022 2927 -13988
rect 2893 -14090 2927 -14056
rect 2991 -14021 3025 -13987
rect 2991 -14089 3025 -14055
rect 3202 -13995 3236 -13961
rect 3202 -14097 3236 -14063
rect 3466 -13995 3500 -13961
rect 3466 -14097 3500 -14063
rect 4398 -13995 4432 -13961
rect 4398 -14097 4432 -14063
rect 5398 -13995 5432 -13961
rect 5398 -14097 5432 -14063
rect 6422 -13995 6456 -13961
rect 6422 -14097 6456 -14063
rect 6686 -13995 6720 -13961
rect 6686 -14097 6720 -14063
rect 6883 -14022 6917 -13988
rect 6883 -14090 6917 -14056
rect 6983 -14022 7017 -13988
rect 6983 -14090 7017 -14056
rect 7141 -14022 7175 -13988
rect 7141 -14090 7175 -14056
rect 7245 -14021 7279 -13987
rect 7245 -14089 7279 -14055
rect 7401 -14022 7435 -13988
rect 7401 -14090 7435 -14056
rect 7499 -14021 7533 -13987
rect 7499 -14089 7533 -14055
rect 7710 -13995 7744 -13961
rect 7710 -14097 7744 -14063
rect 7974 -13995 8008 -13961
rect 7974 -14097 8008 -14063
rect 8171 -14022 8205 -13988
rect 8171 -14090 8205 -14056
rect 8271 -14022 8305 -13988
rect 8271 -14090 8305 -14056
rect 8429 -14022 8463 -13988
rect 8429 -14090 8463 -14056
rect 8533 -14021 8567 -13987
rect 8533 -14089 8567 -14055
rect 8689 -14022 8723 -13988
rect 8689 -14090 8723 -14056
rect 8787 -14021 8821 -13987
rect 8787 -14089 8821 -14055
rect 8998 -13995 9032 -13961
rect 8998 -14097 9032 -14063
rect 9262 -13995 9296 -13961
rect 9262 -14097 9296 -14063
rect 9459 -14022 9493 -13988
rect 9459 -14090 9493 -14056
rect 9559 -14022 9593 -13988
rect 9559 -14090 9593 -14056
rect 9717 -14022 9751 -13988
rect 9717 -14090 9751 -14056
rect 9821 -14021 9855 -13987
rect 9821 -14089 9855 -14055
rect 9977 -14022 10011 -13988
rect 9977 -14090 10011 -14056
rect 10075 -14021 10109 -13987
rect 10075 -14089 10109 -14055
rect 10286 -13995 10320 -13961
rect 10286 -14097 10320 -14063
rect 10550 -13995 10584 -13961
rect 10550 -14097 10584 -14063
rect 10746 -13961 10780 -13927
rect 10746 -14029 10780 -13995
rect 10746 -14097 10780 -14063
rect 10830 -13961 10864 -13927
rect 10830 -14029 10864 -13995
rect 10830 -14097 10864 -14063
rect 10914 -14029 10948 -13995
rect 10914 -14097 10948 -14063
rect 10998 -13961 11032 -13927
rect 10998 -14029 11032 -13995
rect 10998 -14097 11032 -14063
rect 11082 -14029 11116 -13995
rect 11082 -14097 11116 -14063
rect 11166 -13961 11200 -13927
rect 11166 -14029 11200 -13995
rect 11166 -14097 11200 -14063
rect 11250 -14029 11284 -13995
rect 11250 -14097 11284 -14063
rect 11334 -13961 11368 -13927
rect 11334 -14029 11368 -13995
rect 11334 -14097 11368 -14063
rect 11418 -14029 11452 -13995
rect 11418 -14097 11452 -14063
rect 11666 -13995 11700 -13961
rect 11666 -14097 11700 -14063
rect 11930 -13995 11964 -13961
rect 11930 -14097 11964 -14063
rect 13598 -13995 13632 -13961
rect 13598 -14097 13632 -14063
rect 14598 -13995 14632 -13961
rect 14598 -14097 14632 -14063
rect 14794 -13995 14828 -13961
rect 14794 -14097 14828 -14063
rect 15794 -13995 15828 -13961
rect 15794 -14097 15828 -14063
rect 15990 -13995 16024 -13961
rect 15990 -14097 16024 -14063
rect 16622 -13995 16656 -13961
rect 16622 -14097 16656 -14063
<< psubdiff >>
rect -2232 -411 -2198 -387
rect -2232 -492 -2198 -445
rect -1036 -411 -1002 -387
rect -1036 -492 -1002 -445
rect -668 -411 -634 -387
rect -668 -492 -634 -445
rect -208 -411 -174 -387
rect 528 -411 562 -387
rect -208 -492 -174 -445
rect 528 -492 562 -445
rect 988 -411 1022 -387
rect 1356 -411 1390 -387
rect 988 -492 1022 -445
rect 1356 -492 1390 -445
rect 1816 -411 1850 -387
rect 1816 -492 1850 -445
rect 2276 -411 2310 -387
rect 2276 -492 2310 -445
rect 3104 -411 3138 -387
rect 3104 -492 3138 -445
rect 3564 -411 3598 -387
rect 3564 -492 3598 -445
rect 6324 -411 6358 -387
rect 6324 -492 6358 -445
rect 6784 -411 6818 -387
rect 6784 -492 6818 -445
rect 7612 -411 7646 -387
rect 7612 -492 7646 -445
rect 8072 -411 8106 -387
rect 8072 -492 8106 -445
rect 8900 -411 8934 -387
rect 8900 -492 8934 -445
rect 9360 -411 9394 -387
rect 9360 -492 9394 -445
rect 10188 -411 10222 -387
rect 10188 -492 10222 -445
rect 10648 -411 10682 -387
rect 10648 -492 10682 -445
rect 11568 -411 11602 -387
rect 11568 -492 11602 -445
rect 13500 -411 13534 -387
rect 13500 -492 13534 -445
rect 14696 -411 14730 -387
rect 14696 -492 14730 -445
rect 15892 -411 15926 -387
rect 15892 -492 15926 -445
rect -2232 -667 -2198 -620
rect -2232 -725 -2198 -701
rect -116 -667 -82 -620
rect -116 -725 -82 -701
rect 344 -667 378 -620
rect 344 -725 378 -701
rect 1172 -667 1206 -620
rect 1172 -725 1206 -701
rect 1632 -667 1666 -620
rect 1632 -725 1666 -701
rect 2460 -667 2494 -620
rect 2460 -725 2494 -701
rect 2920 -667 2954 -620
rect 2920 -725 2954 -701
rect 3748 -667 3782 -620
rect 3748 -725 3782 -701
rect 4208 -667 4242 -620
rect 4208 -725 4242 -701
rect 5036 -667 5070 -620
rect 5036 -725 5070 -701
rect 5496 -667 5530 -620
rect 5496 -725 5530 -701
rect 6324 -667 6358 -620
rect 6324 -725 6358 -701
rect 6784 -667 6818 -620
rect 6784 -725 6818 -701
rect 7612 -667 7646 -620
rect 7612 -725 7646 -701
rect 8072 -667 8106 -620
rect 8072 -725 8106 -701
rect 8900 -667 8934 -620
rect 8900 -725 8934 -701
rect 9360 -667 9394 -620
rect 9360 -725 9394 -701
rect 10188 -667 10222 -620
rect 10188 -725 10222 -701
rect 11476 -667 11510 -620
rect 11476 -725 11510 -701
rect 13592 -667 13626 -620
rect 15524 -667 15558 -620
rect 13592 -725 13626 -701
rect 15524 -725 15558 -701
rect -2232 -1499 -2198 -1475
rect -2232 -1580 -2198 -1533
rect -116 -1499 -82 -1475
rect -116 -1580 -82 -1533
rect 344 -1499 378 -1475
rect 344 -1580 378 -1533
rect 1172 -1499 1206 -1475
rect 1172 -1580 1206 -1533
rect 1632 -1499 1666 -1475
rect 1632 -1580 1666 -1533
rect 2460 -1499 2494 -1475
rect 2460 -1580 2494 -1533
rect 2920 -1499 2954 -1475
rect 2920 -1580 2954 -1533
rect 3748 -1499 3782 -1475
rect 3748 -1580 3782 -1533
rect 4208 -1499 4242 -1475
rect 4208 -1580 4242 -1533
rect 5036 -1499 5070 -1475
rect 5036 -1580 5070 -1533
rect 5496 -1499 5530 -1475
rect 5496 -1580 5530 -1533
rect 6324 -1499 6358 -1475
rect 6324 -1580 6358 -1533
rect 6784 -1499 6818 -1475
rect 6784 -1580 6818 -1533
rect 7612 -1499 7646 -1475
rect 7612 -1580 7646 -1533
rect 8072 -1499 8106 -1475
rect 8072 -1580 8106 -1533
rect 8900 -1499 8934 -1475
rect 8900 -1580 8934 -1533
rect 9360 -1499 9394 -1475
rect 9360 -1580 9394 -1533
rect 10188 -1499 10222 -1475
rect 10188 -1580 10222 -1533
rect 11476 -1499 11510 -1475
rect 11476 -1580 11510 -1533
rect 12396 -1499 12430 -1475
rect 13132 -1499 13166 -1475
rect 12396 -1580 12430 -1533
rect 13132 -1580 13166 -1533
rect 13592 -1499 13626 -1475
rect 15524 -1499 15558 -1475
rect 13592 -1580 13626 -1533
rect 15524 -1580 15558 -1533
rect -2232 -1755 -2198 -1708
rect -2232 -1813 -2198 -1789
rect -116 -1755 -82 -1708
rect -116 -1813 -82 -1789
rect 344 -1755 378 -1708
rect 344 -1813 378 -1789
rect 1172 -1755 1206 -1708
rect 1172 -1813 1206 -1789
rect 1632 -1755 1666 -1708
rect 1632 -1813 1666 -1789
rect 2460 -1755 2494 -1708
rect 2460 -1813 2494 -1789
rect 2920 -1755 2954 -1708
rect 2920 -1813 2954 -1789
rect 3748 -1755 3782 -1708
rect 3748 -1813 3782 -1789
rect 4208 -1755 4242 -1708
rect 4208 -1813 4242 -1789
rect 5036 -1755 5070 -1708
rect 5036 -1813 5070 -1789
rect 5496 -1755 5530 -1708
rect 5496 -1813 5530 -1789
rect 6324 -1755 6358 -1708
rect 6324 -1813 6358 -1789
rect 6784 -1755 6818 -1708
rect 6784 -1813 6818 -1789
rect 7612 -1755 7646 -1708
rect 7612 -1813 7646 -1789
rect 8072 -1755 8106 -1708
rect 8072 -1813 8106 -1789
rect 8900 -1755 8934 -1708
rect 8900 -1813 8934 -1789
rect 9360 -1755 9394 -1708
rect 9360 -1813 9394 -1789
rect 10188 -1755 10222 -1708
rect 10188 -1813 10222 -1789
rect 11476 -1755 11510 -1708
rect 11476 -1813 11510 -1789
rect 13592 -1755 13626 -1708
rect 15524 -1755 15558 -1708
rect 13592 -1813 13626 -1789
rect 15524 -1813 15558 -1789
rect -2232 -2587 -2198 -2563
rect -2232 -2668 -2198 -2621
rect -116 -2587 -82 -2563
rect -116 -2668 -82 -2621
rect 344 -2587 378 -2563
rect 344 -2668 378 -2621
rect 1172 -2587 1206 -2563
rect 1172 -2668 1206 -2621
rect 1632 -2587 1666 -2563
rect 1632 -2668 1666 -2621
rect 2460 -2587 2494 -2563
rect 2460 -2668 2494 -2621
rect 2920 -2587 2954 -2563
rect 2920 -2668 2954 -2621
rect 3748 -2587 3782 -2563
rect 3748 -2668 3782 -2621
rect 4208 -2587 4242 -2563
rect 4208 -2668 4242 -2621
rect 5036 -2587 5070 -2563
rect 5036 -2668 5070 -2621
rect 5496 -2587 5530 -2563
rect 5496 -2668 5530 -2621
rect 6324 -2587 6358 -2563
rect 6324 -2668 6358 -2621
rect 6784 -2587 6818 -2563
rect 6784 -2668 6818 -2621
rect 7612 -2587 7646 -2563
rect 7612 -2668 7646 -2621
rect 8072 -2587 8106 -2563
rect 8072 -2668 8106 -2621
rect 8900 -2587 8934 -2563
rect 8900 -2668 8934 -2621
rect 9360 -2587 9394 -2563
rect 9360 -2668 9394 -2621
rect 10188 -2587 10222 -2563
rect 10188 -2668 10222 -2621
rect 11476 -2587 11510 -2563
rect 11476 -2668 11510 -2621
rect 12396 -2587 12430 -2563
rect 13132 -2587 13166 -2563
rect 12396 -2668 12430 -2621
rect 13132 -2668 13166 -2621
rect 13592 -2587 13626 -2563
rect 15524 -2587 15558 -2563
rect 13592 -2668 13626 -2621
rect 15524 -2668 15558 -2621
rect -2232 -2843 -2198 -2796
rect -1680 -2843 -1646 -2796
rect -2232 -2901 -2198 -2877
rect -1680 -2901 -1646 -2877
rect -116 -2843 -82 -2796
rect -116 -2901 -82 -2877
rect 344 -2843 378 -2796
rect 344 -2901 378 -2877
rect 1172 -2843 1206 -2796
rect 1172 -2901 1206 -2877
rect 1632 -2843 1666 -2796
rect 1632 -2901 1666 -2877
rect 2460 -2843 2494 -2796
rect 2460 -2901 2494 -2877
rect 2920 -2843 2954 -2796
rect 2920 -2901 2954 -2877
rect 3748 -2843 3782 -2796
rect 3748 -2901 3782 -2877
rect 4208 -2843 4242 -2796
rect 4208 -2901 4242 -2877
rect 5036 -2843 5070 -2796
rect 5036 -2901 5070 -2877
rect 5496 -2843 5530 -2796
rect 5496 -2901 5530 -2877
rect 6324 -2843 6358 -2796
rect 6324 -2901 6358 -2877
rect 6784 -2843 6818 -2796
rect 6784 -2901 6818 -2877
rect 7612 -2843 7646 -2796
rect 7612 -2901 7646 -2877
rect 8072 -2843 8106 -2796
rect 8072 -2901 8106 -2877
rect 8900 -2843 8934 -2796
rect 8900 -2901 8934 -2877
rect 9360 -2843 9394 -2796
rect 9360 -2901 9394 -2877
rect 10188 -2843 10222 -2796
rect 10188 -2901 10222 -2877
rect 11476 -2843 11510 -2796
rect 11476 -2901 11510 -2877
rect 13500 -2843 13534 -2796
rect 13500 -2901 13534 -2877
rect 14696 -2843 14730 -2796
rect 14696 -2901 14730 -2877
rect 15892 -2843 15926 -2796
rect 15892 -2901 15926 -2877
rect -2232 -3675 -2198 -3651
rect -2232 -3756 -2198 -3709
rect -116 -3675 -82 -3651
rect -116 -3756 -82 -3709
rect 344 -3675 378 -3651
rect 344 -3756 378 -3709
rect 1172 -3675 1206 -3651
rect 1172 -3756 1206 -3709
rect 1632 -3675 1666 -3651
rect 1632 -3756 1666 -3709
rect 2460 -3675 2494 -3651
rect 2460 -3756 2494 -3709
rect 2920 -3675 2954 -3651
rect 2920 -3756 2954 -3709
rect 3748 -3675 3782 -3651
rect 3748 -3756 3782 -3709
rect 4208 -3675 4242 -3651
rect 4208 -3756 4242 -3709
rect 5036 -3675 5070 -3651
rect 5036 -3756 5070 -3709
rect 5496 -3675 5530 -3651
rect 5496 -3756 5530 -3709
rect 6324 -3675 6358 -3651
rect 6324 -3756 6358 -3709
rect 6784 -3675 6818 -3651
rect 6784 -3756 6818 -3709
rect 7612 -3675 7646 -3651
rect 7612 -3756 7646 -3709
rect 8072 -3675 8106 -3651
rect 8072 -3756 8106 -3709
rect 8900 -3675 8934 -3651
rect 8900 -3756 8934 -3709
rect 9360 -3675 9394 -3651
rect 9360 -3756 9394 -3709
rect 10188 -3675 10222 -3651
rect 10188 -3756 10222 -3709
rect 11476 -3675 11510 -3651
rect 11476 -3756 11510 -3709
rect 13500 -3675 13534 -3651
rect 13500 -3756 13534 -3709
rect 14696 -3675 14730 -3651
rect 14696 -3756 14730 -3709
rect 15892 -3675 15926 -3651
rect 15892 -3756 15926 -3709
rect -2232 -3931 -2198 -3884
rect -2232 -3989 -2198 -3965
rect -116 -3931 -82 -3884
rect -116 -3989 -82 -3965
rect 344 -3931 378 -3884
rect 344 -3989 378 -3965
rect 1172 -3931 1206 -3884
rect 1172 -3989 1206 -3965
rect 1632 -3931 1666 -3884
rect 1632 -3989 1666 -3965
rect 2460 -3931 2494 -3884
rect 2460 -3989 2494 -3965
rect 2920 -3931 2954 -3884
rect 2920 -3989 2954 -3965
rect 3748 -3931 3782 -3884
rect 3748 -3989 3782 -3965
rect 4208 -3931 4242 -3884
rect 4208 -3989 4242 -3965
rect 5036 -3931 5070 -3884
rect 5036 -3989 5070 -3965
rect 5496 -3931 5530 -3884
rect 5496 -3989 5530 -3965
rect 6324 -3931 6358 -3884
rect 6324 -3989 6358 -3965
rect 6784 -3931 6818 -3884
rect 6784 -3989 6818 -3965
rect 7612 -3931 7646 -3884
rect 7612 -3989 7646 -3965
rect 8072 -3931 8106 -3884
rect 8072 -3989 8106 -3965
rect 8900 -3931 8934 -3884
rect 8900 -3989 8934 -3965
rect 9360 -3931 9394 -3884
rect 9360 -3989 9394 -3965
rect 10188 -3931 10222 -3884
rect 10188 -3989 10222 -3965
rect 11476 -3931 11510 -3884
rect 11476 -3989 11510 -3965
rect 12396 -3931 12430 -3884
rect 13132 -3931 13166 -3884
rect 12396 -3989 12430 -3965
rect 13132 -3989 13166 -3965
rect 13592 -3931 13626 -3884
rect 15524 -3931 15558 -3884
rect 13592 -3989 13626 -3965
rect 15524 -3989 15558 -3965
rect -2232 -4763 -2198 -4739
rect -2232 -4844 -2198 -4797
rect -116 -4763 -82 -4739
rect -116 -4844 -82 -4797
rect 344 -4763 378 -4739
rect 344 -4844 378 -4797
rect 1172 -4763 1206 -4739
rect 1172 -4844 1206 -4797
rect 1632 -4763 1666 -4739
rect 1632 -4844 1666 -4797
rect 2460 -4763 2494 -4739
rect 2460 -4844 2494 -4797
rect 2920 -4763 2954 -4739
rect 2920 -4844 2954 -4797
rect 3748 -4763 3782 -4739
rect 3748 -4844 3782 -4797
rect 4208 -4763 4242 -4739
rect 4208 -4844 4242 -4797
rect 5036 -4763 5070 -4739
rect 5036 -4844 5070 -4797
rect 5496 -4763 5530 -4739
rect 5496 -4844 5530 -4797
rect 6324 -4763 6358 -4739
rect 6324 -4844 6358 -4797
rect 6784 -4763 6818 -4739
rect 6784 -4844 6818 -4797
rect 7612 -4763 7646 -4739
rect 7612 -4844 7646 -4797
rect 8072 -4763 8106 -4739
rect 8072 -4844 8106 -4797
rect 8900 -4763 8934 -4739
rect 8900 -4844 8934 -4797
rect 9360 -4763 9394 -4739
rect 9360 -4844 9394 -4797
rect 10188 -4763 10222 -4739
rect 10188 -4844 10222 -4797
rect 11476 -4763 11510 -4739
rect 11476 -4844 11510 -4797
rect 13592 -4763 13626 -4739
rect 15524 -4763 15558 -4739
rect 13592 -4844 13626 -4797
rect 15524 -4844 15558 -4797
rect -2232 -5019 -2198 -4972
rect -2232 -5077 -2198 -5053
rect -116 -5019 -82 -4972
rect -116 -5077 -82 -5053
rect 344 -5019 378 -4972
rect 344 -5077 378 -5053
rect 1172 -5019 1206 -4972
rect 1172 -5077 1206 -5053
rect 1632 -5019 1666 -4972
rect 1632 -5077 1666 -5053
rect 2460 -5019 2494 -4972
rect 2460 -5077 2494 -5053
rect 2920 -5019 2954 -4972
rect 2920 -5077 2954 -5053
rect 3748 -5019 3782 -4972
rect 3748 -5077 3782 -5053
rect 4208 -5019 4242 -4972
rect 4208 -5077 4242 -5053
rect 5036 -5019 5070 -4972
rect 5036 -5077 5070 -5053
rect 5496 -5019 5530 -4972
rect 5496 -5077 5530 -5053
rect 6324 -5019 6358 -4972
rect 6324 -5077 6358 -5053
rect 6784 -5019 6818 -4972
rect 6784 -5077 6818 -5053
rect 7612 -5019 7646 -4972
rect 7612 -5077 7646 -5053
rect 8072 -5019 8106 -4972
rect 8072 -5077 8106 -5053
rect 8900 -5019 8934 -4972
rect 8900 -5077 8934 -5053
rect 9360 -5019 9394 -4972
rect 9360 -5077 9394 -5053
rect 10188 -5019 10222 -4972
rect 10188 -5077 10222 -5053
rect 11476 -5019 11510 -4972
rect 11476 -5077 11510 -5053
rect 12396 -5019 12430 -4972
rect 13132 -5019 13166 -4972
rect 12396 -5077 12430 -5053
rect 13132 -5077 13166 -5053
rect 13592 -5019 13626 -4972
rect 15524 -5019 15558 -4972
rect 13592 -5077 13626 -5053
rect 15524 -5077 15558 -5053
rect -2232 -5851 -2198 -5827
rect -2232 -5932 -2198 -5885
rect -116 -5851 -82 -5827
rect -116 -5932 -82 -5885
rect 344 -5851 378 -5827
rect 344 -5932 378 -5885
rect 1172 -5851 1206 -5827
rect 1172 -5932 1206 -5885
rect 1632 -5851 1666 -5827
rect 1632 -5932 1666 -5885
rect 2460 -5851 2494 -5827
rect 2460 -5932 2494 -5885
rect 2920 -5851 2954 -5827
rect 2920 -5932 2954 -5885
rect 3748 -5851 3782 -5827
rect 3748 -5932 3782 -5885
rect 4208 -5851 4242 -5827
rect 4208 -5932 4242 -5885
rect 5036 -5851 5070 -5827
rect 5036 -5932 5070 -5885
rect 5496 -5851 5530 -5827
rect 5496 -5932 5530 -5885
rect 6324 -5851 6358 -5827
rect 6324 -5932 6358 -5885
rect 6784 -5851 6818 -5827
rect 6784 -5932 6818 -5885
rect 7612 -5851 7646 -5827
rect 7612 -5932 7646 -5885
rect 8072 -5851 8106 -5827
rect 8072 -5932 8106 -5885
rect 8900 -5851 8934 -5827
rect 8900 -5932 8934 -5885
rect 9360 -5851 9394 -5827
rect 9360 -5932 9394 -5885
rect 10188 -5851 10222 -5827
rect 10188 -5932 10222 -5885
rect 11476 -5851 11510 -5827
rect 11476 -5932 11510 -5885
rect 13592 -5851 13626 -5827
rect 15524 -5851 15558 -5827
rect 13592 -5932 13626 -5885
rect 15524 -5932 15558 -5885
rect -2232 -6107 -2198 -6060
rect -2232 -6165 -2198 -6141
rect -1036 -6107 -1002 -6060
rect -1036 -6165 -1002 -6141
rect -668 -6107 -634 -6060
rect -668 -6165 -634 -6141
rect -208 -6107 -174 -6060
rect 528 -6107 562 -6060
rect -208 -6165 -174 -6141
rect 528 -6165 562 -6141
rect 988 -6107 1022 -6060
rect 1356 -6107 1390 -6060
rect 988 -6165 1022 -6141
rect 1356 -6165 1390 -6141
rect 1816 -6107 1850 -6060
rect 1816 -6165 1850 -6141
rect 2276 -6107 2310 -6060
rect 2276 -6165 2310 -6141
rect 3104 -6107 3138 -6060
rect 3104 -6165 3138 -6141
rect 3564 -6107 3598 -6060
rect 3564 -6165 3598 -6141
rect 6324 -6107 6358 -6060
rect 6324 -6165 6358 -6141
rect 6784 -6107 6818 -6060
rect 6784 -6165 6818 -6141
rect 7612 -6107 7646 -6060
rect 7612 -6165 7646 -6141
rect 8072 -6107 8106 -6060
rect 8072 -6165 8106 -6141
rect 8900 -6107 8934 -6060
rect 8900 -6165 8934 -6141
rect 9360 -6107 9394 -6060
rect 9360 -6165 9394 -6141
rect 10188 -6107 10222 -6060
rect 10188 -6165 10222 -6141
rect 10648 -6107 10682 -6060
rect 10648 -6165 10682 -6141
rect 11568 -6107 11602 -6060
rect 11568 -6165 11602 -6141
rect 13500 -6107 13534 -6060
rect 13500 -6165 13534 -6141
rect 14696 -6107 14730 -6060
rect 14696 -6165 14730 -6141
rect 15892 -6107 15926 -6060
rect 15892 -6165 15926 -6141
rect -2692 -6939 -2658 -6915
rect -2692 -7020 -2658 -6973
rect -116 -6939 -82 -6915
rect -116 -7020 -82 -6973
rect 1448 -6939 1482 -6915
rect 1448 -7020 1482 -6973
rect 3012 -6939 3046 -6915
rect 3012 -7020 3046 -6973
rect 4576 -6939 4610 -6915
rect 4576 -7020 4610 -6973
rect 6140 -6939 6174 -6915
rect 6140 -7020 6174 -6973
rect 7704 -6939 7738 -6915
rect 7704 -7020 7738 -6973
rect 9268 -6939 9302 -6915
rect 9268 -7020 9302 -6973
rect 15892 -6939 15926 -6915
rect 15892 -7020 15926 -6973
rect -2232 -7195 -2198 -7148
rect -2232 -7253 -2198 -7229
rect -116 -7195 -82 -7148
rect -116 -7253 -82 -7229
rect 1448 -7195 1482 -7148
rect 1448 -7253 1482 -7229
rect 2828 -7195 2862 -7148
rect 3196 -7195 3230 -7148
rect 2828 -7253 2862 -7229
rect 3196 -7253 3230 -7229
rect 3656 -7195 3690 -7148
rect 3656 -7253 3690 -7229
rect 4024 -7195 4058 -7148
rect 4024 -7253 4058 -7229
rect 4484 -7195 4518 -7148
rect 4484 -7253 4518 -7229
rect 5404 -7195 5438 -7148
rect 5404 -7253 5438 -7229
rect 5864 -7195 5898 -7148
rect 5864 -7253 5898 -7229
rect 7704 -7195 7738 -7148
rect 7704 -7253 7738 -7229
rect 9268 -7195 9302 -7148
rect 9268 -7253 9302 -7229
rect 15892 -7195 15926 -7148
rect 15892 -7253 15926 -7229
rect -2232 -8027 -2198 -8003
rect -2232 -8108 -2198 -8061
rect -1036 -8027 -1002 -8003
rect -1036 -8108 -1002 -8061
rect -668 -8027 -634 -8003
rect -668 -8108 -634 -8061
rect -208 -8027 -174 -8003
rect 528 -8027 562 -8003
rect -208 -8108 -174 -8061
rect 528 -8108 562 -8061
rect 988 -8027 1022 -8003
rect 1356 -8027 1390 -8003
rect 988 -8108 1022 -8061
rect 1356 -8108 1390 -8061
rect 1816 -8027 1850 -8003
rect 1816 -8108 1850 -8061
rect 2276 -8027 2310 -8003
rect 2276 -8108 2310 -8061
rect 3104 -8027 3138 -8003
rect 3104 -8108 3138 -8061
rect 3564 -8027 3598 -8003
rect 3564 -8108 3598 -8061
rect 6324 -8027 6358 -8003
rect 6324 -8108 6358 -8061
rect 6784 -8027 6818 -8003
rect 6784 -8108 6818 -8061
rect 7612 -8027 7646 -8003
rect 7612 -8108 7646 -8061
rect 8072 -8027 8106 -8003
rect 8072 -8108 8106 -8061
rect 8900 -8027 8934 -8003
rect 8900 -8108 8934 -8061
rect 9360 -8027 9394 -8003
rect 9360 -8108 9394 -8061
rect 10188 -8027 10222 -8003
rect 10188 -8108 10222 -8061
rect 10648 -8027 10682 -8003
rect 10648 -8108 10682 -8061
rect 11568 -8027 11602 -8003
rect 11568 -8108 11602 -8061
rect 13500 -8027 13534 -8003
rect 13500 -8108 13534 -8061
rect 14696 -8027 14730 -8003
rect 14696 -8108 14730 -8061
rect 15892 -8027 15926 -8003
rect 15892 -8108 15926 -8061
rect -2232 -8283 -2198 -8236
rect -2232 -8341 -2198 -8317
rect -116 -8283 -82 -8236
rect -116 -8341 -82 -8317
rect 344 -8283 378 -8236
rect 344 -8341 378 -8317
rect 1172 -8283 1206 -8236
rect 1172 -8341 1206 -8317
rect 1632 -8283 1666 -8236
rect 1632 -8341 1666 -8317
rect 2460 -8283 2494 -8236
rect 2460 -8341 2494 -8317
rect 2920 -8283 2954 -8236
rect 2920 -8341 2954 -8317
rect 3748 -8283 3782 -8236
rect 3748 -8341 3782 -8317
rect 4208 -8283 4242 -8236
rect 4208 -8341 4242 -8317
rect 5036 -8283 5070 -8236
rect 5036 -8341 5070 -8317
rect 5496 -8283 5530 -8236
rect 5496 -8341 5530 -8317
rect 6324 -8283 6358 -8236
rect 6324 -8341 6358 -8317
rect 6784 -8283 6818 -8236
rect 6784 -8341 6818 -8317
rect 7612 -8283 7646 -8236
rect 7612 -8341 7646 -8317
rect 8072 -8283 8106 -8236
rect 8072 -8341 8106 -8317
rect 8900 -8283 8934 -8236
rect 8900 -8341 8934 -8317
rect 9360 -8283 9394 -8236
rect 9360 -8341 9394 -8317
rect 10188 -8283 10222 -8236
rect 10188 -8341 10222 -8317
rect 11476 -8283 11510 -8236
rect 11476 -8341 11510 -8317
rect 13592 -8283 13626 -8236
rect 15524 -8283 15558 -8236
rect 13592 -8341 13626 -8317
rect 15524 -8341 15558 -8317
rect -2232 -9115 -2198 -9091
rect -2232 -9196 -2198 -9149
rect -116 -9115 -82 -9091
rect -116 -9196 -82 -9149
rect 344 -9115 378 -9091
rect 344 -9196 378 -9149
rect 1172 -9115 1206 -9091
rect 1172 -9196 1206 -9149
rect 1632 -9115 1666 -9091
rect 1632 -9196 1666 -9149
rect 2460 -9115 2494 -9091
rect 2460 -9196 2494 -9149
rect 2920 -9115 2954 -9091
rect 2920 -9196 2954 -9149
rect 3748 -9115 3782 -9091
rect 3748 -9196 3782 -9149
rect 4208 -9115 4242 -9091
rect 4208 -9196 4242 -9149
rect 5036 -9115 5070 -9091
rect 5036 -9196 5070 -9149
rect 5496 -9115 5530 -9091
rect 5496 -9196 5530 -9149
rect 6324 -9115 6358 -9091
rect 6324 -9196 6358 -9149
rect 6784 -9115 6818 -9091
rect 6784 -9196 6818 -9149
rect 7612 -9115 7646 -9091
rect 7612 -9196 7646 -9149
rect 8072 -9115 8106 -9091
rect 8072 -9196 8106 -9149
rect 8900 -9115 8934 -9091
rect 8900 -9196 8934 -9149
rect 9360 -9115 9394 -9091
rect 9360 -9196 9394 -9149
rect 10188 -9115 10222 -9091
rect 10188 -9196 10222 -9149
rect 11476 -9115 11510 -9091
rect 11476 -9196 11510 -9149
rect 12396 -9115 12430 -9091
rect 13132 -9115 13166 -9091
rect 12396 -9196 12430 -9149
rect 13132 -9196 13166 -9149
rect 13592 -9115 13626 -9091
rect 15524 -9115 15558 -9091
rect 13592 -9196 13626 -9149
rect 15524 -9196 15558 -9149
rect -2232 -9371 -2198 -9324
rect -2232 -9429 -2198 -9405
rect -116 -9371 -82 -9324
rect -116 -9429 -82 -9405
rect 344 -9371 378 -9324
rect 344 -9429 378 -9405
rect 1172 -9371 1206 -9324
rect 1172 -9429 1206 -9405
rect 1632 -9371 1666 -9324
rect 1632 -9429 1666 -9405
rect 2460 -9371 2494 -9324
rect 2460 -9429 2494 -9405
rect 2920 -9371 2954 -9324
rect 2920 -9429 2954 -9405
rect 3748 -9371 3782 -9324
rect 3748 -9429 3782 -9405
rect 4208 -9371 4242 -9324
rect 4208 -9429 4242 -9405
rect 5036 -9371 5070 -9324
rect 5036 -9429 5070 -9405
rect 5496 -9371 5530 -9324
rect 5496 -9429 5530 -9405
rect 6324 -9371 6358 -9324
rect 6324 -9429 6358 -9405
rect 6784 -9371 6818 -9324
rect 6784 -9429 6818 -9405
rect 7612 -9371 7646 -9324
rect 7612 -9429 7646 -9405
rect 8072 -9371 8106 -9324
rect 8072 -9429 8106 -9405
rect 8900 -9371 8934 -9324
rect 8900 -9429 8934 -9405
rect 9360 -9371 9394 -9324
rect 9360 -9429 9394 -9405
rect 10188 -9371 10222 -9324
rect 10188 -9429 10222 -9405
rect 11476 -9371 11510 -9324
rect 11476 -9429 11510 -9405
rect 13592 -9371 13626 -9324
rect 15524 -9371 15558 -9324
rect 13592 -9429 13626 -9405
rect 15524 -9429 15558 -9405
rect -2232 -10203 -2198 -10179
rect -2232 -10284 -2198 -10237
rect -116 -10203 -82 -10179
rect -116 -10284 -82 -10237
rect 344 -10203 378 -10179
rect 344 -10284 378 -10237
rect 1172 -10203 1206 -10179
rect 1172 -10284 1206 -10237
rect 1632 -10203 1666 -10179
rect 1632 -10284 1666 -10237
rect 2460 -10203 2494 -10179
rect 2460 -10284 2494 -10237
rect 2920 -10203 2954 -10179
rect 2920 -10284 2954 -10237
rect 3748 -10203 3782 -10179
rect 3748 -10284 3782 -10237
rect 4208 -10203 4242 -10179
rect 4208 -10284 4242 -10237
rect 5036 -10203 5070 -10179
rect 5036 -10284 5070 -10237
rect 5496 -10203 5530 -10179
rect 5496 -10284 5530 -10237
rect 6324 -10203 6358 -10179
rect 6324 -10284 6358 -10237
rect 6784 -10203 6818 -10179
rect 6784 -10284 6818 -10237
rect 7612 -10203 7646 -10179
rect 7612 -10284 7646 -10237
rect 8072 -10203 8106 -10179
rect 8072 -10284 8106 -10237
rect 8900 -10203 8934 -10179
rect 8900 -10284 8934 -10237
rect 9360 -10203 9394 -10179
rect 9360 -10284 9394 -10237
rect 10188 -10203 10222 -10179
rect 10188 -10284 10222 -10237
rect 11476 -10203 11510 -10179
rect 11476 -10284 11510 -10237
rect 12396 -10203 12430 -10179
rect 13132 -10203 13166 -10179
rect 12396 -10284 12430 -10237
rect 13132 -10284 13166 -10237
rect 13592 -10203 13626 -10179
rect 15524 -10203 15558 -10179
rect 13592 -10284 13626 -10237
rect 15524 -10284 15558 -10237
rect -2232 -10459 -2198 -10412
rect -1680 -10459 -1646 -10412
rect -2232 -10517 -2198 -10493
rect -1680 -10517 -1646 -10493
rect -116 -10459 -82 -10412
rect -116 -10517 -82 -10493
rect 344 -10459 378 -10412
rect 344 -10517 378 -10493
rect 1172 -10459 1206 -10412
rect 1172 -10517 1206 -10493
rect 1632 -10459 1666 -10412
rect 1632 -10517 1666 -10493
rect 2460 -10459 2494 -10412
rect 2460 -10517 2494 -10493
rect 2920 -10459 2954 -10412
rect 2920 -10517 2954 -10493
rect 3748 -10459 3782 -10412
rect 3748 -10517 3782 -10493
rect 4208 -10459 4242 -10412
rect 4208 -10517 4242 -10493
rect 5036 -10459 5070 -10412
rect 5036 -10517 5070 -10493
rect 5496 -10459 5530 -10412
rect 5496 -10517 5530 -10493
rect 6324 -10459 6358 -10412
rect 6324 -10517 6358 -10493
rect 6784 -10459 6818 -10412
rect 6784 -10517 6818 -10493
rect 7612 -10459 7646 -10412
rect 7612 -10517 7646 -10493
rect 8072 -10459 8106 -10412
rect 8072 -10517 8106 -10493
rect 8900 -10459 8934 -10412
rect 8900 -10517 8934 -10493
rect 9360 -10459 9394 -10412
rect 9360 -10517 9394 -10493
rect 10188 -10459 10222 -10412
rect 10188 -10517 10222 -10493
rect 11476 -10459 11510 -10412
rect 11476 -10517 11510 -10493
rect 13500 -10459 13534 -10412
rect 13500 -10517 13534 -10493
rect 14696 -10459 14730 -10412
rect 14696 -10517 14730 -10493
rect 15892 -10459 15926 -10412
rect 15892 -10517 15926 -10493
rect -2232 -11291 -2198 -11267
rect -2232 -11372 -2198 -11325
rect -116 -11291 -82 -11267
rect -116 -11372 -82 -11325
rect 344 -11291 378 -11267
rect 344 -11372 378 -11325
rect 1172 -11291 1206 -11267
rect 1172 -11372 1206 -11325
rect 1632 -11291 1666 -11267
rect 1632 -11372 1666 -11325
rect 2460 -11291 2494 -11267
rect 2460 -11372 2494 -11325
rect 2920 -11291 2954 -11267
rect 2920 -11372 2954 -11325
rect 3748 -11291 3782 -11267
rect 3748 -11372 3782 -11325
rect 4208 -11291 4242 -11267
rect 4208 -11372 4242 -11325
rect 5036 -11291 5070 -11267
rect 5036 -11372 5070 -11325
rect 5496 -11291 5530 -11267
rect 5496 -11372 5530 -11325
rect 6324 -11291 6358 -11267
rect 6324 -11372 6358 -11325
rect 6784 -11291 6818 -11267
rect 6784 -11372 6818 -11325
rect 7612 -11291 7646 -11267
rect 7612 -11372 7646 -11325
rect 8072 -11291 8106 -11267
rect 8072 -11372 8106 -11325
rect 8900 -11291 8934 -11267
rect 8900 -11372 8934 -11325
rect 9360 -11291 9394 -11267
rect 9360 -11372 9394 -11325
rect 10188 -11291 10222 -11267
rect 10188 -11372 10222 -11325
rect 11476 -11291 11510 -11267
rect 11476 -11372 11510 -11325
rect 13500 -11291 13534 -11267
rect 13500 -11372 13534 -11325
rect 14696 -11291 14730 -11267
rect 14696 -11372 14730 -11325
rect 15892 -11291 15926 -11267
rect 15892 -11372 15926 -11325
rect -2232 -11547 -2198 -11500
rect -2232 -11605 -2198 -11581
rect -116 -11547 -82 -11500
rect -116 -11605 -82 -11581
rect 344 -11547 378 -11500
rect 344 -11605 378 -11581
rect 1172 -11547 1206 -11500
rect 1172 -11605 1206 -11581
rect 1632 -11547 1666 -11500
rect 1632 -11605 1666 -11581
rect 2460 -11547 2494 -11500
rect 2460 -11605 2494 -11581
rect 2920 -11547 2954 -11500
rect 2920 -11605 2954 -11581
rect 3748 -11547 3782 -11500
rect 3748 -11605 3782 -11581
rect 4208 -11547 4242 -11500
rect 4208 -11605 4242 -11581
rect 5036 -11547 5070 -11500
rect 5036 -11605 5070 -11581
rect 5496 -11547 5530 -11500
rect 5496 -11605 5530 -11581
rect 6324 -11547 6358 -11500
rect 6324 -11605 6358 -11581
rect 6784 -11547 6818 -11500
rect 6784 -11605 6818 -11581
rect 7612 -11547 7646 -11500
rect 7612 -11605 7646 -11581
rect 8072 -11547 8106 -11500
rect 8072 -11605 8106 -11581
rect 8900 -11547 8934 -11500
rect 8900 -11605 8934 -11581
rect 9360 -11547 9394 -11500
rect 9360 -11605 9394 -11581
rect 10188 -11547 10222 -11500
rect 10188 -11605 10222 -11581
rect 11476 -11547 11510 -11500
rect 11476 -11605 11510 -11581
rect 12396 -11547 12430 -11500
rect 13132 -11547 13166 -11500
rect 12396 -11605 12430 -11581
rect 13132 -11605 13166 -11581
rect 13592 -11547 13626 -11500
rect 15524 -11547 15558 -11500
rect 13592 -11605 13626 -11581
rect 15524 -11605 15558 -11581
rect -2232 -12379 -2198 -12355
rect -2232 -12460 -2198 -12413
rect -116 -12379 -82 -12355
rect -116 -12460 -82 -12413
rect 344 -12379 378 -12355
rect 344 -12460 378 -12413
rect 1172 -12379 1206 -12355
rect 1172 -12460 1206 -12413
rect 1632 -12379 1666 -12355
rect 1632 -12460 1666 -12413
rect 2460 -12379 2494 -12355
rect 2460 -12460 2494 -12413
rect 2920 -12379 2954 -12355
rect 2920 -12460 2954 -12413
rect 3748 -12379 3782 -12355
rect 3748 -12460 3782 -12413
rect 4208 -12379 4242 -12355
rect 4208 -12460 4242 -12413
rect 5036 -12379 5070 -12355
rect 5036 -12460 5070 -12413
rect 5496 -12379 5530 -12355
rect 5496 -12460 5530 -12413
rect 6324 -12379 6358 -12355
rect 6324 -12460 6358 -12413
rect 6784 -12379 6818 -12355
rect 6784 -12460 6818 -12413
rect 7612 -12379 7646 -12355
rect 7612 -12460 7646 -12413
rect 8072 -12379 8106 -12355
rect 8072 -12460 8106 -12413
rect 8900 -12379 8934 -12355
rect 8900 -12460 8934 -12413
rect 9360 -12379 9394 -12355
rect 9360 -12460 9394 -12413
rect 10188 -12379 10222 -12355
rect 10188 -12460 10222 -12413
rect 11476 -12379 11510 -12355
rect 11476 -12460 11510 -12413
rect 13592 -12379 13626 -12355
rect 15524 -12379 15558 -12355
rect 13592 -12460 13626 -12413
rect 15524 -12460 15558 -12413
rect -2232 -12635 -2198 -12588
rect -2232 -12693 -2198 -12669
rect -116 -12635 -82 -12588
rect -116 -12693 -82 -12669
rect 344 -12635 378 -12588
rect 344 -12693 378 -12669
rect 1172 -12635 1206 -12588
rect 1172 -12693 1206 -12669
rect 1632 -12635 1666 -12588
rect 1632 -12693 1666 -12669
rect 2460 -12635 2494 -12588
rect 2460 -12693 2494 -12669
rect 2920 -12635 2954 -12588
rect 2920 -12693 2954 -12669
rect 3748 -12635 3782 -12588
rect 3748 -12693 3782 -12669
rect 4208 -12635 4242 -12588
rect 4208 -12693 4242 -12669
rect 5036 -12635 5070 -12588
rect 5036 -12693 5070 -12669
rect 5496 -12635 5530 -12588
rect 5496 -12693 5530 -12669
rect 6324 -12635 6358 -12588
rect 6324 -12693 6358 -12669
rect 6784 -12635 6818 -12588
rect 6784 -12693 6818 -12669
rect 7612 -12635 7646 -12588
rect 7612 -12693 7646 -12669
rect 8072 -12635 8106 -12588
rect 8072 -12693 8106 -12669
rect 8900 -12635 8934 -12588
rect 8900 -12693 8934 -12669
rect 9360 -12635 9394 -12588
rect 9360 -12693 9394 -12669
rect 10188 -12635 10222 -12588
rect 10188 -12693 10222 -12669
rect 11476 -12635 11510 -12588
rect 11476 -12693 11510 -12669
rect 12396 -12635 12430 -12588
rect 13132 -12635 13166 -12588
rect 12396 -12693 12430 -12669
rect 13132 -12693 13166 -12669
rect 13592 -12635 13626 -12588
rect 15524 -12635 15558 -12588
rect 13592 -12693 13626 -12669
rect 15524 -12693 15558 -12669
rect -2232 -13467 -2198 -13443
rect -2232 -13548 -2198 -13501
rect -116 -13467 -82 -13443
rect -116 -13548 -82 -13501
rect 344 -13467 378 -13443
rect 344 -13548 378 -13501
rect 1172 -13467 1206 -13443
rect 1172 -13548 1206 -13501
rect 1632 -13467 1666 -13443
rect 1632 -13548 1666 -13501
rect 2460 -13467 2494 -13443
rect 2460 -13548 2494 -13501
rect 2920 -13467 2954 -13443
rect 2920 -13548 2954 -13501
rect 3748 -13467 3782 -13443
rect 3748 -13548 3782 -13501
rect 4208 -13467 4242 -13443
rect 4208 -13548 4242 -13501
rect 5036 -13467 5070 -13443
rect 5036 -13548 5070 -13501
rect 5496 -13467 5530 -13443
rect 5496 -13548 5530 -13501
rect 6324 -13467 6358 -13443
rect 6324 -13548 6358 -13501
rect 6784 -13467 6818 -13443
rect 6784 -13548 6818 -13501
rect 7612 -13467 7646 -13443
rect 7612 -13548 7646 -13501
rect 8072 -13467 8106 -13443
rect 8072 -13548 8106 -13501
rect 8900 -13467 8934 -13443
rect 8900 -13548 8934 -13501
rect 9360 -13467 9394 -13443
rect 9360 -13548 9394 -13501
rect 10188 -13467 10222 -13443
rect 10188 -13548 10222 -13501
rect 11476 -13467 11510 -13443
rect 11476 -13548 11510 -13501
rect 13592 -13467 13626 -13443
rect 15524 -13467 15558 -13443
rect 13592 -13548 13626 -13501
rect 15524 -13548 15558 -13501
rect -2232 -13723 -2198 -13676
rect -2232 -13781 -2198 -13757
rect -1036 -13723 -1002 -13676
rect -1036 -13781 -1002 -13757
rect -668 -13723 -634 -13676
rect -668 -13781 -634 -13757
rect -208 -13723 -174 -13676
rect 528 -13723 562 -13676
rect -208 -13781 -174 -13757
rect 528 -13781 562 -13757
rect 988 -13723 1022 -13676
rect 1356 -13723 1390 -13676
rect 988 -13781 1022 -13757
rect 1356 -13781 1390 -13757
rect 1816 -13723 1850 -13676
rect 1816 -13781 1850 -13757
rect 2276 -13723 2310 -13676
rect 2276 -13781 2310 -13757
rect 3104 -13723 3138 -13676
rect 3104 -13781 3138 -13757
rect 3564 -13723 3598 -13676
rect 3564 -13781 3598 -13757
rect 6324 -13723 6358 -13676
rect 6324 -13781 6358 -13757
rect 6784 -13723 6818 -13676
rect 6784 -13781 6818 -13757
rect 7612 -13723 7646 -13676
rect 7612 -13781 7646 -13757
rect 8072 -13723 8106 -13676
rect 8072 -13781 8106 -13757
rect 8900 -13723 8934 -13676
rect 8900 -13781 8934 -13757
rect 9360 -13723 9394 -13676
rect 9360 -13781 9394 -13757
rect 10188 -13723 10222 -13676
rect 10188 -13781 10222 -13757
rect 10648 -13723 10682 -13676
rect 10648 -13781 10682 -13757
rect 11568 -13723 11602 -13676
rect 11568 -13781 11602 -13757
rect 13500 -13723 13534 -13676
rect 13500 -13781 13534 -13757
rect 14696 -13723 14730 -13676
rect 14696 -13781 14730 -13757
rect 15892 -13723 15926 -13676
rect 15892 -13781 15926 -13757
<< nsubdiff >>
rect -2232 -100 -2198 -76
rect -2232 -193 -2198 -134
rect -2232 -251 -2198 -227
rect -1036 -100 -1002 -76
rect -1036 -193 -1002 -134
rect -1036 -251 -1002 -227
rect -668 -100 -634 -76
rect -668 -193 -634 -134
rect -668 -251 -634 -227
rect -208 -100 -174 -76
rect -208 -193 -174 -134
rect -208 -251 -174 -227
rect 528 -100 562 -76
rect 528 -193 562 -134
rect 528 -251 562 -227
rect 988 -100 1022 -76
rect 988 -193 1022 -134
rect 1356 -100 1390 -76
rect 1356 -193 1390 -134
rect 988 -251 1022 -227
rect 1356 -251 1390 -227
rect 1816 -100 1850 -76
rect 1816 -193 1850 -134
rect 1816 -251 1850 -227
rect 2276 -100 2310 -76
rect 2276 -193 2310 -134
rect 2276 -251 2310 -227
rect 3104 -100 3138 -76
rect 3104 -193 3138 -134
rect 3104 -251 3138 -227
rect 3564 -100 3598 -76
rect 3564 -193 3598 -134
rect 3564 -251 3598 -227
rect 6324 -100 6358 -76
rect 6324 -193 6358 -134
rect 6324 -251 6358 -227
rect 6784 -100 6818 -76
rect 6784 -193 6818 -134
rect 6784 -251 6818 -227
rect 7612 -100 7646 -76
rect 7612 -193 7646 -134
rect 7612 -251 7646 -227
rect 8072 -100 8106 -76
rect 8072 -193 8106 -134
rect 8072 -251 8106 -227
rect 8900 -100 8934 -76
rect 8900 -193 8934 -134
rect 8900 -251 8934 -227
rect 9360 -100 9394 -76
rect 9360 -193 9394 -134
rect 9360 -251 9394 -227
rect 10188 -100 10222 -76
rect 10188 -193 10222 -134
rect 10188 -251 10222 -227
rect 10648 -100 10682 -76
rect 10648 -193 10682 -134
rect 10648 -251 10682 -227
rect 11568 -100 11602 -76
rect 11568 -193 11602 -134
rect 11568 -251 11602 -227
rect 13500 -100 13534 -76
rect 13500 -193 13534 -134
rect 13500 -251 13534 -227
rect 14696 -100 14730 -76
rect 14696 -193 14730 -134
rect 14696 -251 14730 -227
rect 15892 -100 15926 -76
rect 15892 -193 15926 -134
rect 15892 -251 15926 -227
rect -2232 -885 -2198 -861
rect -2232 -978 -2198 -919
rect -2232 -1036 -2198 -1012
rect -116 -885 -82 -861
rect -116 -978 -82 -919
rect -116 -1036 -82 -1012
rect 344 -885 378 -861
rect 344 -978 378 -919
rect 344 -1036 378 -1012
rect 1172 -885 1206 -861
rect 1172 -978 1206 -919
rect 1172 -1036 1206 -1012
rect 1632 -885 1666 -861
rect 1632 -978 1666 -919
rect 1632 -1036 1666 -1012
rect 2460 -885 2494 -861
rect 2460 -978 2494 -919
rect 2460 -1036 2494 -1012
rect 2920 -885 2954 -861
rect 2920 -978 2954 -919
rect 2920 -1036 2954 -1012
rect 3748 -885 3782 -861
rect 3748 -978 3782 -919
rect 3748 -1036 3782 -1012
rect 4208 -885 4242 -861
rect 4208 -978 4242 -919
rect 4208 -1036 4242 -1012
rect 5036 -885 5070 -861
rect 5036 -978 5070 -919
rect 5036 -1036 5070 -1012
rect 5496 -885 5530 -861
rect 5496 -978 5530 -919
rect 5496 -1036 5530 -1012
rect 6324 -885 6358 -861
rect 6324 -978 6358 -919
rect 6324 -1036 6358 -1012
rect 6784 -885 6818 -861
rect 6784 -978 6818 -919
rect 6784 -1036 6818 -1012
rect 7612 -885 7646 -861
rect 7612 -978 7646 -919
rect 7612 -1036 7646 -1012
rect 8072 -885 8106 -861
rect 8072 -978 8106 -919
rect 8072 -1036 8106 -1012
rect 8900 -885 8934 -861
rect 8900 -978 8934 -919
rect 8900 -1036 8934 -1012
rect 9360 -885 9394 -861
rect 9360 -978 9394 -919
rect 9360 -1036 9394 -1012
rect 10188 -885 10222 -861
rect 10188 -978 10222 -919
rect 10188 -1036 10222 -1012
rect 11476 -885 11510 -861
rect 11476 -978 11510 -919
rect 11476 -1036 11510 -1012
rect 13592 -885 13626 -861
rect 13592 -978 13626 -919
rect 13592 -1036 13626 -1012
rect 15524 -885 15558 -861
rect 15524 -978 15558 -919
rect 15524 -1036 15558 -1012
rect -2232 -1188 -2198 -1164
rect -2232 -1281 -2198 -1222
rect -2232 -1339 -2198 -1315
rect -116 -1188 -82 -1164
rect -116 -1281 -82 -1222
rect -116 -1339 -82 -1315
rect 344 -1188 378 -1164
rect 344 -1281 378 -1222
rect 344 -1339 378 -1315
rect 1172 -1188 1206 -1164
rect 1172 -1281 1206 -1222
rect 1172 -1339 1206 -1315
rect 1632 -1188 1666 -1164
rect 1632 -1281 1666 -1222
rect 1632 -1339 1666 -1315
rect 2460 -1188 2494 -1164
rect 2460 -1281 2494 -1222
rect 2460 -1339 2494 -1315
rect 2920 -1188 2954 -1164
rect 2920 -1281 2954 -1222
rect 2920 -1339 2954 -1315
rect 3748 -1188 3782 -1164
rect 3748 -1281 3782 -1222
rect 3748 -1339 3782 -1315
rect 4208 -1188 4242 -1164
rect 4208 -1281 4242 -1222
rect 4208 -1339 4242 -1315
rect 5036 -1188 5070 -1164
rect 5036 -1281 5070 -1222
rect 5036 -1339 5070 -1315
rect 5496 -1188 5530 -1164
rect 5496 -1281 5530 -1222
rect 5496 -1339 5530 -1315
rect 6324 -1188 6358 -1164
rect 6324 -1281 6358 -1222
rect 6324 -1339 6358 -1315
rect 6784 -1188 6818 -1164
rect 6784 -1281 6818 -1222
rect 6784 -1339 6818 -1315
rect 7612 -1188 7646 -1164
rect 7612 -1281 7646 -1222
rect 7612 -1339 7646 -1315
rect 8072 -1188 8106 -1164
rect 8072 -1281 8106 -1222
rect 8072 -1339 8106 -1315
rect 8900 -1188 8934 -1164
rect 8900 -1281 8934 -1222
rect 8900 -1339 8934 -1315
rect 9360 -1188 9394 -1164
rect 9360 -1281 9394 -1222
rect 9360 -1339 9394 -1315
rect 10188 -1188 10222 -1164
rect 10188 -1281 10222 -1222
rect 10188 -1339 10222 -1315
rect 11476 -1188 11510 -1164
rect 11476 -1281 11510 -1222
rect 11476 -1339 11510 -1315
rect 12396 -1188 12430 -1164
rect 12396 -1281 12430 -1222
rect 12396 -1339 12430 -1315
rect 13132 -1188 13166 -1164
rect 13132 -1281 13166 -1222
rect 13132 -1339 13166 -1315
rect 13592 -1188 13626 -1164
rect 13592 -1281 13626 -1222
rect 13592 -1339 13626 -1315
rect 15524 -1188 15558 -1164
rect 15524 -1281 15558 -1222
rect 15524 -1339 15558 -1315
rect -2232 -1973 -2198 -1949
rect -2232 -2066 -2198 -2007
rect -2232 -2124 -2198 -2100
rect -116 -1973 -82 -1949
rect -116 -2066 -82 -2007
rect -116 -2124 -82 -2100
rect 344 -1973 378 -1949
rect 344 -2066 378 -2007
rect 344 -2124 378 -2100
rect 1172 -1973 1206 -1949
rect 1172 -2066 1206 -2007
rect 1172 -2124 1206 -2100
rect 1632 -1973 1666 -1949
rect 1632 -2066 1666 -2007
rect 1632 -2124 1666 -2100
rect 2460 -1973 2494 -1949
rect 2460 -2066 2494 -2007
rect 2460 -2124 2494 -2100
rect 2920 -1973 2954 -1949
rect 2920 -2066 2954 -2007
rect 2920 -2124 2954 -2100
rect 3748 -1973 3782 -1949
rect 3748 -2066 3782 -2007
rect 3748 -2124 3782 -2100
rect 4208 -1973 4242 -1949
rect 4208 -2066 4242 -2007
rect 4208 -2124 4242 -2100
rect 5036 -1973 5070 -1949
rect 5036 -2066 5070 -2007
rect 5036 -2124 5070 -2100
rect 5496 -1973 5530 -1949
rect 5496 -2066 5530 -2007
rect 5496 -2124 5530 -2100
rect 6324 -1973 6358 -1949
rect 6324 -2066 6358 -2007
rect 6324 -2124 6358 -2100
rect 6784 -1973 6818 -1949
rect 6784 -2066 6818 -2007
rect 6784 -2124 6818 -2100
rect 7612 -1973 7646 -1949
rect 7612 -2066 7646 -2007
rect 7612 -2124 7646 -2100
rect 8072 -1973 8106 -1949
rect 8072 -2066 8106 -2007
rect 8072 -2124 8106 -2100
rect 8900 -1973 8934 -1949
rect 8900 -2066 8934 -2007
rect 8900 -2124 8934 -2100
rect 9360 -1973 9394 -1949
rect 9360 -2066 9394 -2007
rect 9360 -2124 9394 -2100
rect 10188 -1973 10222 -1949
rect 10188 -2066 10222 -2007
rect 10188 -2124 10222 -2100
rect 11476 -1973 11510 -1949
rect 11476 -2066 11510 -2007
rect 11476 -2124 11510 -2100
rect 13592 -1973 13626 -1949
rect 13592 -2066 13626 -2007
rect 13592 -2124 13626 -2100
rect 15524 -1973 15558 -1949
rect 15524 -2066 15558 -2007
rect 15524 -2124 15558 -2100
rect -2232 -2276 -2198 -2252
rect -2232 -2369 -2198 -2310
rect -2232 -2427 -2198 -2403
rect -116 -2276 -82 -2252
rect -116 -2369 -82 -2310
rect -116 -2427 -82 -2403
rect 344 -2276 378 -2252
rect 344 -2369 378 -2310
rect 344 -2427 378 -2403
rect 1172 -2276 1206 -2252
rect 1172 -2369 1206 -2310
rect 1172 -2427 1206 -2403
rect 1632 -2276 1666 -2252
rect 1632 -2369 1666 -2310
rect 1632 -2427 1666 -2403
rect 2460 -2276 2494 -2252
rect 2460 -2369 2494 -2310
rect 2460 -2427 2494 -2403
rect 2920 -2276 2954 -2252
rect 2920 -2369 2954 -2310
rect 2920 -2427 2954 -2403
rect 3748 -2276 3782 -2252
rect 3748 -2369 3782 -2310
rect 3748 -2427 3782 -2403
rect 4208 -2276 4242 -2252
rect 4208 -2369 4242 -2310
rect 4208 -2427 4242 -2403
rect 5036 -2276 5070 -2252
rect 5036 -2369 5070 -2310
rect 5036 -2427 5070 -2403
rect 5496 -2276 5530 -2252
rect 5496 -2369 5530 -2310
rect 5496 -2427 5530 -2403
rect 6324 -2276 6358 -2252
rect 6324 -2369 6358 -2310
rect 6324 -2427 6358 -2403
rect 6784 -2276 6818 -2252
rect 6784 -2369 6818 -2310
rect 6784 -2427 6818 -2403
rect 7612 -2276 7646 -2252
rect 7612 -2369 7646 -2310
rect 7612 -2427 7646 -2403
rect 8072 -2276 8106 -2252
rect 8072 -2369 8106 -2310
rect 8072 -2427 8106 -2403
rect 8900 -2276 8934 -2252
rect 8900 -2369 8934 -2310
rect 8900 -2427 8934 -2403
rect 9360 -2276 9394 -2252
rect 9360 -2369 9394 -2310
rect 9360 -2427 9394 -2403
rect 10188 -2276 10222 -2252
rect 10188 -2369 10222 -2310
rect 10188 -2427 10222 -2403
rect 11476 -2276 11510 -2252
rect 11476 -2369 11510 -2310
rect 11476 -2427 11510 -2403
rect 12396 -2276 12430 -2252
rect 12396 -2369 12430 -2310
rect 12396 -2427 12430 -2403
rect 13132 -2276 13166 -2252
rect 13132 -2369 13166 -2310
rect 13132 -2427 13166 -2403
rect 13592 -2276 13626 -2252
rect 13592 -2369 13626 -2310
rect 13592 -2427 13626 -2403
rect 15524 -2276 15558 -2252
rect 15524 -2369 15558 -2310
rect 15524 -2427 15558 -2403
rect -2232 -3061 -2198 -3037
rect -1680 -3061 -1646 -3037
rect -2232 -3154 -2198 -3095
rect -2232 -3212 -2198 -3188
rect -1680 -3154 -1646 -3095
rect -1680 -3212 -1646 -3188
rect -116 -3061 -82 -3037
rect -116 -3154 -82 -3095
rect -116 -3212 -82 -3188
rect 344 -3061 378 -3037
rect 344 -3154 378 -3095
rect 344 -3212 378 -3188
rect 1172 -3061 1206 -3037
rect 1172 -3154 1206 -3095
rect 1172 -3212 1206 -3188
rect 1632 -3061 1666 -3037
rect 1632 -3154 1666 -3095
rect 1632 -3212 1666 -3188
rect 2460 -3061 2494 -3037
rect 2460 -3154 2494 -3095
rect 2460 -3212 2494 -3188
rect 2920 -3061 2954 -3037
rect 2920 -3154 2954 -3095
rect 2920 -3212 2954 -3188
rect 3748 -3061 3782 -3037
rect 3748 -3154 3782 -3095
rect 3748 -3212 3782 -3188
rect 4208 -3061 4242 -3037
rect 4208 -3154 4242 -3095
rect 4208 -3212 4242 -3188
rect 5036 -3061 5070 -3037
rect 5036 -3154 5070 -3095
rect 5036 -3212 5070 -3188
rect 5496 -3061 5530 -3037
rect 5496 -3154 5530 -3095
rect 5496 -3212 5530 -3188
rect 6324 -3061 6358 -3037
rect 6324 -3154 6358 -3095
rect 6324 -3212 6358 -3188
rect 6784 -3061 6818 -3037
rect 6784 -3154 6818 -3095
rect 6784 -3212 6818 -3188
rect 7612 -3061 7646 -3037
rect 7612 -3154 7646 -3095
rect 7612 -3212 7646 -3188
rect 8072 -3061 8106 -3037
rect 8072 -3154 8106 -3095
rect 8072 -3212 8106 -3188
rect 8900 -3061 8934 -3037
rect 8900 -3154 8934 -3095
rect 8900 -3212 8934 -3188
rect 9360 -3061 9394 -3037
rect 9360 -3154 9394 -3095
rect 9360 -3212 9394 -3188
rect 10188 -3061 10222 -3037
rect 10188 -3154 10222 -3095
rect 10188 -3212 10222 -3188
rect 11476 -3061 11510 -3037
rect 11476 -3154 11510 -3095
rect 11476 -3212 11510 -3188
rect 13500 -3061 13534 -3037
rect 13500 -3154 13534 -3095
rect 13500 -3212 13534 -3188
rect 14696 -3061 14730 -3037
rect 14696 -3154 14730 -3095
rect 14696 -3212 14730 -3188
rect 15892 -3061 15926 -3037
rect 15892 -3154 15926 -3095
rect 15892 -3212 15926 -3188
rect -2232 -3364 -2198 -3340
rect -2232 -3457 -2198 -3398
rect -2232 -3515 -2198 -3491
rect -116 -3364 -82 -3340
rect -116 -3457 -82 -3398
rect -116 -3515 -82 -3491
rect 344 -3364 378 -3340
rect 344 -3457 378 -3398
rect 344 -3515 378 -3491
rect 1172 -3364 1206 -3340
rect 1172 -3457 1206 -3398
rect 1172 -3515 1206 -3491
rect 1632 -3364 1666 -3340
rect 1632 -3457 1666 -3398
rect 1632 -3515 1666 -3491
rect 2460 -3364 2494 -3340
rect 2460 -3457 2494 -3398
rect 2460 -3515 2494 -3491
rect 2920 -3364 2954 -3340
rect 2920 -3457 2954 -3398
rect 2920 -3515 2954 -3491
rect 3748 -3364 3782 -3340
rect 3748 -3457 3782 -3398
rect 3748 -3515 3782 -3491
rect 4208 -3364 4242 -3340
rect 4208 -3457 4242 -3398
rect 4208 -3515 4242 -3491
rect 5036 -3364 5070 -3340
rect 5036 -3457 5070 -3398
rect 5036 -3515 5070 -3491
rect 5496 -3364 5530 -3340
rect 5496 -3457 5530 -3398
rect 5496 -3515 5530 -3491
rect 6324 -3364 6358 -3340
rect 6324 -3457 6358 -3398
rect 6324 -3515 6358 -3491
rect 6784 -3364 6818 -3340
rect 6784 -3457 6818 -3398
rect 6784 -3515 6818 -3491
rect 7612 -3364 7646 -3340
rect 7612 -3457 7646 -3398
rect 7612 -3515 7646 -3491
rect 8072 -3364 8106 -3340
rect 8072 -3457 8106 -3398
rect 8072 -3515 8106 -3491
rect 8900 -3364 8934 -3340
rect 8900 -3457 8934 -3398
rect 8900 -3515 8934 -3491
rect 9360 -3364 9394 -3340
rect 9360 -3457 9394 -3398
rect 9360 -3515 9394 -3491
rect 10188 -3364 10222 -3340
rect 10188 -3457 10222 -3398
rect 10188 -3515 10222 -3491
rect 11476 -3364 11510 -3340
rect 11476 -3457 11510 -3398
rect 11476 -3515 11510 -3491
rect 13500 -3364 13534 -3340
rect 13500 -3457 13534 -3398
rect 13500 -3515 13534 -3491
rect 14696 -3364 14730 -3340
rect 14696 -3457 14730 -3398
rect 14696 -3515 14730 -3491
rect 15892 -3364 15926 -3340
rect 15892 -3457 15926 -3398
rect 15892 -3515 15926 -3491
rect -2232 -4149 -2198 -4125
rect -2232 -4242 -2198 -4183
rect -2232 -4300 -2198 -4276
rect -116 -4149 -82 -4125
rect -116 -4242 -82 -4183
rect -116 -4300 -82 -4276
rect 344 -4149 378 -4125
rect 344 -4242 378 -4183
rect 344 -4300 378 -4276
rect 1172 -4149 1206 -4125
rect 1172 -4242 1206 -4183
rect 1172 -4300 1206 -4276
rect 1632 -4149 1666 -4125
rect 1632 -4242 1666 -4183
rect 1632 -4300 1666 -4276
rect 2460 -4149 2494 -4125
rect 2460 -4242 2494 -4183
rect 2460 -4300 2494 -4276
rect 2920 -4149 2954 -4125
rect 2920 -4242 2954 -4183
rect 2920 -4300 2954 -4276
rect 3748 -4149 3782 -4125
rect 3748 -4242 3782 -4183
rect 3748 -4300 3782 -4276
rect 4208 -4149 4242 -4125
rect 4208 -4242 4242 -4183
rect 4208 -4300 4242 -4276
rect 5036 -4149 5070 -4125
rect 5036 -4242 5070 -4183
rect 5036 -4300 5070 -4276
rect 5496 -4149 5530 -4125
rect 5496 -4242 5530 -4183
rect 5496 -4300 5530 -4276
rect 6324 -4149 6358 -4125
rect 6324 -4242 6358 -4183
rect 6324 -4300 6358 -4276
rect 6784 -4149 6818 -4125
rect 6784 -4242 6818 -4183
rect 6784 -4300 6818 -4276
rect 7612 -4149 7646 -4125
rect 7612 -4242 7646 -4183
rect 7612 -4300 7646 -4276
rect 8072 -4149 8106 -4125
rect 8072 -4242 8106 -4183
rect 8072 -4300 8106 -4276
rect 8900 -4149 8934 -4125
rect 8900 -4242 8934 -4183
rect 8900 -4300 8934 -4276
rect 9360 -4149 9394 -4125
rect 9360 -4242 9394 -4183
rect 9360 -4300 9394 -4276
rect 10188 -4149 10222 -4125
rect 10188 -4242 10222 -4183
rect 10188 -4300 10222 -4276
rect 11476 -4149 11510 -4125
rect 11476 -4242 11510 -4183
rect 11476 -4300 11510 -4276
rect 12396 -4149 12430 -4125
rect 12396 -4242 12430 -4183
rect 12396 -4300 12430 -4276
rect 13132 -4149 13166 -4125
rect 13132 -4242 13166 -4183
rect 13132 -4300 13166 -4276
rect 13592 -4149 13626 -4125
rect 13592 -4242 13626 -4183
rect 13592 -4300 13626 -4276
rect 15524 -4149 15558 -4125
rect 15524 -4242 15558 -4183
rect 15524 -4300 15558 -4276
rect -2232 -4452 -2198 -4428
rect -2232 -4545 -2198 -4486
rect -2232 -4603 -2198 -4579
rect -116 -4452 -82 -4428
rect -116 -4545 -82 -4486
rect -116 -4603 -82 -4579
rect 344 -4452 378 -4428
rect 344 -4545 378 -4486
rect 344 -4603 378 -4579
rect 1172 -4452 1206 -4428
rect 1172 -4545 1206 -4486
rect 1172 -4603 1206 -4579
rect 1632 -4452 1666 -4428
rect 1632 -4545 1666 -4486
rect 1632 -4603 1666 -4579
rect 2460 -4452 2494 -4428
rect 2460 -4545 2494 -4486
rect 2460 -4603 2494 -4579
rect 2920 -4452 2954 -4428
rect 2920 -4545 2954 -4486
rect 2920 -4603 2954 -4579
rect 3748 -4452 3782 -4428
rect 3748 -4545 3782 -4486
rect 3748 -4603 3782 -4579
rect 4208 -4452 4242 -4428
rect 4208 -4545 4242 -4486
rect 4208 -4603 4242 -4579
rect 5036 -4452 5070 -4428
rect 5036 -4545 5070 -4486
rect 5036 -4603 5070 -4579
rect 5496 -4452 5530 -4428
rect 5496 -4545 5530 -4486
rect 5496 -4603 5530 -4579
rect 6324 -4452 6358 -4428
rect 6324 -4545 6358 -4486
rect 6324 -4603 6358 -4579
rect 6784 -4452 6818 -4428
rect 6784 -4545 6818 -4486
rect 6784 -4603 6818 -4579
rect 7612 -4452 7646 -4428
rect 7612 -4545 7646 -4486
rect 7612 -4603 7646 -4579
rect 8072 -4452 8106 -4428
rect 8072 -4545 8106 -4486
rect 8072 -4603 8106 -4579
rect 8900 -4452 8934 -4428
rect 8900 -4545 8934 -4486
rect 8900 -4603 8934 -4579
rect 9360 -4452 9394 -4428
rect 9360 -4545 9394 -4486
rect 9360 -4603 9394 -4579
rect 10188 -4452 10222 -4428
rect 10188 -4545 10222 -4486
rect 10188 -4603 10222 -4579
rect 11476 -4452 11510 -4428
rect 11476 -4545 11510 -4486
rect 11476 -4603 11510 -4579
rect 13592 -4452 13626 -4428
rect 13592 -4545 13626 -4486
rect 13592 -4603 13626 -4579
rect 15524 -4452 15558 -4428
rect 15524 -4545 15558 -4486
rect 15524 -4603 15558 -4579
rect -2232 -5237 -2198 -5213
rect -2232 -5330 -2198 -5271
rect -2232 -5388 -2198 -5364
rect -116 -5237 -82 -5213
rect -116 -5330 -82 -5271
rect -116 -5388 -82 -5364
rect 344 -5237 378 -5213
rect 344 -5330 378 -5271
rect 344 -5388 378 -5364
rect 1172 -5237 1206 -5213
rect 1172 -5330 1206 -5271
rect 1172 -5388 1206 -5364
rect 1632 -5237 1666 -5213
rect 1632 -5330 1666 -5271
rect 1632 -5388 1666 -5364
rect 2460 -5237 2494 -5213
rect 2460 -5330 2494 -5271
rect 2460 -5388 2494 -5364
rect 2920 -5237 2954 -5213
rect 2920 -5330 2954 -5271
rect 2920 -5388 2954 -5364
rect 3748 -5237 3782 -5213
rect 3748 -5330 3782 -5271
rect 3748 -5388 3782 -5364
rect 4208 -5237 4242 -5213
rect 4208 -5330 4242 -5271
rect 4208 -5388 4242 -5364
rect 5036 -5237 5070 -5213
rect 5036 -5330 5070 -5271
rect 5036 -5388 5070 -5364
rect 5496 -5237 5530 -5213
rect 5496 -5330 5530 -5271
rect 5496 -5388 5530 -5364
rect 6324 -5237 6358 -5213
rect 6324 -5330 6358 -5271
rect 6324 -5388 6358 -5364
rect 6784 -5237 6818 -5213
rect 6784 -5330 6818 -5271
rect 6784 -5388 6818 -5364
rect 7612 -5237 7646 -5213
rect 7612 -5330 7646 -5271
rect 7612 -5388 7646 -5364
rect 8072 -5237 8106 -5213
rect 8072 -5330 8106 -5271
rect 8072 -5388 8106 -5364
rect 8900 -5237 8934 -5213
rect 8900 -5330 8934 -5271
rect 8900 -5388 8934 -5364
rect 9360 -5237 9394 -5213
rect 9360 -5330 9394 -5271
rect 9360 -5388 9394 -5364
rect 10188 -5237 10222 -5213
rect 10188 -5330 10222 -5271
rect 10188 -5388 10222 -5364
rect 11476 -5237 11510 -5213
rect 11476 -5330 11510 -5271
rect 11476 -5388 11510 -5364
rect 12396 -5237 12430 -5213
rect 12396 -5330 12430 -5271
rect 12396 -5388 12430 -5364
rect 13132 -5237 13166 -5213
rect 13132 -5330 13166 -5271
rect 13132 -5388 13166 -5364
rect 13592 -5237 13626 -5213
rect 13592 -5330 13626 -5271
rect 13592 -5388 13626 -5364
rect 15524 -5237 15558 -5213
rect 15524 -5330 15558 -5271
rect 15524 -5388 15558 -5364
rect -2232 -5540 -2198 -5516
rect -2232 -5633 -2198 -5574
rect -2232 -5691 -2198 -5667
rect -116 -5540 -82 -5516
rect -116 -5633 -82 -5574
rect -116 -5691 -82 -5667
rect 344 -5540 378 -5516
rect 344 -5633 378 -5574
rect 344 -5691 378 -5667
rect 1172 -5540 1206 -5516
rect 1172 -5633 1206 -5574
rect 1172 -5691 1206 -5667
rect 1632 -5540 1666 -5516
rect 1632 -5633 1666 -5574
rect 1632 -5691 1666 -5667
rect 2460 -5540 2494 -5516
rect 2460 -5633 2494 -5574
rect 2460 -5691 2494 -5667
rect 2920 -5540 2954 -5516
rect 2920 -5633 2954 -5574
rect 2920 -5691 2954 -5667
rect 3748 -5540 3782 -5516
rect 3748 -5633 3782 -5574
rect 3748 -5691 3782 -5667
rect 4208 -5540 4242 -5516
rect 4208 -5633 4242 -5574
rect 4208 -5691 4242 -5667
rect 5036 -5540 5070 -5516
rect 5036 -5633 5070 -5574
rect 5036 -5691 5070 -5667
rect 5496 -5540 5530 -5516
rect 5496 -5633 5530 -5574
rect 5496 -5691 5530 -5667
rect 6324 -5540 6358 -5516
rect 6324 -5633 6358 -5574
rect 6324 -5691 6358 -5667
rect 6784 -5540 6818 -5516
rect 6784 -5633 6818 -5574
rect 6784 -5691 6818 -5667
rect 7612 -5540 7646 -5516
rect 7612 -5633 7646 -5574
rect 7612 -5691 7646 -5667
rect 8072 -5540 8106 -5516
rect 8072 -5633 8106 -5574
rect 8072 -5691 8106 -5667
rect 8900 -5540 8934 -5516
rect 8900 -5633 8934 -5574
rect 8900 -5691 8934 -5667
rect 9360 -5540 9394 -5516
rect 9360 -5633 9394 -5574
rect 9360 -5691 9394 -5667
rect 10188 -5540 10222 -5516
rect 10188 -5633 10222 -5574
rect 10188 -5691 10222 -5667
rect 11476 -5540 11510 -5516
rect 11476 -5633 11510 -5574
rect 11476 -5691 11510 -5667
rect 13592 -5540 13626 -5516
rect 13592 -5633 13626 -5574
rect 13592 -5691 13626 -5667
rect 15524 -5540 15558 -5516
rect 15524 -5633 15558 -5574
rect 15524 -5691 15558 -5667
rect -2232 -6325 -2198 -6301
rect -2232 -6418 -2198 -6359
rect -2232 -6476 -2198 -6452
rect -1036 -6325 -1002 -6301
rect -1036 -6418 -1002 -6359
rect -1036 -6476 -1002 -6452
rect -668 -6325 -634 -6301
rect -668 -6418 -634 -6359
rect -668 -6476 -634 -6452
rect -208 -6325 -174 -6301
rect -208 -6418 -174 -6359
rect -208 -6476 -174 -6452
rect 528 -6325 562 -6301
rect 528 -6418 562 -6359
rect 528 -6476 562 -6452
rect 988 -6325 1022 -6301
rect 1356 -6325 1390 -6301
rect 988 -6418 1022 -6359
rect 988 -6476 1022 -6452
rect 1356 -6418 1390 -6359
rect 1356 -6476 1390 -6452
rect 1816 -6325 1850 -6301
rect 1816 -6418 1850 -6359
rect 1816 -6476 1850 -6452
rect 2276 -6325 2310 -6301
rect 2276 -6418 2310 -6359
rect 2276 -6476 2310 -6452
rect 3104 -6325 3138 -6301
rect 3104 -6418 3138 -6359
rect 3104 -6476 3138 -6452
rect 3564 -6325 3598 -6301
rect 3564 -6418 3598 -6359
rect 3564 -6476 3598 -6452
rect 6324 -6325 6358 -6301
rect 6324 -6418 6358 -6359
rect 6324 -6476 6358 -6452
rect 6784 -6325 6818 -6301
rect 6784 -6418 6818 -6359
rect 6784 -6476 6818 -6452
rect 7612 -6325 7646 -6301
rect 7612 -6418 7646 -6359
rect 7612 -6476 7646 -6452
rect 8072 -6325 8106 -6301
rect 8072 -6418 8106 -6359
rect 8072 -6476 8106 -6452
rect 8900 -6325 8934 -6301
rect 8900 -6418 8934 -6359
rect 8900 -6476 8934 -6452
rect 9360 -6325 9394 -6301
rect 9360 -6418 9394 -6359
rect 9360 -6476 9394 -6452
rect 10188 -6325 10222 -6301
rect 10188 -6418 10222 -6359
rect 10188 -6476 10222 -6452
rect 10648 -6325 10682 -6301
rect 10648 -6418 10682 -6359
rect 10648 -6476 10682 -6452
rect 11568 -6325 11602 -6301
rect 11568 -6418 11602 -6359
rect 11568 -6476 11602 -6452
rect 13500 -6325 13534 -6301
rect 13500 -6418 13534 -6359
rect 13500 -6476 13534 -6452
rect 14696 -6325 14730 -6301
rect 14696 -6418 14730 -6359
rect 14696 -6476 14730 -6452
rect 15892 -6325 15926 -6301
rect 15892 -6418 15926 -6359
rect 15892 -6476 15926 -6452
rect -2692 -6628 -2658 -6604
rect -2692 -6721 -2658 -6662
rect -2692 -6779 -2658 -6755
rect -116 -6628 -82 -6604
rect -116 -6721 -82 -6662
rect -116 -6779 -82 -6755
rect 1448 -6628 1482 -6604
rect 1448 -6721 1482 -6662
rect 1448 -6779 1482 -6755
rect 3012 -6628 3046 -6604
rect 3012 -6721 3046 -6662
rect 3012 -6779 3046 -6755
rect 4576 -6628 4610 -6604
rect 4576 -6721 4610 -6662
rect 4576 -6779 4610 -6755
rect 6140 -6628 6174 -6604
rect 6140 -6721 6174 -6662
rect 6140 -6779 6174 -6755
rect 7704 -6628 7738 -6604
rect 7704 -6721 7738 -6662
rect 7704 -6779 7738 -6755
rect 9268 -6628 9302 -6604
rect 9268 -6721 9302 -6662
rect 9268 -6779 9302 -6755
rect 15892 -6628 15926 -6604
rect 15892 -6721 15926 -6662
rect 15892 -6779 15926 -6755
rect -2232 -7413 -2198 -7389
rect -2232 -7506 -2198 -7447
rect -2232 -7564 -2198 -7540
rect -116 -7413 -82 -7389
rect -116 -7506 -82 -7447
rect -116 -7564 -82 -7540
rect 1448 -7413 1482 -7389
rect 1448 -7506 1482 -7447
rect 1448 -7564 1482 -7540
rect 2828 -7413 2862 -7389
rect 3196 -7413 3230 -7389
rect 2828 -7506 2862 -7447
rect 2828 -7564 2862 -7540
rect 3196 -7506 3230 -7447
rect 3196 -7564 3230 -7540
rect 3656 -7413 3690 -7389
rect 3656 -7506 3690 -7447
rect 3656 -7564 3690 -7540
rect 4024 -7413 4058 -7389
rect 4024 -7506 4058 -7447
rect 4024 -7564 4058 -7540
rect 4484 -7413 4518 -7389
rect 4484 -7506 4518 -7447
rect 4484 -7564 4518 -7540
rect 5404 -7413 5438 -7389
rect 5404 -7506 5438 -7447
rect 5404 -7564 5438 -7540
rect 5864 -7413 5898 -7389
rect 5864 -7506 5898 -7447
rect 5864 -7564 5898 -7540
rect 7704 -7413 7738 -7389
rect 7704 -7506 7738 -7447
rect 7704 -7564 7738 -7540
rect 9268 -7413 9302 -7389
rect 9268 -7506 9302 -7447
rect 9268 -7564 9302 -7540
rect 15892 -7413 15926 -7389
rect 15892 -7506 15926 -7447
rect 15892 -7564 15926 -7540
rect -2232 -7716 -2198 -7692
rect -2232 -7809 -2198 -7750
rect -2232 -7867 -2198 -7843
rect -1036 -7716 -1002 -7692
rect -1036 -7809 -1002 -7750
rect -1036 -7867 -1002 -7843
rect -668 -7716 -634 -7692
rect -668 -7809 -634 -7750
rect -668 -7867 -634 -7843
rect -208 -7716 -174 -7692
rect -208 -7809 -174 -7750
rect -208 -7867 -174 -7843
rect 528 -7716 562 -7692
rect 528 -7809 562 -7750
rect 528 -7867 562 -7843
rect 988 -7716 1022 -7692
rect 988 -7809 1022 -7750
rect 1356 -7716 1390 -7692
rect 1356 -7809 1390 -7750
rect 988 -7867 1022 -7843
rect 1356 -7867 1390 -7843
rect 1816 -7716 1850 -7692
rect 1816 -7809 1850 -7750
rect 1816 -7867 1850 -7843
rect 2276 -7716 2310 -7692
rect 2276 -7809 2310 -7750
rect 2276 -7867 2310 -7843
rect 3104 -7716 3138 -7692
rect 3104 -7809 3138 -7750
rect 3104 -7867 3138 -7843
rect 3564 -7716 3598 -7692
rect 3564 -7809 3598 -7750
rect 3564 -7867 3598 -7843
rect 6324 -7716 6358 -7692
rect 6324 -7809 6358 -7750
rect 6324 -7867 6358 -7843
rect 6784 -7716 6818 -7692
rect 6784 -7809 6818 -7750
rect 6784 -7867 6818 -7843
rect 7612 -7716 7646 -7692
rect 7612 -7809 7646 -7750
rect 7612 -7867 7646 -7843
rect 8072 -7716 8106 -7692
rect 8072 -7809 8106 -7750
rect 8072 -7867 8106 -7843
rect 8900 -7716 8934 -7692
rect 8900 -7809 8934 -7750
rect 8900 -7867 8934 -7843
rect 9360 -7716 9394 -7692
rect 9360 -7809 9394 -7750
rect 9360 -7867 9394 -7843
rect 10188 -7716 10222 -7692
rect 10188 -7809 10222 -7750
rect 10188 -7867 10222 -7843
rect 10648 -7716 10682 -7692
rect 10648 -7809 10682 -7750
rect 10648 -7867 10682 -7843
rect 11568 -7716 11602 -7692
rect 11568 -7809 11602 -7750
rect 11568 -7867 11602 -7843
rect 13500 -7716 13534 -7692
rect 13500 -7809 13534 -7750
rect 13500 -7867 13534 -7843
rect 14696 -7716 14730 -7692
rect 14696 -7809 14730 -7750
rect 14696 -7867 14730 -7843
rect 15892 -7716 15926 -7692
rect 15892 -7809 15926 -7750
rect 15892 -7867 15926 -7843
rect -2232 -8501 -2198 -8477
rect -2232 -8594 -2198 -8535
rect -2232 -8652 -2198 -8628
rect -116 -8501 -82 -8477
rect -116 -8594 -82 -8535
rect -116 -8652 -82 -8628
rect 344 -8501 378 -8477
rect 344 -8594 378 -8535
rect 344 -8652 378 -8628
rect 1172 -8501 1206 -8477
rect 1172 -8594 1206 -8535
rect 1172 -8652 1206 -8628
rect 1632 -8501 1666 -8477
rect 1632 -8594 1666 -8535
rect 1632 -8652 1666 -8628
rect 2460 -8501 2494 -8477
rect 2460 -8594 2494 -8535
rect 2460 -8652 2494 -8628
rect 2920 -8501 2954 -8477
rect 2920 -8594 2954 -8535
rect 2920 -8652 2954 -8628
rect 3748 -8501 3782 -8477
rect 3748 -8594 3782 -8535
rect 3748 -8652 3782 -8628
rect 4208 -8501 4242 -8477
rect 4208 -8594 4242 -8535
rect 4208 -8652 4242 -8628
rect 5036 -8501 5070 -8477
rect 5036 -8594 5070 -8535
rect 5036 -8652 5070 -8628
rect 5496 -8501 5530 -8477
rect 5496 -8594 5530 -8535
rect 5496 -8652 5530 -8628
rect 6324 -8501 6358 -8477
rect 6324 -8594 6358 -8535
rect 6324 -8652 6358 -8628
rect 6784 -8501 6818 -8477
rect 6784 -8594 6818 -8535
rect 6784 -8652 6818 -8628
rect 7612 -8501 7646 -8477
rect 7612 -8594 7646 -8535
rect 7612 -8652 7646 -8628
rect 8072 -8501 8106 -8477
rect 8072 -8594 8106 -8535
rect 8072 -8652 8106 -8628
rect 8900 -8501 8934 -8477
rect 8900 -8594 8934 -8535
rect 8900 -8652 8934 -8628
rect 9360 -8501 9394 -8477
rect 9360 -8594 9394 -8535
rect 9360 -8652 9394 -8628
rect 10188 -8501 10222 -8477
rect 10188 -8594 10222 -8535
rect 10188 -8652 10222 -8628
rect 11476 -8501 11510 -8477
rect 11476 -8594 11510 -8535
rect 11476 -8652 11510 -8628
rect 13592 -8501 13626 -8477
rect 13592 -8594 13626 -8535
rect 13592 -8652 13626 -8628
rect 15524 -8501 15558 -8477
rect 15524 -8594 15558 -8535
rect 15524 -8652 15558 -8628
rect -2232 -8804 -2198 -8780
rect -2232 -8897 -2198 -8838
rect -2232 -8955 -2198 -8931
rect -116 -8804 -82 -8780
rect -116 -8897 -82 -8838
rect -116 -8955 -82 -8931
rect 344 -8804 378 -8780
rect 344 -8897 378 -8838
rect 344 -8955 378 -8931
rect 1172 -8804 1206 -8780
rect 1172 -8897 1206 -8838
rect 1172 -8955 1206 -8931
rect 1632 -8804 1666 -8780
rect 1632 -8897 1666 -8838
rect 1632 -8955 1666 -8931
rect 2460 -8804 2494 -8780
rect 2460 -8897 2494 -8838
rect 2460 -8955 2494 -8931
rect 2920 -8804 2954 -8780
rect 2920 -8897 2954 -8838
rect 2920 -8955 2954 -8931
rect 3748 -8804 3782 -8780
rect 3748 -8897 3782 -8838
rect 3748 -8955 3782 -8931
rect 4208 -8804 4242 -8780
rect 4208 -8897 4242 -8838
rect 4208 -8955 4242 -8931
rect 5036 -8804 5070 -8780
rect 5036 -8897 5070 -8838
rect 5036 -8955 5070 -8931
rect 5496 -8804 5530 -8780
rect 5496 -8897 5530 -8838
rect 5496 -8955 5530 -8931
rect 6324 -8804 6358 -8780
rect 6324 -8897 6358 -8838
rect 6324 -8955 6358 -8931
rect 6784 -8804 6818 -8780
rect 6784 -8897 6818 -8838
rect 6784 -8955 6818 -8931
rect 7612 -8804 7646 -8780
rect 7612 -8897 7646 -8838
rect 7612 -8955 7646 -8931
rect 8072 -8804 8106 -8780
rect 8072 -8897 8106 -8838
rect 8072 -8955 8106 -8931
rect 8900 -8804 8934 -8780
rect 8900 -8897 8934 -8838
rect 8900 -8955 8934 -8931
rect 9360 -8804 9394 -8780
rect 9360 -8897 9394 -8838
rect 9360 -8955 9394 -8931
rect 10188 -8804 10222 -8780
rect 10188 -8897 10222 -8838
rect 10188 -8955 10222 -8931
rect 11476 -8804 11510 -8780
rect 11476 -8897 11510 -8838
rect 11476 -8955 11510 -8931
rect 12396 -8804 12430 -8780
rect 12396 -8897 12430 -8838
rect 12396 -8955 12430 -8931
rect 13132 -8804 13166 -8780
rect 13132 -8897 13166 -8838
rect 13132 -8955 13166 -8931
rect 13592 -8804 13626 -8780
rect 13592 -8897 13626 -8838
rect 13592 -8955 13626 -8931
rect 15524 -8804 15558 -8780
rect 15524 -8897 15558 -8838
rect 15524 -8955 15558 -8931
rect -2232 -9589 -2198 -9565
rect -2232 -9682 -2198 -9623
rect -2232 -9740 -2198 -9716
rect -116 -9589 -82 -9565
rect -116 -9682 -82 -9623
rect -116 -9740 -82 -9716
rect 344 -9589 378 -9565
rect 344 -9682 378 -9623
rect 344 -9740 378 -9716
rect 1172 -9589 1206 -9565
rect 1172 -9682 1206 -9623
rect 1172 -9740 1206 -9716
rect 1632 -9589 1666 -9565
rect 1632 -9682 1666 -9623
rect 1632 -9740 1666 -9716
rect 2460 -9589 2494 -9565
rect 2460 -9682 2494 -9623
rect 2460 -9740 2494 -9716
rect 2920 -9589 2954 -9565
rect 2920 -9682 2954 -9623
rect 2920 -9740 2954 -9716
rect 3748 -9589 3782 -9565
rect 3748 -9682 3782 -9623
rect 3748 -9740 3782 -9716
rect 4208 -9589 4242 -9565
rect 4208 -9682 4242 -9623
rect 4208 -9740 4242 -9716
rect 5036 -9589 5070 -9565
rect 5036 -9682 5070 -9623
rect 5036 -9740 5070 -9716
rect 5496 -9589 5530 -9565
rect 5496 -9682 5530 -9623
rect 5496 -9740 5530 -9716
rect 6324 -9589 6358 -9565
rect 6324 -9682 6358 -9623
rect 6324 -9740 6358 -9716
rect 6784 -9589 6818 -9565
rect 6784 -9682 6818 -9623
rect 6784 -9740 6818 -9716
rect 7612 -9589 7646 -9565
rect 7612 -9682 7646 -9623
rect 7612 -9740 7646 -9716
rect 8072 -9589 8106 -9565
rect 8072 -9682 8106 -9623
rect 8072 -9740 8106 -9716
rect 8900 -9589 8934 -9565
rect 8900 -9682 8934 -9623
rect 8900 -9740 8934 -9716
rect 9360 -9589 9394 -9565
rect 9360 -9682 9394 -9623
rect 9360 -9740 9394 -9716
rect 10188 -9589 10222 -9565
rect 10188 -9682 10222 -9623
rect 10188 -9740 10222 -9716
rect 11476 -9589 11510 -9565
rect 11476 -9682 11510 -9623
rect 11476 -9740 11510 -9716
rect 13592 -9589 13626 -9565
rect 13592 -9682 13626 -9623
rect 13592 -9740 13626 -9716
rect 15524 -9589 15558 -9565
rect 15524 -9682 15558 -9623
rect 15524 -9740 15558 -9716
rect -2232 -9892 -2198 -9868
rect -2232 -9985 -2198 -9926
rect -2232 -10043 -2198 -10019
rect -116 -9892 -82 -9868
rect -116 -9985 -82 -9926
rect -116 -10043 -82 -10019
rect 344 -9892 378 -9868
rect 344 -9985 378 -9926
rect 344 -10043 378 -10019
rect 1172 -9892 1206 -9868
rect 1172 -9985 1206 -9926
rect 1172 -10043 1206 -10019
rect 1632 -9892 1666 -9868
rect 1632 -9985 1666 -9926
rect 1632 -10043 1666 -10019
rect 2460 -9892 2494 -9868
rect 2460 -9985 2494 -9926
rect 2460 -10043 2494 -10019
rect 2920 -9892 2954 -9868
rect 2920 -9985 2954 -9926
rect 2920 -10043 2954 -10019
rect 3748 -9892 3782 -9868
rect 3748 -9985 3782 -9926
rect 3748 -10043 3782 -10019
rect 4208 -9892 4242 -9868
rect 4208 -9985 4242 -9926
rect 4208 -10043 4242 -10019
rect 5036 -9892 5070 -9868
rect 5036 -9985 5070 -9926
rect 5036 -10043 5070 -10019
rect 5496 -9892 5530 -9868
rect 5496 -9985 5530 -9926
rect 5496 -10043 5530 -10019
rect 6324 -9892 6358 -9868
rect 6324 -9985 6358 -9926
rect 6324 -10043 6358 -10019
rect 6784 -9892 6818 -9868
rect 6784 -9985 6818 -9926
rect 6784 -10043 6818 -10019
rect 7612 -9892 7646 -9868
rect 7612 -9985 7646 -9926
rect 7612 -10043 7646 -10019
rect 8072 -9892 8106 -9868
rect 8072 -9985 8106 -9926
rect 8072 -10043 8106 -10019
rect 8900 -9892 8934 -9868
rect 8900 -9985 8934 -9926
rect 8900 -10043 8934 -10019
rect 9360 -9892 9394 -9868
rect 9360 -9985 9394 -9926
rect 9360 -10043 9394 -10019
rect 10188 -9892 10222 -9868
rect 10188 -9985 10222 -9926
rect 10188 -10043 10222 -10019
rect 11476 -9892 11510 -9868
rect 11476 -9985 11510 -9926
rect 11476 -10043 11510 -10019
rect 12396 -9892 12430 -9868
rect 12396 -9985 12430 -9926
rect 12396 -10043 12430 -10019
rect 13132 -9892 13166 -9868
rect 13132 -9985 13166 -9926
rect 13132 -10043 13166 -10019
rect 13592 -9892 13626 -9868
rect 13592 -9985 13626 -9926
rect 13592 -10043 13626 -10019
rect 15524 -9892 15558 -9868
rect 15524 -9985 15558 -9926
rect 15524 -10043 15558 -10019
rect -2232 -10677 -2198 -10653
rect -1680 -10677 -1646 -10653
rect -2232 -10770 -2198 -10711
rect -2232 -10828 -2198 -10804
rect -1680 -10770 -1646 -10711
rect -1680 -10828 -1646 -10804
rect -116 -10677 -82 -10653
rect -116 -10770 -82 -10711
rect -116 -10828 -82 -10804
rect 344 -10677 378 -10653
rect 344 -10770 378 -10711
rect 344 -10828 378 -10804
rect 1172 -10677 1206 -10653
rect 1172 -10770 1206 -10711
rect 1172 -10828 1206 -10804
rect 1632 -10677 1666 -10653
rect 1632 -10770 1666 -10711
rect 1632 -10828 1666 -10804
rect 2460 -10677 2494 -10653
rect 2460 -10770 2494 -10711
rect 2460 -10828 2494 -10804
rect 2920 -10677 2954 -10653
rect 2920 -10770 2954 -10711
rect 2920 -10828 2954 -10804
rect 3748 -10677 3782 -10653
rect 3748 -10770 3782 -10711
rect 3748 -10828 3782 -10804
rect 4208 -10677 4242 -10653
rect 4208 -10770 4242 -10711
rect 4208 -10828 4242 -10804
rect 5036 -10677 5070 -10653
rect 5036 -10770 5070 -10711
rect 5036 -10828 5070 -10804
rect 5496 -10677 5530 -10653
rect 5496 -10770 5530 -10711
rect 5496 -10828 5530 -10804
rect 6324 -10677 6358 -10653
rect 6324 -10770 6358 -10711
rect 6324 -10828 6358 -10804
rect 6784 -10677 6818 -10653
rect 6784 -10770 6818 -10711
rect 6784 -10828 6818 -10804
rect 7612 -10677 7646 -10653
rect 7612 -10770 7646 -10711
rect 7612 -10828 7646 -10804
rect 8072 -10677 8106 -10653
rect 8072 -10770 8106 -10711
rect 8072 -10828 8106 -10804
rect 8900 -10677 8934 -10653
rect 8900 -10770 8934 -10711
rect 8900 -10828 8934 -10804
rect 9360 -10677 9394 -10653
rect 9360 -10770 9394 -10711
rect 9360 -10828 9394 -10804
rect 10188 -10677 10222 -10653
rect 10188 -10770 10222 -10711
rect 10188 -10828 10222 -10804
rect 11476 -10677 11510 -10653
rect 11476 -10770 11510 -10711
rect 11476 -10828 11510 -10804
rect 13500 -10677 13534 -10653
rect 13500 -10770 13534 -10711
rect 13500 -10828 13534 -10804
rect 14696 -10677 14730 -10653
rect 14696 -10770 14730 -10711
rect 14696 -10828 14730 -10804
rect 15892 -10677 15926 -10653
rect 15892 -10770 15926 -10711
rect 15892 -10828 15926 -10804
rect -2232 -10980 -2198 -10956
rect -2232 -11073 -2198 -11014
rect -2232 -11131 -2198 -11107
rect -116 -10980 -82 -10956
rect -116 -11073 -82 -11014
rect -116 -11131 -82 -11107
rect 344 -10980 378 -10956
rect 344 -11073 378 -11014
rect 344 -11131 378 -11107
rect 1172 -10980 1206 -10956
rect 1172 -11073 1206 -11014
rect 1172 -11131 1206 -11107
rect 1632 -10980 1666 -10956
rect 1632 -11073 1666 -11014
rect 1632 -11131 1666 -11107
rect 2460 -10980 2494 -10956
rect 2460 -11073 2494 -11014
rect 2460 -11131 2494 -11107
rect 2920 -10980 2954 -10956
rect 2920 -11073 2954 -11014
rect 2920 -11131 2954 -11107
rect 3748 -10980 3782 -10956
rect 3748 -11073 3782 -11014
rect 3748 -11131 3782 -11107
rect 4208 -10980 4242 -10956
rect 4208 -11073 4242 -11014
rect 4208 -11131 4242 -11107
rect 5036 -10980 5070 -10956
rect 5036 -11073 5070 -11014
rect 5036 -11131 5070 -11107
rect 5496 -10980 5530 -10956
rect 5496 -11073 5530 -11014
rect 5496 -11131 5530 -11107
rect 6324 -10980 6358 -10956
rect 6324 -11073 6358 -11014
rect 6324 -11131 6358 -11107
rect 6784 -10980 6818 -10956
rect 6784 -11073 6818 -11014
rect 6784 -11131 6818 -11107
rect 7612 -10980 7646 -10956
rect 7612 -11073 7646 -11014
rect 7612 -11131 7646 -11107
rect 8072 -10980 8106 -10956
rect 8072 -11073 8106 -11014
rect 8072 -11131 8106 -11107
rect 8900 -10980 8934 -10956
rect 8900 -11073 8934 -11014
rect 8900 -11131 8934 -11107
rect 9360 -10980 9394 -10956
rect 9360 -11073 9394 -11014
rect 9360 -11131 9394 -11107
rect 10188 -10980 10222 -10956
rect 10188 -11073 10222 -11014
rect 10188 -11131 10222 -11107
rect 11476 -10980 11510 -10956
rect 11476 -11073 11510 -11014
rect 11476 -11131 11510 -11107
rect 13500 -10980 13534 -10956
rect 13500 -11073 13534 -11014
rect 13500 -11131 13534 -11107
rect 14696 -10980 14730 -10956
rect 14696 -11073 14730 -11014
rect 14696 -11131 14730 -11107
rect 15892 -10980 15926 -10956
rect 15892 -11073 15926 -11014
rect 15892 -11131 15926 -11107
rect -2232 -11765 -2198 -11741
rect -2232 -11858 -2198 -11799
rect -2232 -11916 -2198 -11892
rect -116 -11765 -82 -11741
rect -116 -11858 -82 -11799
rect -116 -11916 -82 -11892
rect 344 -11765 378 -11741
rect 344 -11858 378 -11799
rect 344 -11916 378 -11892
rect 1172 -11765 1206 -11741
rect 1172 -11858 1206 -11799
rect 1172 -11916 1206 -11892
rect 1632 -11765 1666 -11741
rect 1632 -11858 1666 -11799
rect 1632 -11916 1666 -11892
rect 2460 -11765 2494 -11741
rect 2460 -11858 2494 -11799
rect 2460 -11916 2494 -11892
rect 2920 -11765 2954 -11741
rect 2920 -11858 2954 -11799
rect 2920 -11916 2954 -11892
rect 3748 -11765 3782 -11741
rect 3748 -11858 3782 -11799
rect 3748 -11916 3782 -11892
rect 4208 -11765 4242 -11741
rect 4208 -11858 4242 -11799
rect 4208 -11916 4242 -11892
rect 5036 -11765 5070 -11741
rect 5036 -11858 5070 -11799
rect 5036 -11916 5070 -11892
rect 5496 -11765 5530 -11741
rect 5496 -11858 5530 -11799
rect 5496 -11916 5530 -11892
rect 6324 -11765 6358 -11741
rect 6324 -11858 6358 -11799
rect 6324 -11916 6358 -11892
rect 6784 -11765 6818 -11741
rect 6784 -11858 6818 -11799
rect 6784 -11916 6818 -11892
rect 7612 -11765 7646 -11741
rect 7612 -11858 7646 -11799
rect 7612 -11916 7646 -11892
rect 8072 -11765 8106 -11741
rect 8072 -11858 8106 -11799
rect 8072 -11916 8106 -11892
rect 8900 -11765 8934 -11741
rect 8900 -11858 8934 -11799
rect 8900 -11916 8934 -11892
rect 9360 -11765 9394 -11741
rect 9360 -11858 9394 -11799
rect 9360 -11916 9394 -11892
rect 10188 -11765 10222 -11741
rect 10188 -11858 10222 -11799
rect 10188 -11916 10222 -11892
rect 11476 -11765 11510 -11741
rect 11476 -11858 11510 -11799
rect 11476 -11916 11510 -11892
rect 12396 -11765 12430 -11741
rect 12396 -11858 12430 -11799
rect 12396 -11916 12430 -11892
rect 13132 -11765 13166 -11741
rect 13132 -11858 13166 -11799
rect 13132 -11916 13166 -11892
rect 13592 -11765 13626 -11741
rect 13592 -11858 13626 -11799
rect 13592 -11916 13626 -11892
rect 15524 -11765 15558 -11741
rect 15524 -11858 15558 -11799
rect 15524 -11916 15558 -11892
rect -2232 -12068 -2198 -12044
rect -2232 -12161 -2198 -12102
rect -2232 -12219 -2198 -12195
rect -116 -12068 -82 -12044
rect -116 -12161 -82 -12102
rect -116 -12219 -82 -12195
rect 344 -12068 378 -12044
rect 344 -12161 378 -12102
rect 344 -12219 378 -12195
rect 1172 -12068 1206 -12044
rect 1172 -12161 1206 -12102
rect 1172 -12219 1206 -12195
rect 1632 -12068 1666 -12044
rect 1632 -12161 1666 -12102
rect 1632 -12219 1666 -12195
rect 2460 -12068 2494 -12044
rect 2460 -12161 2494 -12102
rect 2460 -12219 2494 -12195
rect 2920 -12068 2954 -12044
rect 2920 -12161 2954 -12102
rect 2920 -12219 2954 -12195
rect 3748 -12068 3782 -12044
rect 3748 -12161 3782 -12102
rect 3748 -12219 3782 -12195
rect 4208 -12068 4242 -12044
rect 4208 -12161 4242 -12102
rect 4208 -12219 4242 -12195
rect 5036 -12068 5070 -12044
rect 5036 -12161 5070 -12102
rect 5036 -12219 5070 -12195
rect 5496 -12068 5530 -12044
rect 5496 -12161 5530 -12102
rect 5496 -12219 5530 -12195
rect 6324 -12068 6358 -12044
rect 6324 -12161 6358 -12102
rect 6324 -12219 6358 -12195
rect 6784 -12068 6818 -12044
rect 6784 -12161 6818 -12102
rect 6784 -12219 6818 -12195
rect 7612 -12068 7646 -12044
rect 7612 -12161 7646 -12102
rect 7612 -12219 7646 -12195
rect 8072 -12068 8106 -12044
rect 8072 -12161 8106 -12102
rect 8072 -12219 8106 -12195
rect 8900 -12068 8934 -12044
rect 8900 -12161 8934 -12102
rect 8900 -12219 8934 -12195
rect 9360 -12068 9394 -12044
rect 9360 -12161 9394 -12102
rect 9360 -12219 9394 -12195
rect 10188 -12068 10222 -12044
rect 10188 -12161 10222 -12102
rect 10188 -12219 10222 -12195
rect 11476 -12068 11510 -12044
rect 11476 -12161 11510 -12102
rect 11476 -12219 11510 -12195
rect 13592 -12068 13626 -12044
rect 13592 -12161 13626 -12102
rect 13592 -12219 13626 -12195
rect 15524 -12068 15558 -12044
rect 15524 -12161 15558 -12102
rect 15524 -12219 15558 -12195
rect -2232 -12853 -2198 -12829
rect -2232 -12946 -2198 -12887
rect -2232 -13004 -2198 -12980
rect -116 -12853 -82 -12829
rect -116 -12946 -82 -12887
rect -116 -13004 -82 -12980
rect 344 -12853 378 -12829
rect 344 -12946 378 -12887
rect 344 -13004 378 -12980
rect 1172 -12853 1206 -12829
rect 1172 -12946 1206 -12887
rect 1172 -13004 1206 -12980
rect 1632 -12853 1666 -12829
rect 1632 -12946 1666 -12887
rect 1632 -13004 1666 -12980
rect 2460 -12853 2494 -12829
rect 2460 -12946 2494 -12887
rect 2460 -13004 2494 -12980
rect 2920 -12853 2954 -12829
rect 2920 -12946 2954 -12887
rect 2920 -13004 2954 -12980
rect 3748 -12853 3782 -12829
rect 3748 -12946 3782 -12887
rect 3748 -13004 3782 -12980
rect 4208 -12853 4242 -12829
rect 4208 -12946 4242 -12887
rect 4208 -13004 4242 -12980
rect 5036 -12853 5070 -12829
rect 5036 -12946 5070 -12887
rect 5036 -13004 5070 -12980
rect 5496 -12853 5530 -12829
rect 5496 -12946 5530 -12887
rect 5496 -13004 5530 -12980
rect 6324 -12853 6358 -12829
rect 6324 -12946 6358 -12887
rect 6324 -13004 6358 -12980
rect 6784 -12853 6818 -12829
rect 6784 -12946 6818 -12887
rect 6784 -13004 6818 -12980
rect 7612 -12853 7646 -12829
rect 7612 -12946 7646 -12887
rect 7612 -13004 7646 -12980
rect 8072 -12853 8106 -12829
rect 8072 -12946 8106 -12887
rect 8072 -13004 8106 -12980
rect 8900 -12853 8934 -12829
rect 8900 -12946 8934 -12887
rect 8900 -13004 8934 -12980
rect 9360 -12853 9394 -12829
rect 9360 -12946 9394 -12887
rect 9360 -13004 9394 -12980
rect 10188 -12853 10222 -12829
rect 10188 -12946 10222 -12887
rect 10188 -13004 10222 -12980
rect 11476 -12853 11510 -12829
rect 11476 -12946 11510 -12887
rect 11476 -13004 11510 -12980
rect 12396 -12853 12430 -12829
rect 12396 -12946 12430 -12887
rect 12396 -13004 12430 -12980
rect 13132 -12853 13166 -12829
rect 13132 -12946 13166 -12887
rect 13132 -13004 13166 -12980
rect 13592 -12853 13626 -12829
rect 13592 -12946 13626 -12887
rect 13592 -13004 13626 -12980
rect 15524 -12853 15558 -12829
rect 15524 -12946 15558 -12887
rect 15524 -13004 15558 -12980
rect -2232 -13156 -2198 -13132
rect -2232 -13249 -2198 -13190
rect -2232 -13307 -2198 -13283
rect -116 -13156 -82 -13132
rect -116 -13249 -82 -13190
rect -116 -13307 -82 -13283
rect 344 -13156 378 -13132
rect 344 -13249 378 -13190
rect 344 -13307 378 -13283
rect 1172 -13156 1206 -13132
rect 1172 -13249 1206 -13190
rect 1172 -13307 1206 -13283
rect 1632 -13156 1666 -13132
rect 1632 -13249 1666 -13190
rect 1632 -13307 1666 -13283
rect 2460 -13156 2494 -13132
rect 2460 -13249 2494 -13190
rect 2460 -13307 2494 -13283
rect 2920 -13156 2954 -13132
rect 2920 -13249 2954 -13190
rect 2920 -13307 2954 -13283
rect 3748 -13156 3782 -13132
rect 3748 -13249 3782 -13190
rect 3748 -13307 3782 -13283
rect 4208 -13156 4242 -13132
rect 4208 -13249 4242 -13190
rect 4208 -13307 4242 -13283
rect 5036 -13156 5070 -13132
rect 5036 -13249 5070 -13190
rect 5036 -13307 5070 -13283
rect 5496 -13156 5530 -13132
rect 5496 -13249 5530 -13190
rect 5496 -13307 5530 -13283
rect 6324 -13156 6358 -13132
rect 6324 -13249 6358 -13190
rect 6324 -13307 6358 -13283
rect 6784 -13156 6818 -13132
rect 6784 -13249 6818 -13190
rect 6784 -13307 6818 -13283
rect 7612 -13156 7646 -13132
rect 7612 -13249 7646 -13190
rect 7612 -13307 7646 -13283
rect 8072 -13156 8106 -13132
rect 8072 -13249 8106 -13190
rect 8072 -13307 8106 -13283
rect 8900 -13156 8934 -13132
rect 8900 -13249 8934 -13190
rect 8900 -13307 8934 -13283
rect 9360 -13156 9394 -13132
rect 9360 -13249 9394 -13190
rect 9360 -13307 9394 -13283
rect 10188 -13156 10222 -13132
rect 10188 -13249 10222 -13190
rect 10188 -13307 10222 -13283
rect 11476 -13156 11510 -13132
rect 11476 -13249 11510 -13190
rect 11476 -13307 11510 -13283
rect 13592 -13156 13626 -13132
rect 13592 -13249 13626 -13190
rect 13592 -13307 13626 -13283
rect 15524 -13156 15558 -13132
rect 15524 -13249 15558 -13190
rect 15524 -13307 15558 -13283
rect -2232 -13941 -2198 -13917
rect -2232 -14034 -2198 -13975
rect -2232 -14092 -2198 -14068
rect -1036 -13941 -1002 -13917
rect -1036 -14034 -1002 -13975
rect -1036 -14092 -1002 -14068
rect -668 -13941 -634 -13917
rect -668 -14034 -634 -13975
rect -668 -14092 -634 -14068
rect -208 -13941 -174 -13917
rect -208 -14034 -174 -13975
rect -208 -14092 -174 -14068
rect 528 -13941 562 -13917
rect 528 -14034 562 -13975
rect 528 -14092 562 -14068
rect 988 -13941 1022 -13917
rect 1356 -13941 1390 -13917
rect 988 -14034 1022 -13975
rect 988 -14092 1022 -14068
rect 1356 -14034 1390 -13975
rect 1356 -14092 1390 -14068
rect 1816 -13941 1850 -13917
rect 1816 -14034 1850 -13975
rect 1816 -14092 1850 -14068
rect 2276 -13941 2310 -13917
rect 2276 -14034 2310 -13975
rect 2276 -14092 2310 -14068
rect 3104 -13941 3138 -13917
rect 3104 -14034 3138 -13975
rect 3104 -14092 3138 -14068
rect 3564 -13941 3598 -13917
rect 3564 -14034 3598 -13975
rect 3564 -14092 3598 -14068
rect 6324 -13941 6358 -13917
rect 6324 -14034 6358 -13975
rect 6324 -14092 6358 -14068
rect 6784 -13941 6818 -13917
rect 6784 -14034 6818 -13975
rect 6784 -14092 6818 -14068
rect 7612 -13941 7646 -13917
rect 7612 -14034 7646 -13975
rect 7612 -14092 7646 -14068
rect 8072 -13941 8106 -13917
rect 8072 -14034 8106 -13975
rect 8072 -14092 8106 -14068
rect 8900 -13941 8934 -13917
rect 8900 -14034 8934 -13975
rect 8900 -14092 8934 -14068
rect 9360 -13941 9394 -13917
rect 9360 -14034 9394 -13975
rect 9360 -14092 9394 -14068
rect 10188 -13941 10222 -13917
rect 10188 -14034 10222 -13975
rect 10188 -14092 10222 -14068
rect 10648 -13941 10682 -13917
rect 10648 -14034 10682 -13975
rect 10648 -14092 10682 -14068
rect 11568 -13941 11602 -13917
rect 11568 -14034 11602 -13975
rect 11568 -14092 11602 -14068
rect 13500 -13941 13534 -13917
rect 13500 -14034 13534 -13975
rect 13500 -14092 13534 -14068
rect 14696 -13941 14730 -13917
rect 14696 -14034 14730 -13975
rect 14696 -14092 14730 -14068
rect 15892 -13941 15926 -13917
rect 15892 -14034 15926 -13975
rect 15892 -14092 15926 -14068
<< psubdiffcont >>
rect -2232 -445 -2198 -411
rect -1036 -445 -1002 -411
rect -668 -445 -634 -411
rect -208 -445 -174 -411
rect 528 -445 562 -411
rect 988 -445 1022 -411
rect 1356 -445 1390 -411
rect 1816 -445 1850 -411
rect 2276 -445 2310 -411
rect 3104 -445 3138 -411
rect 3564 -445 3598 -411
rect 6324 -445 6358 -411
rect 6784 -445 6818 -411
rect 7612 -445 7646 -411
rect 8072 -445 8106 -411
rect 8900 -445 8934 -411
rect 9360 -445 9394 -411
rect 10188 -445 10222 -411
rect 10648 -445 10682 -411
rect 11568 -445 11602 -411
rect 13500 -445 13534 -411
rect 14696 -445 14730 -411
rect 15892 -445 15926 -411
rect -2232 -701 -2198 -667
rect -116 -701 -82 -667
rect 344 -701 378 -667
rect 1172 -701 1206 -667
rect 1632 -701 1666 -667
rect 2460 -701 2494 -667
rect 2920 -701 2954 -667
rect 3748 -701 3782 -667
rect 4208 -701 4242 -667
rect 5036 -701 5070 -667
rect 5496 -701 5530 -667
rect 6324 -701 6358 -667
rect 6784 -701 6818 -667
rect 7612 -701 7646 -667
rect 8072 -701 8106 -667
rect 8900 -701 8934 -667
rect 9360 -701 9394 -667
rect 10188 -701 10222 -667
rect 11476 -701 11510 -667
rect 13592 -701 13626 -667
rect 15524 -701 15558 -667
rect -2232 -1533 -2198 -1499
rect -116 -1533 -82 -1499
rect 344 -1533 378 -1499
rect 1172 -1533 1206 -1499
rect 1632 -1533 1666 -1499
rect 2460 -1533 2494 -1499
rect 2920 -1533 2954 -1499
rect 3748 -1533 3782 -1499
rect 4208 -1533 4242 -1499
rect 5036 -1533 5070 -1499
rect 5496 -1533 5530 -1499
rect 6324 -1533 6358 -1499
rect 6784 -1533 6818 -1499
rect 7612 -1533 7646 -1499
rect 8072 -1533 8106 -1499
rect 8900 -1533 8934 -1499
rect 9360 -1533 9394 -1499
rect 10188 -1533 10222 -1499
rect 11476 -1533 11510 -1499
rect 12396 -1533 12430 -1499
rect 13132 -1533 13166 -1499
rect 13592 -1533 13626 -1499
rect 15524 -1533 15558 -1499
rect -2232 -1789 -2198 -1755
rect -116 -1789 -82 -1755
rect 344 -1789 378 -1755
rect 1172 -1789 1206 -1755
rect 1632 -1789 1666 -1755
rect 2460 -1789 2494 -1755
rect 2920 -1789 2954 -1755
rect 3748 -1789 3782 -1755
rect 4208 -1789 4242 -1755
rect 5036 -1789 5070 -1755
rect 5496 -1789 5530 -1755
rect 6324 -1789 6358 -1755
rect 6784 -1789 6818 -1755
rect 7612 -1789 7646 -1755
rect 8072 -1789 8106 -1755
rect 8900 -1789 8934 -1755
rect 9360 -1789 9394 -1755
rect 10188 -1789 10222 -1755
rect 11476 -1789 11510 -1755
rect 13592 -1789 13626 -1755
rect 15524 -1789 15558 -1755
rect -2232 -2621 -2198 -2587
rect -116 -2621 -82 -2587
rect 344 -2621 378 -2587
rect 1172 -2621 1206 -2587
rect 1632 -2621 1666 -2587
rect 2460 -2621 2494 -2587
rect 2920 -2621 2954 -2587
rect 3748 -2621 3782 -2587
rect 4208 -2621 4242 -2587
rect 5036 -2621 5070 -2587
rect 5496 -2621 5530 -2587
rect 6324 -2621 6358 -2587
rect 6784 -2621 6818 -2587
rect 7612 -2621 7646 -2587
rect 8072 -2621 8106 -2587
rect 8900 -2621 8934 -2587
rect 9360 -2621 9394 -2587
rect 10188 -2621 10222 -2587
rect 11476 -2621 11510 -2587
rect 12396 -2621 12430 -2587
rect 13132 -2621 13166 -2587
rect 13592 -2621 13626 -2587
rect 15524 -2621 15558 -2587
rect -2232 -2877 -2198 -2843
rect -1680 -2877 -1646 -2843
rect -116 -2877 -82 -2843
rect 344 -2877 378 -2843
rect 1172 -2877 1206 -2843
rect 1632 -2877 1666 -2843
rect 2460 -2877 2494 -2843
rect 2920 -2877 2954 -2843
rect 3748 -2877 3782 -2843
rect 4208 -2877 4242 -2843
rect 5036 -2877 5070 -2843
rect 5496 -2877 5530 -2843
rect 6324 -2877 6358 -2843
rect 6784 -2877 6818 -2843
rect 7612 -2877 7646 -2843
rect 8072 -2877 8106 -2843
rect 8900 -2877 8934 -2843
rect 9360 -2877 9394 -2843
rect 10188 -2877 10222 -2843
rect 11476 -2877 11510 -2843
rect 13500 -2877 13534 -2843
rect 14696 -2877 14730 -2843
rect 15892 -2877 15926 -2843
rect -2232 -3709 -2198 -3675
rect -116 -3709 -82 -3675
rect 344 -3709 378 -3675
rect 1172 -3709 1206 -3675
rect 1632 -3709 1666 -3675
rect 2460 -3709 2494 -3675
rect 2920 -3709 2954 -3675
rect 3748 -3709 3782 -3675
rect 4208 -3709 4242 -3675
rect 5036 -3709 5070 -3675
rect 5496 -3709 5530 -3675
rect 6324 -3709 6358 -3675
rect 6784 -3709 6818 -3675
rect 7612 -3709 7646 -3675
rect 8072 -3709 8106 -3675
rect 8900 -3709 8934 -3675
rect 9360 -3709 9394 -3675
rect 10188 -3709 10222 -3675
rect 11476 -3709 11510 -3675
rect 13500 -3709 13534 -3675
rect 14696 -3709 14730 -3675
rect 15892 -3709 15926 -3675
rect -2232 -3965 -2198 -3931
rect -116 -3965 -82 -3931
rect 344 -3965 378 -3931
rect 1172 -3965 1206 -3931
rect 1632 -3965 1666 -3931
rect 2460 -3965 2494 -3931
rect 2920 -3965 2954 -3931
rect 3748 -3965 3782 -3931
rect 4208 -3965 4242 -3931
rect 5036 -3965 5070 -3931
rect 5496 -3965 5530 -3931
rect 6324 -3965 6358 -3931
rect 6784 -3965 6818 -3931
rect 7612 -3965 7646 -3931
rect 8072 -3965 8106 -3931
rect 8900 -3965 8934 -3931
rect 9360 -3965 9394 -3931
rect 10188 -3965 10222 -3931
rect 11476 -3965 11510 -3931
rect 12396 -3965 12430 -3931
rect 13132 -3965 13166 -3931
rect 13592 -3965 13626 -3931
rect 15524 -3965 15558 -3931
rect -2232 -4797 -2198 -4763
rect -116 -4797 -82 -4763
rect 344 -4797 378 -4763
rect 1172 -4797 1206 -4763
rect 1632 -4797 1666 -4763
rect 2460 -4797 2494 -4763
rect 2920 -4797 2954 -4763
rect 3748 -4797 3782 -4763
rect 4208 -4797 4242 -4763
rect 5036 -4797 5070 -4763
rect 5496 -4797 5530 -4763
rect 6324 -4797 6358 -4763
rect 6784 -4797 6818 -4763
rect 7612 -4797 7646 -4763
rect 8072 -4797 8106 -4763
rect 8900 -4797 8934 -4763
rect 9360 -4797 9394 -4763
rect 10188 -4797 10222 -4763
rect 11476 -4797 11510 -4763
rect 13592 -4797 13626 -4763
rect 15524 -4797 15558 -4763
rect -2232 -5053 -2198 -5019
rect -116 -5053 -82 -5019
rect 344 -5053 378 -5019
rect 1172 -5053 1206 -5019
rect 1632 -5053 1666 -5019
rect 2460 -5053 2494 -5019
rect 2920 -5053 2954 -5019
rect 3748 -5053 3782 -5019
rect 4208 -5053 4242 -5019
rect 5036 -5053 5070 -5019
rect 5496 -5053 5530 -5019
rect 6324 -5053 6358 -5019
rect 6784 -5053 6818 -5019
rect 7612 -5053 7646 -5019
rect 8072 -5053 8106 -5019
rect 8900 -5053 8934 -5019
rect 9360 -5053 9394 -5019
rect 10188 -5053 10222 -5019
rect 11476 -5053 11510 -5019
rect 12396 -5053 12430 -5019
rect 13132 -5053 13166 -5019
rect 13592 -5053 13626 -5019
rect 15524 -5053 15558 -5019
rect -2232 -5885 -2198 -5851
rect -116 -5885 -82 -5851
rect 344 -5885 378 -5851
rect 1172 -5885 1206 -5851
rect 1632 -5885 1666 -5851
rect 2460 -5885 2494 -5851
rect 2920 -5885 2954 -5851
rect 3748 -5885 3782 -5851
rect 4208 -5885 4242 -5851
rect 5036 -5885 5070 -5851
rect 5496 -5885 5530 -5851
rect 6324 -5885 6358 -5851
rect 6784 -5885 6818 -5851
rect 7612 -5885 7646 -5851
rect 8072 -5885 8106 -5851
rect 8900 -5885 8934 -5851
rect 9360 -5885 9394 -5851
rect 10188 -5885 10222 -5851
rect 11476 -5885 11510 -5851
rect 13592 -5885 13626 -5851
rect 15524 -5885 15558 -5851
rect -2232 -6141 -2198 -6107
rect -1036 -6141 -1002 -6107
rect -668 -6141 -634 -6107
rect -208 -6141 -174 -6107
rect 528 -6141 562 -6107
rect 988 -6141 1022 -6107
rect 1356 -6141 1390 -6107
rect 1816 -6141 1850 -6107
rect 2276 -6141 2310 -6107
rect 3104 -6141 3138 -6107
rect 3564 -6141 3598 -6107
rect 6324 -6141 6358 -6107
rect 6784 -6141 6818 -6107
rect 7612 -6141 7646 -6107
rect 8072 -6141 8106 -6107
rect 8900 -6141 8934 -6107
rect 9360 -6141 9394 -6107
rect 10188 -6141 10222 -6107
rect 10648 -6141 10682 -6107
rect 11568 -6141 11602 -6107
rect 13500 -6141 13534 -6107
rect 14696 -6141 14730 -6107
rect 15892 -6141 15926 -6107
rect -2692 -6973 -2658 -6939
rect -116 -6973 -82 -6939
rect 1448 -6973 1482 -6939
rect 3012 -6973 3046 -6939
rect 4576 -6973 4610 -6939
rect 6140 -6973 6174 -6939
rect 7704 -6973 7738 -6939
rect 9268 -6973 9302 -6939
rect 15892 -6973 15926 -6939
rect -2232 -7229 -2198 -7195
rect -116 -7229 -82 -7195
rect 1448 -7229 1482 -7195
rect 2828 -7229 2862 -7195
rect 3196 -7229 3230 -7195
rect 3656 -7229 3690 -7195
rect 4024 -7229 4058 -7195
rect 4484 -7229 4518 -7195
rect 5404 -7229 5438 -7195
rect 5864 -7229 5898 -7195
rect 7704 -7229 7738 -7195
rect 9268 -7229 9302 -7195
rect 15892 -7229 15926 -7195
rect -2232 -8061 -2198 -8027
rect -1036 -8061 -1002 -8027
rect -668 -8061 -634 -8027
rect -208 -8061 -174 -8027
rect 528 -8061 562 -8027
rect 988 -8061 1022 -8027
rect 1356 -8061 1390 -8027
rect 1816 -8061 1850 -8027
rect 2276 -8061 2310 -8027
rect 3104 -8061 3138 -8027
rect 3564 -8061 3598 -8027
rect 6324 -8061 6358 -8027
rect 6784 -8061 6818 -8027
rect 7612 -8061 7646 -8027
rect 8072 -8061 8106 -8027
rect 8900 -8061 8934 -8027
rect 9360 -8061 9394 -8027
rect 10188 -8061 10222 -8027
rect 10648 -8061 10682 -8027
rect 11568 -8061 11602 -8027
rect 13500 -8061 13534 -8027
rect 14696 -8061 14730 -8027
rect 15892 -8061 15926 -8027
rect -2232 -8317 -2198 -8283
rect -116 -8317 -82 -8283
rect 344 -8317 378 -8283
rect 1172 -8317 1206 -8283
rect 1632 -8317 1666 -8283
rect 2460 -8317 2494 -8283
rect 2920 -8317 2954 -8283
rect 3748 -8317 3782 -8283
rect 4208 -8317 4242 -8283
rect 5036 -8317 5070 -8283
rect 5496 -8317 5530 -8283
rect 6324 -8317 6358 -8283
rect 6784 -8317 6818 -8283
rect 7612 -8317 7646 -8283
rect 8072 -8317 8106 -8283
rect 8900 -8317 8934 -8283
rect 9360 -8317 9394 -8283
rect 10188 -8317 10222 -8283
rect 11476 -8317 11510 -8283
rect 13592 -8317 13626 -8283
rect 15524 -8317 15558 -8283
rect -2232 -9149 -2198 -9115
rect -116 -9149 -82 -9115
rect 344 -9149 378 -9115
rect 1172 -9149 1206 -9115
rect 1632 -9149 1666 -9115
rect 2460 -9149 2494 -9115
rect 2920 -9149 2954 -9115
rect 3748 -9149 3782 -9115
rect 4208 -9149 4242 -9115
rect 5036 -9149 5070 -9115
rect 5496 -9149 5530 -9115
rect 6324 -9149 6358 -9115
rect 6784 -9149 6818 -9115
rect 7612 -9149 7646 -9115
rect 8072 -9149 8106 -9115
rect 8900 -9149 8934 -9115
rect 9360 -9149 9394 -9115
rect 10188 -9149 10222 -9115
rect 11476 -9149 11510 -9115
rect 12396 -9149 12430 -9115
rect 13132 -9149 13166 -9115
rect 13592 -9149 13626 -9115
rect 15524 -9149 15558 -9115
rect -2232 -9405 -2198 -9371
rect -116 -9405 -82 -9371
rect 344 -9405 378 -9371
rect 1172 -9405 1206 -9371
rect 1632 -9405 1666 -9371
rect 2460 -9405 2494 -9371
rect 2920 -9405 2954 -9371
rect 3748 -9405 3782 -9371
rect 4208 -9405 4242 -9371
rect 5036 -9405 5070 -9371
rect 5496 -9405 5530 -9371
rect 6324 -9405 6358 -9371
rect 6784 -9405 6818 -9371
rect 7612 -9405 7646 -9371
rect 8072 -9405 8106 -9371
rect 8900 -9405 8934 -9371
rect 9360 -9405 9394 -9371
rect 10188 -9405 10222 -9371
rect 11476 -9405 11510 -9371
rect 13592 -9405 13626 -9371
rect 15524 -9405 15558 -9371
rect -2232 -10237 -2198 -10203
rect -116 -10237 -82 -10203
rect 344 -10237 378 -10203
rect 1172 -10237 1206 -10203
rect 1632 -10237 1666 -10203
rect 2460 -10237 2494 -10203
rect 2920 -10237 2954 -10203
rect 3748 -10237 3782 -10203
rect 4208 -10237 4242 -10203
rect 5036 -10237 5070 -10203
rect 5496 -10237 5530 -10203
rect 6324 -10237 6358 -10203
rect 6784 -10237 6818 -10203
rect 7612 -10237 7646 -10203
rect 8072 -10237 8106 -10203
rect 8900 -10237 8934 -10203
rect 9360 -10237 9394 -10203
rect 10188 -10237 10222 -10203
rect 11476 -10237 11510 -10203
rect 12396 -10237 12430 -10203
rect 13132 -10237 13166 -10203
rect 13592 -10237 13626 -10203
rect 15524 -10237 15558 -10203
rect -2232 -10493 -2198 -10459
rect -1680 -10493 -1646 -10459
rect -116 -10493 -82 -10459
rect 344 -10493 378 -10459
rect 1172 -10493 1206 -10459
rect 1632 -10493 1666 -10459
rect 2460 -10493 2494 -10459
rect 2920 -10493 2954 -10459
rect 3748 -10493 3782 -10459
rect 4208 -10493 4242 -10459
rect 5036 -10493 5070 -10459
rect 5496 -10493 5530 -10459
rect 6324 -10493 6358 -10459
rect 6784 -10493 6818 -10459
rect 7612 -10493 7646 -10459
rect 8072 -10493 8106 -10459
rect 8900 -10493 8934 -10459
rect 9360 -10493 9394 -10459
rect 10188 -10493 10222 -10459
rect 11476 -10493 11510 -10459
rect 13500 -10493 13534 -10459
rect 14696 -10493 14730 -10459
rect 15892 -10493 15926 -10459
rect -2232 -11325 -2198 -11291
rect -116 -11325 -82 -11291
rect 344 -11325 378 -11291
rect 1172 -11325 1206 -11291
rect 1632 -11325 1666 -11291
rect 2460 -11325 2494 -11291
rect 2920 -11325 2954 -11291
rect 3748 -11325 3782 -11291
rect 4208 -11325 4242 -11291
rect 5036 -11325 5070 -11291
rect 5496 -11325 5530 -11291
rect 6324 -11325 6358 -11291
rect 6784 -11325 6818 -11291
rect 7612 -11325 7646 -11291
rect 8072 -11325 8106 -11291
rect 8900 -11325 8934 -11291
rect 9360 -11325 9394 -11291
rect 10188 -11325 10222 -11291
rect 11476 -11325 11510 -11291
rect 13500 -11325 13534 -11291
rect 14696 -11325 14730 -11291
rect 15892 -11325 15926 -11291
rect -2232 -11581 -2198 -11547
rect -116 -11581 -82 -11547
rect 344 -11581 378 -11547
rect 1172 -11581 1206 -11547
rect 1632 -11581 1666 -11547
rect 2460 -11581 2494 -11547
rect 2920 -11581 2954 -11547
rect 3748 -11581 3782 -11547
rect 4208 -11581 4242 -11547
rect 5036 -11581 5070 -11547
rect 5496 -11581 5530 -11547
rect 6324 -11581 6358 -11547
rect 6784 -11581 6818 -11547
rect 7612 -11581 7646 -11547
rect 8072 -11581 8106 -11547
rect 8900 -11581 8934 -11547
rect 9360 -11581 9394 -11547
rect 10188 -11581 10222 -11547
rect 11476 -11581 11510 -11547
rect 12396 -11581 12430 -11547
rect 13132 -11581 13166 -11547
rect 13592 -11581 13626 -11547
rect 15524 -11581 15558 -11547
rect -2232 -12413 -2198 -12379
rect -116 -12413 -82 -12379
rect 344 -12413 378 -12379
rect 1172 -12413 1206 -12379
rect 1632 -12413 1666 -12379
rect 2460 -12413 2494 -12379
rect 2920 -12413 2954 -12379
rect 3748 -12413 3782 -12379
rect 4208 -12413 4242 -12379
rect 5036 -12413 5070 -12379
rect 5496 -12413 5530 -12379
rect 6324 -12413 6358 -12379
rect 6784 -12413 6818 -12379
rect 7612 -12413 7646 -12379
rect 8072 -12413 8106 -12379
rect 8900 -12413 8934 -12379
rect 9360 -12413 9394 -12379
rect 10188 -12413 10222 -12379
rect 11476 -12413 11510 -12379
rect 13592 -12413 13626 -12379
rect 15524 -12413 15558 -12379
rect -2232 -12669 -2198 -12635
rect -116 -12669 -82 -12635
rect 344 -12669 378 -12635
rect 1172 -12669 1206 -12635
rect 1632 -12669 1666 -12635
rect 2460 -12669 2494 -12635
rect 2920 -12669 2954 -12635
rect 3748 -12669 3782 -12635
rect 4208 -12669 4242 -12635
rect 5036 -12669 5070 -12635
rect 5496 -12669 5530 -12635
rect 6324 -12669 6358 -12635
rect 6784 -12669 6818 -12635
rect 7612 -12669 7646 -12635
rect 8072 -12669 8106 -12635
rect 8900 -12669 8934 -12635
rect 9360 -12669 9394 -12635
rect 10188 -12669 10222 -12635
rect 11476 -12669 11510 -12635
rect 12396 -12669 12430 -12635
rect 13132 -12669 13166 -12635
rect 13592 -12669 13626 -12635
rect 15524 -12669 15558 -12635
rect -2232 -13501 -2198 -13467
rect -116 -13501 -82 -13467
rect 344 -13501 378 -13467
rect 1172 -13501 1206 -13467
rect 1632 -13501 1666 -13467
rect 2460 -13501 2494 -13467
rect 2920 -13501 2954 -13467
rect 3748 -13501 3782 -13467
rect 4208 -13501 4242 -13467
rect 5036 -13501 5070 -13467
rect 5496 -13501 5530 -13467
rect 6324 -13501 6358 -13467
rect 6784 -13501 6818 -13467
rect 7612 -13501 7646 -13467
rect 8072 -13501 8106 -13467
rect 8900 -13501 8934 -13467
rect 9360 -13501 9394 -13467
rect 10188 -13501 10222 -13467
rect 11476 -13501 11510 -13467
rect 13592 -13501 13626 -13467
rect 15524 -13501 15558 -13467
rect -2232 -13757 -2198 -13723
rect -1036 -13757 -1002 -13723
rect -668 -13757 -634 -13723
rect -208 -13757 -174 -13723
rect 528 -13757 562 -13723
rect 988 -13757 1022 -13723
rect 1356 -13757 1390 -13723
rect 1816 -13757 1850 -13723
rect 2276 -13757 2310 -13723
rect 3104 -13757 3138 -13723
rect 3564 -13757 3598 -13723
rect 6324 -13757 6358 -13723
rect 6784 -13757 6818 -13723
rect 7612 -13757 7646 -13723
rect 8072 -13757 8106 -13723
rect 8900 -13757 8934 -13723
rect 9360 -13757 9394 -13723
rect 10188 -13757 10222 -13723
rect 10648 -13757 10682 -13723
rect 11568 -13757 11602 -13723
rect 13500 -13757 13534 -13723
rect 14696 -13757 14730 -13723
rect 15892 -13757 15926 -13723
<< nsubdiffcont >>
rect -2232 -134 -2198 -100
rect -2232 -227 -2198 -193
rect -1036 -134 -1002 -100
rect -1036 -227 -1002 -193
rect -668 -134 -634 -100
rect -668 -227 -634 -193
rect -208 -134 -174 -100
rect -208 -227 -174 -193
rect 528 -134 562 -100
rect 528 -227 562 -193
rect 988 -134 1022 -100
rect 988 -227 1022 -193
rect 1356 -134 1390 -100
rect 1356 -227 1390 -193
rect 1816 -134 1850 -100
rect 1816 -227 1850 -193
rect 2276 -134 2310 -100
rect 2276 -227 2310 -193
rect 3104 -134 3138 -100
rect 3104 -227 3138 -193
rect 3564 -134 3598 -100
rect 3564 -227 3598 -193
rect 6324 -134 6358 -100
rect 6324 -227 6358 -193
rect 6784 -134 6818 -100
rect 6784 -227 6818 -193
rect 7612 -134 7646 -100
rect 7612 -227 7646 -193
rect 8072 -134 8106 -100
rect 8072 -227 8106 -193
rect 8900 -134 8934 -100
rect 8900 -227 8934 -193
rect 9360 -134 9394 -100
rect 9360 -227 9394 -193
rect 10188 -134 10222 -100
rect 10188 -227 10222 -193
rect 10648 -134 10682 -100
rect 10648 -227 10682 -193
rect 11568 -134 11602 -100
rect 11568 -227 11602 -193
rect 13500 -134 13534 -100
rect 13500 -227 13534 -193
rect 14696 -134 14730 -100
rect 14696 -227 14730 -193
rect 15892 -134 15926 -100
rect 15892 -227 15926 -193
rect -2232 -919 -2198 -885
rect -2232 -1012 -2198 -978
rect -116 -919 -82 -885
rect -116 -1012 -82 -978
rect 344 -919 378 -885
rect 344 -1012 378 -978
rect 1172 -919 1206 -885
rect 1172 -1012 1206 -978
rect 1632 -919 1666 -885
rect 1632 -1012 1666 -978
rect 2460 -919 2494 -885
rect 2460 -1012 2494 -978
rect 2920 -919 2954 -885
rect 2920 -1012 2954 -978
rect 3748 -919 3782 -885
rect 3748 -1012 3782 -978
rect 4208 -919 4242 -885
rect 4208 -1012 4242 -978
rect 5036 -919 5070 -885
rect 5036 -1012 5070 -978
rect 5496 -919 5530 -885
rect 5496 -1012 5530 -978
rect 6324 -919 6358 -885
rect 6324 -1012 6358 -978
rect 6784 -919 6818 -885
rect 6784 -1012 6818 -978
rect 7612 -919 7646 -885
rect 7612 -1012 7646 -978
rect 8072 -919 8106 -885
rect 8072 -1012 8106 -978
rect 8900 -919 8934 -885
rect 8900 -1012 8934 -978
rect 9360 -919 9394 -885
rect 9360 -1012 9394 -978
rect 10188 -919 10222 -885
rect 10188 -1012 10222 -978
rect 11476 -919 11510 -885
rect 11476 -1012 11510 -978
rect 13592 -919 13626 -885
rect 13592 -1012 13626 -978
rect 15524 -919 15558 -885
rect 15524 -1012 15558 -978
rect -2232 -1222 -2198 -1188
rect -2232 -1315 -2198 -1281
rect -116 -1222 -82 -1188
rect -116 -1315 -82 -1281
rect 344 -1222 378 -1188
rect 344 -1315 378 -1281
rect 1172 -1222 1206 -1188
rect 1172 -1315 1206 -1281
rect 1632 -1222 1666 -1188
rect 1632 -1315 1666 -1281
rect 2460 -1222 2494 -1188
rect 2460 -1315 2494 -1281
rect 2920 -1222 2954 -1188
rect 2920 -1315 2954 -1281
rect 3748 -1222 3782 -1188
rect 3748 -1315 3782 -1281
rect 4208 -1222 4242 -1188
rect 4208 -1315 4242 -1281
rect 5036 -1222 5070 -1188
rect 5036 -1315 5070 -1281
rect 5496 -1222 5530 -1188
rect 5496 -1315 5530 -1281
rect 6324 -1222 6358 -1188
rect 6324 -1315 6358 -1281
rect 6784 -1222 6818 -1188
rect 6784 -1315 6818 -1281
rect 7612 -1222 7646 -1188
rect 7612 -1315 7646 -1281
rect 8072 -1222 8106 -1188
rect 8072 -1315 8106 -1281
rect 8900 -1222 8934 -1188
rect 8900 -1315 8934 -1281
rect 9360 -1222 9394 -1188
rect 9360 -1315 9394 -1281
rect 10188 -1222 10222 -1188
rect 10188 -1315 10222 -1281
rect 11476 -1222 11510 -1188
rect 11476 -1315 11510 -1281
rect 12396 -1222 12430 -1188
rect 12396 -1315 12430 -1281
rect 13132 -1222 13166 -1188
rect 13132 -1315 13166 -1281
rect 13592 -1222 13626 -1188
rect 13592 -1315 13626 -1281
rect 15524 -1222 15558 -1188
rect 15524 -1315 15558 -1281
rect -2232 -2007 -2198 -1973
rect -2232 -2100 -2198 -2066
rect -116 -2007 -82 -1973
rect -116 -2100 -82 -2066
rect 344 -2007 378 -1973
rect 344 -2100 378 -2066
rect 1172 -2007 1206 -1973
rect 1172 -2100 1206 -2066
rect 1632 -2007 1666 -1973
rect 1632 -2100 1666 -2066
rect 2460 -2007 2494 -1973
rect 2460 -2100 2494 -2066
rect 2920 -2007 2954 -1973
rect 2920 -2100 2954 -2066
rect 3748 -2007 3782 -1973
rect 3748 -2100 3782 -2066
rect 4208 -2007 4242 -1973
rect 4208 -2100 4242 -2066
rect 5036 -2007 5070 -1973
rect 5036 -2100 5070 -2066
rect 5496 -2007 5530 -1973
rect 5496 -2100 5530 -2066
rect 6324 -2007 6358 -1973
rect 6324 -2100 6358 -2066
rect 6784 -2007 6818 -1973
rect 6784 -2100 6818 -2066
rect 7612 -2007 7646 -1973
rect 7612 -2100 7646 -2066
rect 8072 -2007 8106 -1973
rect 8072 -2100 8106 -2066
rect 8900 -2007 8934 -1973
rect 8900 -2100 8934 -2066
rect 9360 -2007 9394 -1973
rect 9360 -2100 9394 -2066
rect 10188 -2007 10222 -1973
rect 10188 -2100 10222 -2066
rect 11476 -2007 11510 -1973
rect 11476 -2100 11510 -2066
rect 13592 -2007 13626 -1973
rect 13592 -2100 13626 -2066
rect 15524 -2007 15558 -1973
rect 15524 -2100 15558 -2066
rect -2232 -2310 -2198 -2276
rect -2232 -2403 -2198 -2369
rect -116 -2310 -82 -2276
rect -116 -2403 -82 -2369
rect 344 -2310 378 -2276
rect 344 -2403 378 -2369
rect 1172 -2310 1206 -2276
rect 1172 -2403 1206 -2369
rect 1632 -2310 1666 -2276
rect 1632 -2403 1666 -2369
rect 2460 -2310 2494 -2276
rect 2460 -2403 2494 -2369
rect 2920 -2310 2954 -2276
rect 2920 -2403 2954 -2369
rect 3748 -2310 3782 -2276
rect 3748 -2403 3782 -2369
rect 4208 -2310 4242 -2276
rect 4208 -2403 4242 -2369
rect 5036 -2310 5070 -2276
rect 5036 -2403 5070 -2369
rect 5496 -2310 5530 -2276
rect 5496 -2403 5530 -2369
rect 6324 -2310 6358 -2276
rect 6324 -2403 6358 -2369
rect 6784 -2310 6818 -2276
rect 6784 -2403 6818 -2369
rect 7612 -2310 7646 -2276
rect 7612 -2403 7646 -2369
rect 8072 -2310 8106 -2276
rect 8072 -2403 8106 -2369
rect 8900 -2310 8934 -2276
rect 8900 -2403 8934 -2369
rect 9360 -2310 9394 -2276
rect 9360 -2403 9394 -2369
rect 10188 -2310 10222 -2276
rect 10188 -2403 10222 -2369
rect 11476 -2310 11510 -2276
rect 11476 -2403 11510 -2369
rect 12396 -2310 12430 -2276
rect 12396 -2403 12430 -2369
rect 13132 -2310 13166 -2276
rect 13132 -2403 13166 -2369
rect 13592 -2310 13626 -2276
rect 13592 -2403 13626 -2369
rect 15524 -2310 15558 -2276
rect 15524 -2403 15558 -2369
rect -2232 -3095 -2198 -3061
rect -2232 -3188 -2198 -3154
rect -1680 -3095 -1646 -3061
rect -1680 -3188 -1646 -3154
rect -116 -3095 -82 -3061
rect -116 -3188 -82 -3154
rect 344 -3095 378 -3061
rect 344 -3188 378 -3154
rect 1172 -3095 1206 -3061
rect 1172 -3188 1206 -3154
rect 1632 -3095 1666 -3061
rect 1632 -3188 1666 -3154
rect 2460 -3095 2494 -3061
rect 2460 -3188 2494 -3154
rect 2920 -3095 2954 -3061
rect 2920 -3188 2954 -3154
rect 3748 -3095 3782 -3061
rect 3748 -3188 3782 -3154
rect 4208 -3095 4242 -3061
rect 4208 -3188 4242 -3154
rect 5036 -3095 5070 -3061
rect 5036 -3188 5070 -3154
rect 5496 -3095 5530 -3061
rect 5496 -3188 5530 -3154
rect 6324 -3095 6358 -3061
rect 6324 -3188 6358 -3154
rect 6784 -3095 6818 -3061
rect 6784 -3188 6818 -3154
rect 7612 -3095 7646 -3061
rect 7612 -3188 7646 -3154
rect 8072 -3095 8106 -3061
rect 8072 -3188 8106 -3154
rect 8900 -3095 8934 -3061
rect 8900 -3188 8934 -3154
rect 9360 -3095 9394 -3061
rect 9360 -3188 9394 -3154
rect 10188 -3095 10222 -3061
rect 10188 -3188 10222 -3154
rect 11476 -3095 11510 -3061
rect 11476 -3188 11510 -3154
rect 13500 -3095 13534 -3061
rect 13500 -3188 13534 -3154
rect 14696 -3095 14730 -3061
rect 14696 -3188 14730 -3154
rect 15892 -3095 15926 -3061
rect 15892 -3188 15926 -3154
rect -2232 -3398 -2198 -3364
rect -2232 -3491 -2198 -3457
rect -116 -3398 -82 -3364
rect -116 -3491 -82 -3457
rect 344 -3398 378 -3364
rect 344 -3491 378 -3457
rect 1172 -3398 1206 -3364
rect 1172 -3491 1206 -3457
rect 1632 -3398 1666 -3364
rect 1632 -3491 1666 -3457
rect 2460 -3398 2494 -3364
rect 2460 -3491 2494 -3457
rect 2920 -3398 2954 -3364
rect 2920 -3491 2954 -3457
rect 3748 -3398 3782 -3364
rect 3748 -3491 3782 -3457
rect 4208 -3398 4242 -3364
rect 4208 -3491 4242 -3457
rect 5036 -3398 5070 -3364
rect 5036 -3491 5070 -3457
rect 5496 -3398 5530 -3364
rect 5496 -3491 5530 -3457
rect 6324 -3398 6358 -3364
rect 6324 -3491 6358 -3457
rect 6784 -3398 6818 -3364
rect 6784 -3491 6818 -3457
rect 7612 -3398 7646 -3364
rect 7612 -3491 7646 -3457
rect 8072 -3398 8106 -3364
rect 8072 -3491 8106 -3457
rect 8900 -3398 8934 -3364
rect 8900 -3491 8934 -3457
rect 9360 -3398 9394 -3364
rect 9360 -3491 9394 -3457
rect 10188 -3398 10222 -3364
rect 10188 -3491 10222 -3457
rect 11476 -3398 11510 -3364
rect 11476 -3491 11510 -3457
rect 13500 -3398 13534 -3364
rect 13500 -3491 13534 -3457
rect 14696 -3398 14730 -3364
rect 14696 -3491 14730 -3457
rect 15892 -3398 15926 -3364
rect 15892 -3491 15926 -3457
rect -2232 -4183 -2198 -4149
rect -2232 -4276 -2198 -4242
rect -116 -4183 -82 -4149
rect -116 -4276 -82 -4242
rect 344 -4183 378 -4149
rect 344 -4276 378 -4242
rect 1172 -4183 1206 -4149
rect 1172 -4276 1206 -4242
rect 1632 -4183 1666 -4149
rect 1632 -4276 1666 -4242
rect 2460 -4183 2494 -4149
rect 2460 -4276 2494 -4242
rect 2920 -4183 2954 -4149
rect 2920 -4276 2954 -4242
rect 3748 -4183 3782 -4149
rect 3748 -4276 3782 -4242
rect 4208 -4183 4242 -4149
rect 4208 -4276 4242 -4242
rect 5036 -4183 5070 -4149
rect 5036 -4276 5070 -4242
rect 5496 -4183 5530 -4149
rect 5496 -4276 5530 -4242
rect 6324 -4183 6358 -4149
rect 6324 -4276 6358 -4242
rect 6784 -4183 6818 -4149
rect 6784 -4276 6818 -4242
rect 7612 -4183 7646 -4149
rect 7612 -4276 7646 -4242
rect 8072 -4183 8106 -4149
rect 8072 -4276 8106 -4242
rect 8900 -4183 8934 -4149
rect 8900 -4276 8934 -4242
rect 9360 -4183 9394 -4149
rect 9360 -4276 9394 -4242
rect 10188 -4183 10222 -4149
rect 10188 -4276 10222 -4242
rect 11476 -4183 11510 -4149
rect 11476 -4276 11510 -4242
rect 12396 -4183 12430 -4149
rect 12396 -4276 12430 -4242
rect 13132 -4183 13166 -4149
rect 13132 -4276 13166 -4242
rect 13592 -4183 13626 -4149
rect 13592 -4276 13626 -4242
rect 15524 -4183 15558 -4149
rect 15524 -4276 15558 -4242
rect -2232 -4486 -2198 -4452
rect -2232 -4579 -2198 -4545
rect -116 -4486 -82 -4452
rect -116 -4579 -82 -4545
rect 344 -4486 378 -4452
rect 344 -4579 378 -4545
rect 1172 -4486 1206 -4452
rect 1172 -4579 1206 -4545
rect 1632 -4486 1666 -4452
rect 1632 -4579 1666 -4545
rect 2460 -4486 2494 -4452
rect 2460 -4579 2494 -4545
rect 2920 -4486 2954 -4452
rect 2920 -4579 2954 -4545
rect 3748 -4486 3782 -4452
rect 3748 -4579 3782 -4545
rect 4208 -4486 4242 -4452
rect 4208 -4579 4242 -4545
rect 5036 -4486 5070 -4452
rect 5036 -4579 5070 -4545
rect 5496 -4486 5530 -4452
rect 5496 -4579 5530 -4545
rect 6324 -4486 6358 -4452
rect 6324 -4579 6358 -4545
rect 6784 -4486 6818 -4452
rect 6784 -4579 6818 -4545
rect 7612 -4486 7646 -4452
rect 7612 -4579 7646 -4545
rect 8072 -4486 8106 -4452
rect 8072 -4579 8106 -4545
rect 8900 -4486 8934 -4452
rect 8900 -4579 8934 -4545
rect 9360 -4486 9394 -4452
rect 9360 -4579 9394 -4545
rect 10188 -4486 10222 -4452
rect 10188 -4579 10222 -4545
rect 11476 -4486 11510 -4452
rect 11476 -4579 11510 -4545
rect 13592 -4486 13626 -4452
rect 13592 -4579 13626 -4545
rect 15524 -4486 15558 -4452
rect 15524 -4579 15558 -4545
rect -2232 -5271 -2198 -5237
rect -2232 -5364 -2198 -5330
rect -116 -5271 -82 -5237
rect -116 -5364 -82 -5330
rect 344 -5271 378 -5237
rect 344 -5364 378 -5330
rect 1172 -5271 1206 -5237
rect 1172 -5364 1206 -5330
rect 1632 -5271 1666 -5237
rect 1632 -5364 1666 -5330
rect 2460 -5271 2494 -5237
rect 2460 -5364 2494 -5330
rect 2920 -5271 2954 -5237
rect 2920 -5364 2954 -5330
rect 3748 -5271 3782 -5237
rect 3748 -5364 3782 -5330
rect 4208 -5271 4242 -5237
rect 4208 -5364 4242 -5330
rect 5036 -5271 5070 -5237
rect 5036 -5364 5070 -5330
rect 5496 -5271 5530 -5237
rect 5496 -5364 5530 -5330
rect 6324 -5271 6358 -5237
rect 6324 -5364 6358 -5330
rect 6784 -5271 6818 -5237
rect 6784 -5364 6818 -5330
rect 7612 -5271 7646 -5237
rect 7612 -5364 7646 -5330
rect 8072 -5271 8106 -5237
rect 8072 -5364 8106 -5330
rect 8900 -5271 8934 -5237
rect 8900 -5364 8934 -5330
rect 9360 -5271 9394 -5237
rect 9360 -5364 9394 -5330
rect 10188 -5271 10222 -5237
rect 10188 -5364 10222 -5330
rect 11476 -5271 11510 -5237
rect 11476 -5364 11510 -5330
rect 12396 -5271 12430 -5237
rect 12396 -5364 12430 -5330
rect 13132 -5271 13166 -5237
rect 13132 -5364 13166 -5330
rect 13592 -5271 13626 -5237
rect 13592 -5364 13626 -5330
rect 15524 -5271 15558 -5237
rect 15524 -5364 15558 -5330
rect -2232 -5574 -2198 -5540
rect -2232 -5667 -2198 -5633
rect -116 -5574 -82 -5540
rect -116 -5667 -82 -5633
rect 344 -5574 378 -5540
rect 344 -5667 378 -5633
rect 1172 -5574 1206 -5540
rect 1172 -5667 1206 -5633
rect 1632 -5574 1666 -5540
rect 1632 -5667 1666 -5633
rect 2460 -5574 2494 -5540
rect 2460 -5667 2494 -5633
rect 2920 -5574 2954 -5540
rect 2920 -5667 2954 -5633
rect 3748 -5574 3782 -5540
rect 3748 -5667 3782 -5633
rect 4208 -5574 4242 -5540
rect 4208 -5667 4242 -5633
rect 5036 -5574 5070 -5540
rect 5036 -5667 5070 -5633
rect 5496 -5574 5530 -5540
rect 5496 -5667 5530 -5633
rect 6324 -5574 6358 -5540
rect 6324 -5667 6358 -5633
rect 6784 -5574 6818 -5540
rect 6784 -5667 6818 -5633
rect 7612 -5574 7646 -5540
rect 7612 -5667 7646 -5633
rect 8072 -5574 8106 -5540
rect 8072 -5667 8106 -5633
rect 8900 -5574 8934 -5540
rect 8900 -5667 8934 -5633
rect 9360 -5574 9394 -5540
rect 9360 -5667 9394 -5633
rect 10188 -5574 10222 -5540
rect 10188 -5667 10222 -5633
rect 11476 -5574 11510 -5540
rect 11476 -5667 11510 -5633
rect 13592 -5574 13626 -5540
rect 13592 -5667 13626 -5633
rect 15524 -5574 15558 -5540
rect 15524 -5667 15558 -5633
rect -2232 -6359 -2198 -6325
rect -2232 -6452 -2198 -6418
rect -1036 -6359 -1002 -6325
rect -1036 -6452 -1002 -6418
rect -668 -6359 -634 -6325
rect -668 -6452 -634 -6418
rect -208 -6359 -174 -6325
rect -208 -6452 -174 -6418
rect 528 -6359 562 -6325
rect 528 -6452 562 -6418
rect 988 -6359 1022 -6325
rect 988 -6452 1022 -6418
rect 1356 -6359 1390 -6325
rect 1356 -6452 1390 -6418
rect 1816 -6359 1850 -6325
rect 1816 -6452 1850 -6418
rect 2276 -6359 2310 -6325
rect 2276 -6452 2310 -6418
rect 3104 -6359 3138 -6325
rect 3104 -6452 3138 -6418
rect 3564 -6359 3598 -6325
rect 3564 -6452 3598 -6418
rect 6324 -6359 6358 -6325
rect 6324 -6452 6358 -6418
rect 6784 -6359 6818 -6325
rect 6784 -6452 6818 -6418
rect 7612 -6359 7646 -6325
rect 7612 -6452 7646 -6418
rect 8072 -6359 8106 -6325
rect 8072 -6452 8106 -6418
rect 8900 -6359 8934 -6325
rect 8900 -6452 8934 -6418
rect 9360 -6359 9394 -6325
rect 9360 -6452 9394 -6418
rect 10188 -6359 10222 -6325
rect 10188 -6452 10222 -6418
rect 10648 -6359 10682 -6325
rect 10648 -6452 10682 -6418
rect 11568 -6359 11602 -6325
rect 11568 -6452 11602 -6418
rect 13500 -6359 13534 -6325
rect 13500 -6452 13534 -6418
rect 14696 -6359 14730 -6325
rect 14696 -6452 14730 -6418
rect 15892 -6359 15926 -6325
rect 15892 -6452 15926 -6418
rect -2692 -6662 -2658 -6628
rect -2692 -6755 -2658 -6721
rect -116 -6662 -82 -6628
rect -116 -6755 -82 -6721
rect 1448 -6662 1482 -6628
rect 1448 -6755 1482 -6721
rect 3012 -6662 3046 -6628
rect 3012 -6755 3046 -6721
rect 4576 -6662 4610 -6628
rect 4576 -6755 4610 -6721
rect 6140 -6662 6174 -6628
rect 6140 -6755 6174 -6721
rect 7704 -6662 7738 -6628
rect 7704 -6755 7738 -6721
rect 9268 -6662 9302 -6628
rect 9268 -6755 9302 -6721
rect 15892 -6662 15926 -6628
rect 15892 -6755 15926 -6721
rect -2232 -7447 -2198 -7413
rect -2232 -7540 -2198 -7506
rect -116 -7447 -82 -7413
rect -116 -7540 -82 -7506
rect 1448 -7447 1482 -7413
rect 1448 -7540 1482 -7506
rect 2828 -7447 2862 -7413
rect 2828 -7540 2862 -7506
rect 3196 -7447 3230 -7413
rect 3196 -7540 3230 -7506
rect 3656 -7447 3690 -7413
rect 3656 -7540 3690 -7506
rect 4024 -7447 4058 -7413
rect 4024 -7540 4058 -7506
rect 4484 -7447 4518 -7413
rect 4484 -7540 4518 -7506
rect 5404 -7447 5438 -7413
rect 5404 -7540 5438 -7506
rect 5864 -7447 5898 -7413
rect 5864 -7540 5898 -7506
rect 7704 -7447 7738 -7413
rect 7704 -7540 7738 -7506
rect 9268 -7447 9302 -7413
rect 9268 -7540 9302 -7506
rect 15892 -7447 15926 -7413
rect 15892 -7540 15926 -7506
rect -2232 -7750 -2198 -7716
rect -2232 -7843 -2198 -7809
rect -1036 -7750 -1002 -7716
rect -1036 -7843 -1002 -7809
rect -668 -7750 -634 -7716
rect -668 -7843 -634 -7809
rect -208 -7750 -174 -7716
rect -208 -7843 -174 -7809
rect 528 -7750 562 -7716
rect 528 -7843 562 -7809
rect 988 -7750 1022 -7716
rect 988 -7843 1022 -7809
rect 1356 -7750 1390 -7716
rect 1356 -7843 1390 -7809
rect 1816 -7750 1850 -7716
rect 1816 -7843 1850 -7809
rect 2276 -7750 2310 -7716
rect 2276 -7843 2310 -7809
rect 3104 -7750 3138 -7716
rect 3104 -7843 3138 -7809
rect 3564 -7750 3598 -7716
rect 3564 -7843 3598 -7809
rect 6324 -7750 6358 -7716
rect 6324 -7843 6358 -7809
rect 6784 -7750 6818 -7716
rect 6784 -7843 6818 -7809
rect 7612 -7750 7646 -7716
rect 7612 -7843 7646 -7809
rect 8072 -7750 8106 -7716
rect 8072 -7843 8106 -7809
rect 8900 -7750 8934 -7716
rect 8900 -7843 8934 -7809
rect 9360 -7750 9394 -7716
rect 9360 -7843 9394 -7809
rect 10188 -7750 10222 -7716
rect 10188 -7843 10222 -7809
rect 10648 -7750 10682 -7716
rect 10648 -7843 10682 -7809
rect 11568 -7750 11602 -7716
rect 11568 -7843 11602 -7809
rect 13500 -7750 13534 -7716
rect 13500 -7843 13534 -7809
rect 14696 -7750 14730 -7716
rect 14696 -7843 14730 -7809
rect 15892 -7750 15926 -7716
rect 15892 -7843 15926 -7809
rect -2232 -8535 -2198 -8501
rect -2232 -8628 -2198 -8594
rect -116 -8535 -82 -8501
rect -116 -8628 -82 -8594
rect 344 -8535 378 -8501
rect 344 -8628 378 -8594
rect 1172 -8535 1206 -8501
rect 1172 -8628 1206 -8594
rect 1632 -8535 1666 -8501
rect 1632 -8628 1666 -8594
rect 2460 -8535 2494 -8501
rect 2460 -8628 2494 -8594
rect 2920 -8535 2954 -8501
rect 2920 -8628 2954 -8594
rect 3748 -8535 3782 -8501
rect 3748 -8628 3782 -8594
rect 4208 -8535 4242 -8501
rect 4208 -8628 4242 -8594
rect 5036 -8535 5070 -8501
rect 5036 -8628 5070 -8594
rect 5496 -8535 5530 -8501
rect 5496 -8628 5530 -8594
rect 6324 -8535 6358 -8501
rect 6324 -8628 6358 -8594
rect 6784 -8535 6818 -8501
rect 6784 -8628 6818 -8594
rect 7612 -8535 7646 -8501
rect 7612 -8628 7646 -8594
rect 8072 -8535 8106 -8501
rect 8072 -8628 8106 -8594
rect 8900 -8535 8934 -8501
rect 8900 -8628 8934 -8594
rect 9360 -8535 9394 -8501
rect 9360 -8628 9394 -8594
rect 10188 -8535 10222 -8501
rect 10188 -8628 10222 -8594
rect 11476 -8535 11510 -8501
rect 11476 -8628 11510 -8594
rect 13592 -8535 13626 -8501
rect 13592 -8628 13626 -8594
rect 15524 -8535 15558 -8501
rect 15524 -8628 15558 -8594
rect -2232 -8838 -2198 -8804
rect -2232 -8931 -2198 -8897
rect -116 -8838 -82 -8804
rect -116 -8931 -82 -8897
rect 344 -8838 378 -8804
rect 344 -8931 378 -8897
rect 1172 -8838 1206 -8804
rect 1172 -8931 1206 -8897
rect 1632 -8838 1666 -8804
rect 1632 -8931 1666 -8897
rect 2460 -8838 2494 -8804
rect 2460 -8931 2494 -8897
rect 2920 -8838 2954 -8804
rect 2920 -8931 2954 -8897
rect 3748 -8838 3782 -8804
rect 3748 -8931 3782 -8897
rect 4208 -8838 4242 -8804
rect 4208 -8931 4242 -8897
rect 5036 -8838 5070 -8804
rect 5036 -8931 5070 -8897
rect 5496 -8838 5530 -8804
rect 5496 -8931 5530 -8897
rect 6324 -8838 6358 -8804
rect 6324 -8931 6358 -8897
rect 6784 -8838 6818 -8804
rect 6784 -8931 6818 -8897
rect 7612 -8838 7646 -8804
rect 7612 -8931 7646 -8897
rect 8072 -8838 8106 -8804
rect 8072 -8931 8106 -8897
rect 8900 -8838 8934 -8804
rect 8900 -8931 8934 -8897
rect 9360 -8838 9394 -8804
rect 9360 -8931 9394 -8897
rect 10188 -8838 10222 -8804
rect 10188 -8931 10222 -8897
rect 11476 -8838 11510 -8804
rect 11476 -8931 11510 -8897
rect 12396 -8838 12430 -8804
rect 12396 -8931 12430 -8897
rect 13132 -8838 13166 -8804
rect 13132 -8931 13166 -8897
rect 13592 -8838 13626 -8804
rect 13592 -8931 13626 -8897
rect 15524 -8838 15558 -8804
rect 15524 -8931 15558 -8897
rect -2232 -9623 -2198 -9589
rect -2232 -9716 -2198 -9682
rect -116 -9623 -82 -9589
rect -116 -9716 -82 -9682
rect 344 -9623 378 -9589
rect 344 -9716 378 -9682
rect 1172 -9623 1206 -9589
rect 1172 -9716 1206 -9682
rect 1632 -9623 1666 -9589
rect 1632 -9716 1666 -9682
rect 2460 -9623 2494 -9589
rect 2460 -9716 2494 -9682
rect 2920 -9623 2954 -9589
rect 2920 -9716 2954 -9682
rect 3748 -9623 3782 -9589
rect 3748 -9716 3782 -9682
rect 4208 -9623 4242 -9589
rect 4208 -9716 4242 -9682
rect 5036 -9623 5070 -9589
rect 5036 -9716 5070 -9682
rect 5496 -9623 5530 -9589
rect 5496 -9716 5530 -9682
rect 6324 -9623 6358 -9589
rect 6324 -9716 6358 -9682
rect 6784 -9623 6818 -9589
rect 6784 -9716 6818 -9682
rect 7612 -9623 7646 -9589
rect 7612 -9716 7646 -9682
rect 8072 -9623 8106 -9589
rect 8072 -9716 8106 -9682
rect 8900 -9623 8934 -9589
rect 8900 -9716 8934 -9682
rect 9360 -9623 9394 -9589
rect 9360 -9716 9394 -9682
rect 10188 -9623 10222 -9589
rect 10188 -9716 10222 -9682
rect 11476 -9623 11510 -9589
rect 11476 -9716 11510 -9682
rect 13592 -9623 13626 -9589
rect 13592 -9716 13626 -9682
rect 15524 -9623 15558 -9589
rect 15524 -9716 15558 -9682
rect -2232 -9926 -2198 -9892
rect -2232 -10019 -2198 -9985
rect -116 -9926 -82 -9892
rect -116 -10019 -82 -9985
rect 344 -9926 378 -9892
rect 344 -10019 378 -9985
rect 1172 -9926 1206 -9892
rect 1172 -10019 1206 -9985
rect 1632 -9926 1666 -9892
rect 1632 -10019 1666 -9985
rect 2460 -9926 2494 -9892
rect 2460 -10019 2494 -9985
rect 2920 -9926 2954 -9892
rect 2920 -10019 2954 -9985
rect 3748 -9926 3782 -9892
rect 3748 -10019 3782 -9985
rect 4208 -9926 4242 -9892
rect 4208 -10019 4242 -9985
rect 5036 -9926 5070 -9892
rect 5036 -10019 5070 -9985
rect 5496 -9926 5530 -9892
rect 5496 -10019 5530 -9985
rect 6324 -9926 6358 -9892
rect 6324 -10019 6358 -9985
rect 6784 -9926 6818 -9892
rect 6784 -10019 6818 -9985
rect 7612 -9926 7646 -9892
rect 7612 -10019 7646 -9985
rect 8072 -9926 8106 -9892
rect 8072 -10019 8106 -9985
rect 8900 -9926 8934 -9892
rect 8900 -10019 8934 -9985
rect 9360 -9926 9394 -9892
rect 9360 -10019 9394 -9985
rect 10188 -9926 10222 -9892
rect 10188 -10019 10222 -9985
rect 11476 -9926 11510 -9892
rect 11476 -10019 11510 -9985
rect 12396 -9926 12430 -9892
rect 12396 -10019 12430 -9985
rect 13132 -9926 13166 -9892
rect 13132 -10019 13166 -9985
rect 13592 -9926 13626 -9892
rect 13592 -10019 13626 -9985
rect 15524 -9926 15558 -9892
rect 15524 -10019 15558 -9985
rect -2232 -10711 -2198 -10677
rect -2232 -10804 -2198 -10770
rect -1680 -10711 -1646 -10677
rect -1680 -10804 -1646 -10770
rect -116 -10711 -82 -10677
rect -116 -10804 -82 -10770
rect 344 -10711 378 -10677
rect 344 -10804 378 -10770
rect 1172 -10711 1206 -10677
rect 1172 -10804 1206 -10770
rect 1632 -10711 1666 -10677
rect 1632 -10804 1666 -10770
rect 2460 -10711 2494 -10677
rect 2460 -10804 2494 -10770
rect 2920 -10711 2954 -10677
rect 2920 -10804 2954 -10770
rect 3748 -10711 3782 -10677
rect 3748 -10804 3782 -10770
rect 4208 -10711 4242 -10677
rect 4208 -10804 4242 -10770
rect 5036 -10711 5070 -10677
rect 5036 -10804 5070 -10770
rect 5496 -10711 5530 -10677
rect 5496 -10804 5530 -10770
rect 6324 -10711 6358 -10677
rect 6324 -10804 6358 -10770
rect 6784 -10711 6818 -10677
rect 6784 -10804 6818 -10770
rect 7612 -10711 7646 -10677
rect 7612 -10804 7646 -10770
rect 8072 -10711 8106 -10677
rect 8072 -10804 8106 -10770
rect 8900 -10711 8934 -10677
rect 8900 -10804 8934 -10770
rect 9360 -10711 9394 -10677
rect 9360 -10804 9394 -10770
rect 10188 -10711 10222 -10677
rect 10188 -10804 10222 -10770
rect 11476 -10711 11510 -10677
rect 11476 -10804 11510 -10770
rect 13500 -10711 13534 -10677
rect 13500 -10804 13534 -10770
rect 14696 -10711 14730 -10677
rect 14696 -10804 14730 -10770
rect 15892 -10711 15926 -10677
rect 15892 -10804 15926 -10770
rect -2232 -11014 -2198 -10980
rect -2232 -11107 -2198 -11073
rect -116 -11014 -82 -10980
rect -116 -11107 -82 -11073
rect 344 -11014 378 -10980
rect 344 -11107 378 -11073
rect 1172 -11014 1206 -10980
rect 1172 -11107 1206 -11073
rect 1632 -11014 1666 -10980
rect 1632 -11107 1666 -11073
rect 2460 -11014 2494 -10980
rect 2460 -11107 2494 -11073
rect 2920 -11014 2954 -10980
rect 2920 -11107 2954 -11073
rect 3748 -11014 3782 -10980
rect 3748 -11107 3782 -11073
rect 4208 -11014 4242 -10980
rect 4208 -11107 4242 -11073
rect 5036 -11014 5070 -10980
rect 5036 -11107 5070 -11073
rect 5496 -11014 5530 -10980
rect 5496 -11107 5530 -11073
rect 6324 -11014 6358 -10980
rect 6324 -11107 6358 -11073
rect 6784 -11014 6818 -10980
rect 6784 -11107 6818 -11073
rect 7612 -11014 7646 -10980
rect 7612 -11107 7646 -11073
rect 8072 -11014 8106 -10980
rect 8072 -11107 8106 -11073
rect 8900 -11014 8934 -10980
rect 8900 -11107 8934 -11073
rect 9360 -11014 9394 -10980
rect 9360 -11107 9394 -11073
rect 10188 -11014 10222 -10980
rect 10188 -11107 10222 -11073
rect 11476 -11014 11510 -10980
rect 11476 -11107 11510 -11073
rect 13500 -11014 13534 -10980
rect 13500 -11107 13534 -11073
rect 14696 -11014 14730 -10980
rect 14696 -11107 14730 -11073
rect 15892 -11014 15926 -10980
rect 15892 -11107 15926 -11073
rect -2232 -11799 -2198 -11765
rect -2232 -11892 -2198 -11858
rect -116 -11799 -82 -11765
rect -116 -11892 -82 -11858
rect 344 -11799 378 -11765
rect 344 -11892 378 -11858
rect 1172 -11799 1206 -11765
rect 1172 -11892 1206 -11858
rect 1632 -11799 1666 -11765
rect 1632 -11892 1666 -11858
rect 2460 -11799 2494 -11765
rect 2460 -11892 2494 -11858
rect 2920 -11799 2954 -11765
rect 2920 -11892 2954 -11858
rect 3748 -11799 3782 -11765
rect 3748 -11892 3782 -11858
rect 4208 -11799 4242 -11765
rect 4208 -11892 4242 -11858
rect 5036 -11799 5070 -11765
rect 5036 -11892 5070 -11858
rect 5496 -11799 5530 -11765
rect 5496 -11892 5530 -11858
rect 6324 -11799 6358 -11765
rect 6324 -11892 6358 -11858
rect 6784 -11799 6818 -11765
rect 6784 -11892 6818 -11858
rect 7612 -11799 7646 -11765
rect 7612 -11892 7646 -11858
rect 8072 -11799 8106 -11765
rect 8072 -11892 8106 -11858
rect 8900 -11799 8934 -11765
rect 8900 -11892 8934 -11858
rect 9360 -11799 9394 -11765
rect 9360 -11892 9394 -11858
rect 10188 -11799 10222 -11765
rect 10188 -11892 10222 -11858
rect 11476 -11799 11510 -11765
rect 11476 -11892 11510 -11858
rect 12396 -11799 12430 -11765
rect 12396 -11892 12430 -11858
rect 13132 -11799 13166 -11765
rect 13132 -11892 13166 -11858
rect 13592 -11799 13626 -11765
rect 13592 -11892 13626 -11858
rect 15524 -11799 15558 -11765
rect 15524 -11892 15558 -11858
rect -2232 -12102 -2198 -12068
rect -2232 -12195 -2198 -12161
rect -116 -12102 -82 -12068
rect -116 -12195 -82 -12161
rect 344 -12102 378 -12068
rect 344 -12195 378 -12161
rect 1172 -12102 1206 -12068
rect 1172 -12195 1206 -12161
rect 1632 -12102 1666 -12068
rect 1632 -12195 1666 -12161
rect 2460 -12102 2494 -12068
rect 2460 -12195 2494 -12161
rect 2920 -12102 2954 -12068
rect 2920 -12195 2954 -12161
rect 3748 -12102 3782 -12068
rect 3748 -12195 3782 -12161
rect 4208 -12102 4242 -12068
rect 4208 -12195 4242 -12161
rect 5036 -12102 5070 -12068
rect 5036 -12195 5070 -12161
rect 5496 -12102 5530 -12068
rect 5496 -12195 5530 -12161
rect 6324 -12102 6358 -12068
rect 6324 -12195 6358 -12161
rect 6784 -12102 6818 -12068
rect 6784 -12195 6818 -12161
rect 7612 -12102 7646 -12068
rect 7612 -12195 7646 -12161
rect 8072 -12102 8106 -12068
rect 8072 -12195 8106 -12161
rect 8900 -12102 8934 -12068
rect 8900 -12195 8934 -12161
rect 9360 -12102 9394 -12068
rect 9360 -12195 9394 -12161
rect 10188 -12102 10222 -12068
rect 10188 -12195 10222 -12161
rect 11476 -12102 11510 -12068
rect 11476 -12195 11510 -12161
rect 13592 -12102 13626 -12068
rect 13592 -12195 13626 -12161
rect 15524 -12102 15558 -12068
rect 15524 -12195 15558 -12161
rect -2232 -12887 -2198 -12853
rect -2232 -12980 -2198 -12946
rect -116 -12887 -82 -12853
rect -116 -12980 -82 -12946
rect 344 -12887 378 -12853
rect 344 -12980 378 -12946
rect 1172 -12887 1206 -12853
rect 1172 -12980 1206 -12946
rect 1632 -12887 1666 -12853
rect 1632 -12980 1666 -12946
rect 2460 -12887 2494 -12853
rect 2460 -12980 2494 -12946
rect 2920 -12887 2954 -12853
rect 2920 -12980 2954 -12946
rect 3748 -12887 3782 -12853
rect 3748 -12980 3782 -12946
rect 4208 -12887 4242 -12853
rect 4208 -12980 4242 -12946
rect 5036 -12887 5070 -12853
rect 5036 -12980 5070 -12946
rect 5496 -12887 5530 -12853
rect 5496 -12980 5530 -12946
rect 6324 -12887 6358 -12853
rect 6324 -12980 6358 -12946
rect 6784 -12887 6818 -12853
rect 6784 -12980 6818 -12946
rect 7612 -12887 7646 -12853
rect 7612 -12980 7646 -12946
rect 8072 -12887 8106 -12853
rect 8072 -12980 8106 -12946
rect 8900 -12887 8934 -12853
rect 8900 -12980 8934 -12946
rect 9360 -12887 9394 -12853
rect 9360 -12980 9394 -12946
rect 10188 -12887 10222 -12853
rect 10188 -12980 10222 -12946
rect 11476 -12887 11510 -12853
rect 11476 -12980 11510 -12946
rect 12396 -12887 12430 -12853
rect 12396 -12980 12430 -12946
rect 13132 -12887 13166 -12853
rect 13132 -12980 13166 -12946
rect 13592 -12887 13626 -12853
rect 13592 -12980 13626 -12946
rect 15524 -12887 15558 -12853
rect 15524 -12980 15558 -12946
rect -2232 -13190 -2198 -13156
rect -2232 -13283 -2198 -13249
rect -116 -13190 -82 -13156
rect -116 -13283 -82 -13249
rect 344 -13190 378 -13156
rect 344 -13283 378 -13249
rect 1172 -13190 1206 -13156
rect 1172 -13283 1206 -13249
rect 1632 -13190 1666 -13156
rect 1632 -13283 1666 -13249
rect 2460 -13190 2494 -13156
rect 2460 -13283 2494 -13249
rect 2920 -13190 2954 -13156
rect 2920 -13283 2954 -13249
rect 3748 -13190 3782 -13156
rect 3748 -13283 3782 -13249
rect 4208 -13190 4242 -13156
rect 4208 -13283 4242 -13249
rect 5036 -13190 5070 -13156
rect 5036 -13283 5070 -13249
rect 5496 -13190 5530 -13156
rect 5496 -13283 5530 -13249
rect 6324 -13190 6358 -13156
rect 6324 -13283 6358 -13249
rect 6784 -13190 6818 -13156
rect 6784 -13283 6818 -13249
rect 7612 -13190 7646 -13156
rect 7612 -13283 7646 -13249
rect 8072 -13190 8106 -13156
rect 8072 -13283 8106 -13249
rect 8900 -13190 8934 -13156
rect 8900 -13283 8934 -13249
rect 9360 -13190 9394 -13156
rect 9360 -13283 9394 -13249
rect 10188 -13190 10222 -13156
rect 10188 -13283 10222 -13249
rect 11476 -13190 11510 -13156
rect 11476 -13283 11510 -13249
rect 13592 -13190 13626 -13156
rect 13592 -13283 13626 -13249
rect 15524 -13190 15558 -13156
rect 15524 -13283 15558 -13249
rect -2232 -13975 -2198 -13941
rect -2232 -14068 -2198 -14034
rect -1036 -13975 -1002 -13941
rect -1036 -14068 -1002 -14034
rect -668 -13975 -634 -13941
rect -668 -14068 -634 -14034
rect -208 -13975 -174 -13941
rect -208 -14068 -174 -14034
rect 528 -13975 562 -13941
rect 528 -14068 562 -14034
rect 988 -13975 1022 -13941
rect 988 -14068 1022 -14034
rect 1356 -13975 1390 -13941
rect 1356 -14068 1390 -14034
rect 1816 -13975 1850 -13941
rect 1816 -14068 1850 -14034
rect 2276 -13975 2310 -13941
rect 2276 -14068 2310 -14034
rect 3104 -13975 3138 -13941
rect 3104 -14068 3138 -14034
rect 3564 -13975 3598 -13941
rect 3564 -14068 3598 -14034
rect 6324 -13975 6358 -13941
rect 6324 -14068 6358 -14034
rect 6784 -13975 6818 -13941
rect 6784 -14068 6818 -14034
rect 7612 -13975 7646 -13941
rect 7612 -14068 7646 -14034
rect 8072 -13975 8106 -13941
rect 8072 -14068 8106 -14034
rect 8900 -13975 8934 -13941
rect 8900 -14068 8934 -14034
rect 9360 -13975 9394 -13941
rect 9360 -14068 9394 -14034
rect 10188 -13975 10222 -13941
rect 10188 -14068 10222 -14034
rect 10648 -13975 10682 -13941
rect 10648 -14068 10682 -14034
rect 11568 -13975 11602 -13941
rect 11568 -14068 11602 -14034
rect 13500 -13975 13534 -13941
rect 13500 -14068 13534 -14034
rect 14696 -13975 14730 -13941
rect 14696 -14068 14730 -14034
rect 15892 -13975 15926 -13941
rect 15892 -14068 15926 -14034
<< poly >>
rect -2918 -59 -2340 -33
rect -1354 -59 -1144 -33
rect -890 -59 -860 -33
rect -806 -59 -776 -33
rect -526 -59 -316 -33
rect -57 -59 -27 -33
rect 29 -59 59 -33
rect 115 -59 145 -33
rect 201 -59 231 -33
rect 287 -59 317 -33
rect 373 -59 403 -33
rect 670 -59 880 -33
rect 1130 -59 1160 -33
rect 1214 -59 1244 -33
rect 1498 -59 1708 -33
rect 1958 -59 2168 -33
rect 2420 -59 2450 -33
rect 2522 -59 2622 -33
rect 2782 -59 2882 -33
rect 2947 -59 2977 -33
rect 3246 -59 3456 -33
rect 4442 -59 5388 -33
rect 6466 -59 6676 -33
rect 6928 -59 6958 -33
rect 7030 -59 7130 -33
rect 7290 -59 7390 -33
rect 7455 -59 7485 -33
rect 7754 -59 7964 -33
rect 8216 -59 8246 -33
rect 8318 -59 8418 -33
rect 8578 -59 8678 -33
rect 8743 -59 8773 -33
rect 9042 -59 9252 -33
rect 9504 -59 9534 -33
rect 9606 -59 9706 -33
rect 9866 -59 9966 -33
rect 10031 -59 10061 -33
rect 10330 -59 10540 -33
rect 10790 -59 10820 -33
rect 10874 -59 10904 -33
rect 10958 -59 10988 -33
rect 11042 -59 11072 -33
rect 11126 -59 11156 -33
rect 11210 -59 11240 -33
rect 11294 -59 11324 -33
rect 11378 -59 11408 -33
rect 11710 -59 11920 -33
rect 13642 -59 14588 -33
rect 14838 -59 15784 -33
rect 16034 -59 16612 -33
rect -2918 -259 -2340 -233
rect -1354 -259 -1144 -233
rect -526 -259 -316 -233
rect 670 -259 880 -233
rect -2918 -281 -2654 -259
rect -1354 -265 -1270 -259
rect -2918 -315 -2902 -281
rect -2868 -315 -2803 -281
rect -2769 -315 -2704 -281
rect -2670 -315 -2654 -281
rect -1412 -281 -1270 -265
rect -2918 -331 -2654 -315
rect -2612 -317 -2340 -301
rect -2612 -351 -2596 -317
rect -2562 -351 -2493 -317
rect -2459 -351 -2390 -317
rect -2356 -351 -2340 -317
rect -1412 -315 -1396 -281
rect -1362 -315 -1270 -281
rect -890 -291 -860 -259
rect -1412 -331 -1270 -315
rect -1228 -317 -1086 -301
rect -2612 -373 -2340 -351
rect -1228 -351 -1136 -317
rect -1102 -351 -1086 -317
rect -1228 -367 -1086 -351
rect -952 -307 -860 -291
rect -952 -341 -937 -307
rect -903 -341 -860 -307
rect -952 -357 -860 -341
rect -1228 -373 -1144 -367
rect -2918 -399 -2340 -373
rect -1354 -399 -1144 -373
rect -890 -379 -860 -357
rect -806 -291 -776 -259
rect -526 -265 -442 -259
rect -584 -281 -442 -265
rect -806 -307 -718 -291
rect -806 -341 -769 -307
rect -735 -341 -718 -307
rect -584 -315 -568 -281
rect -534 -315 -442 -281
rect -57 -297 -27 -259
rect 29 -297 59 -259
rect 115 -297 145 -259
rect 201 -297 231 -259
rect 287 -297 317 -259
rect 373 -297 403 -259
rect 670 -265 754 -259
rect -584 -331 -442 -315
rect -400 -317 -258 -301
rect -806 -357 -718 -341
rect -400 -351 -308 -317
rect -274 -351 -258 -317
rect -57 -307 403 -297
rect -57 -341 -30 -307
rect 4 -341 38 -307
rect 72 -341 106 -307
rect 140 -341 174 -307
rect 208 -341 242 -307
rect 276 -341 310 -307
rect 344 -341 403 -307
rect 612 -281 754 -265
rect 612 -315 628 -281
rect 662 -315 754 -281
rect 1130 -287 1160 -227
rect 1214 -287 1244 -227
rect 1498 -259 1708 -233
rect 1958 -259 2168 -233
rect 1498 -265 1582 -259
rect 1958 -265 2042 -259
rect 1130 -291 1244 -287
rect 612 -331 754 -315
rect 796 -317 938 -301
rect -57 -351 403 -341
rect 796 -351 888 -317
rect 922 -351 938 -317
rect -806 -379 -776 -357
rect -400 -367 -258 -351
rect -400 -373 -316 -367
rect -526 -399 -316 -373
rect 29 -425 59 -351
rect 115 -425 145 -351
rect 201 -425 231 -351
rect 287 -425 317 -351
rect 796 -367 938 -351
rect 1072 -307 1244 -291
rect 1072 -341 1082 -307
rect 1116 -317 1244 -307
rect 1440 -281 1582 -265
rect 1440 -315 1456 -281
rect 1490 -315 1582 -281
rect 1900 -281 2042 -265
rect 1116 -341 1243 -317
rect 1440 -331 1582 -315
rect 1624 -317 1766 -301
rect 1072 -357 1243 -341
rect 1129 -361 1243 -357
rect 796 -373 880 -367
rect 670 -399 880 -373
rect 1213 -425 1243 -361
rect 1624 -351 1716 -317
rect 1750 -351 1766 -317
rect 1900 -315 1916 -281
rect 1950 -315 2042 -281
rect 2420 -294 2450 -259
rect 1900 -331 2042 -315
rect 2084 -317 2226 -301
rect 1624 -367 1766 -351
rect 2084 -351 2176 -317
rect 2210 -351 2226 -317
rect 2084 -367 2226 -351
rect 2380 -307 2450 -294
rect 2522 -297 2622 -223
rect 2782 -297 2882 -223
rect 3246 -259 3456 -233
rect 4442 -259 5388 -233
rect 6466 -259 6676 -233
rect 2947 -291 2977 -259
rect 3246 -265 3330 -259
rect 3188 -281 3330 -265
rect 2380 -341 2396 -307
rect 2430 -341 2450 -307
rect 2380 -353 2450 -341
rect 2500 -307 2622 -297
rect 2500 -341 2516 -307
rect 2550 -341 2622 -307
rect 2500 -351 2622 -341
rect 2721 -307 2882 -297
rect 2721 -341 2737 -307
rect 2771 -341 2882 -307
rect 2721 -351 2882 -341
rect 1624 -373 1708 -367
rect 2084 -373 2168 -367
rect 1498 -399 1708 -373
rect 1958 -399 2168 -373
rect 2420 -425 2450 -353
rect 2522 -379 2622 -351
rect 2782 -379 2882 -351
rect 2927 -307 2981 -291
rect 2927 -341 2937 -307
rect 2971 -341 2981 -307
rect 3188 -315 3204 -281
rect 3238 -315 3330 -281
rect 4442 -281 4892 -259
rect 6466 -265 6550 -259
rect 3188 -331 3330 -315
rect 3372 -317 3514 -301
rect 2927 -357 2981 -341
rect 3372 -351 3464 -317
rect 3498 -351 3514 -317
rect 4442 -315 4458 -281
rect 4492 -315 4586 -281
rect 4620 -315 4714 -281
rect 4748 -315 4842 -281
rect 4876 -315 4892 -281
rect 6408 -281 6550 -265
rect 4442 -331 4892 -315
rect 4934 -317 5388 -301
rect 2947 -425 2977 -357
rect 3372 -367 3514 -351
rect 4934 -351 4950 -317
rect 4984 -351 5078 -317
rect 5112 -351 5206 -317
rect 5240 -351 5334 -317
rect 5368 -351 5388 -317
rect 6408 -315 6424 -281
rect 6458 -315 6550 -281
rect 6928 -294 6958 -259
rect 6408 -331 6550 -315
rect 6592 -317 6734 -301
rect 3372 -373 3456 -367
rect 4934 -373 5388 -351
rect 6592 -351 6684 -317
rect 6718 -351 6734 -317
rect 6592 -367 6734 -351
rect 6888 -307 6958 -294
rect 7030 -297 7130 -223
rect 7290 -297 7390 -223
rect 7754 -259 7964 -233
rect 7455 -291 7485 -259
rect 7754 -265 7838 -259
rect 7696 -281 7838 -265
rect 6888 -341 6904 -307
rect 6938 -341 6958 -307
rect 6888 -353 6958 -341
rect 7008 -307 7130 -297
rect 7008 -341 7024 -307
rect 7058 -341 7130 -307
rect 7008 -351 7130 -341
rect 7229 -307 7390 -297
rect 7229 -341 7245 -307
rect 7279 -341 7390 -307
rect 7229 -351 7390 -341
rect 6592 -373 6676 -367
rect 3246 -399 3456 -373
rect 4442 -399 5388 -373
rect 6466 -399 6676 -373
rect 6928 -425 6958 -353
rect 7030 -379 7130 -351
rect 7290 -379 7390 -351
rect 7435 -307 7489 -291
rect 7435 -341 7445 -307
rect 7479 -341 7489 -307
rect 7696 -315 7712 -281
rect 7746 -315 7838 -281
rect 8216 -294 8246 -259
rect 7696 -331 7838 -315
rect 7880 -317 8022 -301
rect 7435 -357 7489 -341
rect 7880 -351 7972 -317
rect 8006 -351 8022 -317
rect 7455 -425 7485 -357
rect 7880 -367 8022 -351
rect 8176 -307 8246 -294
rect 8318 -297 8418 -223
rect 8578 -297 8678 -223
rect 9042 -259 9252 -233
rect 8743 -291 8773 -259
rect 9042 -265 9126 -259
rect 8984 -281 9126 -265
rect 8176 -341 8192 -307
rect 8226 -341 8246 -307
rect 8176 -353 8246 -341
rect 8296 -307 8418 -297
rect 8296 -341 8312 -307
rect 8346 -341 8418 -307
rect 8296 -351 8418 -341
rect 8517 -307 8678 -297
rect 8517 -341 8533 -307
rect 8567 -341 8678 -307
rect 8517 -351 8678 -341
rect 7880 -373 7964 -367
rect 7754 -399 7964 -373
rect 8216 -425 8246 -353
rect 8318 -379 8418 -351
rect 8578 -379 8678 -351
rect 8723 -307 8777 -291
rect 8723 -341 8733 -307
rect 8767 -341 8777 -307
rect 8984 -315 9000 -281
rect 9034 -315 9126 -281
rect 9504 -294 9534 -259
rect 8984 -331 9126 -315
rect 9168 -317 9310 -301
rect 8723 -357 8777 -341
rect 9168 -351 9260 -317
rect 9294 -351 9310 -317
rect 8743 -425 8773 -357
rect 9168 -367 9310 -351
rect 9464 -307 9534 -294
rect 9606 -297 9706 -223
rect 9866 -297 9966 -223
rect 10330 -259 10540 -233
rect 11710 -259 11920 -233
rect 13642 -259 14588 -233
rect 14838 -259 15784 -233
rect 16034 -259 16612 -233
rect 10031 -291 10061 -259
rect 10330 -265 10414 -259
rect 10272 -281 10414 -265
rect 9464 -341 9480 -307
rect 9514 -341 9534 -307
rect 9464 -353 9534 -341
rect 9584 -307 9706 -297
rect 9584 -341 9600 -307
rect 9634 -341 9706 -307
rect 9584 -351 9706 -341
rect 9805 -307 9966 -297
rect 9805 -341 9821 -307
rect 9855 -341 9966 -307
rect 9805 -351 9966 -341
rect 9168 -373 9252 -367
rect 9042 -399 9252 -373
rect 9504 -425 9534 -353
rect 9606 -379 9706 -351
rect 9866 -379 9966 -351
rect 10011 -307 10065 -291
rect 10011 -341 10021 -307
rect 10055 -341 10065 -307
rect 10272 -315 10288 -281
rect 10322 -315 10414 -281
rect 10790 -291 10820 -259
rect 10874 -291 10904 -259
rect 10958 -291 10988 -259
rect 11042 -291 11072 -259
rect 10272 -331 10414 -315
rect 10456 -317 10598 -301
rect 10011 -357 10065 -341
rect 10456 -351 10548 -317
rect 10582 -351 10598 -317
rect 10031 -425 10061 -357
rect 10456 -367 10598 -351
rect 10733 -307 11072 -291
rect 10733 -341 10749 -307
rect 10783 -341 10830 -307
rect 10864 -341 10914 -307
rect 10948 -341 10998 -307
rect 11032 -341 11072 -307
rect 10733 -357 11072 -341
rect 10456 -373 10540 -367
rect 10330 -399 10540 -373
rect 10790 -379 10820 -357
rect 10874 -379 10904 -357
rect 10958 -379 10988 -357
rect 11042 -379 11072 -357
rect 11126 -291 11156 -259
rect 11210 -291 11240 -259
rect 11294 -291 11324 -259
rect 11378 -291 11408 -259
rect 11710 -265 11794 -259
rect 11126 -307 11408 -291
rect 11126 -341 11250 -307
rect 11284 -341 11334 -307
rect 11368 -341 11408 -307
rect 11652 -281 11794 -265
rect 11652 -315 11668 -281
rect 11702 -315 11794 -281
rect 13642 -281 14092 -259
rect 11652 -331 11794 -315
rect 11836 -317 11978 -301
rect 11126 -357 11408 -341
rect 11126 -379 11156 -357
rect 11210 -379 11240 -357
rect 11294 -379 11324 -357
rect 11378 -379 11408 -357
rect 11836 -351 11928 -317
rect 11962 -351 11978 -317
rect 13642 -315 13658 -281
rect 13692 -315 13786 -281
rect 13820 -315 13914 -281
rect 13948 -315 14042 -281
rect 14076 -315 14092 -281
rect 14838 -281 15288 -259
rect 13642 -331 14092 -315
rect 14134 -317 14588 -301
rect 11836 -367 11978 -351
rect 14134 -351 14150 -317
rect 14184 -351 14278 -317
rect 14312 -351 14406 -317
rect 14440 -351 14534 -317
rect 14568 -351 14588 -317
rect 14838 -315 14854 -281
rect 14888 -315 14982 -281
rect 15016 -315 15110 -281
rect 15144 -315 15238 -281
rect 15272 -315 15288 -281
rect 16034 -281 16298 -259
rect 14838 -331 15288 -315
rect 15330 -317 15784 -301
rect 11836 -373 11920 -367
rect 14134 -373 14588 -351
rect 15330 -351 15346 -317
rect 15380 -351 15474 -317
rect 15508 -351 15602 -317
rect 15636 -351 15730 -317
rect 15764 -351 15784 -317
rect 16034 -315 16050 -281
rect 16084 -315 16149 -281
rect 16183 -315 16248 -281
rect 16282 -315 16298 -281
rect 16034 -331 16298 -315
rect 16340 -317 16612 -301
rect 15330 -373 15784 -351
rect 16340 -351 16356 -317
rect 16390 -351 16459 -317
rect 16493 -351 16562 -317
rect 16596 -351 16612 -317
rect 16340 -373 16612 -351
rect 11710 -399 11920 -373
rect 13642 -399 14588 -373
rect 14838 -399 15784 -373
rect 16034 -399 16612 -373
rect -2918 -535 -2340 -509
rect -1354 -535 -1144 -509
rect -890 -535 -860 -509
rect -806 -535 -776 -509
rect -526 -535 -316 -509
rect 29 -535 59 -509
rect 115 -535 145 -509
rect 201 -535 231 -509
rect 287 -535 317 -509
rect 670 -535 880 -509
rect 1213 -535 1243 -509
rect 1498 -535 1708 -509
rect 1958 -535 2168 -509
rect 2420 -535 2450 -509
rect 2522 -535 2622 -509
rect 2782 -535 2882 -509
rect 2947 -535 2977 -509
rect 3246 -535 3456 -509
rect 4442 -535 5388 -509
rect 6466 -535 6676 -509
rect 6928 -535 6958 -509
rect 7030 -535 7130 -509
rect 7290 -535 7390 -509
rect 7455 -535 7485 -509
rect 7754 -535 7964 -509
rect 8216 -535 8246 -509
rect 8318 -535 8418 -509
rect 8578 -535 8678 -509
rect 8743 -535 8773 -509
rect 9042 -535 9252 -509
rect 9504 -535 9534 -509
rect 9606 -535 9706 -509
rect 9866 -535 9966 -509
rect 10031 -535 10061 -509
rect 10330 -535 10540 -509
rect 10790 -535 10820 -509
rect 10874 -535 10904 -509
rect 10958 -535 10988 -509
rect 11042 -535 11072 -509
rect 11126 -535 11156 -509
rect 11210 -535 11240 -509
rect 11294 -535 11324 -509
rect 11378 -535 11408 -509
rect 11710 -535 11920 -509
rect 13642 -535 14588 -509
rect 14838 -535 15784 -509
rect 16034 -535 16612 -509
rect -2918 -603 -2340 -577
rect -1538 -603 -960 -577
rect -802 -603 -224 -577
rect 26 -603 236 -577
rect 505 -603 535 -577
rect 600 -603 700 -577
rect 860 -603 960 -577
rect 1032 -603 1062 -577
rect 1314 -603 1524 -577
rect 1774 -603 2352 -577
rect 2602 -603 2812 -577
rect 3081 -603 3111 -577
rect 3176 -603 3276 -577
rect 3436 -603 3536 -577
rect 3608 -603 3638 -577
rect 3890 -603 4100 -577
rect 4350 -603 4928 -577
rect 5178 -603 5388 -577
rect 5657 -603 5687 -577
rect 5752 -603 5852 -577
rect 6012 -603 6112 -577
rect 6184 -603 6214 -577
rect 6466 -603 6676 -577
rect 6926 -603 7504 -577
rect 7754 -603 7964 -577
rect 8233 -603 8263 -577
rect 8328 -603 8428 -577
rect 8588 -603 8688 -577
rect 8760 -603 8790 -577
rect 9042 -603 9252 -577
rect 9502 -603 10080 -577
rect 10422 -603 10632 -577
rect 10809 -603 10839 -577
rect 10904 -603 11004 -577
rect 11164 -603 11264 -577
rect 11336 -603 11366 -577
rect 11710 -603 11920 -577
rect 13735 -603 13765 -577
rect 13821 -603 13851 -577
rect 13907 -603 13937 -577
rect 13993 -603 14023 -577
rect 14079 -603 14109 -577
rect 14165 -603 14195 -577
rect 14251 -603 14281 -577
rect 14337 -603 14367 -577
rect 14423 -603 14453 -577
rect 14509 -603 14539 -577
rect 14595 -603 14625 -577
rect 14681 -603 14711 -577
rect 14766 -603 14796 -577
rect 14852 -603 14882 -577
rect 14938 -603 14968 -577
rect 15024 -603 15054 -577
rect 15110 -603 15140 -577
rect 15196 -603 15226 -577
rect 15282 -603 15312 -577
rect 15368 -603 15398 -577
rect 15666 -603 16612 -577
rect -2918 -739 -2340 -713
rect -1538 -739 -960 -713
rect -802 -739 -224 -713
rect 26 -739 236 -713
rect -2918 -761 -2646 -739
rect -2918 -795 -2902 -761
rect -2868 -795 -2799 -761
rect -2765 -795 -2696 -761
rect -2662 -795 -2646 -761
rect -1538 -761 -1266 -739
rect -2918 -811 -2646 -795
rect -2604 -797 -2340 -781
rect -2604 -831 -2588 -797
rect -2554 -831 -2489 -797
rect -2455 -831 -2390 -797
rect -2356 -831 -2340 -797
rect -1538 -795 -1522 -761
rect -1488 -795 -1419 -761
rect -1385 -795 -1316 -761
rect -1282 -795 -1266 -761
rect -802 -761 -530 -739
rect 26 -745 110 -739
rect -1538 -811 -1266 -795
rect -1224 -797 -960 -781
rect -2604 -853 -2340 -831
rect -1224 -831 -1208 -797
rect -1174 -831 -1109 -797
rect -1075 -831 -1010 -797
rect -976 -831 -960 -797
rect -802 -795 -786 -761
rect -752 -795 -683 -761
rect -649 -795 -580 -761
rect -546 -795 -530 -761
rect -32 -761 110 -745
rect 505 -755 535 -687
rect -802 -811 -530 -795
rect -488 -797 -224 -781
rect -1224 -853 -960 -831
rect -488 -831 -472 -797
rect -438 -831 -373 -797
rect -339 -831 -274 -797
rect -240 -831 -224 -797
rect -32 -795 -16 -761
rect 18 -795 110 -761
rect 501 -771 555 -755
rect -32 -811 110 -795
rect 152 -797 294 -781
rect -488 -853 -224 -831
rect 152 -831 244 -797
rect 278 -831 294 -797
rect 501 -805 511 -771
rect 545 -805 555 -771
rect 501 -821 555 -805
rect 600 -761 700 -733
rect 860 -761 960 -733
rect 1032 -759 1062 -687
rect 1314 -739 1524 -713
rect 1774 -739 2352 -713
rect 2602 -739 2812 -713
rect 1314 -745 1398 -739
rect 600 -771 761 -761
rect 600 -805 711 -771
rect 745 -805 761 -771
rect 600 -815 761 -805
rect 860 -771 982 -761
rect 860 -805 932 -771
rect 966 -805 982 -771
rect 860 -815 982 -805
rect 1032 -771 1102 -759
rect 1032 -805 1052 -771
rect 1086 -805 1102 -771
rect 152 -847 294 -831
rect 152 -853 236 -847
rect 505 -853 535 -821
rect -2918 -879 -2340 -853
rect -1538 -879 -960 -853
rect -802 -879 -224 -853
rect 26 -879 236 -853
rect 600 -889 700 -815
rect 860 -889 960 -815
rect 1032 -818 1102 -805
rect 1256 -761 1398 -745
rect 1256 -795 1272 -761
rect 1306 -795 1398 -761
rect 1774 -761 2046 -739
rect 2602 -745 2686 -739
rect 1256 -811 1398 -795
rect 1440 -797 1582 -781
rect 1032 -853 1062 -818
rect 1440 -831 1532 -797
rect 1566 -831 1582 -797
rect 1774 -795 1790 -761
rect 1824 -795 1893 -761
rect 1927 -795 1996 -761
rect 2030 -795 2046 -761
rect 2544 -761 2686 -745
rect 3081 -755 3111 -687
rect 1774 -811 2046 -795
rect 2088 -797 2352 -781
rect 1440 -847 1582 -831
rect 2088 -831 2104 -797
rect 2138 -831 2203 -797
rect 2237 -831 2302 -797
rect 2336 -831 2352 -797
rect 2544 -795 2560 -761
rect 2594 -795 2686 -761
rect 3077 -771 3131 -755
rect 2544 -811 2686 -795
rect 2728 -797 2870 -781
rect 1440 -853 1524 -847
rect 2088 -853 2352 -831
rect 2728 -831 2820 -797
rect 2854 -831 2870 -797
rect 3077 -805 3087 -771
rect 3121 -805 3131 -771
rect 3077 -821 3131 -805
rect 3176 -761 3276 -733
rect 3436 -761 3536 -733
rect 3608 -759 3638 -687
rect 3890 -739 4100 -713
rect 4350 -739 4928 -713
rect 5178 -739 5388 -713
rect 3890 -745 3974 -739
rect 3176 -771 3337 -761
rect 3176 -805 3287 -771
rect 3321 -805 3337 -771
rect 3176 -815 3337 -805
rect 3436 -771 3558 -761
rect 3436 -805 3508 -771
rect 3542 -805 3558 -771
rect 3436 -815 3558 -805
rect 3608 -771 3678 -759
rect 3608 -805 3628 -771
rect 3662 -805 3678 -771
rect 2728 -847 2870 -831
rect 2728 -853 2812 -847
rect 3081 -853 3111 -821
rect 1314 -879 1524 -853
rect 1774 -879 2352 -853
rect 2602 -879 2812 -853
rect 3176 -889 3276 -815
rect 3436 -889 3536 -815
rect 3608 -818 3678 -805
rect 3832 -761 3974 -745
rect 3832 -795 3848 -761
rect 3882 -795 3974 -761
rect 4350 -761 4622 -739
rect 5178 -745 5262 -739
rect 3832 -811 3974 -795
rect 4016 -797 4158 -781
rect 3608 -853 3638 -818
rect 4016 -831 4108 -797
rect 4142 -831 4158 -797
rect 4350 -795 4366 -761
rect 4400 -795 4469 -761
rect 4503 -795 4572 -761
rect 4606 -795 4622 -761
rect 5120 -761 5262 -745
rect 5657 -755 5687 -687
rect 4350 -811 4622 -795
rect 4664 -797 4928 -781
rect 4016 -847 4158 -831
rect 4664 -831 4680 -797
rect 4714 -831 4779 -797
rect 4813 -831 4878 -797
rect 4912 -831 4928 -797
rect 5120 -795 5136 -761
rect 5170 -795 5262 -761
rect 5653 -771 5707 -755
rect 5120 -811 5262 -795
rect 5304 -797 5446 -781
rect 4016 -853 4100 -847
rect 4664 -853 4928 -831
rect 5304 -831 5396 -797
rect 5430 -831 5446 -797
rect 5653 -805 5663 -771
rect 5697 -805 5707 -771
rect 5653 -821 5707 -805
rect 5752 -761 5852 -733
rect 6012 -761 6112 -733
rect 6184 -759 6214 -687
rect 6466 -739 6676 -713
rect 6926 -739 7504 -713
rect 7754 -739 7964 -713
rect 6466 -745 6550 -739
rect 5752 -771 5913 -761
rect 5752 -805 5863 -771
rect 5897 -805 5913 -771
rect 5752 -815 5913 -805
rect 6012 -771 6134 -761
rect 6012 -805 6084 -771
rect 6118 -805 6134 -771
rect 6012 -815 6134 -805
rect 6184 -771 6254 -759
rect 6184 -805 6204 -771
rect 6238 -805 6254 -771
rect 5304 -847 5446 -831
rect 5304 -853 5388 -847
rect 5657 -853 5687 -821
rect 3890 -879 4100 -853
rect 4350 -879 4928 -853
rect 5178 -879 5388 -853
rect 5752 -889 5852 -815
rect 6012 -889 6112 -815
rect 6184 -818 6254 -805
rect 6408 -761 6550 -745
rect 6408 -795 6424 -761
rect 6458 -795 6550 -761
rect 6926 -761 7198 -739
rect 7754 -745 7838 -739
rect 6408 -811 6550 -795
rect 6592 -797 6734 -781
rect 6184 -853 6214 -818
rect 6592 -831 6684 -797
rect 6718 -831 6734 -797
rect 6926 -795 6942 -761
rect 6976 -795 7045 -761
rect 7079 -795 7148 -761
rect 7182 -795 7198 -761
rect 7696 -761 7838 -745
rect 8233 -755 8263 -687
rect 6926 -811 7198 -795
rect 7240 -797 7504 -781
rect 6592 -847 6734 -831
rect 7240 -831 7256 -797
rect 7290 -831 7355 -797
rect 7389 -831 7454 -797
rect 7488 -831 7504 -797
rect 7696 -795 7712 -761
rect 7746 -795 7838 -761
rect 8229 -771 8283 -755
rect 7696 -811 7838 -795
rect 7880 -797 8022 -781
rect 6592 -853 6676 -847
rect 7240 -853 7504 -831
rect 7880 -831 7972 -797
rect 8006 -831 8022 -797
rect 8229 -805 8239 -771
rect 8273 -805 8283 -771
rect 8229 -821 8283 -805
rect 8328 -761 8428 -733
rect 8588 -761 8688 -733
rect 8760 -759 8790 -687
rect 9042 -739 9252 -713
rect 9502 -739 10080 -713
rect 10422 -739 10632 -713
rect 9042 -745 9126 -739
rect 8328 -771 8489 -761
rect 8328 -805 8439 -771
rect 8473 -805 8489 -771
rect 8328 -815 8489 -805
rect 8588 -771 8710 -761
rect 8588 -805 8660 -771
rect 8694 -805 8710 -771
rect 8588 -815 8710 -805
rect 8760 -771 8830 -759
rect 8760 -805 8780 -771
rect 8814 -805 8830 -771
rect 7880 -847 8022 -831
rect 7880 -853 7964 -847
rect 8233 -853 8263 -821
rect 6466 -879 6676 -853
rect 6926 -879 7504 -853
rect 7754 -879 7964 -853
rect 8328 -889 8428 -815
rect 8588 -889 8688 -815
rect 8760 -818 8830 -805
rect 8984 -761 9126 -745
rect 8984 -795 9000 -761
rect 9034 -795 9126 -761
rect 9502 -761 9774 -739
rect 10422 -745 10506 -739
rect 8984 -811 9126 -795
rect 9168 -797 9310 -781
rect 8760 -853 8790 -818
rect 9168 -831 9260 -797
rect 9294 -831 9310 -797
rect 9502 -795 9518 -761
rect 9552 -795 9621 -761
rect 9655 -795 9724 -761
rect 9758 -795 9774 -761
rect 10364 -761 10506 -745
rect 10809 -755 10839 -687
rect 9502 -811 9774 -795
rect 9816 -797 10080 -781
rect 9168 -847 9310 -831
rect 9816 -831 9832 -797
rect 9866 -831 9931 -797
rect 9965 -831 10030 -797
rect 10064 -831 10080 -797
rect 10364 -795 10380 -761
rect 10414 -795 10506 -761
rect 10805 -771 10859 -755
rect 10364 -811 10506 -795
rect 10548 -797 10690 -781
rect 9168 -853 9252 -847
rect 9816 -853 10080 -831
rect 10548 -831 10640 -797
rect 10674 -831 10690 -797
rect 10805 -805 10815 -771
rect 10849 -805 10859 -771
rect 10805 -821 10859 -805
rect 10904 -761 11004 -733
rect 11164 -761 11264 -733
rect 11336 -759 11366 -687
rect 11710 -739 11920 -713
rect 13735 -736 13765 -687
rect 13821 -736 13851 -687
rect 13907 -736 13937 -687
rect 13993 -736 14023 -687
rect 11710 -745 11794 -739
rect 10904 -771 11065 -761
rect 10904 -805 11015 -771
rect 11049 -805 11065 -771
rect 10904 -815 11065 -805
rect 11164 -771 11286 -761
rect 11164 -805 11236 -771
rect 11270 -805 11286 -771
rect 11164 -815 11286 -805
rect 11336 -771 11406 -759
rect 11336 -805 11356 -771
rect 11390 -805 11406 -771
rect 10548 -847 10690 -831
rect 10548 -853 10632 -847
rect 10809 -853 10839 -821
rect 9042 -879 9252 -853
rect 9502 -879 10080 -853
rect 10422 -879 10632 -853
rect 10904 -889 11004 -815
rect 11164 -889 11264 -815
rect 11336 -818 11406 -805
rect 11652 -761 11794 -745
rect 11652 -795 11668 -761
rect 11702 -795 11794 -761
rect 13676 -771 14023 -736
rect 11652 -811 11794 -795
rect 11836 -797 11978 -781
rect 11336 -853 11366 -818
rect 11836 -831 11928 -797
rect 11962 -831 11978 -797
rect 11836 -847 11978 -831
rect 13676 -805 13692 -771
rect 13726 -805 14023 -771
rect 13676 -838 14023 -805
rect 11836 -853 11920 -847
rect 13735 -853 13765 -838
rect 13821 -853 13851 -838
rect 13907 -853 13937 -838
rect 13993 -853 14023 -838
rect 14079 -746 14109 -687
rect 14165 -746 14195 -687
rect 14251 -746 14281 -687
rect 14337 -746 14367 -687
rect 14423 -746 14453 -687
rect 14509 -746 14539 -687
rect 14595 -746 14625 -687
rect 14681 -746 14711 -687
rect 14766 -746 14796 -687
rect 14852 -746 14882 -687
rect 14938 -746 14968 -687
rect 15024 -746 15054 -687
rect 15110 -746 15140 -687
rect 15196 -746 15226 -687
rect 15282 -746 15312 -687
rect 15368 -746 15398 -687
rect 14079 -771 15398 -746
rect 14079 -805 14119 -771
rect 14153 -805 14187 -771
rect 14221 -805 14255 -771
rect 14289 -805 14323 -771
rect 14357 -805 14391 -771
rect 14425 -805 14459 -771
rect 14493 -805 14527 -771
rect 14561 -805 14595 -771
rect 14629 -805 14663 -771
rect 14697 -805 14731 -771
rect 14765 -805 14799 -771
rect 14833 -805 14867 -771
rect 14901 -805 14935 -771
rect 14969 -805 15003 -771
rect 15037 -805 15071 -771
rect 15105 -805 15139 -771
rect 15173 -805 15398 -771
rect 14079 -821 15398 -805
rect 15666 -739 16612 -713
rect 15666 -761 16120 -739
rect 15666 -795 15686 -761
rect 15720 -795 15814 -761
rect 15848 -795 15942 -761
rect 15976 -795 16070 -761
rect 16104 -795 16120 -761
rect 15666 -811 16120 -795
rect 16162 -797 16612 -781
rect 14079 -853 14109 -821
rect 14165 -853 14195 -821
rect 14251 -853 14281 -821
rect 14337 -853 14367 -821
rect 14423 -853 14453 -821
rect 14509 -853 14539 -821
rect 14595 -853 14625 -821
rect 14681 -853 14711 -821
rect 14766 -853 14796 -821
rect 14852 -853 14882 -821
rect 14938 -853 14968 -821
rect 15024 -853 15054 -821
rect 15110 -853 15140 -821
rect 15196 -853 15226 -821
rect 15282 -853 15312 -821
rect 15368 -853 15398 -821
rect 16162 -831 16178 -797
rect 16212 -831 16306 -797
rect 16340 -831 16434 -797
rect 16468 -831 16562 -797
rect 16596 -831 16612 -797
rect 16162 -853 16612 -831
rect 11710 -879 11920 -853
rect 15666 -879 16612 -853
rect -2918 -1079 -2340 -1053
rect -1538 -1079 -960 -1053
rect -802 -1079 -224 -1053
rect 26 -1079 236 -1053
rect 505 -1079 535 -1053
rect 600 -1079 700 -1053
rect 860 -1079 960 -1053
rect 1032 -1079 1062 -1053
rect 1314 -1079 1524 -1053
rect 1774 -1079 2352 -1053
rect 2602 -1079 2812 -1053
rect 3081 -1079 3111 -1053
rect 3176 -1079 3276 -1053
rect 3436 -1079 3536 -1053
rect 3608 -1079 3638 -1053
rect 3890 -1079 4100 -1053
rect 4350 -1079 4928 -1053
rect 5178 -1079 5388 -1053
rect 5657 -1079 5687 -1053
rect 5752 -1079 5852 -1053
rect 6012 -1079 6112 -1053
rect 6184 -1079 6214 -1053
rect 6466 -1079 6676 -1053
rect 6926 -1079 7504 -1053
rect 7754 -1079 7964 -1053
rect 8233 -1079 8263 -1053
rect 8328 -1079 8428 -1053
rect 8588 -1079 8688 -1053
rect 8760 -1079 8790 -1053
rect 9042 -1079 9252 -1053
rect 9502 -1079 10080 -1053
rect 10422 -1079 10632 -1053
rect 10809 -1079 10839 -1053
rect 10904 -1079 11004 -1053
rect 11164 -1079 11264 -1053
rect 11336 -1079 11366 -1053
rect 11710 -1079 11920 -1053
rect 13735 -1079 13765 -1053
rect 13821 -1079 13851 -1053
rect 13907 -1079 13937 -1053
rect 13993 -1079 14023 -1053
rect 14079 -1079 14109 -1053
rect 14165 -1079 14195 -1053
rect 14251 -1079 14281 -1053
rect 14337 -1079 14367 -1053
rect 14423 -1079 14453 -1053
rect 14509 -1079 14539 -1053
rect 14595 -1079 14625 -1053
rect 14681 -1079 14711 -1053
rect 14766 -1079 14796 -1053
rect 14852 -1079 14882 -1053
rect 14938 -1079 14968 -1053
rect 15024 -1079 15054 -1053
rect 15110 -1079 15140 -1053
rect 15196 -1079 15226 -1053
rect 15282 -1079 15312 -1053
rect 15368 -1079 15398 -1053
rect 15666 -1079 16612 -1053
rect -2918 -1147 -2340 -1121
rect -1538 -1147 -960 -1121
rect -802 -1147 -224 -1121
rect 26 -1147 236 -1121
rect 488 -1147 518 -1121
rect 590 -1147 690 -1121
rect 850 -1147 950 -1121
rect 1015 -1147 1045 -1121
rect 1314 -1147 1524 -1121
rect 1774 -1147 2352 -1121
rect 2602 -1147 2812 -1121
rect 3064 -1147 3094 -1121
rect 3166 -1147 3266 -1121
rect 3426 -1147 3526 -1121
rect 3591 -1147 3621 -1121
rect 3890 -1147 4100 -1121
rect 4350 -1147 4928 -1121
rect 5178 -1147 5388 -1121
rect 5640 -1147 5670 -1121
rect 5742 -1147 5842 -1121
rect 6002 -1147 6102 -1121
rect 6167 -1147 6197 -1121
rect 6466 -1147 6676 -1121
rect 6926 -1147 7504 -1121
rect 7754 -1147 7964 -1121
rect 8216 -1147 8246 -1121
rect 8318 -1147 8418 -1121
rect 8578 -1147 8678 -1121
rect 8743 -1147 8773 -1121
rect 9042 -1147 9252 -1121
rect 9502 -1147 10080 -1121
rect 10422 -1147 10632 -1121
rect 10792 -1147 10822 -1121
rect 10894 -1147 10994 -1121
rect 11154 -1147 11254 -1121
rect 11319 -1147 11349 -1121
rect 11710 -1147 11920 -1121
rect 12547 -1147 12577 -1121
rect 12633 -1147 12663 -1121
rect 12719 -1147 12749 -1121
rect 12805 -1147 12835 -1121
rect 12891 -1147 12921 -1121
rect 12977 -1147 13007 -1121
rect 13274 -1147 13484 -1121
rect 13735 -1147 13765 -1121
rect 13821 -1147 13851 -1121
rect 13907 -1147 13937 -1121
rect 13993 -1147 14023 -1121
rect 14079 -1147 14109 -1121
rect 14165 -1147 14195 -1121
rect 14251 -1147 14281 -1121
rect 14337 -1147 14367 -1121
rect 14423 -1147 14453 -1121
rect 14509 -1147 14539 -1121
rect 14595 -1147 14625 -1121
rect 14681 -1147 14711 -1121
rect 14766 -1147 14796 -1121
rect 14852 -1147 14882 -1121
rect 14938 -1147 14968 -1121
rect 15024 -1147 15054 -1121
rect 15110 -1147 15140 -1121
rect 15196 -1147 15226 -1121
rect 15282 -1147 15312 -1121
rect 15368 -1147 15398 -1121
rect 15666 -1147 16612 -1121
rect -2918 -1347 -2340 -1321
rect -1538 -1347 -960 -1321
rect -802 -1347 -224 -1321
rect 26 -1347 236 -1321
rect -2918 -1369 -2654 -1347
rect -2918 -1403 -2902 -1369
rect -2868 -1403 -2803 -1369
rect -2769 -1403 -2704 -1369
rect -2670 -1403 -2654 -1369
rect -1538 -1369 -1274 -1347
rect -2918 -1419 -2654 -1403
rect -2612 -1405 -2340 -1389
rect -2612 -1439 -2596 -1405
rect -2562 -1439 -2493 -1405
rect -2459 -1439 -2390 -1405
rect -2356 -1439 -2340 -1405
rect -1538 -1403 -1522 -1369
rect -1488 -1403 -1423 -1369
rect -1389 -1403 -1324 -1369
rect -1290 -1403 -1274 -1369
rect -802 -1369 -538 -1347
rect -1538 -1419 -1274 -1403
rect -1232 -1405 -960 -1389
rect -2612 -1461 -2340 -1439
rect -1232 -1439 -1216 -1405
rect -1182 -1439 -1113 -1405
rect -1079 -1439 -1010 -1405
rect -976 -1439 -960 -1405
rect -802 -1403 -786 -1369
rect -752 -1403 -687 -1369
rect -653 -1403 -588 -1369
rect -554 -1403 -538 -1369
rect 152 -1353 236 -1347
rect 152 -1369 294 -1353
rect -802 -1419 -538 -1403
rect -496 -1405 -224 -1389
rect -1232 -1461 -960 -1439
rect -496 -1439 -480 -1405
rect -446 -1439 -377 -1405
rect -343 -1439 -274 -1405
rect -240 -1439 -224 -1405
rect -496 -1461 -224 -1439
rect -32 -1405 110 -1389
rect -32 -1439 -16 -1405
rect 18 -1439 110 -1405
rect 152 -1403 244 -1369
rect 278 -1403 294 -1369
rect 488 -1382 518 -1347
rect 152 -1419 294 -1403
rect 448 -1395 518 -1382
rect 590 -1385 690 -1311
rect 850 -1385 950 -1311
rect 1314 -1347 1524 -1321
rect 1015 -1379 1045 -1347
rect 1440 -1353 1524 -1347
rect 1774 -1347 2352 -1321
rect 2602 -1347 2812 -1321
rect 1440 -1369 1582 -1353
rect -32 -1455 110 -1439
rect 448 -1429 464 -1395
rect 498 -1429 518 -1395
rect 448 -1441 518 -1429
rect 568 -1395 690 -1385
rect 568 -1429 584 -1395
rect 618 -1429 690 -1395
rect 568 -1439 690 -1429
rect 789 -1395 950 -1385
rect 789 -1429 805 -1395
rect 839 -1429 950 -1395
rect 789 -1439 950 -1429
rect -2918 -1487 -2340 -1461
rect -1538 -1487 -960 -1461
rect -802 -1487 -224 -1461
rect 26 -1461 110 -1455
rect 26 -1487 236 -1461
rect 488 -1513 518 -1441
rect 590 -1467 690 -1439
rect 850 -1467 950 -1439
rect 995 -1395 1049 -1379
rect 995 -1429 1005 -1395
rect 1039 -1429 1049 -1395
rect 995 -1445 1049 -1429
rect 1256 -1405 1398 -1389
rect 1256 -1439 1272 -1405
rect 1306 -1439 1398 -1405
rect 1440 -1403 1532 -1369
rect 1566 -1403 1582 -1369
rect 1440 -1419 1582 -1403
rect 1774 -1369 2038 -1347
rect 1774 -1403 1790 -1369
rect 1824 -1403 1889 -1369
rect 1923 -1403 1988 -1369
rect 2022 -1403 2038 -1369
rect 2728 -1353 2812 -1347
rect 2728 -1369 2870 -1353
rect 1774 -1419 2038 -1403
rect 2080 -1405 2352 -1389
rect 1015 -1513 1045 -1445
rect 1256 -1455 1398 -1439
rect 1314 -1461 1398 -1455
rect 2080 -1439 2096 -1405
rect 2130 -1439 2199 -1405
rect 2233 -1439 2302 -1405
rect 2336 -1439 2352 -1405
rect 2080 -1461 2352 -1439
rect 2544 -1405 2686 -1389
rect 2544 -1439 2560 -1405
rect 2594 -1439 2686 -1405
rect 2728 -1403 2820 -1369
rect 2854 -1403 2870 -1369
rect 3064 -1382 3094 -1347
rect 2728 -1419 2870 -1403
rect 3024 -1395 3094 -1382
rect 3166 -1385 3266 -1311
rect 3426 -1385 3526 -1311
rect 3890 -1347 4100 -1321
rect 3591 -1379 3621 -1347
rect 4016 -1353 4100 -1347
rect 4350 -1347 4928 -1321
rect 5178 -1347 5388 -1321
rect 4016 -1369 4158 -1353
rect 2544 -1455 2686 -1439
rect 3024 -1429 3040 -1395
rect 3074 -1429 3094 -1395
rect 3024 -1441 3094 -1429
rect 3144 -1395 3266 -1385
rect 3144 -1429 3160 -1395
rect 3194 -1429 3266 -1395
rect 3144 -1439 3266 -1429
rect 3365 -1395 3526 -1385
rect 3365 -1429 3381 -1395
rect 3415 -1429 3526 -1395
rect 3365 -1439 3526 -1429
rect 1314 -1487 1524 -1461
rect 1774 -1487 2352 -1461
rect 2602 -1461 2686 -1455
rect 2602 -1487 2812 -1461
rect 3064 -1513 3094 -1441
rect 3166 -1467 3266 -1439
rect 3426 -1467 3526 -1439
rect 3571 -1395 3625 -1379
rect 3571 -1429 3581 -1395
rect 3615 -1429 3625 -1395
rect 3571 -1445 3625 -1429
rect 3832 -1405 3974 -1389
rect 3832 -1439 3848 -1405
rect 3882 -1439 3974 -1405
rect 4016 -1403 4108 -1369
rect 4142 -1403 4158 -1369
rect 4016 -1419 4158 -1403
rect 4350 -1369 4614 -1347
rect 4350 -1403 4366 -1369
rect 4400 -1403 4465 -1369
rect 4499 -1403 4564 -1369
rect 4598 -1403 4614 -1369
rect 5304 -1353 5388 -1347
rect 5304 -1369 5446 -1353
rect 4350 -1419 4614 -1403
rect 4656 -1405 4928 -1389
rect 3591 -1513 3621 -1445
rect 3832 -1455 3974 -1439
rect 3890 -1461 3974 -1455
rect 4656 -1439 4672 -1405
rect 4706 -1439 4775 -1405
rect 4809 -1439 4878 -1405
rect 4912 -1439 4928 -1405
rect 4656 -1461 4928 -1439
rect 5120 -1405 5262 -1389
rect 5120 -1439 5136 -1405
rect 5170 -1439 5262 -1405
rect 5304 -1403 5396 -1369
rect 5430 -1403 5446 -1369
rect 5640 -1382 5670 -1347
rect 5304 -1419 5446 -1403
rect 5600 -1395 5670 -1382
rect 5742 -1385 5842 -1311
rect 6002 -1385 6102 -1311
rect 6466 -1347 6676 -1321
rect 6167 -1379 6197 -1347
rect 6592 -1353 6676 -1347
rect 6926 -1347 7504 -1321
rect 7754 -1347 7964 -1321
rect 6592 -1369 6734 -1353
rect 5120 -1455 5262 -1439
rect 5600 -1429 5616 -1395
rect 5650 -1429 5670 -1395
rect 5600 -1441 5670 -1429
rect 5720 -1395 5842 -1385
rect 5720 -1429 5736 -1395
rect 5770 -1429 5842 -1395
rect 5720 -1439 5842 -1429
rect 5941 -1395 6102 -1385
rect 5941 -1429 5957 -1395
rect 5991 -1429 6102 -1395
rect 5941 -1439 6102 -1429
rect 3890 -1487 4100 -1461
rect 4350 -1487 4928 -1461
rect 5178 -1461 5262 -1455
rect 5178 -1487 5388 -1461
rect 5640 -1513 5670 -1441
rect 5742 -1467 5842 -1439
rect 6002 -1467 6102 -1439
rect 6147 -1395 6201 -1379
rect 6147 -1429 6157 -1395
rect 6191 -1429 6201 -1395
rect 6147 -1445 6201 -1429
rect 6408 -1405 6550 -1389
rect 6408 -1439 6424 -1405
rect 6458 -1439 6550 -1405
rect 6592 -1403 6684 -1369
rect 6718 -1403 6734 -1369
rect 6592 -1419 6734 -1403
rect 6926 -1369 7190 -1347
rect 6926 -1403 6942 -1369
rect 6976 -1403 7041 -1369
rect 7075 -1403 7140 -1369
rect 7174 -1403 7190 -1369
rect 7880 -1353 7964 -1347
rect 7880 -1369 8022 -1353
rect 6926 -1419 7190 -1403
rect 7232 -1405 7504 -1389
rect 6167 -1513 6197 -1445
rect 6408 -1455 6550 -1439
rect 6466 -1461 6550 -1455
rect 7232 -1439 7248 -1405
rect 7282 -1439 7351 -1405
rect 7385 -1439 7454 -1405
rect 7488 -1439 7504 -1405
rect 7232 -1461 7504 -1439
rect 7696 -1405 7838 -1389
rect 7696 -1439 7712 -1405
rect 7746 -1439 7838 -1405
rect 7880 -1403 7972 -1369
rect 8006 -1403 8022 -1369
rect 8216 -1382 8246 -1347
rect 7880 -1419 8022 -1403
rect 8176 -1395 8246 -1382
rect 8318 -1385 8418 -1311
rect 8578 -1385 8678 -1311
rect 9042 -1347 9252 -1321
rect 8743 -1379 8773 -1347
rect 9168 -1353 9252 -1347
rect 9502 -1347 10080 -1321
rect 10422 -1347 10632 -1321
rect 9168 -1369 9310 -1353
rect 7696 -1455 7838 -1439
rect 8176 -1429 8192 -1395
rect 8226 -1429 8246 -1395
rect 8176 -1441 8246 -1429
rect 8296 -1395 8418 -1385
rect 8296 -1429 8312 -1395
rect 8346 -1429 8418 -1395
rect 8296 -1439 8418 -1429
rect 8517 -1395 8678 -1385
rect 8517 -1429 8533 -1395
rect 8567 -1429 8678 -1395
rect 8517 -1439 8678 -1429
rect 6466 -1487 6676 -1461
rect 6926 -1487 7504 -1461
rect 7754 -1461 7838 -1455
rect 7754 -1487 7964 -1461
rect 8216 -1513 8246 -1441
rect 8318 -1467 8418 -1439
rect 8578 -1467 8678 -1439
rect 8723 -1395 8777 -1379
rect 8723 -1429 8733 -1395
rect 8767 -1429 8777 -1395
rect 8723 -1445 8777 -1429
rect 8984 -1405 9126 -1389
rect 8984 -1439 9000 -1405
rect 9034 -1439 9126 -1405
rect 9168 -1403 9260 -1369
rect 9294 -1403 9310 -1369
rect 9168 -1419 9310 -1403
rect 9502 -1369 9766 -1347
rect 9502 -1403 9518 -1369
rect 9552 -1403 9617 -1369
rect 9651 -1403 9716 -1369
rect 9750 -1403 9766 -1369
rect 10548 -1353 10632 -1347
rect 10548 -1369 10690 -1353
rect 9502 -1419 9766 -1403
rect 9808 -1405 10080 -1389
rect 8743 -1513 8773 -1445
rect 8984 -1455 9126 -1439
rect 9042 -1461 9126 -1455
rect 9808 -1439 9824 -1405
rect 9858 -1439 9927 -1405
rect 9961 -1439 10030 -1405
rect 10064 -1439 10080 -1405
rect 9808 -1461 10080 -1439
rect 10364 -1405 10506 -1389
rect 10364 -1439 10380 -1405
rect 10414 -1439 10506 -1405
rect 10548 -1403 10640 -1369
rect 10674 -1403 10690 -1369
rect 10792 -1382 10822 -1347
rect 10548 -1419 10690 -1403
rect 10752 -1395 10822 -1382
rect 10894 -1385 10994 -1311
rect 11154 -1385 11254 -1311
rect 11710 -1347 11920 -1321
rect 13274 -1347 13484 -1321
rect 15666 -1347 16612 -1321
rect 11319 -1379 11349 -1347
rect 11836 -1353 11920 -1347
rect 11836 -1369 11978 -1353
rect 10364 -1455 10506 -1439
rect 10752 -1429 10768 -1395
rect 10802 -1429 10822 -1395
rect 10752 -1441 10822 -1429
rect 10872 -1395 10994 -1385
rect 10872 -1429 10888 -1395
rect 10922 -1429 10994 -1395
rect 10872 -1439 10994 -1429
rect 11093 -1395 11254 -1385
rect 11093 -1429 11109 -1395
rect 11143 -1429 11254 -1395
rect 11093 -1439 11254 -1429
rect 9042 -1487 9252 -1461
rect 9502 -1487 10080 -1461
rect 10422 -1461 10506 -1455
rect 10422 -1487 10632 -1461
rect 10792 -1513 10822 -1441
rect 10894 -1467 10994 -1439
rect 11154 -1467 11254 -1439
rect 11299 -1395 11353 -1379
rect 11299 -1429 11309 -1395
rect 11343 -1429 11353 -1395
rect 11299 -1445 11353 -1429
rect 11652 -1405 11794 -1389
rect 11652 -1439 11668 -1405
rect 11702 -1439 11794 -1405
rect 11836 -1403 11928 -1369
rect 11962 -1403 11978 -1369
rect 11836 -1419 11978 -1403
rect 12547 -1385 12577 -1347
rect 12633 -1385 12663 -1347
rect 12719 -1385 12749 -1347
rect 12805 -1385 12835 -1347
rect 12891 -1385 12921 -1347
rect 12977 -1385 13007 -1347
rect 13274 -1353 13358 -1347
rect 12547 -1395 13007 -1385
rect 12547 -1429 12574 -1395
rect 12608 -1429 12642 -1395
rect 12676 -1429 12710 -1395
rect 12744 -1429 12778 -1395
rect 12812 -1429 12846 -1395
rect 12880 -1429 12914 -1395
rect 12948 -1429 13007 -1395
rect 13216 -1369 13358 -1353
rect 13735 -1362 13765 -1347
rect 13821 -1362 13851 -1347
rect 13907 -1362 13937 -1347
rect 13993 -1362 14023 -1347
rect 13216 -1403 13232 -1369
rect 13266 -1403 13358 -1369
rect 13216 -1419 13358 -1403
rect 13400 -1405 13542 -1389
rect 12547 -1439 13007 -1429
rect 13400 -1439 13492 -1405
rect 13526 -1439 13542 -1405
rect 11319 -1513 11349 -1445
rect 11652 -1455 11794 -1439
rect 11710 -1461 11794 -1455
rect 11710 -1487 11920 -1461
rect 12633 -1513 12663 -1439
rect 12719 -1513 12749 -1439
rect 12805 -1513 12835 -1439
rect 12891 -1513 12921 -1439
rect 13400 -1455 13542 -1439
rect 13676 -1395 14023 -1362
rect 13676 -1429 13692 -1395
rect 13726 -1429 14023 -1395
rect 13400 -1461 13484 -1455
rect 13274 -1487 13484 -1461
rect 13676 -1464 14023 -1429
rect 13735 -1513 13765 -1464
rect 13821 -1513 13851 -1464
rect 13907 -1513 13937 -1464
rect 13993 -1513 14023 -1464
rect 14079 -1379 14109 -1347
rect 14165 -1379 14195 -1347
rect 14251 -1379 14281 -1347
rect 14337 -1379 14367 -1347
rect 14423 -1379 14453 -1347
rect 14509 -1379 14539 -1347
rect 14595 -1379 14625 -1347
rect 14681 -1379 14711 -1347
rect 14766 -1379 14796 -1347
rect 14852 -1379 14882 -1347
rect 14938 -1379 14968 -1347
rect 15024 -1379 15054 -1347
rect 15110 -1379 15140 -1347
rect 15196 -1379 15226 -1347
rect 15282 -1379 15312 -1347
rect 15368 -1379 15398 -1347
rect 14079 -1395 15398 -1379
rect 14079 -1429 14119 -1395
rect 14153 -1429 14187 -1395
rect 14221 -1429 14255 -1395
rect 14289 -1429 14323 -1395
rect 14357 -1429 14391 -1395
rect 14425 -1429 14459 -1395
rect 14493 -1429 14527 -1395
rect 14561 -1429 14595 -1395
rect 14629 -1429 14663 -1395
rect 14697 -1429 14731 -1395
rect 14765 -1429 14799 -1395
rect 14833 -1429 14867 -1395
rect 14901 -1429 14935 -1395
rect 14969 -1429 15003 -1395
rect 15037 -1429 15071 -1395
rect 15105 -1429 15139 -1395
rect 15173 -1429 15398 -1395
rect 15666 -1369 16116 -1347
rect 15666 -1403 15682 -1369
rect 15716 -1403 15810 -1369
rect 15844 -1403 15938 -1369
rect 15972 -1403 16066 -1369
rect 16100 -1403 16116 -1369
rect 15666 -1419 16116 -1403
rect 16158 -1405 16612 -1389
rect 14079 -1454 15398 -1429
rect 14079 -1513 14109 -1454
rect 14165 -1513 14195 -1454
rect 14251 -1513 14281 -1454
rect 14337 -1513 14367 -1454
rect 14423 -1513 14453 -1454
rect 14509 -1513 14539 -1454
rect 14595 -1513 14625 -1454
rect 14681 -1513 14711 -1454
rect 14766 -1513 14796 -1454
rect 14852 -1513 14882 -1454
rect 14938 -1513 14968 -1454
rect 15024 -1513 15054 -1454
rect 15110 -1513 15140 -1454
rect 15196 -1513 15226 -1454
rect 15282 -1513 15312 -1454
rect 15368 -1513 15398 -1454
rect 16158 -1439 16174 -1405
rect 16208 -1439 16302 -1405
rect 16336 -1439 16430 -1405
rect 16464 -1439 16558 -1405
rect 16592 -1439 16612 -1405
rect 16158 -1461 16612 -1439
rect 15666 -1487 16612 -1461
rect -2918 -1623 -2340 -1597
rect -1538 -1623 -960 -1597
rect -802 -1623 -224 -1597
rect 26 -1623 236 -1597
rect 488 -1623 518 -1597
rect 590 -1623 690 -1597
rect 850 -1623 950 -1597
rect 1015 -1623 1045 -1597
rect 1314 -1623 1524 -1597
rect 1774 -1623 2352 -1597
rect 2602 -1623 2812 -1597
rect 3064 -1623 3094 -1597
rect 3166 -1623 3266 -1597
rect 3426 -1623 3526 -1597
rect 3591 -1623 3621 -1597
rect 3890 -1623 4100 -1597
rect 4350 -1623 4928 -1597
rect 5178 -1623 5388 -1597
rect 5640 -1623 5670 -1597
rect 5742 -1623 5842 -1597
rect 6002 -1623 6102 -1597
rect 6167 -1623 6197 -1597
rect 6466 -1623 6676 -1597
rect 6926 -1623 7504 -1597
rect 7754 -1623 7964 -1597
rect 8216 -1623 8246 -1597
rect 8318 -1623 8418 -1597
rect 8578 -1623 8678 -1597
rect 8743 -1623 8773 -1597
rect 9042 -1623 9252 -1597
rect 9502 -1623 10080 -1597
rect 10422 -1623 10632 -1597
rect 10792 -1623 10822 -1597
rect 10894 -1623 10994 -1597
rect 11154 -1623 11254 -1597
rect 11319 -1623 11349 -1597
rect 11710 -1623 11920 -1597
rect 12633 -1623 12663 -1597
rect 12719 -1623 12749 -1597
rect 12805 -1623 12835 -1597
rect 12891 -1623 12921 -1597
rect 13274 -1623 13484 -1597
rect 13735 -1623 13765 -1597
rect 13821 -1623 13851 -1597
rect 13907 -1623 13937 -1597
rect 13993 -1623 14023 -1597
rect 14079 -1623 14109 -1597
rect 14165 -1623 14195 -1597
rect 14251 -1623 14281 -1597
rect 14337 -1623 14367 -1597
rect 14423 -1623 14453 -1597
rect 14509 -1623 14539 -1597
rect 14595 -1623 14625 -1597
rect 14681 -1623 14711 -1597
rect 14766 -1623 14796 -1597
rect 14852 -1623 14882 -1597
rect 14938 -1623 14968 -1597
rect 15024 -1623 15054 -1597
rect 15110 -1623 15140 -1597
rect 15196 -1623 15226 -1597
rect 15282 -1623 15312 -1597
rect 15368 -1623 15398 -1597
rect 15666 -1623 16612 -1597
rect -2918 -1691 -2340 -1665
rect -1538 -1691 -960 -1665
rect -783 -1691 -753 -1665
rect -688 -1691 -588 -1665
rect -428 -1691 -328 -1665
rect -256 -1691 -226 -1665
rect 26 -1691 236 -1665
rect 505 -1691 535 -1665
rect 600 -1691 700 -1665
rect 860 -1691 960 -1665
rect 1032 -1691 1062 -1665
rect 1314 -1691 1524 -1665
rect 1774 -1691 2352 -1665
rect 2602 -1691 2812 -1665
rect 3081 -1691 3111 -1665
rect 3176 -1691 3276 -1665
rect 3436 -1691 3536 -1665
rect 3608 -1691 3638 -1665
rect 3890 -1691 4100 -1665
rect 4350 -1691 4928 -1665
rect 5178 -1691 5388 -1665
rect 5657 -1691 5687 -1665
rect 5752 -1691 5852 -1665
rect 6012 -1691 6112 -1665
rect 6184 -1691 6214 -1665
rect 6466 -1691 6676 -1665
rect 6926 -1691 7504 -1665
rect 7754 -1691 7964 -1665
rect 8233 -1691 8263 -1665
rect 8328 -1691 8428 -1665
rect 8588 -1691 8688 -1665
rect 8760 -1691 8790 -1665
rect 9042 -1691 9252 -1665
rect 9502 -1691 10080 -1665
rect 10422 -1691 10632 -1665
rect 10809 -1691 10839 -1665
rect 10904 -1691 11004 -1665
rect 11164 -1691 11264 -1665
rect 11336 -1691 11366 -1665
rect 11710 -1691 11920 -1665
rect 13735 -1691 13765 -1665
rect 13821 -1691 13851 -1665
rect 13907 -1691 13937 -1665
rect 13993 -1691 14023 -1665
rect 14079 -1691 14109 -1665
rect 14165 -1691 14195 -1665
rect 14251 -1691 14281 -1665
rect 14337 -1691 14367 -1665
rect 14423 -1691 14453 -1665
rect 14509 -1691 14539 -1665
rect 14595 -1691 14625 -1665
rect 14681 -1691 14711 -1665
rect 14766 -1691 14796 -1665
rect 14852 -1691 14882 -1665
rect 14938 -1691 14968 -1665
rect 15024 -1691 15054 -1665
rect 15110 -1691 15140 -1665
rect 15196 -1691 15226 -1665
rect 15282 -1691 15312 -1665
rect 15368 -1691 15398 -1665
rect 15666 -1691 16612 -1665
rect -2918 -1827 -2340 -1801
rect -1538 -1827 -960 -1801
rect -2918 -1849 -2646 -1827
rect -2918 -1883 -2902 -1849
rect -2868 -1883 -2799 -1849
rect -2765 -1883 -2696 -1849
rect -2662 -1883 -2646 -1849
rect -1538 -1849 -1266 -1827
rect -783 -1843 -753 -1775
rect -2918 -1899 -2646 -1883
rect -2604 -1885 -2340 -1869
rect -2604 -1919 -2588 -1885
rect -2554 -1919 -2489 -1885
rect -2455 -1919 -2390 -1885
rect -2356 -1919 -2340 -1885
rect -1538 -1883 -1522 -1849
rect -1488 -1883 -1419 -1849
rect -1385 -1883 -1316 -1849
rect -1282 -1883 -1266 -1849
rect -787 -1859 -733 -1843
rect -1538 -1899 -1266 -1883
rect -1224 -1885 -960 -1869
rect -2604 -1941 -2340 -1919
rect -1224 -1919 -1208 -1885
rect -1174 -1919 -1109 -1885
rect -1075 -1919 -1010 -1885
rect -976 -1919 -960 -1885
rect -787 -1893 -777 -1859
rect -743 -1893 -733 -1859
rect -787 -1909 -733 -1893
rect -688 -1849 -588 -1821
rect -428 -1849 -328 -1821
rect -256 -1847 -226 -1775
rect 26 -1827 236 -1801
rect 26 -1833 110 -1827
rect -688 -1859 -527 -1849
rect -688 -1893 -577 -1859
rect -543 -1893 -527 -1859
rect -688 -1903 -527 -1893
rect -428 -1859 -306 -1849
rect -428 -1893 -356 -1859
rect -322 -1893 -306 -1859
rect -428 -1903 -306 -1893
rect -256 -1859 -186 -1847
rect -256 -1893 -236 -1859
rect -202 -1893 -186 -1859
rect -1224 -1941 -960 -1919
rect -783 -1941 -753 -1909
rect -2918 -1967 -2340 -1941
rect -1538 -1967 -960 -1941
rect -688 -1977 -588 -1903
rect -428 -1977 -328 -1903
rect -256 -1906 -186 -1893
rect -32 -1849 110 -1833
rect 505 -1843 535 -1775
rect -32 -1883 -16 -1849
rect 18 -1883 110 -1849
rect 501 -1859 555 -1843
rect -32 -1899 110 -1883
rect 152 -1885 294 -1869
rect -256 -1941 -226 -1906
rect 152 -1919 244 -1885
rect 278 -1919 294 -1885
rect 501 -1893 511 -1859
rect 545 -1893 555 -1859
rect 501 -1909 555 -1893
rect 600 -1849 700 -1821
rect 860 -1849 960 -1821
rect 1032 -1847 1062 -1775
rect 1314 -1827 1524 -1801
rect 1774 -1827 2352 -1801
rect 2602 -1827 2812 -1801
rect 1314 -1833 1398 -1827
rect 600 -1859 761 -1849
rect 600 -1893 711 -1859
rect 745 -1893 761 -1859
rect 600 -1903 761 -1893
rect 860 -1859 982 -1849
rect 860 -1893 932 -1859
rect 966 -1893 982 -1859
rect 860 -1903 982 -1893
rect 1032 -1859 1102 -1847
rect 1032 -1893 1052 -1859
rect 1086 -1893 1102 -1859
rect 152 -1935 294 -1919
rect 152 -1941 236 -1935
rect 505 -1941 535 -1909
rect 26 -1967 236 -1941
rect 600 -1977 700 -1903
rect 860 -1977 960 -1903
rect 1032 -1906 1102 -1893
rect 1256 -1849 1398 -1833
rect 1256 -1883 1272 -1849
rect 1306 -1883 1398 -1849
rect 1774 -1849 2046 -1827
rect 2602 -1833 2686 -1827
rect 1256 -1899 1398 -1883
rect 1440 -1885 1582 -1869
rect 1032 -1941 1062 -1906
rect 1440 -1919 1532 -1885
rect 1566 -1919 1582 -1885
rect 1774 -1883 1790 -1849
rect 1824 -1883 1893 -1849
rect 1927 -1883 1996 -1849
rect 2030 -1883 2046 -1849
rect 2544 -1849 2686 -1833
rect 3081 -1843 3111 -1775
rect 1774 -1899 2046 -1883
rect 2088 -1885 2352 -1869
rect 1440 -1935 1582 -1919
rect 2088 -1919 2104 -1885
rect 2138 -1919 2203 -1885
rect 2237 -1919 2302 -1885
rect 2336 -1919 2352 -1885
rect 2544 -1883 2560 -1849
rect 2594 -1883 2686 -1849
rect 3077 -1859 3131 -1843
rect 2544 -1899 2686 -1883
rect 2728 -1885 2870 -1869
rect 1440 -1941 1524 -1935
rect 2088 -1941 2352 -1919
rect 2728 -1919 2820 -1885
rect 2854 -1919 2870 -1885
rect 3077 -1893 3087 -1859
rect 3121 -1893 3131 -1859
rect 3077 -1909 3131 -1893
rect 3176 -1849 3276 -1821
rect 3436 -1849 3536 -1821
rect 3608 -1847 3638 -1775
rect 3890 -1827 4100 -1801
rect 4350 -1827 4928 -1801
rect 5178 -1827 5388 -1801
rect 3890 -1833 3974 -1827
rect 3176 -1859 3337 -1849
rect 3176 -1893 3287 -1859
rect 3321 -1893 3337 -1859
rect 3176 -1903 3337 -1893
rect 3436 -1859 3558 -1849
rect 3436 -1893 3508 -1859
rect 3542 -1893 3558 -1859
rect 3436 -1903 3558 -1893
rect 3608 -1859 3678 -1847
rect 3608 -1893 3628 -1859
rect 3662 -1893 3678 -1859
rect 2728 -1935 2870 -1919
rect 2728 -1941 2812 -1935
rect 3081 -1941 3111 -1909
rect 1314 -1967 1524 -1941
rect 1774 -1967 2352 -1941
rect 2602 -1967 2812 -1941
rect 3176 -1977 3276 -1903
rect 3436 -1977 3536 -1903
rect 3608 -1906 3678 -1893
rect 3832 -1849 3974 -1833
rect 3832 -1883 3848 -1849
rect 3882 -1883 3974 -1849
rect 4350 -1849 4622 -1827
rect 5178 -1833 5262 -1827
rect 3832 -1899 3974 -1883
rect 4016 -1885 4158 -1869
rect 3608 -1941 3638 -1906
rect 4016 -1919 4108 -1885
rect 4142 -1919 4158 -1885
rect 4350 -1883 4366 -1849
rect 4400 -1883 4469 -1849
rect 4503 -1883 4572 -1849
rect 4606 -1883 4622 -1849
rect 5120 -1849 5262 -1833
rect 5657 -1843 5687 -1775
rect 4350 -1899 4622 -1883
rect 4664 -1885 4928 -1869
rect 4016 -1935 4158 -1919
rect 4664 -1919 4680 -1885
rect 4714 -1919 4779 -1885
rect 4813 -1919 4878 -1885
rect 4912 -1919 4928 -1885
rect 5120 -1883 5136 -1849
rect 5170 -1883 5262 -1849
rect 5653 -1859 5707 -1843
rect 5120 -1899 5262 -1883
rect 5304 -1885 5446 -1869
rect 4016 -1941 4100 -1935
rect 4664 -1941 4928 -1919
rect 5304 -1919 5396 -1885
rect 5430 -1919 5446 -1885
rect 5653 -1893 5663 -1859
rect 5697 -1893 5707 -1859
rect 5653 -1909 5707 -1893
rect 5752 -1849 5852 -1821
rect 6012 -1849 6112 -1821
rect 6184 -1847 6214 -1775
rect 6466 -1827 6676 -1801
rect 6926 -1827 7504 -1801
rect 7754 -1827 7964 -1801
rect 6466 -1833 6550 -1827
rect 5752 -1859 5913 -1849
rect 5752 -1893 5863 -1859
rect 5897 -1893 5913 -1859
rect 5752 -1903 5913 -1893
rect 6012 -1859 6134 -1849
rect 6012 -1893 6084 -1859
rect 6118 -1893 6134 -1859
rect 6012 -1903 6134 -1893
rect 6184 -1859 6254 -1847
rect 6184 -1893 6204 -1859
rect 6238 -1893 6254 -1859
rect 5304 -1935 5446 -1919
rect 5304 -1941 5388 -1935
rect 5657 -1941 5687 -1909
rect 3890 -1967 4100 -1941
rect 4350 -1967 4928 -1941
rect 5178 -1967 5388 -1941
rect 5752 -1977 5852 -1903
rect 6012 -1977 6112 -1903
rect 6184 -1906 6254 -1893
rect 6408 -1849 6550 -1833
rect 6408 -1883 6424 -1849
rect 6458 -1883 6550 -1849
rect 6926 -1849 7198 -1827
rect 7754 -1833 7838 -1827
rect 6408 -1899 6550 -1883
rect 6592 -1885 6734 -1869
rect 6184 -1941 6214 -1906
rect 6592 -1919 6684 -1885
rect 6718 -1919 6734 -1885
rect 6926 -1883 6942 -1849
rect 6976 -1883 7045 -1849
rect 7079 -1883 7148 -1849
rect 7182 -1883 7198 -1849
rect 7696 -1849 7838 -1833
rect 8233 -1843 8263 -1775
rect 6926 -1899 7198 -1883
rect 7240 -1885 7504 -1869
rect 6592 -1935 6734 -1919
rect 7240 -1919 7256 -1885
rect 7290 -1919 7355 -1885
rect 7389 -1919 7454 -1885
rect 7488 -1919 7504 -1885
rect 7696 -1883 7712 -1849
rect 7746 -1883 7838 -1849
rect 8229 -1859 8283 -1843
rect 7696 -1899 7838 -1883
rect 7880 -1885 8022 -1869
rect 6592 -1941 6676 -1935
rect 7240 -1941 7504 -1919
rect 7880 -1919 7972 -1885
rect 8006 -1919 8022 -1885
rect 8229 -1893 8239 -1859
rect 8273 -1893 8283 -1859
rect 8229 -1909 8283 -1893
rect 8328 -1849 8428 -1821
rect 8588 -1849 8688 -1821
rect 8760 -1847 8790 -1775
rect 9042 -1827 9252 -1801
rect 9502 -1827 10080 -1801
rect 10422 -1827 10632 -1801
rect 9042 -1833 9126 -1827
rect 8328 -1859 8489 -1849
rect 8328 -1893 8439 -1859
rect 8473 -1893 8489 -1859
rect 8328 -1903 8489 -1893
rect 8588 -1859 8710 -1849
rect 8588 -1893 8660 -1859
rect 8694 -1893 8710 -1859
rect 8588 -1903 8710 -1893
rect 8760 -1859 8830 -1847
rect 8760 -1893 8780 -1859
rect 8814 -1893 8830 -1859
rect 7880 -1935 8022 -1919
rect 7880 -1941 7964 -1935
rect 8233 -1941 8263 -1909
rect 6466 -1967 6676 -1941
rect 6926 -1967 7504 -1941
rect 7754 -1967 7964 -1941
rect 8328 -1977 8428 -1903
rect 8588 -1977 8688 -1903
rect 8760 -1906 8830 -1893
rect 8984 -1849 9126 -1833
rect 8984 -1883 9000 -1849
rect 9034 -1883 9126 -1849
rect 9502 -1849 9774 -1827
rect 10422 -1833 10506 -1827
rect 8984 -1899 9126 -1883
rect 9168 -1885 9310 -1869
rect 8760 -1941 8790 -1906
rect 9168 -1919 9260 -1885
rect 9294 -1919 9310 -1885
rect 9502 -1883 9518 -1849
rect 9552 -1883 9621 -1849
rect 9655 -1883 9724 -1849
rect 9758 -1883 9774 -1849
rect 10364 -1849 10506 -1833
rect 10809 -1843 10839 -1775
rect 9502 -1899 9774 -1883
rect 9816 -1885 10080 -1869
rect 9168 -1935 9310 -1919
rect 9816 -1919 9832 -1885
rect 9866 -1919 9931 -1885
rect 9965 -1919 10030 -1885
rect 10064 -1919 10080 -1885
rect 10364 -1883 10380 -1849
rect 10414 -1883 10506 -1849
rect 10805 -1859 10859 -1843
rect 10364 -1899 10506 -1883
rect 10548 -1885 10690 -1869
rect 9168 -1941 9252 -1935
rect 9816 -1941 10080 -1919
rect 10548 -1919 10640 -1885
rect 10674 -1919 10690 -1885
rect 10805 -1893 10815 -1859
rect 10849 -1893 10859 -1859
rect 10805 -1909 10859 -1893
rect 10904 -1849 11004 -1821
rect 11164 -1849 11264 -1821
rect 11336 -1847 11366 -1775
rect 11710 -1827 11920 -1801
rect 13735 -1824 13765 -1775
rect 13821 -1824 13851 -1775
rect 13907 -1824 13937 -1775
rect 13993 -1824 14023 -1775
rect 11710 -1833 11794 -1827
rect 10904 -1859 11065 -1849
rect 10904 -1893 11015 -1859
rect 11049 -1893 11065 -1859
rect 10904 -1903 11065 -1893
rect 11164 -1859 11286 -1849
rect 11164 -1893 11236 -1859
rect 11270 -1893 11286 -1859
rect 11164 -1903 11286 -1893
rect 11336 -1859 11406 -1847
rect 11336 -1893 11356 -1859
rect 11390 -1893 11406 -1859
rect 10548 -1935 10690 -1919
rect 10548 -1941 10632 -1935
rect 10809 -1941 10839 -1909
rect 9042 -1967 9252 -1941
rect 9502 -1967 10080 -1941
rect 10422 -1967 10632 -1941
rect 10904 -1977 11004 -1903
rect 11164 -1977 11264 -1903
rect 11336 -1906 11406 -1893
rect 11652 -1849 11794 -1833
rect 11652 -1883 11668 -1849
rect 11702 -1883 11794 -1849
rect 13676 -1859 14023 -1824
rect 11652 -1899 11794 -1883
rect 11836 -1885 11978 -1869
rect 11336 -1941 11366 -1906
rect 11836 -1919 11928 -1885
rect 11962 -1919 11978 -1885
rect 11836 -1935 11978 -1919
rect 13676 -1893 13692 -1859
rect 13726 -1893 14023 -1859
rect 13676 -1926 14023 -1893
rect 11836 -1941 11920 -1935
rect 13735 -1941 13765 -1926
rect 13821 -1941 13851 -1926
rect 13907 -1941 13937 -1926
rect 13993 -1941 14023 -1926
rect 14079 -1834 14109 -1775
rect 14165 -1834 14195 -1775
rect 14251 -1834 14281 -1775
rect 14337 -1834 14367 -1775
rect 14423 -1834 14453 -1775
rect 14509 -1834 14539 -1775
rect 14595 -1834 14625 -1775
rect 14681 -1834 14711 -1775
rect 14766 -1834 14796 -1775
rect 14852 -1834 14882 -1775
rect 14938 -1834 14968 -1775
rect 15024 -1834 15054 -1775
rect 15110 -1834 15140 -1775
rect 15196 -1834 15226 -1775
rect 15282 -1834 15312 -1775
rect 15368 -1834 15398 -1775
rect 14079 -1859 15398 -1834
rect 14079 -1893 14119 -1859
rect 14153 -1893 14187 -1859
rect 14221 -1893 14255 -1859
rect 14289 -1893 14323 -1859
rect 14357 -1893 14391 -1859
rect 14425 -1893 14459 -1859
rect 14493 -1893 14527 -1859
rect 14561 -1893 14595 -1859
rect 14629 -1893 14663 -1859
rect 14697 -1893 14731 -1859
rect 14765 -1893 14799 -1859
rect 14833 -1893 14867 -1859
rect 14901 -1893 14935 -1859
rect 14969 -1893 15003 -1859
rect 15037 -1893 15071 -1859
rect 15105 -1893 15139 -1859
rect 15173 -1893 15398 -1859
rect 14079 -1909 15398 -1893
rect 15666 -1827 16612 -1801
rect 15666 -1849 16120 -1827
rect 15666 -1883 15686 -1849
rect 15720 -1883 15814 -1849
rect 15848 -1883 15942 -1849
rect 15976 -1883 16070 -1849
rect 16104 -1883 16120 -1849
rect 15666 -1899 16120 -1883
rect 16162 -1885 16612 -1869
rect 14079 -1941 14109 -1909
rect 14165 -1941 14195 -1909
rect 14251 -1941 14281 -1909
rect 14337 -1941 14367 -1909
rect 14423 -1941 14453 -1909
rect 14509 -1941 14539 -1909
rect 14595 -1941 14625 -1909
rect 14681 -1941 14711 -1909
rect 14766 -1941 14796 -1909
rect 14852 -1941 14882 -1909
rect 14938 -1941 14968 -1909
rect 15024 -1941 15054 -1909
rect 15110 -1941 15140 -1909
rect 15196 -1941 15226 -1909
rect 15282 -1941 15312 -1909
rect 15368 -1941 15398 -1909
rect 16162 -1919 16178 -1885
rect 16212 -1919 16306 -1885
rect 16340 -1919 16434 -1885
rect 16468 -1919 16562 -1885
rect 16596 -1919 16612 -1885
rect 16162 -1941 16612 -1919
rect 11710 -1967 11920 -1941
rect 15666 -1967 16612 -1941
rect -2918 -2167 -2340 -2141
rect -1538 -2167 -960 -2141
rect -783 -2167 -753 -2141
rect -688 -2167 -588 -2141
rect -428 -2167 -328 -2141
rect -256 -2167 -226 -2141
rect 26 -2167 236 -2141
rect 505 -2167 535 -2141
rect 600 -2167 700 -2141
rect 860 -2167 960 -2141
rect 1032 -2167 1062 -2141
rect 1314 -2167 1524 -2141
rect 1774 -2167 2352 -2141
rect 2602 -2167 2812 -2141
rect 3081 -2167 3111 -2141
rect 3176 -2167 3276 -2141
rect 3436 -2167 3536 -2141
rect 3608 -2167 3638 -2141
rect 3890 -2167 4100 -2141
rect 4350 -2167 4928 -2141
rect 5178 -2167 5388 -2141
rect 5657 -2167 5687 -2141
rect 5752 -2167 5852 -2141
rect 6012 -2167 6112 -2141
rect 6184 -2167 6214 -2141
rect 6466 -2167 6676 -2141
rect 6926 -2167 7504 -2141
rect 7754 -2167 7964 -2141
rect 8233 -2167 8263 -2141
rect 8328 -2167 8428 -2141
rect 8588 -2167 8688 -2141
rect 8760 -2167 8790 -2141
rect 9042 -2167 9252 -2141
rect 9502 -2167 10080 -2141
rect 10422 -2167 10632 -2141
rect 10809 -2167 10839 -2141
rect 10904 -2167 11004 -2141
rect 11164 -2167 11264 -2141
rect 11336 -2167 11366 -2141
rect 11710 -2167 11920 -2141
rect 13735 -2167 13765 -2141
rect 13821 -2167 13851 -2141
rect 13907 -2167 13937 -2141
rect 13993 -2167 14023 -2141
rect 14079 -2167 14109 -2141
rect 14165 -2167 14195 -2141
rect 14251 -2167 14281 -2141
rect 14337 -2167 14367 -2141
rect 14423 -2167 14453 -2141
rect 14509 -2167 14539 -2141
rect 14595 -2167 14625 -2141
rect 14681 -2167 14711 -2141
rect 14766 -2167 14796 -2141
rect 14852 -2167 14882 -2141
rect 14938 -2167 14968 -2141
rect 15024 -2167 15054 -2141
rect 15110 -2167 15140 -2141
rect 15196 -2167 15226 -2141
rect 15282 -2167 15312 -2141
rect 15368 -2167 15398 -2141
rect 15666 -2167 16612 -2141
rect -2918 -2235 -2340 -2209
rect -1538 -2235 -960 -2209
rect -802 -2235 -224 -2209
rect 26 -2235 236 -2209
rect 488 -2235 518 -2209
rect 590 -2235 690 -2209
rect 850 -2235 950 -2209
rect 1015 -2235 1045 -2209
rect 1314 -2235 1524 -2209
rect 1774 -2235 2352 -2209
rect 2602 -2235 2812 -2209
rect 3064 -2235 3094 -2209
rect 3166 -2235 3266 -2209
rect 3426 -2235 3526 -2209
rect 3591 -2235 3621 -2209
rect 3890 -2235 4100 -2209
rect 4350 -2235 4928 -2209
rect 5178 -2235 5388 -2209
rect 5640 -2235 5670 -2209
rect 5742 -2235 5842 -2209
rect 6002 -2235 6102 -2209
rect 6167 -2235 6197 -2209
rect 6466 -2235 6676 -2209
rect 6926 -2235 7504 -2209
rect 7754 -2235 7964 -2209
rect 8216 -2235 8246 -2209
rect 8318 -2235 8418 -2209
rect 8578 -2235 8678 -2209
rect 8743 -2235 8773 -2209
rect 9042 -2235 9252 -2209
rect 9502 -2235 10080 -2209
rect 10422 -2235 10632 -2209
rect 10792 -2235 10822 -2209
rect 10894 -2235 10994 -2209
rect 11154 -2235 11254 -2209
rect 11319 -2235 11349 -2209
rect 11710 -2235 11920 -2209
rect 12547 -2235 12577 -2209
rect 12633 -2235 12663 -2209
rect 12719 -2235 12749 -2209
rect 12805 -2235 12835 -2209
rect 12891 -2235 12921 -2209
rect 12977 -2235 13007 -2209
rect 13274 -2235 13484 -2209
rect 13735 -2235 13765 -2209
rect 13821 -2235 13851 -2209
rect 13907 -2235 13937 -2209
rect 13993 -2235 14023 -2209
rect 14079 -2235 14109 -2209
rect 14165 -2235 14195 -2209
rect 14251 -2235 14281 -2209
rect 14337 -2235 14367 -2209
rect 14423 -2235 14453 -2209
rect 14509 -2235 14539 -2209
rect 14595 -2235 14625 -2209
rect 14681 -2235 14711 -2209
rect 14766 -2235 14796 -2209
rect 14852 -2235 14882 -2209
rect 14938 -2235 14968 -2209
rect 15024 -2235 15054 -2209
rect 15110 -2235 15140 -2209
rect 15196 -2235 15226 -2209
rect 15282 -2235 15312 -2209
rect 15368 -2235 15398 -2209
rect 15666 -2235 16612 -2209
rect -2918 -2435 -2340 -2409
rect -1538 -2435 -960 -2409
rect -802 -2435 -224 -2409
rect 26 -2435 236 -2409
rect -2918 -2457 -2654 -2435
rect -2918 -2491 -2902 -2457
rect -2868 -2491 -2803 -2457
rect -2769 -2491 -2704 -2457
rect -2670 -2491 -2654 -2457
rect -1538 -2457 -1274 -2435
rect -2918 -2507 -2654 -2491
rect -2612 -2493 -2340 -2477
rect -2612 -2527 -2596 -2493
rect -2562 -2527 -2493 -2493
rect -2459 -2527 -2390 -2493
rect -2356 -2527 -2340 -2493
rect -1538 -2491 -1522 -2457
rect -1488 -2491 -1423 -2457
rect -1389 -2491 -1324 -2457
rect -1290 -2491 -1274 -2457
rect -802 -2457 -538 -2435
rect -1538 -2507 -1274 -2491
rect -1232 -2493 -960 -2477
rect -2612 -2549 -2340 -2527
rect -1232 -2527 -1216 -2493
rect -1182 -2527 -1113 -2493
rect -1079 -2527 -1010 -2493
rect -976 -2527 -960 -2493
rect -802 -2491 -786 -2457
rect -752 -2491 -687 -2457
rect -653 -2491 -588 -2457
rect -554 -2491 -538 -2457
rect 152 -2441 236 -2435
rect 152 -2457 294 -2441
rect -802 -2507 -538 -2491
rect -496 -2493 -224 -2477
rect -1232 -2549 -960 -2527
rect -496 -2527 -480 -2493
rect -446 -2527 -377 -2493
rect -343 -2527 -274 -2493
rect -240 -2527 -224 -2493
rect -496 -2549 -224 -2527
rect -32 -2493 110 -2477
rect -32 -2527 -16 -2493
rect 18 -2527 110 -2493
rect 152 -2491 244 -2457
rect 278 -2491 294 -2457
rect 488 -2470 518 -2435
rect 152 -2507 294 -2491
rect 448 -2483 518 -2470
rect 590 -2473 690 -2399
rect 850 -2473 950 -2399
rect 1314 -2435 1524 -2409
rect 1015 -2467 1045 -2435
rect 1440 -2441 1524 -2435
rect 1774 -2435 2352 -2409
rect 2602 -2435 2812 -2409
rect 1440 -2457 1582 -2441
rect -32 -2543 110 -2527
rect 448 -2517 464 -2483
rect 498 -2517 518 -2483
rect 448 -2529 518 -2517
rect 568 -2483 690 -2473
rect 568 -2517 584 -2483
rect 618 -2517 690 -2483
rect 568 -2527 690 -2517
rect 789 -2483 950 -2473
rect 789 -2517 805 -2483
rect 839 -2517 950 -2483
rect 789 -2527 950 -2517
rect -2918 -2575 -2340 -2549
rect -1538 -2575 -960 -2549
rect -802 -2575 -224 -2549
rect 26 -2549 110 -2543
rect 26 -2575 236 -2549
rect 488 -2601 518 -2529
rect 590 -2555 690 -2527
rect 850 -2555 950 -2527
rect 995 -2483 1049 -2467
rect 995 -2517 1005 -2483
rect 1039 -2517 1049 -2483
rect 995 -2533 1049 -2517
rect 1256 -2493 1398 -2477
rect 1256 -2527 1272 -2493
rect 1306 -2527 1398 -2493
rect 1440 -2491 1532 -2457
rect 1566 -2491 1582 -2457
rect 1440 -2507 1582 -2491
rect 1774 -2457 2038 -2435
rect 1774 -2491 1790 -2457
rect 1824 -2491 1889 -2457
rect 1923 -2491 1988 -2457
rect 2022 -2491 2038 -2457
rect 2728 -2441 2812 -2435
rect 2728 -2457 2870 -2441
rect 1774 -2507 2038 -2491
rect 2080 -2493 2352 -2477
rect 1015 -2601 1045 -2533
rect 1256 -2543 1398 -2527
rect 1314 -2549 1398 -2543
rect 2080 -2527 2096 -2493
rect 2130 -2527 2199 -2493
rect 2233 -2527 2302 -2493
rect 2336 -2527 2352 -2493
rect 2080 -2549 2352 -2527
rect 2544 -2493 2686 -2477
rect 2544 -2527 2560 -2493
rect 2594 -2527 2686 -2493
rect 2728 -2491 2820 -2457
rect 2854 -2491 2870 -2457
rect 3064 -2470 3094 -2435
rect 2728 -2507 2870 -2491
rect 3024 -2483 3094 -2470
rect 3166 -2473 3266 -2399
rect 3426 -2473 3526 -2399
rect 3890 -2435 4100 -2409
rect 3591 -2467 3621 -2435
rect 4016 -2441 4100 -2435
rect 4350 -2435 4928 -2409
rect 5178 -2435 5388 -2409
rect 4016 -2457 4158 -2441
rect 2544 -2543 2686 -2527
rect 3024 -2517 3040 -2483
rect 3074 -2517 3094 -2483
rect 3024 -2529 3094 -2517
rect 3144 -2483 3266 -2473
rect 3144 -2517 3160 -2483
rect 3194 -2517 3266 -2483
rect 3144 -2527 3266 -2517
rect 3365 -2483 3526 -2473
rect 3365 -2517 3381 -2483
rect 3415 -2517 3526 -2483
rect 3365 -2527 3526 -2517
rect 1314 -2575 1524 -2549
rect 1774 -2575 2352 -2549
rect 2602 -2549 2686 -2543
rect 2602 -2575 2812 -2549
rect 3064 -2601 3094 -2529
rect 3166 -2555 3266 -2527
rect 3426 -2555 3526 -2527
rect 3571 -2483 3625 -2467
rect 3571 -2517 3581 -2483
rect 3615 -2517 3625 -2483
rect 3571 -2533 3625 -2517
rect 3832 -2493 3974 -2477
rect 3832 -2527 3848 -2493
rect 3882 -2527 3974 -2493
rect 4016 -2491 4108 -2457
rect 4142 -2491 4158 -2457
rect 4016 -2507 4158 -2491
rect 4350 -2457 4614 -2435
rect 4350 -2491 4366 -2457
rect 4400 -2491 4465 -2457
rect 4499 -2491 4564 -2457
rect 4598 -2491 4614 -2457
rect 5304 -2441 5388 -2435
rect 5304 -2457 5446 -2441
rect 4350 -2507 4614 -2491
rect 4656 -2493 4928 -2477
rect 3591 -2601 3621 -2533
rect 3832 -2543 3974 -2527
rect 3890 -2549 3974 -2543
rect 4656 -2527 4672 -2493
rect 4706 -2527 4775 -2493
rect 4809 -2527 4878 -2493
rect 4912 -2527 4928 -2493
rect 4656 -2549 4928 -2527
rect 5120 -2493 5262 -2477
rect 5120 -2527 5136 -2493
rect 5170 -2527 5262 -2493
rect 5304 -2491 5396 -2457
rect 5430 -2491 5446 -2457
rect 5640 -2470 5670 -2435
rect 5304 -2507 5446 -2491
rect 5600 -2483 5670 -2470
rect 5742 -2473 5842 -2399
rect 6002 -2473 6102 -2399
rect 6466 -2435 6676 -2409
rect 6167 -2467 6197 -2435
rect 6592 -2441 6676 -2435
rect 6926 -2435 7504 -2409
rect 7754 -2435 7964 -2409
rect 6592 -2457 6734 -2441
rect 5120 -2543 5262 -2527
rect 5600 -2517 5616 -2483
rect 5650 -2517 5670 -2483
rect 5600 -2529 5670 -2517
rect 5720 -2483 5842 -2473
rect 5720 -2517 5736 -2483
rect 5770 -2517 5842 -2483
rect 5720 -2527 5842 -2517
rect 5941 -2483 6102 -2473
rect 5941 -2517 5957 -2483
rect 5991 -2517 6102 -2483
rect 5941 -2527 6102 -2517
rect 3890 -2575 4100 -2549
rect 4350 -2575 4928 -2549
rect 5178 -2549 5262 -2543
rect 5178 -2575 5388 -2549
rect 5640 -2601 5670 -2529
rect 5742 -2555 5842 -2527
rect 6002 -2555 6102 -2527
rect 6147 -2483 6201 -2467
rect 6147 -2517 6157 -2483
rect 6191 -2517 6201 -2483
rect 6147 -2533 6201 -2517
rect 6408 -2493 6550 -2477
rect 6408 -2527 6424 -2493
rect 6458 -2527 6550 -2493
rect 6592 -2491 6684 -2457
rect 6718 -2491 6734 -2457
rect 6592 -2507 6734 -2491
rect 6926 -2457 7190 -2435
rect 6926 -2491 6942 -2457
rect 6976 -2491 7041 -2457
rect 7075 -2491 7140 -2457
rect 7174 -2491 7190 -2457
rect 7880 -2441 7964 -2435
rect 7880 -2457 8022 -2441
rect 6926 -2507 7190 -2491
rect 7232 -2493 7504 -2477
rect 6167 -2601 6197 -2533
rect 6408 -2543 6550 -2527
rect 6466 -2549 6550 -2543
rect 7232 -2527 7248 -2493
rect 7282 -2527 7351 -2493
rect 7385 -2527 7454 -2493
rect 7488 -2527 7504 -2493
rect 7232 -2549 7504 -2527
rect 7696 -2493 7838 -2477
rect 7696 -2527 7712 -2493
rect 7746 -2527 7838 -2493
rect 7880 -2491 7972 -2457
rect 8006 -2491 8022 -2457
rect 8216 -2470 8246 -2435
rect 7880 -2507 8022 -2491
rect 8176 -2483 8246 -2470
rect 8318 -2473 8418 -2399
rect 8578 -2473 8678 -2399
rect 9042 -2435 9252 -2409
rect 8743 -2467 8773 -2435
rect 9168 -2441 9252 -2435
rect 9502 -2435 10080 -2409
rect 10422 -2435 10632 -2409
rect 9168 -2457 9310 -2441
rect 7696 -2543 7838 -2527
rect 8176 -2517 8192 -2483
rect 8226 -2517 8246 -2483
rect 8176 -2529 8246 -2517
rect 8296 -2483 8418 -2473
rect 8296 -2517 8312 -2483
rect 8346 -2517 8418 -2483
rect 8296 -2527 8418 -2517
rect 8517 -2483 8678 -2473
rect 8517 -2517 8533 -2483
rect 8567 -2517 8678 -2483
rect 8517 -2527 8678 -2517
rect 6466 -2575 6676 -2549
rect 6926 -2575 7504 -2549
rect 7754 -2549 7838 -2543
rect 7754 -2575 7964 -2549
rect 8216 -2601 8246 -2529
rect 8318 -2555 8418 -2527
rect 8578 -2555 8678 -2527
rect 8723 -2483 8777 -2467
rect 8723 -2517 8733 -2483
rect 8767 -2517 8777 -2483
rect 8723 -2533 8777 -2517
rect 8984 -2493 9126 -2477
rect 8984 -2527 9000 -2493
rect 9034 -2527 9126 -2493
rect 9168 -2491 9260 -2457
rect 9294 -2491 9310 -2457
rect 9168 -2507 9310 -2491
rect 9502 -2457 9766 -2435
rect 9502 -2491 9518 -2457
rect 9552 -2491 9617 -2457
rect 9651 -2491 9716 -2457
rect 9750 -2491 9766 -2457
rect 10548 -2441 10632 -2435
rect 10548 -2457 10690 -2441
rect 9502 -2507 9766 -2491
rect 9808 -2493 10080 -2477
rect 8743 -2601 8773 -2533
rect 8984 -2543 9126 -2527
rect 9042 -2549 9126 -2543
rect 9808 -2527 9824 -2493
rect 9858 -2527 9927 -2493
rect 9961 -2527 10030 -2493
rect 10064 -2527 10080 -2493
rect 9808 -2549 10080 -2527
rect 10364 -2493 10506 -2477
rect 10364 -2527 10380 -2493
rect 10414 -2527 10506 -2493
rect 10548 -2491 10640 -2457
rect 10674 -2491 10690 -2457
rect 10792 -2470 10822 -2435
rect 10548 -2507 10690 -2491
rect 10752 -2483 10822 -2470
rect 10894 -2473 10994 -2399
rect 11154 -2473 11254 -2399
rect 11710 -2435 11920 -2409
rect 13274 -2435 13484 -2409
rect 15666 -2435 16612 -2409
rect 11319 -2467 11349 -2435
rect 11836 -2441 11920 -2435
rect 11836 -2457 11978 -2441
rect 10364 -2543 10506 -2527
rect 10752 -2517 10768 -2483
rect 10802 -2517 10822 -2483
rect 10752 -2529 10822 -2517
rect 10872 -2483 10994 -2473
rect 10872 -2517 10888 -2483
rect 10922 -2517 10994 -2483
rect 10872 -2527 10994 -2517
rect 11093 -2483 11254 -2473
rect 11093 -2517 11109 -2483
rect 11143 -2517 11254 -2483
rect 11093 -2527 11254 -2517
rect 9042 -2575 9252 -2549
rect 9502 -2575 10080 -2549
rect 10422 -2549 10506 -2543
rect 10422 -2575 10632 -2549
rect 10792 -2601 10822 -2529
rect 10894 -2555 10994 -2527
rect 11154 -2555 11254 -2527
rect 11299 -2483 11353 -2467
rect 11299 -2517 11309 -2483
rect 11343 -2517 11353 -2483
rect 11299 -2533 11353 -2517
rect 11652 -2493 11794 -2477
rect 11652 -2527 11668 -2493
rect 11702 -2527 11794 -2493
rect 11836 -2491 11928 -2457
rect 11962 -2491 11978 -2457
rect 11836 -2507 11978 -2491
rect 12547 -2473 12577 -2435
rect 12633 -2473 12663 -2435
rect 12719 -2473 12749 -2435
rect 12805 -2473 12835 -2435
rect 12891 -2473 12921 -2435
rect 12977 -2473 13007 -2435
rect 13274 -2441 13358 -2435
rect 12547 -2483 13007 -2473
rect 12547 -2517 12574 -2483
rect 12608 -2517 12642 -2483
rect 12676 -2517 12710 -2483
rect 12744 -2517 12778 -2483
rect 12812 -2517 12846 -2483
rect 12880 -2517 12914 -2483
rect 12948 -2517 13007 -2483
rect 13216 -2457 13358 -2441
rect 13735 -2450 13765 -2435
rect 13821 -2450 13851 -2435
rect 13907 -2450 13937 -2435
rect 13993 -2450 14023 -2435
rect 13216 -2491 13232 -2457
rect 13266 -2491 13358 -2457
rect 13216 -2507 13358 -2491
rect 13400 -2493 13542 -2477
rect 12547 -2527 13007 -2517
rect 13400 -2527 13492 -2493
rect 13526 -2527 13542 -2493
rect 11319 -2601 11349 -2533
rect 11652 -2543 11794 -2527
rect 11710 -2549 11794 -2543
rect 11710 -2575 11920 -2549
rect 12633 -2601 12663 -2527
rect 12719 -2601 12749 -2527
rect 12805 -2601 12835 -2527
rect 12891 -2601 12921 -2527
rect 13400 -2543 13542 -2527
rect 13676 -2483 14023 -2450
rect 13676 -2517 13692 -2483
rect 13726 -2517 14023 -2483
rect 13400 -2549 13484 -2543
rect 13274 -2575 13484 -2549
rect 13676 -2552 14023 -2517
rect 13735 -2601 13765 -2552
rect 13821 -2601 13851 -2552
rect 13907 -2601 13937 -2552
rect 13993 -2601 14023 -2552
rect 14079 -2467 14109 -2435
rect 14165 -2467 14195 -2435
rect 14251 -2467 14281 -2435
rect 14337 -2467 14367 -2435
rect 14423 -2467 14453 -2435
rect 14509 -2467 14539 -2435
rect 14595 -2467 14625 -2435
rect 14681 -2467 14711 -2435
rect 14766 -2467 14796 -2435
rect 14852 -2467 14882 -2435
rect 14938 -2467 14968 -2435
rect 15024 -2467 15054 -2435
rect 15110 -2467 15140 -2435
rect 15196 -2467 15226 -2435
rect 15282 -2467 15312 -2435
rect 15368 -2467 15398 -2435
rect 14079 -2483 15398 -2467
rect 14079 -2517 14119 -2483
rect 14153 -2517 14187 -2483
rect 14221 -2517 14255 -2483
rect 14289 -2517 14323 -2483
rect 14357 -2517 14391 -2483
rect 14425 -2517 14459 -2483
rect 14493 -2517 14527 -2483
rect 14561 -2517 14595 -2483
rect 14629 -2517 14663 -2483
rect 14697 -2517 14731 -2483
rect 14765 -2517 14799 -2483
rect 14833 -2517 14867 -2483
rect 14901 -2517 14935 -2483
rect 14969 -2517 15003 -2483
rect 15037 -2517 15071 -2483
rect 15105 -2517 15139 -2483
rect 15173 -2517 15398 -2483
rect 15666 -2457 16116 -2435
rect 15666 -2491 15682 -2457
rect 15716 -2491 15810 -2457
rect 15844 -2491 15938 -2457
rect 15972 -2491 16066 -2457
rect 16100 -2491 16116 -2457
rect 15666 -2507 16116 -2491
rect 16158 -2493 16612 -2477
rect 14079 -2542 15398 -2517
rect 14079 -2601 14109 -2542
rect 14165 -2601 14195 -2542
rect 14251 -2601 14281 -2542
rect 14337 -2601 14367 -2542
rect 14423 -2601 14453 -2542
rect 14509 -2601 14539 -2542
rect 14595 -2601 14625 -2542
rect 14681 -2601 14711 -2542
rect 14766 -2601 14796 -2542
rect 14852 -2601 14882 -2542
rect 14938 -2601 14968 -2542
rect 15024 -2601 15054 -2542
rect 15110 -2601 15140 -2542
rect 15196 -2601 15226 -2542
rect 15282 -2601 15312 -2542
rect 15368 -2601 15398 -2542
rect 16158 -2527 16174 -2493
rect 16208 -2527 16302 -2493
rect 16336 -2527 16430 -2493
rect 16464 -2527 16558 -2493
rect 16592 -2527 16612 -2493
rect 16158 -2549 16612 -2527
rect 15666 -2575 16612 -2549
rect -2918 -2711 -2340 -2685
rect -1538 -2711 -960 -2685
rect -802 -2711 -224 -2685
rect 26 -2711 236 -2685
rect 488 -2711 518 -2685
rect 590 -2711 690 -2685
rect 850 -2711 950 -2685
rect 1015 -2711 1045 -2685
rect 1314 -2711 1524 -2685
rect 1774 -2711 2352 -2685
rect 2602 -2711 2812 -2685
rect 3064 -2711 3094 -2685
rect 3166 -2711 3266 -2685
rect 3426 -2711 3526 -2685
rect 3591 -2711 3621 -2685
rect 3890 -2711 4100 -2685
rect 4350 -2711 4928 -2685
rect 5178 -2711 5388 -2685
rect 5640 -2711 5670 -2685
rect 5742 -2711 5842 -2685
rect 6002 -2711 6102 -2685
rect 6167 -2711 6197 -2685
rect 6466 -2711 6676 -2685
rect 6926 -2711 7504 -2685
rect 7754 -2711 7964 -2685
rect 8216 -2711 8246 -2685
rect 8318 -2711 8418 -2685
rect 8578 -2711 8678 -2685
rect 8743 -2711 8773 -2685
rect 9042 -2711 9252 -2685
rect 9502 -2711 10080 -2685
rect 10422 -2711 10632 -2685
rect 10792 -2711 10822 -2685
rect 10894 -2711 10994 -2685
rect 11154 -2711 11254 -2685
rect 11319 -2711 11349 -2685
rect 11710 -2711 11920 -2685
rect 12633 -2711 12663 -2685
rect 12719 -2711 12749 -2685
rect 12805 -2711 12835 -2685
rect 12891 -2711 12921 -2685
rect 13274 -2711 13484 -2685
rect 13735 -2711 13765 -2685
rect 13821 -2711 13851 -2685
rect 13907 -2711 13937 -2685
rect 13993 -2711 14023 -2685
rect 14079 -2711 14109 -2685
rect 14165 -2711 14195 -2685
rect 14251 -2711 14281 -2685
rect 14337 -2711 14367 -2685
rect 14423 -2711 14453 -2685
rect 14509 -2711 14539 -2685
rect 14595 -2711 14625 -2685
rect 14681 -2711 14711 -2685
rect 14766 -2711 14796 -2685
rect 14852 -2711 14882 -2685
rect 14938 -2711 14968 -2685
rect 15024 -2711 15054 -2685
rect 15110 -2711 15140 -2685
rect 15196 -2711 15226 -2685
rect 15282 -2711 15312 -2685
rect 15368 -2711 15398 -2685
rect 15666 -2711 16612 -2685
rect -2918 -2779 -2340 -2753
rect -1823 -2779 -1793 -2753
rect -1538 -2779 -960 -2753
rect -802 -2779 -224 -2753
rect 26 -2779 236 -2753
rect 505 -2779 535 -2753
rect 600 -2779 700 -2753
rect 860 -2779 960 -2753
rect 1032 -2779 1062 -2753
rect 1314 -2779 1524 -2753
rect 1774 -2779 2352 -2753
rect 2602 -2779 2812 -2753
rect 3081 -2779 3111 -2753
rect 3176 -2779 3276 -2753
rect 3436 -2779 3536 -2753
rect 3608 -2779 3638 -2753
rect 3890 -2779 4100 -2753
rect 4350 -2779 4928 -2753
rect 5178 -2779 5388 -2753
rect 5657 -2779 5687 -2753
rect 5752 -2779 5852 -2753
rect 6012 -2779 6112 -2753
rect 6184 -2779 6214 -2753
rect 6466 -2779 6676 -2753
rect 6926 -2779 7504 -2753
rect 7754 -2779 7964 -2753
rect 8233 -2779 8263 -2753
rect 8328 -2779 8428 -2753
rect 8588 -2779 8688 -2753
rect 8760 -2779 8790 -2753
rect 9042 -2779 9252 -2753
rect 9502 -2779 10080 -2753
rect 10422 -2779 10632 -2753
rect 10809 -2779 10839 -2753
rect 10904 -2779 11004 -2753
rect 11164 -2779 11264 -2753
rect 11336 -2779 11366 -2753
rect 11710 -2779 11920 -2753
rect 13642 -2779 14588 -2753
rect 14838 -2779 15784 -2753
rect 16034 -2779 16612 -2753
rect -2918 -2915 -2340 -2889
rect -2918 -2937 -2646 -2915
rect -1823 -2927 -1793 -2863
rect -1907 -2931 -1793 -2927
rect -2918 -2971 -2902 -2937
rect -2868 -2971 -2799 -2937
rect -2765 -2971 -2696 -2937
rect -2662 -2971 -2646 -2937
rect -1964 -2947 -1793 -2931
rect -2918 -2987 -2646 -2971
rect -2604 -2973 -2340 -2957
rect -2604 -3007 -2588 -2973
rect -2554 -3007 -2489 -2973
rect -2455 -3007 -2390 -2973
rect -2356 -3007 -2340 -2973
rect -1964 -2981 -1954 -2947
rect -1920 -2971 -1793 -2947
rect -1538 -2915 -960 -2889
rect -802 -2915 -224 -2889
rect 26 -2915 236 -2889
rect -1538 -2937 -1266 -2915
rect -1538 -2971 -1522 -2937
rect -1488 -2971 -1419 -2937
rect -1385 -2971 -1316 -2937
rect -1282 -2971 -1266 -2937
rect -802 -2937 -530 -2915
rect 26 -2921 110 -2915
rect -1920 -2981 -1792 -2971
rect -1964 -2997 -1792 -2981
rect -1538 -2987 -1266 -2971
rect -1224 -2973 -960 -2957
rect -2604 -3029 -2340 -3007
rect -2918 -3055 -2340 -3029
rect -1906 -3001 -1792 -2997
rect -1906 -3061 -1876 -3001
rect -1822 -3061 -1792 -3001
rect -1224 -3007 -1208 -2973
rect -1174 -3007 -1109 -2973
rect -1075 -3007 -1010 -2973
rect -976 -3007 -960 -2973
rect -802 -2971 -786 -2937
rect -752 -2971 -683 -2937
rect -649 -2971 -580 -2937
rect -546 -2971 -530 -2937
rect -32 -2937 110 -2921
rect 505 -2931 535 -2863
rect -802 -2987 -530 -2971
rect -488 -2973 -224 -2957
rect -1224 -3029 -960 -3007
rect -488 -3007 -472 -2973
rect -438 -3007 -373 -2973
rect -339 -3007 -274 -2973
rect -240 -3007 -224 -2973
rect -32 -2971 -16 -2937
rect 18 -2971 110 -2937
rect 501 -2947 555 -2931
rect -32 -2987 110 -2971
rect 152 -2973 294 -2957
rect -488 -3029 -224 -3007
rect 152 -3007 244 -2973
rect 278 -3007 294 -2973
rect 501 -2981 511 -2947
rect 545 -2981 555 -2947
rect 501 -2997 555 -2981
rect 600 -2937 700 -2909
rect 860 -2937 960 -2909
rect 1032 -2935 1062 -2863
rect 1314 -2915 1524 -2889
rect 1774 -2915 2352 -2889
rect 2602 -2915 2812 -2889
rect 1314 -2921 1398 -2915
rect 600 -2947 761 -2937
rect 600 -2981 711 -2947
rect 745 -2981 761 -2947
rect 600 -2991 761 -2981
rect 860 -2947 982 -2937
rect 860 -2981 932 -2947
rect 966 -2981 982 -2947
rect 860 -2991 982 -2981
rect 1032 -2947 1102 -2935
rect 1032 -2981 1052 -2947
rect 1086 -2981 1102 -2947
rect 152 -3023 294 -3007
rect 152 -3029 236 -3023
rect 505 -3029 535 -2997
rect -1538 -3055 -960 -3029
rect -802 -3055 -224 -3029
rect 26 -3055 236 -3029
rect 600 -3065 700 -2991
rect 860 -3065 960 -2991
rect 1032 -2994 1102 -2981
rect 1256 -2937 1398 -2921
rect 1256 -2971 1272 -2937
rect 1306 -2971 1398 -2937
rect 1774 -2937 2046 -2915
rect 2602 -2921 2686 -2915
rect 1256 -2987 1398 -2971
rect 1440 -2973 1582 -2957
rect 1032 -3029 1062 -2994
rect 1440 -3007 1532 -2973
rect 1566 -3007 1582 -2973
rect 1774 -2971 1790 -2937
rect 1824 -2971 1893 -2937
rect 1927 -2971 1996 -2937
rect 2030 -2971 2046 -2937
rect 2544 -2937 2686 -2921
rect 3081 -2931 3111 -2863
rect 1774 -2987 2046 -2971
rect 2088 -2973 2352 -2957
rect 1440 -3023 1582 -3007
rect 2088 -3007 2104 -2973
rect 2138 -3007 2203 -2973
rect 2237 -3007 2302 -2973
rect 2336 -3007 2352 -2973
rect 2544 -2971 2560 -2937
rect 2594 -2971 2686 -2937
rect 3077 -2947 3131 -2931
rect 2544 -2987 2686 -2971
rect 2728 -2973 2870 -2957
rect 1440 -3029 1524 -3023
rect 2088 -3029 2352 -3007
rect 2728 -3007 2820 -2973
rect 2854 -3007 2870 -2973
rect 3077 -2981 3087 -2947
rect 3121 -2981 3131 -2947
rect 3077 -2997 3131 -2981
rect 3176 -2937 3276 -2909
rect 3436 -2937 3536 -2909
rect 3608 -2935 3638 -2863
rect 3890 -2915 4100 -2889
rect 4350 -2915 4928 -2889
rect 5178 -2915 5388 -2889
rect 3890 -2921 3974 -2915
rect 3176 -2947 3337 -2937
rect 3176 -2981 3287 -2947
rect 3321 -2981 3337 -2947
rect 3176 -2991 3337 -2981
rect 3436 -2947 3558 -2937
rect 3436 -2981 3508 -2947
rect 3542 -2981 3558 -2947
rect 3436 -2991 3558 -2981
rect 3608 -2947 3678 -2935
rect 3608 -2981 3628 -2947
rect 3662 -2981 3678 -2947
rect 2728 -3023 2870 -3007
rect 2728 -3029 2812 -3023
rect 3081 -3029 3111 -2997
rect 1314 -3055 1524 -3029
rect 1774 -3055 2352 -3029
rect 2602 -3055 2812 -3029
rect 3176 -3065 3276 -2991
rect 3436 -3065 3536 -2991
rect 3608 -2994 3678 -2981
rect 3832 -2937 3974 -2921
rect 3832 -2971 3848 -2937
rect 3882 -2971 3974 -2937
rect 4350 -2937 4622 -2915
rect 5178 -2921 5262 -2915
rect 3832 -2987 3974 -2971
rect 4016 -2973 4158 -2957
rect 3608 -3029 3638 -2994
rect 4016 -3007 4108 -2973
rect 4142 -3007 4158 -2973
rect 4350 -2971 4366 -2937
rect 4400 -2971 4469 -2937
rect 4503 -2971 4572 -2937
rect 4606 -2971 4622 -2937
rect 5120 -2937 5262 -2921
rect 5657 -2931 5687 -2863
rect 4350 -2987 4622 -2971
rect 4664 -2973 4928 -2957
rect 4016 -3023 4158 -3007
rect 4664 -3007 4680 -2973
rect 4714 -3007 4779 -2973
rect 4813 -3007 4878 -2973
rect 4912 -3007 4928 -2973
rect 5120 -2971 5136 -2937
rect 5170 -2971 5262 -2937
rect 5653 -2947 5707 -2931
rect 5120 -2987 5262 -2971
rect 5304 -2973 5446 -2957
rect 4016 -3029 4100 -3023
rect 4664 -3029 4928 -3007
rect 5304 -3007 5396 -2973
rect 5430 -3007 5446 -2973
rect 5653 -2981 5663 -2947
rect 5697 -2981 5707 -2947
rect 5653 -2997 5707 -2981
rect 5752 -2937 5852 -2909
rect 6012 -2937 6112 -2909
rect 6184 -2935 6214 -2863
rect 6466 -2915 6676 -2889
rect 6926 -2915 7504 -2889
rect 7754 -2915 7964 -2889
rect 6466 -2921 6550 -2915
rect 5752 -2947 5913 -2937
rect 5752 -2981 5863 -2947
rect 5897 -2981 5913 -2947
rect 5752 -2991 5913 -2981
rect 6012 -2947 6134 -2937
rect 6012 -2981 6084 -2947
rect 6118 -2981 6134 -2947
rect 6012 -2991 6134 -2981
rect 6184 -2947 6254 -2935
rect 6184 -2981 6204 -2947
rect 6238 -2981 6254 -2947
rect 5304 -3023 5446 -3007
rect 5304 -3029 5388 -3023
rect 5657 -3029 5687 -2997
rect 3890 -3055 4100 -3029
rect 4350 -3055 4928 -3029
rect 5178 -3055 5388 -3029
rect 5752 -3065 5852 -2991
rect 6012 -3065 6112 -2991
rect 6184 -2994 6254 -2981
rect 6408 -2937 6550 -2921
rect 6408 -2971 6424 -2937
rect 6458 -2971 6550 -2937
rect 6926 -2937 7198 -2915
rect 7754 -2921 7838 -2915
rect 6408 -2987 6550 -2971
rect 6592 -2973 6734 -2957
rect 6184 -3029 6214 -2994
rect 6592 -3007 6684 -2973
rect 6718 -3007 6734 -2973
rect 6926 -2971 6942 -2937
rect 6976 -2971 7045 -2937
rect 7079 -2971 7148 -2937
rect 7182 -2971 7198 -2937
rect 7696 -2937 7838 -2921
rect 8233 -2931 8263 -2863
rect 6926 -2987 7198 -2971
rect 7240 -2973 7504 -2957
rect 6592 -3023 6734 -3007
rect 7240 -3007 7256 -2973
rect 7290 -3007 7355 -2973
rect 7389 -3007 7454 -2973
rect 7488 -3007 7504 -2973
rect 7696 -2971 7712 -2937
rect 7746 -2971 7838 -2937
rect 8229 -2947 8283 -2931
rect 7696 -2987 7838 -2971
rect 7880 -2973 8022 -2957
rect 6592 -3029 6676 -3023
rect 7240 -3029 7504 -3007
rect 7880 -3007 7972 -2973
rect 8006 -3007 8022 -2973
rect 8229 -2981 8239 -2947
rect 8273 -2981 8283 -2947
rect 8229 -2997 8283 -2981
rect 8328 -2937 8428 -2909
rect 8588 -2937 8688 -2909
rect 8760 -2935 8790 -2863
rect 9042 -2915 9252 -2889
rect 9502 -2915 10080 -2889
rect 10422 -2915 10632 -2889
rect 9042 -2921 9126 -2915
rect 8328 -2947 8489 -2937
rect 8328 -2981 8439 -2947
rect 8473 -2981 8489 -2947
rect 8328 -2991 8489 -2981
rect 8588 -2947 8710 -2937
rect 8588 -2981 8660 -2947
rect 8694 -2981 8710 -2947
rect 8588 -2991 8710 -2981
rect 8760 -2947 8830 -2935
rect 8760 -2981 8780 -2947
rect 8814 -2981 8830 -2947
rect 7880 -3023 8022 -3007
rect 7880 -3029 7964 -3023
rect 8233 -3029 8263 -2997
rect 6466 -3055 6676 -3029
rect 6926 -3055 7504 -3029
rect 7754 -3055 7964 -3029
rect 8328 -3065 8428 -2991
rect 8588 -3065 8688 -2991
rect 8760 -2994 8830 -2981
rect 8984 -2937 9126 -2921
rect 8984 -2971 9000 -2937
rect 9034 -2971 9126 -2937
rect 9502 -2937 9774 -2915
rect 10422 -2921 10506 -2915
rect 8984 -2987 9126 -2971
rect 9168 -2973 9310 -2957
rect 8760 -3029 8790 -2994
rect 9168 -3007 9260 -2973
rect 9294 -3007 9310 -2973
rect 9502 -2971 9518 -2937
rect 9552 -2971 9621 -2937
rect 9655 -2971 9724 -2937
rect 9758 -2971 9774 -2937
rect 10364 -2937 10506 -2921
rect 10809 -2931 10839 -2863
rect 9502 -2987 9774 -2971
rect 9816 -2973 10080 -2957
rect 9168 -3023 9310 -3007
rect 9816 -3007 9832 -2973
rect 9866 -3007 9931 -2973
rect 9965 -3007 10030 -2973
rect 10064 -3007 10080 -2973
rect 10364 -2971 10380 -2937
rect 10414 -2971 10506 -2937
rect 10805 -2947 10859 -2931
rect 10364 -2987 10506 -2971
rect 10548 -2973 10690 -2957
rect 9168 -3029 9252 -3023
rect 9816 -3029 10080 -3007
rect 10548 -3007 10640 -2973
rect 10674 -3007 10690 -2973
rect 10805 -2981 10815 -2947
rect 10849 -2981 10859 -2947
rect 10805 -2997 10859 -2981
rect 10904 -2937 11004 -2909
rect 11164 -2937 11264 -2909
rect 11336 -2935 11366 -2863
rect 11710 -2915 11920 -2889
rect 13642 -2915 14588 -2889
rect 14838 -2915 15784 -2889
rect 16034 -2915 16612 -2889
rect 11710 -2921 11794 -2915
rect 10904 -2947 11065 -2937
rect 10904 -2981 11015 -2947
rect 11049 -2981 11065 -2947
rect 10904 -2991 11065 -2981
rect 11164 -2947 11286 -2937
rect 11164 -2981 11236 -2947
rect 11270 -2981 11286 -2947
rect 11164 -2991 11286 -2981
rect 11336 -2947 11406 -2935
rect 11336 -2981 11356 -2947
rect 11390 -2981 11406 -2947
rect 10548 -3023 10690 -3007
rect 10548 -3029 10632 -3023
rect 10809 -3029 10839 -2997
rect 9042 -3055 9252 -3029
rect 9502 -3055 10080 -3029
rect 10422 -3055 10632 -3029
rect 10904 -3065 11004 -2991
rect 11164 -3065 11264 -2991
rect 11336 -2994 11406 -2981
rect 11652 -2937 11794 -2921
rect 11652 -2971 11668 -2937
rect 11702 -2971 11794 -2937
rect 13642 -2937 14096 -2915
rect 11652 -2987 11794 -2971
rect 11836 -2973 11978 -2957
rect 11336 -3029 11366 -2994
rect 11836 -3007 11928 -2973
rect 11962 -3007 11978 -2973
rect 13642 -2971 13662 -2937
rect 13696 -2971 13790 -2937
rect 13824 -2971 13918 -2937
rect 13952 -2971 14046 -2937
rect 14080 -2971 14096 -2937
rect 14838 -2937 15292 -2915
rect 13642 -2987 14096 -2971
rect 14138 -2973 14588 -2957
rect 11836 -3023 11978 -3007
rect 14138 -3007 14154 -2973
rect 14188 -3007 14282 -2973
rect 14316 -3007 14410 -2973
rect 14444 -3007 14538 -2973
rect 14572 -3007 14588 -2973
rect 14838 -2971 14858 -2937
rect 14892 -2971 14986 -2937
rect 15020 -2971 15114 -2937
rect 15148 -2971 15242 -2937
rect 15276 -2971 15292 -2937
rect 16034 -2937 16306 -2915
rect 14838 -2987 15292 -2971
rect 15334 -2973 15784 -2957
rect 11836 -3029 11920 -3023
rect 14138 -3029 14588 -3007
rect 15334 -3007 15350 -2973
rect 15384 -3007 15478 -2973
rect 15512 -3007 15606 -2973
rect 15640 -3007 15734 -2973
rect 15768 -3007 15784 -2973
rect 16034 -2971 16050 -2937
rect 16084 -2971 16153 -2937
rect 16187 -2971 16256 -2937
rect 16290 -2971 16306 -2937
rect 16034 -2987 16306 -2971
rect 16348 -2973 16612 -2957
rect 15334 -3029 15784 -3007
rect 16348 -3007 16364 -2973
rect 16398 -3007 16463 -2973
rect 16497 -3007 16562 -2973
rect 16596 -3007 16612 -2973
rect 16348 -3029 16612 -3007
rect 11710 -3055 11920 -3029
rect 13642 -3055 14588 -3029
rect 14838 -3055 15784 -3029
rect 16034 -3055 16612 -3029
rect -2918 -3255 -2340 -3229
rect -1906 -3255 -1876 -3229
rect -1822 -3255 -1792 -3229
rect -1538 -3255 -960 -3229
rect -802 -3255 -224 -3229
rect 26 -3255 236 -3229
rect 505 -3255 535 -3229
rect 600 -3255 700 -3229
rect 860 -3255 960 -3229
rect 1032 -3255 1062 -3229
rect 1314 -3255 1524 -3229
rect 1774 -3255 2352 -3229
rect 2602 -3255 2812 -3229
rect 3081 -3255 3111 -3229
rect 3176 -3255 3276 -3229
rect 3436 -3255 3536 -3229
rect 3608 -3255 3638 -3229
rect 3890 -3255 4100 -3229
rect 4350 -3255 4928 -3229
rect 5178 -3255 5388 -3229
rect 5657 -3255 5687 -3229
rect 5752 -3255 5852 -3229
rect 6012 -3255 6112 -3229
rect 6184 -3255 6214 -3229
rect 6466 -3255 6676 -3229
rect 6926 -3255 7504 -3229
rect 7754 -3255 7964 -3229
rect 8233 -3255 8263 -3229
rect 8328 -3255 8428 -3229
rect 8588 -3255 8688 -3229
rect 8760 -3255 8790 -3229
rect 9042 -3255 9252 -3229
rect 9502 -3255 10080 -3229
rect 10422 -3255 10632 -3229
rect 10809 -3255 10839 -3229
rect 10904 -3255 11004 -3229
rect 11164 -3255 11264 -3229
rect 11336 -3255 11366 -3229
rect 11710 -3255 11920 -3229
rect 13642 -3255 14588 -3229
rect 14838 -3255 15784 -3229
rect 16034 -3255 16612 -3229
rect -2918 -3323 -2340 -3297
rect -1538 -3323 -960 -3297
rect -802 -3323 -224 -3297
rect 26 -3323 236 -3297
rect 505 -3323 535 -3297
rect 600 -3323 700 -3297
rect 860 -3323 960 -3297
rect 1032 -3323 1062 -3297
rect 1314 -3323 1524 -3297
rect 1774 -3323 2352 -3297
rect 2602 -3323 2812 -3297
rect 3081 -3323 3111 -3297
rect 3176 -3323 3276 -3297
rect 3436 -3323 3536 -3297
rect 3608 -3323 3638 -3297
rect 3890 -3323 4100 -3297
rect 4350 -3323 4928 -3297
rect 5178 -3323 5388 -3297
rect 5657 -3323 5687 -3297
rect 5752 -3323 5852 -3297
rect 6012 -3323 6112 -3297
rect 6184 -3323 6214 -3297
rect 6466 -3323 6676 -3297
rect 6926 -3323 7504 -3297
rect 7754 -3323 7964 -3297
rect 8233 -3323 8263 -3297
rect 8328 -3323 8428 -3297
rect 8588 -3323 8688 -3297
rect 8760 -3323 8790 -3297
rect 9042 -3323 9252 -3297
rect 9502 -3323 10080 -3297
rect 10422 -3323 10632 -3297
rect 10809 -3323 10839 -3297
rect 10904 -3323 11004 -3297
rect 11164 -3323 11264 -3297
rect 11336 -3323 11366 -3297
rect 11710 -3323 11920 -3297
rect 13642 -3323 14588 -3297
rect 14838 -3323 15784 -3297
rect 16034 -3323 16612 -3297
rect -2918 -3523 -2340 -3497
rect -1538 -3523 -960 -3497
rect -802 -3523 -224 -3497
rect 26 -3523 236 -3497
rect -2918 -3545 -2654 -3523
rect -2918 -3579 -2902 -3545
rect -2868 -3579 -2803 -3545
rect -2769 -3579 -2704 -3545
rect -2670 -3579 -2654 -3545
rect -1224 -3545 -960 -3523
rect -2918 -3595 -2654 -3579
rect -2612 -3581 -2340 -3565
rect -2612 -3615 -2596 -3581
rect -2562 -3615 -2493 -3581
rect -2459 -3615 -2390 -3581
rect -2356 -3615 -2340 -3581
rect -2612 -3637 -2340 -3615
rect -2918 -3663 -2340 -3637
rect -1538 -3581 -1266 -3565
rect -1538 -3615 -1522 -3581
rect -1488 -3615 -1419 -3581
rect -1385 -3615 -1316 -3581
rect -1282 -3615 -1266 -3581
rect -1224 -3579 -1208 -3545
rect -1174 -3579 -1109 -3545
rect -1075 -3579 -1010 -3545
rect -976 -3579 -960 -3545
rect -488 -3545 -224 -3523
rect -1224 -3595 -960 -3579
rect -802 -3581 -530 -3565
rect -1538 -3637 -1266 -3615
rect -802 -3615 -786 -3581
rect -752 -3615 -683 -3581
rect -649 -3615 -580 -3581
rect -546 -3615 -530 -3581
rect -488 -3579 -472 -3545
rect -438 -3579 -373 -3545
rect -339 -3579 -274 -3545
rect -240 -3579 -224 -3545
rect 152 -3529 236 -3523
rect 152 -3545 294 -3529
rect -488 -3595 -224 -3579
rect -32 -3581 110 -3565
rect -802 -3637 -530 -3615
rect -32 -3615 -16 -3581
rect 18 -3615 110 -3581
rect 152 -3579 244 -3545
rect 278 -3579 294 -3545
rect 505 -3555 535 -3523
rect 152 -3595 294 -3579
rect 501 -3571 555 -3555
rect -32 -3631 110 -3615
rect 501 -3605 511 -3571
rect 545 -3605 555 -3571
rect 501 -3621 555 -3605
rect 600 -3561 700 -3487
rect 860 -3561 960 -3487
rect 1314 -3523 1524 -3497
rect 1032 -3558 1062 -3523
rect 1440 -3529 1524 -3523
rect 1774 -3523 2352 -3497
rect 2602 -3523 2812 -3497
rect 1440 -3545 1582 -3529
rect 600 -3571 761 -3561
rect 600 -3605 711 -3571
rect 745 -3605 761 -3571
rect 600 -3615 761 -3605
rect 860 -3571 982 -3561
rect 860 -3605 932 -3571
rect 966 -3605 982 -3571
rect 860 -3615 982 -3605
rect 1032 -3571 1102 -3558
rect 1032 -3605 1052 -3571
rect 1086 -3605 1102 -3571
rect 26 -3637 110 -3631
rect -1538 -3663 -960 -3637
rect -802 -3663 -224 -3637
rect 26 -3663 236 -3637
rect 505 -3689 535 -3621
rect 600 -3643 700 -3615
rect 860 -3643 960 -3615
rect 1032 -3617 1102 -3605
rect 1256 -3581 1398 -3565
rect 1256 -3615 1272 -3581
rect 1306 -3615 1398 -3581
rect 1440 -3579 1532 -3545
rect 1566 -3579 1582 -3545
rect 1440 -3595 1582 -3579
rect 1774 -3545 2038 -3523
rect 1774 -3579 1790 -3545
rect 1824 -3579 1889 -3545
rect 1923 -3579 1988 -3545
rect 2022 -3579 2038 -3545
rect 2728 -3529 2812 -3523
rect 2728 -3545 2870 -3529
rect 1774 -3595 2038 -3579
rect 2080 -3581 2352 -3565
rect 1032 -3689 1062 -3617
rect 1256 -3631 1398 -3615
rect 1314 -3637 1398 -3631
rect 2080 -3615 2096 -3581
rect 2130 -3615 2199 -3581
rect 2233 -3615 2302 -3581
rect 2336 -3615 2352 -3581
rect 2080 -3637 2352 -3615
rect 2544 -3581 2686 -3565
rect 2544 -3615 2560 -3581
rect 2594 -3615 2686 -3581
rect 2728 -3579 2820 -3545
rect 2854 -3579 2870 -3545
rect 3081 -3555 3111 -3523
rect 2728 -3595 2870 -3579
rect 3077 -3571 3131 -3555
rect 2544 -3631 2686 -3615
rect 3077 -3605 3087 -3571
rect 3121 -3605 3131 -3571
rect 3077 -3621 3131 -3605
rect 3176 -3561 3276 -3487
rect 3436 -3561 3536 -3487
rect 3890 -3523 4100 -3497
rect 3608 -3558 3638 -3523
rect 4016 -3529 4100 -3523
rect 4350 -3523 4928 -3497
rect 5178 -3523 5388 -3497
rect 4016 -3545 4158 -3529
rect 3176 -3571 3337 -3561
rect 3176 -3605 3287 -3571
rect 3321 -3605 3337 -3571
rect 3176 -3615 3337 -3605
rect 3436 -3571 3558 -3561
rect 3436 -3605 3508 -3571
rect 3542 -3605 3558 -3571
rect 3436 -3615 3558 -3605
rect 3608 -3571 3678 -3558
rect 3608 -3605 3628 -3571
rect 3662 -3605 3678 -3571
rect 1314 -3663 1524 -3637
rect 1774 -3663 2352 -3637
rect 2602 -3637 2686 -3631
rect 2602 -3663 2812 -3637
rect 3081 -3689 3111 -3621
rect 3176 -3643 3276 -3615
rect 3436 -3643 3536 -3615
rect 3608 -3617 3678 -3605
rect 3832 -3581 3974 -3565
rect 3832 -3615 3848 -3581
rect 3882 -3615 3974 -3581
rect 4016 -3579 4108 -3545
rect 4142 -3579 4158 -3545
rect 4016 -3595 4158 -3579
rect 4350 -3545 4614 -3523
rect 4350 -3579 4366 -3545
rect 4400 -3579 4465 -3545
rect 4499 -3579 4564 -3545
rect 4598 -3579 4614 -3545
rect 5304 -3529 5388 -3523
rect 5304 -3545 5446 -3529
rect 4350 -3595 4614 -3579
rect 4656 -3581 4928 -3565
rect 3608 -3689 3638 -3617
rect 3832 -3631 3974 -3615
rect 3890 -3637 3974 -3631
rect 4656 -3615 4672 -3581
rect 4706 -3615 4775 -3581
rect 4809 -3615 4878 -3581
rect 4912 -3615 4928 -3581
rect 4656 -3637 4928 -3615
rect 5120 -3581 5262 -3565
rect 5120 -3615 5136 -3581
rect 5170 -3615 5262 -3581
rect 5304 -3579 5396 -3545
rect 5430 -3579 5446 -3545
rect 5657 -3555 5687 -3523
rect 5304 -3595 5446 -3579
rect 5653 -3571 5707 -3555
rect 5120 -3631 5262 -3615
rect 5653 -3605 5663 -3571
rect 5697 -3605 5707 -3571
rect 5653 -3621 5707 -3605
rect 5752 -3561 5852 -3487
rect 6012 -3561 6112 -3487
rect 6466 -3523 6676 -3497
rect 6184 -3558 6214 -3523
rect 6592 -3529 6676 -3523
rect 6926 -3523 7504 -3497
rect 7754 -3523 7964 -3497
rect 6592 -3545 6734 -3529
rect 5752 -3571 5913 -3561
rect 5752 -3605 5863 -3571
rect 5897 -3605 5913 -3571
rect 5752 -3615 5913 -3605
rect 6012 -3571 6134 -3561
rect 6012 -3605 6084 -3571
rect 6118 -3605 6134 -3571
rect 6012 -3615 6134 -3605
rect 6184 -3571 6254 -3558
rect 6184 -3605 6204 -3571
rect 6238 -3605 6254 -3571
rect 3890 -3663 4100 -3637
rect 4350 -3663 4928 -3637
rect 5178 -3637 5262 -3631
rect 5178 -3663 5388 -3637
rect 5657 -3689 5687 -3621
rect 5752 -3643 5852 -3615
rect 6012 -3643 6112 -3615
rect 6184 -3617 6254 -3605
rect 6408 -3581 6550 -3565
rect 6408 -3615 6424 -3581
rect 6458 -3615 6550 -3581
rect 6592 -3579 6684 -3545
rect 6718 -3579 6734 -3545
rect 6592 -3595 6734 -3579
rect 6926 -3545 7190 -3523
rect 6926 -3579 6942 -3545
rect 6976 -3579 7041 -3545
rect 7075 -3579 7140 -3545
rect 7174 -3579 7190 -3545
rect 7880 -3529 7964 -3523
rect 7880 -3545 8022 -3529
rect 6926 -3595 7190 -3579
rect 7232 -3581 7504 -3565
rect 6184 -3689 6214 -3617
rect 6408 -3631 6550 -3615
rect 6466 -3637 6550 -3631
rect 7232 -3615 7248 -3581
rect 7282 -3615 7351 -3581
rect 7385 -3615 7454 -3581
rect 7488 -3615 7504 -3581
rect 7232 -3637 7504 -3615
rect 7696 -3581 7838 -3565
rect 7696 -3615 7712 -3581
rect 7746 -3615 7838 -3581
rect 7880 -3579 7972 -3545
rect 8006 -3579 8022 -3545
rect 8233 -3555 8263 -3523
rect 7880 -3595 8022 -3579
rect 8229 -3571 8283 -3555
rect 7696 -3631 7838 -3615
rect 8229 -3605 8239 -3571
rect 8273 -3605 8283 -3571
rect 8229 -3621 8283 -3605
rect 8328 -3561 8428 -3487
rect 8588 -3561 8688 -3487
rect 9042 -3523 9252 -3497
rect 8760 -3558 8790 -3523
rect 9168 -3529 9252 -3523
rect 9502 -3523 10080 -3497
rect 10422 -3523 10632 -3497
rect 9168 -3545 9310 -3529
rect 8328 -3571 8489 -3561
rect 8328 -3605 8439 -3571
rect 8473 -3605 8489 -3571
rect 8328 -3615 8489 -3605
rect 8588 -3571 8710 -3561
rect 8588 -3605 8660 -3571
rect 8694 -3605 8710 -3571
rect 8588 -3615 8710 -3605
rect 8760 -3571 8830 -3558
rect 8760 -3605 8780 -3571
rect 8814 -3605 8830 -3571
rect 6466 -3663 6676 -3637
rect 6926 -3663 7504 -3637
rect 7754 -3637 7838 -3631
rect 7754 -3663 7964 -3637
rect 8233 -3689 8263 -3621
rect 8328 -3643 8428 -3615
rect 8588 -3643 8688 -3615
rect 8760 -3617 8830 -3605
rect 8984 -3581 9126 -3565
rect 8984 -3615 9000 -3581
rect 9034 -3615 9126 -3581
rect 9168 -3579 9260 -3545
rect 9294 -3579 9310 -3545
rect 9168 -3595 9310 -3579
rect 9502 -3545 9766 -3523
rect 9502 -3579 9518 -3545
rect 9552 -3579 9617 -3545
rect 9651 -3579 9716 -3545
rect 9750 -3579 9766 -3545
rect 10548 -3529 10632 -3523
rect 10548 -3545 10690 -3529
rect 9502 -3595 9766 -3579
rect 9808 -3581 10080 -3565
rect 8760 -3689 8790 -3617
rect 8984 -3631 9126 -3615
rect 9042 -3637 9126 -3631
rect 9808 -3615 9824 -3581
rect 9858 -3615 9927 -3581
rect 9961 -3615 10030 -3581
rect 10064 -3615 10080 -3581
rect 9808 -3637 10080 -3615
rect 10364 -3581 10506 -3565
rect 10364 -3615 10380 -3581
rect 10414 -3615 10506 -3581
rect 10548 -3579 10640 -3545
rect 10674 -3579 10690 -3545
rect 10809 -3555 10839 -3523
rect 10548 -3595 10690 -3579
rect 10805 -3571 10859 -3555
rect 10364 -3631 10506 -3615
rect 10805 -3605 10815 -3571
rect 10849 -3605 10859 -3571
rect 10805 -3621 10859 -3605
rect 10904 -3561 11004 -3487
rect 11164 -3561 11264 -3487
rect 11710 -3523 11920 -3497
rect 13642 -3523 14588 -3497
rect 14838 -3523 15784 -3497
rect 16034 -3523 16612 -3497
rect 11336 -3558 11366 -3523
rect 11836 -3529 11920 -3523
rect 11836 -3545 11978 -3529
rect 10904 -3571 11065 -3561
rect 10904 -3605 11015 -3571
rect 11049 -3605 11065 -3571
rect 10904 -3615 11065 -3605
rect 11164 -3571 11286 -3561
rect 11164 -3605 11236 -3571
rect 11270 -3605 11286 -3571
rect 11164 -3615 11286 -3605
rect 11336 -3571 11406 -3558
rect 11336 -3605 11356 -3571
rect 11390 -3605 11406 -3571
rect 9042 -3663 9252 -3637
rect 9502 -3663 10080 -3637
rect 10422 -3637 10506 -3631
rect 10422 -3663 10632 -3637
rect 10809 -3689 10839 -3621
rect 10904 -3643 11004 -3615
rect 11164 -3643 11264 -3615
rect 11336 -3617 11406 -3605
rect 11652 -3581 11794 -3565
rect 11652 -3615 11668 -3581
rect 11702 -3615 11794 -3581
rect 11836 -3579 11928 -3545
rect 11962 -3579 11978 -3545
rect 14138 -3545 14588 -3523
rect 11836 -3595 11978 -3579
rect 13642 -3581 14096 -3565
rect 11336 -3689 11366 -3617
rect 11652 -3631 11794 -3615
rect 11710 -3637 11794 -3631
rect 13642 -3615 13662 -3581
rect 13696 -3615 13790 -3581
rect 13824 -3615 13918 -3581
rect 13952 -3615 14046 -3581
rect 14080 -3615 14096 -3581
rect 14138 -3579 14154 -3545
rect 14188 -3579 14282 -3545
rect 14316 -3579 14410 -3545
rect 14444 -3579 14538 -3545
rect 14572 -3579 14588 -3545
rect 15334 -3545 15784 -3523
rect 14138 -3595 14588 -3579
rect 14838 -3581 15292 -3565
rect 13642 -3637 14096 -3615
rect 14838 -3615 14858 -3581
rect 14892 -3615 14986 -3581
rect 15020 -3615 15114 -3581
rect 15148 -3615 15242 -3581
rect 15276 -3615 15292 -3581
rect 15334 -3579 15350 -3545
rect 15384 -3579 15478 -3545
rect 15512 -3579 15606 -3545
rect 15640 -3579 15734 -3545
rect 15768 -3579 15784 -3545
rect 16348 -3545 16612 -3523
rect 15334 -3595 15784 -3579
rect 16034 -3581 16306 -3565
rect 14838 -3637 15292 -3615
rect 16034 -3615 16050 -3581
rect 16084 -3615 16153 -3581
rect 16187 -3615 16256 -3581
rect 16290 -3615 16306 -3581
rect 16348 -3579 16364 -3545
rect 16398 -3579 16463 -3545
rect 16497 -3579 16562 -3545
rect 16596 -3579 16612 -3545
rect 16348 -3595 16612 -3579
rect 16034 -3637 16306 -3615
rect 11710 -3663 11920 -3637
rect 13642 -3663 14588 -3637
rect 14838 -3663 15784 -3637
rect 16034 -3663 16612 -3637
rect -2918 -3799 -2340 -3773
rect -1538 -3799 -960 -3773
rect -802 -3799 -224 -3773
rect 26 -3799 236 -3773
rect 505 -3799 535 -3773
rect 600 -3799 700 -3773
rect 860 -3799 960 -3773
rect 1032 -3799 1062 -3773
rect 1314 -3799 1524 -3773
rect 1774 -3799 2352 -3773
rect 2602 -3799 2812 -3773
rect 3081 -3799 3111 -3773
rect 3176 -3799 3276 -3773
rect 3436 -3799 3536 -3773
rect 3608 -3799 3638 -3773
rect 3890 -3799 4100 -3773
rect 4350 -3799 4928 -3773
rect 5178 -3799 5388 -3773
rect 5657 -3799 5687 -3773
rect 5752 -3799 5852 -3773
rect 6012 -3799 6112 -3773
rect 6184 -3799 6214 -3773
rect 6466 -3799 6676 -3773
rect 6926 -3799 7504 -3773
rect 7754 -3799 7964 -3773
rect 8233 -3799 8263 -3773
rect 8328 -3799 8428 -3773
rect 8588 -3799 8688 -3773
rect 8760 -3799 8790 -3773
rect 9042 -3799 9252 -3773
rect 9502 -3799 10080 -3773
rect 10422 -3799 10632 -3773
rect 10809 -3799 10839 -3773
rect 10904 -3799 11004 -3773
rect 11164 -3799 11264 -3773
rect 11336 -3799 11366 -3773
rect 11710 -3799 11920 -3773
rect 13642 -3799 14588 -3773
rect 14838 -3799 15784 -3773
rect 16034 -3799 16612 -3773
rect -2918 -3867 -2340 -3841
rect -1538 -3867 -960 -3841
rect -802 -3867 -224 -3841
rect 26 -3867 236 -3841
rect 488 -3867 518 -3841
rect 590 -3867 690 -3841
rect 850 -3867 950 -3841
rect 1015 -3867 1045 -3841
rect 1314 -3867 1524 -3841
rect 1774 -3867 2352 -3841
rect 2602 -3867 2812 -3841
rect 3064 -3867 3094 -3841
rect 3166 -3867 3266 -3841
rect 3426 -3867 3526 -3841
rect 3591 -3867 3621 -3841
rect 3890 -3867 4100 -3841
rect 4350 -3867 4928 -3841
rect 5178 -3867 5388 -3841
rect 5640 -3867 5670 -3841
rect 5742 -3867 5842 -3841
rect 6002 -3867 6102 -3841
rect 6167 -3867 6197 -3841
rect 6466 -3867 6676 -3841
rect 6926 -3867 7504 -3841
rect 7754 -3867 7964 -3841
rect 8216 -3867 8246 -3841
rect 8318 -3867 8418 -3841
rect 8578 -3867 8678 -3841
rect 8743 -3867 8773 -3841
rect 9042 -3867 9252 -3841
rect 9502 -3867 10080 -3841
rect 10422 -3867 10632 -3841
rect 10792 -3867 10822 -3841
rect 10894 -3867 10994 -3841
rect 11154 -3867 11254 -3841
rect 11319 -3867 11349 -3841
rect 11710 -3867 11920 -3841
rect 12633 -3867 12663 -3841
rect 12719 -3867 12749 -3841
rect 12805 -3867 12835 -3841
rect 12891 -3867 12921 -3841
rect 13274 -3867 13484 -3841
rect 13735 -3867 13765 -3841
rect 13821 -3867 13851 -3841
rect 13907 -3867 13937 -3841
rect 13993 -3867 14023 -3841
rect 14079 -3867 14109 -3841
rect 14165 -3867 14195 -3841
rect 14251 -3867 14281 -3841
rect 14337 -3867 14367 -3841
rect 14423 -3867 14453 -3841
rect 14509 -3867 14539 -3841
rect 14595 -3867 14625 -3841
rect 14681 -3867 14711 -3841
rect 14766 -3867 14796 -3841
rect 14852 -3867 14882 -3841
rect 14938 -3867 14968 -3841
rect 15024 -3867 15054 -3841
rect 15110 -3867 15140 -3841
rect 15196 -3867 15226 -3841
rect 15282 -3867 15312 -3841
rect 15368 -3867 15398 -3841
rect 15666 -3867 16612 -3841
rect -2918 -4003 -2340 -3977
rect -1538 -4003 -960 -3977
rect -802 -4003 -224 -3977
rect -2918 -4025 -2646 -4003
rect -2918 -4059 -2902 -4025
rect -2868 -4059 -2799 -4025
rect -2765 -4059 -2696 -4025
rect -2662 -4059 -2646 -4025
rect -1232 -4025 -960 -4003
rect -2918 -4075 -2646 -4059
rect -2604 -4061 -2340 -4045
rect -2604 -4095 -2588 -4061
rect -2554 -4095 -2489 -4061
rect -2455 -4095 -2390 -4061
rect -2356 -4095 -2340 -4061
rect -2604 -4117 -2340 -4095
rect -2918 -4143 -2340 -4117
rect -1538 -4061 -1274 -4045
rect -1538 -4095 -1522 -4061
rect -1488 -4095 -1423 -4061
rect -1389 -4095 -1324 -4061
rect -1290 -4095 -1274 -4061
rect -1232 -4059 -1216 -4025
rect -1182 -4059 -1113 -4025
rect -1079 -4059 -1010 -4025
rect -976 -4059 -960 -4025
rect -496 -4025 -224 -4003
rect 26 -4003 236 -3977
rect 26 -4009 110 -4003
rect -1232 -4075 -960 -4059
rect -802 -4061 -538 -4045
rect -1538 -4117 -1274 -4095
rect -802 -4095 -786 -4061
rect -752 -4095 -687 -4061
rect -653 -4095 -588 -4061
rect -554 -4095 -538 -4061
rect -496 -4059 -480 -4025
rect -446 -4059 -377 -4025
rect -343 -4059 -274 -4025
rect -240 -4059 -224 -4025
rect -496 -4075 -224 -4059
rect -32 -4025 110 -4009
rect 488 -4023 518 -3951
rect -32 -4059 -16 -4025
rect 18 -4059 110 -4025
rect 448 -4035 518 -4023
rect 590 -4025 690 -3997
rect 850 -4025 950 -3997
rect 1015 -4019 1045 -3951
rect 1314 -4003 1524 -3977
rect 1774 -4003 2352 -3977
rect 2602 -4003 2812 -3977
rect 1314 -4009 1398 -4003
rect -32 -4075 110 -4059
rect 152 -4061 294 -4045
rect -802 -4117 -538 -4095
rect 152 -4095 244 -4061
rect 278 -4095 294 -4061
rect 448 -4069 464 -4035
rect 498 -4069 518 -4035
rect 448 -4082 518 -4069
rect 568 -4035 690 -4025
rect 568 -4069 584 -4035
rect 618 -4069 690 -4035
rect 568 -4079 690 -4069
rect 789 -4035 950 -4025
rect 789 -4069 805 -4035
rect 839 -4069 950 -4035
rect 789 -4079 950 -4069
rect 152 -4111 294 -4095
rect 152 -4117 236 -4111
rect 488 -4117 518 -4082
rect -1538 -4143 -960 -4117
rect -802 -4143 -224 -4117
rect 26 -4143 236 -4117
rect 590 -4153 690 -4079
rect 850 -4153 950 -4079
rect 995 -4035 1049 -4019
rect 995 -4069 1005 -4035
rect 1039 -4069 1049 -4035
rect 995 -4085 1049 -4069
rect 1256 -4025 1398 -4009
rect 1256 -4059 1272 -4025
rect 1306 -4059 1398 -4025
rect 1774 -4025 2046 -4003
rect 2602 -4009 2686 -4003
rect 1256 -4075 1398 -4059
rect 1440 -4061 1582 -4045
rect 1015 -4117 1045 -4085
rect 1440 -4095 1532 -4061
rect 1566 -4095 1582 -4061
rect 1774 -4059 1790 -4025
rect 1824 -4059 1893 -4025
rect 1927 -4059 1996 -4025
rect 2030 -4059 2046 -4025
rect 2544 -4025 2686 -4009
rect 3064 -4023 3094 -3951
rect 1774 -4075 2046 -4059
rect 2088 -4061 2352 -4045
rect 1440 -4111 1582 -4095
rect 2088 -4095 2104 -4061
rect 2138 -4095 2203 -4061
rect 2237 -4095 2302 -4061
rect 2336 -4095 2352 -4061
rect 2544 -4059 2560 -4025
rect 2594 -4059 2686 -4025
rect 3024 -4035 3094 -4023
rect 3166 -4025 3266 -3997
rect 3426 -4025 3526 -3997
rect 3591 -4019 3621 -3951
rect 3890 -4003 4100 -3977
rect 4350 -4003 4928 -3977
rect 5178 -4003 5388 -3977
rect 3890 -4009 3974 -4003
rect 2544 -4075 2686 -4059
rect 2728 -4061 2870 -4045
rect 1440 -4117 1524 -4111
rect 2088 -4117 2352 -4095
rect 2728 -4095 2820 -4061
rect 2854 -4095 2870 -4061
rect 3024 -4069 3040 -4035
rect 3074 -4069 3094 -4035
rect 3024 -4082 3094 -4069
rect 3144 -4035 3266 -4025
rect 3144 -4069 3160 -4035
rect 3194 -4069 3266 -4035
rect 3144 -4079 3266 -4069
rect 3365 -4035 3526 -4025
rect 3365 -4069 3381 -4035
rect 3415 -4069 3526 -4035
rect 3365 -4079 3526 -4069
rect 2728 -4111 2870 -4095
rect 2728 -4117 2812 -4111
rect 3064 -4117 3094 -4082
rect 1314 -4143 1524 -4117
rect 1774 -4143 2352 -4117
rect 2602 -4143 2812 -4117
rect 3166 -4153 3266 -4079
rect 3426 -4153 3526 -4079
rect 3571 -4035 3625 -4019
rect 3571 -4069 3581 -4035
rect 3615 -4069 3625 -4035
rect 3571 -4085 3625 -4069
rect 3832 -4025 3974 -4009
rect 3832 -4059 3848 -4025
rect 3882 -4059 3974 -4025
rect 4350 -4025 4622 -4003
rect 5178 -4009 5262 -4003
rect 3832 -4075 3974 -4059
rect 4016 -4061 4158 -4045
rect 3591 -4117 3621 -4085
rect 4016 -4095 4108 -4061
rect 4142 -4095 4158 -4061
rect 4350 -4059 4366 -4025
rect 4400 -4059 4469 -4025
rect 4503 -4059 4572 -4025
rect 4606 -4059 4622 -4025
rect 5120 -4025 5262 -4009
rect 5640 -4023 5670 -3951
rect 4350 -4075 4622 -4059
rect 4664 -4061 4928 -4045
rect 4016 -4111 4158 -4095
rect 4664 -4095 4680 -4061
rect 4714 -4095 4779 -4061
rect 4813 -4095 4878 -4061
rect 4912 -4095 4928 -4061
rect 5120 -4059 5136 -4025
rect 5170 -4059 5262 -4025
rect 5600 -4035 5670 -4023
rect 5742 -4025 5842 -3997
rect 6002 -4025 6102 -3997
rect 6167 -4019 6197 -3951
rect 6466 -4003 6676 -3977
rect 6926 -4003 7504 -3977
rect 7754 -4003 7964 -3977
rect 6466 -4009 6550 -4003
rect 5120 -4075 5262 -4059
rect 5304 -4061 5446 -4045
rect 4016 -4117 4100 -4111
rect 4664 -4117 4928 -4095
rect 5304 -4095 5396 -4061
rect 5430 -4095 5446 -4061
rect 5600 -4069 5616 -4035
rect 5650 -4069 5670 -4035
rect 5600 -4082 5670 -4069
rect 5720 -4035 5842 -4025
rect 5720 -4069 5736 -4035
rect 5770 -4069 5842 -4035
rect 5720 -4079 5842 -4069
rect 5941 -4035 6102 -4025
rect 5941 -4069 5957 -4035
rect 5991 -4069 6102 -4035
rect 5941 -4079 6102 -4069
rect 5304 -4111 5446 -4095
rect 5304 -4117 5388 -4111
rect 5640 -4117 5670 -4082
rect 3890 -4143 4100 -4117
rect 4350 -4143 4928 -4117
rect 5178 -4143 5388 -4117
rect 5742 -4153 5842 -4079
rect 6002 -4153 6102 -4079
rect 6147 -4035 6201 -4019
rect 6147 -4069 6157 -4035
rect 6191 -4069 6201 -4035
rect 6147 -4085 6201 -4069
rect 6408 -4025 6550 -4009
rect 6408 -4059 6424 -4025
rect 6458 -4059 6550 -4025
rect 6926 -4025 7198 -4003
rect 7754 -4009 7838 -4003
rect 6408 -4075 6550 -4059
rect 6592 -4061 6734 -4045
rect 6167 -4117 6197 -4085
rect 6592 -4095 6684 -4061
rect 6718 -4095 6734 -4061
rect 6926 -4059 6942 -4025
rect 6976 -4059 7045 -4025
rect 7079 -4059 7148 -4025
rect 7182 -4059 7198 -4025
rect 7696 -4025 7838 -4009
rect 8216 -4023 8246 -3951
rect 6926 -4075 7198 -4059
rect 7240 -4061 7504 -4045
rect 6592 -4111 6734 -4095
rect 7240 -4095 7256 -4061
rect 7290 -4095 7355 -4061
rect 7389 -4095 7454 -4061
rect 7488 -4095 7504 -4061
rect 7696 -4059 7712 -4025
rect 7746 -4059 7838 -4025
rect 8176 -4035 8246 -4023
rect 8318 -4025 8418 -3997
rect 8578 -4025 8678 -3997
rect 8743 -4019 8773 -3951
rect 9042 -4003 9252 -3977
rect 9502 -4003 10080 -3977
rect 10422 -4003 10632 -3977
rect 9042 -4009 9126 -4003
rect 7696 -4075 7838 -4059
rect 7880 -4061 8022 -4045
rect 6592 -4117 6676 -4111
rect 7240 -4117 7504 -4095
rect 7880 -4095 7972 -4061
rect 8006 -4095 8022 -4061
rect 8176 -4069 8192 -4035
rect 8226 -4069 8246 -4035
rect 8176 -4082 8246 -4069
rect 8296 -4035 8418 -4025
rect 8296 -4069 8312 -4035
rect 8346 -4069 8418 -4035
rect 8296 -4079 8418 -4069
rect 8517 -4035 8678 -4025
rect 8517 -4069 8533 -4035
rect 8567 -4069 8678 -4035
rect 8517 -4079 8678 -4069
rect 7880 -4111 8022 -4095
rect 7880 -4117 7964 -4111
rect 8216 -4117 8246 -4082
rect 6466 -4143 6676 -4117
rect 6926 -4143 7504 -4117
rect 7754 -4143 7964 -4117
rect 8318 -4153 8418 -4079
rect 8578 -4153 8678 -4079
rect 8723 -4035 8777 -4019
rect 8723 -4069 8733 -4035
rect 8767 -4069 8777 -4035
rect 8723 -4085 8777 -4069
rect 8984 -4025 9126 -4009
rect 8984 -4059 9000 -4025
rect 9034 -4059 9126 -4025
rect 9502 -4025 9774 -4003
rect 10422 -4009 10506 -4003
rect 8984 -4075 9126 -4059
rect 9168 -4061 9310 -4045
rect 8743 -4117 8773 -4085
rect 9168 -4095 9260 -4061
rect 9294 -4095 9310 -4061
rect 9502 -4059 9518 -4025
rect 9552 -4059 9621 -4025
rect 9655 -4059 9724 -4025
rect 9758 -4059 9774 -4025
rect 10364 -4025 10506 -4009
rect 10792 -4023 10822 -3951
rect 9502 -4075 9774 -4059
rect 9816 -4061 10080 -4045
rect 9168 -4111 9310 -4095
rect 9816 -4095 9832 -4061
rect 9866 -4095 9931 -4061
rect 9965 -4095 10030 -4061
rect 10064 -4095 10080 -4061
rect 10364 -4059 10380 -4025
rect 10414 -4059 10506 -4025
rect 10752 -4035 10822 -4023
rect 10894 -4025 10994 -3997
rect 11154 -4025 11254 -3997
rect 11319 -4019 11349 -3951
rect 11710 -4003 11920 -3977
rect 11710 -4009 11794 -4003
rect 10364 -4075 10506 -4059
rect 10548 -4061 10690 -4045
rect 9168 -4117 9252 -4111
rect 9816 -4117 10080 -4095
rect 10548 -4095 10640 -4061
rect 10674 -4095 10690 -4061
rect 10752 -4069 10768 -4035
rect 10802 -4069 10822 -4035
rect 10752 -4082 10822 -4069
rect 10872 -4035 10994 -4025
rect 10872 -4069 10888 -4035
rect 10922 -4069 10994 -4035
rect 10872 -4079 10994 -4069
rect 11093 -4035 11254 -4025
rect 11093 -4069 11109 -4035
rect 11143 -4069 11254 -4035
rect 11093 -4079 11254 -4069
rect 10548 -4111 10690 -4095
rect 10548 -4117 10632 -4111
rect 10792 -4117 10822 -4082
rect 9042 -4143 9252 -4117
rect 9502 -4143 10080 -4117
rect 10422 -4143 10632 -4117
rect 10894 -4153 10994 -4079
rect 11154 -4153 11254 -4079
rect 11299 -4035 11353 -4019
rect 11299 -4069 11309 -4035
rect 11343 -4069 11353 -4035
rect 11299 -4085 11353 -4069
rect 11652 -4025 11794 -4009
rect 12633 -4025 12663 -3951
rect 12719 -4025 12749 -3951
rect 12805 -4025 12835 -3951
rect 12891 -4025 12921 -3951
rect 13274 -4003 13484 -3977
rect 13735 -4000 13765 -3951
rect 13821 -4000 13851 -3951
rect 13907 -4000 13937 -3951
rect 13993 -4000 14023 -3951
rect 13400 -4009 13484 -4003
rect 13400 -4025 13542 -4009
rect 11652 -4059 11668 -4025
rect 11702 -4059 11794 -4025
rect 12547 -4035 13007 -4025
rect 11652 -4075 11794 -4059
rect 11836 -4061 11978 -4045
rect 11319 -4117 11349 -4085
rect 11836 -4095 11928 -4061
rect 11962 -4095 11978 -4061
rect 11836 -4111 11978 -4095
rect 12547 -4069 12574 -4035
rect 12608 -4069 12642 -4035
rect 12676 -4069 12710 -4035
rect 12744 -4069 12778 -4035
rect 12812 -4069 12846 -4035
rect 12880 -4069 12914 -4035
rect 12948 -4069 13007 -4035
rect 12547 -4079 13007 -4069
rect 11836 -4117 11920 -4111
rect 12547 -4117 12577 -4079
rect 12633 -4117 12663 -4079
rect 12719 -4117 12749 -4079
rect 12805 -4117 12835 -4079
rect 12891 -4117 12921 -4079
rect 12977 -4117 13007 -4079
rect 13216 -4061 13358 -4045
rect 13216 -4095 13232 -4061
rect 13266 -4095 13358 -4061
rect 13400 -4059 13492 -4025
rect 13526 -4059 13542 -4025
rect 13400 -4075 13542 -4059
rect 13676 -4035 14023 -4000
rect 13676 -4069 13692 -4035
rect 13726 -4069 14023 -4035
rect 13216 -4111 13358 -4095
rect 13676 -4102 14023 -4069
rect 13274 -4117 13358 -4111
rect 13735 -4117 13765 -4102
rect 13821 -4117 13851 -4102
rect 13907 -4117 13937 -4102
rect 13993 -4117 14023 -4102
rect 14079 -4010 14109 -3951
rect 14165 -4010 14195 -3951
rect 14251 -4010 14281 -3951
rect 14337 -4010 14367 -3951
rect 14423 -4010 14453 -3951
rect 14509 -4010 14539 -3951
rect 14595 -4010 14625 -3951
rect 14681 -4010 14711 -3951
rect 14766 -4010 14796 -3951
rect 14852 -4010 14882 -3951
rect 14938 -4010 14968 -3951
rect 15024 -4010 15054 -3951
rect 15110 -4010 15140 -3951
rect 15196 -4010 15226 -3951
rect 15282 -4010 15312 -3951
rect 15368 -4010 15398 -3951
rect 15666 -4003 16612 -3977
rect 14079 -4035 15398 -4010
rect 14079 -4069 14119 -4035
rect 14153 -4069 14187 -4035
rect 14221 -4069 14255 -4035
rect 14289 -4069 14323 -4035
rect 14357 -4069 14391 -4035
rect 14425 -4069 14459 -4035
rect 14493 -4069 14527 -4035
rect 14561 -4069 14595 -4035
rect 14629 -4069 14663 -4035
rect 14697 -4069 14731 -4035
rect 14765 -4069 14799 -4035
rect 14833 -4069 14867 -4035
rect 14901 -4069 14935 -4035
rect 14969 -4069 15003 -4035
rect 15037 -4069 15071 -4035
rect 15105 -4069 15139 -4035
rect 15173 -4069 15398 -4035
rect 16158 -4025 16612 -4003
rect 14079 -4085 15398 -4069
rect 14079 -4117 14109 -4085
rect 14165 -4117 14195 -4085
rect 14251 -4117 14281 -4085
rect 14337 -4117 14367 -4085
rect 14423 -4117 14453 -4085
rect 14509 -4117 14539 -4085
rect 14595 -4117 14625 -4085
rect 14681 -4117 14711 -4085
rect 14766 -4117 14796 -4085
rect 14852 -4117 14882 -4085
rect 14938 -4117 14968 -4085
rect 15024 -4117 15054 -4085
rect 15110 -4117 15140 -4085
rect 15196 -4117 15226 -4085
rect 15282 -4117 15312 -4085
rect 15368 -4117 15398 -4085
rect 15666 -4061 16116 -4045
rect 15666 -4095 15682 -4061
rect 15716 -4095 15810 -4061
rect 15844 -4095 15938 -4061
rect 15972 -4095 16066 -4061
rect 16100 -4095 16116 -4061
rect 16158 -4059 16174 -4025
rect 16208 -4059 16302 -4025
rect 16336 -4059 16430 -4025
rect 16464 -4059 16558 -4025
rect 16592 -4059 16612 -4025
rect 16158 -4075 16612 -4059
rect 15666 -4117 16116 -4095
rect 11710 -4143 11920 -4117
rect 13274 -4143 13484 -4117
rect 15666 -4143 16612 -4117
rect -2918 -4343 -2340 -4317
rect -1538 -4343 -960 -4317
rect -802 -4343 -224 -4317
rect 26 -4343 236 -4317
rect 488 -4343 518 -4317
rect 590 -4343 690 -4317
rect 850 -4343 950 -4317
rect 1015 -4343 1045 -4317
rect 1314 -4343 1524 -4317
rect 1774 -4343 2352 -4317
rect 2602 -4343 2812 -4317
rect 3064 -4343 3094 -4317
rect 3166 -4343 3266 -4317
rect 3426 -4343 3526 -4317
rect 3591 -4343 3621 -4317
rect 3890 -4343 4100 -4317
rect 4350 -4343 4928 -4317
rect 5178 -4343 5388 -4317
rect 5640 -4343 5670 -4317
rect 5742 -4343 5842 -4317
rect 6002 -4343 6102 -4317
rect 6167 -4343 6197 -4317
rect 6466 -4343 6676 -4317
rect 6926 -4343 7504 -4317
rect 7754 -4343 7964 -4317
rect 8216 -4343 8246 -4317
rect 8318 -4343 8418 -4317
rect 8578 -4343 8678 -4317
rect 8743 -4343 8773 -4317
rect 9042 -4343 9252 -4317
rect 9502 -4343 10080 -4317
rect 10422 -4343 10632 -4317
rect 10792 -4343 10822 -4317
rect 10894 -4343 10994 -4317
rect 11154 -4343 11254 -4317
rect 11319 -4343 11349 -4317
rect 11710 -4343 11920 -4317
rect 12547 -4343 12577 -4317
rect 12633 -4343 12663 -4317
rect 12719 -4343 12749 -4317
rect 12805 -4343 12835 -4317
rect 12891 -4343 12921 -4317
rect 12977 -4343 13007 -4317
rect 13274 -4343 13484 -4317
rect 13735 -4343 13765 -4317
rect 13821 -4343 13851 -4317
rect 13907 -4343 13937 -4317
rect 13993 -4343 14023 -4317
rect 14079 -4343 14109 -4317
rect 14165 -4343 14195 -4317
rect 14251 -4343 14281 -4317
rect 14337 -4343 14367 -4317
rect 14423 -4343 14453 -4317
rect 14509 -4343 14539 -4317
rect 14595 -4343 14625 -4317
rect 14681 -4343 14711 -4317
rect 14766 -4343 14796 -4317
rect 14852 -4343 14882 -4317
rect 14938 -4343 14968 -4317
rect 15024 -4343 15054 -4317
rect 15110 -4343 15140 -4317
rect 15196 -4343 15226 -4317
rect 15282 -4343 15312 -4317
rect 15368 -4343 15398 -4317
rect 15666 -4343 16612 -4317
rect -2918 -4411 -2340 -4385
rect -1538 -4411 -960 -4385
rect -783 -4411 -753 -4385
rect -688 -4411 -588 -4385
rect -428 -4411 -328 -4385
rect -256 -4411 -226 -4385
rect 26 -4411 236 -4385
rect 505 -4411 535 -4385
rect 600 -4411 700 -4385
rect 860 -4411 960 -4385
rect 1032 -4411 1062 -4385
rect 1314 -4411 1524 -4385
rect 1774 -4411 2352 -4385
rect 2602 -4411 2812 -4385
rect 3081 -4411 3111 -4385
rect 3176 -4411 3276 -4385
rect 3436 -4411 3536 -4385
rect 3608 -4411 3638 -4385
rect 3890 -4411 4100 -4385
rect 4350 -4411 4928 -4385
rect 5178 -4411 5388 -4385
rect 5657 -4411 5687 -4385
rect 5752 -4411 5852 -4385
rect 6012 -4411 6112 -4385
rect 6184 -4411 6214 -4385
rect 6466 -4411 6676 -4385
rect 6926 -4411 7504 -4385
rect 7754 -4411 7964 -4385
rect 8233 -4411 8263 -4385
rect 8328 -4411 8428 -4385
rect 8588 -4411 8688 -4385
rect 8760 -4411 8790 -4385
rect 9042 -4411 9252 -4385
rect 9502 -4411 10080 -4385
rect 10422 -4411 10632 -4385
rect 10809 -4411 10839 -4385
rect 10904 -4411 11004 -4385
rect 11164 -4411 11264 -4385
rect 11336 -4411 11366 -4385
rect 11710 -4411 11920 -4385
rect 13735 -4411 13765 -4385
rect 13821 -4411 13851 -4385
rect 13907 -4411 13937 -4385
rect 13993 -4411 14023 -4385
rect 14079 -4411 14109 -4385
rect 14165 -4411 14195 -4385
rect 14251 -4411 14281 -4385
rect 14337 -4411 14367 -4385
rect 14423 -4411 14453 -4385
rect 14509 -4411 14539 -4385
rect 14595 -4411 14625 -4385
rect 14681 -4411 14711 -4385
rect 14766 -4411 14796 -4385
rect 14852 -4411 14882 -4385
rect 14938 -4411 14968 -4385
rect 15024 -4411 15054 -4385
rect 15110 -4411 15140 -4385
rect 15196 -4411 15226 -4385
rect 15282 -4411 15312 -4385
rect 15368 -4411 15398 -4385
rect 15666 -4411 16612 -4385
rect -2918 -4611 -2340 -4585
rect -1538 -4611 -960 -4585
rect -2918 -4633 -2654 -4611
rect -2918 -4667 -2902 -4633
rect -2868 -4667 -2803 -4633
rect -2769 -4667 -2704 -4633
rect -2670 -4667 -2654 -4633
rect -1224 -4633 -960 -4611
rect -2918 -4683 -2654 -4667
rect -2612 -4669 -2340 -4653
rect -2612 -4703 -2596 -4669
rect -2562 -4703 -2493 -4669
rect -2459 -4703 -2390 -4669
rect -2356 -4703 -2340 -4669
rect -2612 -4725 -2340 -4703
rect -2918 -4751 -2340 -4725
rect -1538 -4669 -1266 -4653
rect -1538 -4703 -1522 -4669
rect -1488 -4703 -1419 -4669
rect -1385 -4703 -1316 -4669
rect -1282 -4703 -1266 -4669
rect -1224 -4667 -1208 -4633
rect -1174 -4667 -1109 -4633
rect -1075 -4667 -1010 -4633
rect -976 -4667 -960 -4633
rect -783 -4643 -753 -4611
rect -1224 -4683 -960 -4667
rect -787 -4659 -733 -4643
rect -1538 -4725 -1266 -4703
rect -787 -4693 -777 -4659
rect -743 -4693 -733 -4659
rect -787 -4709 -733 -4693
rect -688 -4649 -588 -4575
rect -428 -4649 -328 -4575
rect 26 -4611 236 -4585
rect -256 -4646 -226 -4611
rect 152 -4617 236 -4611
rect 152 -4633 294 -4617
rect -688 -4659 -527 -4649
rect -688 -4693 -577 -4659
rect -543 -4693 -527 -4659
rect -688 -4703 -527 -4693
rect -428 -4659 -306 -4649
rect -428 -4693 -356 -4659
rect -322 -4693 -306 -4659
rect -428 -4703 -306 -4693
rect -256 -4659 -186 -4646
rect -256 -4693 -236 -4659
rect -202 -4693 -186 -4659
rect -1538 -4751 -960 -4725
rect -783 -4777 -753 -4709
rect -688 -4731 -588 -4703
rect -428 -4731 -328 -4703
rect -256 -4705 -186 -4693
rect -32 -4669 110 -4653
rect -32 -4703 -16 -4669
rect 18 -4703 110 -4669
rect 152 -4667 244 -4633
rect 278 -4667 294 -4633
rect 505 -4643 535 -4611
rect 152 -4683 294 -4667
rect 501 -4659 555 -4643
rect -256 -4777 -226 -4705
rect -32 -4719 110 -4703
rect 501 -4693 511 -4659
rect 545 -4693 555 -4659
rect 501 -4709 555 -4693
rect 600 -4649 700 -4575
rect 860 -4649 960 -4575
rect 1314 -4611 1524 -4585
rect 1032 -4646 1062 -4611
rect 1440 -4617 1524 -4611
rect 1774 -4611 2352 -4585
rect 2602 -4611 2812 -4585
rect 1440 -4633 1582 -4617
rect 600 -4659 761 -4649
rect 600 -4693 711 -4659
rect 745 -4693 761 -4659
rect 600 -4703 761 -4693
rect 860 -4659 982 -4649
rect 860 -4693 932 -4659
rect 966 -4693 982 -4659
rect 860 -4703 982 -4693
rect 1032 -4659 1102 -4646
rect 1032 -4693 1052 -4659
rect 1086 -4693 1102 -4659
rect 26 -4725 110 -4719
rect 26 -4751 236 -4725
rect 505 -4777 535 -4709
rect 600 -4731 700 -4703
rect 860 -4731 960 -4703
rect 1032 -4705 1102 -4693
rect 1256 -4669 1398 -4653
rect 1256 -4703 1272 -4669
rect 1306 -4703 1398 -4669
rect 1440 -4667 1532 -4633
rect 1566 -4667 1582 -4633
rect 1440 -4683 1582 -4667
rect 1774 -4633 2038 -4611
rect 1774 -4667 1790 -4633
rect 1824 -4667 1889 -4633
rect 1923 -4667 1988 -4633
rect 2022 -4667 2038 -4633
rect 2728 -4617 2812 -4611
rect 2728 -4633 2870 -4617
rect 1774 -4683 2038 -4667
rect 2080 -4669 2352 -4653
rect 1032 -4777 1062 -4705
rect 1256 -4719 1398 -4703
rect 1314 -4725 1398 -4719
rect 2080 -4703 2096 -4669
rect 2130 -4703 2199 -4669
rect 2233 -4703 2302 -4669
rect 2336 -4703 2352 -4669
rect 2080 -4725 2352 -4703
rect 2544 -4669 2686 -4653
rect 2544 -4703 2560 -4669
rect 2594 -4703 2686 -4669
rect 2728 -4667 2820 -4633
rect 2854 -4667 2870 -4633
rect 3081 -4643 3111 -4611
rect 2728 -4683 2870 -4667
rect 3077 -4659 3131 -4643
rect 2544 -4719 2686 -4703
rect 3077 -4693 3087 -4659
rect 3121 -4693 3131 -4659
rect 3077 -4709 3131 -4693
rect 3176 -4649 3276 -4575
rect 3436 -4649 3536 -4575
rect 3890 -4611 4100 -4585
rect 3608 -4646 3638 -4611
rect 4016 -4617 4100 -4611
rect 4350 -4611 4928 -4585
rect 5178 -4611 5388 -4585
rect 4016 -4633 4158 -4617
rect 3176 -4659 3337 -4649
rect 3176 -4693 3287 -4659
rect 3321 -4693 3337 -4659
rect 3176 -4703 3337 -4693
rect 3436 -4659 3558 -4649
rect 3436 -4693 3508 -4659
rect 3542 -4693 3558 -4659
rect 3436 -4703 3558 -4693
rect 3608 -4659 3678 -4646
rect 3608 -4693 3628 -4659
rect 3662 -4693 3678 -4659
rect 1314 -4751 1524 -4725
rect 1774 -4751 2352 -4725
rect 2602 -4725 2686 -4719
rect 2602 -4751 2812 -4725
rect 3081 -4777 3111 -4709
rect 3176 -4731 3276 -4703
rect 3436 -4731 3536 -4703
rect 3608 -4705 3678 -4693
rect 3832 -4669 3974 -4653
rect 3832 -4703 3848 -4669
rect 3882 -4703 3974 -4669
rect 4016 -4667 4108 -4633
rect 4142 -4667 4158 -4633
rect 4016 -4683 4158 -4667
rect 4350 -4633 4614 -4611
rect 4350 -4667 4366 -4633
rect 4400 -4667 4465 -4633
rect 4499 -4667 4564 -4633
rect 4598 -4667 4614 -4633
rect 5304 -4617 5388 -4611
rect 5304 -4633 5446 -4617
rect 4350 -4683 4614 -4667
rect 4656 -4669 4928 -4653
rect 3608 -4777 3638 -4705
rect 3832 -4719 3974 -4703
rect 3890 -4725 3974 -4719
rect 4656 -4703 4672 -4669
rect 4706 -4703 4775 -4669
rect 4809 -4703 4878 -4669
rect 4912 -4703 4928 -4669
rect 4656 -4725 4928 -4703
rect 5120 -4669 5262 -4653
rect 5120 -4703 5136 -4669
rect 5170 -4703 5262 -4669
rect 5304 -4667 5396 -4633
rect 5430 -4667 5446 -4633
rect 5657 -4643 5687 -4611
rect 5304 -4683 5446 -4667
rect 5653 -4659 5707 -4643
rect 5120 -4719 5262 -4703
rect 5653 -4693 5663 -4659
rect 5697 -4693 5707 -4659
rect 5653 -4709 5707 -4693
rect 5752 -4649 5852 -4575
rect 6012 -4649 6112 -4575
rect 6466 -4611 6676 -4585
rect 6184 -4646 6214 -4611
rect 6592 -4617 6676 -4611
rect 6926 -4611 7504 -4585
rect 7754 -4611 7964 -4585
rect 6592 -4633 6734 -4617
rect 5752 -4659 5913 -4649
rect 5752 -4693 5863 -4659
rect 5897 -4693 5913 -4659
rect 5752 -4703 5913 -4693
rect 6012 -4659 6134 -4649
rect 6012 -4693 6084 -4659
rect 6118 -4693 6134 -4659
rect 6012 -4703 6134 -4693
rect 6184 -4659 6254 -4646
rect 6184 -4693 6204 -4659
rect 6238 -4693 6254 -4659
rect 3890 -4751 4100 -4725
rect 4350 -4751 4928 -4725
rect 5178 -4725 5262 -4719
rect 5178 -4751 5388 -4725
rect 5657 -4777 5687 -4709
rect 5752 -4731 5852 -4703
rect 6012 -4731 6112 -4703
rect 6184 -4705 6254 -4693
rect 6408 -4669 6550 -4653
rect 6408 -4703 6424 -4669
rect 6458 -4703 6550 -4669
rect 6592 -4667 6684 -4633
rect 6718 -4667 6734 -4633
rect 6592 -4683 6734 -4667
rect 6926 -4633 7190 -4611
rect 6926 -4667 6942 -4633
rect 6976 -4667 7041 -4633
rect 7075 -4667 7140 -4633
rect 7174 -4667 7190 -4633
rect 7880 -4617 7964 -4611
rect 7880 -4633 8022 -4617
rect 6926 -4683 7190 -4667
rect 7232 -4669 7504 -4653
rect 6184 -4777 6214 -4705
rect 6408 -4719 6550 -4703
rect 6466 -4725 6550 -4719
rect 7232 -4703 7248 -4669
rect 7282 -4703 7351 -4669
rect 7385 -4703 7454 -4669
rect 7488 -4703 7504 -4669
rect 7232 -4725 7504 -4703
rect 7696 -4669 7838 -4653
rect 7696 -4703 7712 -4669
rect 7746 -4703 7838 -4669
rect 7880 -4667 7972 -4633
rect 8006 -4667 8022 -4633
rect 8233 -4643 8263 -4611
rect 7880 -4683 8022 -4667
rect 8229 -4659 8283 -4643
rect 7696 -4719 7838 -4703
rect 8229 -4693 8239 -4659
rect 8273 -4693 8283 -4659
rect 8229 -4709 8283 -4693
rect 8328 -4649 8428 -4575
rect 8588 -4649 8688 -4575
rect 9042 -4611 9252 -4585
rect 8760 -4646 8790 -4611
rect 9168 -4617 9252 -4611
rect 9502 -4611 10080 -4585
rect 10422 -4611 10632 -4585
rect 9168 -4633 9310 -4617
rect 8328 -4659 8489 -4649
rect 8328 -4693 8439 -4659
rect 8473 -4693 8489 -4659
rect 8328 -4703 8489 -4693
rect 8588 -4659 8710 -4649
rect 8588 -4693 8660 -4659
rect 8694 -4693 8710 -4659
rect 8588 -4703 8710 -4693
rect 8760 -4659 8830 -4646
rect 8760 -4693 8780 -4659
rect 8814 -4693 8830 -4659
rect 6466 -4751 6676 -4725
rect 6926 -4751 7504 -4725
rect 7754 -4725 7838 -4719
rect 7754 -4751 7964 -4725
rect 8233 -4777 8263 -4709
rect 8328 -4731 8428 -4703
rect 8588 -4731 8688 -4703
rect 8760 -4705 8830 -4693
rect 8984 -4669 9126 -4653
rect 8984 -4703 9000 -4669
rect 9034 -4703 9126 -4669
rect 9168 -4667 9260 -4633
rect 9294 -4667 9310 -4633
rect 9168 -4683 9310 -4667
rect 9502 -4633 9766 -4611
rect 9502 -4667 9518 -4633
rect 9552 -4667 9617 -4633
rect 9651 -4667 9716 -4633
rect 9750 -4667 9766 -4633
rect 10548 -4617 10632 -4611
rect 10548 -4633 10690 -4617
rect 9502 -4683 9766 -4667
rect 9808 -4669 10080 -4653
rect 8760 -4777 8790 -4705
rect 8984 -4719 9126 -4703
rect 9042 -4725 9126 -4719
rect 9808 -4703 9824 -4669
rect 9858 -4703 9927 -4669
rect 9961 -4703 10030 -4669
rect 10064 -4703 10080 -4669
rect 9808 -4725 10080 -4703
rect 10364 -4669 10506 -4653
rect 10364 -4703 10380 -4669
rect 10414 -4703 10506 -4669
rect 10548 -4667 10640 -4633
rect 10674 -4667 10690 -4633
rect 10809 -4643 10839 -4611
rect 10548 -4683 10690 -4667
rect 10805 -4659 10859 -4643
rect 10364 -4719 10506 -4703
rect 10805 -4693 10815 -4659
rect 10849 -4693 10859 -4659
rect 10805 -4709 10859 -4693
rect 10904 -4649 11004 -4575
rect 11164 -4649 11264 -4575
rect 11710 -4611 11920 -4585
rect 15666 -4611 16612 -4585
rect 11336 -4646 11366 -4611
rect 11836 -4617 11920 -4611
rect 11836 -4633 11978 -4617
rect 13735 -4626 13765 -4611
rect 13821 -4626 13851 -4611
rect 13907 -4626 13937 -4611
rect 13993 -4626 14023 -4611
rect 10904 -4659 11065 -4649
rect 10904 -4693 11015 -4659
rect 11049 -4693 11065 -4659
rect 10904 -4703 11065 -4693
rect 11164 -4659 11286 -4649
rect 11164 -4693 11236 -4659
rect 11270 -4693 11286 -4659
rect 11164 -4703 11286 -4693
rect 11336 -4659 11406 -4646
rect 11336 -4693 11356 -4659
rect 11390 -4693 11406 -4659
rect 9042 -4751 9252 -4725
rect 9502 -4751 10080 -4725
rect 10422 -4725 10506 -4719
rect 10422 -4751 10632 -4725
rect 10809 -4777 10839 -4709
rect 10904 -4731 11004 -4703
rect 11164 -4731 11264 -4703
rect 11336 -4705 11406 -4693
rect 11652 -4669 11794 -4653
rect 11652 -4703 11668 -4669
rect 11702 -4703 11794 -4669
rect 11836 -4667 11928 -4633
rect 11962 -4667 11978 -4633
rect 11836 -4683 11978 -4667
rect 13676 -4659 14023 -4626
rect 11336 -4777 11366 -4705
rect 11652 -4719 11794 -4703
rect 11710 -4725 11794 -4719
rect 13676 -4693 13692 -4659
rect 13726 -4693 14023 -4659
rect 11710 -4751 11920 -4725
rect 13676 -4728 14023 -4693
rect 13735 -4777 13765 -4728
rect 13821 -4777 13851 -4728
rect 13907 -4777 13937 -4728
rect 13993 -4777 14023 -4728
rect 14079 -4643 14109 -4611
rect 14165 -4643 14195 -4611
rect 14251 -4643 14281 -4611
rect 14337 -4643 14367 -4611
rect 14423 -4643 14453 -4611
rect 14509 -4643 14539 -4611
rect 14595 -4643 14625 -4611
rect 14681 -4643 14711 -4611
rect 14766 -4643 14796 -4611
rect 14852 -4643 14882 -4611
rect 14938 -4643 14968 -4611
rect 15024 -4643 15054 -4611
rect 15110 -4643 15140 -4611
rect 15196 -4643 15226 -4611
rect 15282 -4643 15312 -4611
rect 15368 -4643 15398 -4611
rect 14079 -4659 15398 -4643
rect 16162 -4633 16612 -4611
rect 14079 -4693 14119 -4659
rect 14153 -4693 14187 -4659
rect 14221 -4693 14255 -4659
rect 14289 -4693 14323 -4659
rect 14357 -4693 14391 -4659
rect 14425 -4693 14459 -4659
rect 14493 -4693 14527 -4659
rect 14561 -4693 14595 -4659
rect 14629 -4693 14663 -4659
rect 14697 -4693 14731 -4659
rect 14765 -4693 14799 -4659
rect 14833 -4693 14867 -4659
rect 14901 -4693 14935 -4659
rect 14969 -4693 15003 -4659
rect 15037 -4693 15071 -4659
rect 15105 -4693 15139 -4659
rect 15173 -4693 15398 -4659
rect 14079 -4718 15398 -4693
rect 14079 -4777 14109 -4718
rect 14165 -4777 14195 -4718
rect 14251 -4777 14281 -4718
rect 14337 -4777 14367 -4718
rect 14423 -4777 14453 -4718
rect 14509 -4777 14539 -4718
rect 14595 -4777 14625 -4718
rect 14681 -4777 14711 -4718
rect 14766 -4777 14796 -4718
rect 14852 -4777 14882 -4718
rect 14938 -4777 14968 -4718
rect 15024 -4777 15054 -4718
rect 15110 -4777 15140 -4718
rect 15196 -4777 15226 -4718
rect 15282 -4777 15312 -4718
rect 15368 -4777 15398 -4718
rect 15666 -4669 16120 -4653
rect 15666 -4703 15686 -4669
rect 15720 -4703 15814 -4669
rect 15848 -4703 15942 -4669
rect 15976 -4703 16070 -4669
rect 16104 -4703 16120 -4669
rect 16162 -4667 16178 -4633
rect 16212 -4667 16306 -4633
rect 16340 -4667 16434 -4633
rect 16468 -4667 16562 -4633
rect 16596 -4667 16612 -4633
rect 16162 -4683 16612 -4667
rect 15666 -4725 16120 -4703
rect 15666 -4751 16612 -4725
rect -2918 -4887 -2340 -4861
rect -1538 -4887 -960 -4861
rect -783 -4887 -753 -4861
rect -688 -4887 -588 -4861
rect -428 -4887 -328 -4861
rect -256 -4887 -226 -4861
rect 26 -4887 236 -4861
rect 505 -4887 535 -4861
rect 600 -4887 700 -4861
rect 860 -4887 960 -4861
rect 1032 -4887 1062 -4861
rect 1314 -4887 1524 -4861
rect 1774 -4887 2352 -4861
rect 2602 -4887 2812 -4861
rect 3081 -4887 3111 -4861
rect 3176 -4887 3276 -4861
rect 3436 -4887 3536 -4861
rect 3608 -4887 3638 -4861
rect 3890 -4887 4100 -4861
rect 4350 -4887 4928 -4861
rect 5178 -4887 5388 -4861
rect 5657 -4887 5687 -4861
rect 5752 -4887 5852 -4861
rect 6012 -4887 6112 -4861
rect 6184 -4887 6214 -4861
rect 6466 -4887 6676 -4861
rect 6926 -4887 7504 -4861
rect 7754 -4887 7964 -4861
rect 8233 -4887 8263 -4861
rect 8328 -4887 8428 -4861
rect 8588 -4887 8688 -4861
rect 8760 -4887 8790 -4861
rect 9042 -4887 9252 -4861
rect 9502 -4887 10080 -4861
rect 10422 -4887 10632 -4861
rect 10809 -4887 10839 -4861
rect 10904 -4887 11004 -4861
rect 11164 -4887 11264 -4861
rect 11336 -4887 11366 -4861
rect 11710 -4887 11920 -4861
rect 13735 -4887 13765 -4861
rect 13821 -4887 13851 -4861
rect 13907 -4887 13937 -4861
rect 13993 -4887 14023 -4861
rect 14079 -4887 14109 -4861
rect 14165 -4887 14195 -4861
rect 14251 -4887 14281 -4861
rect 14337 -4887 14367 -4861
rect 14423 -4887 14453 -4861
rect 14509 -4887 14539 -4861
rect 14595 -4887 14625 -4861
rect 14681 -4887 14711 -4861
rect 14766 -4887 14796 -4861
rect 14852 -4887 14882 -4861
rect 14938 -4887 14968 -4861
rect 15024 -4887 15054 -4861
rect 15110 -4887 15140 -4861
rect 15196 -4887 15226 -4861
rect 15282 -4887 15312 -4861
rect 15368 -4887 15398 -4861
rect 15666 -4887 16612 -4861
rect -2918 -4955 -2340 -4929
rect -1538 -4955 -960 -4929
rect -802 -4955 -224 -4929
rect 26 -4955 236 -4929
rect 488 -4955 518 -4929
rect 590 -4955 690 -4929
rect 850 -4955 950 -4929
rect 1015 -4955 1045 -4929
rect 1314 -4955 1524 -4929
rect 1774 -4955 2352 -4929
rect 2602 -4955 2812 -4929
rect 3064 -4955 3094 -4929
rect 3166 -4955 3266 -4929
rect 3426 -4955 3526 -4929
rect 3591 -4955 3621 -4929
rect 3890 -4955 4100 -4929
rect 4350 -4955 4928 -4929
rect 5178 -4955 5388 -4929
rect 5640 -4955 5670 -4929
rect 5742 -4955 5842 -4929
rect 6002 -4955 6102 -4929
rect 6167 -4955 6197 -4929
rect 6466 -4955 6676 -4929
rect 6926 -4955 7504 -4929
rect 7754 -4955 7964 -4929
rect 8216 -4955 8246 -4929
rect 8318 -4955 8418 -4929
rect 8578 -4955 8678 -4929
rect 8743 -4955 8773 -4929
rect 9042 -4955 9252 -4929
rect 9502 -4955 10080 -4929
rect 10422 -4955 10632 -4929
rect 10792 -4955 10822 -4929
rect 10894 -4955 10994 -4929
rect 11154 -4955 11254 -4929
rect 11319 -4955 11349 -4929
rect 11710 -4955 11920 -4929
rect 12633 -4955 12663 -4929
rect 12719 -4955 12749 -4929
rect 12805 -4955 12835 -4929
rect 12891 -4955 12921 -4929
rect 13274 -4955 13484 -4929
rect 13735 -4955 13765 -4929
rect 13821 -4955 13851 -4929
rect 13907 -4955 13937 -4929
rect 13993 -4955 14023 -4929
rect 14079 -4955 14109 -4929
rect 14165 -4955 14195 -4929
rect 14251 -4955 14281 -4929
rect 14337 -4955 14367 -4929
rect 14423 -4955 14453 -4929
rect 14509 -4955 14539 -4929
rect 14595 -4955 14625 -4929
rect 14681 -4955 14711 -4929
rect 14766 -4955 14796 -4929
rect 14852 -4955 14882 -4929
rect 14938 -4955 14968 -4929
rect 15024 -4955 15054 -4929
rect 15110 -4955 15140 -4929
rect 15196 -4955 15226 -4929
rect 15282 -4955 15312 -4929
rect 15368 -4955 15398 -4929
rect 15666 -4955 16612 -4929
rect -2918 -5091 -2340 -5065
rect -1538 -5091 -960 -5065
rect -802 -5091 -224 -5065
rect -2918 -5113 -2646 -5091
rect -2918 -5147 -2902 -5113
rect -2868 -5147 -2799 -5113
rect -2765 -5147 -2696 -5113
rect -2662 -5147 -2646 -5113
rect -1232 -5113 -960 -5091
rect -2918 -5163 -2646 -5147
rect -2604 -5149 -2340 -5133
rect -2604 -5183 -2588 -5149
rect -2554 -5183 -2489 -5149
rect -2455 -5183 -2390 -5149
rect -2356 -5183 -2340 -5149
rect -2604 -5205 -2340 -5183
rect -2918 -5231 -2340 -5205
rect -1538 -5149 -1274 -5133
rect -1538 -5183 -1522 -5149
rect -1488 -5183 -1423 -5149
rect -1389 -5183 -1324 -5149
rect -1290 -5183 -1274 -5149
rect -1232 -5147 -1216 -5113
rect -1182 -5147 -1113 -5113
rect -1079 -5147 -1010 -5113
rect -976 -5147 -960 -5113
rect -496 -5113 -224 -5091
rect 26 -5091 236 -5065
rect 26 -5097 110 -5091
rect -1232 -5163 -960 -5147
rect -802 -5149 -538 -5133
rect -1538 -5205 -1274 -5183
rect -802 -5183 -786 -5149
rect -752 -5183 -687 -5149
rect -653 -5183 -588 -5149
rect -554 -5183 -538 -5149
rect -496 -5147 -480 -5113
rect -446 -5147 -377 -5113
rect -343 -5147 -274 -5113
rect -240 -5147 -224 -5113
rect -496 -5163 -224 -5147
rect -32 -5113 110 -5097
rect 488 -5111 518 -5039
rect -32 -5147 -16 -5113
rect 18 -5147 110 -5113
rect 448 -5123 518 -5111
rect 590 -5113 690 -5085
rect 850 -5113 950 -5085
rect 1015 -5107 1045 -5039
rect 1314 -5091 1524 -5065
rect 1774 -5091 2352 -5065
rect 2602 -5091 2812 -5065
rect 1314 -5097 1398 -5091
rect -32 -5163 110 -5147
rect 152 -5149 294 -5133
rect -802 -5205 -538 -5183
rect 152 -5183 244 -5149
rect 278 -5183 294 -5149
rect 448 -5157 464 -5123
rect 498 -5157 518 -5123
rect 448 -5170 518 -5157
rect 568 -5123 690 -5113
rect 568 -5157 584 -5123
rect 618 -5157 690 -5123
rect 568 -5167 690 -5157
rect 789 -5123 950 -5113
rect 789 -5157 805 -5123
rect 839 -5157 950 -5123
rect 789 -5167 950 -5157
rect 152 -5199 294 -5183
rect 152 -5205 236 -5199
rect 488 -5205 518 -5170
rect -1538 -5231 -960 -5205
rect -802 -5231 -224 -5205
rect 26 -5231 236 -5205
rect 590 -5241 690 -5167
rect 850 -5241 950 -5167
rect 995 -5123 1049 -5107
rect 995 -5157 1005 -5123
rect 1039 -5157 1049 -5123
rect 995 -5173 1049 -5157
rect 1256 -5113 1398 -5097
rect 1256 -5147 1272 -5113
rect 1306 -5147 1398 -5113
rect 1774 -5113 2046 -5091
rect 2602 -5097 2686 -5091
rect 1256 -5163 1398 -5147
rect 1440 -5149 1582 -5133
rect 1015 -5205 1045 -5173
rect 1440 -5183 1532 -5149
rect 1566 -5183 1582 -5149
rect 1774 -5147 1790 -5113
rect 1824 -5147 1893 -5113
rect 1927 -5147 1996 -5113
rect 2030 -5147 2046 -5113
rect 2544 -5113 2686 -5097
rect 3064 -5111 3094 -5039
rect 1774 -5163 2046 -5147
rect 2088 -5149 2352 -5133
rect 1440 -5199 1582 -5183
rect 2088 -5183 2104 -5149
rect 2138 -5183 2203 -5149
rect 2237 -5183 2302 -5149
rect 2336 -5183 2352 -5149
rect 2544 -5147 2560 -5113
rect 2594 -5147 2686 -5113
rect 3024 -5123 3094 -5111
rect 3166 -5113 3266 -5085
rect 3426 -5113 3526 -5085
rect 3591 -5107 3621 -5039
rect 3890 -5091 4100 -5065
rect 4350 -5091 4928 -5065
rect 5178 -5091 5388 -5065
rect 3890 -5097 3974 -5091
rect 2544 -5163 2686 -5147
rect 2728 -5149 2870 -5133
rect 1440 -5205 1524 -5199
rect 2088 -5205 2352 -5183
rect 2728 -5183 2820 -5149
rect 2854 -5183 2870 -5149
rect 3024 -5157 3040 -5123
rect 3074 -5157 3094 -5123
rect 3024 -5170 3094 -5157
rect 3144 -5123 3266 -5113
rect 3144 -5157 3160 -5123
rect 3194 -5157 3266 -5123
rect 3144 -5167 3266 -5157
rect 3365 -5123 3526 -5113
rect 3365 -5157 3381 -5123
rect 3415 -5157 3526 -5123
rect 3365 -5167 3526 -5157
rect 2728 -5199 2870 -5183
rect 2728 -5205 2812 -5199
rect 3064 -5205 3094 -5170
rect 1314 -5231 1524 -5205
rect 1774 -5231 2352 -5205
rect 2602 -5231 2812 -5205
rect 3166 -5241 3266 -5167
rect 3426 -5241 3526 -5167
rect 3571 -5123 3625 -5107
rect 3571 -5157 3581 -5123
rect 3615 -5157 3625 -5123
rect 3571 -5173 3625 -5157
rect 3832 -5113 3974 -5097
rect 3832 -5147 3848 -5113
rect 3882 -5147 3974 -5113
rect 4350 -5113 4622 -5091
rect 5178 -5097 5262 -5091
rect 3832 -5163 3974 -5147
rect 4016 -5149 4158 -5133
rect 3591 -5205 3621 -5173
rect 4016 -5183 4108 -5149
rect 4142 -5183 4158 -5149
rect 4350 -5147 4366 -5113
rect 4400 -5147 4469 -5113
rect 4503 -5147 4572 -5113
rect 4606 -5147 4622 -5113
rect 5120 -5113 5262 -5097
rect 5640 -5111 5670 -5039
rect 4350 -5163 4622 -5147
rect 4664 -5149 4928 -5133
rect 4016 -5199 4158 -5183
rect 4664 -5183 4680 -5149
rect 4714 -5183 4779 -5149
rect 4813 -5183 4878 -5149
rect 4912 -5183 4928 -5149
rect 5120 -5147 5136 -5113
rect 5170 -5147 5262 -5113
rect 5600 -5123 5670 -5111
rect 5742 -5113 5842 -5085
rect 6002 -5113 6102 -5085
rect 6167 -5107 6197 -5039
rect 6466 -5091 6676 -5065
rect 6926 -5091 7504 -5065
rect 7754 -5091 7964 -5065
rect 6466 -5097 6550 -5091
rect 5120 -5163 5262 -5147
rect 5304 -5149 5446 -5133
rect 4016 -5205 4100 -5199
rect 4664 -5205 4928 -5183
rect 5304 -5183 5396 -5149
rect 5430 -5183 5446 -5149
rect 5600 -5157 5616 -5123
rect 5650 -5157 5670 -5123
rect 5600 -5170 5670 -5157
rect 5720 -5123 5842 -5113
rect 5720 -5157 5736 -5123
rect 5770 -5157 5842 -5123
rect 5720 -5167 5842 -5157
rect 5941 -5123 6102 -5113
rect 5941 -5157 5957 -5123
rect 5991 -5157 6102 -5123
rect 5941 -5167 6102 -5157
rect 5304 -5199 5446 -5183
rect 5304 -5205 5388 -5199
rect 5640 -5205 5670 -5170
rect 3890 -5231 4100 -5205
rect 4350 -5231 4928 -5205
rect 5178 -5231 5388 -5205
rect 5742 -5241 5842 -5167
rect 6002 -5241 6102 -5167
rect 6147 -5123 6201 -5107
rect 6147 -5157 6157 -5123
rect 6191 -5157 6201 -5123
rect 6147 -5173 6201 -5157
rect 6408 -5113 6550 -5097
rect 6408 -5147 6424 -5113
rect 6458 -5147 6550 -5113
rect 6926 -5113 7198 -5091
rect 7754 -5097 7838 -5091
rect 6408 -5163 6550 -5147
rect 6592 -5149 6734 -5133
rect 6167 -5205 6197 -5173
rect 6592 -5183 6684 -5149
rect 6718 -5183 6734 -5149
rect 6926 -5147 6942 -5113
rect 6976 -5147 7045 -5113
rect 7079 -5147 7148 -5113
rect 7182 -5147 7198 -5113
rect 7696 -5113 7838 -5097
rect 8216 -5111 8246 -5039
rect 6926 -5163 7198 -5147
rect 7240 -5149 7504 -5133
rect 6592 -5199 6734 -5183
rect 7240 -5183 7256 -5149
rect 7290 -5183 7355 -5149
rect 7389 -5183 7454 -5149
rect 7488 -5183 7504 -5149
rect 7696 -5147 7712 -5113
rect 7746 -5147 7838 -5113
rect 8176 -5123 8246 -5111
rect 8318 -5113 8418 -5085
rect 8578 -5113 8678 -5085
rect 8743 -5107 8773 -5039
rect 9042 -5091 9252 -5065
rect 9502 -5091 10080 -5065
rect 10422 -5091 10632 -5065
rect 9042 -5097 9126 -5091
rect 7696 -5163 7838 -5147
rect 7880 -5149 8022 -5133
rect 6592 -5205 6676 -5199
rect 7240 -5205 7504 -5183
rect 7880 -5183 7972 -5149
rect 8006 -5183 8022 -5149
rect 8176 -5157 8192 -5123
rect 8226 -5157 8246 -5123
rect 8176 -5170 8246 -5157
rect 8296 -5123 8418 -5113
rect 8296 -5157 8312 -5123
rect 8346 -5157 8418 -5123
rect 8296 -5167 8418 -5157
rect 8517 -5123 8678 -5113
rect 8517 -5157 8533 -5123
rect 8567 -5157 8678 -5123
rect 8517 -5167 8678 -5157
rect 7880 -5199 8022 -5183
rect 7880 -5205 7964 -5199
rect 8216 -5205 8246 -5170
rect 6466 -5231 6676 -5205
rect 6926 -5231 7504 -5205
rect 7754 -5231 7964 -5205
rect 8318 -5241 8418 -5167
rect 8578 -5241 8678 -5167
rect 8723 -5123 8777 -5107
rect 8723 -5157 8733 -5123
rect 8767 -5157 8777 -5123
rect 8723 -5173 8777 -5157
rect 8984 -5113 9126 -5097
rect 8984 -5147 9000 -5113
rect 9034 -5147 9126 -5113
rect 9502 -5113 9774 -5091
rect 10422 -5097 10506 -5091
rect 8984 -5163 9126 -5147
rect 9168 -5149 9310 -5133
rect 8743 -5205 8773 -5173
rect 9168 -5183 9260 -5149
rect 9294 -5183 9310 -5149
rect 9502 -5147 9518 -5113
rect 9552 -5147 9621 -5113
rect 9655 -5147 9724 -5113
rect 9758 -5147 9774 -5113
rect 10364 -5113 10506 -5097
rect 10792 -5111 10822 -5039
rect 9502 -5163 9774 -5147
rect 9816 -5149 10080 -5133
rect 9168 -5199 9310 -5183
rect 9816 -5183 9832 -5149
rect 9866 -5183 9931 -5149
rect 9965 -5183 10030 -5149
rect 10064 -5183 10080 -5149
rect 10364 -5147 10380 -5113
rect 10414 -5147 10506 -5113
rect 10752 -5123 10822 -5111
rect 10894 -5113 10994 -5085
rect 11154 -5113 11254 -5085
rect 11319 -5107 11349 -5039
rect 11710 -5091 11920 -5065
rect 11710 -5097 11794 -5091
rect 10364 -5163 10506 -5147
rect 10548 -5149 10690 -5133
rect 9168 -5205 9252 -5199
rect 9816 -5205 10080 -5183
rect 10548 -5183 10640 -5149
rect 10674 -5183 10690 -5149
rect 10752 -5157 10768 -5123
rect 10802 -5157 10822 -5123
rect 10752 -5170 10822 -5157
rect 10872 -5123 10994 -5113
rect 10872 -5157 10888 -5123
rect 10922 -5157 10994 -5123
rect 10872 -5167 10994 -5157
rect 11093 -5123 11254 -5113
rect 11093 -5157 11109 -5123
rect 11143 -5157 11254 -5123
rect 11093 -5167 11254 -5157
rect 10548 -5199 10690 -5183
rect 10548 -5205 10632 -5199
rect 10792 -5205 10822 -5170
rect 9042 -5231 9252 -5205
rect 9502 -5231 10080 -5205
rect 10422 -5231 10632 -5205
rect 10894 -5241 10994 -5167
rect 11154 -5241 11254 -5167
rect 11299 -5123 11353 -5107
rect 11299 -5157 11309 -5123
rect 11343 -5157 11353 -5123
rect 11299 -5173 11353 -5157
rect 11652 -5113 11794 -5097
rect 12633 -5113 12663 -5039
rect 12719 -5113 12749 -5039
rect 12805 -5113 12835 -5039
rect 12891 -5113 12921 -5039
rect 13274 -5091 13484 -5065
rect 13735 -5088 13765 -5039
rect 13821 -5088 13851 -5039
rect 13907 -5088 13937 -5039
rect 13993 -5088 14023 -5039
rect 13400 -5097 13484 -5091
rect 13400 -5113 13542 -5097
rect 11652 -5147 11668 -5113
rect 11702 -5147 11794 -5113
rect 12547 -5123 13007 -5113
rect 11652 -5163 11794 -5147
rect 11836 -5149 11978 -5133
rect 11319 -5205 11349 -5173
rect 11836 -5183 11928 -5149
rect 11962 -5183 11978 -5149
rect 11836 -5199 11978 -5183
rect 12547 -5157 12574 -5123
rect 12608 -5157 12642 -5123
rect 12676 -5157 12710 -5123
rect 12744 -5157 12778 -5123
rect 12812 -5157 12846 -5123
rect 12880 -5157 12914 -5123
rect 12948 -5157 13007 -5123
rect 12547 -5167 13007 -5157
rect 11836 -5205 11920 -5199
rect 12547 -5205 12577 -5167
rect 12633 -5205 12663 -5167
rect 12719 -5205 12749 -5167
rect 12805 -5205 12835 -5167
rect 12891 -5205 12921 -5167
rect 12977 -5205 13007 -5167
rect 13216 -5149 13358 -5133
rect 13216 -5183 13232 -5149
rect 13266 -5183 13358 -5149
rect 13400 -5147 13492 -5113
rect 13526 -5147 13542 -5113
rect 13400 -5163 13542 -5147
rect 13676 -5123 14023 -5088
rect 13676 -5157 13692 -5123
rect 13726 -5157 14023 -5123
rect 13216 -5199 13358 -5183
rect 13676 -5190 14023 -5157
rect 13274 -5205 13358 -5199
rect 13735 -5205 13765 -5190
rect 13821 -5205 13851 -5190
rect 13907 -5205 13937 -5190
rect 13993 -5205 14023 -5190
rect 14079 -5098 14109 -5039
rect 14165 -5098 14195 -5039
rect 14251 -5098 14281 -5039
rect 14337 -5098 14367 -5039
rect 14423 -5098 14453 -5039
rect 14509 -5098 14539 -5039
rect 14595 -5098 14625 -5039
rect 14681 -5098 14711 -5039
rect 14766 -5098 14796 -5039
rect 14852 -5098 14882 -5039
rect 14938 -5098 14968 -5039
rect 15024 -5098 15054 -5039
rect 15110 -5098 15140 -5039
rect 15196 -5098 15226 -5039
rect 15282 -5098 15312 -5039
rect 15368 -5098 15398 -5039
rect 15666 -5091 16612 -5065
rect 14079 -5123 15398 -5098
rect 14079 -5157 14119 -5123
rect 14153 -5157 14187 -5123
rect 14221 -5157 14255 -5123
rect 14289 -5157 14323 -5123
rect 14357 -5157 14391 -5123
rect 14425 -5157 14459 -5123
rect 14493 -5157 14527 -5123
rect 14561 -5157 14595 -5123
rect 14629 -5157 14663 -5123
rect 14697 -5157 14731 -5123
rect 14765 -5157 14799 -5123
rect 14833 -5157 14867 -5123
rect 14901 -5157 14935 -5123
rect 14969 -5157 15003 -5123
rect 15037 -5157 15071 -5123
rect 15105 -5157 15139 -5123
rect 15173 -5157 15398 -5123
rect 16158 -5113 16612 -5091
rect 14079 -5173 15398 -5157
rect 14079 -5205 14109 -5173
rect 14165 -5205 14195 -5173
rect 14251 -5205 14281 -5173
rect 14337 -5205 14367 -5173
rect 14423 -5205 14453 -5173
rect 14509 -5205 14539 -5173
rect 14595 -5205 14625 -5173
rect 14681 -5205 14711 -5173
rect 14766 -5205 14796 -5173
rect 14852 -5205 14882 -5173
rect 14938 -5205 14968 -5173
rect 15024 -5205 15054 -5173
rect 15110 -5205 15140 -5173
rect 15196 -5205 15226 -5173
rect 15282 -5205 15312 -5173
rect 15368 -5205 15398 -5173
rect 15666 -5149 16116 -5133
rect 15666 -5183 15682 -5149
rect 15716 -5183 15810 -5149
rect 15844 -5183 15938 -5149
rect 15972 -5183 16066 -5149
rect 16100 -5183 16116 -5149
rect 16158 -5147 16174 -5113
rect 16208 -5147 16302 -5113
rect 16336 -5147 16430 -5113
rect 16464 -5147 16558 -5113
rect 16592 -5147 16612 -5113
rect 16158 -5163 16612 -5147
rect 15666 -5205 16116 -5183
rect 11710 -5231 11920 -5205
rect 13274 -5231 13484 -5205
rect 15666 -5231 16612 -5205
rect -2918 -5431 -2340 -5405
rect -1538 -5431 -960 -5405
rect -802 -5431 -224 -5405
rect 26 -5431 236 -5405
rect 488 -5431 518 -5405
rect 590 -5431 690 -5405
rect 850 -5431 950 -5405
rect 1015 -5431 1045 -5405
rect 1314 -5431 1524 -5405
rect 1774 -5431 2352 -5405
rect 2602 -5431 2812 -5405
rect 3064 -5431 3094 -5405
rect 3166 -5431 3266 -5405
rect 3426 -5431 3526 -5405
rect 3591 -5431 3621 -5405
rect 3890 -5431 4100 -5405
rect 4350 -5431 4928 -5405
rect 5178 -5431 5388 -5405
rect 5640 -5431 5670 -5405
rect 5742 -5431 5842 -5405
rect 6002 -5431 6102 -5405
rect 6167 -5431 6197 -5405
rect 6466 -5431 6676 -5405
rect 6926 -5431 7504 -5405
rect 7754 -5431 7964 -5405
rect 8216 -5431 8246 -5405
rect 8318 -5431 8418 -5405
rect 8578 -5431 8678 -5405
rect 8743 -5431 8773 -5405
rect 9042 -5431 9252 -5405
rect 9502 -5431 10080 -5405
rect 10422 -5431 10632 -5405
rect 10792 -5431 10822 -5405
rect 10894 -5431 10994 -5405
rect 11154 -5431 11254 -5405
rect 11319 -5431 11349 -5405
rect 11710 -5431 11920 -5405
rect 12547 -5431 12577 -5405
rect 12633 -5431 12663 -5405
rect 12719 -5431 12749 -5405
rect 12805 -5431 12835 -5405
rect 12891 -5431 12921 -5405
rect 12977 -5431 13007 -5405
rect 13274 -5431 13484 -5405
rect 13735 -5431 13765 -5405
rect 13821 -5431 13851 -5405
rect 13907 -5431 13937 -5405
rect 13993 -5431 14023 -5405
rect 14079 -5431 14109 -5405
rect 14165 -5431 14195 -5405
rect 14251 -5431 14281 -5405
rect 14337 -5431 14367 -5405
rect 14423 -5431 14453 -5405
rect 14509 -5431 14539 -5405
rect 14595 -5431 14625 -5405
rect 14681 -5431 14711 -5405
rect 14766 -5431 14796 -5405
rect 14852 -5431 14882 -5405
rect 14938 -5431 14968 -5405
rect 15024 -5431 15054 -5405
rect 15110 -5431 15140 -5405
rect 15196 -5431 15226 -5405
rect 15282 -5431 15312 -5405
rect 15368 -5431 15398 -5405
rect 15666 -5431 16612 -5405
rect -2918 -5499 -2340 -5473
rect -1538 -5499 -960 -5473
rect -802 -5499 -224 -5473
rect 26 -5499 236 -5473
rect 505 -5499 535 -5473
rect 600 -5499 700 -5473
rect 860 -5499 960 -5473
rect 1032 -5499 1062 -5473
rect 1314 -5499 1524 -5473
rect 1774 -5499 2352 -5473
rect 2602 -5499 2812 -5473
rect 3081 -5499 3111 -5473
rect 3176 -5499 3276 -5473
rect 3436 -5499 3536 -5473
rect 3608 -5499 3638 -5473
rect 3890 -5499 4100 -5473
rect 4350 -5499 4928 -5473
rect 5178 -5499 5388 -5473
rect 5657 -5499 5687 -5473
rect 5752 -5499 5852 -5473
rect 6012 -5499 6112 -5473
rect 6184 -5499 6214 -5473
rect 6466 -5499 6676 -5473
rect 6926 -5499 7504 -5473
rect 7754 -5499 7964 -5473
rect 8233 -5499 8263 -5473
rect 8328 -5499 8428 -5473
rect 8588 -5499 8688 -5473
rect 8760 -5499 8790 -5473
rect 9042 -5499 9252 -5473
rect 9502 -5499 10080 -5473
rect 10422 -5499 10632 -5473
rect 10809 -5499 10839 -5473
rect 10904 -5499 11004 -5473
rect 11164 -5499 11264 -5473
rect 11336 -5499 11366 -5473
rect 11710 -5499 11920 -5473
rect 13735 -5499 13765 -5473
rect 13821 -5499 13851 -5473
rect 13907 -5499 13937 -5473
rect 13993 -5499 14023 -5473
rect 14079 -5499 14109 -5473
rect 14165 -5499 14195 -5473
rect 14251 -5499 14281 -5473
rect 14337 -5499 14367 -5473
rect 14423 -5499 14453 -5473
rect 14509 -5499 14539 -5473
rect 14595 -5499 14625 -5473
rect 14681 -5499 14711 -5473
rect 14766 -5499 14796 -5473
rect 14852 -5499 14882 -5473
rect 14938 -5499 14968 -5473
rect 15024 -5499 15054 -5473
rect 15110 -5499 15140 -5473
rect 15196 -5499 15226 -5473
rect 15282 -5499 15312 -5473
rect 15368 -5499 15398 -5473
rect 15666 -5499 16612 -5473
rect -2918 -5699 -2340 -5673
rect -1538 -5699 -960 -5673
rect -802 -5699 -224 -5673
rect 26 -5699 236 -5673
rect -2918 -5721 -2654 -5699
rect -2918 -5755 -2902 -5721
rect -2868 -5755 -2803 -5721
rect -2769 -5755 -2704 -5721
rect -2670 -5755 -2654 -5721
rect -1224 -5721 -960 -5699
rect -2918 -5771 -2654 -5755
rect -2612 -5757 -2340 -5741
rect -2612 -5791 -2596 -5757
rect -2562 -5791 -2493 -5757
rect -2459 -5791 -2390 -5757
rect -2356 -5791 -2340 -5757
rect -2612 -5813 -2340 -5791
rect -2918 -5839 -2340 -5813
rect -1538 -5757 -1266 -5741
rect -1538 -5791 -1522 -5757
rect -1488 -5791 -1419 -5757
rect -1385 -5791 -1316 -5757
rect -1282 -5791 -1266 -5757
rect -1224 -5755 -1208 -5721
rect -1174 -5755 -1109 -5721
rect -1075 -5755 -1010 -5721
rect -976 -5755 -960 -5721
rect -488 -5721 -224 -5699
rect -1224 -5771 -960 -5755
rect -802 -5757 -530 -5741
rect -1538 -5813 -1266 -5791
rect -802 -5791 -786 -5757
rect -752 -5791 -683 -5757
rect -649 -5791 -580 -5757
rect -546 -5791 -530 -5757
rect -488 -5755 -472 -5721
rect -438 -5755 -373 -5721
rect -339 -5755 -274 -5721
rect -240 -5755 -224 -5721
rect 152 -5705 236 -5699
rect 152 -5721 294 -5705
rect -488 -5771 -224 -5755
rect -32 -5757 110 -5741
rect -802 -5813 -530 -5791
rect -32 -5791 -16 -5757
rect 18 -5791 110 -5757
rect 152 -5755 244 -5721
rect 278 -5755 294 -5721
rect 505 -5731 535 -5699
rect 152 -5771 294 -5755
rect 501 -5747 555 -5731
rect -32 -5807 110 -5791
rect 501 -5781 511 -5747
rect 545 -5781 555 -5747
rect 501 -5797 555 -5781
rect 600 -5737 700 -5663
rect 860 -5737 960 -5663
rect 1314 -5699 1524 -5673
rect 1032 -5734 1062 -5699
rect 1440 -5705 1524 -5699
rect 1774 -5699 2352 -5673
rect 2602 -5699 2812 -5673
rect 1440 -5721 1582 -5705
rect 600 -5747 761 -5737
rect 600 -5781 711 -5747
rect 745 -5781 761 -5747
rect 600 -5791 761 -5781
rect 860 -5747 982 -5737
rect 860 -5781 932 -5747
rect 966 -5781 982 -5747
rect 860 -5791 982 -5781
rect 1032 -5747 1102 -5734
rect 1032 -5781 1052 -5747
rect 1086 -5781 1102 -5747
rect 26 -5813 110 -5807
rect -1538 -5839 -960 -5813
rect -802 -5839 -224 -5813
rect 26 -5839 236 -5813
rect 505 -5865 535 -5797
rect 600 -5819 700 -5791
rect 860 -5819 960 -5791
rect 1032 -5793 1102 -5781
rect 1256 -5757 1398 -5741
rect 1256 -5791 1272 -5757
rect 1306 -5791 1398 -5757
rect 1440 -5755 1532 -5721
rect 1566 -5755 1582 -5721
rect 1440 -5771 1582 -5755
rect 1774 -5721 2038 -5699
rect 1774 -5755 1790 -5721
rect 1824 -5755 1889 -5721
rect 1923 -5755 1988 -5721
rect 2022 -5755 2038 -5721
rect 2728 -5705 2812 -5699
rect 2728 -5721 2870 -5705
rect 1774 -5771 2038 -5755
rect 2080 -5757 2352 -5741
rect 1032 -5865 1062 -5793
rect 1256 -5807 1398 -5791
rect 1314 -5813 1398 -5807
rect 2080 -5791 2096 -5757
rect 2130 -5791 2199 -5757
rect 2233 -5791 2302 -5757
rect 2336 -5791 2352 -5757
rect 2080 -5813 2352 -5791
rect 2544 -5757 2686 -5741
rect 2544 -5791 2560 -5757
rect 2594 -5791 2686 -5757
rect 2728 -5755 2820 -5721
rect 2854 -5755 2870 -5721
rect 3081 -5731 3111 -5699
rect 2728 -5771 2870 -5755
rect 3077 -5747 3131 -5731
rect 2544 -5807 2686 -5791
rect 3077 -5781 3087 -5747
rect 3121 -5781 3131 -5747
rect 3077 -5797 3131 -5781
rect 3176 -5737 3276 -5663
rect 3436 -5737 3536 -5663
rect 3890 -5699 4100 -5673
rect 3608 -5734 3638 -5699
rect 4016 -5705 4100 -5699
rect 4350 -5699 4928 -5673
rect 5178 -5699 5388 -5673
rect 4016 -5721 4158 -5705
rect 3176 -5747 3337 -5737
rect 3176 -5781 3287 -5747
rect 3321 -5781 3337 -5747
rect 3176 -5791 3337 -5781
rect 3436 -5747 3558 -5737
rect 3436 -5781 3508 -5747
rect 3542 -5781 3558 -5747
rect 3436 -5791 3558 -5781
rect 3608 -5747 3678 -5734
rect 3608 -5781 3628 -5747
rect 3662 -5781 3678 -5747
rect 1314 -5839 1524 -5813
rect 1774 -5839 2352 -5813
rect 2602 -5813 2686 -5807
rect 2602 -5839 2812 -5813
rect 3081 -5865 3111 -5797
rect 3176 -5819 3276 -5791
rect 3436 -5819 3536 -5791
rect 3608 -5793 3678 -5781
rect 3832 -5757 3974 -5741
rect 3832 -5791 3848 -5757
rect 3882 -5791 3974 -5757
rect 4016 -5755 4108 -5721
rect 4142 -5755 4158 -5721
rect 4016 -5771 4158 -5755
rect 4350 -5721 4614 -5699
rect 4350 -5755 4366 -5721
rect 4400 -5755 4465 -5721
rect 4499 -5755 4564 -5721
rect 4598 -5755 4614 -5721
rect 5304 -5705 5388 -5699
rect 5304 -5721 5446 -5705
rect 4350 -5771 4614 -5755
rect 4656 -5757 4928 -5741
rect 3608 -5865 3638 -5793
rect 3832 -5807 3974 -5791
rect 3890 -5813 3974 -5807
rect 4656 -5791 4672 -5757
rect 4706 -5791 4775 -5757
rect 4809 -5791 4878 -5757
rect 4912 -5791 4928 -5757
rect 4656 -5813 4928 -5791
rect 5120 -5757 5262 -5741
rect 5120 -5791 5136 -5757
rect 5170 -5791 5262 -5757
rect 5304 -5755 5396 -5721
rect 5430 -5755 5446 -5721
rect 5657 -5731 5687 -5699
rect 5304 -5771 5446 -5755
rect 5653 -5747 5707 -5731
rect 5120 -5807 5262 -5791
rect 5653 -5781 5663 -5747
rect 5697 -5781 5707 -5747
rect 5653 -5797 5707 -5781
rect 5752 -5737 5852 -5663
rect 6012 -5737 6112 -5663
rect 6466 -5699 6676 -5673
rect 6184 -5734 6214 -5699
rect 6592 -5705 6676 -5699
rect 6926 -5699 7504 -5673
rect 7754 -5699 7964 -5673
rect 6592 -5721 6734 -5705
rect 5752 -5747 5913 -5737
rect 5752 -5781 5863 -5747
rect 5897 -5781 5913 -5747
rect 5752 -5791 5913 -5781
rect 6012 -5747 6134 -5737
rect 6012 -5781 6084 -5747
rect 6118 -5781 6134 -5747
rect 6012 -5791 6134 -5781
rect 6184 -5747 6254 -5734
rect 6184 -5781 6204 -5747
rect 6238 -5781 6254 -5747
rect 3890 -5839 4100 -5813
rect 4350 -5839 4928 -5813
rect 5178 -5813 5262 -5807
rect 5178 -5839 5388 -5813
rect 5657 -5865 5687 -5797
rect 5752 -5819 5852 -5791
rect 6012 -5819 6112 -5791
rect 6184 -5793 6254 -5781
rect 6408 -5757 6550 -5741
rect 6408 -5791 6424 -5757
rect 6458 -5791 6550 -5757
rect 6592 -5755 6684 -5721
rect 6718 -5755 6734 -5721
rect 6592 -5771 6734 -5755
rect 6926 -5721 7190 -5699
rect 6926 -5755 6942 -5721
rect 6976 -5755 7041 -5721
rect 7075 -5755 7140 -5721
rect 7174 -5755 7190 -5721
rect 7880 -5705 7964 -5699
rect 7880 -5721 8022 -5705
rect 6926 -5771 7190 -5755
rect 7232 -5757 7504 -5741
rect 6184 -5865 6214 -5793
rect 6408 -5807 6550 -5791
rect 6466 -5813 6550 -5807
rect 7232 -5791 7248 -5757
rect 7282 -5791 7351 -5757
rect 7385 -5791 7454 -5757
rect 7488 -5791 7504 -5757
rect 7232 -5813 7504 -5791
rect 7696 -5757 7838 -5741
rect 7696 -5791 7712 -5757
rect 7746 -5791 7838 -5757
rect 7880 -5755 7972 -5721
rect 8006 -5755 8022 -5721
rect 8233 -5731 8263 -5699
rect 7880 -5771 8022 -5755
rect 8229 -5747 8283 -5731
rect 7696 -5807 7838 -5791
rect 8229 -5781 8239 -5747
rect 8273 -5781 8283 -5747
rect 8229 -5797 8283 -5781
rect 8328 -5737 8428 -5663
rect 8588 -5737 8688 -5663
rect 9042 -5699 9252 -5673
rect 8760 -5734 8790 -5699
rect 9168 -5705 9252 -5699
rect 9502 -5699 10080 -5673
rect 10422 -5699 10632 -5673
rect 9168 -5721 9310 -5705
rect 8328 -5747 8489 -5737
rect 8328 -5781 8439 -5747
rect 8473 -5781 8489 -5747
rect 8328 -5791 8489 -5781
rect 8588 -5747 8710 -5737
rect 8588 -5781 8660 -5747
rect 8694 -5781 8710 -5747
rect 8588 -5791 8710 -5781
rect 8760 -5747 8830 -5734
rect 8760 -5781 8780 -5747
rect 8814 -5781 8830 -5747
rect 6466 -5839 6676 -5813
rect 6926 -5839 7504 -5813
rect 7754 -5813 7838 -5807
rect 7754 -5839 7964 -5813
rect 8233 -5865 8263 -5797
rect 8328 -5819 8428 -5791
rect 8588 -5819 8688 -5791
rect 8760 -5793 8830 -5781
rect 8984 -5757 9126 -5741
rect 8984 -5791 9000 -5757
rect 9034 -5791 9126 -5757
rect 9168 -5755 9260 -5721
rect 9294 -5755 9310 -5721
rect 9168 -5771 9310 -5755
rect 9502 -5721 9766 -5699
rect 9502 -5755 9518 -5721
rect 9552 -5755 9617 -5721
rect 9651 -5755 9716 -5721
rect 9750 -5755 9766 -5721
rect 10548 -5705 10632 -5699
rect 10548 -5721 10690 -5705
rect 9502 -5771 9766 -5755
rect 9808 -5757 10080 -5741
rect 8760 -5865 8790 -5793
rect 8984 -5807 9126 -5791
rect 9042 -5813 9126 -5807
rect 9808 -5791 9824 -5757
rect 9858 -5791 9927 -5757
rect 9961 -5791 10030 -5757
rect 10064 -5791 10080 -5757
rect 9808 -5813 10080 -5791
rect 10364 -5757 10506 -5741
rect 10364 -5791 10380 -5757
rect 10414 -5791 10506 -5757
rect 10548 -5755 10640 -5721
rect 10674 -5755 10690 -5721
rect 10809 -5731 10839 -5699
rect 10548 -5771 10690 -5755
rect 10805 -5747 10859 -5731
rect 10364 -5807 10506 -5791
rect 10805 -5781 10815 -5747
rect 10849 -5781 10859 -5747
rect 10805 -5797 10859 -5781
rect 10904 -5737 11004 -5663
rect 11164 -5737 11264 -5663
rect 11710 -5699 11920 -5673
rect 15666 -5699 16612 -5673
rect 11336 -5734 11366 -5699
rect 11836 -5705 11920 -5699
rect 11836 -5721 11978 -5705
rect 13735 -5714 13765 -5699
rect 13821 -5714 13851 -5699
rect 13907 -5714 13937 -5699
rect 13993 -5714 14023 -5699
rect 10904 -5747 11065 -5737
rect 10904 -5781 11015 -5747
rect 11049 -5781 11065 -5747
rect 10904 -5791 11065 -5781
rect 11164 -5747 11286 -5737
rect 11164 -5781 11236 -5747
rect 11270 -5781 11286 -5747
rect 11164 -5791 11286 -5781
rect 11336 -5747 11406 -5734
rect 11336 -5781 11356 -5747
rect 11390 -5781 11406 -5747
rect 9042 -5839 9252 -5813
rect 9502 -5839 10080 -5813
rect 10422 -5813 10506 -5807
rect 10422 -5839 10632 -5813
rect 10809 -5865 10839 -5797
rect 10904 -5819 11004 -5791
rect 11164 -5819 11264 -5791
rect 11336 -5793 11406 -5781
rect 11652 -5757 11794 -5741
rect 11652 -5791 11668 -5757
rect 11702 -5791 11794 -5757
rect 11836 -5755 11928 -5721
rect 11962 -5755 11978 -5721
rect 11836 -5771 11978 -5755
rect 13676 -5747 14023 -5714
rect 11336 -5865 11366 -5793
rect 11652 -5807 11794 -5791
rect 11710 -5813 11794 -5807
rect 13676 -5781 13692 -5747
rect 13726 -5781 14023 -5747
rect 11710 -5839 11920 -5813
rect 13676 -5816 14023 -5781
rect 13735 -5865 13765 -5816
rect 13821 -5865 13851 -5816
rect 13907 -5865 13937 -5816
rect 13993 -5865 14023 -5816
rect 14079 -5731 14109 -5699
rect 14165 -5731 14195 -5699
rect 14251 -5731 14281 -5699
rect 14337 -5731 14367 -5699
rect 14423 -5731 14453 -5699
rect 14509 -5731 14539 -5699
rect 14595 -5731 14625 -5699
rect 14681 -5731 14711 -5699
rect 14766 -5731 14796 -5699
rect 14852 -5731 14882 -5699
rect 14938 -5731 14968 -5699
rect 15024 -5731 15054 -5699
rect 15110 -5731 15140 -5699
rect 15196 -5731 15226 -5699
rect 15282 -5731 15312 -5699
rect 15368 -5731 15398 -5699
rect 14079 -5747 15398 -5731
rect 16162 -5721 16612 -5699
rect 14079 -5781 14119 -5747
rect 14153 -5781 14187 -5747
rect 14221 -5781 14255 -5747
rect 14289 -5781 14323 -5747
rect 14357 -5781 14391 -5747
rect 14425 -5781 14459 -5747
rect 14493 -5781 14527 -5747
rect 14561 -5781 14595 -5747
rect 14629 -5781 14663 -5747
rect 14697 -5781 14731 -5747
rect 14765 -5781 14799 -5747
rect 14833 -5781 14867 -5747
rect 14901 -5781 14935 -5747
rect 14969 -5781 15003 -5747
rect 15037 -5781 15071 -5747
rect 15105 -5781 15139 -5747
rect 15173 -5781 15398 -5747
rect 14079 -5806 15398 -5781
rect 14079 -5865 14109 -5806
rect 14165 -5865 14195 -5806
rect 14251 -5865 14281 -5806
rect 14337 -5865 14367 -5806
rect 14423 -5865 14453 -5806
rect 14509 -5865 14539 -5806
rect 14595 -5865 14625 -5806
rect 14681 -5865 14711 -5806
rect 14766 -5865 14796 -5806
rect 14852 -5865 14882 -5806
rect 14938 -5865 14968 -5806
rect 15024 -5865 15054 -5806
rect 15110 -5865 15140 -5806
rect 15196 -5865 15226 -5806
rect 15282 -5865 15312 -5806
rect 15368 -5865 15398 -5806
rect 15666 -5757 16120 -5741
rect 15666 -5791 15686 -5757
rect 15720 -5791 15814 -5757
rect 15848 -5791 15942 -5757
rect 15976 -5791 16070 -5757
rect 16104 -5791 16120 -5757
rect 16162 -5755 16178 -5721
rect 16212 -5755 16306 -5721
rect 16340 -5755 16434 -5721
rect 16468 -5755 16562 -5721
rect 16596 -5755 16612 -5721
rect 16162 -5771 16612 -5755
rect 15666 -5813 16120 -5791
rect 15666 -5839 16612 -5813
rect -2918 -5975 -2340 -5949
rect -1538 -5975 -960 -5949
rect -802 -5975 -224 -5949
rect 26 -5975 236 -5949
rect 505 -5975 535 -5949
rect 600 -5975 700 -5949
rect 860 -5975 960 -5949
rect 1032 -5975 1062 -5949
rect 1314 -5975 1524 -5949
rect 1774 -5975 2352 -5949
rect 2602 -5975 2812 -5949
rect 3081 -5975 3111 -5949
rect 3176 -5975 3276 -5949
rect 3436 -5975 3536 -5949
rect 3608 -5975 3638 -5949
rect 3890 -5975 4100 -5949
rect 4350 -5975 4928 -5949
rect 5178 -5975 5388 -5949
rect 5657 -5975 5687 -5949
rect 5752 -5975 5852 -5949
rect 6012 -5975 6112 -5949
rect 6184 -5975 6214 -5949
rect 6466 -5975 6676 -5949
rect 6926 -5975 7504 -5949
rect 7754 -5975 7964 -5949
rect 8233 -5975 8263 -5949
rect 8328 -5975 8428 -5949
rect 8588 -5975 8688 -5949
rect 8760 -5975 8790 -5949
rect 9042 -5975 9252 -5949
rect 9502 -5975 10080 -5949
rect 10422 -5975 10632 -5949
rect 10809 -5975 10839 -5949
rect 10904 -5975 11004 -5949
rect 11164 -5975 11264 -5949
rect 11336 -5975 11366 -5949
rect 11710 -5975 11920 -5949
rect 13735 -5975 13765 -5949
rect 13821 -5975 13851 -5949
rect 13907 -5975 13937 -5949
rect 13993 -5975 14023 -5949
rect 14079 -5975 14109 -5949
rect 14165 -5975 14195 -5949
rect 14251 -5975 14281 -5949
rect 14337 -5975 14367 -5949
rect 14423 -5975 14453 -5949
rect 14509 -5975 14539 -5949
rect 14595 -5975 14625 -5949
rect 14681 -5975 14711 -5949
rect 14766 -5975 14796 -5949
rect 14852 -5975 14882 -5949
rect 14938 -5975 14968 -5949
rect 15024 -5975 15054 -5949
rect 15110 -5975 15140 -5949
rect 15196 -5975 15226 -5949
rect 15282 -5975 15312 -5949
rect 15368 -5975 15398 -5949
rect 15666 -5975 16612 -5949
rect -2918 -6043 -2340 -6017
rect -1354 -6043 -1144 -6017
rect -890 -6043 -860 -6017
rect -806 -6043 -776 -6017
rect -526 -6043 -316 -6017
rect 29 -6043 59 -6017
rect 115 -6043 145 -6017
rect 201 -6043 231 -6017
rect 287 -6043 317 -6017
rect 670 -6043 880 -6017
rect 1213 -6043 1243 -6017
rect 1498 -6043 1708 -6017
rect 1958 -6043 2168 -6017
rect 2420 -6043 2450 -6017
rect 2522 -6043 2622 -6017
rect 2782 -6043 2882 -6017
rect 2947 -6043 2977 -6017
rect 3246 -6043 3456 -6017
rect 4442 -6043 5388 -6017
rect 6466 -6043 6676 -6017
rect 6928 -6043 6958 -6017
rect 7030 -6043 7130 -6017
rect 7290 -6043 7390 -6017
rect 7455 -6043 7485 -6017
rect 7754 -6043 7964 -6017
rect 8216 -6043 8246 -6017
rect 8318 -6043 8418 -6017
rect 8578 -6043 8678 -6017
rect 8743 -6043 8773 -6017
rect 9042 -6043 9252 -6017
rect 9504 -6043 9534 -6017
rect 9606 -6043 9706 -6017
rect 9866 -6043 9966 -6017
rect 10031 -6043 10061 -6017
rect 10330 -6043 10540 -6017
rect 10790 -6043 10820 -6017
rect 10874 -6043 10904 -6017
rect 10958 -6043 10988 -6017
rect 11042 -6043 11072 -6017
rect 11126 -6043 11156 -6017
rect 11210 -6043 11240 -6017
rect 11294 -6043 11324 -6017
rect 11378 -6043 11408 -6017
rect 11710 -6043 11920 -6017
rect 13642 -6043 14588 -6017
rect 14838 -6043 15784 -6017
rect 16034 -6043 16612 -6017
rect -2918 -6179 -2340 -6153
rect -1354 -6179 -1144 -6153
rect -2918 -6201 -2646 -6179
rect -2918 -6235 -2902 -6201
rect -2868 -6235 -2799 -6201
rect -2765 -6235 -2696 -6201
rect -2662 -6235 -2646 -6201
rect -1228 -6185 -1144 -6179
rect -1228 -6201 -1086 -6185
rect -890 -6195 -860 -6173
rect -2918 -6251 -2646 -6235
rect -2604 -6237 -2340 -6221
rect -2604 -6271 -2588 -6237
rect -2554 -6271 -2489 -6237
rect -2455 -6271 -2390 -6237
rect -2356 -6271 -2340 -6237
rect -2604 -6293 -2340 -6271
rect -1412 -6237 -1270 -6221
rect -1412 -6271 -1396 -6237
rect -1362 -6271 -1270 -6237
rect -1228 -6235 -1136 -6201
rect -1102 -6235 -1086 -6201
rect -1228 -6251 -1086 -6235
rect -952 -6211 -860 -6195
rect -952 -6245 -937 -6211
rect -903 -6245 -860 -6211
rect -952 -6261 -860 -6245
rect -1412 -6287 -1270 -6271
rect -2918 -6319 -2340 -6293
rect -1354 -6293 -1270 -6287
rect -890 -6293 -860 -6261
rect -806 -6195 -776 -6173
rect -526 -6179 -316 -6153
rect -400 -6185 -316 -6179
rect -806 -6211 -718 -6195
rect -806 -6245 -769 -6211
rect -735 -6245 -718 -6211
rect -400 -6201 -258 -6185
rect 29 -6201 59 -6127
rect 115 -6201 145 -6127
rect 201 -6201 231 -6127
rect 287 -6201 317 -6127
rect 670 -6179 880 -6153
rect 796 -6185 880 -6179
rect 796 -6201 938 -6185
rect 1213 -6191 1243 -6127
rect 1498 -6179 1708 -6153
rect 1958 -6179 2168 -6153
rect 1129 -6195 1243 -6191
rect -806 -6261 -718 -6245
rect -584 -6237 -442 -6221
rect -806 -6293 -776 -6261
rect -584 -6271 -568 -6237
rect -534 -6271 -442 -6237
rect -400 -6235 -308 -6201
rect -274 -6235 -258 -6201
rect -400 -6251 -258 -6235
rect -57 -6211 403 -6201
rect -57 -6245 -30 -6211
rect 4 -6245 38 -6211
rect 72 -6245 106 -6211
rect 140 -6245 174 -6211
rect 208 -6245 242 -6211
rect 276 -6245 310 -6211
rect 344 -6245 403 -6211
rect -584 -6287 -442 -6271
rect -526 -6293 -442 -6287
rect -57 -6255 403 -6245
rect -57 -6293 -27 -6255
rect 29 -6293 59 -6255
rect 115 -6293 145 -6255
rect 201 -6293 231 -6255
rect 287 -6293 317 -6255
rect 373 -6293 403 -6255
rect 612 -6237 754 -6221
rect 612 -6271 628 -6237
rect 662 -6271 754 -6237
rect 796 -6235 888 -6201
rect 922 -6235 938 -6201
rect 796 -6251 938 -6235
rect 1072 -6211 1243 -6195
rect 1072 -6245 1082 -6211
rect 1116 -6235 1243 -6211
rect 1624 -6185 1708 -6179
rect 2084 -6185 2168 -6179
rect 1624 -6201 1766 -6185
rect 1116 -6245 1244 -6235
rect 1072 -6261 1244 -6245
rect 612 -6287 754 -6271
rect 670 -6293 754 -6287
rect 1130 -6265 1244 -6261
rect -1354 -6319 -1144 -6293
rect -526 -6319 -316 -6293
rect 670 -6319 880 -6293
rect 1130 -6325 1160 -6265
rect 1214 -6325 1244 -6265
rect 1440 -6237 1582 -6221
rect 1440 -6271 1456 -6237
rect 1490 -6271 1582 -6237
rect 1624 -6235 1716 -6201
rect 1750 -6235 1766 -6201
rect 2084 -6201 2226 -6185
rect 2420 -6199 2450 -6127
rect 1624 -6251 1766 -6235
rect 1900 -6237 2042 -6221
rect 1440 -6287 1582 -6271
rect 1900 -6271 1916 -6237
rect 1950 -6271 2042 -6237
rect 2084 -6235 2176 -6201
rect 2210 -6235 2226 -6201
rect 2084 -6251 2226 -6235
rect 2380 -6211 2450 -6199
rect 2522 -6201 2622 -6173
rect 2782 -6201 2882 -6173
rect 2947 -6195 2977 -6127
rect 3246 -6179 3456 -6153
rect 4442 -6179 5388 -6153
rect 6466 -6179 6676 -6153
rect 3372 -6185 3456 -6179
rect 2380 -6245 2396 -6211
rect 2430 -6245 2450 -6211
rect 2380 -6258 2450 -6245
rect 2500 -6211 2622 -6201
rect 2500 -6245 2516 -6211
rect 2550 -6245 2622 -6211
rect 2500 -6255 2622 -6245
rect 2721 -6211 2882 -6201
rect 2721 -6245 2737 -6211
rect 2771 -6245 2882 -6211
rect 2721 -6255 2882 -6245
rect 1900 -6287 2042 -6271
rect 1498 -6293 1582 -6287
rect 1958 -6293 2042 -6287
rect 2420 -6293 2450 -6258
rect 1498 -6319 1708 -6293
rect 1958 -6319 2168 -6293
rect 2522 -6329 2622 -6255
rect 2782 -6329 2882 -6255
rect 2927 -6211 2981 -6195
rect 2927 -6245 2937 -6211
rect 2971 -6245 2981 -6211
rect 3372 -6201 3514 -6185
rect 2927 -6261 2981 -6245
rect 3188 -6237 3330 -6221
rect 2947 -6293 2977 -6261
rect 3188 -6271 3204 -6237
rect 3238 -6271 3330 -6237
rect 3372 -6235 3464 -6201
rect 3498 -6235 3514 -6201
rect 4934 -6201 5388 -6179
rect 3372 -6251 3514 -6235
rect 4442 -6237 4892 -6221
rect 3188 -6287 3330 -6271
rect 3246 -6293 3330 -6287
rect 4442 -6271 4458 -6237
rect 4492 -6271 4586 -6237
rect 4620 -6271 4714 -6237
rect 4748 -6271 4842 -6237
rect 4876 -6271 4892 -6237
rect 4934 -6235 4950 -6201
rect 4984 -6235 5078 -6201
rect 5112 -6235 5206 -6201
rect 5240 -6235 5334 -6201
rect 5368 -6235 5388 -6201
rect 6592 -6185 6676 -6179
rect 6592 -6201 6734 -6185
rect 6928 -6199 6958 -6127
rect 4934 -6251 5388 -6235
rect 6408 -6237 6550 -6221
rect 4442 -6293 4892 -6271
rect 6408 -6271 6424 -6237
rect 6458 -6271 6550 -6237
rect 6592 -6235 6684 -6201
rect 6718 -6235 6734 -6201
rect 6592 -6251 6734 -6235
rect 6888 -6211 6958 -6199
rect 7030 -6201 7130 -6173
rect 7290 -6201 7390 -6173
rect 7455 -6195 7485 -6127
rect 7754 -6179 7964 -6153
rect 7880 -6185 7964 -6179
rect 6888 -6245 6904 -6211
rect 6938 -6245 6958 -6211
rect 6888 -6258 6958 -6245
rect 7008 -6211 7130 -6201
rect 7008 -6245 7024 -6211
rect 7058 -6245 7130 -6211
rect 7008 -6255 7130 -6245
rect 7229 -6211 7390 -6201
rect 7229 -6245 7245 -6211
rect 7279 -6245 7390 -6211
rect 7229 -6255 7390 -6245
rect 6408 -6287 6550 -6271
rect 6466 -6293 6550 -6287
rect 6928 -6293 6958 -6258
rect 3246 -6319 3456 -6293
rect 4442 -6319 5388 -6293
rect 6466 -6319 6676 -6293
rect 7030 -6329 7130 -6255
rect 7290 -6329 7390 -6255
rect 7435 -6211 7489 -6195
rect 7435 -6245 7445 -6211
rect 7479 -6245 7489 -6211
rect 7880 -6201 8022 -6185
rect 8216 -6199 8246 -6127
rect 7435 -6261 7489 -6245
rect 7696 -6237 7838 -6221
rect 7455 -6293 7485 -6261
rect 7696 -6271 7712 -6237
rect 7746 -6271 7838 -6237
rect 7880 -6235 7972 -6201
rect 8006 -6235 8022 -6201
rect 7880 -6251 8022 -6235
rect 8176 -6211 8246 -6199
rect 8318 -6201 8418 -6173
rect 8578 -6201 8678 -6173
rect 8743 -6195 8773 -6127
rect 9042 -6179 9252 -6153
rect 9168 -6185 9252 -6179
rect 8176 -6245 8192 -6211
rect 8226 -6245 8246 -6211
rect 8176 -6258 8246 -6245
rect 8296 -6211 8418 -6201
rect 8296 -6245 8312 -6211
rect 8346 -6245 8418 -6211
rect 8296 -6255 8418 -6245
rect 8517 -6211 8678 -6201
rect 8517 -6245 8533 -6211
rect 8567 -6245 8678 -6211
rect 8517 -6255 8678 -6245
rect 7696 -6287 7838 -6271
rect 7754 -6293 7838 -6287
rect 8216 -6293 8246 -6258
rect 7754 -6319 7964 -6293
rect 8318 -6329 8418 -6255
rect 8578 -6329 8678 -6255
rect 8723 -6211 8777 -6195
rect 8723 -6245 8733 -6211
rect 8767 -6245 8777 -6211
rect 9168 -6201 9310 -6185
rect 9504 -6199 9534 -6127
rect 8723 -6261 8777 -6245
rect 8984 -6237 9126 -6221
rect 8743 -6293 8773 -6261
rect 8984 -6271 9000 -6237
rect 9034 -6271 9126 -6237
rect 9168 -6235 9260 -6201
rect 9294 -6235 9310 -6201
rect 9168 -6251 9310 -6235
rect 9464 -6211 9534 -6199
rect 9606 -6201 9706 -6173
rect 9866 -6201 9966 -6173
rect 10031 -6195 10061 -6127
rect 10330 -6179 10540 -6153
rect 10456 -6185 10540 -6179
rect 9464 -6245 9480 -6211
rect 9514 -6245 9534 -6211
rect 9464 -6258 9534 -6245
rect 9584 -6211 9706 -6201
rect 9584 -6245 9600 -6211
rect 9634 -6245 9706 -6211
rect 9584 -6255 9706 -6245
rect 9805 -6211 9966 -6201
rect 9805 -6245 9821 -6211
rect 9855 -6245 9966 -6211
rect 9805 -6255 9966 -6245
rect 8984 -6287 9126 -6271
rect 9042 -6293 9126 -6287
rect 9504 -6293 9534 -6258
rect 9042 -6319 9252 -6293
rect 9606 -6329 9706 -6255
rect 9866 -6329 9966 -6255
rect 10011 -6211 10065 -6195
rect 10011 -6245 10021 -6211
rect 10055 -6245 10065 -6211
rect 10456 -6201 10598 -6185
rect 10790 -6195 10820 -6173
rect 10874 -6195 10904 -6173
rect 10958 -6195 10988 -6173
rect 11042 -6195 11072 -6173
rect 10011 -6261 10065 -6245
rect 10272 -6237 10414 -6221
rect 10031 -6293 10061 -6261
rect 10272 -6271 10288 -6237
rect 10322 -6271 10414 -6237
rect 10456 -6235 10548 -6201
rect 10582 -6235 10598 -6201
rect 10456 -6251 10598 -6235
rect 10733 -6211 11072 -6195
rect 10733 -6245 10749 -6211
rect 10783 -6245 10830 -6211
rect 10864 -6245 10914 -6211
rect 10948 -6245 10998 -6211
rect 11032 -6245 11072 -6211
rect 10733 -6261 11072 -6245
rect 10272 -6287 10414 -6271
rect 10330 -6293 10414 -6287
rect 10790 -6293 10820 -6261
rect 10874 -6293 10904 -6261
rect 10958 -6293 10988 -6261
rect 11042 -6293 11072 -6261
rect 11126 -6195 11156 -6173
rect 11210 -6195 11240 -6173
rect 11294 -6195 11324 -6173
rect 11378 -6195 11408 -6173
rect 11710 -6179 11920 -6153
rect 13642 -6179 14588 -6153
rect 14838 -6179 15784 -6153
rect 16034 -6179 16612 -6153
rect 11126 -6211 11408 -6195
rect 11126 -6245 11250 -6211
rect 11284 -6245 11334 -6211
rect 11368 -6245 11408 -6211
rect 11836 -6185 11920 -6179
rect 11836 -6201 11978 -6185
rect 11126 -6261 11408 -6245
rect 11126 -6293 11156 -6261
rect 11210 -6293 11240 -6261
rect 11294 -6293 11324 -6261
rect 11378 -6293 11408 -6261
rect 11652 -6237 11794 -6221
rect 11652 -6271 11668 -6237
rect 11702 -6271 11794 -6237
rect 11836 -6235 11928 -6201
rect 11962 -6235 11978 -6201
rect 14134 -6201 14588 -6179
rect 11836 -6251 11978 -6235
rect 13642 -6237 14092 -6221
rect 11652 -6287 11794 -6271
rect 11710 -6293 11794 -6287
rect 13642 -6271 13658 -6237
rect 13692 -6271 13786 -6237
rect 13820 -6271 13914 -6237
rect 13948 -6271 14042 -6237
rect 14076 -6271 14092 -6237
rect 14134 -6235 14150 -6201
rect 14184 -6235 14278 -6201
rect 14312 -6235 14406 -6201
rect 14440 -6235 14534 -6201
rect 14568 -6235 14588 -6201
rect 15330 -6201 15784 -6179
rect 14134 -6251 14588 -6235
rect 14838 -6237 15288 -6221
rect 13642 -6293 14092 -6271
rect 14838 -6271 14854 -6237
rect 14888 -6271 14982 -6237
rect 15016 -6271 15110 -6237
rect 15144 -6271 15238 -6237
rect 15272 -6271 15288 -6237
rect 15330 -6235 15346 -6201
rect 15380 -6235 15474 -6201
rect 15508 -6235 15602 -6201
rect 15636 -6235 15730 -6201
rect 15764 -6235 15784 -6201
rect 16340 -6201 16612 -6179
rect 15330 -6251 15784 -6235
rect 16034 -6237 16298 -6221
rect 14838 -6293 15288 -6271
rect 16034 -6271 16050 -6237
rect 16084 -6271 16149 -6237
rect 16183 -6271 16248 -6237
rect 16282 -6271 16298 -6237
rect 16340 -6235 16356 -6201
rect 16390 -6235 16459 -6201
rect 16493 -6235 16562 -6201
rect 16596 -6235 16612 -6201
rect 16340 -6251 16612 -6235
rect 16034 -6293 16298 -6271
rect 10330 -6319 10540 -6293
rect 11710 -6319 11920 -6293
rect 13642 -6319 14588 -6293
rect 14838 -6319 15784 -6293
rect 16034 -6319 16612 -6293
rect -2918 -6519 -2340 -6493
rect -1354 -6519 -1144 -6493
rect -890 -6519 -860 -6493
rect -806 -6519 -776 -6493
rect -526 -6519 -316 -6493
rect -57 -6519 -27 -6493
rect 29 -6519 59 -6493
rect 115 -6519 145 -6493
rect 201 -6519 231 -6493
rect 287 -6519 317 -6493
rect 373 -6519 403 -6493
rect 670 -6519 880 -6493
rect 1130 -6519 1160 -6493
rect 1214 -6519 1244 -6493
rect 1498 -6519 1708 -6493
rect 1958 -6519 2168 -6493
rect 2420 -6519 2450 -6493
rect 2522 -6519 2622 -6493
rect 2782 -6519 2882 -6493
rect 2947 -6519 2977 -6493
rect 3246 -6519 3456 -6493
rect 4442 -6519 5388 -6493
rect 6466 -6519 6676 -6493
rect 6928 -6519 6958 -6493
rect 7030 -6519 7130 -6493
rect 7290 -6519 7390 -6493
rect 7455 -6519 7485 -6493
rect 7754 -6519 7964 -6493
rect 8216 -6519 8246 -6493
rect 8318 -6519 8418 -6493
rect 8578 -6519 8678 -6493
rect 8743 -6519 8773 -6493
rect 9042 -6519 9252 -6493
rect 9504 -6519 9534 -6493
rect 9606 -6519 9706 -6493
rect 9866 -6519 9966 -6493
rect 10031 -6519 10061 -6493
rect 10330 -6519 10540 -6493
rect 10790 -6519 10820 -6493
rect 10874 -6519 10904 -6493
rect 10958 -6519 10988 -6493
rect 11042 -6519 11072 -6493
rect 11126 -6519 11156 -6493
rect 11210 -6519 11240 -6493
rect 11294 -6519 11324 -6493
rect 11378 -6519 11408 -6493
rect 11710 -6519 11920 -6493
rect 13642 -6519 14588 -6493
rect 14838 -6519 15784 -6493
rect 16034 -6519 16612 -6493
rect -2918 -6587 -2800 -6561
rect -2550 -6593 -2520 -6567
rect -2466 -6593 -2436 -6567
rect -2278 -6587 -2248 -6561
rect -2193 -6587 -2163 -6561
rect -2098 -6587 -2068 -6561
rect -1995 -6587 -1965 -6561
rect -1863 -6587 -1833 -6561
rect -1768 -6587 -1738 -6561
rect -1684 -6587 -1654 -6561
rect -1570 -6587 -1540 -6561
rect -1359 -6587 -1329 -6561
rect -1275 -6587 -1245 -6561
rect -1087 -6587 -1057 -6561
rect -990 -6587 -960 -6561
rect -802 -6587 -224 -6561
rect 26 -6587 604 -6561
rect 762 -6587 1340 -6561
rect 1590 -6587 2168 -6561
rect 2326 -6587 2904 -6561
rect 3154 -6587 3732 -6561
rect 3890 -6587 4468 -6561
rect 4718 -6587 5296 -6561
rect 5454 -6587 6032 -6561
rect 6282 -6587 6860 -6561
rect 7018 -6587 7596 -6561
rect 7846 -6587 8424 -6561
rect 8582 -6587 9160 -6561
rect 16034 -6587 16612 -6561
rect -2550 -6736 -2520 -6721
rect -2918 -6791 -2800 -6761
rect -2583 -6766 -2520 -6736
rect -2918 -6793 -2880 -6791
rect -2946 -6809 -2880 -6793
rect -2946 -6843 -2930 -6809
rect -2896 -6843 -2880 -6809
rect -2583 -6819 -2553 -6766
rect -2466 -6810 -2436 -6721
rect -2278 -6751 -2248 -6671
rect -2946 -6859 -2880 -6843
rect -2838 -6849 -2772 -6833
rect -2838 -6883 -2822 -6849
rect -2788 -6883 -2772 -6849
rect -2838 -6899 -2772 -6883
rect -2607 -6835 -2553 -6819
rect -2607 -6869 -2597 -6835
rect -2563 -6869 -2553 -6835
rect -2511 -6820 -2436 -6810
rect -2343 -6767 -2248 -6751
rect -2343 -6801 -2333 -6767
rect -2299 -6801 -2248 -6767
rect -2193 -6787 -2163 -6671
rect -2098 -6703 -2068 -6671
rect -2098 -6719 -2037 -6703
rect -2098 -6753 -2081 -6719
rect -2047 -6753 -2037 -6719
rect -2098 -6769 -2037 -6753
rect -2343 -6817 -2248 -6801
rect -2511 -6854 -2495 -6820
rect -2461 -6854 -2436 -6820
rect -2511 -6864 -2436 -6854
rect -2607 -6885 -2553 -6869
rect -2838 -6901 -2800 -6899
rect -2918 -6927 -2800 -6901
rect -2583 -6908 -2553 -6885
rect -2583 -6938 -2520 -6908
rect -2550 -6953 -2520 -6938
rect -2466 -6953 -2436 -6864
rect -2278 -6953 -2248 -6817
rect -2206 -6797 -2140 -6787
rect -2206 -6831 -2190 -6797
rect -2156 -6811 -2140 -6797
rect -2156 -6831 -2037 -6811
rect -2206 -6841 -2037 -6831
rect -2186 -6893 -2120 -6883
rect -2186 -6927 -2170 -6893
rect -2136 -6927 -2120 -6893
rect -2186 -6937 -2120 -6927
rect -2166 -6965 -2136 -6937
rect -2067 -6965 -2037 -6841
rect -1995 -6871 -1965 -6671
rect -1863 -6775 -1833 -6737
rect -1768 -6769 -1738 -6671
rect -1684 -6709 -1654 -6671
rect -1570 -6703 -1540 -6671
rect -1685 -6719 -1619 -6709
rect -1685 -6753 -1669 -6719
rect -1635 -6753 -1619 -6719
rect -1685 -6763 -1619 -6753
rect -1570 -6719 -1489 -6703
rect -1570 -6753 -1533 -6719
rect -1499 -6753 -1489 -6719
rect -1570 -6769 -1489 -6753
rect -1923 -6785 -1833 -6775
rect -1923 -6819 -1907 -6785
rect -1873 -6819 -1833 -6785
rect -1923 -6829 -1833 -6819
rect -1863 -6864 -1833 -6829
rect -1781 -6785 -1727 -6769
rect -1781 -6819 -1771 -6785
rect -1737 -6805 -1727 -6785
rect -1737 -6819 -1612 -6805
rect -1781 -6835 -1612 -6819
rect -1995 -6881 -1921 -6871
rect -1995 -6915 -1971 -6881
rect -1937 -6915 -1921 -6881
rect -1863 -6894 -1819 -6864
rect -1849 -6909 -1819 -6894
rect -1748 -6893 -1684 -6877
rect -1995 -6925 -1921 -6915
rect -1968 -6953 -1938 -6925
rect -1748 -6927 -1728 -6893
rect -1694 -6927 -1684 -6893
rect -1748 -6943 -1684 -6927
rect -1748 -6965 -1718 -6943
rect -1642 -6965 -1612 -6835
rect -1547 -6953 -1517 -6769
rect -1087 -6751 -1057 -6715
rect -1096 -6781 -1057 -6751
rect -1359 -6819 -1329 -6787
rect -1275 -6819 -1245 -6787
rect -1096 -6819 -1066 -6781
rect -802 -6787 -224 -6761
rect 26 -6787 604 -6761
rect 762 -6787 1340 -6761
rect 1590 -6787 2168 -6761
rect 2326 -6787 2904 -6761
rect 3154 -6787 3732 -6761
rect 3890 -6787 4468 -6761
rect 4718 -6787 5296 -6761
rect 5454 -6787 6032 -6761
rect 6282 -6787 6860 -6761
rect 7018 -6787 7596 -6761
rect 7846 -6787 8424 -6761
rect 8582 -6787 9160 -6761
rect 16034 -6787 16612 -6761
rect -990 -6819 -960 -6787
rect -1469 -6835 -1327 -6819
rect -1469 -6869 -1459 -6835
rect -1425 -6869 -1327 -6835
rect -1469 -6885 -1327 -6869
rect -1285 -6835 -1066 -6819
rect -1285 -6869 -1275 -6835
rect -1241 -6869 -1066 -6835
rect -1285 -6885 -1066 -6869
rect -1024 -6835 -960 -6819
rect -488 -6809 -224 -6787
rect -1024 -6869 -1014 -6835
rect -980 -6869 -960 -6835
rect -1024 -6885 -960 -6869
rect -1357 -6907 -1327 -6885
rect -1273 -6907 -1243 -6885
rect -1096 -6914 -1066 -6885
rect -990 -6907 -960 -6885
rect -802 -6845 -530 -6829
rect -802 -6879 -786 -6845
rect -752 -6879 -683 -6845
rect -649 -6879 -580 -6845
rect -546 -6879 -530 -6845
rect -488 -6843 -472 -6809
rect -438 -6843 -373 -6809
rect -339 -6843 -274 -6809
rect -240 -6843 -224 -6809
rect 340 -6809 604 -6787
rect -488 -6859 -224 -6843
rect 26 -6845 298 -6829
rect -802 -6901 -530 -6879
rect 26 -6879 42 -6845
rect 76 -6879 145 -6845
rect 179 -6879 248 -6845
rect 282 -6879 298 -6845
rect 340 -6843 356 -6809
rect 390 -6843 455 -6809
rect 489 -6843 554 -6809
rect 588 -6843 604 -6809
rect 1076 -6809 1340 -6787
rect 340 -6859 604 -6843
rect 762 -6845 1034 -6829
rect 26 -6901 298 -6879
rect 762 -6879 778 -6845
rect 812 -6879 881 -6845
rect 915 -6879 984 -6845
rect 1018 -6879 1034 -6845
rect 1076 -6843 1092 -6809
rect 1126 -6843 1191 -6809
rect 1225 -6843 1290 -6809
rect 1324 -6843 1340 -6809
rect 1904 -6809 2168 -6787
rect 1076 -6859 1340 -6843
rect 1590 -6845 1862 -6829
rect 762 -6901 1034 -6879
rect 1590 -6879 1606 -6845
rect 1640 -6879 1709 -6845
rect 1743 -6879 1812 -6845
rect 1846 -6879 1862 -6845
rect 1904 -6843 1920 -6809
rect 1954 -6843 2019 -6809
rect 2053 -6843 2118 -6809
rect 2152 -6843 2168 -6809
rect 2640 -6809 2904 -6787
rect 1904 -6859 2168 -6843
rect 2326 -6845 2598 -6829
rect 1590 -6901 1862 -6879
rect 2326 -6879 2342 -6845
rect 2376 -6879 2445 -6845
rect 2479 -6879 2548 -6845
rect 2582 -6879 2598 -6845
rect 2640 -6843 2656 -6809
rect 2690 -6843 2755 -6809
rect 2789 -6843 2854 -6809
rect 2888 -6843 2904 -6809
rect 3468 -6809 3732 -6787
rect 2640 -6859 2904 -6843
rect 3154 -6845 3426 -6829
rect 2326 -6901 2598 -6879
rect 3154 -6879 3170 -6845
rect 3204 -6879 3273 -6845
rect 3307 -6879 3376 -6845
rect 3410 -6879 3426 -6845
rect 3468 -6843 3484 -6809
rect 3518 -6843 3583 -6809
rect 3617 -6843 3682 -6809
rect 3716 -6843 3732 -6809
rect 4204 -6809 4468 -6787
rect 3468 -6859 3732 -6843
rect 3890 -6845 4162 -6829
rect 3154 -6901 3426 -6879
rect 3890 -6879 3906 -6845
rect 3940 -6879 4009 -6845
rect 4043 -6879 4112 -6845
rect 4146 -6879 4162 -6845
rect 4204 -6843 4220 -6809
rect 4254 -6843 4319 -6809
rect 4353 -6843 4418 -6809
rect 4452 -6843 4468 -6809
rect 5032 -6809 5296 -6787
rect 4204 -6859 4468 -6843
rect 4718 -6845 4990 -6829
rect 3890 -6901 4162 -6879
rect 4718 -6879 4734 -6845
rect 4768 -6879 4837 -6845
rect 4871 -6879 4940 -6845
rect 4974 -6879 4990 -6845
rect 5032 -6843 5048 -6809
rect 5082 -6843 5147 -6809
rect 5181 -6843 5246 -6809
rect 5280 -6843 5296 -6809
rect 5768 -6809 6032 -6787
rect 5032 -6859 5296 -6843
rect 5454 -6845 5726 -6829
rect 4718 -6901 4990 -6879
rect 5454 -6879 5470 -6845
rect 5504 -6879 5573 -6845
rect 5607 -6879 5676 -6845
rect 5710 -6879 5726 -6845
rect 5768 -6843 5784 -6809
rect 5818 -6843 5883 -6809
rect 5917 -6843 5982 -6809
rect 6016 -6843 6032 -6809
rect 6596 -6809 6860 -6787
rect 5768 -6859 6032 -6843
rect 6282 -6845 6554 -6829
rect 5454 -6901 5726 -6879
rect 6282 -6879 6298 -6845
rect 6332 -6879 6401 -6845
rect 6435 -6879 6504 -6845
rect 6538 -6879 6554 -6845
rect 6596 -6843 6612 -6809
rect 6646 -6843 6711 -6809
rect 6745 -6843 6810 -6809
rect 6844 -6843 6860 -6809
rect 7332 -6809 7596 -6787
rect 6596 -6859 6860 -6843
rect 7018 -6845 7290 -6829
rect 6282 -6901 6554 -6879
rect 7018 -6879 7034 -6845
rect 7068 -6879 7137 -6845
rect 7171 -6879 7240 -6845
rect 7274 -6879 7290 -6845
rect 7332 -6843 7348 -6809
rect 7382 -6843 7447 -6809
rect 7481 -6843 7546 -6809
rect 7580 -6843 7596 -6809
rect 8160 -6809 8424 -6787
rect 7332 -6859 7596 -6843
rect 7846 -6845 8118 -6829
rect 7018 -6901 7290 -6879
rect 7846 -6879 7862 -6845
rect 7896 -6879 7965 -6845
rect 7999 -6879 8068 -6845
rect 8102 -6879 8118 -6845
rect 8160 -6843 8176 -6809
rect 8210 -6843 8275 -6809
rect 8309 -6843 8374 -6809
rect 8408 -6843 8424 -6809
rect 8896 -6809 9160 -6787
rect 8160 -6859 8424 -6843
rect 8582 -6845 8854 -6829
rect 7846 -6901 8118 -6879
rect 8582 -6879 8598 -6845
rect 8632 -6879 8701 -6845
rect 8735 -6879 8804 -6845
rect 8838 -6879 8854 -6845
rect 8896 -6843 8912 -6809
rect 8946 -6843 9011 -6809
rect 9045 -6843 9110 -6809
rect 9144 -6843 9160 -6809
rect 16348 -6809 16612 -6787
rect 8896 -6859 9160 -6843
rect 16034 -6845 16306 -6829
rect 8582 -6901 8854 -6879
rect 16034 -6879 16050 -6845
rect 16084 -6879 16153 -6845
rect 16187 -6879 16256 -6845
rect 16290 -6879 16306 -6845
rect 16348 -6843 16364 -6809
rect 16398 -6843 16463 -6809
rect 16497 -6843 16562 -6809
rect 16596 -6843 16612 -6809
rect 16348 -6859 16612 -6843
rect 16034 -6901 16306 -6879
rect -1096 -6938 -1055 -6914
rect -1085 -6953 -1055 -6938
rect -802 -6927 -224 -6901
rect 26 -6927 604 -6901
rect 762 -6927 1340 -6901
rect 1590 -6927 2168 -6901
rect 2326 -6927 2904 -6901
rect 3154 -6927 3732 -6901
rect 3890 -6927 4468 -6901
rect 4718 -6927 5296 -6901
rect 5454 -6927 6032 -6901
rect 6282 -6927 6860 -6901
rect 7018 -6927 7596 -6901
rect 7846 -6927 8424 -6901
rect 8582 -6927 9160 -6901
rect 16034 -6927 16612 -6901
rect -2918 -7063 -2800 -7037
rect -2550 -7063 -2520 -7037
rect -2466 -7063 -2436 -7037
rect -2278 -7063 -2248 -7037
rect -2166 -7063 -2136 -7037
rect -2067 -7063 -2037 -7037
rect -1968 -7063 -1938 -7037
rect -1849 -7063 -1819 -7037
rect -1748 -7063 -1718 -7037
rect -1642 -7063 -1612 -7037
rect -1547 -7063 -1517 -7037
rect -1357 -7063 -1327 -7037
rect -1273 -7063 -1243 -7037
rect -1085 -7063 -1055 -7037
rect -990 -7063 -960 -7037
rect -802 -7063 -224 -7037
rect 26 -7063 604 -7037
rect 762 -7063 1340 -7037
rect 1590 -7063 2168 -7037
rect 2326 -7063 2904 -7037
rect 3154 -7063 3732 -7037
rect 3890 -7063 4468 -7037
rect 4718 -7063 5296 -7037
rect 5454 -7063 6032 -7037
rect 6282 -7063 6860 -7037
rect 7018 -7063 7596 -7037
rect 7846 -7063 8424 -7037
rect 8582 -7063 9160 -7037
rect 16034 -7063 16612 -7037
rect -2918 -7131 -2340 -7105
rect -1538 -7131 -960 -7105
rect -802 -7131 -224 -7105
rect 26 -7131 604 -7105
rect 762 -7131 1340 -7105
rect 1590 -7131 2168 -7105
rect 2326 -7131 2536 -7105
rect 2975 -7131 3005 -7105
rect 3338 -7131 3548 -7105
rect 3802 -7131 3832 -7105
rect 3886 -7131 3916 -7105
rect 4166 -7131 4376 -7105
rect 4626 -7131 4656 -7105
rect 4735 -7131 4765 -7105
rect 4831 -7131 4861 -7105
rect 4956 -7131 4986 -7105
rect 5052 -7131 5082 -7105
rect 5220 -7131 5250 -7105
rect 5546 -7131 5756 -7105
rect 6006 -7131 6036 -7105
rect 6101 -7131 6131 -7105
rect 6289 -7131 6319 -7105
rect 6373 -7131 6403 -7105
rect 6563 -7131 6593 -7105
rect 6658 -7131 6688 -7105
rect 6764 -7131 6794 -7105
rect 6865 -7131 6895 -7105
rect 6984 -7131 7014 -7105
rect 7083 -7131 7113 -7105
rect 7182 -7131 7212 -7105
rect 7294 -7131 7324 -7105
rect 7482 -7131 7512 -7105
rect 7566 -7131 7596 -7105
rect 7846 -7131 8424 -7105
rect 8582 -7131 9160 -7105
rect 16034 -7131 16612 -7105
rect -2918 -7267 -2340 -7241
rect -1538 -7267 -960 -7241
rect -802 -7267 -224 -7241
rect 26 -7267 604 -7241
rect 762 -7267 1340 -7241
rect 1590 -7267 2168 -7241
rect -2918 -7289 -2646 -7267
rect -2918 -7323 -2902 -7289
rect -2868 -7323 -2799 -7289
rect -2765 -7323 -2696 -7289
rect -2662 -7323 -2646 -7289
rect -1232 -7289 -960 -7267
rect -2918 -7339 -2646 -7323
rect -2604 -7325 -2340 -7309
rect -2604 -7359 -2588 -7325
rect -2554 -7359 -2489 -7325
rect -2455 -7359 -2390 -7325
rect -2356 -7359 -2340 -7325
rect -2604 -7381 -2340 -7359
rect -2918 -7407 -2340 -7381
rect -1538 -7325 -1274 -7309
rect -1538 -7359 -1522 -7325
rect -1488 -7359 -1423 -7325
rect -1389 -7359 -1324 -7325
rect -1290 -7359 -1274 -7325
rect -1232 -7323 -1216 -7289
rect -1182 -7323 -1113 -7289
rect -1079 -7323 -1010 -7289
rect -976 -7323 -960 -7289
rect -496 -7289 -224 -7267
rect -1232 -7339 -960 -7323
rect -802 -7325 -538 -7309
rect -1538 -7381 -1274 -7359
rect -802 -7359 -786 -7325
rect -752 -7359 -687 -7325
rect -653 -7359 -588 -7325
rect -554 -7359 -538 -7325
rect -496 -7323 -480 -7289
rect -446 -7323 -377 -7289
rect -343 -7323 -274 -7289
rect -240 -7323 -224 -7289
rect 332 -7289 604 -7267
rect -496 -7339 -224 -7323
rect 26 -7325 290 -7309
rect -802 -7381 -538 -7359
rect 26 -7359 42 -7325
rect 76 -7359 141 -7325
rect 175 -7359 240 -7325
rect 274 -7359 290 -7325
rect 332 -7323 348 -7289
rect 382 -7323 451 -7289
rect 485 -7323 554 -7289
rect 588 -7323 604 -7289
rect 1068 -7289 1340 -7267
rect 332 -7339 604 -7323
rect 762 -7325 1026 -7309
rect 26 -7381 290 -7359
rect 762 -7359 778 -7325
rect 812 -7359 877 -7325
rect 911 -7359 976 -7325
rect 1010 -7359 1026 -7325
rect 1068 -7323 1084 -7289
rect 1118 -7323 1187 -7289
rect 1221 -7323 1290 -7289
rect 1324 -7323 1340 -7289
rect 1896 -7289 2168 -7267
rect 2326 -7267 2536 -7241
rect 2326 -7273 2410 -7267
rect 1068 -7339 1340 -7323
rect 1590 -7325 1854 -7309
rect 762 -7381 1026 -7359
rect 1590 -7359 1606 -7325
rect 1640 -7359 1705 -7325
rect 1739 -7359 1804 -7325
rect 1838 -7359 1854 -7325
rect 1896 -7323 1912 -7289
rect 1946 -7323 2015 -7289
rect 2049 -7323 2118 -7289
rect 2152 -7323 2168 -7289
rect 1896 -7339 2168 -7323
rect 2268 -7289 2410 -7273
rect 2268 -7323 2284 -7289
rect 2318 -7323 2410 -7289
rect 2975 -7279 3005 -7215
rect 3338 -7267 3548 -7241
rect 3338 -7273 3422 -7267
rect 2975 -7283 3089 -7279
rect 2975 -7299 3146 -7283
rect 2268 -7339 2410 -7323
rect 2452 -7325 2594 -7309
rect 2975 -7323 3102 -7299
rect 1590 -7381 1854 -7359
rect 2452 -7359 2544 -7325
rect 2578 -7359 2594 -7325
rect 2452 -7375 2594 -7359
rect 2974 -7333 3102 -7323
rect 3136 -7333 3146 -7299
rect 2974 -7349 3146 -7333
rect 3280 -7289 3422 -7273
rect 3802 -7283 3832 -7261
rect 3280 -7323 3296 -7289
rect 3330 -7323 3422 -7289
rect 3740 -7299 3832 -7283
rect 3280 -7339 3422 -7323
rect 3464 -7325 3606 -7309
rect 2974 -7353 3088 -7349
rect 2452 -7381 2536 -7375
rect -1538 -7407 -960 -7381
rect -802 -7407 -224 -7381
rect 26 -7407 604 -7381
rect 762 -7407 1340 -7381
rect 1590 -7407 2168 -7381
rect 2326 -7407 2536 -7381
rect 2974 -7413 3004 -7353
rect 3058 -7413 3088 -7353
rect 3464 -7359 3556 -7325
rect 3590 -7359 3606 -7325
rect 3740 -7333 3755 -7299
rect 3789 -7333 3832 -7299
rect 3740 -7349 3832 -7333
rect 3464 -7375 3606 -7359
rect 3464 -7381 3548 -7375
rect 3802 -7381 3832 -7349
rect 3886 -7283 3916 -7261
rect 4166 -7267 4376 -7241
rect 4166 -7273 4250 -7267
rect 3886 -7299 3974 -7283
rect 3886 -7333 3923 -7299
rect 3957 -7333 3974 -7299
rect 3886 -7349 3974 -7333
rect 4108 -7289 4250 -7273
rect 4626 -7283 4656 -7261
rect 4735 -7283 4765 -7215
rect 4831 -7247 4861 -7215
rect 4956 -7247 4986 -7215
rect 4831 -7263 4914 -7247
rect 4108 -7323 4124 -7289
rect 4158 -7323 4250 -7289
rect 4623 -7299 4677 -7283
rect 4108 -7339 4250 -7323
rect 4292 -7325 4434 -7309
rect 3886 -7381 3916 -7349
rect 4292 -7359 4384 -7325
rect 4418 -7359 4434 -7325
rect 4623 -7333 4633 -7299
rect 4667 -7333 4677 -7299
rect 4623 -7349 4677 -7333
rect 4719 -7299 4773 -7283
rect 4719 -7333 4729 -7299
rect 4763 -7333 4773 -7299
rect 4831 -7297 4870 -7263
rect 4904 -7297 4914 -7263
rect 4831 -7313 4914 -7297
rect 4956 -7263 5010 -7247
rect 4956 -7297 4966 -7263
rect 5000 -7297 5010 -7263
rect 5052 -7253 5082 -7215
rect 5052 -7263 5178 -7253
rect 5052 -7283 5128 -7263
rect 4956 -7313 5010 -7297
rect 5112 -7297 5128 -7283
rect 5162 -7297 5178 -7263
rect 5112 -7307 5178 -7297
rect 4719 -7349 4773 -7333
rect 4292 -7375 4434 -7359
rect 4292 -7381 4376 -7375
rect 4626 -7381 4656 -7349
rect 3338 -7407 3548 -7381
rect 4166 -7407 4376 -7381
rect 4735 -7458 4765 -7349
rect 4956 -7413 4986 -7313
rect 4838 -7443 4986 -7413
rect 5028 -7376 5082 -7360
rect 5028 -7410 5038 -7376
rect 5072 -7410 5082 -7376
rect 5028 -7426 5082 -7410
rect 4838 -7458 4868 -7443
rect 5052 -7458 5082 -7426
rect 5124 -7458 5154 -7307
rect 5220 -7360 5250 -7215
rect 5546 -7267 5756 -7241
rect 6101 -7230 6131 -7215
rect 6101 -7254 6142 -7230
rect 5546 -7273 5630 -7267
rect 5488 -7289 5630 -7273
rect 5488 -7323 5504 -7289
rect 5538 -7323 5630 -7289
rect 6006 -7283 6036 -7261
rect 6112 -7283 6142 -7254
rect 6289 -7283 6319 -7261
rect 6373 -7283 6403 -7261
rect 6006 -7299 6070 -7283
rect 5488 -7339 5630 -7323
rect 5672 -7325 5814 -7309
rect 5196 -7376 5250 -7360
rect 5196 -7410 5206 -7376
rect 5240 -7410 5250 -7376
rect 5672 -7359 5764 -7325
rect 5798 -7359 5814 -7325
rect 5672 -7375 5814 -7359
rect 6006 -7333 6026 -7299
rect 6060 -7333 6070 -7299
rect 6006 -7349 6070 -7333
rect 6112 -7299 6331 -7283
rect 6112 -7333 6287 -7299
rect 6321 -7333 6331 -7299
rect 6112 -7349 6331 -7333
rect 6373 -7299 6515 -7283
rect 6373 -7333 6471 -7299
rect 6505 -7333 6515 -7299
rect 6373 -7349 6515 -7333
rect 5672 -7381 5756 -7375
rect 6006 -7381 6036 -7349
rect 5196 -7426 5250 -7410
rect 5220 -7458 5250 -7426
rect 5546 -7407 5756 -7381
rect 4735 -7568 4765 -7542
rect 4838 -7568 4868 -7542
rect 5052 -7568 5082 -7542
rect 5124 -7568 5154 -7542
rect 5220 -7568 5250 -7542
rect 6112 -7387 6142 -7349
rect 6291 -7381 6321 -7349
rect 6375 -7381 6405 -7349
rect 6103 -7417 6142 -7387
rect 6103 -7453 6133 -7417
rect 6563 -7399 6593 -7215
rect 6658 -7333 6688 -7203
rect 6764 -7225 6794 -7203
rect 6730 -7241 6794 -7225
rect 6730 -7275 6740 -7241
rect 6774 -7275 6794 -7241
rect 6984 -7243 7014 -7215
rect 6967 -7253 7041 -7243
rect 6730 -7291 6794 -7275
rect 6865 -7274 6895 -7259
rect 6865 -7304 6909 -7274
rect 6967 -7287 6983 -7253
rect 7017 -7287 7041 -7253
rect 6967 -7297 7041 -7287
rect 6658 -7349 6827 -7333
rect 6658 -7363 6783 -7349
rect 6773 -7383 6783 -7363
rect 6817 -7383 6827 -7349
rect 6773 -7399 6827 -7383
rect 6879 -7339 6909 -7304
rect 6879 -7349 6969 -7339
rect 6879 -7383 6919 -7349
rect 6953 -7383 6969 -7349
rect 6879 -7393 6969 -7383
rect 6535 -7415 6616 -7399
rect 6535 -7449 6545 -7415
rect 6579 -7449 6616 -7415
rect 6535 -7465 6616 -7449
rect 6665 -7415 6731 -7405
rect 6665 -7449 6681 -7415
rect 6715 -7449 6731 -7415
rect 6665 -7459 6731 -7449
rect 6586 -7497 6616 -7465
rect 6700 -7497 6730 -7459
rect 6784 -7497 6814 -7399
rect 6879 -7431 6909 -7393
rect 7011 -7497 7041 -7297
rect 7083 -7327 7113 -7203
rect 7182 -7231 7212 -7203
rect 7166 -7241 7232 -7231
rect 7166 -7275 7182 -7241
rect 7216 -7275 7232 -7241
rect 7166 -7285 7232 -7275
rect 7083 -7337 7252 -7327
rect 7083 -7357 7202 -7337
rect 7186 -7371 7202 -7357
rect 7236 -7371 7252 -7337
rect 7186 -7381 7252 -7371
rect 7294 -7351 7324 -7215
rect 7482 -7304 7512 -7215
rect 7566 -7230 7596 -7215
rect 7566 -7260 7629 -7230
rect 7599 -7283 7629 -7260
rect 7846 -7267 8424 -7241
rect 8582 -7267 9160 -7241
rect 16034 -7267 16612 -7241
rect 7599 -7299 7653 -7283
rect 7482 -7314 7557 -7304
rect 7482 -7348 7507 -7314
rect 7541 -7348 7557 -7314
rect 7294 -7367 7389 -7351
rect 7083 -7415 7144 -7399
rect 7083 -7449 7093 -7415
rect 7127 -7449 7144 -7415
rect 7083 -7465 7144 -7449
rect 7114 -7497 7144 -7465
rect 7209 -7497 7239 -7381
rect 7294 -7401 7345 -7367
rect 7379 -7401 7389 -7367
rect 7294 -7417 7389 -7401
rect 7482 -7358 7557 -7348
rect 7599 -7333 7609 -7299
rect 7643 -7333 7653 -7299
rect 8152 -7289 8424 -7267
rect 7599 -7349 7653 -7333
rect 7846 -7325 8110 -7309
rect 7294 -7497 7324 -7417
rect 7482 -7447 7512 -7358
rect 7599 -7402 7629 -7349
rect 7846 -7359 7862 -7325
rect 7896 -7359 7961 -7325
rect 7995 -7359 8060 -7325
rect 8094 -7359 8110 -7325
rect 8152 -7323 8168 -7289
rect 8202 -7323 8271 -7289
rect 8305 -7323 8374 -7289
rect 8408 -7323 8424 -7289
rect 8888 -7289 9160 -7267
rect 8152 -7339 8424 -7323
rect 8582 -7325 8846 -7309
rect 7846 -7381 8110 -7359
rect 8582 -7359 8598 -7325
rect 8632 -7359 8697 -7325
rect 8731 -7359 8796 -7325
rect 8830 -7359 8846 -7325
rect 8888 -7323 8904 -7289
rect 8938 -7323 9007 -7289
rect 9041 -7323 9110 -7289
rect 9144 -7323 9160 -7289
rect 16340 -7289 16612 -7267
rect 8888 -7339 9160 -7323
rect 16034 -7325 16298 -7309
rect 8582 -7381 8846 -7359
rect 16034 -7359 16050 -7325
rect 16084 -7359 16149 -7325
rect 16183 -7359 16248 -7325
rect 16282 -7359 16298 -7325
rect 16340 -7323 16356 -7289
rect 16390 -7323 16459 -7289
rect 16493 -7323 16562 -7289
rect 16596 -7323 16612 -7289
rect 16340 -7339 16612 -7323
rect 16034 -7381 16298 -7359
rect 7566 -7432 7629 -7402
rect 7846 -7407 8424 -7381
rect 8582 -7407 9160 -7381
rect 7566 -7447 7596 -7432
rect -2918 -7607 -2340 -7581
rect -1538 -7607 -960 -7581
rect -802 -7607 -224 -7581
rect 26 -7607 604 -7581
rect 762 -7607 1340 -7581
rect 1590 -7607 2168 -7581
rect 2326 -7607 2536 -7581
rect 2974 -7607 3004 -7581
rect 3058 -7607 3088 -7581
rect 3338 -7607 3548 -7581
rect 3802 -7607 3832 -7581
rect 3886 -7607 3916 -7581
rect 4166 -7607 4376 -7581
rect 4626 -7607 4656 -7581
rect 5546 -7607 5756 -7581
rect 6006 -7607 6036 -7581
rect 6103 -7607 6133 -7581
rect 6291 -7607 6321 -7581
rect 6375 -7607 6405 -7581
rect 6586 -7607 6616 -7581
rect 6700 -7607 6730 -7581
rect 6784 -7607 6814 -7581
rect 6879 -7607 6909 -7581
rect 7011 -7607 7041 -7581
rect 7114 -7607 7144 -7581
rect 7209 -7607 7239 -7581
rect 7294 -7607 7324 -7581
rect 7482 -7601 7512 -7575
rect 7566 -7601 7596 -7575
rect 16034 -7407 16612 -7381
rect 7846 -7607 8424 -7581
rect 8582 -7607 9160 -7581
rect 16034 -7607 16612 -7581
rect -2918 -7675 -2340 -7649
rect -1354 -7675 -1144 -7649
rect -890 -7675 -860 -7649
rect -806 -7675 -776 -7649
rect -526 -7675 -316 -7649
rect -57 -7675 -27 -7649
rect 29 -7675 59 -7649
rect 115 -7675 145 -7649
rect 201 -7675 231 -7649
rect 287 -7675 317 -7649
rect 373 -7675 403 -7649
rect 670 -7675 880 -7649
rect 1130 -7675 1160 -7649
rect 1214 -7675 1244 -7649
rect 1498 -7675 1708 -7649
rect 1958 -7675 2168 -7649
rect 2420 -7675 2450 -7649
rect 2522 -7675 2622 -7649
rect 2782 -7675 2882 -7649
rect 2947 -7675 2977 -7649
rect 3246 -7675 3456 -7649
rect 4442 -7675 5388 -7649
rect 6466 -7675 6676 -7649
rect 6928 -7675 6958 -7649
rect 7030 -7675 7130 -7649
rect 7290 -7675 7390 -7649
rect 7455 -7675 7485 -7649
rect 7754 -7675 7964 -7649
rect 8216 -7675 8246 -7649
rect 8318 -7675 8418 -7649
rect 8578 -7675 8678 -7649
rect 8743 -7675 8773 -7649
rect 9042 -7675 9252 -7649
rect 9504 -7675 9534 -7649
rect 9606 -7675 9706 -7649
rect 9866 -7675 9966 -7649
rect 10031 -7675 10061 -7649
rect 10330 -7675 10540 -7649
rect 10790 -7675 10820 -7649
rect 10874 -7675 10904 -7649
rect 10958 -7675 10988 -7649
rect 11042 -7675 11072 -7649
rect 11126 -7675 11156 -7649
rect 11210 -7675 11240 -7649
rect 11294 -7675 11324 -7649
rect 11378 -7675 11408 -7649
rect 11710 -7675 11920 -7649
rect 13642 -7675 14588 -7649
rect 14838 -7675 15784 -7649
rect 16034 -7675 16612 -7649
rect -2918 -7875 -2340 -7849
rect -1354 -7875 -1144 -7849
rect -526 -7875 -316 -7849
rect 670 -7875 880 -7849
rect -2918 -7897 -2654 -7875
rect -1354 -7881 -1270 -7875
rect -2918 -7931 -2902 -7897
rect -2868 -7931 -2803 -7897
rect -2769 -7931 -2704 -7897
rect -2670 -7931 -2654 -7897
rect -1412 -7897 -1270 -7881
rect -2918 -7947 -2654 -7931
rect -2612 -7933 -2340 -7917
rect -2612 -7967 -2596 -7933
rect -2562 -7967 -2493 -7933
rect -2459 -7967 -2390 -7933
rect -2356 -7967 -2340 -7933
rect -1412 -7931 -1396 -7897
rect -1362 -7931 -1270 -7897
rect -890 -7907 -860 -7875
rect -1412 -7947 -1270 -7931
rect -1228 -7933 -1086 -7917
rect -2612 -7989 -2340 -7967
rect -1228 -7967 -1136 -7933
rect -1102 -7967 -1086 -7933
rect -1228 -7983 -1086 -7967
rect -952 -7923 -860 -7907
rect -952 -7957 -937 -7923
rect -903 -7957 -860 -7923
rect -952 -7973 -860 -7957
rect -1228 -7989 -1144 -7983
rect -2918 -8015 -2340 -7989
rect -1354 -8015 -1144 -7989
rect -890 -7995 -860 -7973
rect -806 -7907 -776 -7875
rect -526 -7881 -442 -7875
rect -584 -7897 -442 -7881
rect -806 -7923 -718 -7907
rect -806 -7957 -769 -7923
rect -735 -7957 -718 -7923
rect -584 -7931 -568 -7897
rect -534 -7931 -442 -7897
rect -57 -7913 -27 -7875
rect 29 -7913 59 -7875
rect 115 -7913 145 -7875
rect 201 -7913 231 -7875
rect 287 -7913 317 -7875
rect 373 -7913 403 -7875
rect 670 -7881 754 -7875
rect -584 -7947 -442 -7931
rect -400 -7933 -258 -7917
rect -806 -7973 -718 -7957
rect -400 -7967 -308 -7933
rect -274 -7967 -258 -7933
rect -57 -7923 403 -7913
rect -57 -7957 -30 -7923
rect 4 -7957 38 -7923
rect 72 -7957 106 -7923
rect 140 -7957 174 -7923
rect 208 -7957 242 -7923
rect 276 -7957 310 -7923
rect 344 -7957 403 -7923
rect 612 -7897 754 -7881
rect 612 -7931 628 -7897
rect 662 -7931 754 -7897
rect 1130 -7903 1160 -7843
rect 1214 -7903 1244 -7843
rect 1498 -7875 1708 -7849
rect 1958 -7875 2168 -7849
rect 1498 -7881 1582 -7875
rect 1958 -7881 2042 -7875
rect 1130 -7907 1244 -7903
rect 612 -7947 754 -7931
rect 796 -7933 938 -7917
rect -57 -7967 403 -7957
rect 796 -7967 888 -7933
rect 922 -7967 938 -7933
rect -806 -7995 -776 -7973
rect -400 -7983 -258 -7967
rect -400 -7989 -316 -7983
rect -526 -8015 -316 -7989
rect 29 -8041 59 -7967
rect 115 -8041 145 -7967
rect 201 -8041 231 -7967
rect 287 -8041 317 -7967
rect 796 -7983 938 -7967
rect 1072 -7923 1244 -7907
rect 1072 -7957 1082 -7923
rect 1116 -7933 1244 -7923
rect 1440 -7897 1582 -7881
rect 1440 -7931 1456 -7897
rect 1490 -7931 1582 -7897
rect 1900 -7897 2042 -7881
rect 1116 -7957 1243 -7933
rect 1440 -7947 1582 -7931
rect 1624 -7933 1766 -7917
rect 1072 -7973 1243 -7957
rect 1129 -7977 1243 -7973
rect 796 -7989 880 -7983
rect 670 -8015 880 -7989
rect 1213 -8041 1243 -7977
rect 1624 -7967 1716 -7933
rect 1750 -7967 1766 -7933
rect 1900 -7931 1916 -7897
rect 1950 -7931 2042 -7897
rect 2420 -7910 2450 -7875
rect 1900 -7947 2042 -7931
rect 2084 -7933 2226 -7917
rect 1624 -7983 1766 -7967
rect 2084 -7967 2176 -7933
rect 2210 -7967 2226 -7933
rect 2084 -7983 2226 -7967
rect 2380 -7923 2450 -7910
rect 2522 -7913 2622 -7839
rect 2782 -7913 2882 -7839
rect 3246 -7875 3456 -7849
rect 4442 -7875 5388 -7849
rect 6466 -7875 6676 -7849
rect 2947 -7907 2977 -7875
rect 3246 -7881 3330 -7875
rect 3188 -7897 3330 -7881
rect 2380 -7957 2396 -7923
rect 2430 -7957 2450 -7923
rect 2380 -7969 2450 -7957
rect 2500 -7923 2622 -7913
rect 2500 -7957 2516 -7923
rect 2550 -7957 2622 -7923
rect 2500 -7967 2622 -7957
rect 2721 -7923 2882 -7913
rect 2721 -7957 2737 -7923
rect 2771 -7957 2882 -7923
rect 2721 -7967 2882 -7957
rect 1624 -7989 1708 -7983
rect 2084 -7989 2168 -7983
rect 1498 -8015 1708 -7989
rect 1958 -8015 2168 -7989
rect 2420 -8041 2450 -7969
rect 2522 -7995 2622 -7967
rect 2782 -7995 2882 -7967
rect 2927 -7923 2981 -7907
rect 2927 -7957 2937 -7923
rect 2971 -7957 2981 -7923
rect 3188 -7931 3204 -7897
rect 3238 -7931 3330 -7897
rect 4442 -7897 4892 -7875
rect 6466 -7881 6550 -7875
rect 3188 -7947 3330 -7931
rect 3372 -7933 3514 -7917
rect 2927 -7973 2981 -7957
rect 3372 -7967 3464 -7933
rect 3498 -7967 3514 -7933
rect 4442 -7931 4458 -7897
rect 4492 -7931 4586 -7897
rect 4620 -7931 4714 -7897
rect 4748 -7931 4842 -7897
rect 4876 -7931 4892 -7897
rect 6408 -7897 6550 -7881
rect 4442 -7947 4892 -7931
rect 4934 -7933 5388 -7917
rect 2947 -8041 2977 -7973
rect 3372 -7983 3514 -7967
rect 4934 -7967 4950 -7933
rect 4984 -7967 5078 -7933
rect 5112 -7967 5206 -7933
rect 5240 -7967 5334 -7933
rect 5368 -7967 5388 -7933
rect 6408 -7931 6424 -7897
rect 6458 -7931 6550 -7897
rect 6928 -7910 6958 -7875
rect 6408 -7947 6550 -7931
rect 6592 -7933 6734 -7917
rect 3372 -7989 3456 -7983
rect 4934 -7989 5388 -7967
rect 6592 -7967 6684 -7933
rect 6718 -7967 6734 -7933
rect 6592 -7983 6734 -7967
rect 6888 -7923 6958 -7910
rect 7030 -7913 7130 -7839
rect 7290 -7913 7390 -7839
rect 7754 -7875 7964 -7849
rect 7455 -7907 7485 -7875
rect 7754 -7881 7838 -7875
rect 7696 -7897 7838 -7881
rect 6888 -7957 6904 -7923
rect 6938 -7957 6958 -7923
rect 6888 -7969 6958 -7957
rect 7008 -7923 7130 -7913
rect 7008 -7957 7024 -7923
rect 7058 -7957 7130 -7923
rect 7008 -7967 7130 -7957
rect 7229 -7923 7390 -7913
rect 7229 -7957 7245 -7923
rect 7279 -7957 7390 -7923
rect 7229 -7967 7390 -7957
rect 6592 -7989 6676 -7983
rect 3246 -8015 3456 -7989
rect 4442 -8015 5388 -7989
rect 6466 -8015 6676 -7989
rect 6928 -8041 6958 -7969
rect 7030 -7995 7130 -7967
rect 7290 -7995 7390 -7967
rect 7435 -7923 7489 -7907
rect 7435 -7957 7445 -7923
rect 7479 -7957 7489 -7923
rect 7696 -7931 7712 -7897
rect 7746 -7931 7838 -7897
rect 8216 -7910 8246 -7875
rect 7696 -7947 7838 -7931
rect 7880 -7933 8022 -7917
rect 7435 -7973 7489 -7957
rect 7880 -7967 7972 -7933
rect 8006 -7967 8022 -7933
rect 7455 -8041 7485 -7973
rect 7880 -7983 8022 -7967
rect 8176 -7923 8246 -7910
rect 8318 -7913 8418 -7839
rect 8578 -7913 8678 -7839
rect 9042 -7875 9252 -7849
rect 8743 -7907 8773 -7875
rect 9042 -7881 9126 -7875
rect 8984 -7897 9126 -7881
rect 8176 -7957 8192 -7923
rect 8226 -7957 8246 -7923
rect 8176 -7969 8246 -7957
rect 8296 -7923 8418 -7913
rect 8296 -7957 8312 -7923
rect 8346 -7957 8418 -7923
rect 8296 -7967 8418 -7957
rect 8517 -7923 8678 -7913
rect 8517 -7957 8533 -7923
rect 8567 -7957 8678 -7923
rect 8517 -7967 8678 -7957
rect 7880 -7989 7964 -7983
rect 7754 -8015 7964 -7989
rect 8216 -8041 8246 -7969
rect 8318 -7995 8418 -7967
rect 8578 -7995 8678 -7967
rect 8723 -7923 8777 -7907
rect 8723 -7957 8733 -7923
rect 8767 -7957 8777 -7923
rect 8984 -7931 9000 -7897
rect 9034 -7931 9126 -7897
rect 9504 -7910 9534 -7875
rect 8984 -7947 9126 -7931
rect 9168 -7933 9310 -7917
rect 8723 -7973 8777 -7957
rect 9168 -7967 9260 -7933
rect 9294 -7967 9310 -7933
rect 8743 -8041 8773 -7973
rect 9168 -7983 9310 -7967
rect 9464 -7923 9534 -7910
rect 9606 -7913 9706 -7839
rect 9866 -7913 9966 -7839
rect 10330 -7875 10540 -7849
rect 11710 -7875 11920 -7849
rect 13642 -7875 14588 -7849
rect 14838 -7875 15784 -7849
rect 16034 -7875 16612 -7849
rect 10031 -7907 10061 -7875
rect 10330 -7881 10414 -7875
rect 10272 -7897 10414 -7881
rect 9464 -7957 9480 -7923
rect 9514 -7957 9534 -7923
rect 9464 -7969 9534 -7957
rect 9584 -7923 9706 -7913
rect 9584 -7957 9600 -7923
rect 9634 -7957 9706 -7923
rect 9584 -7967 9706 -7957
rect 9805 -7923 9966 -7913
rect 9805 -7957 9821 -7923
rect 9855 -7957 9966 -7923
rect 9805 -7967 9966 -7957
rect 9168 -7989 9252 -7983
rect 9042 -8015 9252 -7989
rect 9504 -8041 9534 -7969
rect 9606 -7995 9706 -7967
rect 9866 -7995 9966 -7967
rect 10011 -7923 10065 -7907
rect 10011 -7957 10021 -7923
rect 10055 -7957 10065 -7923
rect 10272 -7931 10288 -7897
rect 10322 -7931 10414 -7897
rect 10790 -7907 10820 -7875
rect 10874 -7907 10904 -7875
rect 10958 -7907 10988 -7875
rect 11042 -7907 11072 -7875
rect 10272 -7947 10414 -7931
rect 10456 -7933 10598 -7917
rect 10011 -7973 10065 -7957
rect 10456 -7967 10548 -7933
rect 10582 -7967 10598 -7933
rect 10031 -8041 10061 -7973
rect 10456 -7983 10598 -7967
rect 10733 -7923 11072 -7907
rect 10733 -7957 10749 -7923
rect 10783 -7957 10830 -7923
rect 10864 -7957 10914 -7923
rect 10948 -7957 10998 -7923
rect 11032 -7957 11072 -7923
rect 10733 -7973 11072 -7957
rect 10456 -7989 10540 -7983
rect 10330 -8015 10540 -7989
rect 10790 -7995 10820 -7973
rect 10874 -7995 10904 -7973
rect 10958 -7995 10988 -7973
rect 11042 -7995 11072 -7973
rect 11126 -7907 11156 -7875
rect 11210 -7907 11240 -7875
rect 11294 -7907 11324 -7875
rect 11378 -7907 11408 -7875
rect 11710 -7881 11794 -7875
rect 11126 -7923 11408 -7907
rect 11126 -7957 11250 -7923
rect 11284 -7957 11334 -7923
rect 11368 -7957 11408 -7923
rect 11652 -7897 11794 -7881
rect 11652 -7931 11668 -7897
rect 11702 -7931 11794 -7897
rect 13642 -7897 14092 -7875
rect 11652 -7947 11794 -7931
rect 11836 -7933 11978 -7917
rect 11126 -7973 11408 -7957
rect 11126 -7995 11156 -7973
rect 11210 -7995 11240 -7973
rect 11294 -7995 11324 -7973
rect 11378 -7995 11408 -7973
rect 11836 -7967 11928 -7933
rect 11962 -7967 11978 -7933
rect 13642 -7931 13658 -7897
rect 13692 -7931 13786 -7897
rect 13820 -7931 13914 -7897
rect 13948 -7931 14042 -7897
rect 14076 -7931 14092 -7897
rect 14838 -7897 15288 -7875
rect 13642 -7947 14092 -7931
rect 14134 -7933 14588 -7917
rect 11836 -7983 11978 -7967
rect 14134 -7967 14150 -7933
rect 14184 -7967 14278 -7933
rect 14312 -7967 14406 -7933
rect 14440 -7967 14534 -7933
rect 14568 -7967 14588 -7933
rect 14838 -7931 14854 -7897
rect 14888 -7931 14982 -7897
rect 15016 -7931 15110 -7897
rect 15144 -7931 15238 -7897
rect 15272 -7931 15288 -7897
rect 16034 -7897 16298 -7875
rect 14838 -7947 15288 -7931
rect 15330 -7933 15784 -7917
rect 11836 -7989 11920 -7983
rect 14134 -7989 14588 -7967
rect 15330 -7967 15346 -7933
rect 15380 -7967 15474 -7933
rect 15508 -7967 15602 -7933
rect 15636 -7967 15730 -7933
rect 15764 -7967 15784 -7933
rect 16034 -7931 16050 -7897
rect 16084 -7931 16149 -7897
rect 16183 -7931 16248 -7897
rect 16282 -7931 16298 -7897
rect 16034 -7947 16298 -7931
rect 16340 -7933 16612 -7917
rect 15330 -7989 15784 -7967
rect 16340 -7967 16356 -7933
rect 16390 -7967 16459 -7933
rect 16493 -7967 16562 -7933
rect 16596 -7967 16612 -7933
rect 16340 -7989 16612 -7967
rect 11710 -8015 11920 -7989
rect 13642 -8015 14588 -7989
rect 14838 -8015 15784 -7989
rect 16034 -8015 16612 -7989
rect -2918 -8151 -2340 -8125
rect -1354 -8151 -1144 -8125
rect -890 -8151 -860 -8125
rect -806 -8151 -776 -8125
rect -526 -8151 -316 -8125
rect 29 -8151 59 -8125
rect 115 -8151 145 -8125
rect 201 -8151 231 -8125
rect 287 -8151 317 -8125
rect 670 -8151 880 -8125
rect 1213 -8151 1243 -8125
rect 1498 -8151 1708 -8125
rect 1958 -8151 2168 -8125
rect 2420 -8151 2450 -8125
rect 2522 -8151 2622 -8125
rect 2782 -8151 2882 -8125
rect 2947 -8151 2977 -8125
rect 3246 -8151 3456 -8125
rect 4442 -8151 5388 -8125
rect 6466 -8151 6676 -8125
rect 6928 -8151 6958 -8125
rect 7030 -8151 7130 -8125
rect 7290 -8151 7390 -8125
rect 7455 -8151 7485 -8125
rect 7754 -8151 7964 -8125
rect 8216 -8151 8246 -8125
rect 8318 -8151 8418 -8125
rect 8578 -8151 8678 -8125
rect 8743 -8151 8773 -8125
rect 9042 -8151 9252 -8125
rect 9504 -8151 9534 -8125
rect 9606 -8151 9706 -8125
rect 9866 -8151 9966 -8125
rect 10031 -8151 10061 -8125
rect 10330 -8151 10540 -8125
rect 10790 -8151 10820 -8125
rect 10874 -8151 10904 -8125
rect 10958 -8151 10988 -8125
rect 11042 -8151 11072 -8125
rect 11126 -8151 11156 -8125
rect 11210 -8151 11240 -8125
rect 11294 -8151 11324 -8125
rect 11378 -8151 11408 -8125
rect 11710 -8151 11920 -8125
rect 13642 -8151 14588 -8125
rect 14838 -8151 15784 -8125
rect 16034 -8151 16612 -8125
rect -2918 -8219 -2340 -8193
rect -1538 -8219 -960 -8193
rect -802 -8219 -224 -8193
rect 26 -8219 236 -8193
rect 505 -8219 535 -8193
rect 600 -8219 700 -8193
rect 860 -8219 960 -8193
rect 1032 -8219 1062 -8193
rect 1314 -8219 1524 -8193
rect 1774 -8219 2352 -8193
rect 2602 -8219 2812 -8193
rect 3081 -8219 3111 -8193
rect 3176 -8219 3276 -8193
rect 3436 -8219 3536 -8193
rect 3608 -8219 3638 -8193
rect 3890 -8219 4100 -8193
rect 4350 -8219 4928 -8193
rect 5178 -8219 5388 -8193
rect 5657 -8219 5687 -8193
rect 5752 -8219 5852 -8193
rect 6012 -8219 6112 -8193
rect 6184 -8219 6214 -8193
rect 6466 -8219 6676 -8193
rect 6926 -8219 7504 -8193
rect 7754 -8219 7964 -8193
rect 8233 -8219 8263 -8193
rect 8328 -8219 8428 -8193
rect 8588 -8219 8688 -8193
rect 8760 -8219 8790 -8193
rect 9042 -8219 9252 -8193
rect 9502 -8219 10080 -8193
rect 10422 -8219 10632 -8193
rect 10809 -8219 10839 -8193
rect 10904 -8219 11004 -8193
rect 11164 -8219 11264 -8193
rect 11336 -8219 11366 -8193
rect 11710 -8219 11920 -8193
rect 13735 -8219 13765 -8193
rect 13821 -8219 13851 -8193
rect 13907 -8219 13937 -8193
rect 13993 -8219 14023 -8193
rect 14079 -8219 14109 -8193
rect 14165 -8219 14195 -8193
rect 14251 -8219 14281 -8193
rect 14337 -8219 14367 -8193
rect 14423 -8219 14453 -8193
rect 14509 -8219 14539 -8193
rect 14595 -8219 14625 -8193
rect 14681 -8219 14711 -8193
rect 14766 -8219 14796 -8193
rect 14852 -8219 14882 -8193
rect 14938 -8219 14968 -8193
rect 15024 -8219 15054 -8193
rect 15110 -8219 15140 -8193
rect 15196 -8219 15226 -8193
rect 15282 -8219 15312 -8193
rect 15368 -8219 15398 -8193
rect 15666 -8219 16612 -8193
rect -2918 -8355 -2340 -8329
rect -1538 -8355 -960 -8329
rect -802 -8355 -224 -8329
rect 26 -8355 236 -8329
rect -2918 -8377 -2646 -8355
rect -2918 -8411 -2902 -8377
rect -2868 -8411 -2799 -8377
rect -2765 -8411 -2696 -8377
rect -2662 -8411 -2646 -8377
rect -1538 -8377 -1266 -8355
rect -2918 -8427 -2646 -8411
rect -2604 -8413 -2340 -8397
rect -2604 -8447 -2588 -8413
rect -2554 -8447 -2489 -8413
rect -2455 -8447 -2390 -8413
rect -2356 -8447 -2340 -8413
rect -1538 -8411 -1522 -8377
rect -1488 -8411 -1419 -8377
rect -1385 -8411 -1316 -8377
rect -1282 -8411 -1266 -8377
rect -802 -8377 -530 -8355
rect 26 -8361 110 -8355
rect -1538 -8427 -1266 -8411
rect -1224 -8413 -960 -8397
rect -2604 -8469 -2340 -8447
rect -1224 -8447 -1208 -8413
rect -1174 -8447 -1109 -8413
rect -1075 -8447 -1010 -8413
rect -976 -8447 -960 -8413
rect -802 -8411 -786 -8377
rect -752 -8411 -683 -8377
rect -649 -8411 -580 -8377
rect -546 -8411 -530 -8377
rect -32 -8377 110 -8361
rect 505 -8371 535 -8303
rect -802 -8427 -530 -8411
rect -488 -8413 -224 -8397
rect -1224 -8469 -960 -8447
rect -488 -8447 -472 -8413
rect -438 -8447 -373 -8413
rect -339 -8447 -274 -8413
rect -240 -8447 -224 -8413
rect -32 -8411 -16 -8377
rect 18 -8411 110 -8377
rect 501 -8387 555 -8371
rect -32 -8427 110 -8411
rect 152 -8413 294 -8397
rect -488 -8469 -224 -8447
rect 152 -8447 244 -8413
rect 278 -8447 294 -8413
rect 501 -8421 511 -8387
rect 545 -8421 555 -8387
rect 501 -8437 555 -8421
rect 600 -8377 700 -8349
rect 860 -8377 960 -8349
rect 1032 -8375 1062 -8303
rect 1314 -8355 1524 -8329
rect 1774 -8355 2352 -8329
rect 2602 -8355 2812 -8329
rect 1314 -8361 1398 -8355
rect 600 -8387 761 -8377
rect 600 -8421 711 -8387
rect 745 -8421 761 -8387
rect 600 -8431 761 -8421
rect 860 -8387 982 -8377
rect 860 -8421 932 -8387
rect 966 -8421 982 -8387
rect 860 -8431 982 -8421
rect 1032 -8387 1102 -8375
rect 1032 -8421 1052 -8387
rect 1086 -8421 1102 -8387
rect 152 -8463 294 -8447
rect 152 -8469 236 -8463
rect 505 -8469 535 -8437
rect -2918 -8495 -2340 -8469
rect -1538 -8495 -960 -8469
rect -802 -8495 -224 -8469
rect 26 -8495 236 -8469
rect 600 -8505 700 -8431
rect 860 -8505 960 -8431
rect 1032 -8434 1102 -8421
rect 1256 -8377 1398 -8361
rect 1256 -8411 1272 -8377
rect 1306 -8411 1398 -8377
rect 1774 -8377 2046 -8355
rect 2602 -8361 2686 -8355
rect 1256 -8427 1398 -8411
rect 1440 -8413 1582 -8397
rect 1032 -8469 1062 -8434
rect 1440 -8447 1532 -8413
rect 1566 -8447 1582 -8413
rect 1774 -8411 1790 -8377
rect 1824 -8411 1893 -8377
rect 1927 -8411 1996 -8377
rect 2030 -8411 2046 -8377
rect 2544 -8377 2686 -8361
rect 3081 -8371 3111 -8303
rect 1774 -8427 2046 -8411
rect 2088 -8413 2352 -8397
rect 1440 -8463 1582 -8447
rect 2088 -8447 2104 -8413
rect 2138 -8447 2203 -8413
rect 2237 -8447 2302 -8413
rect 2336 -8447 2352 -8413
rect 2544 -8411 2560 -8377
rect 2594 -8411 2686 -8377
rect 3077 -8387 3131 -8371
rect 2544 -8427 2686 -8411
rect 2728 -8413 2870 -8397
rect 1440 -8469 1524 -8463
rect 2088 -8469 2352 -8447
rect 2728 -8447 2820 -8413
rect 2854 -8447 2870 -8413
rect 3077 -8421 3087 -8387
rect 3121 -8421 3131 -8387
rect 3077 -8437 3131 -8421
rect 3176 -8377 3276 -8349
rect 3436 -8377 3536 -8349
rect 3608 -8375 3638 -8303
rect 3890 -8355 4100 -8329
rect 4350 -8355 4928 -8329
rect 5178 -8355 5388 -8329
rect 3890 -8361 3974 -8355
rect 3176 -8387 3337 -8377
rect 3176 -8421 3287 -8387
rect 3321 -8421 3337 -8387
rect 3176 -8431 3337 -8421
rect 3436 -8387 3558 -8377
rect 3436 -8421 3508 -8387
rect 3542 -8421 3558 -8387
rect 3436 -8431 3558 -8421
rect 3608 -8387 3678 -8375
rect 3608 -8421 3628 -8387
rect 3662 -8421 3678 -8387
rect 2728 -8463 2870 -8447
rect 2728 -8469 2812 -8463
rect 3081 -8469 3111 -8437
rect 1314 -8495 1524 -8469
rect 1774 -8495 2352 -8469
rect 2602 -8495 2812 -8469
rect 3176 -8505 3276 -8431
rect 3436 -8505 3536 -8431
rect 3608 -8434 3678 -8421
rect 3832 -8377 3974 -8361
rect 3832 -8411 3848 -8377
rect 3882 -8411 3974 -8377
rect 4350 -8377 4622 -8355
rect 5178 -8361 5262 -8355
rect 3832 -8427 3974 -8411
rect 4016 -8413 4158 -8397
rect 3608 -8469 3638 -8434
rect 4016 -8447 4108 -8413
rect 4142 -8447 4158 -8413
rect 4350 -8411 4366 -8377
rect 4400 -8411 4469 -8377
rect 4503 -8411 4572 -8377
rect 4606 -8411 4622 -8377
rect 5120 -8377 5262 -8361
rect 5657 -8371 5687 -8303
rect 4350 -8427 4622 -8411
rect 4664 -8413 4928 -8397
rect 4016 -8463 4158 -8447
rect 4664 -8447 4680 -8413
rect 4714 -8447 4779 -8413
rect 4813 -8447 4878 -8413
rect 4912 -8447 4928 -8413
rect 5120 -8411 5136 -8377
rect 5170 -8411 5262 -8377
rect 5653 -8387 5707 -8371
rect 5120 -8427 5262 -8411
rect 5304 -8413 5446 -8397
rect 4016 -8469 4100 -8463
rect 4664 -8469 4928 -8447
rect 5304 -8447 5396 -8413
rect 5430 -8447 5446 -8413
rect 5653 -8421 5663 -8387
rect 5697 -8421 5707 -8387
rect 5653 -8437 5707 -8421
rect 5752 -8377 5852 -8349
rect 6012 -8377 6112 -8349
rect 6184 -8375 6214 -8303
rect 6466 -8355 6676 -8329
rect 6926 -8355 7504 -8329
rect 7754 -8355 7964 -8329
rect 6466 -8361 6550 -8355
rect 5752 -8387 5913 -8377
rect 5752 -8421 5863 -8387
rect 5897 -8421 5913 -8387
rect 5752 -8431 5913 -8421
rect 6012 -8387 6134 -8377
rect 6012 -8421 6084 -8387
rect 6118 -8421 6134 -8387
rect 6012 -8431 6134 -8421
rect 6184 -8387 6254 -8375
rect 6184 -8421 6204 -8387
rect 6238 -8421 6254 -8387
rect 5304 -8463 5446 -8447
rect 5304 -8469 5388 -8463
rect 5657 -8469 5687 -8437
rect 3890 -8495 4100 -8469
rect 4350 -8495 4928 -8469
rect 5178 -8495 5388 -8469
rect 5752 -8505 5852 -8431
rect 6012 -8505 6112 -8431
rect 6184 -8434 6254 -8421
rect 6408 -8377 6550 -8361
rect 6408 -8411 6424 -8377
rect 6458 -8411 6550 -8377
rect 6926 -8377 7198 -8355
rect 7754 -8361 7838 -8355
rect 6408 -8427 6550 -8411
rect 6592 -8413 6734 -8397
rect 6184 -8469 6214 -8434
rect 6592 -8447 6684 -8413
rect 6718 -8447 6734 -8413
rect 6926 -8411 6942 -8377
rect 6976 -8411 7045 -8377
rect 7079 -8411 7148 -8377
rect 7182 -8411 7198 -8377
rect 7696 -8377 7838 -8361
rect 8233 -8371 8263 -8303
rect 6926 -8427 7198 -8411
rect 7240 -8413 7504 -8397
rect 6592 -8463 6734 -8447
rect 7240 -8447 7256 -8413
rect 7290 -8447 7355 -8413
rect 7389 -8447 7454 -8413
rect 7488 -8447 7504 -8413
rect 7696 -8411 7712 -8377
rect 7746 -8411 7838 -8377
rect 8229 -8387 8283 -8371
rect 7696 -8427 7838 -8411
rect 7880 -8413 8022 -8397
rect 6592 -8469 6676 -8463
rect 7240 -8469 7504 -8447
rect 7880 -8447 7972 -8413
rect 8006 -8447 8022 -8413
rect 8229 -8421 8239 -8387
rect 8273 -8421 8283 -8387
rect 8229 -8437 8283 -8421
rect 8328 -8377 8428 -8349
rect 8588 -8377 8688 -8349
rect 8760 -8375 8790 -8303
rect 9042 -8355 9252 -8329
rect 9502 -8355 10080 -8329
rect 10422 -8355 10632 -8329
rect 9042 -8361 9126 -8355
rect 8328 -8387 8489 -8377
rect 8328 -8421 8439 -8387
rect 8473 -8421 8489 -8387
rect 8328 -8431 8489 -8421
rect 8588 -8387 8710 -8377
rect 8588 -8421 8660 -8387
rect 8694 -8421 8710 -8387
rect 8588 -8431 8710 -8421
rect 8760 -8387 8830 -8375
rect 8760 -8421 8780 -8387
rect 8814 -8421 8830 -8387
rect 7880 -8463 8022 -8447
rect 7880 -8469 7964 -8463
rect 8233 -8469 8263 -8437
rect 6466 -8495 6676 -8469
rect 6926 -8495 7504 -8469
rect 7754 -8495 7964 -8469
rect 8328 -8505 8428 -8431
rect 8588 -8505 8688 -8431
rect 8760 -8434 8830 -8421
rect 8984 -8377 9126 -8361
rect 8984 -8411 9000 -8377
rect 9034 -8411 9126 -8377
rect 9502 -8377 9774 -8355
rect 10422 -8361 10506 -8355
rect 8984 -8427 9126 -8411
rect 9168 -8413 9310 -8397
rect 8760 -8469 8790 -8434
rect 9168 -8447 9260 -8413
rect 9294 -8447 9310 -8413
rect 9502 -8411 9518 -8377
rect 9552 -8411 9621 -8377
rect 9655 -8411 9724 -8377
rect 9758 -8411 9774 -8377
rect 10364 -8377 10506 -8361
rect 10809 -8371 10839 -8303
rect 9502 -8427 9774 -8411
rect 9816 -8413 10080 -8397
rect 9168 -8463 9310 -8447
rect 9816 -8447 9832 -8413
rect 9866 -8447 9931 -8413
rect 9965 -8447 10030 -8413
rect 10064 -8447 10080 -8413
rect 10364 -8411 10380 -8377
rect 10414 -8411 10506 -8377
rect 10805 -8387 10859 -8371
rect 10364 -8427 10506 -8411
rect 10548 -8413 10690 -8397
rect 9168 -8469 9252 -8463
rect 9816 -8469 10080 -8447
rect 10548 -8447 10640 -8413
rect 10674 -8447 10690 -8413
rect 10805 -8421 10815 -8387
rect 10849 -8421 10859 -8387
rect 10805 -8437 10859 -8421
rect 10904 -8377 11004 -8349
rect 11164 -8377 11264 -8349
rect 11336 -8375 11366 -8303
rect 11710 -8355 11920 -8329
rect 13735 -8352 13765 -8303
rect 13821 -8352 13851 -8303
rect 13907 -8352 13937 -8303
rect 13993 -8352 14023 -8303
rect 11710 -8361 11794 -8355
rect 10904 -8387 11065 -8377
rect 10904 -8421 11015 -8387
rect 11049 -8421 11065 -8387
rect 10904 -8431 11065 -8421
rect 11164 -8387 11286 -8377
rect 11164 -8421 11236 -8387
rect 11270 -8421 11286 -8387
rect 11164 -8431 11286 -8421
rect 11336 -8387 11406 -8375
rect 11336 -8421 11356 -8387
rect 11390 -8421 11406 -8387
rect 10548 -8463 10690 -8447
rect 10548 -8469 10632 -8463
rect 10809 -8469 10839 -8437
rect 9042 -8495 9252 -8469
rect 9502 -8495 10080 -8469
rect 10422 -8495 10632 -8469
rect 10904 -8505 11004 -8431
rect 11164 -8505 11264 -8431
rect 11336 -8434 11406 -8421
rect 11652 -8377 11794 -8361
rect 11652 -8411 11668 -8377
rect 11702 -8411 11794 -8377
rect 13676 -8387 14023 -8352
rect 11652 -8427 11794 -8411
rect 11836 -8413 11978 -8397
rect 11336 -8469 11366 -8434
rect 11836 -8447 11928 -8413
rect 11962 -8447 11978 -8413
rect 11836 -8463 11978 -8447
rect 13676 -8421 13692 -8387
rect 13726 -8421 14023 -8387
rect 13676 -8454 14023 -8421
rect 11836 -8469 11920 -8463
rect 13735 -8469 13765 -8454
rect 13821 -8469 13851 -8454
rect 13907 -8469 13937 -8454
rect 13993 -8469 14023 -8454
rect 14079 -8362 14109 -8303
rect 14165 -8362 14195 -8303
rect 14251 -8362 14281 -8303
rect 14337 -8362 14367 -8303
rect 14423 -8362 14453 -8303
rect 14509 -8362 14539 -8303
rect 14595 -8362 14625 -8303
rect 14681 -8362 14711 -8303
rect 14766 -8362 14796 -8303
rect 14852 -8362 14882 -8303
rect 14938 -8362 14968 -8303
rect 15024 -8362 15054 -8303
rect 15110 -8362 15140 -8303
rect 15196 -8362 15226 -8303
rect 15282 -8362 15312 -8303
rect 15368 -8362 15398 -8303
rect 14079 -8387 15398 -8362
rect 14079 -8421 14119 -8387
rect 14153 -8421 14187 -8387
rect 14221 -8421 14255 -8387
rect 14289 -8421 14323 -8387
rect 14357 -8421 14391 -8387
rect 14425 -8421 14459 -8387
rect 14493 -8421 14527 -8387
rect 14561 -8421 14595 -8387
rect 14629 -8421 14663 -8387
rect 14697 -8421 14731 -8387
rect 14765 -8421 14799 -8387
rect 14833 -8421 14867 -8387
rect 14901 -8421 14935 -8387
rect 14969 -8421 15003 -8387
rect 15037 -8421 15071 -8387
rect 15105 -8421 15139 -8387
rect 15173 -8421 15398 -8387
rect 14079 -8437 15398 -8421
rect 15666 -8355 16612 -8329
rect 15666 -8377 16120 -8355
rect 15666 -8411 15686 -8377
rect 15720 -8411 15814 -8377
rect 15848 -8411 15942 -8377
rect 15976 -8411 16070 -8377
rect 16104 -8411 16120 -8377
rect 15666 -8427 16120 -8411
rect 16162 -8413 16612 -8397
rect 14079 -8469 14109 -8437
rect 14165 -8469 14195 -8437
rect 14251 -8469 14281 -8437
rect 14337 -8469 14367 -8437
rect 14423 -8469 14453 -8437
rect 14509 -8469 14539 -8437
rect 14595 -8469 14625 -8437
rect 14681 -8469 14711 -8437
rect 14766 -8469 14796 -8437
rect 14852 -8469 14882 -8437
rect 14938 -8469 14968 -8437
rect 15024 -8469 15054 -8437
rect 15110 -8469 15140 -8437
rect 15196 -8469 15226 -8437
rect 15282 -8469 15312 -8437
rect 15368 -8469 15398 -8437
rect 16162 -8447 16178 -8413
rect 16212 -8447 16306 -8413
rect 16340 -8447 16434 -8413
rect 16468 -8447 16562 -8413
rect 16596 -8447 16612 -8413
rect 16162 -8469 16612 -8447
rect 11710 -8495 11920 -8469
rect 15666 -8495 16612 -8469
rect -2918 -8695 -2340 -8669
rect -1538 -8695 -960 -8669
rect -802 -8695 -224 -8669
rect 26 -8695 236 -8669
rect 505 -8695 535 -8669
rect 600 -8695 700 -8669
rect 860 -8695 960 -8669
rect 1032 -8695 1062 -8669
rect 1314 -8695 1524 -8669
rect 1774 -8695 2352 -8669
rect 2602 -8695 2812 -8669
rect 3081 -8695 3111 -8669
rect 3176 -8695 3276 -8669
rect 3436 -8695 3536 -8669
rect 3608 -8695 3638 -8669
rect 3890 -8695 4100 -8669
rect 4350 -8695 4928 -8669
rect 5178 -8695 5388 -8669
rect 5657 -8695 5687 -8669
rect 5752 -8695 5852 -8669
rect 6012 -8695 6112 -8669
rect 6184 -8695 6214 -8669
rect 6466 -8695 6676 -8669
rect 6926 -8695 7504 -8669
rect 7754 -8695 7964 -8669
rect 8233 -8695 8263 -8669
rect 8328 -8695 8428 -8669
rect 8588 -8695 8688 -8669
rect 8760 -8695 8790 -8669
rect 9042 -8695 9252 -8669
rect 9502 -8695 10080 -8669
rect 10422 -8695 10632 -8669
rect 10809 -8695 10839 -8669
rect 10904 -8695 11004 -8669
rect 11164 -8695 11264 -8669
rect 11336 -8695 11366 -8669
rect 11710 -8695 11920 -8669
rect 13735 -8695 13765 -8669
rect 13821 -8695 13851 -8669
rect 13907 -8695 13937 -8669
rect 13993 -8695 14023 -8669
rect 14079 -8695 14109 -8669
rect 14165 -8695 14195 -8669
rect 14251 -8695 14281 -8669
rect 14337 -8695 14367 -8669
rect 14423 -8695 14453 -8669
rect 14509 -8695 14539 -8669
rect 14595 -8695 14625 -8669
rect 14681 -8695 14711 -8669
rect 14766 -8695 14796 -8669
rect 14852 -8695 14882 -8669
rect 14938 -8695 14968 -8669
rect 15024 -8695 15054 -8669
rect 15110 -8695 15140 -8669
rect 15196 -8695 15226 -8669
rect 15282 -8695 15312 -8669
rect 15368 -8695 15398 -8669
rect 15666 -8695 16612 -8669
rect -2918 -8763 -2340 -8737
rect -1538 -8763 -960 -8737
rect -802 -8763 -224 -8737
rect 26 -8763 236 -8737
rect 488 -8763 518 -8737
rect 590 -8763 690 -8737
rect 850 -8763 950 -8737
rect 1015 -8763 1045 -8737
rect 1314 -8763 1524 -8737
rect 1774 -8763 2352 -8737
rect 2602 -8763 2812 -8737
rect 3064 -8763 3094 -8737
rect 3166 -8763 3266 -8737
rect 3426 -8763 3526 -8737
rect 3591 -8763 3621 -8737
rect 3890 -8763 4100 -8737
rect 4350 -8763 4928 -8737
rect 5178 -8763 5388 -8737
rect 5640 -8763 5670 -8737
rect 5742 -8763 5842 -8737
rect 6002 -8763 6102 -8737
rect 6167 -8763 6197 -8737
rect 6466 -8763 6676 -8737
rect 6926 -8763 7504 -8737
rect 7754 -8763 7964 -8737
rect 8216 -8763 8246 -8737
rect 8318 -8763 8418 -8737
rect 8578 -8763 8678 -8737
rect 8743 -8763 8773 -8737
rect 9042 -8763 9252 -8737
rect 9502 -8763 10080 -8737
rect 10422 -8763 10632 -8737
rect 10792 -8763 10822 -8737
rect 10894 -8763 10994 -8737
rect 11154 -8763 11254 -8737
rect 11319 -8763 11349 -8737
rect 11710 -8763 11920 -8737
rect 12547 -8763 12577 -8737
rect 12633 -8763 12663 -8737
rect 12719 -8763 12749 -8737
rect 12805 -8763 12835 -8737
rect 12891 -8763 12921 -8737
rect 12977 -8763 13007 -8737
rect 13274 -8763 13484 -8737
rect 13735 -8763 13765 -8737
rect 13821 -8763 13851 -8737
rect 13907 -8763 13937 -8737
rect 13993 -8763 14023 -8737
rect 14079 -8763 14109 -8737
rect 14165 -8763 14195 -8737
rect 14251 -8763 14281 -8737
rect 14337 -8763 14367 -8737
rect 14423 -8763 14453 -8737
rect 14509 -8763 14539 -8737
rect 14595 -8763 14625 -8737
rect 14681 -8763 14711 -8737
rect 14766 -8763 14796 -8737
rect 14852 -8763 14882 -8737
rect 14938 -8763 14968 -8737
rect 15024 -8763 15054 -8737
rect 15110 -8763 15140 -8737
rect 15196 -8763 15226 -8737
rect 15282 -8763 15312 -8737
rect 15368 -8763 15398 -8737
rect 15666 -8763 16612 -8737
rect -2918 -8963 -2340 -8937
rect -1538 -8963 -960 -8937
rect -802 -8963 -224 -8937
rect 26 -8963 236 -8937
rect -2918 -8985 -2654 -8963
rect -2918 -9019 -2902 -8985
rect -2868 -9019 -2803 -8985
rect -2769 -9019 -2704 -8985
rect -2670 -9019 -2654 -8985
rect -1538 -8985 -1274 -8963
rect -2918 -9035 -2654 -9019
rect -2612 -9021 -2340 -9005
rect -2612 -9055 -2596 -9021
rect -2562 -9055 -2493 -9021
rect -2459 -9055 -2390 -9021
rect -2356 -9055 -2340 -9021
rect -1538 -9019 -1522 -8985
rect -1488 -9019 -1423 -8985
rect -1389 -9019 -1324 -8985
rect -1290 -9019 -1274 -8985
rect -802 -8985 -538 -8963
rect -1538 -9035 -1274 -9019
rect -1232 -9021 -960 -9005
rect -2612 -9077 -2340 -9055
rect -1232 -9055 -1216 -9021
rect -1182 -9055 -1113 -9021
rect -1079 -9055 -1010 -9021
rect -976 -9055 -960 -9021
rect -802 -9019 -786 -8985
rect -752 -9019 -687 -8985
rect -653 -9019 -588 -8985
rect -554 -9019 -538 -8985
rect 152 -8969 236 -8963
rect 152 -8985 294 -8969
rect -802 -9035 -538 -9019
rect -496 -9021 -224 -9005
rect -1232 -9077 -960 -9055
rect -496 -9055 -480 -9021
rect -446 -9055 -377 -9021
rect -343 -9055 -274 -9021
rect -240 -9055 -224 -9021
rect -496 -9077 -224 -9055
rect -32 -9021 110 -9005
rect -32 -9055 -16 -9021
rect 18 -9055 110 -9021
rect 152 -9019 244 -8985
rect 278 -9019 294 -8985
rect 488 -8998 518 -8963
rect 152 -9035 294 -9019
rect 448 -9011 518 -8998
rect 590 -9001 690 -8927
rect 850 -9001 950 -8927
rect 1314 -8963 1524 -8937
rect 1015 -8995 1045 -8963
rect 1440 -8969 1524 -8963
rect 1774 -8963 2352 -8937
rect 2602 -8963 2812 -8937
rect 1440 -8985 1582 -8969
rect -32 -9071 110 -9055
rect 448 -9045 464 -9011
rect 498 -9045 518 -9011
rect 448 -9057 518 -9045
rect 568 -9011 690 -9001
rect 568 -9045 584 -9011
rect 618 -9045 690 -9011
rect 568 -9055 690 -9045
rect 789 -9011 950 -9001
rect 789 -9045 805 -9011
rect 839 -9045 950 -9011
rect 789 -9055 950 -9045
rect -2918 -9103 -2340 -9077
rect -1538 -9103 -960 -9077
rect -802 -9103 -224 -9077
rect 26 -9077 110 -9071
rect 26 -9103 236 -9077
rect 488 -9129 518 -9057
rect 590 -9083 690 -9055
rect 850 -9083 950 -9055
rect 995 -9011 1049 -8995
rect 995 -9045 1005 -9011
rect 1039 -9045 1049 -9011
rect 995 -9061 1049 -9045
rect 1256 -9021 1398 -9005
rect 1256 -9055 1272 -9021
rect 1306 -9055 1398 -9021
rect 1440 -9019 1532 -8985
rect 1566 -9019 1582 -8985
rect 1440 -9035 1582 -9019
rect 1774 -8985 2038 -8963
rect 1774 -9019 1790 -8985
rect 1824 -9019 1889 -8985
rect 1923 -9019 1988 -8985
rect 2022 -9019 2038 -8985
rect 2728 -8969 2812 -8963
rect 2728 -8985 2870 -8969
rect 1774 -9035 2038 -9019
rect 2080 -9021 2352 -9005
rect 1015 -9129 1045 -9061
rect 1256 -9071 1398 -9055
rect 1314 -9077 1398 -9071
rect 2080 -9055 2096 -9021
rect 2130 -9055 2199 -9021
rect 2233 -9055 2302 -9021
rect 2336 -9055 2352 -9021
rect 2080 -9077 2352 -9055
rect 2544 -9021 2686 -9005
rect 2544 -9055 2560 -9021
rect 2594 -9055 2686 -9021
rect 2728 -9019 2820 -8985
rect 2854 -9019 2870 -8985
rect 3064 -8998 3094 -8963
rect 2728 -9035 2870 -9019
rect 3024 -9011 3094 -8998
rect 3166 -9001 3266 -8927
rect 3426 -9001 3526 -8927
rect 3890 -8963 4100 -8937
rect 3591 -8995 3621 -8963
rect 4016 -8969 4100 -8963
rect 4350 -8963 4928 -8937
rect 5178 -8963 5388 -8937
rect 4016 -8985 4158 -8969
rect 2544 -9071 2686 -9055
rect 3024 -9045 3040 -9011
rect 3074 -9045 3094 -9011
rect 3024 -9057 3094 -9045
rect 3144 -9011 3266 -9001
rect 3144 -9045 3160 -9011
rect 3194 -9045 3266 -9011
rect 3144 -9055 3266 -9045
rect 3365 -9011 3526 -9001
rect 3365 -9045 3381 -9011
rect 3415 -9045 3526 -9011
rect 3365 -9055 3526 -9045
rect 1314 -9103 1524 -9077
rect 1774 -9103 2352 -9077
rect 2602 -9077 2686 -9071
rect 2602 -9103 2812 -9077
rect 3064 -9129 3094 -9057
rect 3166 -9083 3266 -9055
rect 3426 -9083 3526 -9055
rect 3571 -9011 3625 -8995
rect 3571 -9045 3581 -9011
rect 3615 -9045 3625 -9011
rect 3571 -9061 3625 -9045
rect 3832 -9021 3974 -9005
rect 3832 -9055 3848 -9021
rect 3882 -9055 3974 -9021
rect 4016 -9019 4108 -8985
rect 4142 -9019 4158 -8985
rect 4016 -9035 4158 -9019
rect 4350 -8985 4614 -8963
rect 4350 -9019 4366 -8985
rect 4400 -9019 4465 -8985
rect 4499 -9019 4564 -8985
rect 4598 -9019 4614 -8985
rect 5304 -8969 5388 -8963
rect 5304 -8985 5446 -8969
rect 4350 -9035 4614 -9019
rect 4656 -9021 4928 -9005
rect 3591 -9129 3621 -9061
rect 3832 -9071 3974 -9055
rect 3890 -9077 3974 -9071
rect 4656 -9055 4672 -9021
rect 4706 -9055 4775 -9021
rect 4809 -9055 4878 -9021
rect 4912 -9055 4928 -9021
rect 4656 -9077 4928 -9055
rect 5120 -9021 5262 -9005
rect 5120 -9055 5136 -9021
rect 5170 -9055 5262 -9021
rect 5304 -9019 5396 -8985
rect 5430 -9019 5446 -8985
rect 5640 -8998 5670 -8963
rect 5304 -9035 5446 -9019
rect 5600 -9011 5670 -8998
rect 5742 -9001 5842 -8927
rect 6002 -9001 6102 -8927
rect 6466 -8963 6676 -8937
rect 6167 -8995 6197 -8963
rect 6592 -8969 6676 -8963
rect 6926 -8963 7504 -8937
rect 7754 -8963 7964 -8937
rect 6592 -8985 6734 -8969
rect 5120 -9071 5262 -9055
rect 5600 -9045 5616 -9011
rect 5650 -9045 5670 -9011
rect 5600 -9057 5670 -9045
rect 5720 -9011 5842 -9001
rect 5720 -9045 5736 -9011
rect 5770 -9045 5842 -9011
rect 5720 -9055 5842 -9045
rect 5941 -9011 6102 -9001
rect 5941 -9045 5957 -9011
rect 5991 -9045 6102 -9011
rect 5941 -9055 6102 -9045
rect 3890 -9103 4100 -9077
rect 4350 -9103 4928 -9077
rect 5178 -9077 5262 -9071
rect 5178 -9103 5388 -9077
rect 5640 -9129 5670 -9057
rect 5742 -9083 5842 -9055
rect 6002 -9083 6102 -9055
rect 6147 -9011 6201 -8995
rect 6147 -9045 6157 -9011
rect 6191 -9045 6201 -9011
rect 6147 -9061 6201 -9045
rect 6408 -9021 6550 -9005
rect 6408 -9055 6424 -9021
rect 6458 -9055 6550 -9021
rect 6592 -9019 6684 -8985
rect 6718 -9019 6734 -8985
rect 6592 -9035 6734 -9019
rect 6926 -8985 7190 -8963
rect 6926 -9019 6942 -8985
rect 6976 -9019 7041 -8985
rect 7075 -9019 7140 -8985
rect 7174 -9019 7190 -8985
rect 7880 -8969 7964 -8963
rect 7880 -8985 8022 -8969
rect 6926 -9035 7190 -9019
rect 7232 -9021 7504 -9005
rect 6167 -9129 6197 -9061
rect 6408 -9071 6550 -9055
rect 6466 -9077 6550 -9071
rect 7232 -9055 7248 -9021
rect 7282 -9055 7351 -9021
rect 7385 -9055 7454 -9021
rect 7488 -9055 7504 -9021
rect 7232 -9077 7504 -9055
rect 7696 -9021 7838 -9005
rect 7696 -9055 7712 -9021
rect 7746 -9055 7838 -9021
rect 7880 -9019 7972 -8985
rect 8006 -9019 8022 -8985
rect 8216 -8998 8246 -8963
rect 7880 -9035 8022 -9019
rect 8176 -9011 8246 -8998
rect 8318 -9001 8418 -8927
rect 8578 -9001 8678 -8927
rect 9042 -8963 9252 -8937
rect 8743 -8995 8773 -8963
rect 9168 -8969 9252 -8963
rect 9502 -8963 10080 -8937
rect 10422 -8963 10632 -8937
rect 9168 -8985 9310 -8969
rect 7696 -9071 7838 -9055
rect 8176 -9045 8192 -9011
rect 8226 -9045 8246 -9011
rect 8176 -9057 8246 -9045
rect 8296 -9011 8418 -9001
rect 8296 -9045 8312 -9011
rect 8346 -9045 8418 -9011
rect 8296 -9055 8418 -9045
rect 8517 -9011 8678 -9001
rect 8517 -9045 8533 -9011
rect 8567 -9045 8678 -9011
rect 8517 -9055 8678 -9045
rect 6466 -9103 6676 -9077
rect 6926 -9103 7504 -9077
rect 7754 -9077 7838 -9071
rect 7754 -9103 7964 -9077
rect 8216 -9129 8246 -9057
rect 8318 -9083 8418 -9055
rect 8578 -9083 8678 -9055
rect 8723 -9011 8777 -8995
rect 8723 -9045 8733 -9011
rect 8767 -9045 8777 -9011
rect 8723 -9061 8777 -9045
rect 8984 -9021 9126 -9005
rect 8984 -9055 9000 -9021
rect 9034 -9055 9126 -9021
rect 9168 -9019 9260 -8985
rect 9294 -9019 9310 -8985
rect 9168 -9035 9310 -9019
rect 9502 -8985 9766 -8963
rect 9502 -9019 9518 -8985
rect 9552 -9019 9617 -8985
rect 9651 -9019 9716 -8985
rect 9750 -9019 9766 -8985
rect 10548 -8969 10632 -8963
rect 10548 -8985 10690 -8969
rect 9502 -9035 9766 -9019
rect 9808 -9021 10080 -9005
rect 8743 -9129 8773 -9061
rect 8984 -9071 9126 -9055
rect 9042 -9077 9126 -9071
rect 9808 -9055 9824 -9021
rect 9858 -9055 9927 -9021
rect 9961 -9055 10030 -9021
rect 10064 -9055 10080 -9021
rect 9808 -9077 10080 -9055
rect 10364 -9021 10506 -9005
rect 10364 -9055 10380 -9021
rect 10414 -9055 10506 -9021
rect 10548 -9019 10640 -8985
rect 10674 -9019 10690 -8985
rect 10792 -8998 10822 -8963
rect 10548 -9035 10690 -9019
rect 10752 -9011 10822 -8998
rect 10894 -9001 10994 -8927
rect 11154 -9001 11254 -8927
rect 11710 -8963 11920 -8937
rect 13274 -8963 13484 -8937
rect 15666 -8963 16612 -8937
rect 11319 -8995 11349 -8963
rect 11836 -8969 11920 -8963
rect 11836 -8985 11978 -8969
rect 10364 -9071 10506 -9055
rect 10752 -9045 10768 -9011
rect 10802 -9045 10822 -9011
rect 10752 -9057 10822 -9045
rect 10872 -9011 10994 -9001
rect 10872 -9045 10888 -9011
rect 10922 -9045 10994 -9011
rect 10872 -9055 10994 -9045
rect 11093 -9011 11254 -9001
rect 11093 -9045 11109 -9011
rect 11143 -9045 11254 -9011
rect 11093 -9055 11254 -9045
rect 9042 -9103 9252 -9077
rect 9502 -9103 10080 -9077
rect 10422 -9077 10506 -9071
rect 10422 -9103 10632 -9077
rect 10792 -9129 10822 -9057
rect 10894 -9083 10994 -9055
rect 11154 -9083 11254 -9055
rect 11299 -9011 11353 -8995
rect 11299 -9045 11309 -9011
rect 11343 -9045 11353 -9011
rect 11299 -9061 11353 -9045
rect 11652 -9021 11794 -9005
rect 11652 -9055 11668 -9021
rect 11702 -9055 11794 -9021
rect 11836 -9019 11928 -8985
rect 11962 -9019 11978 -8985
rect 11836 -9035 11978 -9019
rect 12547 -9001 12577 -8963
rect 12633 -9001 12663 -8963
rect 12719 -9001 12749 -8963
rect 12805 -9001 12835 -8963
rect 12891 -9001 12921 -8963
rect 12977 -9001 13007 -8963
rect 13274 -8969 13358 -8963
rect 12547 -9011 13007 -9001
rect 12547 -9045 12574 -9011
rect 12608 -9045 12642 -9011
rect 12676 -9045 12710 -9011
rect 12744 -9045 12778 -9011
rect 12812 -9045 12846 -9011
rect 12880 -9045 12914 -9011
rect 12948 -9045 13007 -9011
rect 13216 -8985 13358 -8969
rect 13735 -8978 13765 -8963
rect 13821 -8978 13851 -8963
rect 13907 -8978 13937 -8963
rect 13993 -8978 14023 -8963
rect 13216 -9019 13232 -8985
rect 13266 -9019 13358 -8985
rect 13216 -9035 13358 -9019
rect 13400 -9021 13542 -9005
rect 12547 -9055 13007 -9045
rect 13400 -9055 13492 -9021
rect 13526 -9055 13542 -9021
rect 11319 -9129 11349 -9061
rect 11652 -9071 11794 -9055
rect 11710 -9077 11794 -9071
rect 11710 -9103 11920 -9077
rect 12633 -9129 12663 -9055
rect 12719 -9129 12749 -9055
rect 12805 -9129 12835 -9055
rect 12891 -9129 12921 -9055
rect 13400 -9071 13542 -9055
rect 13676 -9011 14023 -8978
rect 13676 -9045 13692 -9011
rect 13726 -9045 14023 -9011
rect 13400 -9077 13484 -9071
rect 13274 -9103 13484 -9077
rect 13676 -9080 14023 -9045
rect 13735 -9129 13765 -9080
rect 13821 -9129 13851 -9080
rect 13907 -9129 13937 -9080
rect 13993 -9129 14023 -9080
rect 14079 -8995 14109 -8963
rect 14165 -8995 14195 -8963
rect 14251 -8995 14281 -8963
rect 14337 -8995 14367 -8963
rect 14423 -8995 14453 -8963
rect 14509 -8995 14539 -8963
rect 14595 -8995 14625 -8963
rect 14681 -8995 14711 -8963
rect 14766 -8995 14796 -8963
rect 14852 -8995 14882 -8963
rect 14938 -8995 14968 -8963
rect 15024 -8995 15054 -8963
rect 15110 -8995 15140 -8963
rect 15196 -8995 15226 -8963
rect 15282 -8995 15312 -8963
rect 15368 -8995 15398 -8963
rect 14079 -9011 15398 -8995
rect 14079 -9045 14119 -9011
rect 14153 -9045 14187 -9011
rect 14221 -9045 14255 -9011
rect 14289 -9045 14323 -9011
rect 14357 -9045 14391 -9011
rect 14425 -9045 14459 -9011
rect 14493 -9045 14527 -9011
rect 14561 -9045 14595 -9011
rect 14629 -9045 14663 -9011
rect 14697 -9045 14731 -9011
rect 14765 -9045 14799 -9011
rect 14833 -9045 14867 -9011
rect 14901 -9045 14935 -9011
rect 14969 -9045 15003 -9011
rect 15037 -9045 15071 -9011
rect 15105 -9045 15139 -9011
rect 15173 -9045 15398 -9011
rect 15666 -8985 16116 -8963
rect 15666 -9019 15682 -8985
rect 15716 -9019 15810 -8985
rect 15844 -9019 15938 -8985
rect 15972 -9019 16066 -8985
rect 16100 -9019 16116 -8985
rect 15666 -9035 16116 -9019
rect 16158 -9021 16612 -9005
rect 14079 -9070 15398 -9045
rect 14079 -9129 14109 -9070
rect 14165 -9129 14195 -9070
rect 14251 -9129 14281 -9070
rect 14337 -9129 14367 -9070
rect 14423 -9129 14453 -9070
rect 14509 -9129 14539 -9070
rect 14595 -9129 14625 -9070
rect 14681 -9129 14711 -9070
rect 14766 -9129 14796 -9070
rect 14852 -9129 14882 -9070
rect 14938 -9129 14968 -9070
rect 15024 -9129 15054 -9070
rect 15110 -9129 15140 -9070
rect 15196 -9129 15226 -9070
rect 15282 -9129 15312 -9070
rect 15368 -9129 15398 -9070
rect 16158 -9055 16174 -9021
rect 16208 -9055 16302 -9021
rect 16336 -9055 16430 -9021
rect 16464 -9055 16558 -9021
rect 16592 -9055 16612 -9021
rect 16158 -9077 16612 -9055
rect 15666 -9103 16612 -9077
rect -2918 -9239 -2340 -9213
rect -1538 -9239 -960 -9213
rect -802 -9239 -224 -9213
rect 26 -9239 236 -9213
rect 488 -9239 518 -9213
rect 590 -9239 690 -9213
rect 850 -9239 950 -9213
rect 1015 -9239 1045 -9213
rect 1314 -9239 1524 -9213
rect 1774 -9239 2352 -9213
rect 2602 -9239 2812 -9213
rect 3064 -9239 3094 -9213
rect 3166 -9239 3266 -9213
rect 3426 -9239 3526 -9213
rect 3591 -9239 3621 -9213
rect 3890 -9239 4100 -9213
rect 4350 -9239 4928 -9213
rect 5178 -9239 5388 -9213
rect 5640 -9239 5670 -9213
rect 5742 -9239 5842 -9213
rect 6002 -9239 6102 -9213
rect 6167 -9239 6197 -9213
rect 6466 -9239 6676 -9213
rect 6926 -9239 7504 -9213
rect 7754 -9239 7964 -9213
rect 8216 -9239 8246 -9213
rect 8318 -9239 8418 -9213
rect 8578 -9239 8678 -9213
rect 8743 -9239 8773 -9213
rect 9042 -9239 9252 -9213
rect 9502 -9239 10080 -9213
rect 10422 -9239 10632 -9213
rect 10792 -9239 10822 -9213
rect 10894 -9239 10994 -9213
rect 11154 -9239 11254 -9213
rect 11319 -9239 11349 -9213
rect 11710 -9239 11920 -9213
rect 12633 -9239 12663 -9213
rect 12719 -9239 12749 -9213
rect 12805 -9239 12835 -9213
rect 12891 -9239 12921 -9213
rect 13274 -9239 13484 -9213
rect 13735 -9239 13765 -9213
rect 13821 -9239 13851 -9213
rect 13907 -9239 13937 -9213
rect 13993 -9239 14023 -9213
rect 14079 -9239 14109 -9213
rect 14165 -9239 14195 -9213
rect 14251 -9239 14281 -9213
rect 14337 -9239 14367 -9213
rect 14423 -9239 14453 -9213
rect 14509 -9239 14539 -9213
rect 14595 -9239 14625 -9213
rect 14681 -9239 14711 -9213
rect 14766 -9239 14796 -9213
rect 14852 -9239 14882 -9213
rect 14938 -9239 14968 -9213
rect 15024 -9239 15054 -9213
rect 15110 -9239 15140 -9213
rect 15196 -9239 15226 -9213
rect 15282 -9239 15312 -9213
rect 15368 -9239 15398 -9213
rect 15666 -9239 16612 -9213
rect -2918 -9307 -2340 -9281
rect -1538 -9307 -960 -9281
rect -783 -9307 -753 -9281
rect -688 -9307 -588 -9281
rect -428 -9307 -328 -9281
rect -256 -9307 -226 -9281
rect 26 -9307 236 -9281
rect 505 -9307 535 -9281
rect 600 -9307 700 -9281
rect 860 -9307 960 -9281
rect 1032 -9307 1062 -9281
rect 1314 -9307 1524 -9281
rect 1774 -9307 2352 -9281
rect 2602 -9307 2812 -9281
rect 3081 -9307 3111 -9281
rect 3176 -9307 3276 -9281
rect 3436 -9307 3536 -9281
rect 3608 -9307 3638 -9281
rect 3890 -9307 4100 -9281
rect 4350 -9307 4928 -9281
rect 5178 -9307 5388 -9281
rect 5657 -9307 5687 -9281
rect 5752 -9307 5852 -9281
rect 6012 -9307 6112 -9281
rect 6184 -9307 6214 -9281
rect 6466 -9307 6676 -9281
rect 6926 -9307 7504 -9281
rect 7754 -9307 7964 -9281
rect 8233 -9307 8263 -9281
rect 8328 -9307 8428 -9281
rect 8588 -9307 8688 -9281
rect 8760 -9307 8790 -9281
rect 9042 -9307 9252 -9281
rect 9502 -9307 10080 -9281
rect 10422 -9307 10632 -9281
rect 10809 -9307 10839 -9281
rect 10904 -9307 11004 -9281
rect 11164 -9307 11264 -9281
rect 11336 -9307 11366 -9281
rect 11710 -9307 11920 -9281
rect 13735 -9307 13765 -9281
rect 13821 -9307 13851 -9281
rect 13907 -9307 13937 -9281
rect 13993 -9307 14023 -9281
rect 14079 -9307 14109 -9281
rect 14165 -9307 14195 -9281
rect 14251 -9307 14281 -9281
rect 14337 -9307 14367 -9281
rect 14423 -9307 14453 -9281
rect 14509 -9307 14539 -9281
rect 14595 -9307 14625 -9281
rect 14681 -9307 14711 -9281
rect 14766 -9307 14796 -9281
rect 14852 -9307 14882 -9281
rect 14938 -9307 14968 -9281
rect 15024 -9307 15054 -9281
rect 15110 -9307 15140 -9281
rect 15196 -9307 15226 -9281
rect 15282 -9307 15312 -9281
rect 15368 -9307 15398 -9281
rect 15666 -9307 16612 -9281
rect -2918 -9443 -2340 -9417
rect -1538 -9443 -960 -9417
rect -2918 -9465 -2646 -9443
rect -2918 -9499 -2902 -9465
rect -2868 -9499 -2799 -9465
rect -2765 -9499 -2696 -9465
rect -2662 -9499 -2646 -9465
rect -1538 -9465 -1266 -9443
rect -783 -9459 -753 -9391
rect -2918 -9515 -2646 -9499
rect -2604 -9501 -2340 -9485
rect -2604 -9535 -2588 -9501
rect -2554 -9535 -2489 -9501
rect -2455 -9535 -2390 -9501
rect -2356 -9535 -2340 -9501
rect -1538 -9499 -1522 -9465
rect -1488 -9499 -1419 -9465
rect -1385 -9499 -1316 -9465
rect -1282 -9499 -1266 -9465
rect -787 -9475 -733 -9459
rect -1538 -9515 -1266 -9499
rect -1224 -9501 -960 -9485
rect -2604 -9557 -2340 -9535
rect -1224 -9535 -1208 -9501
rect -1174 -9535 -1109 -9501
rect -1075 -9535 -1010 -9501
rect -976 -9535 -960 -9501
rect -787 -9509 -777 -9475
rect -743 -9509 -733 -9475
rect -787 -9525 -733 -9509
rect -688 -9465 -588 -9437
rect -428 -9465 -328 -9437
rect -256 -9463 -226 -9391
rect 26 -9443 236 -9417
rect 26 -9449 110 -9443
rect -688 -9475 -527 -9465
rect -688 -9509 -577 -9475
rect -543 -9509 -527 -9475
rect -688 -9519 -527 -9509
rect -428 -9475 -306 -9465
rect -428 -9509 -356 -9475
rect -322 -9509 -306 -9475
rect -428 -9519 -306 -9509
rect -256 -9475 -186 -9463
rect -256 -9509 -236 -9475
rect -202 -9509 -186 -9475
rect -1224 -9557 -960 -9535
rect -783 -9557 -753 -9525
rect -2918 -9583 -2340 -9557
rect -1538 -9583 -960 -9557
rect -688 -9593 -588 -9519
rect -428 -9593 -328 -9519
rect -256 -9522 -186 -9509
rect -32 -9465 110 -9449
rect 505 -9459 535 -9391
rect -32 -9499 -16 -9465
rect 18 -9499 110 -9465
rect 501 -9475 555 -9459
rect -32 -9515 110 -9499
rect 152 -9501 294 -9485
rect -256 -9557 -226 -9522
rect 152 -9535 244 -9501
rect 278 -9535 294 -9501
rect 501 -9509 511 -9475
rect 545 -9509 555 -9475
rect 501 -9525 555 -9509
rect 600 -9465 700 -9437
rect 860 -9465 960 -9437
rect 1032 -9463 1062 -9391
rect 1314 -9443 1524 -9417
rect 1774 -9443 2352 -9417
rect 2602 -9443 2812 -9417
rect 1314 -9449 1398 -9443
rect 600 -9475 761 -9465
rect 600 -9509 711 -9475
rect 745 -9509 761 -9475
rect 600 -9519 761 -9509
rect 860 -9475 982 -9465
rect 860 -9509 932 -9475
rect 966 -9509 982 -9475
rect 860 -9519 982 -9509
rect 1032 -9475 1102 -9463
rect 1032 -9509 1052 -9475
rect 1086 -9509 1102 -9475
rect 152 -9551 294 -9535
rect 152 -9557 236 -9551
rect 505 -9557 535 -9525
rect 26 -9583 236 -9557
rect 600 -9593 700 -9519
rect 860 -9593 960 -9519
rect 1032 -9522 1102 -9509
rect 1256 -9465 1398 -9449
rect 1256 -9499 1272 -9465
rect 1306 -9499 1398 -9465
rect 1774 -9465 2046 -9443
rect 2602 -9449 2686 -9443
rect 1256 -9515 1398 -9499
rect 1440 -9501 1582 -9485
rect 1032 -9557 1062 -9522
rect 1440 -9535 1532 -9501
rect 1566 -9535 1582 -9501
rect 1774 -9499 1790 -9465
rect 1824 -9499 1893 -9465
rect 1927 -9499 1996 -9465
rect 2030 -9499 2046 -9465
rect 2544 -9465 2686 -9449
rect 3081 -9459 3111 -9391
rect 1774 -9515 2046 -9499
rect 2088 -9501 2352 -9485
rect 1440 -9551 1582 -9535
rect 2088 -9535 2104 -9501
rect 2138 -9535 2203 -9501
rect 2237 -9535 2302 -9501
rect 2336 -9535 2352 -9501
rect 2544 -9499 2560 -9465
rect 2594 -9499 2686 -9465
rect 3077 -9475 3131 -9459
rect 2544 -9515 2686 -9499
rect 2728 -9501 2870 -9485
rect 1440 -9557 1524 -9551
rect 2088 -9557 2352 -9535
rect 2728 -9535 2820 -9501
rect 2854 -9535 2870 -9501
rect 3077 -9509 3087 -9475
rect 3121 -9509 3131 -9475
rect 3077 -9525 3131 -9509
rect 3176 -9465 3276 -9437
rect 3436 -9465 3536 -9437
rect 3608 -9463 3638 -9391
rect 3890 -9443 4100 -9417
rect 4350 -9443 4928 -9417
rect 5178 -9443 5388 -9417
rect 3890 -9449 3974 -9443
rect 3176 -9475 3337 -9465
rect 3176 -9509 3287 -9475
rect 3321 -9509 3337 -9475
rect 3176 -9519 3337 -9509
rect 3436 -9475 3558 -9465
rect 3436 -9509 3508 -9475
rect 3542 -9509 3558 -9475
rect 3436 -9519 3558 -9509
rect 3608 -9475 3678 -9463
rect 3608 -9509 3628 -9475
rect 3662 -9509 3678 -9475
rect 2728 -9551 2870 -9535
rect 2728 -9557 2812 -9551
rect 3081 -9557 3111 -9525
rect 1314 -9583 1524 -9557
rect 1774 -9583 2352 -9557
rect 2602 -9583 2812 -9557
rect 3176 -9593 3276 -9519
rect 3436 -9593 3536 -9519
rect 3608 -9522 3678 -9509
rect 3832 -9465 3974 -9449
rect 3832 -9499 3848 -9465
rect 3882 -9499 3974 -9465
rect 4350 -9465 4622 -9443
rect 5178 -9449 5262 -9443
rect 3832 -9515 3974 -9499
rect 4016 -9501 4158 -9485
rect 3608 -9557 3638 -9522
rect 4016 -9535 4108 -9501
rect 4142 -9535 4158 -9501
rect 4350 -9499 4366 -9465
rect 4400 -9499 4469 -9465
rect 4503 -9499 4572 -9465
rect 4606 -9499 4622 -9465
rect 5120 -9465 5262 -9449
rect 5657 -9459 5687 -9391
rect 4350 -9515 4622 -9499
rect 4664 -9501 4928 -9485
rect 4016 -9551 4158 -9535
rect 4664 -9535 4680 -9501
rect 4714 -9535 4779 -9501
rect 4813 -9535 4878 -9501
rect 4912 -9535 4928 -9501
rect 5120 -9499 5136 -9465
rect 5170 -9499 5262 -9465
rect 5653 -9475 5707 -9459
rect 5120 -9515 5262 -9499
rect 5304 -9501 5446 -9485
rect 4016 -9557 4100 -9551
rect 4664 -9557 4928 -9535
rect 5304 -9535 5396 -9501
rect 5430 -9535 5446 -9501
rect 5653 -9509 5663 -9475
rect 5697 -9509 5707 -9475
rect 5653 -9525 5707 -9509
rect 5752 -9465 5852 -9437
rect 6012 -9465 6112 -9437
rect 6184 -9463 6214 -9391
rect 6466 -9443 6676 -9417
rect 6926 -9443 7504 -9417
rect 7754 -9443 7964 -9417
rect 6466 -9449 6550 -9443
rect 5752 -9475 5913 -9465
rect 5752 -9509 5863 -9475
rect 5897 -9509 5913 -9475
rect 5752 -9519 5913 -9509
rect 6012 -9475 6134 -9465
rect 6012 -9509 6084 -9475
rect 6118 -9509 6134 -9475
rect 6012 -9519 6134 -9509
rect 6184 -9475 6254 -9463
rect 6184 -9509 6204 -9475
rect 6238 -9509 6254 -9475
rect 5304 -9551 5446 -9535
rect 5304 -9557 5388 -9551
rect 5657 -9557 5687 -9525
rect 3890 -9583 4100 -9557
rect 4350 -9583 4928 -9557
rect 5178 -9583 5388 -9557
rect 5752 -9593 5852 -9519
rect 6012 -9593 6112 -9519
rect 6184 -9522 6254 -9509
rect 6408 -9465 6550 -9449
rect 6408 -9499 6424 -9465
rect 6458 -9499 6550 -9465
rect 6926 -9465 7198 -9443
rect 7754 -9449 7838 -9443
rect 6408 -9515 6550 -9499
rect 6592 -9501 6734 -9485
rect 6184 -9557 6214 -9522
rect 6592 -9535 6684 -9501
rect 6718 -9535 6734 -9501
rect 6926 -9499 6942 -9465
rect 6976 -9499 7045 -9465
rect 7079 -9499 7148 -9465
rect 7182 -9499 7198 -9465
rect 7696 -9465 7838 -9449
rect 8233 -9459 8263 -9391
rect 6926 -9515 7198 -9499
rect 7240 -9501 7504 -9485
rect 6592 -9551 6734 -9535
rect 7240 -9535 7256 -9501
rect 7290 -9535 7355 -9501
rect 7389 -9535 7454 -9501
rect 7488 -9535 7504 -9501
rect 7696 -9499 7712 -9465
rect 7746 -9499 7838 -9465
rect 8229 -9475 8283 -9459
rect 7696 -9515 7838 -9499
rect 7880 -9501 8022 -9485
rect 6592 -9557 6676 -9551
rect 7240 -9557 7504 -9535
rect 7880 -9535 7972 -9501
rect 8006 -9535 8022 -9501
rect 8229 -9509 8239 -9475
rect 8273 -9509 8283 -9475
rect 8229 -9525 8283 -9509
rect 8328 -9465 8428 -9437
rect 8588 -9465 8688 -9437
rect 8760 -9463 8790 -9391
rect 9042 -9443 9252 -9417
rect 9502 -9443 10080 -9417
rect 10422 -9443 10632 -9417
rect 9042 -9449 9126 -9443
rect 8328 -9475 8489 -9465
rect 8328 -9509 8439 -9475
rect 8473 -9509 8489 -9475
rect 8328 -9519 8489 -9509
rect 8588 -9475 8710 -9465
rect 8588 -9509 8660 -9475
rect 8694 -9509 8710 -9475
rect 8588 -9519 8710 -9509
rect 8760 -9475 8830 -9463
rect 8760 -9509 8780 -9475
rect 8814 -9509 8830 -9475
rect 7880 -9551 8022 -9535
rect 7880 -9557 7964 -9551
rect 8233 -9557 8263 -9525
rect 6466 -9583 6676 -9557
rect 6926 -9583 7504 -9557
rect 7754 -9583 7964 -9557
rect 8328 -9593 8428 -9519
rect 8588 -9593 8688 -9519
rect 8760 -9522 8830 -9509
rect 8984 -9465 9126 -9449
rect 8984 -9499 9000 -9465
rect 9034 -9499 9126 -9465
rect 9502 -9465 9774 -9443
rect 10422 -9449 10506 -9443
rect 8984 -9515 9126 -9499
rect 9168 -9501 9310 -9485
rect 8760 -9557 8790 -9522
rect 9168 -9535 9260 -9501
rect 9294 -9535 9310 -9501
rect 9502 -9499 9518 -9465
rect 9552 -9499 9621 -9465
rect 9655 -9499 9724 -9465
rect 9758 -9499 9774 -9465
rect 10364 -9465 10506 -9449
rect 10809 -9459 10839 -9391
rect 9502 -9515 9774 -9499
rect 9816 -9501 10080 -9485
rect 9168 -9551 9310 -9535
rect 9816 -9535 9832 -9501
rect 9866 -9535 9931 -9501
rect 9965 -9535 10030 -9501
rect 10064 -9535 10080 -9501
rect 10364 -9499 10380 -9465
rect 10414 -9499 10506 -9465
rect 10805 -9475 10859 -9459
rect 10364 -9515 10506 -9499
rect 10548 -9501 10690 -9485
rect 9168 -9557 9252 -9551
rect 9816 -9557 10080 -9535
rect 10548 -9535 10640 -9501
rect 10674 -9535 10690 -9501
rect 10805 -9509 10815 -9475
rect 10849 -9509 10859 -9475
rect 10805 -9525 10859 -9509
rect 10904 -9465 11004 -9437
rect 11164 -9465 11264 -9437
rect 11336 -9463 11366 -9391
rect 11710 -9443 11920 -9417
rect 13735 -9440 13765 -9391
rect 13821 -9440 13851 -9391
rect 13907 -9440 13937 -9391
rect 13993 -9440 14023 -9391
rect 11710 -9449 11794 -9443
rect 10904 -9475 11065 -9465
rect 10904 -9509 11015 -9475
rect 11049 -9509 11065 -9475
rect 10904 -9519 11065 -9509
rect 11164 -9475 11286 -9465
rect 11164 -9509 11236 -9475
rect 11270 -9509 11286 -9475
rect 11164 -9519 11286 -9509
rect 11336 -9475 11406 -9463
rect 11336 -9509 11356 -9475
rect 11390 -9509 11406 -9475
rect 10548 -9551 10690 -9535
rect 10548 -9557 10632 -9551
rect 10809 -9557 10839 -9525
rect 9042 -9583 9252 -9557
rect 9502 -9583 10080 -9557
rect 10422 -9583 10632 -9557
rect 10904 -9593 11004 -9519
rect 11164 -9593 11264 -9519
rect 11336 -9522 11406 -9509
rect 11652 -9465 11794 -9449
rect 11652 -9499 11668 -9465
rect 11702 -9499 11794 -9465
rect 13676 -9475 14023 -9440
rect 11652 -9515 11794 -9499
rect 11836 -9501 11978 -9485
rect 11336 -9557 11366 -9522
rect 11836 -9535 11928 -9501
rect 11962 -9535 11978 -9501
rect 11836 -9551 11978 -9535
rect 13676 -9509 13692 -9475
rect 13726 -9509 14023 -9475
rect 13676 -9542 14023 -9509
rect 11836 -9557 11920 -9551
rect 13735 -9557 13765 -9542
rect 13821 -9557 13851 -9542
rect 13907 -9557 13937 -9542
rect 13993 -9557 14023 -9542
rect 14079 -9450 14109 -9391
rect 14165 -9450 14195 -9391
rect 14251 -9450 14281 -9391
rect 14337 -9450 14367 -9391
rect 14423 -9450 14453 -9391
rect 14509 -9450 14539 -9391
rect 14595 -9450 14625 -9391
rect 14681 -9450 14711 -9391
rect 14766 -9450 14796 -9391
rect 14852 -9450 14882 -9391
rect 14938 -9450 14968 -9391
rect 15024 -9450 15054 -9391
rect 15110 -9450 15140 -9391
rect 15196 -9450 15226 -9391
rect 15282 -9450 15312 -9391
rect 15368 -9450 15398 -9391
rect 14079 -9475 15398 -9450
rect 14079 -9509 14119 -9475
rect 14153 -9509 14187 -9475
rect 14221 -9509 14255 -9475
rect 14289 -9509 14323 -9475
rect 14357 -9509 14391 -9475
rect 14425 -9509 14459 -9475
rect 14493 -9509 14527 -9475
rect 14561 -9509 14595 -9475
rect 14629 -9509 14663 -9475
rect 14697 -9509 14731 -9475
rect 14765 -9509 14799 -9475
rect 14833 -9509 14867 -9475
rect 14901 -9509 14935 -9475
rect 14969 -9509 15003 -9475
rect 15037 -9509 15071 -9475
rect 15105 -9509 15139 -9475
rect 15173 -9509 15398 -9475
rect 14079 -9525 15398 -9509
rect 15666 -9443 16612 -9417
rect 15666 -9465 16120 -9443
rect 15666 -9499 15686 -9465
rect 15720 -9499 15814 -9465
rect 15848 -9499 15942 -9465
rect 15976 -9499 16070 -9465
rect 16104 -9499 16120 -9465
rect 15666 -9515 16120 -9499
rect 16162 -9501 16612 -9485
rect 14079 -9557 14109 -9525
rect 14165 -9557 14195 -9525
rect 14251 -9557 14281 -9525
rect 14337 -9557 14367 -9525
rect 14423 -9557 14453 -9525
rect 14509 -9557 14539 -9525
rect 14595 -9557 14625 -9525
rect 14681 -9557 14711 -9525
rect 14766 -9557 14796 -9525
rect 14852 -9557 14882 -9525
rect 14938 -9557 14968 -9525
rect 15024 -9557 15054 -9525
rect 15110 -9557 15140 -9525
rect 15196 -9557 15226 -9525
rect 15282 -9557 15312 -9525
rect 15368 -9557 15398 -9525
rect 16162 -9535 16178 -9501
rect 16212 -9535 16306 -9501
rect 16340 -9535 16434 -9501
rect 16468 -9535 16562 -9501
rect 16596 -9535 16612 -9501
rect 16162 -9557 16612 -9535
rect 11710 -9583 11920 -9557
rect 15666 -9583 16612 -9557
rect -2918 -9783 -2340 -9757
rect -1538 -9783 -960 -9757
rect -783 -9783 -753 -9757
rect -688 -9783 -588 -9757
rect -428 -9783 -328 -9757
rect -256 -9783 -226 -9757
rect 26 -9783 236 -9757
rect 505 -9783 535 -9757
rect 600 -9783 700 -9757
rect 860 -9783 960 -9757
rect 1032 -9783 1062 -9757
rect 1314 -9783 1524 -9757
rect 1774 -9783 2352 -9757
rect 2602 -9783 2812 -9757
rect 3081 -9783 3111 -9757
rect 3176 -9783 3276 -9757
rect 3436 -9783 3536 -9757
rect 3608 -9783 3638 -9757
rect 3890 -9783 4100 -9757
rect 4350 -9783 4928 -9757
rect 5178 -9783 5388 -9757
rect 5657 -9783 5687 -9757
rect 5752 -9783 5852 -9757
rect 6012 -9783 6112 -9757
rect 6184 -9783 6214 -9757
rect 6466 -9783 6676 -9757
rect 6926 -9783 7504 -9757
rect 7754 -9783 7964 -9757
rect 8233 -9783 8263 -9757
rect 8328 -9783 8428 -9757
rect 8588 -9783 8688 -9757
rect 8760 -9783 8790 -9757
rect 9042 -9783 9252 -9757
rect 9502 -9783 10080 -9757
rect 10422 -9783 10632 -9757
rect 10809 -9783 10839 -9757
rect 10904 -9783 11004 -9757
rect 11164 -9783 11264 -9757
rect 11336 -9783 11366 -9757
rect 11710 -9783 11920 -9757
rect 13735 -9783 13765 -9757
rect 13821 -9783 13851 -9757
rect 13907 -9783 13937 -9757
rect 13993 -9783 14023 -9757
rect 14079 -9783 14109 -9757
rect 14165 -9783 14195 -9757
rect 14251 -9783 14281 -9757
rect 14337 -9783 14367 -9757
rect 14423 -9783 14453 -9757
rect 14509 -9783 14539 -9757
rect 14595 -9783 14625 -9757
rect 14681 -9783 14711 -9757
rect 14766 -9783 14796 -9757
rect 14852 -9783 14882 -9757
rect 14938 -9783 14968 -9757
rect 15024 -9783 15054 -9757
rect 15110 -9783 15140 -9757
rect 15196 -9783 15226 -9757
rect 15282 -9783 15312 -9757
rect 15368 -9783 15398 -9757
rect 15666 -9783 16612 -9757
rect -2918 -9851 -2340 -9825
rect -1538 -9851 -960 -9825
rect -802 -9851 -224 -9825
rect 26 -9851 236 -9825
rect 488 -9851 518 -9825
rect 590 -9851 690 -9825
rect 850 -9851 950 -9825
rect 1015 -9851 1045 -9825
rect 1314 -9851 1524 -9825
rect 1774 -9851 2352 -9825
rect 2602 -9851 2812 -9825
rect 3064 -9851 3094 -9825
rect 3166 -9851 3266 -9825
rect 3426 -9851 3526 -9825
rect 3591 -9851 3621 -9825
rect 3890 -9851 4100 -9825
rect 4350 -9851 4928 -9825
rect 5178 -9851 5388 -9825
rect 5640 -9851 5670 -9825
rect 5742 -9851 5842 -9825
rect 6002 -9851 6102 -9825
rect 6167 -9851 6197 -9825
rect 6466 -9851 6676 -9825
rect 6926 -9851 7504 -9825
rect 7754 -9851 7964 -9825
rect 8216 -9851 8246 -9825
rect 8318 -9851 8418 -9825
rect 8578 -9851 8678 -9825
rect 8743 -9851 8773 -9825
rect 9042 -9851 9252 -9825
rect 9502 -9851 10080 -9825
rect 10422 -9851 10632 -9825
rect 10792 -9851 10822 -9825
rect 10894 -9851 10994 -9825
rect 11154 -9851 11254 -9825
rect 11319 -9851 11349 -9825
rect 11710 -9851 11920 -9825
rect 12547 -9851 12577 -9825
rect 12633 -9851 12663 -9825
rect 12719 -9851 12749 -9825
rect 12805 -9851 12835 -9825
rect 12891 -9851 12921 -9825
rect 12977 -9851 13007 -9825
rect 13274 -9851 13484 -9825
rect 13735 -9851 13765 -9825
rect 13821 -9851 13851 -9825
rect 13907 -9851 13937 -9825
rect 13993 -9851 14023 -9825
rect 14079 -9851 14109 -9825
rect 14165 -9851 14195 -9825
rect 14251 -9851 14281 -9825
rect 14337 -9851 14367 -9825
rect 14423 -9851 14453 -9825
rect 14509 -9851 14539 -9825
rect 14595 -9851 14625 -9825
rect 14681 -9851 14711 -9825
rect 14766 -9851 14796 -9825
rect 14852 -9851 14882 -9825
rect 14938 -9851 14968 -9825
rect 15024 -9851 15054 -9825
rect 15110 -9851 15140 -9825
rect 15196 -9851 15226 -9825
rect 15282 -9851 15312 -9825
rect 15368 -9851 15398 -9825
rect 15666 -9851 16612 -9825
rect -2918 -10051 -2340 -10025
rect -1538 -10051 -960 -10025
rect -802 -10051 -224 -10025
rect 26 -10051 236 -10025
rect -2918 -10073 -2654 -10051
rect -2918 -10107 -2902 -10073
rect -2868 -10107 -2803 -10073
rect -2769 -10107 -2704 -10073
rect -2670 -10107 -2654 -10073
rect -1538 -10073 -1274 -10051
rect -2918 -10123 -2654 -10107
rect -2612 -10109 -2340 -10093
rect -2612 -10143 -2596 -10109
rect -2562 -10143 -2493 -10109
rect -2459 -10143 -2390 -10109
rect -2356 -10143 -2340 -10109
rect -1538 -10107 -1522 -10073
rect -1488 -10107 -1423 -10073
rect -1389 -10107 -1324 -10073
rect -1290 -10107 -1274 -10073
rect -802 -10073 -538 -10051
rect -1538 -10123 -1274 -10107
rect -1232 -10109 -960 -10093
rect -2612 -10165 -2340 -10143
rect -1232 -10143 -1216 -10109
rect -1182 -10143 -1113 -10109
rect -1079 -10143 -1010 -10109
rect -976 -10143 -960 -10109
rect -802 -10107 -786 -10073
rect -752 -10107 -687 -10073
rect -653 -10107 -588 -10073
rect -554 -10107 -538 -10073
rect 152 -10057 236 -10051
rect 152 -10073 294 -10057
rect -802 -10123 -538 -10107
rect -496 -10109 -224 -10093
rect -1232 -10165 -960 -10143
rect -496 -10143 -480 -10109
rect -446 -10143 -377 -10109
rect -343 -10143 -274 -10109
rect -240 -10143 -224 -10109
rect -496 -10165 -224 -10143
rect -32 -10109 110 -10093
rect -32 -10143 -16 -10109
rect 18 -10143 110 -10109
rect 152 -10107 244 -10073
rect 278 -10107 294 -10073
rect 488 -10086 518 -10051
rect 152 -10123 294 -10107
rect 448 -10099 518 -10086
rect 590 -10089 690 -10015
rect 850 -10089 950 -10015
rect 1314 -10051 1524 -10025
rect 1015 -10083 1045 -10051
rect 1440 -10057 1524 -10051
rect 1774 -10051 2352 -10025
rect 2602 -10051 2812 -10025
rect 1440 -10073 1582 -10057
rect -32 -10159 110 -10143
rect 448 -10133 464 -10099
rect 498 -10133 518 -10099
rect 448 -10145 518 -10133
rect 568 -10099 690 -10089
rect 568 -10133 584 -10099
rect 618 -10133 690 -10099
rect 568 -10143 690 -10133
rect 789 -10099 950 -10089
rect 789 -10133 805 -10099
rect 839 -10133 950 -10099
rect 789 -10143 950 -10133
rect -2918 -10191 -2340 -10165
rect -1538 -10191 -960 -10165
rect -802 -10191 -224 -10165
rect 26 -10165 110 -10159
rect 26 -10191 236 -10165
rect 488 -10217 518 -10145
rect 590 -10171 690 -10143
rect 850 -10171 950 -10143
rect 995 -10099 1049 -10083
rect 995 -10133 1005 -10099
rect 1039 -10133 1049 -10099
rect 995 -10149 1049 -10133
rect 1256 -10109 1398 -10093
rect 1256 -10143 1272 -10109
rect 1306 -10143 1398 -10109
rect 1440 -10107 1532 -10073
rect 1566 -10107 1582 -10073
rect 1440 -10123 1582 -10107
rect 1774 -10073 2038 -10051
rect 1774 -10107 1790 -10073
rect 1824 -10107 1889 -10073
rect 1923 -10107 1988 -10073
rect 2022 -10107 2038 -10073
rect 2728 -10057 2812 -10051
rect 2728 -10073 2870 -10057
rect 1774 -10123 2038 -10107
rect 2080 -10109 2352 -10093
rect 1015 -10217 1045 -10149
rect 1256 -10159 1398 -10143
rect 1314 -10165 1398 -10159
rect 2080 -10143 2096 -10109
rect 2130 -10143 2199 -10109
rect 2233 -10143 2302 -10109
rect 2336 -10143 2352 -10109
rect 2080 -10165 2352 -10143
rect 2544 -10109 2686 -10093
rect 2544 -10143 2560 -10109
rect 2594 -10143 2686 -10109
rect 2728 -10107 2820 -10073
rect 2854 -10107 2870 -10073
rect 3064 -10086 3094 -10051
rect 2728 -10123 2870 -10107
rect 3024 -10099 3094 -10086
rect 3166 -10089 3266 -10015
rect 3426 -10089 3526 -10015
rect 3890 -10051 4100 -10025
rect 3591 -10083 3621 -10051
rect 4016 -10057 4100 -10051
rect 4350 -10051 4928 -10025
rect 5178 -10051 5388 -10025
rect 4016 -10073 4158 -10057
rect 2544 -10159 2686 -10143
rect 3024 -10133 3040 -10099
rect 3074 -10133 3094 -10099
rect 3024 -10145 3094 -10133
rect 3144 -10099 3266 -10089
rect 3144 -10133 3160 -10099
rect 3194 -10133 3266 -10099
rect 3144 -10143 3266 -10133
rect 3365 -10099 3526 -10089
rect 3365 -10133 3381 -10099
rect 3415 -10133 3526 -10099
rect 3365 -10143 3526 -10133
rect 1314 -10191 1524 -10165
rect 1774 -10191 2352 -10165
rect 2602 -10165 2686 -10159
rect 2602 -10191 2812 -10165
rect 3064 -10217 3094 -10145
rect 3166 -10171 3266 -10143
rect 3426 -10171 3526 -10143
rect 3571 -10099 3625 -10083
rect 3571 -10133 3581 -10099
rect 3615 -10133 3625 -10099
rect 3571 -10149 3625 -10133
rect 3832 -10109 3974 -10093
rect 3832 -10143 3848 -10109
rect 3882 -10143 3974 -10109
rect 4016 -10107 4108 -10073
rect 4142 -10107 4158 -10073
rect 4016 -10123 4158 -10107
rect 4350 -10073 4614 -10051
rect 4350 -10107 4366 -10073
rect 4400 -10107 4465 -10073
rect 4499 -10107 4564 -10073
rect 4598 -10107 4614 -10073
rect 5304 -10057 5388 -10051
rect 5304 -10073 5446 -10057
rect 4350 -10123 4614 -10107
rect 4656 -10109 4928 -10093
rect 3591 -10217 3621 -10149
rect 3832 -10159 3974 -10143
rect 3890 -10165 3974 -10159
rect 4656 -10143 4672 -10109
rect 4706 -10143 4775 -10109
rect 4809 -10143 4878 -10109
rect 4912 -10143 4928 -10109
rect 4656 -10165 4928 -10143
rect 5120 -10109 5262 -10093
rect 5120 -10143 5136 -10109
rect 5170 -10143 5262 -10109
rect 5304 -10107 5396 -10073
rect 5430 -10107 5446 -10073
rect 5640 -10086 5670 -10051
rect 5304 -10123 5446 -10107
rect 5600 -10099 5670 -10086
rect 5742 -10089 5842 -10015
rect 6002 -10089 6102 -10015
rect 6466 -10051 6676 -10025
rect 6167 -10083 6197 -10051
rect 6592 -10057 6676 -10051
rect 6926 -10051 7504 -10025
rect 7754 -10051 7964 -10025
rect 6592 -10073 6734 -10057
rect 5120 -10159 5262 -10143
rect 5600 -10133 5616 -10099
rect 5650 -10133 5670 -10099
rect 5600 -10145 5670 -10133
rect 5720 -10099 5842 -10089
rect 5720 -10133 5736 -10099
rect 5770 -10133 5842 -10099
rect 5720 -10143 5842 -10133
rect 5941 -10099 6102 -10089
rect 5941 -10133 5957 -10099
rect 5991 -10133 6102 -10099
rect 5941 -10143 6102 -10133
rect 3890 -10191 4100 -10165
rect 4350 -10191 4928 -10165
rect 5178 -10165 5262 -10159
rect 5178 -10191 5388 -10165
rect 5640 -10217 5670 -10145
rect 5742 -10171 5842 -10143
rect 6002 -10171 6102 -10143
rect 6147 -10099 6201 -10083
rect 6147 -10133 6157 -10099
rect 6191 -10133 6201 -10099
rect 6147 -10149 6201 -10133
rect 6408 -10109 6550 -10093
rect 6408 -10143 6424 -10109
rect 6458 -10143 6550 -10109
rect 6592 -10107 6684 -10073
rect 6718 -10107 6734 -10073
rect 6592 -10123 6734 -10107
rect 6926 -10073 7190 -10051
rect 6926 -10107 6942 -10073
rect 6976 -10107 7041 -10073
rect 7075 -10107 7140 -10073
rect 7174 -10107 7190 -10073
rect 7880 -10057 7964 -10051
rect 7880 -10073 8022 -10057
rect 6926 -10123 7190 -10107
rect 7232 -10109 7504 -10093
rect 6167 -10217 6197 -10149
rect 6408 -10159 6550 -10143
rect 6466 -10165 6550 -10159
rect 7232 -10143 7248 -10109
rect 7282 -10143 7351 -10109
rect 7385 -10143 7454 -10109
rect 7488 -10143 7504 -10109
rect 7232 -10165 7504 -10143
rect 7696 -10109 7838 -10093
rect 7696 -10143 7712 -10109
rect 7746 -10143 7838 -10109
rect 7880 -10107 7972 -10073
rect 8006 -10107 8022 -10073
rect 8216 -10086 8246 -10051
rect 7880 -10123 8022 -10107
rect 8176 -10099 8246 -10086
rect 8318 -10089 8418 -10015
rect 8578 -10089 8678 -10015
rect 9042 -10051 9252 -10025
rect 8743 -10083 8773 -10051
rect 9168 -10057 9252 -10051
rect 9502 -10051 10080 -10025
rect 10422 -10051 10632 -10025
rect 9168 -10073 9310 -10057
rect 7696 -10159 7838 -10143
rect 8176 -10133 8192 -10099
rect 8226 -10133 8246 -10099
rect 8176 -10145 8246 -10133
rect 8296 -10099 8418 -10089
rect 8296 -10133 8312 -10099
rect 8346 -10133 8418 -10099
rect 8296 -10143 8418 -10133
rect 8517 -10099 8678 -10089
rect 8517 -10133 8533 -10099
rect 8567 -10133 8678 -10099
rect 8517 -10143 8678 -10133
rect 6466 -10191 6676 -10165
rect 6926 -10191 7504 -10165
rect 7754 -10165 7838 -10159
rect 7754 -10191 7964 -10165
rect 8216 -10217 8246 -10145
rect 8318 -10171 8418 -10143
rect 8578 -10171 8678 -10143
rect 8723 -10099 8777 -10083
rect 8723 -10133 8733 -10099
rect 8767 -10133 8777 -10099
rect 8723 -10149 8777 -10133
rect 8984 -10109 9126 -10093
rect 8984 -10143 9000 -10109
rect 9034 -10143 9126 -10109
rect 9168 -10107 9260 -10073
rect 9294 -10107 9310 -10073
rect 9168 -10123 9310 -10107
rect 9502 -10073 9766 -10051
rect 9502 -10107 9518 -10073
rect 9552 -10107 9617 -10073
rect 9651 -10107 9716 -10073
rect 9750 -10107 9766 -10073
rect 10548 -10057 10632 -10051
rect 10548 -10073 10690 -10057
rect 9502 -10123 9766 -10107
rect 9808 -10109 10080 -10093
rect 8743 -10217 8773 -10149
rect 8984 -10159 9126 -10143
rect 9042 -10165 9126 -10159
rect 9808 -10143 9824 -10109
rect 9858 -10143 9927 -10109
rect 9961 -10143 10030 -10109
rect 10064 -10143 10080 -10109
rect 9808 -10165 10080 -10143
rect 10364 -10109 10506 -10093
rect 10364 -10143 10380 -10109
rect 10414 -10143 10506 -10109
rect 10548 -10107 10640 -10073
rect 10674 -10107 10690 -10073
rect 10792 -10086 10822 -10051
rect 10548 -10123 10690 -10107
rect 10752 -10099 10822 -10086
rect 10894 -10089 10994 -10015
rect 11154 -10089 11254 -10015
rect 11710 -10051 11920 -10025
rect 13274 -10051 13484 -10025
rect 15666 -10051 16612 -10025
rect 11319 -10083 11349 -10051
rect 11836 -10057 11920 -10051
rect 11836 -10073 11978 -10057
rect 10364 -10159 10506 -10143
rect 10752 -10133 10768 -10099
rect 10802 -10133 10822 -10099
rect 10752 -10145 10822 -10133
rect 10872 -10099 10994 -10089
rect 10872 -10133 10888 -10099
rect 10922 -10133 10994 -10099
rect 10872 -10143 10994 -10133
rect 11093 -10099 11254 -10089
rect 11093 -10133 11109 -10099
rect 11143 -10133 11254 -10099
rect 11093 -10143 11254 -10133
rect 9042 -10191 9252 -10165
rect 9502 -10191 10080 -10165
rect 10422 -10165 10506 -10159
rect 10422 -10191 10632 -10165
rect 10792 -10217 10822 -10145
rect 10894 -10171 10994 -10143
rect 11154 -10171 11254 -10143
rect 11299 -10099 11353 -10083
rect 11299 -10133 11309 -10099
rect 11343 -10133 11353 -10099
rect 11299 -10149 11353 -10133
rect 11652 -10109 11794 -10093
rect 11652 -10143 11668 -10109
rect 11702 -10143 11794 -10109
rect 11836 -10107 11928 -10073
rect 11962 -10107 11978 -10073
rect 11836 -10123 11978 -10107
rect 12547 -10089 12577 -10051
rect 12633 -10089 12663 -10051
rect 12719 -10089 12749 -10051
rect 12805 -10089 12835 -10051
rect 12891 -10089 12921 -10051
rect 12977 -10089 13007 -10051
rect 13274 -10057 13358 -10051
rect 12547 -10099 13007 -10089
rect 12547 -10133 12574 -10099
rect 12608 -10133 12642 -10099
rect 12676 -10133 12710 -10099
rect 12744 -10133 12778 -10099
rect 12812 -10133 12846 -10099
rect 12880 -10133 12914 -10099
rect 12948 -10133 13007 -10099
rect 13216 -10073 13358 -10057
rect 13735 -10066 13765 -10051
rect 13821 -10066 13851 -10051
rect 13907 -10066 13937 -10051
rect 13993 -10066 14023 -10051
rect 13216 -10107 13232 -10073
rect 13266 -10107 13358 -10073
rect 13216 -10123 13358 -10107
rect 13400 -10109 13542 -10093
rect 12547 -10143 13007 -10133
rect 13400 -10143 13492 -10109
rect 13526 -10143 13542 -10109
rect 11319 -10217 11349 -10149
rect 11652 -10159 11794 -10143
rect 11710 -10165 11794 -10159
rect 11710 -10191 11920 -10165
rect 12633 -10217 12663 -10143
rect 12719 -10217 12749 -10143
rect 12805 -10217 12835 -10143
rect 12891 -10217 12921 -10143
rect 13400 -10159 13542 -10143
rect 13676 -10099 14023 -10066
rect 13676 -10133 13692 -10099
rect 13726 -10133 14023 -10099
rect 13400 -10165 13484 -10159
rect 13274 -10191 13484 -10165
rect 13676 -10168 14023 -10133
rect 13735 -10217 13765 -10168
rect 13821 -10217 13851 -10168
rect 13907 -10217 13937 -10168
rect 13993 -10217 14023 -10168
rect 14079 -10083 14109 -10051
rect 14165 -10083 14195 -10051
rect 14251 -10083 14281 -10051
rect 14337 -10083 14367 -10051
rect 14423 -10083 14453 -10051
rect 14509 -10083 14539 -10051
rect 14595 -10083 14625 -10051
rect 14681 -10083 14711 -10051
rect 14766 -10083 14796 -10051
rect 14852 -10083 14882 -10051
rect 14938 -10083 14968 -10051
rect 15024 -10083 15054 -10051
rect 15110 -10083 15140 -10051
rect 15196 -10083 15226 -10051
rect 15282 -10083 15312 -10051
rect 15368 -10083 15398 -10051
rect 14079 -10099 15398 -10083
rect 14079 -10133 14119 -10099
rect 14153 -10133 14187 -10099
rect 14221 -10133 14255 -10099
rect 14289 -10133 14323 -10099
rect 14357 -10133 14391 -10099
rect 14425 -10133 14459 -10099
rect 14493 -10133 14527 -10099
rect 14561 -10133 14595 -10099
rect 14629 -10133 14663 -10099
rect 14697 -10133 14731 -10099
rect 14765 -10133 14799 -10099
rect 14833 -10133 14867 -10099
rect 14901 -10133 14935 -10099
rect 14969 -10133 15003 -10099
rect 15037 -10133 15071 -10099
rect 15105 -10133 15139 -10099
rect 15173 -10133 15398 -10099
rect 15666 -10073 16116 -10051
rect 15666 -10107 15682 -10073
rect 15716 -10107 15810 -10073
rect 15844 -10107 15938 -10073
rect 15972 -10107 16066 -10073
rect 16100 -10107 16116 -10073
rect 15666 -10123 16116 -10107
rect 16158 -10109 16612 -10093
rect 14079 -10158 15398 -10133
rect 14079 -10217 14109 -10158
rect 14165 -10217 14195 -10158
rect 14251 -10217 14281 -10158
rect 14337 -10217 14367 -10158
rect 14423 -10217 14453 -10158
rect 14509 -10217 14539 -10158
rect 14595 -10217 14625 -10158
rect 14681 -10217 14711 -10158
rect 14766 -10217 14796 -10158
rect 14852 -10217 14882 -10158
rect 14938 -10217 14968 -10158
rect 15024 -10217 15054 -10158
rect 15110 -10217 15140 -10158
rect 15196 -10217 15226 -10158
rect 15282 -10217 15312 -10158
rect 15368 -10217 15398 -10158
rect 16158 -10143 16174 -10109
rect 16208 -10143 16302 -10109
rect 16336 -10143 16430 -10109
rect 16464 -10143 16558 -10109
rect 16592 -10143 16612 -10109
rect 16158 -10165 16612 -10143
rect 15666 -10191 16612 -10165
rect -2918 -10327 -2340 -10301
rect -1538 -10327 -960 -10301
rect -802 -10327 -224 -10301
rect 26 -10327 236 -10301
rect 488 -10327 518 -10301
rect 590 -10327 690 -10301
rect 850 -10327 950 -10301
rect 1015 -10327 1045 -10301
rect 1314 -10327 1524 -10301
rect 1774 -10327 2352 -10301
rect 2602 -10327 2812 -10301
rect 3064 -10327 3094 -10301
rect 3166 -10327 3266 -10301
rect 3426 -10327 3526 -10301
rect 3591 -10327 3621 -10301
rect 3890 -10327 4100 -10301
rect 4350 -10327 4928 -10301
rect 5178 -10327 5388 -10301
rect 5640 -10327 5670 -10301
rect 5742 -10327 5842 -10301
rect 6002 -10327 6102 -10301
rect 6167 -10327 6197 -10301
rect 6466 -10327 6676 -10301
rect 6926 -10327 7504 -10301
rect 7754 -10327 7964 -10301
rect 8216 -10327 8246 -10301
rect 8318 -10327 8418 -10301
rect 8578 -10327 8678 -10301
rect 8743 -10327 8773 -10301
rect 9042 -10327 9252 -10301
rect 9502 -10327 10080 -10301
rect 10422 -10327 10632 -10301
rect 10792 -10327 10822 -10301
rect 10894 -10327 10994 -10301
rect 11154 -10327 11254 -10301
rect 11319 -10327 11349 -10301
rect 11710 -10327 11920 -10301
rect 12633 -10327 12663 -10301
rect 12719 -10327 12749 -10301
rect 12805 -10327 12835 -10301
rect 12891 -10327 12921 -10301
rect 13274 -10327 13484 -10301
rect 13735 -10327 13765 -10301
rect 13821 -10327 13851 -10301
rect 13907 -10327 13937 -10301
rect 13993 -10327 14023 -10301
rect 14079 -10327 14109 -10301
rect 14165 -10327 14195 -10301
rect 14251 -10327 14281 -10301
rect 14337 -10327 14367 -10301
rect 14423 -10327 14453 -10301
rect 14509 -10327 14539 -10301
rect 14595 -10327 14625 -10301
rect 14681 -10327 14711 -10301
rect 14766 -10327 14796 -10301
rect 14852 -10327 14882 -10301
rect 14938 -10327 14968 -10301
rect 15024 -10327 15054 -10301
rect 15110 -10327 15140 -10301
rect 15196 -10327 15226 -10301
rect 15282 -10327 15312 -10301
rect 15368 -10327 15398 -10301
rect 15666 -10327 16612 -10301
rect -2918 -10395 -2340 -10369
rect -1823 -10395 -1793 -10369
rect -1538 -10395 -960 -10369
rect -802 -10395 -224 -10369
rect 26 -10395 236 -10369
rect 505 -10395 535 -10369
rect 600 -10395 700 -10369
rect 860 -10395 960 -10369
rect 1032 -10395 1062 -10369
rect 1314 -10395 1524 -10369
rect 1774 -10395 2352 -10369
rect 2602 -10395 2812 -10369
rect 3081 -10395 3111 -10369
rect 3176 -10395 3276 -10369
rect 3436 -10395 3536 -10369
rect 3608 -10395 3638 -10369
rect 3890 -10395 4100 -10369
rect 4350 -10395 4928 -10369
rect 5178 -10395 5388 -10369
rect 5657 -10395 5687 -10369
rect 5752 -10395 5852 -10369
rect 6012 -10395 6112 -10369
rect 6184 -10395 6214 -10369
rect 6466 -10395 6676 -10369
rect 6926 -10395 7504 -10369
rect 7754 -10395 7964 -10369
rect 8233 -10395 8263 -10369
rect 8328 -10395 8428 -10369
rect 8588 -10395 8688 -10369
rect 8760 -10395 8790 -10369
rect 9042 -10395 9252 -10369
rect 9502 -10395 10080 -10369
rect 10422 -10395 10632 -10369
rect 10809 -10395 10839 -10369
rect 10904 -10395 11004 -10369
rect 11164 -10395 11264 -10369
rect 11336 -10395 11366 -10369
rect 11710 -10395 11920 -10369
rect 13642 -10395 14588 -10369
rect 14838 -10395 15784 -10369
rect 16034 -10395 16612 -10369
rect -2918 -10531 -2340 -10505
rect -2918 -10553 -2646 -10531
rect -1823 -10543 -1793 -10479
rect -1907 -10547 -1793 -10543
rect -2918 -10587 -2902 -10553
rect -2868 -10587 -2799 -10553
rect -2765 -10587 -2696 -10553
rect -2662 -10587 -2646 -10553
rect -1964 -10563 -1793 -10547
rect -2918 -10603 -2646 -10587
rect -2604 -10589 -2340 -10573
rect -2604 -10623 -2588 -10589
rect -2554 -10623 -2489 -10589
rect -2455 -10623 -2390 -10589
rect -2356 -10623 -2340 -10589
rect -1964 -10597 -1954 -10563
rect -1920 -10587 -1793 -10563
rect -1538 -10531 -960 -10505
rect -802 -10531 -224 -10505
rect 26 -10531 236 -10505
rect -1538 -10553 -1266 -10531
rect -1538 -10587 -1522 -10553
rect -1488 -10587 -1419 -10553
rect -1385 -10587 -1316 -10553
rect -1282 -10587 -1266 -10553
rect -802 -10553 -530 -10531
rect 26 -10537 110 -10531
rect -1920 -10597 -1792 -10587
rect -1964 -10613 -1792 -10597
rect -1538 -10603 -1266 -10587
rect -1224 -10589 -960 -10573
rect -2604 -10645 -2340 -10623
rect -2918 -10671 -2340 -10645
rect -1906 -10617 -1792 -10613
rect -1906 -10677 -1876 -10617
rect -1822 -10677 -1792 -10617
rect -1224 -10623 -1208 -10589
rect -1174 -10623 -1109 -10589
rect -1075 -10623 -1010 -10589
rect -976 -10623 -960 -10589
rect -802 -10587 -786 -10553
rect -752 -10587 -683 -10553
rect -649 -10587 -580 -10553
rect -546 -10587 -530 -10553
rect -32 -10553 110 -10537
rect 505 -10547 535 -10479
rect -802 -10603 -530 -10587
rect -488 -10589 -224 -10573
rect -1224 -10645 -960 -10623
rect -488 -10623 -472 -10589
rect -438 -10623 -373 -10589
rect -339 -10623 -274 -10589
rect -240 -10623 -224 -10589
rect -32 -10587 -16 -10553
rect 18 -10587 110 -10553
rect 501 -10563 555 -10547
rect -32 -10603 110 -10587
rect 152 -10589 294 -10573
rect -488 -10645 -224 -10623
rect 152 -10623 244 -10589
rect 278 -10623 294 -10589
rect 501 -10597 511 -10563
rect 545 -10597 555 -10563
rect 501 -10613 555 -10597
rect 600 -10553 700 -10525
rect 860 -10553 960 -10525
rect 1032 -10551 1062 -10479
rect 1314 -10531 1524 -10505
rect 1774 -10531 2352 -10505
rect 2602 -10531 2812 -10505
rect 1314 -10537 1398 -10531
rect 600 -10563 761 -10553
rect 600 -10597 711 -10563
rect 745 -10597 761 -10563
rect 600 -10607 761 -10597
rect 860 -10563 982 -10553
rect 860 -10597 932 -10563
rect 966 -10597 982 -10563
rect 860 -10607 982 -10597
rect 1032 -10563 1102 -10551
rect 1032 -10597 1052 -10563
rect 1086 -10597 1102 -10563
rect 152 -10639 294 -10623
rect 152 -10645 236 -10639
rect 505 -10645 535 -10613
rect -1538 -10671 -960 -10645
rect -802 -10671 -224 -10645
rect 26 -10671 236 -10645
rect 600 -10681 700 -10607
rect 860 -10681 960 -10607
rect 1032 -10610 1102 -10597
rect 1256 -10553 1398 -10537
rect 1256 -10587 1272 -10553
rect 1306 -10587 1398 -10553
rect 1774 -10553 2046 -10531
rect 2602 -10537 2686 -10531
rect 1256 -10603 1398 -10587
rect 1440 -10589 1582 -10573
rect 1032 -10645 1062 -10610
rect 1440 -10623 1532 -10589
rect 1566 -10623 1582 -10589
rect 1774 -10587 1790 -10553
rect 1824 -10587 1893 -10553
rect 1927 -10587 1996 -10553
rect 2030 -10587 2046 -10553
rect 2544 -10553 2686 -10537
rect 3081 -10547 3111 -10479
rect 1774 -10603 2046 -10587
rect 2088 -10589 2352 -10573
rect 1440 -10639 1582 -10623
rect 2088 -10623 2104 -10589
rect 2138 -10623 2203 -10589
rect 2237 -10623 2302 -10589
rect 2336 -10623 2352 -10589
rect 2544 -10587 2560 -10553
rect 2594 -10587 2686 -10553
rect 3077 -10563 3131 -10547
rect 2544 -10603 2686 -10587
rect 2728 -10589 2870 -10573
rect 1440 -10645 1524 -10639
rect 2088 -10645 2352 -10623
rect 2728 -10623 2820 -10589
rect 2854 -10623 2870 -10589
rect 3077 -10597 3087 -10563
rect 3121 -10597 3131 -10563
rect 3077 -10613 3131 -10597
rect 3176 -10553 3276 -10525
rect 3436 -10553 3536 -10525
rect 3608 -10551 3638 -10479
rect 3890 -10531 4100 -10505
rect 4350 -10531 4928 -10505
rect 5178 -10531 5388 -10505
rect 3890 -10537 3974 -10531
rect 3176 -10563 3337 -10553
rect 3176 -10597 3287 -10563
rect 3321 -10597 3337 -10563
rect 3176 -10607 3337 -10597
rect 3436 -10563 3558 -10553
rect 3436 -10597 3508 -10563
rect 3542 -10597 3558 -10563
rect 3436 -10607 3558 -10597
rect 3608 -10563 3678 -10551
rect 3608 -10597 3628 -10563
rect 3662 -10597 3678 -10563
rect 2728 -10639 2870 -10623
rect 2728 -10645 2812 -10639
rect 3081 -10645 3111 -10613
rect 1314 -10671 1524 -10645
rect 1774 -10671 2352 -10645
rect 2602 -10671 2812 -10645
rect 3176 -10681 3276 -10607
rect 3436 -10681 3536 -10607
rect 3608 -10610 3678 -10597
rect 3832 -10553 3974 -10537
rect 3832 -10587 3848 -10553
rect 3882 -10587 3974 -10553
rect 4350 -10553 4622 -10531
rect 5178 -10537 5262 -10531
rect 3832 -10603 3974 -10587
rect 4016 -10589 4158 -10573
rect 3608 -10645 3638 -10610
rect 4016 -10623 4108 -10589
rect 4142 -10623 4158 -10589
rect 4350 -10587 4366 -10553
rect 4400 -10587 4469 -10553
rect 4503 -10587 4572 -10553
rect 4606 -10587 4622 -10553
rect 5120 -10553 5262 -10537
rect 5657 -10547 5687 -10479
rect 4350 -10603 4622 -10587
rect 4664 -10589 4928 -10573
rect 4016 -10639 4158 -10623
rect 4664 -10623 4680 -10589
rect 4714 -10623 4779 -10589
rect 4813 -10623 4878 -10589
rect 4912 -10623 4928 -10589
rect 5120 -10587 5136 -10553
rect 5170 -10587 5262 -10553
rect 5653 -10563 5707 -10547
rect 5120 -10603 5262 -10587
rect 5304 -10589 5446 -10573
rect 4016 -10645 4100 -10639
rect 4664 -10645 4928 -10623
rect 5304 -10623 5396 -10589
rect 5430 -10623 5446 -10589
rect 5653 -10597 5663 -10563
rect 5697 -10597 5707 -10563
rect 5653 -10613 5707 -10597
rect 5752 -10553 5852 -10525
rect 6012 -10553 6112 -10525
rect 6184 -10551 6214 -10479
rect 6466 -10531 6676 -10505
rect 6926 -10531 7504 -10505
rect 7754 -10531 7964 -10505
rect 6466 -10537 6550 -10531
rect 5752 -10563 5913 -10553
rect 5752 -10597 5863 -10563
rect 5897 -10597 5913 -10563
rect 5752 -10607 5913 -10597
rect 6012 -10563 6134 -10553
rect 6012 -10597 6084 -10563
rect 6118 -10597 6134 -10563
rect 6012 -10607 6134 -10597
rect 6184 -10563 6254 -10551
rect 6184 -10597 6204 -10563
rect 6238 -10597 6254 -10563
rect 5304 -10639 5446 -10623
rect 5304 -10645 5388 -10639
rect 5657 -10645 5687 -10613
rect 3890 -10671 4100 -10645
rect 4350 -10671 4928 -10645
rect 5178 -10671 5388 -10645
rect 5752 -10681 5852 -10607
rect 6012 -10681 6112 -10607
rect 6184 -10610 6254 -10597
rect 6408 -10553 6550 -10537
rect 6408 -10587 6424 -10553
rect 6458 -10587 6550 -10553
rect 6926 -10553 7198 -10531
rect 7754 -10537 7838 -10531
rect 6408 -10603 6550 -10587
rect 6592 -10589 6734 -10573
rect 6184 -10645 6214 -10610
rect 6592 -10623 6684 -10589
rect 6718 -10623 6734 -10589
rect 6926 -10587 6942 -10553
rect 6976 -10587 7045 -10553
rect 7079 -10587 7148 -10553
rect 7182 -10587 7198 -10553
rect 7696 -10553 7838 -10537
rect 8233 -10547 8263 -10479
rect 6926 -10603 7198 -10587
rect 7240 -10589 7504 -10573
rect 6592 -10639 6734 -10623
rect 7240 -10623 7256 -10589
rect 7290 -10623 7355 -10589
rect 7389 -10623 7454 -10589
rect 7488 -10623 7504 -10589
rect 7696 -10587 7712 -10553
rect 7746 -10587 7838 -10553
rect 8229 -10563 8283 -10547
rect 7696 -10603 7838 -10587
rect 7880 -10589 8022 -10573
rect 6592 -10645 6676 -10639
rect 7240 -10645 7504 -10623
rect 7880 -10623 7972 -10589
rect 8006 -10623 8022 -10589
rect 8229 -10597 8239 -10563
rect 8273 -10597 8283 -10563
rect 8229 -10613 8283 -10597
rect 8328 -10553 8428 -10525
rect 8588 -10553 8688 -10525
rect 8760 -10551 8790 -10479
rect 9042 -10531 9252 -10505
rect 9502 -10531 10080 -10505
rect 10422 -10531 10632 -10505
rect 9042 -10537 9126 -10531
rect 8328 -10563 8489 -10553
rect 8328 -10597 8439 -10563
rect 8473 -10597 8489 -10563
rect 8328 -10607 8489 -10597
rect 8588 -10563 8710 -10553
rect 8588 -10597 8660 -10563
rect 8694 -10597 8710 -10563
rect 8588 -10607 8710 -10597
rect 8760 -10563 8830 -10551
rect 8760 -10597 8780 -10563
rect 8814 -10597 8830 -10563
rect 7880 -10639 8022 -10623
rect 7880 -10645 7964 -10639
rect 8233 -10645 8263 -10613
rect 6466 -10671 6676 -10645
rect 6926 -10671 7504 -10645
rect 7754 -10671 7964 -10645
rect 8328 -10681 8428 -10607
rect 8588 -10681 8688 -10607
rect 8760 -10610 8830 -10597
rect 8984 -10553 9126 -10537
rect 8984 -10587 9000 -10553
rect 9034 -10587 9126 -10553
rect 9502 -10553 9774 -10531
rect 10422 -10537 10506 -10531
rect 8984 -10603 9126 -10587
rect 9168 -10589 9310 -10573
rect 8760 -10645 8790 -10610
rect 9168 -10623 9260 -10589
rect 9294 -10623 9310 -10589
rect 9502 -10587 9518 -10553
rect 9552 -10587 9621 -10553
rect 9655 -10587 9724 -10553
rect 9758 -10587 9774 -10553
rect 10364 -10553 10506 -10537
rect 10809 -10547 10839 -10479
rect 9502 -10603 9774 -10587
rect 9816 -10589 10080 -10573
rect 9168 -10639 9310 -10623
rect 9816 -10623 9832 -10589
rect 9866 -10623 9931 -10589
rect 9965 -10623 10030 -10589
rect 10064 -10623 10080 -10589
rect 10364 -10587 10380 -10553
rect 10414 -10587 10506 -10553
rect 10805 -10563 10859 -10547
rect 10364 -10603 10506 -10587
rect 10548 -10589 10690 -10573
rect 9168 -10645 9252 -10639
rect 9816 -10645 10080 -10623
rect 10548 -10623 10640 -10589
rect 10674 -10623 10690 -10589
rect 10805 -10597 10815 -10563
rect 10849 -10597 10859 -10563
rect 10805 -10613 10859 -10597
rect 10904 -10553 11004 -10525
rect 11164 -10553 11264 -10525
rect 11336 -10551 11366 -10479
rect 11710 -10531 11920 -10505
rect 13642 -10531 14588 -10505
rect 14838 -10531 15784 -10505
rect 16034 -10531 16612 -10505
rect 11710 -10537 11794 -10531
rect 10904 -10563 11065 -10553
rect 10904 -10597 11015 -10563
rect 11049 -10597 11065 -10563
rect 10904 -10607 11065 -10597
rect 11164 -10563 11286 -10553
rect 11164 -10597 11236 -10563
rect 11270 -10597 11286 -10563
rect 11164 -10607 11286 -10597
rect 11336 -10563 11406 -10551
rect 11336 -10597 11356 -10563
rect 11390 -10597 11406 -10563
rect 10548 -10639 10690 -10623
rect 10548 -10645 10632 -10639
rect 10809 -10645 10839 -10613
rect 9042 -10671 9252 -10645
rect 9502 -10671 10080 -10645
rect 10422 -10671 10632 -10645
rect 10904 -10681 11004 -10607
rect 11164 -10681 11264 -10607
rect 11336 -10610 11406 -10597
rect 11652 -10553 11794 -10537
rect 11652 -10587 11668 -10553
rect 11702 -10587 11794 -10553
rect 13642 -10553 14096 -10531
rect 11652 -10603 11794 -10587
rect 11836 -10589 11978 -10573
rect 11336 -10645 11366 -10610
rect 11836 -10623 11928 -10589
rect 11962 -10623 11978 -10589
rect 13642 -10587 13662 -10553
rect 13696 -10587 13790 -10553
rect 13824 -10587 13918 -10553
rect 13952 -10587 14046 -10553
rect 14080 -10587 14096 -10553
rect 14838 -10553 15292 -10531
rect 13642 -10603 14096 -10587
rect 14138 -10589 14588 -10573
rect 11836 -10639 11978 -10623
rect 14138 -10623 14154 -10589
rect 14188 -10623 14282 -10589
rect 14316 -10623 14410 -10589
rect 14444 -10623 14538 -10589
rect 14572 -10623 14588 -10589
rect 14838 -10587 14858 -10553
rect 14892 -10587 14986 -10553
rect 15020 -10587 15114 -10553
rect 15148 -10587 15242 -10553
rect 15276 -10587 15292 -10553
rect 16034 -10553 16306 -10531
rect 14838 -10603 15292 -10587
rect 15334 -10589 15784 -10573
rect 11836 -10645 11920 -10639
rect 14138 -10645 14588 -10623
rect 15334 -10623 15350 -10589
rect 15384 -10623 15478 -10589
rect 15512 -10623 15606 -10589
rect 15640 -10623 15734 -10589
rect 15768 -10623 15784 -10589
rect 16034 -10587 16050 -10553
rect 16084 -10587 16153 -10553
rect 16187 -10587 16256 -10553
rect 16290 -10587 16306 -10553
rect 16034 -10603 16306 -10587
rect 16348 -10589 16612 -10573
rect 15334 -10645 15784 -10623
rect 16348 -10623 16364 -10589
rect 16398 -10623 16463 -10589
rect 16497 -10623 16562 -10589
rect 16596 -10623 16612 -10589
rect 16348 -10645 16612 -10623
rect 11710 -10671 11920 -10645
rect 13642 -10671 14588 -10645
rect 14838 -10671 15784 -10645
rect 16034 -10671 16612 -10645
rect -2918 -10871 -2340 -10845
rect -1906 -10871 -1876 -10845
rect -1822 -10871 -1792 -10845
rect -1538 -10871 -960 -10845
rect -802 -10871 -224 -10845
rect 26 -10871 236 -10845
rect 505 -10871 535 -10845
rect 600 -10871 700 -10845
rect 860 -10871 960 -10845
rect 1032 -10871 1062 -10845
rect 1314 -10871 1524 -10845
rect 1774 -10871 2352 -10845
rect 2602 -10871 2812 -10845
rect 3081 -10871 3111 -10845
rect 3176 -10871 3276 -10845
rect 3436 -10871 3536 -10845
rect 3608 -10871 3638 -10845
rect 3890 -10871 4100 -10845
rect 4350 -10871 4928 -10845
rect 5178 -10871 5388 -10845
rect 5657 -10871 5687 -10845
rect 5752 -10871 5852 -10845
rect 6012 -10871 6112 -10845
rect 6184 -10871 6214 -10845
rect 6466 -10871 6676 -10845
rect 6926 -10871 7504 -10845
rect 7754 -10871 7964 -10845
rect 8233 -10871 8263 -10845
rect 8328 -10871 8428 -10845
rect 8588 -10871 8688 -10845
rect 8760 -10871 8790 -10845
rect 9042 -10871 9252 -10845
rect 9502 -10871 10080 -10845
rect 10422 -10871 10632 -10845
rect 10809 -10871 10839 -10845
rect 10904 -10871 11004 -10845
rect 11164 -10871 11264 -10845
rect 11336 -10871 11366 -10845
rect 11710 -10871 11920 -10845
rect 13642 -10871 14588 -10845
rect 14838 -10871 15784 -10845
rect 16034 -10871 16612 -10845
rect -2918 -10939 -2340 -10913
rect -1538 -10939 -960 -10913
rect -802 -10939 -224 -10913
rect 26 -10939 236 -10913
rect 505 -10939 535 -10913
rect 600 -10939 700 -10913
rect 860 -10939 960 -10913
rect 1032 -10939 1062 -10913
rect 1314 -10939 1524 -10913
rect 1774 -10939 2352 -10913
rect 2602 -10939 2812 -10913
rect 3081 -10939 3111 -10913
rect 3176 -10939 3276 -10913
rect 3436 -10939 3536 -10913
rect 3608 -10939 3638 -10913
rect 3890 -10939 4100 -10913
rect 4350 -10939 4928 -10913
rect 5178 -10939 5388 -10913
rect 5657 -10939 5687 -10913
rect 5752 -10939 5852 -10913
rect 6012 -10939 6112 -10913
rect 6184 -10939 6214 -10913
rect 6466 -10939 6676 -10913
rect 6926 -10939 7504 -10913
rect 7754 -10939 7964 -10913
rect 8233 -10939 8263 -10913
rect 8328 -10939 8428 -10913
rect 8588 -10939 8688 -10913
rect 8760 -10939 8790 -10913
rect 9042 -10939 9252 -10913
rect 9502 -10939 10080 -10913
rect 10422 -10939 10632 -10913
rect 10809 -10939 10839 -10913
rect 10904 -10939 11004 -10913
rect 11164 -10939 11264 -10913
rect 11336 -10939 11366 -10913
rect 11710 -10939 11920 -10913
rect 13642 -10939 14588 -10913
rect 14838 -10939 15784 -10913
rect 16034 -10939 16612 -10913
rect -2918 -11139 -2340 -11113
rect -1538 -11139 -960 -11113
rect -802 -11139 -224 -11113
rect 26 -11139 236 -11113
rect -2918 -11161 -2654 -11139
rect -2918 -11195 -2902 -11161
rect -2868 -11195 -2803 -11161
rect -2769 -11195 -2704 -11161
rect -2670 -11195 -2654 -11161
rect -1224 -11161 -960 -11139
rect -2918 -11211 -2654 -11195
rect -2612 -11197 -2340 -11181
rect -2612 -11231 -2596 -11197
rect -2562 -11231 -2493 -11197
rect -2459 -11231 -2390 -11197
rect -2356 -11231 -2340 -11197
rect -2612 -11253 -2340 -11231
rect -2918 -11279 -2340 -11253
rect -1538 -11197 -1266 -11181
rect -1538 -11231 -1522 -11197
rect -1488 -11231 -1419 -11197
rect -1385 -11231 -1316 -11197
rect -1282 -11231 -1266 -11197
rect -1224 -11195 -1208 -11161
rect -1174 -11195 -1109 -11161
rect -1075 -11195 -1010 -11161
rect -976 -11195 -960 -11161
rect -488 -11161 -224 -11139
rect -1224 -11211 -960 -11195
rect -802 -11197 -530 -11181
rect -1538 -11253 -1266 -11231
rect -802 -11231 -786 -11197
rect -752 -11231 -683 -11197
rect -649 -11231 -580 -11197
rect -546 -11231 -530 -11197
rect -488 -11195 -472 -11161
rect -438 -11195 -373 -11161
rect -339 -11195 -274 -11161
rect -240 -11195 -224 -11161
rect 152 -11145 236 -11139
rect 152 -11161 294 -11145
rect -488 -11211 -224 -11195
rect -32 -11197 110 -11181
rect -802 -11253 -530 -11231
rect -32 -11231 -16 -11197
rect 18 -11231 110 -11197
rect 152 -11195 244 -11161
rect 278 -11195 294 -11161
rect 505 -11171 535 -11139
rect 152 -11211 294 -11195
rect 501 -11187 555 -11171
rect -32 -11247 110 -11231
rect 501 -11221 511 -11187
rect 545 -11221 555 -11187
rect 501 -11237 555 -11221
rect 600 -11177 700 -11103
rect 860 -11177 960 -11103
rect 1314 -11139 1524 -11113
rect 1032 -11174 1062 -11139
rect 1440 -11145 1524 -11139
rect 1774 -11139 2352 -11113
rect 2602 -11139 2812 -11113
rect 1440 -11161 1582 -11145
rect 600 -11187 761 -11177
rect 600 -11221 711 -11187
rect 745 -11221 761 -11187
rect 600 -11231 761 -11221
rect 860 -11187 982 -11177
rect 860 -11221 932 -11187
rect 966 -11221 982 -11187
rect 860 -11231 982 -11221
rect 1032 -11187 1102 -11174
rect 1032 -11221 1052 -11187
rect 1086 -11221 1102 -11187
rect 26 -11253 110 -11247
rect -1538 -11279 -960 -11253
rect -802 -11279 -224 -11253
rect 26 -11279 236 -11253
rect 505 -11305 535 -11237
rect 600 -11259 700 -11231
rect 860 -11259 960 -11231
rect 1032 -11233 1102 -11221
rect 1256 -11197 1398 -11181
rect 1256 -11231 1272 -11197
rect 1306 -11231 1398 -11197
rect 1440 -11195 1532 -11161
rect 1566 -11195 1582 -11161
rect 1440 -11211 1582 -11195
rect 1774 -11161 2038 -11139
rect 1774 -11195 1790 -11161
rect 1824 -11195 1889 -11161
rect 1923 -11195 1988 -11161
rect 2022 -11195 2038 -11161
rect 2728 -11145 2812 -11139
rect 2728 -11161 2870 -11145
rect 1774 -11211 2038 -11195
rect 2080 -11197 2352 -11181
rect 1032 -11305 1062 -11233
rect 1256 -11247 1398 -11231
rect 1314 -11253 1398 -11247
rect 2080 -11231 2096 -11197
rect 2130 -11231 2199 -11197
rect 2233 -11231 2302 -11197
rect 2336 -11231 2352 -11197
rect 2080 -11253 2352 -11231
rect 2544 -11197 2686 -11181
rect 2544 -11231 2560 -11197
rect 2594 -11231 2686 -11197
rect 2728 -11195 2820 -11161
rect 2854 -11195 2870 -11161
rect 3081 -11171 3111 -11139
rect 2728 -11211 2870 -11195
rect 3077 -11187 3131 -11171
rect 2544 -11247 2686 -11231
rect 3077 -11221 3087 -11187
rect 3121 -11221 3131 -11187
rect 3077 -11237 3131 -11221
rect 3176 -11177 3276 -11103
rect 3436 -11177 3536 -11103
rect 3890 -11139 4100 -11113
rect 3608 -11174 3638 -11139
rect 4016 -11145 4100 -11139
rect 4350 -11139 4928 -11113
rect 5178 -11139 5388 -11113
rect 4016 -11161 4158 -11145
rect 3176 -11187 3337 -11177
rect 3176 -11221 3287 -11187
rect 3321 -11221 3337 -11187
rect 3176 -11231 3337 -11221
rect 3436 -11187 3558 -11177
rect 3436 -11221 3508 -11187
rect 3542 -11221 3558 -11187
rect 3436 -11231 3558 -11221
rect 3608 -11187 3678 -11174
rect 3608 -11221 3628 -11187
rect 3662 -11221 3678 -11187
rect 1314 -11279 1524 -11253
rect 1774 -11279 2352 -11253
rect 2602 -11253 2686 -11247
rect 2602 -11279 2812 -11253
rect 3081 -11305 3111 -11237
rect 3176 -11259 3276 -11231
rect 3436 -11259 3536 -11231
rect 3608 -11233 3678 -11221
rect 3832 -11197 3974 -11181
rect 3832 -11231 3848 -11197
rect 3882 -11231 3974 -11197
rect 4016 -11195 4108 -11161
rect 4142 -11195 4158 -11161
rect 4016 -11211 4158 -11195
rect 4350 -11161 4614 -11139
rect 4350 -11195 4366 -11161
rect 4400 -11195 4465 -11161
rect 4499 -11195 4564 -11161
rect 4598 -11195 4614 -11161
rect 5304 -11145 5388 -11139
rect 5304 -11161 5446 -11145
rect 4350 -11211 4614 -11195
rect 4656 -11197 4928 -11181
rect 3608 -11305 3638 -11233
rect 3832 -11247 3974 -11231
rect 3890 -11253 3974 -11247
rect 4656 -11231 4672 -11197
rect 4706 -11231 4775 -11197
rect 4809 -11231 4878 -11197
rect 4912 -11231 4928 -11197
rect 4656 -11253 4928 -11231
rect 5120 -11197 5262 -11181
rect 5120 -11231 5136 -11197
rect 5170 -11231 5262 -11197
rect 5304 -11195 5396 -11161
rect 5430 -11195 5446 -11161
rect 5657 -11171 5687 -11139
rect 5304 -11211 5446 -11195
rect 5653 -11187 5707 -11171
rect 5120 -11247 5262 -11231
rect 5653 -11221 5663 -11187
rect 5697 -11221 5707 -11187
rect 5653 -11237 5707 -11221
rect 5752 -11177 5852 -11103
rect 6012 -11177 6112 -11103
rect 6466 -11139 6676 -11113
rect 6184 -11174 6214 -11139
rect 6592 -11145 6676 -11139
rect 6926 -11139 7504 -11113
rect 7754 -11139 7964 -11113
rect 6592 -11161 6734 -11145
rect 5752 -11187 5913 -11177
rect 5752 -11221 5863 -11187
rect 5897 -11221 5913 -11187
rect 5752 -11231 5913 -11221
rect 6012 -11187 6134 -11177
rect 6012 -11221 6084 -11187
rect 6118 -11221 6134 -11187
rect 6012 -11231 6134 -11221
rect 6184 -11187 6254 -11174
rect 6184 -11221 6204 -11187
rect 6238 -11221 6254 -11187
rect 3890 -11279 4100 -11253
rect 4350 -11279 4928 -11253
rect 5178 -11253 5262 -11247
rect 5178 -11279 5388 -11253
rect 5657 -11305 5687 -11237
rect 5752 -11259 5852 -11231
rect 6012 -11259 6112 -11231
rect 6184 -11233 6254 -11221
rect 6408 -11197 6550 -11181
rect 6408 -11231 6424 -11197
rect 6458 -11231 6550 -11197
rect 6592 -11195 6684 -11161
rect 6718 -11195 6734 -11161
rect 6592 -11211 6734 -11195
rect 6926 -11161 7190 -11139
rect 6926 -11195 6942 -11161
rect 6976 -11195 7041 -11161
rect 7075 -11195 7140 -11161
rect 7174 -11195 7190 -11161
rect 7880 -11145 7964 -11139
rect 7880 -11161 8022 -11145
rect 6926 -11211 7190 -11195
rect 7232 -11197 7504 -11181
rect 6184 -11305 6214 -11233
rect 6408 -11247 6550 -11231
rect 6466 -11253 6550 -11247
rect 7232 -11231 7248 -11197
rect 7282 -11231 7351 -11197
rect 7385 -11231 7454 -11197
rect 7488 -11231 7504 -11197
rect 7232 -11253 7504 -11231
rect 7696 -11197 7838 -11181
rect 7696 -11231 7712 -11197
rect 7746 -11231 7838 -11197
rect 7880 -11195 7972 -11161
rect 8006 -11195 8022 -11161
rect 8233 -11171 8263 -11139
rect 7880 -11211 8022 -11195
rect 8229 -11187 8283 -11171
rect 7696 -11247 7838 -11231
rect 8229 -11221 8239 -11187
rect 8273 -11221 8283 -11187
rect 8229 -11237 8283 -11221
rect 8328 -11177 8428 -11103
rect 8588 -11177 8688 -11103
rect 9042 -11139 9252 -11113
rect 8760 -11174 8790 -11139
rect 9168 -11145 9252 -11139
rect 9502 -11139 10080 -11113
rect 10422 -11139 10632 -11113
rect 9168 -11161 9310 -11145
rect 8328 -11187 8489 -11177
rect 8328 -11221 8439 -11187
rect 8473 -11221 8489 -11187
rect 8328 -11231 8489 -11221
rect 8588 -11187 8710 -11177
rect 8588 -11221 8660 -11187
rect 8694 -11221 8710 -11187
rect 8588 -11231 8710 -11221
rect 8760 -11187 8830 -11174
rect 8760 -11221 8780 -11187
rect 8814 -11221 8830 -11187
rect 6466 -11279 6676 -11253
rect 6926 -11279 7504 -11253
rect 7754 -11253 7838 -11247
rect 7754 -11279 7964 -11253
rect 8233 -11305 8263 -11237
rect 8328 -11259 8428 -11231
rect 8588 -11259 8688 -11231
rect 8760 -11233 8830 -11221
rect 8984 -11197 9126 -11181
rect 8984 -11231 9000 -11197
rect 9034 -11231 9126 -11197
rect 9168 -11195 9260 -11161
rect 9294 -11195 9310 -11161
rect 9168 -11211 9310 -11195
rect 9502 -11161 9766 -11139
rect 9502 -11195 9518 -11161
rect 9552 -11195 9617 -11161
rect 9651 -11195 9716 -11161
rect 9750 -11195 9766 -11161
rect 10548 -11145 10632 -11139
rect 10548 -11161 10690 -11145
rect 9502 -11211 9766 -11195
rect 9808 -11197 10080 -11181
rect 8760 -11305 8790 -11233
rect 8984 -11247 9126 -11231
rect 9042 -11253 9126 -11247
rect 9808 -11231 9824 -11197
rect 9858 -11231 9927 -11197
rect 9961 -11231 10030 -11197
rect 10064 -11231 10080 -11197
rect 9808 -11253 10080 -11231
rect 10364 -11197 10506 -11181
rect 10364 -11231 10380 -11197
rect 10414 -11231 10506 -11197
rect 10548 -11195 10640 -11161
rect 10674 -11195 10690 -11161
rect 10809 -11171 10839 -11139
rect 10548 -11211 10690 -11195
rect 10805 -11187 10859 -11171
rect 10364 -11247 10506 -11231
rect 10805 -11221 10815 -11187
rect 10849 -11221 10859 -11187
rect 10805 -11237 10859 -11221
rect 10904 -11177 11004 -11103
rect 11164 -11177 11264 -11103
rect 11710 -11139 11920 -11113
rect 13642 -11139 14588 -11113
rect 14838 -11139 15784 -11113
rect 16034 -11139 16612 -11113
rect 11336 -11174 11366 -11139
rect 11836 -11145 11920 -11139
rect 11836 -11161 11978 -11145
rect 10904 -11187 11065 -11177
rect 10904 -11221 11015 -11187
rect 11049 -11221 11065 -11187
rect 10904 -11231 11065 -11221
rect 11164 -11187 11286 -11177
rect 11164 -11221 11236 -11187
rect 11270 -11221 11286 -11187
rect 11164 -11231 11286 -11221
rect 11336 -11187 11406 -11174
rect 11336 -11221 11356 -11187
rect 11390 -11221 11406 -11187
rect 9042 -11279 9252 -11253
rect 9502 -11279 10080 -11253
rect 10422 -11253 10506 -11247
rect 10422 -11279 10632 -11253
rect 10809 -11305 10839 -11237
rect 10904 -11259 11004 -11231
rect 11164 -11259 11264 -11231
rect 11336 -11233 11406 -11221
rect 11652 -11197 11794 -11181
rect 11652 -11231 11668 -11197
rect 11702 -11231 11794 -11197
rect 11836 -11195 11928 -11161
rect 11962 -11195 11978 -11161
rect 14138 -11161 14588 -11139
rect 11836 -11211 11978 -11195
rect 13642 -11197 14096 -11181
rect 11336 -11305 11366 -11233
rect 11652 -11247 11794 -11231
rect 11710 -11253 11794 -11247
rect 13642 -11231 13662 -11197
rect 13696 -11231 13790 -11197
rect 13824 -11231 13918 -11197
rect 13952 -11231 14046 -11197
rect 14080 -11231 14096 -11197
rect 14138 -11195 14154 -11161
rect 14188 -11195 14282 -11161
rect 14316 -11195 14410 -11161
rect 14444 -11195 14538 -11161
rect 14572 -11195 14588 -11161
rect 15334 -11161 15784 -11139
rect 14138 -11211 14588 -11195
rect 14838 -11197 15292 -11181
rect 13642 -11253 14096 -11231
rect 14838 -11231 14858 -11197
rect 14892 -11231 14986 -11197
rect 15020 -11231 15114 -11197
rect 15148 -11231 15242 -11197
rect 15276 -11231 15292 -11197
rect 15334 -11195 15350 -11161
rect 15384 -11195 15478 -11161
rect 15512 -11195 15606 -11161
rect 15640 -11195 15734 -11161
rect 15768 -11195 15784 -11161
rect 16348 -11161 16612 -11139
rect 15334 -11211 15784 -11195
rect 16034 -11197 16306 -11181
rect 14838 -11253 15292 -11231
rect 16034 -11231 16050 -11197
rect 16084 -11231 16153 -11197
rect 16187 -11231 16256 -11197
rect 16290 -11231 16306 -11197
rect 16348 -11195 16364 -11161
rect 16398 -11195 16463 -11161
rect 16497 -11195 16562 -11161
rect 16596 -11195 16612 -11161
rect 16348 -11211 16612 -11195
rect 16034 -11253 16306 -11231
rect 11710 -11279 11920 -11253
rect 13642 -11279 14588 -11253
rect 14838 -11279 15784 -11253
rect 16034 -11279 16612 -11253
rect -2918 -11415 -2340 -11389
rect -1538 -11415 -960 -11389
rect -802 -11415 -224 -11389
rect 26 -11415 236 -11389
rect 505 -11415 535 -11389
rect 600 -11415 700 -11389
rect 860 -11415 960 -11389
rect 1032 -11415 1062 -11389
rect 1314 -11415 1524 -11389
rect 1774 -11415 2352 -11389
rect 2602 -11415 2812 -11389
rect 3081 -11415 3111 -11389
rect 3176 -11415 3276 -11389
rect 3436 -11415 3536 -11389
rect 3608 -11415 3638 -11389
rect 3890 -11415 4100 -11389
rect 4350 -11415 4928 -11389
rect 5178 -11415 5388 -11389
rect 5657 -11415 5687 -11389
rect 5752 -11415 5852 -11389
rect 6012 -11415 6112 -11389
rect 6184 -11415 6214 -11389
rect 6466 -11415 6676 -11389
rect 6926 -11415 7504 -11389
rect 7754 -11415 7964 -11389
rect 8233 -11415 8263 -11389
rect 8328 -11415 8428 -11389
rect 8588 -11415 8688 -11389
rect 8760 -11415 8790 -11389
rect 9042 -11415 9252 -11389
rect 9502 -11415 10080 -11389
rect 10422 -11415 10632 -11389
rect 10809 -11415 10839 -11389
rect 10904 -11415 11004 -11389
rect 11164 -11415 11264 -11389
rect 11336 -11415 11366 -11389
rect 11710 -11415 11920 -11389
rect 13642 -11415 14588 -11389
rect 14838 -11415 15784 -11389
rect 16034 -11415 16612 -11389
rect -2918 -11483 -2340 -11457
rect -1538 -11483 -960 -11457
rect -802 -11483 -224 -11457
rect 26 -11483 236 -11457
rect 488 -11483 518 -11457
rect 590 -11483 690 -11457
rect 850 -11483 950 -11457
rect 1015 -11483 1045 -11457
rect 1314 -11483 1524 -11457
rect 1774 -11483 2352 -11457
rect 2602 -11483 2812 -11457
rect 3064 -11483 3094 -11457
rect 3166 -11483 3266 -11457
rect 3426 -11483 3526 -11457
rect 3591 -11483 3621 -11457
rect 3890 -11483 4100 -11457
rect 4350 -11483 4928 -11457
rect 5178 -11483 5388 -11457
rect 5640 -11483 5670 -11457
rect 5742 -11483 5842 -11457
rect 6002 -11483 6102 -11457
rect 6167 -11483 6197 -11457
rect 6466 -11483 6676 -11457
rect 6926 -11483 7504 -11457
rect 7754 -11483 7964 -11457
rect 8216 -11483 8246 -11457
rect 8318 -11483 8418 -11457
rect 8578 -11483 8678 -11457
rect 8743 -11483 8773 -11457
rect 9042 -11483 9252 -11457
rect 9502 -11483 10080 -11457
rect 10422 -11483 10632 -11457
rect 10792 -11483 10822 -11457
rect 10894 -11483 10994 -11457
rect 11154 -11483 11254 -11457
rect 11319 -11483 11349 -11457
rect 11710 -11483 11920 -11457
rect 12633 -11483 12663 -11457
rect 12719 -11483 12749 -11457
rect 12805 -11483 12835 -11457
rect 12891 -11483 12921 -11457
rect 13274 -11483 13484 -11457
rect 13735 -11483 13765 -11457
rect 13821 -11483 13851 -11457
rect 13907 -11483 13937 -11457
rect 13993 -11483 14023 -11457
rect 14079 -11483 14109 -11457
rect 14165 -11483 14195 -11457
rect 14251 -11483 14281 -11457
rect 14337 -11483 14367 -11457
rect 14423 -11483 14453 -11457
rect 14509 -11483 14539 -11457
rect 14595 -11483 14625 -11457
rect 14681 -11483 14711 -11457
rect 14766 -11483 14796 -11457
rect 14852 -11483 14882 -11457
rect 14938 -11483 14968 -11457
rect 15024 -11483 15054 -11457
rect 15110 -11483 15140 -11457
rect 15196 -11483 15226 -11457
rect 15282 -11483 15312 -11457
rect 15368 -11483 15398 -11457
rect 15666 -11483 16612 -11457
rect -2918 -11619 -2340 -11593
rect -1538 -11619 -960 -11593
rect -802 -11619 -224 -11593
rect -2918 -11641 -2646 -11619
rect -2918 -11675 -2902 -11641
rect -2868 -11675 -2799 -11641
rect -2765 -11675 -2696 -11641
rect -2662 -11675 -2646 -11641
rect -1232 -11641 -960 -11619
rect -2918 -11691 -2646 -11675
rect -2604 -11677 -2340 -11661
rect -2604 -11711 -2588 -11677
rect -2554 -11711 -2489 -11677
rect -2455 -11711 -2390 -11677
rect -2356 -11711 -2340 -11677
rect -2604 -11733 -2340 -11711
rect -2918 -11759 -2340 -11733
rect -1538 -11677 -1274 -11661
rect -1538 -11711 -1522 -11677
rect -1488 -11711 -1423 -11677
rect -1389 -11711 -1324 -11677
rect -1290 -11711 -1274 -11677
rect -1232 -11675 -1216 -11641
rect -1182 -11675 -1113 -11641
rect -1079 -11675 -1010 -11641
rect -976 -11675 -960 -11641
rect -496 -11641 -224 -11619
rect 26 -11619 236 -11593
rect 26 -11625 110 -11619
rect -1232 -11691 -960 -11675
rect -802 -11677 -538 -11661
rect -1538 -11733 -1274 -11711
rect -802 -11711 -786 -11677
rect -752 -11711 -687 -11677
rect -653 -11711 -588 -11677
rect -554 -11711 -538 -11677
rect -496 -11675 -480 -11641
rect -446 -11675 -377 -11641
rect -343 -11675 -274 -11641
rect -240 -11675 -224 -11641
rect -496 -11691 -224 -11675
rect -32 -11641 110 -11625
rect 488 -11639 518 -11567
rect -32 -11675 -16 -11641
rect 18 -11675 110 -11641
rect 448 -11651 518 -11639
rect 590 -11641 690 -11613
rect 850 -11641 950 -11613
rect 1015 -11635 1045 -11567
rect 1314 -11619 1524 -11593
rect 1774 -11619 2352 -11593
rect 2602 -11619 2812 -11593
rect 1314 -11625 1398 -11619
rect -32 -11691 110 -11675
rect 152 -11677 294 -11661
rect -802 -11733 -538 -11711
rect 152 -11711 244 -11677
rect 278 -11711 294 -11677
rect 448 -11685 464 -11651
rect 498 -11685 518 -11651
rect 448 -11698 518 -11685
rect 568 -11651 690 -11641
rect 568 -11685 584 -11651
rect 618 -11685 690 -11651
rect 568 -11695 690 -11685
rect 789 -11651 950 -11641
rect 789 -11685 805 -11651
rect 839 -11685 950 -11651
rect 789 -11695 950 -11685
rect 152 -11727 294 -11711
rect 152 -11733 236 -11727
rect 488 -11733 518 -11698
rect -1538 -11759 -960 -11733
rect -802 -11759 -224 -11733
rect 26 -11759 236 -11733
rect 590 -11769 690 -11695
rect 850 -11769 950 -11695
rect 995 -11651 1049 -11635
rect 995 -11685 1005 -11651
rect 1039 -11685 1049 -11651
rect 995 -11701 1049 -11685
rect 1256 -11641 1398 -11625
rect 1256 -11675 1272 -11641
rect 1306 -11675 1398 -11641
rect 1774 -11641 2046 -11619
rect 2602 -11625 2686 -11619
rect 1256 -11691 1398 -11675
rect 1440 -11677 1582 -11661
rect 1015 -11733 1045 -11701
rect 1440 -11711 1532 -11677
rect 1566 -11711 1582 -11677
rect 1774 -11675 1790 -11641
rect 1824 -11675 1893 -11641
rect 1927 -11675 1996 -11641
rect 2030 -11675 2046 -11641
rect 2544 -11641 2686 -11625
rect 3064 -11639 3094 -11567
rect 1774 -11691 2046 -11675
rect 2088 -11677 2352 -11661
rect 1440 -11727 1582 -11711
rect 2088 -11711 2104 -11677
rect 2138 -11711 2203 -11677
rect 2237 -11711 2302 -11677
rect 2336 -11711 2352 -11677
rect 2544 -11675 2560 -11641
rect 2594 -11675 2686 -11641
rect 3024 -11651 3094 -11639
rect 3166 -11641 3266 -11613
rect 3426 -11641 3526 -11613
rect 3591 -11635 3621 -11567
rect 3890 -11619 4100 -11593
rect 4350 -11619 4928 -11593
rect 5178 -11619 5388 -11593
rect 3890 -11625 3974 -11619
rect 2544 -11691 2686 -11675
rect 2728 -11677 2870 -11661
rect 1440 -11733 1524 -11727
rect 2088 -11733 2352 -11711
rect 2728 -11711 2820 -11677
rect 2854 -11711 2870 -11677
rect 3024 -11685 3040 -11651
rect 3074 -11685 3094 -11651
rect 3024 -11698 3094 -11685
rect 3144 -11651 3266 -11641
rect 3144 -11685 3160 -11651
rect 3194 -11685 3266 -11651
rect 3144 -11695 3266 -11685
rect 3365 -11651 3526 -11641
rect 3365 -11685 3381 -11651
rect 3415 -11685 3526 -11651
rect 3365 -11695 3526 -11685
rect 2728 -11727 2870 -11711
rect 2728 -11733 2812 -11727
rect 3064 -11733 3094 -11698
rect 1314 -11759 1524 -11733
rect 1774 -11759 2352 -11733
rect 2602 -11759 2812 -11733
rect 3166 -11769 3266 -11695
rect 3426 -11769 3526 -11695
rect 3571 -11651 3625 -11635
rect 3571 -11685 3581 -11651
rect 3615 -11685 3625 -11651
rect 3571 -11701 3625 -11685
rect 3832 -11641 3974 -11625
rect 3832 -11675 3848 -11641
rect 3882 -11675 3974 -11641
rect 4350 -11641 4622 -11619
rect 5178 -11625 5262 -11619
rect 3832 -11691 3974 -11675
rect 4016 -11677 4158 -11661
rect 3591 -11733 3621 -11701
rect 4016 -11711 4108 -11677
rect 4142 -11711 4158 -11677
rect 4350 -11675 4366 -11641
rect 4400 -11675 4469 -11641
rect 4503 -11675 4572 -11641
rect 4606 -11675 4622 -11641
rect 5120 -11641 5262 -11625
rect 5640 -11639 5670 -11567
rect 4350 -11691 4622 -11675
rect 4664 -11677 4928 -11661
rect 4016 -11727 4158 -11711
rect 4664 -11711 4680 -11677
rect 4714 -11711 4779 -11677
rect 4813 -11711 4878 -11677
rect 4912 -11711 4928 -11677
rect 5120 -11675 5136 -11641
rect 5170 -11675 5262 -11641
rect 5600 -11651 5670 -11639
rect 5742 -11641 5842 -11613
rect 6002 -11641 6102 -11613
rect 6167 -11635 6197 -11567
rect 6466 -11619 6676 -11593
rect 6926 -11619 7504 -11593
rect 7754 -11619 7964 -11593
rect 6466 -11625 6550 -11619
rect 5120 -11691 5262 -11675
rect 5304 -11677 5446 -11661
rect 4016 -11733 4100 -11727
rect 4664 -11733 4928 -11711
rect 5304 -11711 5396 -11677
rect 5430 -11711 5446 -11677
rect 5600 -11685 5616 -11651
rect 5650 -11685 5670 -11651
rect 5600 -11698 5670 -11685
rect 5720 -11651 5842 -11641
rect 5720 -11685 5736 -11651
rect 5770 -11685 5842 -11651
rect 5720 -11695 5842 -11685
rect 5941 -11651 6102 -11641
rect 5941 -11685 5957 -11651
rect 5991 -11685 6102 -11651
rect 5941 -11695 6102 -11685
rect 5304 -11727 5446 -11711
rect 5304 -11733 5388 -11727
rect 5640 -11733 5670 -11698
rect 3890 -11759 4100 -11733
rect 4350 -11759 4928 -11733
rect 5178 -11759 5388 -11733
rect 5742 -11769 5842 -11695
rect 6002 -11769 6102 -11695
rect 6147 -11651 6201 -11635
rect 6147 -11685 6157 -11651
rect 6191 -11685 6201 -11651
rect 6147 -11701 6201 -11685
rect 6408 -11641 6550 -11625
rect 6408 -11675 6424 -11641
rect 6458 -11675 6550 -11641
rect 6926 -11641 7198 -11619
rect 7754 -11625 7838 -11619
rect 6408 -11691 6550 -11675
rect 6592 -11677 6734 -11661
rect 6167 -11733 6197 -11701
rect 6592 -11711 6684 -11677
rect 6718 -11711 6734 -11677
rect 6926 -11675 6942 -11641
rect 6976 -11675 7045 -11641
rect 7079 -11675 7148 -11641
rect 7182 -11675 7198 -11641
rect 7696 -11641 7838 -11625
rect 8216 -11639 8246 -11567
rect 6926 -11691 7198 -11675
rect 7240 -11677 7504 -11661
rect 6592 -11727 6734 -11711
rect 7240 -11711 7256 -11677
rect 7290 -11711 7355 -11677
rect 7389 -11711 7454 -11677
rect 7488 -11711 7504 -11677
rect 7696 -11675 7712 -11641
rect 7746 -11675 7838 -11641
rect 8176 -11651 8246 -11639
rect 8318 -11641 8418 -11613
rect 8578 -11641 8678 -11613
rect 8743 -11635 8773 -11567
rect 9042 -11619 9252 -11593
rect 9502 -11619 10080 -11593
rect 10422 -11619 10632 -11593
rect 9042 -11625 9126 -11619
rect 7696 -11691 7838 -11675
rect 7880 -11677 8022 -11661
rect 6592 -11733 6676 -11727
rect 7240 -11733 7504 -11711
rect 7880 -11711 7972 -11677
rect 8006 -11711 8022 -11677
rect 8176 -11685 8192 -11651
rect 8226 -11685 8246 -11651
rect 8176 -11698 8246 -11685
rect 8296 -11651 8418 -11641
rect 8296 -11685 8312 -11651
rect 8346 -11685 8418 -11651
rect 8296 -11695 8418 -11685
rect 8517 -11651 8678 -11641
rect 8517 -11685 8533 -11651
rect 8567 -11685 8678 -11651
rect 8517 -11695 8678 -11685
rect 7880 -11727 8022 -11711
rect 7880 -11733 7964 -11727
rect 8216 -11733 8246 -11698
rect 6466 -11759 6676 -11733
rect 6926 -11759 7504 -11733
rect 7754 -11759 7964 -11733
rect 8318 -11769 8418 -11695
rect 8578 -11769 8678 -11695
rect 8723 -11651 8777 -11635
rect 8723 -11685 8733 -11651
rect 8767 -11685 8777 -11651
rect 8723 -11701 8777 -11685
rect 8984 -11641 9126 -11625
rect 8984 -11675 9000 -11641
rect 9034 -11675 9126 -11641
rect 9502 -11641 9774 -11619
rect 10422 -11625 10506 -11619
rect 8984 -11691 9126 -11675
rect 9168 -11677 9310 -11661
rect 8743 -11733 8773 -11701
rect 9168 -11711 9260 -11677
rect 9294 -11711 9310 -11677
rect 9502 -11675 9518 -11641
rect 9552 -11675 9621 -11641
rect 9655 -11675 9724 -11641
rect 9758 -11675 9774 -11641
rect 10364 -11641 10506 -11625
rect 10792 -11639 10822 -11567
rect 9502 -11691 9774 -11675
rect 9816 -11677 10080 -11661
rect 9168 -11727 9310 -11711
rect 9816 -11711 9832 -11677
rect 9866 -11711 9931 -11677
rect 9965 -11711 10030 -11677
rect 10064 -11711 10080 -11677
rect 10364 -11675 10380 -11641
rect 10414 -11675 10506 -11641
rect 10752 -11651 10822 -11639
rect 10894 -11641 10994 -11613
rect 11154 -11641 11254 -11613
rect 11319 -11635 11349 -11567
rect 11710 -11619 11920 -11593
rect 11710 -11625 11794 -11619
rect 10364 -11691 10506 -11675
rect 10548 -11677 10690 -11661
rect 9168 -11733 9252 -11727
rect 9816 -11733 10080 -11711
rect 10548 -11711 10640 -11677
rect 10674 -11711 10690 -11677
rect 10752 -11685 10768 -11651
rect 10802 -11685 10822 -11651
rect 10752 -11698 10822 -11685
rect 10872 -11651 10994 -11641
rect 10872 -11685 10888 -11651
rect 10922 -11685 10994 -11651
rect 10872 -11695 10994 -11685
rect 11093 -11651 11254 -11641
rect 11093 -11685 11109 -11651
rect 11143 -11685 11254 -11651
rect 11093 -11695 11254 -11685
rect 10548 -11727 10690 -11711
rect 10548 -11733 10632 -11727
rect 10792 -11733 10822 -11698
rect 9042 -11759 9252 -11733
rect 9502 -11759 10080 -11733
rect 10422 -11759 10632 -11733
rect 10894 -11769 10994 -11695
rect 11154 -11769 11254 -11695
rect 11299 -11651 11353 -11635
rect 11299 -11685 11309 -11651
rect 11343 -11685 11353 -11651
rect 11299 -11701 11353 -11685
rect 11652 -11641 11794 -11625
rect 12633 -11641 12663 -11567
rect 12719 -11641 12749 -11567
rect 12805 -11641 12835 -11567
rect 12891 -11641 12921 -11567
rect 13274 -11619 13484 -11593
rect 13735 -11616 13765 -11567
rect 13821 -11616 13851 -11567
rect 13907 -11616 13937 -11567
rect 13993 -11616 14023 -11567
rect 13400 -11625 13484 -11619
rect 13400 -11641 13542 -11625
rect 11652 -11675 11668 -11641
rect 11702 -11675 11794 -11641
rect 12547 -11651 13007 -11641
rect 11652 -11691 11794 -11675
rect 11836 -11677 11978 -11661
rect 11319 -11733 11349 -11701
rect 11836 -11711 11928 -11677
rect 11962 -11711 11978 -11677
rect 11836 -11727 11978 -11711
rect 12547 -11685 12574 -11651
rect 12608 -11685 12642 -11651
rect 12676 -11685 12710 -11651
rect 12744 -11685 12778 -11651
rect 12812 -11685 12846 -11651
rect 12880 -11685 12914 -11651
rect 12948 -11685 13007 -11651
rect 12547 -11695 13007 -11685
rect 11836 -11733 11920 -11727
rect 12547 -11733 12577 -11695
rect 12633 -11733 12663 -11695
rect 12719 -11733 12749 -11695
rect 12805 -11733 12835 -11695
rect 12891 -11733 12921 -11695
rect 12977 -11733 13007 -11695
rect 13216 -11677 13358 -11661
rect 13216 -11711 13232 -11677
rect 13266 -11711 13358 -11677
rect 13400 -11675 13492 -11641
rect 13526 -11675 13542 -11641
rect 13400 -11691 13542 -11675
rect 13676 -11651 14023 -11616
rect 13676 -11685 13692 -11651
rect 13726 -11685 14023 -11651
rect 13216 -11727 13358 -11711
rect 13676 -11718 14023 -11685
rect 13274 -11733 13358 -11727
rect 13735 -11733 13765 -11718
rect 13821 -11733 13851 -11718
rect 13907 -11733 13937 -11718
rect 13993 -11733 14023 -11718
rect 14079 -11626 14109 -11567
rect 14165 -11626 14195 -11567
rect 14251 -11626 14281 -11567
rect 14337 -11626 14367 -11567
rect 14423 -11626 14453 -11567
rect 14509 -11626 14539 -11567
rect 14595 -11626 14625 -11567
rect 14681 -11626 14711 -11567
rect 14766 -11626 14796 -11567
rect 14852 -11626 14882 -11567
rect 14938 -11626 14968 -11567
rect 15024 -11626 15054 -11567
rect 15110 -11626 15140 -11567
rect 15196 -11626 15226 -11567
rect 15282 -11626 15312 -11567
rect 15368 -11626 15398 -11567
rect 15666 -11619 16612 -11593
rect 14079 -11651 15398 -11626
rect 14079 -11685 14119 -11651
rect 14153 -11685 14187 -11651
rect 14221 -11685 14255 -11651
rect 14289 -11685 14323 -11651
rect 14357 -11685 14391 -11651
rect 14425 -11685 14459 -11651
rect 14493 -11685 14527 -11651
rect 14561 -11685 14595 -11651
rect 14629 -11685 14663 -11651
rect 14697 -11685 14731 -11651
rect 14765 -11685 14799 -11651
rect 14833 -11685 14867 -11651
rect 14901 -11685 14935 -11651
rect 14969 -11685 15003 -11651
rect 15037 -11685 15071 -11651
rect 15105 -11685 15139 -11651
rect 15173 -11685 15398 -11651
rect 16158 -11641 16612 -11619
rect 14079 -11701 15398 -11685
rect 14079 -11733 14109 -11701
rect 14165 -11733 14195 -11701
rect 14251 -11733 14281 -11701
rect 14337 -11733 14367 -11701
rect 14423 -11733 14453 -11701
rect 14509 -11733 14539 -11701
rect 14595 -11733 14625 -11701
rect 14681 -11733 14711 -11701
rect 14766 -11733 14796 -11701
rect 14852 -11733 14882 -11701
rect 14938 -11733 14968 -11701
rect 15024 -11733 15054 -11701
rect 15110 -11733 15140 -11701
rect 15196 -11733 15226 -11701
rect 15282 -11733 15312 -11701
rect 15368 -11733 15398 -11701
rect 15666 -11677 16116 -11661
rect 15666 -11711 15682 -11677
rect 15716 -11711 15810 -11677
rect 15844 -11711 15938 -11677
rect 15972 -11711 16066 -11677
rect 16100 -11711 16116 -11677
rect 16158 -11675 16174 -11641
rect 16208 -11675 16302 -11641
rect 16336 -11675 16430 -11641
rect 16464 -11675 16558 -11641
rect 16592 -11675 16612 -11641
rect 16158 -11691 16612 -11675
rect 15666 -11733 16116 -11711
rect 11710 -11759 11920 -11733
rect 13274 -11759 13484 -11733
rect 15666 -11759 16612 -11733
rect -2918 -11959 -2340 -11933
rect -1538 -11959 -960 -11933
rect -802 -11959 -224 -11933
rect 26 -11959 236 -11933
rect 488 -11959 518 -11933
rect 590 -11959 690 -11933
rect 850 -11959 950 -11933
rect 1015 -11959 1045 -11933
rect 1314 -11959 1524 -11933
rect 1774 -11959 2352 -11933
rect 2602 -11959 2812 -11933
rect 3064 -11959 3094 -11933
rect 3166 -11959 3266 -11933
rect 3426 -11959 3526 -11933
rect 3591 -11959 3621 -11933
rect 3890 -11959 4100 -11933
rect 4350 -11959 4928 -11933
rect 5178 -11959 5388 -11933
rect 5640 -11959 5670 -11933
rect 5742 -11959 5842 -11933
rect 6002 -11959 6102 -11933
rect 6167 -11959 6197 -11933
rect 6466 -11959 6676 -11933
rect 6926 -11959 7504 -11933
rect 7754 -11959 7964 -11933
rect 8216 -11959 8246 -11933
rect 8318 -11959 8418 -11933
rect 8578 -11959 8678 -11933
rect 8743 -11959 8773 -11933
rect 9042 -11959 9252 -11933
rect 9502 -11959 10080 -11933
rect 10422 -11959 10632 -11933
rect 10792 -11959 10822 -11933
rect 10894 -11959 10994 -11933
rect 11154 -11959 11254 -11933
rect 11319 -11959 11349 -11933
rect 11710 -11959 11920 -11933
rect 12547 -11959 12577 -11933
rect 12633 -11959 12663 -11933
rect 12719 -11959 12749 -11933
rect 12805 -11959 12835 -11933
rect 12891 -11959 12921 -11933
rect 12977 -11959 13007 -11933
rect 13274 -11959 13484 -11933
rect 13735 -11959 13765 -11933
rect 13821 -11959 13851 -11933
rect 13907 -11959 13937 -11933
rect 13993 -11959 14023 -11933
rect 14079 -11959 14109 -11933
rect 14165 -11959 14195 -11933
rect 14251 -11959 14281 -11933
rect 14337 -11959 14367 -11933
rect 14423 -11959 14453 -11933
rect 14509 -11959 14539 -11933
rect 14595 -11959 14625 -11933
rect 14681 -11959 14711 -11933
rect 14766 -11959 14796 -11933
rect 14852 -11959 14882 -11933
rect 14938 -11959 14968 -11933
rect 15024 -11959 15054 -11933
rect 15110 -11959 15140 -11933
rect 15196 -11959 15226 -11933
rect 15282 -11959 15312 -11933
rect 15368 -11959 15398 -11933
rect 15666 -11959 16612 -11933
rect -2918 -12027 -2340 -12001
rect -1538 -12027 -960 -12001
rect -783 -12027 -753 -12001
rect -688 -12027 -588 -12001
rect -428 -12027 -328 -12001
rect -256 -12027 -226 -12001
rect 26 -12027 236 -12001
rect 505 -12027 535 -12001
rect 600 -12027 700 -12001
rect 860 -12027 960 -12001
rect 1032 -12027 1062 -12001
rect 1314 -12027 1524 -12001
rect 1774 -12027 2352 -12001
rect 2602 -12027 2812 -12001
rect 3081 -12027 3111 -12001
rect 3176 -12027 3276 -12001
rect 3436 -12027 3536 -12001
rect 3608 -12027 3638 -12001
rect 3890 -12027 4100 -12001
rect 4350 -12027 4928 -12001
rect 5178 -12027 5388 -12001
rect 5657 -12027 5687 -12001
rect 5752 -12027 5852 -12001
rect 6012 -12027 6112 -12001
rect 6184 -12027 6214 -12001
rect 6466 -12027 6676 -12001
rect 6926 -12027 7504 -12001
rect 7754 -12027 7964 -12001
rect 8233 -12027 8263 -12001
rect 8328 -12027 8428 -12001
rect 8588 -12027 8688 -12001
rect 8760 -12027 8790 -12001
rect 9042 -12027 9252 -12001
rect 9502 -12027 10080 -12001
rect 10422 -12027 10632 -12001
rect 10809 -12027 10839 -12001
rect 10904 -12027 11004 -12001
rect 11164 -12027 11264 -12001
rect 11336 -12027 11366 -12001
rect 11710 -12027 11920 -12001
rect 13735 -12027 13765 -12001
rect 13821 -12027 13851 -12001
rect 13907 -12027 13937 -12001
rect 13993 -12027 14023 -12001
rect 14079 -12027 14109 -12001
rect 14165 -12027 14195 -12001
rect 14251 -12027 14281 -12001
rect 14337 -12027 14367 -12001
rect 14423 -12027 14453 -12001
rect 14509 -12027 14539 -12001
rect 14595 -12027 14625 -12001
rect 14681 -12027 14711 -12001
rect 14766 -12027 14796 -12001
rect 14852 -12027 14882 -12001
rect 14938 -12027 14968 -12001
rect 15024 -12027 15054 -12001
rect 15110 -12027 15140 -12001
rect 15196 -12027 15226 -12001
rect 15282 -12027 15312 -12001
rect 15368 -12027 15398 -12001
rect 15666 -12027 16612 -12001
rect -2918 -12227 -2340 -12201
rect -1538 -12227 -960 -12201
rect -2918 -12249 -2654 -12227
rect -2918 -12283 -2902 -12249
rect -2868 -12283 -2803 -12249
rect -2769 -12283 -2704 -12249
rect -2670 -12283 -2654 -12249
rect -1224 -12249 -960 -12227
rect -2918 -12299 -2654 -12283
rect -2612 -12285 -2340 -12269
rect -2612 -12319 -2596 -12285
rect -2562 -12319 -2493 -12285
rect -2459 -12319 -2390 -12285
rect -2356 -12319 -2340 -12285
rect -2612 -12341 -2340 -12319
rect -2918 -12367 -2340 -12341
rect -1538 -12285 -1266 -12269
rect -1538 -12319 -1522 -12285
rect -1488 -12319 -1419 -12285
rect -1385 -12319 -1316 -12285
rect -1282 -12319 -1266 -12285
rect -1224 -12283 -1208 -12249
rect -1174 -12283 -1109 -12249
rect -1075 -12283 -1010 -12249
rect -976 -12283 -960 -12249
rect -783 -12259 -753 -12227
rect -1224 -12299 -960 -12283
rect -787 -12275 -733 -12259
rect -1538 -12341 -1266 -12319
rect -787 -12309 -777 -12275
rect -743 -12309 -733 -12275
rect -787 -12325 -733 -12309
rect -688 -12265 -588 -12191
rect -428 -12265 -328 -12191
rect 26 -12227 236 -12201
rect -256 -12262 -226 -12227
rect 152 -12233 236 -12227
rect 152 -12249 294 -12233
rect -688 -12275 -527 -12265
rect -688 -12309 -577 -12275
rect -543 -12309 -527 -12275
rect -688 -12319 -527 -12309
rect -428 -12275 -306 -12265
rect -428 -12309 -356 -12275
rect -322 -12309 -306 -12275
rect -428 -12319 -306 -12309
rect -256 -12275 -186 -12262
rect -256 -12309 -236 -12275
rect -202 -12309 -186 -12275
rect -1538 -12367 -960 -12341
rect -783 -12393 -753 -12325
rect -688 -12347 -588 -12319
rect -428 -12347 -328 -12319
rect -256 -12321 -186 -12309
rect -32 -12285 110 -12269
rect -32 -12319 -16 -12285
rect 18 -12319 110 -12285
rect 152 -12283 244 -12249
rect 278 -12283 294 -12249
rect 505 -12259 535 -12227
rect 152 -12299 294 -12283
rect 501 -12275 555 -12259
rect -256 -12393 -226 -12321
rect -32 -12335 110 -12319
rect 501 -12309 511 -12275
rect 545 -12309 555 -12275
rect 501 -12325 555 -12309
rect 600 -12265 700 -12191
rect 860 -12265 960 -12191
rect 1314 -12227 1524 -12201
rect 1032 -12262 1062 -12227
rect 1440 -12233 1524 -12227
rect 1774 -12227 2352 -12201
rect 2602 -12227 2812 -12201
rect 1440 -12249 1582 -12233
rect 600 -12275 761 -12265
rect 600 -12309 711 -12275
rect 745 -12309 761 -12275
rect 600 -12319 761 -12309
rect 860 -12275 982 -12265
rect 860 -12309 932 -12275
rect 966 -12309 982 -12275
rect 860 -12319 982 -12309
rect 1032 -12275 1102 -12262
rect 1032 -12309 1052 -12275
rect 1086 -12309 1102 -12275
rect 26 -12341 110 -12335
rect 26 -12367 236 -12341
rect 505 -12393 535 -12325
rect 600 -12347 700 -12319
rect 860 -12347 960 -12319
rect 1032 -12321 1102 -12309
rect 1256 -12285 1398 -12269
rect 1256 -12319 1272 -12285
rect 1306 -12319 1398 -12285
rect 1440 -12283 1532 -12249
rect 1566 -12283 1582 -12249
rect 1440 -12299 1582 -12283
rect 1774 -12249 2038 -12227
rect 1774 -12283 1790 -12249
rect 1824 -12283 1889 -12249
rect 1923 -12283 1988 -12249
rect 2022 -12283 2038 -12249
rect 2728 -12233 2812 -12227
rect 2728 -12249 2870 -12233
rect 1774 -12299 2038 -12283
rect 2080 -12285 2352 -12269
rect 1032 -12393 1062 -12321
rect 1256 -12335 1398 -12319
rect 1314 -12341 1398 -12335
rect 2080 -12319 2096 -12285
rect 2130 -12319 2199 -12285
rect 2233 -12319 2302 -12285
rect 2336 -12319 2352 -12285
rect 2080 -12341 2352 -12319
rect 2544 -12285 2686 -12269
rect 2544 -12319 2560 -12285
rect 2594 -12319 2686 -12285
rect 2728 -12283 2820 -12249
rect 2854 -12283 2870 -12249
rect 3081 -12259 3111 -12227
rect 2728 -12299 2870 -12283
rect 3077 -12275 3131 -12259
rect 2544 -12335 2686 -12319
rect 3077 -12309 3087 -12275
rect 3121 -12309 3131 -12275
rect 3077 -12325 3131 -12309
rect 3176 -12265 3276 -12191
rect 3436 -12265 3536 -12191
rect 3890 -12227 4100 -12201
rect 3608 -12262 3638 -12227
rect 4016 -12233 4100 -12227
rect 4350 -12227 4928 -12201
rect 5178 -12227 5388 -12201
rect 4016 -12249 4158 -12233
rect 3176 -12275 3337 -12265
rect 3176 -12309 3287 -12275
rect 3321 -12309 3337 -12275
rect 3176 -12319 3337 -12309
rect 3436 -12275 3558 -12265
rect 3436 -12309 3508 -12275
rect 3542 -12309 3558 -12275
rect 3436 -12319 3558 -12309
rect 3608 -12275 3678 -12262
rect 3608 -12309 3628 -12275
rect 3662 -12309 3678 -12275
rect 1314 -12367 1524 -12341
rect 1774 -12367 2352 -12341
rect 2602 -12341 2686 -12335
rect 2602 -12367 2812 -12341
rect 3081 -12393 3111 -12325
rect 3176 -12347 3276 -12319
rect 3436 -12347 3536 -12319
rect 3608 -12321 3678 -12309
rect 3832 -12285 3974 -12269
rect 3832 -12319 3848 -12285
rect 3882 -12319 3974 -12285
rect 4016 -12283 4108 -12249
rect 4142 -12283 4158 -12249
rect 4016 -12299 4158 -12283
rect 4350 -12249 4614 -12227
rect 4350 -12283 4366 -12249
rect 4400 -12283 4465 -12249
rect 4499 -12283 4564 -12249
rect 4598 -12283 4614 -12249
rect 5304 -12233 5388 -12227
rect 5304 -12249 5446 -12233
rect 4350 -12299 4614 -12283
rect 4656 -12285 4928 -12269
rect 3608 -12393 3638 -12321
rect 3832 -12335 3974 -12319
rect 3890 -12341 3974 -12335
rect 4656 -12319 4672 -12285
rect 4706 -12319 4775 -12285
rect 4809 -12319 4878 -12285
rect 4912 -12319 4928 -12285
rect 4656 -12341 4928 -12319
rect 5120 -12285 5262 -12269
rect 5120 -12319 5136 -12285
rect 5170 -12319 5262 -12285
rect 5304 -12283 5396 -12249
rect 5430 -12283 5446 -12249
rect 5657 -12259 5687 -12227
rect 5304 -12299 5446 -12283
rect 5653 -12275 5707 -12259
rect 5120 -12335 5262 -12319
rect 5653 -12309 5663 -12275
rect 5697 -12309 5707 -12275
rect 5653 -12325 5707 -12309
rect 5752 -12265 5852 -12191
rect 6012 -12265 6112 -12191
rect 6466 -12227 6676 -12201
rect 6184 -12262 6214 -12227
rect 6592 -12233 6676 -12227
rect 6926 -12227 7504 -12201
rect 7754 -12227 7964 -12201
rect 6592 -12249 6734 -12233
rect 5752 -12275 5913 -12265
rect 5752 -12309 5863 -12275
rect 5897 -12309 5913 -12275
rect 5752 -12319 5913 -12309
rect 6012 -12275 6134 -12265
rect 6012 -12309 6084 -12275
rect 6118 -12309 6134 -12275
rect 6012 -12319 6134 -12309
rect 6184 -12275 6254 -12262
rect 6184 -12309 6204 -12275
rect 6238 -12309 6254 -12275
rect 3890 -12367 4100 -12341
rect 4350 -12367 4928 -12341
rect 5178 -12341 5262 -12335
rect 5178 -12367 5388 -12341
rect 5657 -12393 5687 -12325
rect 5752 -12347 5852 -12319
rect 6012 -12347 6112 -12319
rect 6184 -12321 6254 -12309
rect 6408 -12285 6550 -12269
rect 6408 -12319 6424 -12285
rect 6458 -12319 6550 -12285
rect 6592 -12283 6684 -12249
rect 6718 -12283 6734 -12249
rect 6592 -12299 6734 -12283
rect 6926 -12249 7190 -12227
rect 6926 -12283 6942 -12249
rect 6976 -12283 7041 -12249
rect 7075 -12283 7140 -12249
rect 7174 -12283 7190 -12249
rect 7880 -12233 7964 -12227
rect 7880 -12249 8022 -12233
rect 6926 -12299 7190 -12283
rect 7232 -12285 7504 -12269
rect 6184 -12393 6214 -12321
rect 6408 -12335 6550 -12319
rect 6466 -12341 6550 -12335
rect 7232 -12319 7248 -12285
rect 7282 -12319 7351 -12285
rect 7385 -12319 7454 -12285
rect 7488 -12319 7504 -12285
rect 7232 -12341 7504 -12319
rect 7696 -12285 7838 -12269
rect 7696 -12319 7712 -12285
rect 7746 -12319 7838 -12285
rect 7880 -12283 7972 -12249
rect 8006 -12283 8022 -12249
rect 8233 -12259 8263 -12227
rect 7880 -12299 8022 -12283
rect 8229 -12275 8283 -12259
rect 7696 -12335 7838 -12319
rect 8229 -12309 8239 -12275
rect 8273 -12309 8283 -12275
rect 8229 -12325 8283 -12309
rect 8328 -12265 8428 -12191
rect 8588 -12265 8688 -12191
rect 9042 -12227 9252 -12201
rect 8760 -12262 8790 -12227
rect 9168 -12233 9252 -12227
rect 9502 -12227 10080 -12201
rect 10422 -12227 10632 -12201
rect 9168 -12249 9310 -12233
rect 8328 -12275 8489 -12265
rect 8328 -12309 8439 -12275
rect 8473 -12309 8489 -12275
rect 8328 -12319 8489 -12309
rect 8588 -12275 8710 -12265
rect 8588 -12309 8660 -12275
rect 8694 -12309 8710 -12275
rect 8588 -12319 8710 -12309
rect 8760 -12275 8830 -12262
rect 8760 -12309 8780 -12275
rect 8814 -12309 8830 -12275
rect 6466 -12367 6676 -12341
rect 6926 -12367 7504 -12341
rect 7754 -12341 7838 -12335
rect 7754 -12367 7964 -12341
rect 8233 -12393 8263 -12325
rect 8328 -12347 8428 -12319
rect 8588 -12347 8688 -12319
rect 8760 -12321 8830 -12309
rect 8984 -12285 9126 -12269
rect 8984 -12319 9000 -12285
rect 9034 -12319 9126 -12285
rect 9168 -12283 9260 -12249
rect 9294 -12283 9310 -12249
rect 9168 -12299 9310 -12283
rect 9502 -12249 9766 -12227
rect 9502 -12283 9518 -12249
rect 9552 -12283 9617 -12249
rect 9651 -12283 9716 -12249
rect 9750 -12283 9766 -12249
rect 10548 -12233 10632 -12227
rect 10548 -12249 10690 -12233
rect 9502 -12299 9766 -12283
rect 9808 -12285 10080 -12269
rect 8760 -12393 8790 -12321
rect 8984 -12335 9126 -12319
rect 9042 -12341 9126 -12335
rect 9808 -12319 9824 -12285
rect 9858 -12319 9927 -12285
rect 9961 -12319 10030 -12285
rect 10064 -12319 10080 -12285
rect 9808 -12341 10080 -12319
rect 10364 -12285 10506 -12269
rect 10364 -12319 10380 -12285
rect 10414 -12319 10506 -12285
rect 10548 -12283 10640 -12249
rect 10674 -12283 10690 -12249
rect 10809 -12259 10839 -12227
rect 10548 -12299 10690 -12283
rect 10805 -12275 10859 -12259
rect 10364 -12335 10506 -12319
rect 10805 -12309 10815 -12275
rect 10849 -12309 10859 -12275
rect 10805 -12325 10859 -12309
rect 10904 -12265 11004 -12191
rect 11164 -12265 11264 -12191
rect 11710 -12227 11920 -12201
rect 15666 -12227 16612 -12201
rect 11336 -12262 11366 -12227
rect 11836 -12233 11920 -12227
rect 11836 -12249 11978 -12233
rect 13735 -12242 13765 -12227
rect 13821 -12242 13851 -12227
rect 13907 -12242 13937 -12227
rect 13993 -12242 14023 -12227
rect 10904 -12275 11065 -12265
rect 10904 -12309 11015 -12275
rect 11049 -12309 11065 -12275
rect 10904 -12319 11065 -12309
rect 11164 -12275 11286 -12265
rect 11164 -12309 11236 -12275
rect 11270 -12309 11286 -12275
rect 11164 -12319 11286 -12309
rect 11336 -12275 11406 -12262
rect 11336 -12309 11356 -12275
rect 11390 -12309 11406 -12275
rect 9042 -12367 9252 -12341
rect 9502 -12367 10080 -12341
rect 10422 -12341 10506 -12335
rect 10422 -12367 10632 -12341
rect 10809 -12393 10839 -12325
rect 10904 -12347 11004 -12319
rect 11164 -12347 11264 -12319
rect 11336 -12321 11406 -12309
rect 11652 -12285 11794 -12269
rect 11652 -12319 11668 -12285
rect 11702 -12319 11794 -12285
rect 11836 -12283 11928 -12249
rect 11962 -12283 11978 -12249
rect 11836 -12299 11978 -12283
rect 13676 -12275 14023 -12242
rect 11336 -12393 11366 -12321
rect 11652 -12335 11794 -12319
rect 11710 -12341 11794 -12335
rect 13676 -12309 13692 -12275
rect 13726 -12309 14023 -12275
rect 11710 -12367 11920 -12341
rect 13676 -12344 14023 -12309
rect 13735 -12393 13765 -12344
rect 13821 -12393 13851 -12344
rect 13907 -12393 13937 -12344
rect 13993 -12393 14023 -12344
rect 14079 -12259 14109 -12227
rect 14165 -12259 14195 -12227
rect 14251 -12259 14281 -12227
rect 14337 -12259 14367 -12227
rect 14423 -12259 14453 -12227
rect 14509 -12259 14539 -12227
rect 14595 -12259 14625 -12227
rect 14681 -12259 14711 -12227
rect 14766 -12259 14796 -12227
rect 14852 -12259 14882 -12227
rect 14938 -12259 14968 -12227
rect 15024 -12259 15054 -12227
rect 15110 -12259 15140 -12227
rect 15196 -12259 15226 -12227
rect 15282 -12259 15312 -12227
rect 15368 -12259 15398 -12227
rect 14079 -12275 15398 -12259
rect 16162 -12249 16612 -12227
rect 14079 -12309 14119 -12275
rect 14153 -12309 14187 -12275
rect 14221 -12309 14255 -12275
rect 14289 -12309 14323 -12275
rect 14357 -12309 14391 -12275
rect 14425 -12309 14459 -12275
rect 14493 -12309 14527 -12275
rect 14561 -12309 14595 -12275
rect 14629 -12309 14663 -12275
rect 14697 -12309 14731 -12275
rect 14765 -12309 14799 -12275
rect 14833 -12309 14867 -12275
rect 14901 -12309 14935 -12275
rect 14969 -12309 15003 -12275
rect 15037 -12309 15071 -12275
rect 15105 -12309 15139 -12275
rect 15173 -12309 15398 -12275
rect 14079 -12334 15398 -12309
rect 14079 -12393 14109 -12334
rect 14165 -12393 14195 -12334
rect 14251 -12393 14281 -12334
rect 14337 -12393 14367 -12334
rect 14423 -12393 14453 -12334
rect 14509 -12393 14539 -12334
rect 14595 -12393 14625 -12334
rect 14681 -12393 14711 -12334
rect 14766 -12393 14796 -12334
rect 14852 -12393 14882 -12334
rect 14938 -12393 14968 -12334
rect 15024 -12393 15054 -12334
rect 15110 -12393 15140 -12334
rect 15196 -12393 15226 -12334
rect 15282 -12393 15312 -12334
rect 15368 -12393 15398 -12334
rect 15666 -12285 16120 -12269
rect 15666 -12319 15686 -12285
rect 15720 -12319 15814 -12285
rect 15848 -12319 15942 -12285
rect 15976 -12319 16070 -12285
rect 16104 -12319 16120 -12285
rect 16162 -12283 16178 -12249
rect 16212 -12283 16306 -12249
rect 16340 -12283 16434 -12249
rect 16468 -12283 16562 -12249
rect 16596 -12283 16612 -12249
rect 16162 -12299 16612 -12283
rect 15666 -12341 16120 -12319
rect 15666 -12367 16612 -12341
rect -2918 -12503 -2340 -12477
rect -1538 -12503 -960 -12477
rect -783 -12503 -753 -12477
rect -688 -12503 -588 -12477
rect -428 -12503 -328 -12477
rect -256 -12503 -226 -12477
rect 26 -12503 236 -12477
rect 505 -12503 535 -12477
rect 600 -12503 700 -12477
rect 860 -12503 960 -12477
rect 1032 -12503 1062 -12477
rect 1314 -12503 1524 -12477
rect 1774 -12503 2352 -12477
rect 2602 -12503 2812 -12477
rect 3081 -12503 3111 -12477
rect 3176 -12503 3276 -12477
rect 3436 -12503 3536 -12477
rect 3608 -12503 3638 -12477
rect 3890 -12503 4100 -12477
rect 4350 -12503 4928 -12477
rect 5178 -12503 5388 -12477
rect 5657 -12503 5687 -12477
rect 5752 -12503 5852 -12477
rect 6012 -12503 6112 -12477
rect 6184 -12503 6214 -12477
rect 6466 -12503 6676 -12477
rect 6926 -12503 7504 -12477
rect 7754 -12503 7964 -12477
rect 8233 -12503 8263 -12477
rect 8328 -12503 8428 -12477
rect 8588 -12503 8688 -12477
rect 8760 -12503 8790 -12477
rect 9042 -12503 9252 -12477
rect 9502 -12503 10080 -12477
rect 10422 -12503 10632 -12477
rect 10809 -12503 10839 -12477
rect 10904 -12503 11004 -12477
rect 11164 -12503 11264 -12477
rect 11336 -12503 11366 -12477
rect 11710 -12503 11920 -12477
rect 13735 -12503 13765 -12477
rect 13821 -12503 13851 -12477
rect 13907 -12503 13937 -12477
rect 13993 -12503 14023 -12477
rect 14079 -12503 14109 -12477
rect 14165 -12503 14195 -12477
rect 14251 -12503 14281 -12477
rect 14337 -12503 14367 -12477
rect 14423 -12503 14453 -12477
rect 14509 -12503 14539 -12477
rect 14595 -12503 14625 -12477
rect 14681 -12503 14711 -12477
rect 14766 -12503 14796 -12477
rect 14852 -12503 14882 -12477
rect 14938 -12503 14968 -12477
rect 15024 -12503 15054 -12477
rect 15110 -12503 15140 -12477
rect 15196 -12503 15226 -12477
rect 15282 -12503 15312 -12477
rect 15368 -12503 15398 -12477
rect 15666 -12503 16612 -12477
rect -2918 -12571 -2340 -12545
rect -1538 -12571 -960 -12545
rect -802 -12571 -224 -12545
rect 26 -12571 236 -12545
rect 488 -12571 518 -12545
rect 590 -12571 690 -12545
rect 850 -12571 950 -12545
rect 1015 -12571 1045 -12545
rect 1314 -12571 1524 -12545
rect 1774 -12571 2352 -12545
rect 2602 -12571 2812 -12545
rect 3064 -12571 3094 -12545
rect 3166 -12571 3266 -12545
rect 3426 -12571 3526 -12545
rect 3591 -12571 3621 -12545
rect 3890 -12571 4100 -12545
rect 4350 -12571 4928 -12545
rect 5178 -12571 5388 -12545
rect 5640 -12571 5670 -12545
rect 5742 -12571 5842 -12545
rect 6002 -12571 6102 -12545
rect 6167 -12571 6197 -12545
rect 6466 -12571 6676 -12545
rect 6926 -12571 7504 -12545
rect 7754 -12571 7964 -12545
rect 8216 -12571 8246 -12545
rect 8318 -12571 8418 -12545
rect 8578 -12571 8678 -12545
rect 8743 -12571 8773 -12545
rect 9042 -12571 9252 -12545
rect 9502 -12571 10080 -12545
rect 10422 -12571 10632 -12545
rect 10792 -12571 10822 -12545
rect 10894 -12571 10994 -12545
rect 11154 -12571 11254 -12545
rect 11319 -12571 11349 -12545
rect 11710 -12571 11920 -12545
rect 12633 -12571 12663 -12545
rect 12719 -12571 12749 -12545
rect 12805 -12571 12835 -12545
rect 12891 -12571 12921 -12545
rect 13274 -12571 13484 -12545
rect 13735 -12571 13765 -12545
rect 13821 -12571 13851 -12545
rect 13907 -12571 13937 -12545
rect 13993 -12571 14023 -12545
rect 14079 -12571 14109 -12545
rect 14165 -12571 14195 -12545
rect 14251 -12571 14281 -12545
rect 14337 -12571 14367 -12545
rect 14423 -12571 14453 -12545
rect 14509 -12571 14539 -12545
rect 14595 -12571 14625 -12545
rect 14681 -12571 14711 -12545
rect 14766 -12571 14796 -12545
rect 14852 -12571 14882 -12545
rect 14938 -12571 14968 -12545
rect 15024 -12571 15054 -12545
rect 15110 -12571 15140 -12545
rect 15196 -12571 15226 -12545
rect 15282 -12571 15312 -12545
rect 15368 -12571 15398 -12545
rect 15666 -12571 16612 -12545
rect -2918 -12707 -2340 -12681
rect -1538 -12707 -960 -12681
rect -802 -12707 -224 -12681
rect -2918 -12729 -2646 -12707
rect -2918 -12763 -2902 -12729
rect -2868 -12763 -2799 -12729
rect -2765 -12763 -2696 -12729
rect -2662 -12763 -2646 -12729
rect -1232 -12729 -960 -12707
rect -2918 -12779 -2646 -12763
rect -2604 -12765 -2340 -12749
rect -2604 -12799 -2588 -12765
rect -2554 -12799 -2489 -12765
rect -2455 -12799 -2390 -12765
rect -2356 -12799 -2340 -12765
rect -2604 -12821 -2340 -12799
rect -2918 -12847 -2340 -12821
rect -1538 -12765 -1274 -12749
rect -1538 -12799 -1522 -12765
rect -1488 -12799 -1423 -12765
rect -1389 -12799 -1324 -12765
rect -1290 -12799 -1274 -12765
rect -1232 -12763 -1216 -12729
rect -1182 -12763 -1113 -12729
rect -1079 -12763 -1010 -12729
rect -976 -12763 -960 -12729
rect -496 -12729 -224 -12707
rect 26 -12707 236 -12681
rect 26 -12713 110 -12707
rect -1232 -12779 -960 -12763
rect -802 -12765 -538 -12749
rect -1538 -12821 -1274 -12799
rect -802 -12799 -786 -12765
rect -752 -12799 -687 -12765
rect -653 -12799 -588 -12765
rect -554 -12799 -538 -12765
rect -496 -12763 -480 -12729
rect -446 -12763 -377 -12729
rect -343 -12763 -274 -12729
rect -240 -12763 -224 -12729
rect -496 -12779 -224 -12763
rect -32 -12729 110 -12713
rect 488 -12727 518 -12655
rect -32 -12763 -16 -12729
rect 18 -12763 110 -12729
rect 448 -12739 518 -12727
rect 590 -12729 690 -12701
rect 850 -12729 950 -12701
rect 1015 -12723 1045 -12655
rect 1314 -12707 1524 -12681
rect 1774 -12707 2352 -12681
rect 2602 -12707 2812 -12681
rect 1314 -12713 1398 -12707
rect -32 -12779 110 -12763
rect 152 -12765 294 -12749
rect -802 -12821 -538 -12799
rect 152 -12799 244 -12765
rect 278 -12799 294 -12765
rect 448 -12773 464 -12739
rect 498 -12773 518 -12739
rect 448 -12786 518 -12773
rect 568 -12739 690 -12729
rect 568 -12773 584 -12739
rect 618 -12773 690 -12739
rect 568 -12783 690 -12773
rect 789 -12739 950 -12729
rect 789 -12773 805 -12739
rect 839 -12773 950 -12739
rect 789 -12783 950 -12773
rect 152 -12815 294 -12799
rect 152 -12821 236 -12815
rect 488 -12821 518 -12786
rect -1538 -12847 -960 -12821
rect -802 -12847 -224 -12821
rect 26 -12847 236 -12821
rect 590 -12857 690 -12783
rect 850 -12857 950 -12783
rect 995 -12739 1049 -12723
rect 995 -12773 1005 -12739
rect 1039 -12773 1049 -12739
rect 995 -12789 1049 -12773
rect 1256 -12729 1398 -12713
rect 1256 -12763 1272 -12729
rect 1306 -12763 1398 -12729
rect 1774 -12729 2046 -12707
rect 2602 -12713 2686 -12707
rect 1256 -12779 1398 -12763
rect 1440 -12765 1582 -12749
rect 1015 -12821 1045 -12789
rect 1440 -12799 1532 -12765
rect 1566 -12799 1582 -12765
rect 1774 -12763 1790 -12729
rect 1824 -12763 1893 -12729
rect 1927 -12763 1996 -12729
rect 2030 -12763 2046 -12729
rect 2544 -12729 2686 -12713
rect 3064 -12727 3094 -12655
rect 1774 -12779 2046 -12763
rect 2088 -12765 2352 -12749
rect 1440 -12815 1582 -12799
rect 2088 -12799 2104 -12765
rect 2138 -12799 2203 -12765
rect 2237 -12799 2302 -12765
rect 2336 -12799 2352 -12765
rect 2544 -12763 2560 -12729
rect 2594 -12763 2686 -12729
rect 3024 -12739 3094 -12727
rect 3166 -12729 3266 -12701
rect 3426 -12729 3526 -12701
rect 3591 -12723 3621 -12655
rect 3890 -12707 4100 -12681
rect 4350 -12707 4928 -12681
rect 5178 -12707 5388 -12681
rect 3890 -12713 3974 -12707
rect 2544 -12779 2686 -12763
rect 2728 -12765 2870 -12749
rect 1440 -12821 1524 -12815
rect 2088 -12821 2352 -12799
rect 2728 -12799 2820 -12765
rect 2854 -12799 2870 -12765
rect 3024 -12773 3040 -12739
rect 3074 -12773 3094 -12739
rect 3024 -12786 3094 -12773
rect 3144 -12739 3266 -12729
rect 3144 -12773 3160 -12739
rect 3194 -12773 3266 -12739
rect 3144 -12783 3266 -12773
rect 3365 -12739 3526 -12729
rect 3365 -12773 3381 -12739
rect 3415 -12773 3526 -12739
rect 3365 -12783 3526 -12773
rect 2728 -12815 2870 -12799
rect 2728 -12821 2812 -12815
rect 3064 -12821 3094 -12786
rect 1314 -12847 1524 -12821
rect 1774 -12847 2352 -12821
rect 2602 -12847 2812 -12821
rect 3166 -12857 3266 -12783
rect 3426 -12857 3526 -12783
rect 3571 -12739 3625 -12723
rect 3571 -12773 3581 -12739
rect 3615 -12773 3625 -12739
rect 3571 -12789 3625 -12773
rect 3832 -12729 3974 -12713
rect 3832 -12763 3848 -12729
rect 3882 -12763 3974 -12729
rect 4350 -12729 4622 -12707
rect 5178 -12713 5262 -12707
rect 3832 -12779 3974 -12763
rect 4016 -12765 4158 -12749
rect 3591 -12821 3621 -12789
rect 4016 -12799 4108 -12765
rect 4142 -12799 4158 -12765
rect 4350 -12763 4366 -12729
rect 4400 -12763 4469 -12729
rect 4503 -12763 4572 -12729
rect 4606 -12763 4622 -12729
rect 5120 -12729 5262 -12713
rect 5640 -12727 5670 -12655
rect 4350 -12779 4622 -12763
rect 4664 -12765 4928 -12749
rect 4016 -12815 4158 -12799
rect 4664 -12799 4680 -12765
rect 4714 -12799 4779 -12765
rect 4813 -12799 4878 -12765
rect 4912 -12799 4928 -12765
rect 5120 -12763 5136 -12729
rect 5170 -12763 5262 -12729
rect 5600 -12739 5670 -12727
rect 5742 -12729 5842 -12701
rect 6002 -12729 6102 -12701
rect 6167 -12723 6197 -12655
rect 6466 -12707 6676 -12681
rect 6926 -12707 7504 -12681
rect 7754 -12707 7964 -12681
rect 6466 -12713 6550 -12707
rect 5120 -12779 5262 -12763
rect 5304 -12765 5446 -12749
rect 4016 -12821 4100 -12815
rect 4664 -12821 4928 -12799
rect 5304 -12799 5396 -12765
rect 5430 -12799 5446 -12765
rect 5600 -12773 5616 -12739
rect 5650 -12773 5670 -12739
rect 5600 -12786 5670 -12773
rect 5720 -12739 5842 -12729
rect 5720 -12773 5736 -12739
rect 5770 -12773 5842 -12739
rect 5720 -12783 5842 -12773
rect 5941 -12739 6102 -12729
rect 5941 -12773 5957 -12739
rect 5991 -12773 6102 -12739
rect 5941 -12783 6102 -12773
rect 5304 -12815 5446 -12799
rect 5304 -12821 5388 -12815
rect 5640 -12821 5670 -12786
rect 3890 -12847 4100 -12821
rect 4350 -12847 4928 -12821
rect 5178 -12847 5388 -12821
rect 5742 -12857 5842 -12783
rect 6002 -12857 6102 -12783
rect 6147 -12739 6201 -12723
rect 6147 -12773 6157 -12739
rect 6191 -12773 6201 -12739
rect 6147 -12789 6201 -12773
rect 6408 -12729 6550 -12713
rect 6408 -12763 6424 -12729
rect 6458 -12763 6550 -12729
rect 6926 -12729 7198 -12707
rect 7754 -12713 7838 -12707
rect 6408 -12779 6550 -12763
rect 6592 -12765 6734 -12749
rect 6167 -12821 6197 -12789
rect 6592 -12799 6684 -12765
rect 6718 -12799 6734 -12765
rect 6926 -12763 6942 -12729
rect 6976 -12763 7045 -12729
rect 7079 -12763 7148 -12729
rect 7182 -12763 7198 -12729
rect 7696 -12729 7838 -12713
rect 8216 -12727 8246 -12655
rect 6926 -12779 7198 -12763
rect 7240 -12765 7504 -12749
rect 6592 -12815 6734 -12799
rect 7240 -12799 7256 -12765
rect 7290 -12799 7355 -12765
rect 7389 -12799 7454 -12765
rect 7488 -12799 7504 -12765
rect 7696 -12763 7712 -12729
rect 7746 -12763 7838 -12729
rect 8176 -12739 8246 -12727
rect 8318 -12729 8418 -12701
rect 8578 -12729 8678 -12701
rect 8743 -12723 8773 -12655
rect 9042 -12707 9252 -12681
rect 9502 -12707 10080 -12681
rect 10422 -12707 10632 -12681
rect 9042 -12713 9126 -12707
rect 7696 -12779 7838 -12763
rect 7880 -12765 8022 -12749
rect 6592 -12821 6676 -12815
rect 7240 -12821 7504 -12799
rect 7880 -12799 7972 -12765
rect 8006 -12799 8022 -12765
rect 8176 -12773 8192 -12739
rect 8226 -12773 8246 -12739
rect 8176 -12786 8246 -12773
rect 8296 -12739 8418 -12729
rect 8296 -12773 8312 -12739
rect 8346 -12773 8418 -12739
rect 8296 -12783 8418 -12773
rect 8517 -12739 8678 -12729
rect 8517 -12773 8533 -12739
rect 8567 -12773 8678 -12739
rect 8517 -12783 8678 -12773
rect 7880 -12815 8022 -12799
rect 7880 -12821 7964 -12815
rect 8216 -12821 8246 -12786
rect 6466 -12847 6676 -12821
rect 6926 -12847 7504 -12821
rect 7754 -12847 7964 -12821
rect 8318 -12857 8418 -12783
rect 8578 -12857 8678 -12783
rect 8723 -12739 8777 -12723
rect 8723 -12773 8733 -12739
rect 8767 -12773 8777 -12739
rect 8723 -12789 8777 -12773
rect 8984 -12729 9126 -12713
rect 8984 -12763 9000 -12729
rect 9034 -12763 9126 -12729
rect 9502 -12729 9774 -12707
rect 10422 -12713 10506 -12707
rect 8984 -12779 9126 -12763
rect 9168 -12765 9310 -12749
rect 8743 -12821 8773 -12789
rect 9168 -12799 9260 -12765
rect 9294 -12799 9310 -12765
rect 9502 -12763 9518 -12729
rect 9552 -12763 9621 -12729
rect 9655 -12763 9724 -12729
rect 9758 -12763 9774 -12729
rect 10364 -12729 10506 -12713
rect 10792 -12727 10822 -12655
rect 9502 -12779 9774 -12763
rect 9816 -12765 10080 -12749
rect 9168 -12815 9310 -12799
rect 9816 -12799 9832 -12765
rect 9866 -12799 9931 -12765
rect 9965 -12799 10030 -12765
rect 10064 -12799 10080 -12765
rect 10364 -12763 10380 -12729
rect 10414 -12763 10506 -12729
rect 10752 -12739 10822 -12727
rect 10894 -12729 10994 -12701
rect 11154 -12729 11254 -12701
rect 11319 -12723 11349 -12655
rect 11710 -12707 11920 -12681
rect 11710 -12713 11794 -12707
rect 10364 -12779 10506 -12763
rect 10548 -12765 10690 -12749
rect 9168 -12821 9252 -12815
rect 9816 -12821 10080 -12799
rect 10548 -12799 10640 -12765
rect 10674 -12799 10690 -12765
rect 10752 -12773 10768 -12739
rect 10802 -12773 10822 -12739
rect 10752 -12786 10822 -12773
rect 10872 -12739 10994 -12729
rect 10872 -12773 10888 -12739
rect 10922 -12773 10994 -12739
rect 10872 -12783 10994 -12773
rect 11093 -12739 11254 -12729
rect 11093 -12773 11109 -12739
rect 11143 -12773 11254 -12739
rect 11093 -12783 11254 -12773
rect 10548 -12815 10690 -12799
rect 10548 -12821 10632 -12815
rect 10792 -12821 10822 -12786
rect 9042 -12847 9252 -12821
rect 9502 -12847 10080 -12821
rect 10422 -12847 10632 -12821
rect 10894 -12857 10994 -12783
rect 11154 -12857 11254 -12783
rect 11299 -12739 11353 -12723
rect 11299 -12773 11309 -12739
rect 11343 -12773 11353 -12739
rect 11299 -12789 11353 -12773
rect 11652 -12729 11794 -12713
rect 12633 -12729 12663 -12655
rect 12719 -12729 12749 -12655
rect 12805 -12729 12835 -12655
rect 12891 -12729 12921 -12655
rect 13274 -12707 13484 -12681
rect 13735 -12704 13765 -12655
rect 13821 -12704 13851 -12655
rect 13907 -12704 13937 -12655
rect 13993 -12704 14023 -12655
rect 13400 -12713 13484 -12707
rect 13400 -12729 13542 -12713
rect 11652 -12763 11668 -12729
rect 11702 -12763 11794 -12729
rect 12547 -12739 13007 -12729
rect 11652 -12779 11794 -12763
rect 11836 -12765 11978 -12749
rect 11319 -12821 11349 -12789
rect 11836 -12799 11928 -12765
rect 11962 -12799 11978 -12765
rect 11836 -12815 11978 -12799
rect 12547 -12773 12574 -12739
rect 12608 -12773 12642 -12739
rect 12676 -12773 12710 -12739
rect 12744 -12773 12778 -12739
rect 12812 -12773 12846 -12739
rect 12880 -12773 12914 -12739
rect 12948 -12773 13007 -12739
rect 12547 -12783 13007 -12773
rect 11836 -12821 11920 -12815
rect 12547 -12821 12577 -12783
rect 12633 -12821 12663 -12783
rect 12719 -12821 12749 -12783
rect 12805 -12821 12835 -12783
rect 12891 -12821 12921 -12783
rect 12977 -12821 13007 -12783
rect 13216 -12765 13358 -12749
rect 13216 -12799 13232 -12765
rect 13266 -12799 13358 -12765
rect 13400 -12763 13492 -12729
rect 13526 -12763 13542 -12729
rect 13400 -12779 13542 -12763
rect 13676 -12739 14023 -12704
rect 13676 -12773 13692 -12739
rect 13726 -12773 14023 -12739
rect 13216 -12815 13358 -12799
rect 13676 -12806 14023 -12773
rect 13274 -12821 13358 -12815
rect 13735 -12821 13765 -12806
rect 13821 -12821 13851 -12806
rect 13907 -12821 13937 -12806
rect 13993 -12821 14023 -12806
rect 14079 -12714 14109 -12655
rect 14165 -12714 14195 -12655
rect 14251 -12714 14281 -12655
rect 14337 -12714 14367 -12655
rect 14423 -12714 14453 -12655
rect 14509 -12714 14539 -12655
rect 14595 -12714 14625 -12655
rect 14681 -12714 14711 -12655
rect 14766 -12714 14796 -12655
rect 14852 -12714 14882 -12655
rect 14938 -12714 14968 -12655
rect 15024 -12714 15054 -12655
rect 15110 -12714 15140 -12655
rect 15196 -12714 15226 -12655
rect 15282 -12714 15312 -12655
rect 15368 -12714 15398 -12655
rect 15666 -12707 16612 -12681
rect 14079 -12739 15398 -12714
rect 14079 -12773 14119 -12739
rect 14153 -12773 14187 -12739
rect 14221 -12773 14255 -12739
rect 14289 -12773 14323 -12739
rect 14357 -12773 14391 -12739
rect 14425 -12773 14459 -12739
rect 14493 -12773 14527 -12739
rect 14561 -12773 14595 -12739
rect 14629 -12773 14663 -12739
rect 14697 -12773 14731 -12739
rect 14765 -12773 14799 -12739
rect 14833 -12773 14867 -12739
rect 14901 -12773 14935 -12739
rect 14969 -12773 15003 -12739
rect 15037 -12773 15071 -12739
rect 15105 -12773 15139 -12739
rect 15173 -12773 15398 -12739
rect 16158 -12729 16612 -12707
rect 14079 -12789 15398 -12773
rect 14079 -12821 14109 -12789
rect 14165 -12821 14195 -12789
rect 14251 -12821 14281 -12789
rect 14337 -12821 14367 -12789
rect 14423 -12821 14453 -12789
rect 14509 -12821 14539 -12789
rect 14595 -12821 14625 -12789
rect 14681 -12821 14711 -12789
rect 14766 -12821 14796 -12789
rect 14852 -12821 14882 -12789
rect 14938 -12821 14968 -12789
rect 15024 -12821 15054 -12789
rect 15110 -12821 15140 -12789
rect 15196 -12821 15226 -12789
rect 15282 -12821 15312 -12789
rect 15368 -12821 15398 -12789
rect 15666 -12765 16116 -12749
rect 15666 -12799 15682 -12765
rect 15716 -12799 15810 -12765
rect 15844 -12799 15938 -12765
rect 15972 -12799 16066 -12765
rect 16100 -12799 16116 -12765
rect 16158 -12763 16174 -12729
rect 16208 -12763 16302 -12729
rect 16336 -12763 16430 -12729
rect 16464 -12763 16558 -12729
rect 16592 -12763 16612 -12729
rect 16158 -12779 16612 -12763
rect 15666 -12821 16116 -12799
rect 11710 -12847 11920 -12821
rect 13274 -12847 13484 -12821
rect 15666 -12847 16612 -12821
rect -2918 -13047 -2340 -13021
rect -1538 -13047 -960 -13021
rect -802 -13047 -224 -13021
rect 26 -13047 236 -13021
rect 488 -13047 518 -13021
rect 590 -13047 690 -13021
rect 850 -13047 950 -13021
rect 1015 -13047 1045 -13021
rect 1314 -13047 1524 -13021
rect 1774 -13047 2352 -13021
rect 2602 -13047 2812 -13021
rect 3064 -13047 3094 -13021
rect 3166 -13047 3266 -13021
rect 3426 -13047 3526 -13021
rect 3591 -13047 3621 -13021
rect 3890 -13047 4100 -13021
rect 4350 -13047 4928 -13021
rect 5178 -13047 5388 -13021
rect 5640 -13047 5670 -13021
rect 5742 -13047 5842 -13021
rect 6002 -13047 6102 -13021
rect 6167 -13047 6197 -13021
rect 6466 -13047 6676 -13021
rect 6926 -13047 7504 -13021
rect 7754 -13047 7964 -13021
rect 8216 -13047 8246 -13021
rect 8318 -13047 8418 -13021
rect 8578 -13047 8678 -13021
rect 8743 -13047 8773 -13021
rect 9042 -13047 9252 -13021
rect 9502 -13047 10080 -13021
rect 10422 -13047 10632 -13021
rect 10792 -13047 10822 -13021
rect 10894 -13047 10994 -13021
rect 11154 -13047 11254 -13021
rect 11319 -13047 11349 -13021
rect 11710 -13047 11920 -13021
rect 12547 -13047 12577 -13021
rect 12633 -13047 12663 -13021
rect 12719 -13047 12749 -13021
rect 12805 -13047 12835 -13021
rect 12891 -13047 12921 -13021
rect 12977 -13047 13007 -13021
rect 13274 -13047 13484 -13021
rect 13735 -13047 13765 -13021
rect 13821 -13047 13851 -13021
rect 13907 -13047 13937 -13021
rect 13993 -13047 14023 -13021
rect 14079 -13047 14109 -13021
rect 14165 -13047 14195 -13021
rect 14251 -13047 14281 -13021
rect 14337 -13047 14367 -13021
rect 14423 -13047 14453 -13021
rect 14509 -13047 14539 -13021
rect 14595 -13047 14625 -13021
rect 14681 -13047 14711 -13021
rect 14766 -13047 14796 -13021
rect 14852 -13047 14882 -13021
rect 14938 -13047 14968 -13021
rect 15024 -13047 15054 -13021
rect 15110 -13047 15140 -13021
rect 15196 -13047 15226 -13021
rect 15282 -13047 15312 -13021
rect 15368 -13047 15398 -13021
rect 15666 -13047 16612 -13021
rect -2918 -13115 -2340 -13089
rect -1538 -13115 -960 -13089
rect -802 -13115 -224 -13089
rect 26 -13115 236 -13089
rect 505 -13115 535 -13089
rect 600 -13115 700 -13089
rect 860 -13115 960 -13089
rect 1032 -13115 1062 -13089
rect 1314 -13115 1524 -13089
rect 1774 -13115 2352 -13089
rect 2602 -13115 2812 -13089
rect 3081 -13115 3111 -13089
rect 3176 -13115 3276 -13089
rect 3436 -13115 3536 -13089
rect 3608 -13115 3638 -13089
rect 3890 -13115 4100 -13089
rect 4350 -13115 4928 -13089
rect 5178 -13115 5388 -13089
rect 5657 -13115 5687 -13089
rect 5752 -13115 5852 -13089
rect 6012 -13115 6112 -13089
rect 6184 -13115 6214 -13089
rect 6466 -13115 6676 -13089
rect 6926 -13115 7504 -13089
rect 7754 -13115 7964 -13089
rect 8233 -13115 8263 -13089
rect 8328 -13115 8428 -13089
rect 8588 -13115 8688 -13089
rect 8760 -13115 8790 -13089
rect 9042 -13115 9252 -13089
rect 9502 -13115 10080 -13089
rect 10422 -13115 10632 -13089
rect 10809 -13115 10839 -13089
rect 10904 -13115 11004 -13089
rect 11164 -13115 11264 -13089
rect 11336 -13115 11366 -13089
rect 11710 -13115 11920 -13089
rect 13735 -13115 13765 -13089
rect 13821 -13115 13851 -13089
rect 13907 -13115 13937 -13089
rect 13993 -13115 14023 -13089
rect 14079 -13115 14109 -13089
rect 14165 -13115 14195 -13089
rect 14251 -13115 14281 -13089
rect 14337 -13115 14367 -13089
rect 14423 -13115 14453 -13089
rect 14509 -13115 14539 -13089
rect 14595 -13115 14625 -13089
rect 14681 -13115 14711 -13089
rect 14766 -13115 14796 -13089
rect 14852 -13115 14882 -13089
rect 14938 -13115 14968 -13089
rect 15024 -13115 15054 -13089
rect 15110 -13115 15140 -13089
rect 15196 -13115 15226 -13089
rect 15282 -13115 15312 -13089
rect 15368 -13115 15398 -13089
rect 15666 -13115 16612 -13089
rect -2918 -13315 -2340 -13289
rect -1538 -13315 -960 -13289
rect -802 -13315 -224 -13289
rect 26 -13315 236 -13289
rect -2918 -13337 -2654 -13315
rect -2918 -13371 -2902 -13337
rect -2868 -13371 -2803 -13337
rect -2769 -13371 -2704 -13337
rect -2670 -13371 -2654 -13337
rect -1224 -13337 -960 -13315
rect -2918 -13387 -2654 -13371
rect -2612 -13373 -2340 -13357
rect -2612 -13407 -2596 -13373
rect -2562 -13407 -2493 -13373
rect -2459 -13407 -2390 -13373
rect -2356 -13407 -2340 -13373
rect -2612 -13429 -2340 -13407
rect -2918 -13455 -2340 -13429
rect -1538 -13373 -1266 -13357
rect -1538 -13407 -1522 -13373
rect -1488 -13407 -1419 -13373
rect -1385 -13407 -1316 -13373
rect -1282 -13407 -1266 -13373
rect -1224 -13371 -1208 -13337
rect -1174 -13371 -1109 -13337
rect -1075 -13371 -1010 -13337
rect -976 -13371 -960 -13337
rect -488 -13337 -224 -13315
rect -1224 -13387 -960 -13371
rect -802 -13373 -530 -13357
rect -1538 -13429 -1266 -13407
rect -802 -13407 -786 -13373
rect -752 -13407 -683 -13373
rect -649 -13407 -580 -13373
rect -546 -13407 -530 -13373
rect -488 -13371 -472 -13337
rect -438 -13371 -373 -13337
rect -339 -13371 -274 -13337
rect -240 -13371 -224 -13337
rect 152 -13321 236 -13315
rect 152 -13337 294 -13321
rect -488 -13387 -224 -13371
rect -32 -13373 110 -13357
rect -802 -13429 -530 -13407
rect -32 -13407 -16 -13373
rect 18 -13407 110 -13373
rect 152 -13371 244 -13337
rect 278 -13371 294 -13337
rect 505 -13347 535 -13315
rect 152 -13387 294 -13371
rect 501 -13363 555 -13347
rect -32 -13423 110 -13407
rect 501 -13397 511 -13363
rect 545 -13397 555 -13363
rect 501 -13413 555 -13397
rect 600 -13353 700 -13279
rect 860 -13353 960 -13279
rect 1314 -13315 1524 -13289
rect 1032 -13350 1062 -13315
rect 1440 -13321 1524 -13315
rect 1774 -13315 2352 -13289
rect 2602 -13315 2812 -13289
rect 1440 -13337 1582 -13321
rect 600 -13363 761 -13353
rect 600 -13397 711 -13363
rect 745 -13397 761 -13363
rect 600 -13407 761 -13397
rect 860 -13363 982 -13353
rect 860 -13397 932 -13363
rect 966 -13397 982 -13363
rect 860 -13407 982 -13397
rect 1032 -13363 1102 -13350
rect 1032 -13397 1052 -13363
rect 1086 -13397 1102 -13363
rect 26 -13429 110 -13423
rect -1538 -13455 -960 -13429
rect -802 -13455 -224 -13429
rect 26 -13455 236 -13429
rect 505 -13481 535 -13413
rect 600 -13435 700 -13407
rect 860 -13435 960 -13407
rect 1032 -13409 1102 -13397
rect 1256 -13373 1398 -13357
rect 1256 -13407 1272 -13373
rect 1306 -13407 1398 -13373
rect 1440 -13371 1532 -13337
rect 1566 -13371 1582 -13337
rect 1440 -13387 1582 -13371
rect 1774 -13337 2038 -13315
rect 1774 -13371 1790 -13337
rect 1824 -13371 1889 -13337
rect 1923 -13371 1988 -13337
rect 2022 -13371 2038 -13337
rect 2728 -13321 2812 -13315
rect 2728 -13337 2870 -13321
rect 1774 -13387 2038 -13371
rect 2080 -13373 2352 -13357
rect 1032 -13481 1062 -13409
rect 1256 -13423 1398 -13407
rect 1314 -13429 1398 -13423
rect 2080 -13407 2096 -13373
rect 2130 -13407 2199 -13373
rect 2233 -13407 2302 -13373
rect 2336 -13407 2352 -13373
rect 2080 -13429 2352 -13407
rect 2544 -13373 2686 -13357
rect 2544 -13407 2560 -13373
rect 2594 -13407 2686 -13373
rect 2728 -13371 2820 -13337
rect 2854 -13371 2870 -13337
rect 3081 -13347 3111 -13315
rect 2728 -13387 2870 -13371
rect 3077 -13363 3131 -13347
rect 2544 -13423 2686 -13407
rect 3077 -13397 3087 -13363
rect 3121 -13397 3131 -13363
rect 3077 -13413 3131 -13397
rect 3176 -13353 3276 -13279
rect 3436 -13353 3536 -13279
rect 3890 -13315 4100 -13289
rect 3608 -13350 3638 -13315
rect 4016 -13321 4100 -13315
rect 4350 -13315 4928 -13289
rect 5178 -13315 5388 -13289
rect 4016 -13337 4158 -13321
rect 3176 -13363 3337 -13353
rect 3176 -13397 3287 -13363
rect 3321 -13397 3337 -13363
rect 3176 -13407 3337 -13397
rect 3436 -13363 3558 -13353
rect 3436 -13397 3508 -13363
rect 3542 -13397 3558 -13363
rect 3436 -13407 3558 -13397
rect 3608 -13363 3678 -13350
rect 3608 -13397 3628 -13363
rect 3662 -13397 3678 -13363
rect 1314 -13455 1524 -13429
rect 1774 -13455 2352 -13429
rect 2602 -13429 2686 -13423
rect 2602 -13455 2812 -13429
rect 3081 -13481 3111 -13413
rect 3176 -13435 3276 -13407
rect 3436 -13435 3536 -13407
rect 3608 -13409 3678 -13397
rect 3832 -13373 3974 -13357
rect 3832 -13407 3848 -13373
rect 3882 -13407 3974 -13373
rect 4016 -13371 4108 -13337
rect 4142 -13371 4158 -13337
rect 4016 -13387 4158 -13371
rect 4350 -13337 4614 -13315
rect 4350 -13371 4366 -13337
rect 4400 -13371 4465 -13337
rect 4499 -13371 4564 -13337
rect 4598 -13371 4614 -13337
rect 5304 -13321 5388 -13315
rect 5304 -13337 5446 -13321
rect 4350 -13387 4614 -13371
rect 4656 -13373 4928 -13357
rect 3608 -13481 3638 -13409
rect 3832 -13423 3974 -13407
rect 3890 -13429 3974 -13423
rect 4656 -13407 4672 -13373
rect 4706 -13407 4775 -13373
rect 4809 -13407 4878 -13373
rect 4912 -13407 4928 -13373
rect 4656 -13429 4928 -13407
rect 5120 -13373 5262 -13357
rect 5120 -13407 5136 -13373
rect 5170 -13407 5262 -13373
rect 5304 -13371 5396 -13337
rect 5430 -13371 5446 -13337
rect 5657 -13347 5687 -13315
rect 5304 -13387 5446 -13371
rect 5653 -13363 5707 -13347
rect 5120 -13423 5262 -13407
rect 5653 -13397 5663 -13363
rect 5697 -13397 5707 -13363
rect 5653 -13413 5707 -13397
rect 5752 -13353 5852 -13279
rect 6012 -13353 6112 -13279
rect 6466 -13315 6676 -13289
rect 6184 -13350 6214 -13315
rect 6592 -13321 6676 -13315
rect 6926 -13315 7504 -13289
rect 7754 -13315 7964 -13289
rect 6592 -13337 6734 -13321
rect 5752 -13363 5913 -13353
rect 5752 -13397 5863 -13363
rect 5897 -13397 5913 -13363
rect 5752 -13407 5913 -13397
rect 6012 -13363 6134 -13353
rect 6012 -13397 6084 -13363
rect 6118 -13397 6134 -13363
rect 6012 -13407 6134 -13397
rect 6184 -13363 6254 -13350
rect 6184 -13397 6204 -13363
rect 6238 -13397 6254 -13363
rect 3890 -13455 4100 -13429
rect 4350 -13455 4928 -13429
rect 5178 -13429 5262 -13423
rect 5178 -13455 5388 -13429
rect 5657 -13481 5687 -13413
rect 5752 -13435 5852 -13407
rect 6012 -13435 6112 -13407
rect 6184 -13409 6254 -13397
rect 6408 -13373 6550 -13357
rect 6408 -13407 6424 -13373
rect 6458 -13407 6550 -13373
rect 6592 -13371 6684 -13337
rect 6718 -13371 6734 -13337
rect 6592 -13387 6734 -13371
rect 6926 -13337 7190 -13315
rect 6926 -13371 6942 -13337
rect 6976 -13371 7041 -13337
rect 7075 -13371 7140 -13337
rect 7174 -13371 7190 -13337
rect 7880 -13321 7964 -13315
rect 7880 -13337 8022 -13321
rect 6926 -13387 7190 -13371
rect 7232 -13373 7504 -13357
rect 6184 -13481 6214 -13409
rect 6408 -13423 6550 -13407
rect 6466 -13429 6550 -13423
rect 7232 -13407 7248 -13373
rect 7282 -13407 7351 -13373
rect 7385 -13407 7454 -13373
rect 7488 -13407 7504 -13373
rect 7232 -13429 7504 -13407
rect 7696 -13373 7838 -13357
rect 7696 -13407 7712 -13373
rect 7746 -13407 7838 -13373
rect 7880 -13371 7972 -13337
rect 8006 -13371 8022 -13337
rect 8233 -13347 8263 -13315
rect 7880 -13387 8022 -13371
rect 8229 -13363 8283 -13347
rect 7696 -13423 7838 -13407
rect 8229 -13397 8239 -13363
rect 8273 -13397 8283 -13363
rect 8229 -13413 8283 -13397
rect 8328 -13353 8428 -13279
rect 8588 -13353 8688 -13279
rect 9042 -13315 9252 -13289
rect 8760 -13350 8790 -13315
rect 9168 -13321 9252 -13315
rect 9502 -13315 10080 -13289
rect 10422 -13315 10632 -13289
rect 9168 -13337 9310 -13321
rect 8328 -13363 8489 -13353
rect 8328 -13397 8439 -13363
rect 8473 -13397 8489 -13363
rect 8328 -13407 8489 -13397
rect 8588 -13363 8710 -13353
rect 8588 -13397 8660 -13363
rect 8694 -13397 8710 -13363
rect 8588 -13407 8710 -13397
rect 8760 -13363 8830 -13350
rect 8760 -13397 8780 -13363
rect 8814 -13397 8830 -13363
rect 6466 -13455 6676 -13429
rect 6926 -13455 7504 -13429
rect 7754 -13429 7838 -13423
rect 7754 -13455 7964 -13429
rect 8233 -13481 8263 -13413
rect 8328 -13435 8428 -13407
rect 8588 -13435 8688 -13407
rect 8760 -13409 8830 -13397
rect 8984 -13373 9126 -13357
rect 8984 -13407 9000 -13373
rect 9034 -13407 9126 -13373
rect 9168 -13371 9260 -13337
rect 9294 -13371 9310 -13337
rect 9168 -13387 9310 -13371
rect 9502 -13337 9766 -13315
rect 9502 -13371 9518 -13337
rect 9552 -13371 9617 -13337
rect 9651 -13371 9716 -13337
rect 9750 -13371 9766 -13337
rect 10548 -13321 10632 -13315
rect 10548 -13337 10690 -13321
rect 9502 -13387 9766 -13371
rect 9808 -13373 10080 -13357
rect 8760 -13481 8790 -13409
rect 8984 -13423 9126 -13407
rect 9042 -13429 9126 -13423
rect 9808 -13407 9824 -13373
rect 9858 -13407 9927 -13373
rect 9961 -13407 10030 -13373
rect 10064 -13407 10080 -13373
rect 9808 -13429 10080 -13407
rect 10364 -13373 10506 -13357
rect 10364 -13407 10380 -13373
rect 10414 -13407 10506 -13373
rect 10548 -13371 10640 -13337
rect 10674 -13371 10690 -13337
rect 10809 -13347 10839 -13315
rect 10548 -13387 10690 -13371
rect 10805 -13363 10859 -13347
rect 10364 -13423 10506 -13407
rect 10805 -13397 10815 -13363
rect 10849 -13397 10859 -13363
rect 10805 -13413 10859 -13397
rect 10904 -13353 11004 -13279
rect 11164 -13353 11264 -13279
rect 11710 -13315 11920 -13289
rect 15666 -13315 16612 -13289
rect 11336 -13350 11366 -13315
rect 11836 -13321 11920 -13315
rect 11836 -13337 11978 -13321
rect 13735 -13330 13765 -13315
rect 13821 -13330 13851 -13315
rect 13907 -13330 13937 -13315
rect 13993 -13330 14023 -13315
rect 10904 -13363 11065 -13353
rect 10904 -13397 11015 -13363
rect 11049 -13397 11065 -13363
rect 10904 -13407 11065 -13397
rect 11164 -13363 11286 -13353
rect 11164 -13397 11236 -13363
rect 11270 -13397 11286 -13363
rect 11164 -13407 11286 -13397
rect 11336 -13363 11406 -13350
rect 11336 -13397 11356 -13363
rect 11390 -13397 11406 -13363
rect 9042 -13455 9252 -13429
rect 9502 -13455 10080 -13429
rect 10422 -13429 10506 -13423
rect 10422 -13455 10632 -13429
rect 10809 -13481 10839 -13413
rect 10904 -13435 11004 -13407
rect 11164 -13435 11264 -13407
rect 11336 -13409 11406 -13397
rect 11652 -13373 11794 -13357
rect 11652 -13407 11668 -13373
rect 11702 -13407 11794 -13373
rect 11836 -13371 11928 -13337
rect 11962 -13371 11978 -13337
rect 11836 -13387 11978 -13371
rect 13676 -13363 14023 -13330
rect 11336 -13481 11366 -13409
rect 11652 -13423 11794 -13407
rect 11710 -13429 11794 -13423
rect 13676 -13397 13692 -13363
rect 13726 -13397 14023 -13363
rect 11710 -13455 11920 -13429
rect 13676 -13432 14023 -13397
rect 13735 -13481 13765 -13432
rect 13821 -13481 13851 -13432
rect 13907 -13481 13937 -13432
rect 13993 -13481 14023 -13432
rect 14079 -13347 14109 -13315
rect 14165 -13347 14195 -13315
rect 14251 -13347 14281 -13315
rect 14337 -13347 14367 -13315
rect 14423 -13347 14453 -13315
rect 14509 -13347 14539 -13315
rect 14595 -13347 14625 -13315
rect 14681 -13347 14711 -13315
rect 14766 -13347 14796 -13315
rect 14852 -13347 14882 -13315
rect 14938 -13347 14968 -13315
rect 15024 -13347 15054 -13315
rect 15110 -13347 15140 -13315
rect 15196 -13347 15226 -13315
rect 15282 -13347 15312 -13315
rect 15368 -13347 15398 -13315
rect 14079 -13363 15398 -13347
rect 16162 -13337 16612 -13315
rect 14079 -13397 14119 -13363
rect 14153 -13397 14187 -13363
rect 14221 -13397 14255 -13363
rect 14289 -13397 14323 -13363
rect 14357 -13397 14391 -13363
rect 14425 -13397 14459 -13363
rect 14493 -13397 14527 -13363
rect 14561 -13397 14595 -13363
rect 14629 -13397 14663 -13363
rect 14697 -13397 14731 -13363
rect 14765 -13397 14799 -13363
rect 14833 -13397 14867 -13363
rect 14901 -13397 14935 -13363
rect 14969 -13397 15003 -13363
rect 15037 -13397 15071 -13363
rect 15105 -13397 15139 -13363
rect 15173 -13397 15398 -13363
rect 14079 -13422 15398 -13397
rect 14079 -13481 14109 -13422
rect 14165 -13481 14195 -13422
rect 14251 -13481 14281 -13422
rect 14337 -13481 14367 -13422
rect 14423 -13481 14453 -13422
rect 14509 -13481 14539 -13422
rect 14595 -13481 14625 -13422
rect 14681 -13481 14711 -13422
rect 14766 -13481 14796 -13422
rect 14852 -13481 14882 -13422
rect 14938 -13481 14968 -13422
rect 15024 -13481 15054 -13422
rect 15110 -13481 15140 -13422
rect 15196 -13481 15226 -13422
rect 15282 -13481 15312 -13422
rect 15368 -13481 15398 -13422
rect 15666 -13373 16120 -13357
rect 15666 -13407 15686 -13373
rect 15720 -13407 15814 -13373
rect 15848 -13407 15942 -13373
rect 15976 -13407 16070 -13373
rect 16104 -13407 16120 -13373
rect 16162 -13371 16178 -13337
rect 16212 -13371 16306 -13337
rect 16340 -13371 16434 -13337
rect 16468 -13371 16562 -13337
rect 16596 -13371 16612 -13337
rect 16162 -13387 16612 -13371
rect 15666 -13429 16120 -13407
rect 15666 -13455 16612 -13429
rect -2918 -13591 -2340 -13565
rect -1538 -13591 -960 -13565
rect -802 -13591 -224 -13565
rect 26 -13591 236 -13565
rect 505 -13591 535 -13565
rect 600 -13591 700 -13565
rect 860 -13591 960 -13565
rect 1032 -13591 1062 -13565
rect 1314 -13591 1524 -13565
rect 1774 -13591 2352 -13565
rect 2602 -13591 2812 -13565
rect 3081 -13591 3111 -13565
rect 3176 -13591 3276 -13565
rect 3436 -13591 3536 -13565
rect 3608 -13591 3638 -13565
rect 3890 -13591 4100 -13565
rect 4350 -13591 4928 -13565
rect 5178 -13591 5388 -13565
rect 5657 -13591 5687 -13565
rect 5752 -13591 5852 -13565
rect 6012 -13591 6112 -13565
rect 6184 -13591 6214 -13565
rect 6466 -13591 6676 -13565
rect 6926 -13591 7504 -13565
rect 7754 -13591 7964 -13565
rect 8233 -13591 8263 -13565
rect 8328 -13591 8428 -13565
rect 8588 -13591 8688 -13565
rect 8760 -13591 8790 -13565
rect 9042 -13591 9252 -13565
rect 9502 -13591 10080 -13565
rect 10422 -13591 10632 -13565
rect 10809 -13591 10839 -13565
rect 10904 -13591 11004 -13565
rect 11164 -13591 11264 -13565
rect 11336 -13591 11366 -13565
rect 11710 -13591 11920 -13565
rect 13735 -13591 13765 -13565
rect 13821 -13591 13851 -13565
rect 13907 -13591 13937 -13565
rect 13993 -13591 14023 -13565
rect 14079 -13591 14109 -13565
rect 14165 -13591 14195 -13565
rect 14251 -13591 14281 -13565
rect 14337 -13591 14367 -13565
rect 14423 -13591 14453 -13565
rect 14509 -13591 14539 -13565
rect 14595 -13591 14625 -13565
rect 14681 -13591 14711 -13565
rect 14766 -13591 14796 -13565
rect 14852 -13591 14882 -13565
rect 14938 -13591 14968 -13565
rect 15024 -13591 15054 -13565
rect 15110 -13591 15140 -13565
rect 15196 -13591 15226 -13565
rect 15282 -13591 15312 -13565
rect 15368 -13591 15398 -13565
rect 15666 -13591 16612 -13565
rect -2918 -13659 -2340 -13633
rect -1354 -13659 -1144 -13633
rect -890 -13659 -860 -13633
rect -806 -13659 -776 -13633
rect -526 -13659 -316 -13633
rect 29 -13659 59 -13633
rect 115 -13659 145 -13633
rect 201 -13659 231 -13633
rect 287 -13659 317 -13633
rect 670 -13659 880 -13633
rect 1213 -13659 1243 -13633
rect 1498 -13659 1708 -13633
rect 1958 -13659 2168 -13633
rect 2420 -13659 2450 -13633
rect 2522 -13659 2622 -13633
rect 2782 -13659 2882 -13633
rect 2947 -13659 2977 -13633
rect 3246 -13659 3456 -13633
rect 4442 -13659 5388 -13633
rect 6466 -13659 6676 -13633
rect 6928 -13659 6958 -13633
rect 7030 -13659 7130 -13633
rect 7290 -13659 7390 -13633
rect 7455 -13659 7485 -13633
rect 7754 -13659 7964 -13633
rect 8216 -13659 8246 -13633
rect 8318 -13659 8418 -13633
rect 8578 -13659 8678 -13633
rect 8743 -13659 8773 -13633
rect 9042 -13659 9252 -13633
rect 9504 -13659 9534 -13633
rect 9606 -13659 9706 -13633
rect 9866 -13659 9966 -13633
rect 10031 -13659 10061 -13633
rect 10330 -13659 10540 -13633
rect 10790 -13659 10820 -13633
rect 10874 -13659 10904 -13633
rect 10958 -13659 10988 -13633
rect 11042 -13659 11072 -13633
rect 11126 -13659 11156 -13633
rect 11210 -13659 11240 -13633
rect 11294 -13659 11324 -13633
rect 11378 -13659 11408 -13633
rect 11710 -13659 11920 -13633
rect 13642 -13659 14588 -13633
rect 14838 -13659 15784 -13633
rect 16034 -13659 16612 -13633
rect -2918 -13795 -2340 -13769
rect -1354 -13795 -1144 -13769
rect -2918 -13817 -2646 -13795
rect -2918 -13851 -2902 -13817
rect -2868 -13851 -2799 -13817
rect -2765 -13851 -2696 -13817
rect -2662 -13851 -2646 -13817
rect -1228 -13801 -1144 -13795
rect -1228 -13817 -1086 -13801
rect -890 -13811 -860 -13789
rect -2918 -13867 -2646 -13851
rect -2604 -13853 -2340 -13837
rect -2604 -13887 -2588 -13853
rect -2554 -13887 -2489 -13853
rect -2455 -13887 -2390 -13853
rect -2356 -13887 -2340 -13853
rect -2604 -13909 -2340 -13887
rect -1412 -13853 -1270 -13837
rect -1412 -13887 -1396 -13853
rect -1362 -13887 -1270 -13853
rect -1228 -13851 -1136 -13817
rect -1102 -13851 -1086 -13817
rect -1228 -13867 -1086 -13851
rect -952 -13827 -860 -13811
rect -952 -13861 -937 -13827
rect -903 -13861 -860 -13827
rect -952 -13877 -860 -13861
rect -1412 -13903 -1270 -13887
rect -2918 -13935 -2340 -13909
rect -1354 -13909 -1270 -13903
rect -890 -13909 -860 -13877
rect -806 -13811 -776 -13789
rect -526 -13795 -316 -13769
rect -400 -13801 -316 -13795
rect -806 -13827 -718 -13811
rect -806 -13861 -769 -13827
rect -735 -13861 -718 -13827
rect -400 -13817 -258 -13801
rect 29 -13817 59 -13743
rect 115 -13817 145 -13743
rect 201 -13817 231 -13743
rect 287 -13817 317 -13743
rect 670 -13795 880 -13769
rect 796 -13801 880 -13795
rect 796 -13817 938 -13801
rect 1213 -13807 1243 -13743
rect 1498 -13795 1708 -13769
rect 1958 -13795 2168 -13769
rect 1129 -13811 1243 -13807
rect -806 -13877 -718 -13861
rect -584 -13853 -442 -13837
rect -806 -13909 -776 -13877
rect -584 -13887 -568 -13853
rect -534 -13887 -442 -13853
rect -400 -13851 -308 -13817
rect -274 -13851 -258 -13817
rect -400 -13867 -258 -13851
rect -57 -13827 403 -13817
rect -57 -13861 -30 -13827
rect 4 -13861 38 -13827
rect 72 -13861 106 -13827
rect 140 -13861 174 -13827
rect 208 -13861 242 -13827
rect 276 -13861 310 -13827
rect 344 -13861 403 -13827
rect -584 -13903 -442 -13887
rect -526 -13909 -442 -13903
rect -57 -13871 403 -13861
rect -57 -13909 -27 -13871
rect 29 -13909 59 -13871
rect 115 -13909 145 -13871
rect 201 -13909 231 -13871
rect 287 -13909 317 -13871
rect 373 -13909 403 -13871
rect 612 -13853 754 -13837
rect 612 -13887 628 -13853
rect 662 -13887 754 -13853
rect 796 -13851 888 -13817
rect 922 -13851 938 -13817
rect 796 -13867 938 -13851
rect 1072 -13827 1243 -13811
rect 1072 -13861 1082 -13827
rect 1116 -13851 1243 -13827
rect 1624 -13801 1708 -13795
rect 2084 -13801 2168 -13795
rect 1624 -13817 1766 -13801
rect 1116 -13861 1244 -13851
rect 1072 -13877 1244 -13861
rect 612 -13903 754 -13887
rect 670 -13909 754 -13903
rect 1130 -13881 1244 -13877
rect -1354 -13935 -1144 -13909
rect -526 -13935 -316 -13909
rect 670 -13935 880 -13909
rect 1130 -13941 1160 -13881
rect 1214 -13941 1244 -13881
rect 1440 -13853 1582 -13837
rect 1440 -13887 1456 -13853
rect 1490 -13887 1582 -13853
rect 1624 -13851 1716 -13817
rect 1750 -13851 1766 -13817
rect 2084 -13817 2226 -13801
rect 2420 -13815 2450 -13743
rect 1624 -13867 1766 -13851
rect 1900 -13853 2042 -13837
rect 1440 -13903 1582 -13887
rect 1900 -13887 1916 -13853
rect 1950 -13887 2042 -13853
rect 2084 -13851 2176 -13817
rect 2210 -13851 2226 -13817
rect 2084 -13867 2226 -13851
rect 2380 -13827 2450 -13815
rect 2522 -13817 2622 -13789
rect 2782 -13817 2882 -13789
rect 2947 -13811 2977 -13743
rect 3246 -13795 3456 -13769
rect 4442 -13795 5388 -13769
rect 6466 -13795 6676 -13769
rect 3372 -13801 3456 -13795
rect 2380 -13861 2396 -13827
rect 2430 -13861 2450 -13827
rect 2380 -13874 2450 -13861
rect 2500 -13827 2622 -13817
rect 2500 -13861 2516 -13827
rect 2550 -13861 2622 -13827
rect 2500 -13871 2622 -13861
rect 2721 -13827 2882 -13817
rect 2721 -13861 2737 -13827
rect 2771 -13861 2882 -13827
rect 2721 -13871 2882 -13861
rect 1900 -13903 2042 -13887
rect 1498 -13909 1582 -13903
rect 1958 -13909 2042 -13903
rect 2420 -13909 2450 -13874
rect 1498 -13935 1708 -13909
rect 1958 -13935 2168 -13909
rect 2522 -13945 2622 -13871
rect 2782 -13945 2882 -13871
rect 2927 -13827 2981 -13811
rect 2927 -13861 2937 -13827
rect 2971 -13861 2981 -13827
rect 3372 -13817 3514 -13801
rect 2927 -13877 2981 -13861
rect 3188 -13853 3330 -13837
rect 2947 -13909 2977 -13877
rect 3188 -13887 3204 -13853
rect 3238 -13887 3330 -13853
rect 3372 -13851 3464 -13817
rect 3498 -13851 3514 -13817
rect 4934 -13817 5388 -13795
rect 3372 -13867 3514 -13851
rect 4442 -13853 4892 -13837
rect 3188 -13903 3330 -13887
rect 3246 -13909 3330 -13903
rect 4442 -13887 4458 -13853
rect 4492 -13887 4586 -13853
rect 4620 -13887 4714 -13853
rect 4748 -13887 4842 -13853
rect 4876 -13887 4892 -13853
rect 4934 -13851 4950 -13817
rect 4984 -13851 5078 -13817
rect 5112 -13851 5206 -13817
rect 5240 -13851 5334 -13817
rect 5368 -13851 5388 -13817
rect 6592 -13801 6676 -13795
rect 6592 -13817 6734 -13801
rect 6928 -13815 6958 -13743
rect 4934 -13867 5388 -13851
rect 6408 -13853 6550 -13837
rect 4442 -13909 4892 -13887
rect 6408 -13887 6424 -13853
rect 6458 -13887 6550 -13853
rect 6592 -13851 6684 -13817
rect 6718 -13851 6734 -13817
rect 6592 -13867 6734 -13851
rect 6888 -13827 6958 -13815
rect 7030 -13817 7130 -13789
rect 7290 -13817 7390 -13789
rect 7455 -13811 7485 -13743
rect 7754 -13795 7964 -13769
rect 7880 -13801 7964 -13795
rect 6888 -13861 6904 -13827
rect 6938 -13861 6958 -13827
rect 6888 -13874 6958 -13861
rect 7008 -13827 7130 -13817
rect 7008 -13861 7024 -13827
rect 7058 -13861 7130 -13827
rect 7008 -13871 7130 -13861
rect 7229 -13827 7390 -13817
rect 7229 -13861 7245 -13827
rect 7279 -13861 7390 -13827
rect 7229 -13871 7390 -13861
rect 6408 -13903 6550 -13887
rect 6466 -13909 6550 -13903
rect 6928 -13909 6958 -13874
rect 3246 -13935 3456 -13909
rect 4442 -13935 5388 -13909
rect 6466 -13935 6676 -13909
rect 7030 -13945 7130 -13871
rect 7290 -13945 7390 -13871
rect 7435 -13827 7489 -13811
rect 7435 -13861 7445 -13827
rect 7479 -13861 7489 -13827
rect 7880 -13817 8022 -13801
rect 8216 -13815 8246 -13743
rect 7435 -13877 7489 -13861
rect 7696 -13853 7838 -13837
rect 7455 -13909 7485 -13877
rect 7696 -13887 7712 -13853
rect 7746 -13887 7838 -13853
rect 7880 -13851 7972 -13817
rect 8006 -13851 8022 -13817
rect 7880 -13867 8022 -13851
rect 8176 -13827 8246 -13815
rect 8318 -13817 8418 -13789
rect 8578 -13817 8678 -13789
rect 8743 -13811 8773 -13743
rect 9042 -13795 9252 -13769
rect 9168 -13801 9252 -13795
rect 8176 -13861 8192 -13827
rect 8226 -13861 8246 -13827
rect 8176 -13874 8246 -13861
rect 8296 -13827 8418 -13817
rect 8296 -13861 8312 -13827
rect 8346 -13861 8418 -13827
rect 8296 -13871 8418 -13861
rect 8517 -13827 8678 -13817
rect 8517 -13861 8533 -13827
rect 8567 -13861 8678 -13827
rect 8517 -13871 8678 -13861
rect 7696 -13903 7838 -13887
rect 7754 -13909 7838 -13903
rect 8216 -13909 8246 -13874
rect 7754 -13935 7964 -13909
rect 8318 -13945 8418 -13871
rect 8578 -13945 8678 -13871
rect 8723 -13827 8777 -13811
rect 8723 -13861 8733 -13827
rect 8767 -13861 8777 -13827
rect 9168 -13817 9310 -13801
rect 9504 -13815 9534 -13743
rect 8723 -13877 8777 -13861
rect 8984 -13853 9126 -13837
rect 8743 -13909 8773 -13877
rect 8984 -13887 9000 -13853
rect 9034 -13887 9126 -13853
rect 9168 -13851 9260 -13817
rect 9294 -13851 9310 -13817
rect 9168 -13867 9310 -13851
rect 9464 -13827 9534 -13815
rect 9606 -13817 9706 -13789
rect 9866 -13817 9966 -13789
rect 10031 -13811 10061 -13743
rect 10330 -13795 10540 -13769
rect 10456 -13801 10540 -13795
rect 9464 -13861 9480 -13827
rect 9514 -13861 9534 -13827
rect 9464 -13874 9534 -13861
rect 9584 -13827 9706 -13817
rect 9584 -13861 9600 -13827
rect 9634 -13861 9706 -13827
rect 9584 -13871 9706 -13861
rect 9805 -13827 9966 -13817
rect 9805 -13861 9821 -13827
rect 9855 -13861 9966 -13827
rect 9805 -13871 9966 -13861
rect 8984 -13903 9126 -13887
rect 9042 -13909 9126 -13903
rect 9504 -13909 9534 -13874
rect 9042 -13935 9252 -13909
rect 9606 -13945 9706 -13871
rect 9866 -13945 9966 -13871
rect 10011 -13827 10065 -13811
rect 10011 -13861 10021 -13827
rect 10055 -13861 10065 -13827
rect 10456 -13817 10598 -13801
rect 10790 -13811 10820 -13789
rect 10874 -13811 10904 -13789
rect 10958 -13811 10988 -13789
rect 11042 -13811 11072 -13789
rect 10011 -13877 10065 -13861
rect 10272 -13853 10414 -13837
rect 10031 -13909 10061 -13877
rect 10272 -13887 10288 -13853
rect 10322 -13887 10414 -13853
rect 10456 -13851 10548 -13817
rect 10582 -13851 10598 -13817
rect 10456 -13867 10598 -13851
rect 10733 -13827 11072 -13811
rect 10733 -13861 10749 -13827
rect 10783 -13861 10830 -13827
rect 10864 -13861 10914 -13827
rect 10948 -13861 10998 -13827
rect 11032 -13861 11072 -13827
rect 10733 -13877 11072 -13861
rect 10272 -13903 10414 -13887
rect 10330 -13909 10414 -13903
rect 10790 -13909 10820 -13877
rect 10874 -13909 10904 -13877
rect 10958 -13909 10988 -13877
rect 11042 -13909 11072 -13877
rect 11126 -13811 11156 -13789
rect 11210 -13811 11240 -13789
rect 11294 -13811 11324 -13789
rect 11378 -13811 11408 -13789
rect 11710 -13795 11920 -13769
rect 13642 -13795 14588 -13769
rect 14838 -13795 15784 -13769
rect 16034 -13795 16612 -13769
rect 11126 -13827 11408 -13811
rect 11126 -13861 11250 -13827
rect 11284 -13861 11334 -13827
rect 11368 -13861 11408 -13827
rect 11836 -13801 11920 -13795
rect 11836 -13817 11978 -13801
rect 11126 -13877 11408 -13861
rect 11126 -13909 11156 -13877
rect 11210 -13909 11240 -13877
rect 11294 -13909 11324 -13877
rect 11378 -13909 11408 -13877
rect 11652 -13853 11794 -13837
rect 11652 -13887 11668 -13853
rect 11702 -13887 11794 -13853
rect 11836 -13851 11928 -13817
rect 11962 -13851 11978 -13817
rect 14134 -13817 14588 -13795
rect 11836 -13867 11978 -13851
rect 13642 -13853 14092 -13837
rect 11652 -13903 11794 -13887
rect 11710 -13909 11794 -13903
rect 13642 -13887 13658 -13853
rect 13692 -13887 13786 -13853
rect 13820 -13887 13914 -13853
rect 13948 -13887 14042 -13853
rect 14076 -13887 14092 -13853
rect 14134 -13851 14150 -13817
rect 14184 -13851 14278 -13817
rect 14312 -13851 14406 -13817
rect 14440 -13851 14534 -13817
rect 14568 -13851 14588 -13817
rect 15330 -13817 15784 -13795
rect 14134 -13867 14588 -13851
rect 14838 -13853 15288 -13837
rect 13642 -13909 14092 -13887
rect 14838 -13887 14854 -13853
rect 14888 -13887 14982 -13853
rect 15016 -13887 15110 -13853
rect 15144 -13887 15238 -13853
rect 15272 -13887 15288 -13853
rect 15330 -13851 15346 -13817
rect 15380 -13851 15474 -13817
rect 15508 -13851 15602 -13817
rect 15636 -13851 15730 -13817
rect 15764 -13851 15784 -13817
rect 16340 -13817 16612 -13795
rect 15330 -13867 15784 -13851
rect 16034 -13853 16298 -13837
rect 14838 -13909 15288 -13887
rect 16034 -13887 16050 -13853
rect 16084 -13887 16149 -13853
rect 16183 -13887 16248 -13853
rect 16282 -13887 16298 -13853
rect 16340 -13851 16356 -13817
rect 16390 -13851 16459 -13817
rect 16493 -13851 16562 -13817
rect 16596 -13851 16612 -13817
rect 16340 -13867 16612 -13851
rect 16034 -13909 16298 -13887
rect 10330 -13935 10540 -13909
rect 11710 -13935 11920 -13909
rect 13642 -13935 14588 -13909
rect 14838 -13935 15784 -13909
rect 16034 -13935 16612 -13909
rect -2918 -14135 -2340 -14109
rect -1354 -14135 -1144 -14109
rect -890 -14135 -860 -14109
rect -806 -14135 -776 -14109
rect -526 -14135 -316 -14109
rect -57 -14135 -27 -14109
rect 29 -14135 59 -14109
rect 115 -14135 145 -14109
rect 201 -14135 231 -14109
rect 287 -14135 317 -14109
rect 373 -14135 403 -14109
rect 670 -14135 880 -14109
rect 1130 -14135 1160 -14109
rect 1214 -14135 1244 -14109
rect 1498 -14135 1708 -14109
rect 1958 -14135 2168 -14109
rect 2420 -14135 2450 -14109
rect 2522 -14135 2622 -14109
rect 2782 -14135 2882 -14109
rect 2947 -14135 2977 -14109
rect 3246 -14135 3456 -14109
rect 4442 -14135 5388 -14109
rect 6466 -14135 6676 -14109
rect 6928 -14135 6958 -14109
rect 7030 -14135 7130 -14109
rect 7290 -14135 7390 -14109
rect 7455 -14135 7485 -14109
rect 7754 -14135 7964 -14109
rect 8216 -14135 8246 -14109
rect 8318 -14135 8418 -14109
rect 8578 -14135 8678 -14109
rect 8743 -14135 8773 -14109
rect 9042 -14135 9252 -14109
rect 9504 -14135 9534 -14109
rect 9606 -14135 9706 -14109
rect 9866 -14135 9966 -14109
rect 10031 -14135 10061 -14109
rect 10330 -14135 10540 -14109
rect 10790 -14135 10820 -14109
rect 10874 -14135 10904 -14109
rect 10958 -14135 10988 -14109
rect 11042 -14135 11072 -14109
rect 11126 -14135 11156 -14109
rect 11210 -14135 11240 -14109
rect 11294 -14135 11324 -14109
rect 11378 -14135 11408 -14109
rect 11710 -14135 11920 -14109
rect 13642 -14135 14588 -14109
rect 14838 -14135 15784 -14109
rect 16034 -14135 16612 -14109
<< polycont >>
rect -2902 -315 -2868 -281
rect -2803 -315 -2769 -281
rect -2704 -315 -2670 -281
rect -2596 -351 -2562 -317
rect -2493 -351 -2459 -317
rect -2390 -351 -2356 -317
rect -1396 -315 -1362 -281
rect -1136 -351 -1102 -317
rect -937 -341 -903 -307
rect -769 -341 -735 -307
rect -568 -315 -534 -281
rect -308 -351 -274 -317
rect -30 -341 4 -307
rect 38 -341 72 -307
rect 106 -341 140 -307
rect 174 -341 208 -307
rect 242 -341 276 -307
rect 310 -341 344 -307
rect 628 -315 662 -281
rect 888 -351 922 -317
rect 1082 -341 1116 -307
rect 1456 -315 1490 -281
rect 1716 -351 1750 -317
rect 1916 -315 1950 -281
rect 2176 -351 2210 -317
rect 2396 -341 2430 -307
rect 2516 -341 2550 -307
rect 2737 -341 2771 -307
rect 2937 -341 2971 -307
rect 3204 -315 3238 -281
rect 3464 -351 3498 -317
rect 4458 -315 4492 -281
rect 4586 -315 4620 -281
rect 4714 -315 4748 -281
rect 4842 -315 4876 -281
rect 4950 -351 4984 -317
rect 5078 -351 5112 -317
rect 5206 -351 5240 -317
rect 5334 -351 5368 -317
rect 6424 -315 6458 -281
rect 6684 -351 6718 -317
rect 6904 -341 6938 -307
rect 7024 -341 7058 -307
rect 7245 -341 7279 -307
rect 7445 -341 7479 -307
rect 7712 -315 7746 -281
rect 7972 -351 8006 -317
rect 8192 -341 8226 -307
rect 8312 -341 8346 -307
rect 8533 -341 8567 -307
rect 8733 -341 8767 -307
rect 9000 -315 9034 -281
rect 9260 -351 9294 -317
rect 9480 -341 9514 -307
rect 9600 -341 9634 -307
rect 9821 -341 9855 -307
rect 10021 -341 10055 -307
rect 10288 -315 10322 -281
rect 10548 -351 10582 -317
rect 10749 -341 10783 -307
rect 10830 -341 10864 -307
rect 10914 -341 10948 -307
rect 10998 -341 11032 -307
rect 11250 -341 11284 -307
rect 11334 -341 11368 -307
rect 11668 -315 11702 -281
rect 11928 -351 11962 -317
rect 13658 -315 13692 -281
rect 13786 -315 13820 -281
rect 13914 -315 13948 -281
rect 14042 -315 14076 -281
rect 14150 -351 14184 -317
rect 14278 -351 14312 -317
rect 14406 -351 14440 -317
rect 14534 -351 14568 -317
rect 14854 -315 14888 -281
rect 14982 -315 15016 -281
rect 15110 -315 15144 -281
rect 15238 -315 15272 -281
rect 15346 -351 15380 -317
rect 15474 -351 15508 -317
rect 15602 -351 15636 -317
rect 15730 -351 15764 -317
rect 16050 -315 16084 -281
rect 16149 -315 16183 -281
rect 16248 -315 16282 -281
rect 16356 -351 16390 -317
rect 16459 -351 16493 -317
rect 16562 -351 16596 -317
rect -2902 -795 -2868 -761
rect -2799 -795 -2765 -761
rect -2696 -795 -2662 -761
rect -2588 -831 -2554 -797
rect -2489 -831 -2455 -797
rect -2390 -831 -2356 -797
rect -1522 -795 -1488 -761
rect -1419 -795 -1385 -761
rect -1316 -795 -1282 -761
rect -1208 -831 -1174 -797
rect -1109 -831 -1075 -797
rect -1010 -831 -976 -797
rect -786 -795 -752 -761
rect -683 -795 -649 -761
rect -580 -795 -546 -761
rect -472 -831 -438 -797
rect -373 -831 -339 -797
rect -274 -831 -240 -797
rect -16 -795 18 -761
rect 244 -831 278 -797
rect 511 -805 545 -771
rect 711 -805 745 -771
rect 932 -805 966 -771
rect 1052 -805 1086 -771
rect 1272 -795 1306 -761
rect 1532 -831 1566 -797
rect 1790 -795 1824 -761
rect 1893 -795 1927 -761
rect 1996 -795 2030 -761
rect 2104 -831 2138 -797
rect 2203 -831 2237 -797
rect 2302 -831 2336 -797
rect 2560 -795 2594 -761
rect 2820 -831 2854 -797
rect 3087 -805 3121 -771
rect 3287 -805 3321 -771
rect 3508 -805 3542 -771
rect 3628 -805 3662 -771
rect 3848 -795 3882 -761
rect 4108 -831 4142 -797
rect 4366 -795 4400 -761
rect 4469 -795 4503 -761
rect 4572 -795 4606 -761
rect 4680 -831 4714 -797
rect 4779 -831 4813 -797
rect 4878 -831 4912 -797
rect 5136 -795 5170 -761
rect 5396 -831 5430 -797
rect 5663 -805 5697 -771
rect 5863 -805 5897 -771
rect 6084 -805 6118 -771
rect 6204 -805 6238 -771
rect 6424 -795 6458 -761
rect 6684 -831 6718 -797
rect 6942 -795 6976 -761
rect 7045 -795 7079 -761
rect 7148 -795 7182 -761
rect 7256 -831 7290 -797
rect 7355 -831 7389 -797
rect 7454 -831 7488 -797
rect 7712 -795 7746 -761
rect 7972 -831 8006 -797
rect 8239 -805 8273 -771
rect 8439 -805 8473 -771
rect 8660 -805 8694 -771
rect 8780 -805 8814 -771
rect 9000 -795 9034 -761
rect 9260 -831 9294 -797
rect 9518 -795 9552 -761
rect 9621 -795 9655 -761
rect 9724 -795 9758 -761
rect 9832 -831 9866 -797
rect 9931 -831 9965 -797
rect 10030 -831 10064 -797
rect 10380 -795 10414 -761
rect 10640 -831 10674 -797
rect 10815 -805 10849 -771
rect 11015 -805 11049 -771
rect 11236 -805 11270 -771
rect 11356 -805 11390 -771
rect 11668 -795 11702 -761
rect 11928 -831 11962 -797
rect 13692 -805 13726 -771
rect 14119 -805 14153 -771
rect 14187 -805 14221 -771
rect 14255 -805 14289 -771
rect 14323 -805 14357 -771
rect 14391 -805 14425 -771
rect 14459 -805 14493 -771
rect 14527 -805 14561 -771
rect 14595 -805 14629 -771
rect 14663 -805 14697 -771
rect 14731 -805 14765 -771
rect 14799 -805 14833 -771
rect 14867 -805 14901 -771
rect 14935 -805 14969 -771
rect 15003 -805 15037 -771
rect 15071 -805 15105 -771
rect 15139 -805 15173 -771
rect 15686 -795 15720 -761
rect 15814 -795 15848 -761
rect 15942 -795 15976 -761
rect 16070 -795 16104 -761
rect 16178 -831 16212 -797
rect 16306 -831 16340 -797
rect 16434 -831 16468 -797
rect 16562 -831 16596 -797
rect -2902 -1403 -2868 -1369
rect -2803 -1403 -2769 -1369
rect -2704 -1403 -2670 -1369
rect -2596 -1439 -2562 -1405
rect -2493 -1439 -2459 -1405
rect -2390 -1439 -2356 -1405
rect -1522 -1403 -1488 -1369
rect -1423 -1403 -1389 -1369
rect -1324 -1403 -1290 -1369
rect -1216 -1439 -1182 -1405
rect -1113 -1439 -1079 -1405
rect -1010 -1439 -976 -1405
rect -786 -1403 -752 -1369
rect -687 -1403 -653 -1369
rect -588 -1403 -554 -1369
rect -480 -1439 -446 -1405
rect -377 -1439 -343 -1405
rect -274 -1439 -240 -1405
rect -16 -1439 18 -1405
rect 244 -1403 278 -1369
rect 464 -1429 498 -1395
rect 584 -1429 618 -1395
rect 805 -1429 839 -1395
rect 1005 -1429 1039 -1395
rect 1272 -1439 1306 -1405
rect 1532 -1403 1566 -1369
rect 1790 -1403 1824 -1369
rect 1889 -1403 1923 -1369
rect 1988 -1403 2022 -1369
rect 2096 -1439 2130 -1405
rect 2199 -1439 2233 -1405
rect 2302 -1439 2336 -1405
rect 2560 -1439 2594 -1405
rect 2820 -1403 2854 -1369
rect 3040 -1429 3074 -1395
rect 3160 -1429 3194 -1395
rect 3381 -1429 3415 -1395
rect 3581 -1429 3615 -1395
rect 3848 -1439 3882 -1405
rect 4108 -1403 4142 -1369
rect 4366 -1403 4400 -1369
rect 4465 -1403 4499 -1369
rect 4564 -1403 4598 -1369
rect 4672 -1439 4706 -1405
rect 4775 -1439 4809 -1405
rect 4878 -1439 4912 -1405
rect 5136 -1439 5170 -1405
rect 5396 -1403 5430 -1369
rect 5616 -1429 5650 -1395
rect 5736 -1429 5770 -1395
rect 5957 -1429 5991 -1395
rect 6157 -1429 6191 -1395
rect 6424 -1439 6458 -1405
rect 6684 -1403 6718 -1369
rect 6942 -1403 6976 -1369
rect 7041 -1403 7075 -1369
rect 7140 -1403 7174 -1369
rect 7248 -1439 7282 -1405
rect 7351 -1439 7385 -1405
rect 7454 -1439 7488 -1405
rect 7712 -1439 7746 -1405
rect 7972 -1403 8006 -1369
rect 8192 -1429 8226 -1395
rect 8312 -1429 8346 -1395
rect 8533 -1429 8567 -1395
rect 8733 -1429 8767 -1395
rect 9000 -1439 9034 -1405
rect 9260 -1403 9294 -1369
rect 9518 -1403 9552 -1369
rect 9617 -1403 9651 -1369
rect 9716 -1403 9750 -1369
rect 9824 -1439 9858 -1405
rect 9927 -1439 9961 -1405
rect 10030 -1439 10064 -1405
rect 10380 -1439 10414 -1405
rect 10640 -1403 10674 -1369
rect 10768 -1429 10802 -1395
rect 10888 -1429 10922 -1395
rect 11109 -1429 11143 -1395
rect 11309 -1429 11343 -1395
rect 11668 -1439 11702 -1405
rect 11928 -1403 11962 -1369
rect 12574 -1429 12608 -1395
rect 12642 -1429 12676 -1395
rect 12710 -1429 12744 -1395
rect 12778 -1429 12812 -1395
rect 12846 -1429 12880 -1395
rect 12914 -1429 12948 -1395
rect 13232 -1403 13266 -1369
rect 13492 -1439 13526 -1405
rect 13692 -1429 13726 -1395
rect 14119 -1429 14153 -1395
rect 14187 -1429 14221 -1395
rect 14255 -1429 14289 -1395
rect 14323 -1429 14357 -1395
rect 14391 -1429 14425 -1395
rect 14459 -1429 14493 -1395
rect 14527 -1429 14561 -1395
rect 14595 -1429 14629 -1395
rect 14663 -1429 14697 -1395
rect 14731 -1429 14765 -1395
rect 14799 -1429 14833 -1395
rect 14867 -1429 14901 -1395
rect 14935 -1429 14969 -1395
rect 15003 -1429 15037 -1395
rect 15071 -1429 15105 -1395
rect 15139 -1429 15173 -1395
rect 15682 -1403 15716 -1369
rect 15810 -1403 15844 -1369
rect 15938 -1403 15972 -1369
rect 16066 -1403 16100 -1369
rect 16174 -1439 16208 -1405
rect 16302 -1439 16336 -1405
rect 16430 -1439 16464 -1405
rect 16558 -1439 16592 -1405
rect -2902 -1883 -2868 -1849
rect -2799 -1883 -2765 -1849
rect -2696 -1883 -2662 -1849
rect -2588 -1919 -2554 -1885
rect -2489 -1919 -2455 -1885
rect -2390 -1919 -2356 -1885
rect -1522 -1883 -1488 -1849
rect -1419 -1883 -1385 -1849
rect -1316 -1883 -1282 -1849
rect -1208 -1919 -1174 -1885
rect -1109 -1919 -1075 -1885
rect -1010 -1919 -976 -1885
rect -777 -1893 -743 -1859
rect -577 -1893 -543 -1859
rect -356 -1893 -322 -1859
rect -236 -1893 -202 -1859
rect -16 -1883 18 -1849
rect 244 -1919 278 -1885
rect 511 -1893 545 -1859
rect 711 -1893 745 -1859
rect 932 -1893 966 -1859
rect 1052 -1893 1086 -1859
rect 1272 -1883 1306 -1849
rect 1532 -1919 1566 -1885
rect 1790 -1883 1824 -1849
rect 1893 -1883 1927 -1849
rect 1996 -1883 2030 -1849
rect 2104 -1919 2138 -1885
rect 2203 -1919 2237 -1885
rect 2302 -1919 2336 -1885
rect 2560 -1883 2594 -1849
rect 2820 -1919 2854 -1885
rect 3087 -1893 3121 -1859
rect 3287 -1893 3321 -1859
rect 3508 -1893 3542 -1859
rect 3628 -1893 3662 -1859
rect 3848 -1883 3882 -1849
rect 4108 -1919 4142 -1885
rect 4366 -1883 4400 -1849
rect 4469 -1883 4503 -1849
rect 4572 -1883 4606 -1849
rect 4680 -1919 4714 -1885
rect 4779 -1919 4813 -1885
rect 4878 -1919 4912 -1885
rect 5136 -1883 5170 -1849
rect 5396 -1919 5430 -1885
rect 5663 -1893 5697 -1859
rect 5863 -1893 5897 -1859
rect 6084 -1893 6118 -1859
rect 6204 -1893 6238 -1859
rect 6424 -1883 6458 -1849
rect 6684 -1919 6718 -1885
rect 6942 -1883 6976 -1849
rect 7045 -1883 7079 -1849
rect 7148 -1883 7182 -1849
rect 7256 -1919 7290 -1885
rect 7355 -1919 7389 -1885
rect 7454 -1919 7488 -1885
rect 7712 -1883 7746 -1849
rect 7972 -1919 8006 -1885
rect 8239 -1893 8273 -1859
rect 8439 -1893 8473 -1859
rect 8660 -1893 8694 -1859
rect 8780 -1893 8814 -1859
rect 9000 -1883 9034 -1849
rect 9260 -1919 9294 -1885
rect 9518 -1883 9552 -1849
rect 9621 -1883 9655 -1849
rect 9724 -1883 9758 -1849
rect 9832 -1919 9866 -1885
rect 9931 -1919 9965 -1885
rect 10030 -1919 10064 -1885
rect 10380 -1883 10414 -1849
rect 10640 -1919 10674 -1885
rect 10815 -1893 10849 -1859
rect 11015 -1893 11049 -1859
rect 11236 -1893 11270 -1859
rect 11356 -1893 11390 -1859
rect 11668 -1883 11702 -1849
rect 11928 -1919 11962 -1885
rect 13692 -1893 13726 -1859
rect 14119 -1893 14153 -1859
rect 14187 -1893 14221 -1859
rect 14255 -1893 14289 -1859
rect 14323 -1893 14357 -1859
rect 14391 -1893 14425 -1859
rect 14459 -1893 14493 -1859
rect 14527 -1893 14561 -1859
rect 14595 -1893 14629 -1859
rect 14663 -1893 14697 -1859
rect 14731 -1893 14765 -1859
rect 14799 -1893 14833 -1859
rect 14867 -1893 14901 -1859
rect 14935 -1893 14969 -1859
rect 15003 -1893 15037 -1859
rect 15071 -1893 15105 -1859
rect 15139 -1893 15173 -1859
rect 15686 -1883 15720 -1849
rect 15814 -1883 15848 -1849
rect 15942 -1883 15976 -1849
rect 16070 -1883 16104 -1849
rect 16178 -1919 16212 -1885
rect 16306 -1919 16340 -1885
rect 16434 -1919 16468 -1885
rect 16562 -1919 16596 -1885
rect -2902 -2491 -2868 -2457
rect -2803 -2491 -2769 -2457
rect -2704 -2491 -2670 -2457
rect -2596 -2527 -2562 -2493
rect -2493 -2527 -2459 -2493
rect -2390 -2527 -2356 -2493
rect -1522 -2491 -1488 -2457
rect -1423 -2491 -1389 -2457
rect -1324 -2491 -1290 -2457
rect -1216 -2527 -1182 -2493
rect -1113 -2527 -1079 -2493
rect -1010 -2527 -976 -2493
rect -786 -2491 -752 -2457
rect -687 -2491 -653 -2457
rect -588 -2491 -554 -2457
rect -480 -2527 -446 -2493
rect -377 -2527 -343 -2493
rect -274 -2527 -240 -2493
rect -16 -2527 18 -2493
rect 244 -2491 278 -2457
rect 464 -2517 498 -2483
rect 584 -2517 618 -2483
rect 805 -2517 839 -2483
rect 1005 -2517 1039 -2483
rect 1272 -2527 1306 -2493
rect 1532 -2491 1566 -2457
rect 1790 -2491 1824 -2457
rect 1889 -2491 1923 -2457
rect 1988 -2491 2022 -2457
rect 2096 -2527 2130 -2493
rect 2199 -2527 2233 -2493
rect 2302 -2527 2336 -2493
rect 2560 -2527 2594 -2493
rect 2820 -2491 2854 -2457
rect 3040 -2517 3074 -2483
rect 3160 -2517 3194 -2483
rect 3381 -2517 3415 -2483
rect 3581 -2517 3615 -2483
rect 3848 -2527 3882 -2493
rect 4108 -2491 4142 -2457
rect 4366 -2491 4400 -2457
rect 4465 -2491 4499 -2457
rect 4564 -2491 4598 -2457
rect 4672 -2527 4706 -2493
rect 4775 -2527 4809 -2493
rect 4878 -2527 4912 -2493
rect 5136 -2527 5170 -2493
rect 5396 -2491 5430 -2457
rect 5616 -2517 5650 -2483
rect 5736 -2517 5770 -2483
rect 5957 -2517 5991 -2483
rect 6157 -2517 6191 -2483
rect 6424 -2527 6458 -2493
rect 6684 -2491 6718 -2457
rect 6942 -2491 6976 -2457
rect 7041 -2491 7075 -2457
rect 7140 -2491 7174 -2457
rect 7248 -2527 7282 -2493
rect 7351 -2527 7385 -2493
rect 7454 -2527 7488 -2493
rect 7712 -2527 7746 -2493
rect 7972 -2491 8006 -2457
rect 8192 -2517 8226 -2483
rect 8312 -2517 8346 -2483
rect 8533 -2517 8567 -2483
rect 8733 -2517 8767 -2483
rect 9000 -2527 9034 -2493
rect 9260 -2491 9294 -2457
rect 9518 -2491 9552 -2457
rect 9617 -2491 9651 -2457
rect 9716 -2491 9750 -2457
rect 9824 -2527 9858 -2493
rect 9927 -2527 9961 -2493
rect 10030 -2527 10064 -2493
rect 10380 -2527 10414 -2493
rect 10640 -2491 10674 -2457
rect 10768 -2517 10802 -2483
rect 10888 -2517 10922 -2483
rect 11109 -2517 11143 -2483
rect 11309 -2517 11343 -2483
rect 11668 -2527 11702 -2493
rect 11928 -2491 11962 -2457
rect 12574 -2517 12608 -2483
rect 12642 -2517 12676 -2483
rect 12710 -2517 12744 -2483
rect 12778 -2517 12812 -2483
rect 12846 -2517 12880 -2483
rect 12914 -2517 12948 -2483
rect 13232 -2491 13266 -2457
rect 13492 -2527 13526 -2493
rect 13692 -2517 13726 -2483
rect 14119 -2517 14153 -2483
rect 14187 -2517 14221 -2483
rect 14255 -2517 14289 -2483
rect 14323 -2517 14357 -2483
rect 14391 -2517 14425 -2483
rect 14459 -2517 14493 -2483
rect 14527 -2517 14561 -2483
rect 14595 -2517 14629 -2483
rect 14663 -2517 14697 -2483
rect 14731 -2517 14765 -2483
rect 14799 -2517 14833 -2483
rect 14867 -2517 14901 -2483
rect 14935 -2517 14969 -2483
rect 15003 -2517 15037 -2483
rect 15071 -2517 15105 -2483
rect 15139 -2517 15173 -2483
rect 15682 -2491 15716 -2457
rect 15810 -2491 15844 -2457
rect 15938 -2491 15972 -2457
rect 16066 -2491 16100 -2457
rect 16174 -2527 16208 -2493
rect 16302 -2527 16336 -2493
rect 16430 -2527 16464 -2493
rect 16558 -2527 16592 -2493
rect -2902 -2971 -2868 -2937
rect -2799 -2971 -2765 -2937
rect -2696 -2971 -2662 -2937
rect -2588 -3007 -2554 -2973
rect -2489 -3007 -2455 -2973
rect -2390 -3007 -2356 -2973
rect -1954 -2981 -1920 -2947
rect -1522 -2971 -1488 -2937
rect -1419 -2971 -1385 -2937
rect -1316 -2971 -1282 -2937
rect -1208 -3007 -1174 -2973
rect -1109 -3007 -1075 -2973
rect -1010 -3007 -976 -2973
rect -786 -2971 -752 -2937
rect -683 -2971 -649 -2937
rect -580 -2971 -546 -2937
rect -472 -3007 -438 -2973
rect -373 -3007 -339 -2973
rect -274 -3007 -240 -2973
rect -16 -2971 18 -2937
rect 244 -3007 278 -2973
rect 511 -2981 545 -2947
rect 711 -2981 745 -2947
rect 932 -2981 966 -2947
rect 1052 -2981 1086 -2947
rect 1272 -2971 1306 -2937
rect 1532 -3007 1566 -2973
rect 1790 -2971 1824 -2937
rect 1893 -2971 1927 -2937
rect 1996 -2971 2030 -2937
rect 2104 -3007 2138 -2973
rect 2203 -3007 2237 -2973
rect 2302 -3007 2336 -2973
rect 2560 -2971 2594 -2937
rect 2820 -3007 2854 -2973
rect 3087 -2981 3121 -2947
rect 3287 -2981 3321 -2947
rect 3508 -2981 3542 -2947
rect 3628 -2981 3662 -2947
rect 3848 -2971 3882 -2937
rect 4108 -3007 4142 -2973
rect 4366 -2971 4400 -2937
rect 4469 -2971 4503 -2937
rect 4572 -2971 4606 -2937
rect 4680 -3007 4714 -2973
rect 4779 -3007 4813 -2973
rect 4878 -3007 4912 -2973
rect 5136 -2971 5170 -2937
rect 5396 -3007 5430 -2973
rect 5663 -2981 5697 -2947
rect 5863 -2981 5897 -2947
rect 6084 -2981 6118 -2947
rect 6204 -2981 6238 -2947
rect 6424 -2971 6458 -2937
rect 6684 -3007 6718 -2973
rect 6942 -2971 6976 -2937
rect 7045 -2971 7079 -2937
rect 7148 -2971 7182 -2937
rect 7256 -3007 7290 -2973
rect 7355 -3007 7389 -2973
rect 7454 -3007 7488 -2973
rect 7712 -2971 7746 -2937
rect 7972 -3007 8006 -2973
rect 8239 -2981 8273 -2947
rect 8439 -2981 8473 -2947
rect 8660 -2981 8694 -2947
rect 8780 -2981 8814 -2947
rect 9000 -2971 9034 -2937
rect 9260 -3007 9294 -2973
rect 9518 -2971 9552 -2937
rect 9621 -2971 9655 -2937
rect 9724 -2971 9758 -2937
rect 9832 -3007 9866 -2973
rect 9931 -3007 9965 -2973
rect 10030 -3007 10064 -2973
rect 10380 -2971 10414 -2937
rect 10640 -3007 10674 -2973
rect 10815 -2981 10849 -2947
rect 11015 -2981 11049 -2947
rect 11236 -2981 11270 -2947
rect 11356 -2981 11390 -2947
rect 11668 -2971 11702 -2937
rect 11928 -3007 11962 -2973
rect 13662 -2971 13696 -2937
rect 13790 -2971 13824 -2937
rect 13918 -2971 13952 -2937
rect 14046 -2971 14080 -2937
rect 14154 -3007 14188 -2973
rect 14282 -3007 14316 -2973
rect 14410 -3007 14444 -2973
rect 14538 -3007 14572 -2973
rect 14858 -2971 14892 -2937
rect 14986 -2971 15020 -2937
rect 15114 -2971 15148 -2937
rect 15242 -2971 15276 -2937
rect 15350 -3007 15384 -2973
rect 15478 -3007 15512 -2973
rect 15606 -3007 15640 -2973
rect 15734 -3007 15768 -2973
rect 16050 -2971 16084 -2937
rect 16153 -2971 16187 -2937
rect 16256 -2971 16290 -2937
rect 16364 -3007 16398 -2973
rect 16463 -3007 16497 -2973
rect 16562 -3007 16596 -2973
rect -2902 -3579 -2868 -3545
rect -2803 -3579 -2769 -3545
rect -2704 -3579 -2670 -3545
rect -2596 -3615 -2562 -3581
rect -2493 -3615 -2459 -3581
rect -2390 -3615 -2356 -3581
rect -1522 -3615 -1488 -3581
rect -1419 -3615 -1385 -3581
rect -1316 -3615 -1282 -3581
rect -1208 -3579 -1174 -3545
rect -1109 -3579 -1075 -3545
rect -1010 -3579 -976 -3545
rect -786 -3615 -752 -3581
rect -683 -3615 -649 -3581
rect -580 -3615 -546 -3581
rect -472 -3579 -438 -3545
rect -373 -3579 -339 -3545
rect -274 -3579 -240 -3545
rect -16 -3615 18 -3581
rect 244 -3579 278 -3545
rect 511 -3605 545 -3571
rect 711 -3605 745 -3571
rect 932 -3605 966 -3571
rect 1052 -3605 1086 -3571
rect 1272 -3615 1306 -3581
rect 1532 -3579 1566 -3545
rect 1790 -3579 1824 -3545
rect 1889 -3579 1923 -3545
rect 1988 -3579 2022 -3545
rect 2096 -3615 2130 -3581
rect 2199 -3615 2233 -3581
rect 2302 -3615 2336 -3581
rect 2560 -3615 2594 -3581
rect 2820 -3579 2854 -3545
rect 3087 -3605 3121 -3571
rect 3287 -3605 3321 -3571
rect 3508 -3605 3542 -3571
rect 3628 -3605 3662 -3571
rect 3848 -3615 3882 -3581
rect 4108 -3579 4142 -3545
rect 4366 -3579 4400 -3545
rect 4465 -3579 4499 -3545
rect 4564 -3579 4598 -3545
rect 4672 -3615 4706 -3581
rect 4775 -3615 4809 -3581
rect 4878 -3615 4912 -3581
rect 5136 -3615 5170 -3581
rect 5396 -3579 5430 -3545
rect 5663 -3605 5697 -3571
rect 5863 -3605 5897 -3571
rect 6084 -3605 6118 -3571
rect 6204 -3605 6238 -3571
rect 6424 -3615 6458 -3581
rect 6684 -3579 6718 -3545
rect 6942 -3579 6976 -3545
rect 7041 -3579 7075 -3545
rect 7140 -3579 7174 -3545
rect 7248 -3615 7282 -3581
rect 7351 -3615 7385 -3581
rect 7454 -3615 7488 -3581
rect 7712 -3615 7746 -3581
rect 7972 -3579 8006 -3545
rect 8239 -3605 8273 -3571
rect 8439 -3605 8473 -3571
rect 8660 -3605 8694 -3571
rect 8780 -3605 8814 -3571
rect 9000 -3615 9034 -3581
rect 9260 -3579 9294 -3545
rect 9518 -3579 9552 -3545
rect 9617 -3579 9651 -3545
rect 9716 -3579 9750 -3545
rect 9824 -3615 9858 -3581
rect 9927 -3615 9961 -3581
rect 10030 -3615 10064 -3581
rect 10380 -3615 10414 -3581
rect 10640 -3579 10674 -3545
rect 10815 -3605 10849 -3571
rect 11015 -3605 11049 -3571
rect 11236 -3605 11270 -3571
rect 11356 -3605 11390 -3571
rect 11668 -3615 11702 -3581
rect 11928 -3579 11962 -3545
rect 13662 -3615 13696 -3581
rect 13790 -3615 13824 -3581
rect 13918 -3615 13952 -3581
rect 14046 -3615 14080 -3581
rect 14154 -3579 14188 -3545
rect 14282 -3579 14316 -3545
rect 14410 -3579 14444 -3545
rect 14538 -3579 14572 -3545
rect 14858 -3615 14892 -3581
rect 14986 -3615 15020 -3581
rect 15114 -3615 15148 -3581
rect 15242 -3615 15276 -3581
rect 15350 -3579 15384 -3545
rect 15478 -3579 15512 -3545
rect 15606 -3579 15640 -3545
rect 15734 -3579 15768 -3545
rect 16050 -3615 16084 -3581
rect 16153 -3615 16187 -3581
rect 16256 -3615 16290 -3581
rect 16364 -3579 16398 -3545
rect 16463 -3579 16497 -3545
rect 16562 -3579 16596 -3545
rect -2902 -4059 -2868 -4025
rect -2799 -4059 -2765 -4025
rect -2696 -4059 -2662 -4025
rect -2588 -4095 -2554 -4061
rect -2489 -4095 -2455 -4061
rect -2390 -4095 -2356 -4061
rect -1522 -4095 -1488 -4061
rect -1423 -4095 -1389 -4061
rect -1324 -4095 -1290 -4061
rect -1216 -4059 -1182 -4025
rect -1113 -4059 -1079 -4025
rect -1010 -4059 -976 -4025
rect -786 -4095 -752 -4061
rect -687 -4095 -653 -4061
rect -588 -4095 -554 -4061
rect -480 -4059 -446 -4025
rect -377 -4059 -343 -4025
rect -274 -4059 -240 -4025
rect -16 -4059 18 -4025
rect 244 -4095 278 -4061
rect 464 -4069 498 -4035
rect 584 -4069 618 -4035
rect 805 -4069 839 -4035
rect 1005 -4069 1039 -4035
rect 1272 -4059 1306 -4025
rect 1532 -4095 1566 -4061
rect 1790 -4059 1824 -4025
rect 1893 -4059 1927 -4025
rect 1996 -4059 2030 -4025
rect 2104 -4095 2138 -4061
rect 2203 -4095 2237 -4061
rect 2302 -4095 2336 -4061
rect 2560 -4059 2594 -4025
rect 2820 -4095 2854 -4061
rect 3040 -4069 3074 -4035
rect 3160 -4069 3194 -4035
rect 3381 -4069 3415 -4035
rect 3581 -4069 3615 -4035
rect 3848 -4059 3882 -4025
rect 4108 -4095 4142 -4061
rect 4366 -4059 4400 -4025
rect 4469 -4059 4503 -4025
rect 4572 -4059 4606 -4025
rect 4680 -4095 4714 -4061
rect 4779 -4095 4813 -4061
rect 4878 -4095 4912 -4061
rect 5136 -4059 5170 -4025
rect 5396 -4095 5430 -4061
rect 5616 -4069 5650 -4035
rect 5736 -4069 5770 -4035
rect 5957 -4069 5991 -4035
rect 6157 -4069 6191 -4035
rect 6424 -4059 6458 -4025
rect 6684 -4095 6718 -4061
rect 6942 -4059 6976 -4025
rect 7045 -4059 7079 -4025
rect 7148 -4059 7182 -4025
rect 7256 -4095 7290 -4061
rect 7355 -4095 7389 -4061
rect 7454 -4095 7488 -4061
rect 7712 -4059 7746 -4025
rect 7972 -4095 8006 -4061
rect 8192 -4069 8226 -4035
rect 8312 -4069 8346 -4035
rect 8533 -4069 8567 -4035
rect 8733 -4069 8767 -4035
rect 9000 -4059 9034 -4025
rect 9260 -4095 9294 -4061
rect 9518 -4059 9552 -4025
rect 9621 -4059 9655 -4025
rect 9724 -4059 9758 -4025
rect 9832 -4095 9866 -4061
rect 9931 -4095 9965 -4061
rect 10030 -4095 10064 -4061
rect 10380 -4059 10414 -4025
rect 10640 -4095 10674 -4061
rect 10768 -4069 10802 -4035
rect 10888 -4069 10922 -4035
rect 11109 -4069 11143 -4035
rect 11309 -4069 11343 -4035
rect 11668 -4059 11702 -4025
rect 11928 -4095 11962 -4061
rect 12574 -4069 12608 -4035
rect 12642 -4069 12676 -4035
rect 12710 -4069 12744 -4035
rect 12778 -4069 12812 -4035
rect 12846 -4069 12880 -4035
rect 12914 -4069 12948 -4035
rect 13232 -4095 13266 -4061
rect 13492 -4059 13526 -4025
rect 13692 -4069 13726 -4035
rect 14119 -4069 14153 -4035
rect 14187 -4069 14221 -4035
rect 14255 -4069 14289 -4035
rect 14323 -4069 14357 -4035
rect 14391 -4069 14425 -4035
rect 14459 -4069 14493 -4035
rect 14527 -4069 14561 -4035
rect 14595 -4069 14629 -4035
rect 14663 -4069 14697 -4035
rect 14731 -4069 14765 -4035
rect 14799 -4069 14833 -4035
rect 14867 -4069 14901 -4035
rect 14935 -4069 14969 -4035
rect 15003 -4069 15037 -4035
rect 15071 -4069 15105 -4035
rect 15139 -4069 15173 -4035
rect 15682 -4095 15716 -4061
rect 15810 -4095 15844 -4061
rect 15938 -4095 15972 -4061
rect 16066 -4095 16100 -4061
rect 16174 -4059 16208 -4025
rect 16302 -4059 16336 -4025
rect 16430 -4059 16464 -4025
rect 16558 -4059 16592 -4025
rect -2902 -4667 -2868 -4633
rect -2803 -4667 -2769 -4633
rect -2704 -4667 -2670 -4633
rect -2596 -4703 -2562 -4669
rect -2493 -4703 -2459 -4669
rect -2390 -4703 -2356 -4669
rect -1522 -4703 -1488 -4669
rect -1419 -4703 -1385 -4669
rect -1316 -4703 -1282 -4669
rect -1208 -4667 -1174 -4633
rect -1109 -4667 -1075 -4633
rect -1010 -4667 -976 -4633
rect -777 -4693 -743 -4659
rect -577 -4693 -543 -4659
rect -356 -4693 -322 -4659
rect -236 -4693 -202 -4659
rect -16 -4703 18 -4669
rect 244 -4667 278 -4633
rect 511 -4693 545 -4659
rect 711 -4693 745 -4659
rect 932 -4693 966 -4659
rect 1052 -4693 1086 -4659
rect 1272 -4703 1306 -4669
rect 1532 -4667 1566 -4633
rect 1790 -4667 1824 -4633
rect 1889 -4667 1923 -4633
rect 1988 -4667 2022 -4633
rect 2096 -4703 2130 -4669
rect 2199 -4703 2233 -4669
rect 2302 -4703 2336 -4669
rect 2560 -4703 2594 -4669
rect 2820 -4667 2854 -4633
rect 3087 -4693 3121 -4659
rect 3287 -4693 3321 -4659
rect 3508 -4693 3542 -4659
rect 3628 -4693 3662 -4659
rect 3848 -4703 3882 -4669
rect 4108 -4667 4142 -4633
rect 4366 -4667 4400 -4633
rect 4465 -4667 4499 -4633
rect 4564 -4667 4598 -4633
rect 4672 -4703 4706 -4669
rect 4775 -4703 4809 -4669
rect 4878 -4703 4912 -4669
rect 5136 -4703 5170 -4669
rect 5396 -4667 5430 -4633
rect 5663 -4693 5697 -4659
rect 5863 -4693 5897 -4659
rect 6084 -4693 6118 -4659
rect 6204 -4693 6238 -4659
rect 6424 -4703 6458 -4669
rect 6684 -4667 6718 -4633
rect 6942 -4667 6976 -4633
rect 7041 -4667 7075 -4633
rect 7140 -4667 7174 -4633
rect 7248 -4703 7282 -4669
rect 7351 -4703 7385 -4669
rect 7454 -4703 7488 -4669
rect 7712 -4703 7746 -4669
rect 7972 -4667 8006 -4633
rect 8239 -4693 8273 -4659
rect 8439 -4693 8473 -4659
rect 8660 -4693 8694 -4659
rect 8780 -4693 8814 -4659
rect 9000 -4703 9034 -4669
rect 9260 -4667 9294 -4633
rect 9518 -4667 9552 -4633
rect 9617 -4667 9651 -4633
rect 9716 -4667 9750 -4633
rect 9824 -4703 9858 -4669
rect 9927 -4703 9961 -4669
rect 10030 -4703 10064 -4669
rect 10380 -4703 10414 -4669
rect 10640 -4667 10674 -4633
rect 10815 -4693 10849 -4659
rect 11015 -4693 11049 -4659
rect 11236 -4693 11270 -4659
rect 11356 -4693 11390 -4659
rect 11668 -4703 11702 -4669
rect 11928 -4667 11962 -4633
rect 13692 -4693 13726 -4659
rect 14119 -4693 14153 -4659
rect 14187 -4693 14221 -4659
rect 14255 -4693 14289 -4659
rect 14323 -4693 14357 -4659
rect 14391 -4693 14425 -4659
rect 14459 -4693 14493 -4659
rect 14527 -4693 14561 -4659
rect 14595 -4693 14629 -4659
rect 14663 -4693 14697 -4659
rect 14731 -4693 14765 -4659
rect 14799 -4693 14833 -4659
rect 14867 -4693 14901 -4659
rect 14935 -4693 14969 -4659
rect 15003 -4693 15037 -4659
rect 15071 -4693 15105 -4659
rect 15139 -4693 15173 -4659
rect 15686 -4703 15720 -4669
rect 15814 -4703 15848 -4669
rect 15942 -4703 15976 -4669
rect 16070 -4703 16104 -4669
rect 16178 -4667 16212 -4633
rect 16306 -4667 16340 -4633
rect 16434 -4667 16468 -4633
rect 16562 -4667 16596 -4633
rect -2902 -5147 -2868 -5113
rect -2799 -5147 -2765 -5113
rect -2696 -5147 -2662 -5113
rect -2588 -5183 -2554 -5149
rect -2489 -5183 -2455 -5149
rect -2390 -5183 -2356 -5149
rect -1522 -5183 -1488 -5149
rect -1423 -5183 -1389 -5149
rect -1324 -5183 -1290 -5149
rect -1216 -5147 -1182 -5113
rect -1113 -5147 -1079 -5113
rect -1010 -5147 -976 -5113
rect -786 -5183 -752 -5149
rect -687 -5183 -653 -5149
rect -588 -5183 -554 -5149
rect -480 -5147 -446 -5113
rect -377 -5147 -343 -5113
rect -274 -5147 -240 -5113
rect -16 -5147 18 -5113
rect 244 -5183 278 -5149
rect 464 -5157 498 -5123
rect 584 -5157 618 -5123
rect 805 -5157 839 -5123
rect 1005 -5157 1039 -5123
rect 1272 -5147 1306 -5113
rect 1532 -5183 1566 -5149
rect 1790 -5147 1824 -5113
rect 1893 -5147 1927 -5113
rect 1996 -5147 2030 -5113
rect 2104 -5183 2138 -5149
rect 2203 -5183 2237 -5149
rect 2302 -5183 2336 -5149
rect 2560 -5147 2594 -5113
rect 2820 -5183 2854 -5149
rect 3040 -5157 3074 -5123
rect 3160 -5157 3194 -5123
rect 3381 -5157 3415 -5123
rect 3581 -5157 3615 -5123
rect 3848 -5147 3882 -5113
rect 4108 -5183 4142 -5149
rect 4366 -5147 4400 -5113
rect 4469 -5147 4503 -5113
rect 4572 -5147 4606 -5113
rect 4680 -5183 4714 -5149
rect 4779 -5183 4813 -5149
rect 4878 -5183 4912 -5149
rect 5136 -5147 5170 -5113
rect 5396 -5183 5430 -5149
rect 5616 -5157 5650 -5123
rect 5736 -5157 5770 -5123
rect 5957 -5157 5991 -5123
rect 6157 -5157 6191 -5123
rect 6424 -5147 6458 -5113
rect 6684 -5183 6718 -5149
rect 6942 -5147 6976 -5113
rect 7045 -5147 7079 -5113
rect 7148 -5147 7182 -5113
rect 7256 -5183 7290 -5149
rect 7355 -5183 7389 -5149
rect 7454 -5183 7488 -5149
rect 7712 -5147 7746 -5113
rect 7972 -5183 8006 -5149
rect 8192 -5157 8226 -5123
rect 8312 -5157 8346 -5123
rect 8533 -5157 8567 -5123
rect 8733 -5157 8767 -5123
rect 9000 -5147 9034 -5113
rect 9260 -5183 9294 -5149
rect 9518 -5147 9552 -5113
rect 9621 -5147 9655 -5113
rect 9724 -5147 9758 -5113
rect 9832 -5183 9866 -5149
rect 9931 -5183 9965 -5149
rect 10030 -5183 10064 -5149
rect 10380 -5147 10414 -5113
rect 10640 -5183 10674 -5149
rect 10768 -5157 10802 -5123
rect 10888 -5157 10922 -5123
rect 11109 -5157 11143 -5123
rect 11309 -5157 11343 -5123
rect 11668 -5147 11702 -5113
rect 11928 -5183 11962 -5149
rect 12574 -5157 12608 -5123
rect 12642 -5157 12676 -5123
rect 12710 -5157 12744 -5123
rect 12778 -5157 12812 -5123
rect 12846 -5157 12880 -5123
rect 12914 -5157 12948 -5123
rect 13232 -5183 13266 -5149
rect 13492 -5147 13526 -5113
rect 13692 -5157 13726 -5123
rect 14119 -5157 14153 -5123
rect 14187 -5157 14221 -5123
rect 14255 -5157 14289 -5123
rect 14323 -5157 14357 -5123
rect 14391 -5157 14425 -5123
rect 14459 -5157 14493 -5123
rect 14527 -5157 14561 -5123
rect 14595 -5157 14629 -5123
rect 14663 -5157 14697 -5123
rect 14731 -5157 14765 -5123
rect 14799 -5157 14833 -5123
rect 14867 -5157 14901 -5123
rect 14935 -5157 14969 -5123
rect 15003 -5157 15037 -5123
rect 15071 -5157 15105 -5123
rect 15139 -5157 15173 -5123
rect 15682 -5183 15716 -5149
rect 15810 -5183 15844 -5149
rect 15938 -5183 15972 -5149
rect 16066 -5183 16100 -5149
rect 16174 -5147 16208 -5113
rect 16302 -5147 16336 -5113
rect 16430 -5147 16464 -5113
rect 16558 -5147 16592 -5113
rect -2902 -5755 -2868 -5721
rect -2803 -5755 -2769 -5721
rect -2704 -5755 -2670 -5721
rect -2596 -5791 -2562 -5757
rect -2493 -5791 -2459 -5757
rect -2390 -5791 -2356 -5757
rect -1522 -5791 -1488 -5757
rect -1419 -5791 -1385 -5757
rect -1316 -5791 -1282 -5757
rect -1208 -5755 -1174 -5721
rect -1109 -5755 -1075 -5721
rect -1010 -5755 -976 -5721
rect -786 -5791 -752 -5757
rect -683 -5791 -649 -5757
rect -580 -5791 -546 -5757
rect -472 -5755 -438 -5721
rect -373 -5755 -339 -5721
rect -274 -5755 -240 -5721
rect -16 -5791 18 -5757
rect 244 -5755 278 -5721
rect 511 -5781 545 -5747
rect 711 -5781 745 -5747
rect 932 -5781 966 -5747
rect 1052 -5781 1086 -5747
rect 1272 -5791 1306 -5757
rect 1532 -5755 1566 -5721
rect 1790 -5755 1824 -5721
rect 1889 -5755 1923 -5721
rect 1988 -5755 2022 -5721
rect 2096 -5791 2130 -5757
rect 2199 -5791 2233 -5757
rect 2302 -5791 2336 -5757
rect 2560 -5791 2594 -5757
rect 2820 -5755 2854 -5721
rect 3087 -5781 3121 -5747
rect 3287 -5781 3321 -5747
rect 3508 -5781 3542 -5747
rect 3628 -5781 3662 -5747
rect 3848 -5791 3882 -5757
rect 4108 -5755 4142 -5721
rect 4366 -5755 4400 -5721
rect 4465 -5755 4499 -5721
rect 4564 -5755 4598 -5721
rect 4672 -5791 4706 -5757
rect 4775 -5791 4809 -5757
rect 4878 -5791 4912 -5757
rect 5136 -5791 5170 -5757
rect 5396 -5755 5430 -5721
rect 5663 -5781 5697 -5747
rect 5863 -5781 5897 -5747
rect 6084 -5781 6118 -5747
rect 6204 -5781 6238 -5747
rect 6424 -5791 6458 -5757
rect 6684 -5755 6718 -5721
rect 6942 -5755 6976 -5721
rect 7041 -5755 7075 -5721
rect 7140 -5755 7174 -5721
rect 7248 -5791 7282 -5757
rect 7351 -5791 7385 -5757
rect 7454 -5791 7488 -5757
rect 7712 -5791 7746 -5757
rect 7972 -5755 8006 -5721
rect 8239 -5781 8273 -5747
rect 8439 -5781 8473 -5747
rect 8660 -5781 8694 -5747
rect 8780 -5781 8814 -5747
rect 9000 -5791 9034 -5757
rect 9260 -5755 9294 -5721
rect 9518 -5755 9552 -5721
rect 9617 -5755 9651 -5721
rect 9716 -5755 9750 -5721
rect 9824 -5791 9858 -5757
rect 9927 -5791 9961 -5757
rect 10030 -5791 10064 -5757
rect 10380 -5791 10414 -5757
rect 10640 -5755 10674 -5721
rect 10815 -5781 10849 -5747
rect 11015 -5781 11049 -5747
rect 11236 -5781 11270 -5747
rect 11356 -5781 11390 -5747
rect 11668 -5791 11702 -5757
rect 11928 -5755 11962 -5721
rect 13692 -5781 13726 -5747
rect 14119 -5781 14153 -5747
rect 14187 -5781 14221 -5747
rect 14255 -5781 14289 -5747
rect 14323 -5781 14357 -5747
rect 14391 -5781 14425 -5747
rect 14459 -5781 14493 -5747
rect 14527 -5781 14561 -5747
rect 14595 -5781 14629 -5747
rect 14663 -5781 14697 -5747
rect 14731 -5781 14765 -5747
rect 14799 -5781 14833 -5747
rect 14867 -5781 14901 -5747
rect 14935 -5781 14969 -5747
rect 15003 -5781 15037 -5747
rect 15071 -5781 15105 -5747
rect 15139 -5781 15173 -5747
rect 15686 -5791 15720 -5757
rect 15814 -5791 15848 -5757
rect 15942 -5791 15976 -5757
rect 16070 -5791 16104 -5757
rect 16178 -5755 16212 -5721
rect 16306 -5755 16340 -5721
rect 16434 -5755 16468 -5721
rect 16562 -5755 16596 -5721
rect -2902 -6235 -2868 -6201
rect -2799 -6235 -2765 -6201
rect -2696 -6235 -2662 -6201
rect -2588 -6271 -2554 -6237
rect -2489 -6271 -2455 -6237
rect -2390 -6271 -2356 -6237
rect -1396 -6271 -1362 -6237
rect -1136 -6235 -1102 -6201
rect -937 -6245 -903 -6211
rect -769 -6245 -735 -6211
rect -568 -6271 -534 -6237
rect -308 -6235 -274 -6201
rect -30 -6245 4 -6211
rect 38 -6245 72 -6211
rect 106 -6245 140 -6211
rect 174 -6245 208 -6211
rect 242 -6245 276 -6211
rect 310 -6245 344 -6211
rect 628 -6271 662 -6237
rect 888 -6235 922 -6201
rect 1082 -6245 1116 -6211
rect 1456 -6271 1490 -6237
rect 1716 -6235 1750 -6201
rect 1916 -6271 1950 -6237
rect 2176 -6235 2210 -6201
rect 2396 -6245 2430 -6211
rect 2516 -6245 2550 -6211
rect 2737 -6245 2771 -6211
rect 2937 -6245 2971 -6211
rect 3204 -6271 3238 -6237
rect 3464 -6235 3498 -6201
rect 4458 -6271 4492 -6237
rect 4586 -6271 4620 -6237
rect 4714 -6271 4748 -6237
rect 4842 -6271 4876 -6237
rect 4950 -6235 4984 -6201
rect 5078 -6235 5112 -6201
rect 5206 -6235 5240 -6201
rect 5334 -6235 5368 -6201
rect 6424 -6271 6458 -6237
rect 6684 -6235 6718 -6201
rect 6904 -6245 6938 -6211
rect 7024 -6245 7058 -6211
rect 7245 -6245 7279 -6211
rect 7445 -6245 7479 -6211
rect 7712 -6271 7746 -6237
rect 7972 -6235 8006 -6201
rect 8192 -6245 8226 -6211
rect 8312 -6245 8346 -6211
rect 8533 -6245 8567 -6211
rect 8733 -6245 8767 -6211
rect 9000 -6271 9034 -6237
rect 9260 -6235 9294 -6201
rect 9480 -6245 9514 -6211
rect 9600 -6245 9634 -6211
rect 9821 -6245 9855 -6211
rect 10021 -6245 10055 -6211
rect 10288 -6271 10322 -6237
rect 10548 -6235 10582 -6201
rect 10749 -6245 10783 -6211
rect 10830 -6245 10864 -6211
rect 10914 -6245 10948 -6211
rect 10998 -6245 11032 -6211
rect 11250 -6245 11284 -6211
rect 11334 -6245 11368 -6211
rect 11668 -6271 11702 -6237
rect 11928 -6235 11962 -6201
rect 13658 -6271 13692 -6237
rect 13786 -6271 13820 -6237
rect 13914 -6271 13948 -6237
rect 14042 -6271 14076 -6237
rect 14150 -6235 14184 -6201
rect 14278 -6235 14312 -6201
rect 14406 -6235 14440 -6201
rect 14534 -6235 14568 -6201
rect 14854 -6271 14888 -6237
rect 14982 -6271 15016 -6237
rect 15110 -6271 15144 -6237
rect 15238 -6271 15272 -6237
rect 15346 -6235 15380 -6201
rect 15474 -6235 15508 -6201
rect 15602 -6235 15636 -6201
rect 15730 -6235 15764 -6201
rect 16050 -6271 16084 -6237
rect 16149 -6271 16183 -6237
rect 16248 -6271 16282 -6237
rect 16356 -6235 16390 -6201
rect 16459 -6235 16493 -6201
rect 16562 -6235 16596 -6201
rect -2930 -6843 -2896 -6809
rect -2822 -6883 -2788 -6849
rect -2597 -6869 -2563 -6835
rect -2333 -6801 -2299 -6767
rect -2081 -6753 -2047 -6719
rect -2495 -6854 -2461 -6820
rect -2190 -6831 -2156 -6797
rect -2170 -6927 -2136 -6893
rect -1669 -6753 -1635 -6719
rect -1533 -6753 -1499 -6719
rect -1907 -6819 -1873 -6785
rect -1771 -6819 -1737 -6785
rect -1971 -6915 -1937 -6881
rect -1728 -6927 -1694 -6893
rect -1459 -6869 -1425 -6835
rect -1275 -6869 -1241 -6835
rect -1014 -6869 -980 -6835
rect -786 -6879 -752 -6845
rect -683 -6879 -649 -6845
rect -580 -6879 -546 -6845
rect -472 -6843 -438 -6809
rect -373 -6843 -339 -6809
rect -274 -6843 -240 -6809
rect 42 -6879 76 -6845
rect 145 -6879 179 -6845
rect 248 -6879 282 -6845
rect 356 -6843 390 -6809
rect 455 -6843 489 -6809
rect 554 -6843 588 -6809
rect 778 -6879 812 -6845
rect 881 -6879 915 -6845
rect 984 -6879 1018 -6845
rect 1092 -6843 1126 -6809
rect 1191 -6843 1225 -6809
rect 1290 -6843 1324 -6809
rect 1606 -6879 1640 -6845
rect 1709 -6879 1743 -6845
rect 1812 -6879 1846 -6845
rect 1920 -6843 1954 -6809
rect 2019 -6843 2053 -6809
rect 2118 -6843 2152 -6809
rect 2342 -6879 2376 -6845
rect 2445 -6879 2479 -6845
rect 2548 -6879 2582 -6845
rect 2656 -6843 2690 -6809
rect 2755 -6843 2789 -6809
rect 2854 -6843 2888 -6809
rect 3170 -6879 3204 -6845
rect 3273 -6879 3307 -6845
rect 3376 -6879 3410 -6845
rect 3484 -6843 3518 -6809
rect 3583 -6843 3617 -6809
rect 3682 -6843 3716 -6809
rect 3906 -6879 3940 -6845
rect 4009 -6879 4043 -6845
rect 4112 -6879 4146 -6845
rect 4220 -6843 4254 -6809
rect 4319 -6843 4353 -6809
rect 4418 -6843 4452 -6809
rect 4734 -6879 4768 -6845
rect 4837 -6879 4871 -6845
rect 4940 -6879 4974 -6845
rect 5048 -6843 5082 -6809
rect 5147 -6843 5181 -6809
rect 5246 -6843 5280 -6809
rect 5470 -6879 5504 -6845
rect 5573 -6879 5607 -6845
rect 5676 -6879 5710 -6845
rect 5784 -6843 5818 -6809
rect 5883 -6843 5917 -6809
rect 5982 -6843 6016 -6809
rect 6298 -6879 6332 -6845
rect 6401 -6879 6435 -6845
rect 6504 -6879 6538 -6845
rect 6612 -6843 6646 -6809
rect 6711 -6843 6745 -6809
rect 6810 -6843 6844 -6809
rect 7034 -6879 7068 -6845
rect 7137 -6879 7171 -6845
rect 7240 -6879 7274 -6845
rect 7348 -6843 7382 -6809
rect 7447 -6843 7481 -6809
rect 7546 -6843 7580 -6809
rect 7862 -6879 7896 -6845
rect 7965 -6879 7999 -6845
rect 8068 -6879 8102 -6845
rect 8176 -6843 8210 -6809
rect 8275 -6843 8309 -6809
rect 8374 -6843 8408 -6809
rect 8598 -6879 8632 -6845
rect 8701 -6879 8735 -6845
rect 8804 -6879 8838 -6845
rect 8912 -6843 8946 -6809
rect 9011 -6843 9045 -6809
rect 9110 -6843 9144 -6809
rect 16050 -6879 16084 -6845
rect 16153 -6879 16187 -6845
rect 16256 -6879 16290 -6845
rect 16364 -6843 16398 -6809
rect 16463 -6843 16497 -6809
rect 16562 -6843 16596 -6809
rect -2902 -7323 -2868 -7289
rect -2799 -7323 -2765 -7289
rect -2696 -7323 -2662 -7289
rect -2588 -7359 -2554 -7325
rect -2489 -7359 -2455 -7325
rect -2390 -7359 -2356 -7325
rect -1522 -7359 -1488 -7325
rect -1423 -7359 -1389 -7325
rect -1324 -7359 -1290 -7325
rect -1216 -7323 -1182 -7289
rect -1113 -7323 -1079 -7289
rect -1010 -7323 -976 -7289
rect -786 -7359 -752 -7325
rect -687 -7359 -653 -7325
rect -588 -7359 -554 -7325
rect -480 -7323 -446 -7289
rect -377 -7323 -343 -7289
rect -274 -7323 -240 -7289
rect 42 -7359 76 -7325
rect 141 -7359 175 -7325
rect 240 -7359 274 -7325
rect 348 -7323 382 -7289
rect 451 -7323 485 -7289
rect 554 -7323 588 -7289
rect 778 -7359 812 -7325
rect 877 -7359 911 -7325
rect 976 -7359 1010 -7325
rect 1084 -7323 1118 -7289
rect 1187 -7323 1221 -7289
rect 1290 -7323 1324 -7289
rect 1606 -7359 1640 -7325
rect 1705 -7359 1739 -7325
rect 1804 -7359 1838 -7325
rect 1912 -7323 1946 -7289
rect 2015 -7323 2049 -7289
rect 2118 -7323 2152 -7289
rect 2284 -7323 2318 -7289
rect 2544 -7359 2578 -7325
rect 3102 -7333 3136 -7299
rect 3296 -7323 3330 -7289
rect 3556 -7359 3590 -7325
rect 3755 -7333 3789 -7299
rect 3923 -7333 3957 -7299
rect 4124 -7323 4158 -7289
rect 4384 -7359 4418 -7325
rect 4633 -7333 4667 -7299
rect 4729 -7333 4763 -7299
rect 4870 -7297 4904 -7263
rect 4966 -7297 5000 -7263
rect 5128 -7297 5162 -7263
rect 5038 -7410 5072 -7376
rect 5504 -7323 5538 -7289
rect 5206 -7410 5240 -7376
rect 5764 -7359 5798 -7325
rect 6026 -7333 6060 -7299
rect 6287 -7333 6321 -7299
rect 6471 -7333 6505 -7299
rect 6740 -7275 6774 -7241
rect 6983 -7287 7017 -7253
rect 6783 -7383 6817 -7349
rect 6919 -7383 6953 -7349
rect 6545 -7449 6579 -7415
rect 6681 -7449 6715 -7415
rect 7182 -7275 7216 -7241
rect 7202 -7371 7236 -7337
rect 7507 -7348 7541 -7314
rect 7093 -7449 7127 -7415
rect 7345 -7401 7379 -7367
rect 7609 -7333 7643 -7299
rect 7862 -7359 7896 -7325
rect 7961 -7359 7995 -7325
rect 8060 -7359 8094 -7325
rect 8168 -7323 8202 -7289
rect 8271 -7323 8305 -7289
rect 8374 -7323 8408 -7289
rect 8598 -7359 8632 -7325
rect 8697 -7359 8731 -7325
rect 8796 -7359 8830 -7325
rect 8904 -7323 8938 -7289
rect 9007 -7323 9041 -7289
rect 9110 -7323 9144 -7289
rect 16050 -7359 16084 -7325
rect 16149 -7359 16183 -7325
rect 16248 -7359 16282 -7325
rect 16356 -7323 16390 -7289
rect 16459 -7323 16493 -7289
rect 16562 -7323 16596 -7289
rect -2902 -7931 -2868 -7897
rect -2803 -7931 -2769 -7897
rect -2704 -7931 -2670 -7897
rect -2596 -7967 -2562 -7933
rect -2493 -7967 -2459 -7933
rect -2390 -7967 -2356 -7933
rect -1396 -7931 -1362 -7897
rect -1136 -7967 -1102 -7933
rect -937 -7957 -903 -7923
rect -769 -7957 -735 -7923
rect -568 -7931 -534 -7897
rect -308 -7967 -274 -7933
rect -30 -7957 4 -7923
rect 38 -7957 72 -7923
rect 106 -7957 140 -7923
rect 174 -7957 208 -7923
rect 242 -7957 276 -7923
rect 310 -7957 344 -7923
rect 628 -7931 662 -7897
rect 888 -7967 922 -7933
rect 1082 -7957 1116 -7923
rect 1456 -7931 1490 -7897
rect 1716 -7967 1750 -7933
rect 1916 -7931 1950 -7897
rect 2176 -7967 2210 -7933
rect 2396 -7957 2430 -7923
rect 2516 -7957 2550 -7923
rect 2737 -7957 2771 -7923
rect 2937 -7957 2971 -7923
rect 3204 -7931 3238 -7897
rect 3464 -7967 3498 -7933
rect 4458 -7931 4492 -7897
rect 4586 -7931 4620 -7897
rect 4714 -7931 4748 -7897
rect 4842 -7931 4876 -7897
rect 4950 -7967 4984 -7933
rect 5078 -7967 5112 -7933
rect 5206 -7967 5240 -7933
rect 5334 -7967 5368 -7933
rect 6424 -7931 6458 -7897
rect 6684 -7967 6718 -7933
rect 6904 -7957 6938 -7923
rect 7024 -7957 7058 -7923
rect 7245 -7957 7279 -7923
rect 7445 -7957 7479 -7923
rect 7712 -7931 7746 -7897
rect 7972 -7967 8006 -7933
rect 8192 -7957 8226 -7923
rect 8312 -7957 8346 -7923
rect 8533 -7957 8567 -7923
rect 8733 -7957 8767 -7923
rect 9000 -7931 9034 -7897
rect 9260 -7967 9294 -7933
rect 9480 -7957 9514 -7923
rect 9600 -7957 9634 -7923
rect 9821 -7957 9855 -7923
rect 10021 -7957 10055 -7923
rect 10288 -7931 10322 -7897
rect 10548 -7967 10582 -7933
rect 10749 -7957 10783 -7923
rect 10830 -7957 10864 -7923
rect 10914 -7957 10948 -7923
rect 10998 -7957 11032 -7923
rect 11250 -7957 11284 -7923
rect 11334 -7957 11368 -7923
rect 11668 -7931 11702 -7897
rect 11928 -7967 11962 -7933
rect 13658 -7931 13692 -7897
rect 13786 -7931 13820 -7897
rect 13914 -7931 13948 -7897
rect 14042 -7931 14076 -7897
rect 14150 -7967 14184 -7933
rect 14278 -7967 14312 -7933
rect 14406 -7967 14440 -7933
rect 14534 -7967 14568 -7933
rect 14854 -7931 14888 -7897
rect 14982 -7931 15016 -7897
rect 15110 -7931 15144 -7897
rect 15238 -7931 15272 -7897
rect 15346 -7967 15380 -7933
rect 15474 -7967 15508 -7933
rect 15602 -7967 15636 -7933
rect 15730 -7967 15764 -7933
rect 16050 -7931 16084 -7897
rect 16149 -7931 16183 -7897
rect 16248 -7931 16282 -7897
rect 16356 -7967 16390 -7933
rect 16459 -7967 16493 -7933
rect 16562 -7967 16596 -7933
rect -2902 -8411 -2868 -8377
rect -2799 -8411 -2765 -8377
rect -2696 -8411 -2662 -8377
rect -2588 -8447 -2554 -8413
rect -2489 -8447 -2455 -8413
rect -2390 -8447 -2356 -8413
rect -1522 -8411 -1488 -8377
rect -1419 -8411 -1385 -8377
rect -1316 -8411 -1282 -8377
rect -1208 -8447 -1174 -8413
rect -1109 -8447 -1075 -8413
rect -1010 -8447 -976 -8413
rect -786 -8411 -752 -8377
rect -683 -8411 -649 -8377
rect -580 -8411 -546 -8377
rect -472 -8447 -438 -8413
rect -373 -8447 -339 -8413
rect -274 -8447 -240 -8413
rect -16 -8411 18 -8377
rect 244 -8447 278 -8413
rect 511 -8421 545 -8387
rect 711 -8421 745 -8387
rect 932 -8421 966 -8387
rect 1052 -8421 1086 -8387
rect 1272 -8411 1306 -8377
rect 1532 -8447 1566 -8413
rect 1790 -8411 1824 -8377
rect 1893 -8411 1927 -8377
rect 1996 -8411 2030 -8377
rect 2104 -8447 2138 -8413
rect 2203 -8447 2237 -8413
rect 2302 -8447 2336 -8413
rect 2560 -8411 2594 -8377
rect 2820 -8447 2854 -8413
rect 3087 -8421 3121 -8387
rect 3287 -8421 3321 -8387
rect 3508 -8421 3542 -8387
rect 3628 -8421 3662 -8387
rect 3848 -8411 3882 -8377
rect 4108 -8447 4142 -8413
rect 4366 -8411 4400 -8377
rect 4469 -8411 4503 -8377
rect 4572 -8411 4606 -8377
rect 4680 -8447 4714 -8413
rect 4779 -8447 4813 -8413
rect 4878 -8447 4912 -8413
rect 5136 -8411 5170 -8377
rect 5396 -8447 5430 -8413
rect 5663 -8421 5697 -8387
rect 5863 -8421 5897 -8387
rect 6084 -8421 6118 -8387
rect 6204 -8421 6238 -8387
rect 6424 -8411 6458 -8377
rect 6684 -8447 6718 -8413
rect 6942 -8411 6976 -8377
rect 7045 -8411 7079 -8377
rect 7148 -8411 7182 -8377
rect 7256 -8447 7290 -8413
rect 7355 -8447 7389 -8413
rect 7454 -8447 7488 -8413
rect 7712 -8411 7746 -8377
rect 7972 -8447 8006 -8413
rect 8239 -8421 8273 -8387
rect 8439 -8421 8473 -8387
rect 8660 -8421 8694 -8387
rect 8780 -8421 8814 -8387
rect 9000 -8411 9034 -8377
rect 9260 -8447 9294 -8413
rect 9518 -8411 9552 -8377
rect 9621 -8411 9655 -8377
rect 9724 -8411 9758 -8377
rect 9832 -8447 9866 -8413
rect 9931 -8447 9965 -8413
rect 10030 -8447 10064 -8413
rect 10380 -8411 10414 -8377
rect 10640 -8447 10674 -8413
rect 10815 -8421 10849 -8387
rect 11015 -8421 11049 -8387
rect 11236 -8421 11270 -8387
rect 11356 -8421 11390 -8387
rect 11668 -8411 11702 -8377
rect 11928 -8447 11962 -8413
rect 13692 -8421 13726 -8387
rect 14119 -8421 14153 -8387
rect 14187 -8421 14221 -8387
rect 14255 -8421 14289 -8387
rect 14323 -8421 14357 -8387
rect 14391 -8421 14425 -8387
rect 14459 -8421 14493 -8387
rect 14527 -8421 14561 -8387
rect 14595 -8421 14629 -8387
rect 14663 -8421 14697 -8387
rect 14731 -8421 14765 -8387
rect 14799 -8421 14833 -8387
rect 14867 -8421 14901 -8387
rect 14935 -8421 14969 -8387
rect 15003 -8421 15037 -8387
rect 15071 -8421 15105 -8387
rect 15139 -8421 15173 -8387
rect 15686 -8411 15720 -8377
rect 15814 -8411 15848 -8377
rect 15942 -8411 15976 -8377
rect 16070 -8411 16104 -8377
rect 16178 -8447 16212 -8413
rect 16306 -8447 16340 -8413
rect 16434 -8447 16468 -8413
rect 16562 -8447 16596 -8413
rect -2902 -9019 -2868 -8985
rect -2803 -9019 -2769 -8985
rect -2704 -9019 -2670 -8985
rect -2596 -9055 -2562 -9021
rect -2493 -9055 -2459 -9021
rect -2390 -9055 -2356 -9021
rect -1522 -9019 -1488 -8985
rect -1423 -9019 -1389 -8985
rect -1324 -9019 -1290 -8985
rect -1216 -9055 -1182 -9021
rect -1113 -9055 -1079 -9021
rect -1010 -9055 -976 -9021
rect -786 -9019 -752 -8985
rect -687 -9019 -653 -8985
rect -588 -9019 -554 -8985
rect -480 -9055 -446 -9021
rect -377 -9055 -343 -9021
rect -274 -9055 -240 -9021
rect -16 -9055 18 -9021
rect 244 -9019 278 -8985
rect 464 -9045 498 -9011
rect 584 -9045 618 -9011
rect 805 -9045 839 -9011
rect 1005 -9045 1039 -9011
rect 1272 -9055 1306 -9021
rect 1532 -9019 1566 -8985
rect 1790 -9019 1824 -8985
rect 1889 -9019 1923 -8985
rect 1988 -9019 2022 -8985
rect 2096 -9055 2130 -9021
rect 2199 -9055 2233 -9021
rect 2302 -9055 2336 -9021
rect 2560 -9055 2594 -9021
rect 2820 -9019 2854 -8985
rect 3040 -9045 3074 -9011
rect 3160 -9045 3194 -9011
rect 3381 -9045 3415 -9011
rect 3581 -9045 3615 -9011
rect 3848 -9055 3882 -9021
rect 4108 -9019 4142 -8985
rect 4366 -9019 4400 -8985
rect 4465 -9019 4499 -8985
rect 4564 -9019 4598 -8985
rect 4672 -9055 4706 -9021
rect 4775 -9055 4809 -9021
rect 4878 -9055 4912 -9021
rect 5136 -9055 5170 -9021
rect 5396 -9019 5430 -8985
rect 5616 -9045 5650 -9011
rect 5736 -9045 5770 -9011
rect 5957 -9045 5991 -9011
rect 6157 -9045 6191 -9011
rect 6424 -9055 6458 -9021
rect 6684 -9019 6718 -8985
rect 6942 -9019 6976 -8985
rect 7041 -9019 7075 -8985
rect 7140 -9019 7174 -8985
rect 7248 -9055 7282 -9021
rect 7351 -9055 7385 -9021
rect 7454 -9055 7488 -9021
rect 7712 -9055 7746 -9021
rect 7972 -9019 8006 -8985
rect 8192 -9045 8226 -9011
rect 8312 -9045 8346 -9011
rect 8533 -9045 8567 -9011
rect 8733 -9045 8767 -9011
rect 9000 -9055 9034 -9021
rect 9260 -9019 9294 -8985
rect 9518 -9019 9552 -8985
rect 9617 -9019 9651 -8985
rect 9716 -9019 9750 -8985
rect 9824 -9055 9858 -9021
rect 9927 -9055 9961 -9021
rect 10030 -9055 10064 -9021
rect 10380 -9055 10414 -9021
rect 10640 -9019 10674 -8985
rect 10768 -9045 10802 -9011
rect 10888 -9045 10922 -9011
rect 11109 -9045 11143 -9011
rect 11309 -9045 11343 -9011
rect 11668 -9055 11702 -9021
rect 11928 -9019 11962 -8985
rect 12574 -9045 12608 -9011
rect 12642 -9045 12676 -9011
rect 12710 -9045 12744 -9011
rect 12778 -9045 12812 -9011
rect 12846 -9045 12880 -9011
rect 12914 -9045 12948 -9011
rect 13232 -9019 13266 -8985
rect 13492 -9055 13526 -9021
rect 13692 -9045 13726 -9011
rect 14119 -9045 14153 -9011
rect 14187 -9045 14221 -9011
rect 14255 -9045 14289 -9011
rect 14323 -9045 14357 -9011
rect 14391 -9045 14425 -9011
rect 14459 -9045 14493 -9011
rect 14527 -9045 14561 -9011
rect 14595 -9045 14629 -9011
rect 14663 -9045 14697 -9011
rect 14731 -9045 14765 -9011
rect 14799 -9045 14833 -9011
rect 14867 -9045 14901 -9011
rect 14935 -9045 14969 -9011
rect 15003 -9045 15037 -9011
rect 15071 -9045 15105 -9011
rect 15139 -9045 15173 -9011
rect 15682 -9019 15716 -8985
rect 15810 -9019 15844 -8985
rect 15938 -9019 15972 -8985
rect 16066 -9019 16100 -8985
rect 16174 -9055 16208 -9021
rect 16302 -9055 16336 -9021
rect 16430 -9055 16464 -9021
rect 16558 -9055 16592 -9021
rect -2902 -9499 -2868 -9465
rect -2799 -9499 -2765 -9465
rect -2696 -9499 -2662 -9465
rect -2588 -9535 -2554 -9501
rect -2489 -9535 -2455 -9501
rect -2390 -9535 -2356 -9501
rect -1522 -9499 -1488 -9465
rect -1419 -9499 -1385 -9465
rect -1316 -9499 -1282 -9465
rect -1208 -9535 -1174 -9501
rect -1109 -9535 -1075 -9501
rect -1010 -9535 -976 -9501
rect -777 -9509 -743 -9475
rect -577 -9509 -543 -9475
rect -356 -9509 -322 -9475
rect -236 -9509 -202 -9475
rect -16 -9499 18 -9465
rect 244 -9535 278 -9501
rect 511 -9509 545 -9475
rect 711 -9509 745 -9475
rect 932 -9509 966 -9475
rect 1052 -9509 1086 -9475
rect 1272 -9499 1306 -9465
rect 1532 -9535 1566 -9501
rect 1790 -9499 1824 -9465
rect 1893 -9499 1927 -9465
rect 1996 -9499 2030 -9465
rect 2104 -9535 2138 -9501
rect 2203 -9535 2237 -9501
rect 2302 -9535 2336 -9501
rect 2560 -9499 2594 -9465
rect 2820 -9535 2854 -9501
rect 3087 -9509 3121 -9475
rect 3287 -9509 3321 -9475
rect 3508 -9509 3542 -9475
rect 3628 -9509 3662 -9475
rect 3848 -9499 3882 -9465
rect 4108 -9535 4142 -9501
rect 4366 -9499 4400 -9465
rect 4469 -9499 4503 -9465
rect 4572 -9499 4606 -9465
rect 4680 -9535 4714 -9501
rect 4779 -9535 4813 -9501
rect 4878 -9535 4912 -9501
rect 5136 -9499 5170 -9465
rect 5396 -9535 5430 -9501
rect 5663 -9509 5697 -9475
rect 5863 -9509 5897 -9475
rect 6084 -9509 6118 -9475
rect 6204 -9509 6238 -9475
rect 6424 -9499 6458 -9465
rect 6684 -9535 6718 -9501
rect 6942 -9499 6976 -9465
rect 7045 -9499 7079 -9465
rect 7148 -9499 7182 -9465
rect 7256 -9535 7290 -9501
rect 7355 -9535 7389 -9501
rect 7454 -9535 7488 -9501
rect 7712 -9499 7746 -9465
rect 7972 -9535 8006 -9501
rect 8239 -9509 8273 -9475
rect 8439 -9509 8473 -9475
rect 8660 -9509 8694 -9475
rect 8780 -9509 8814 -9475
rect 9000 -9499 9034 -9465
rect 9260 -9535 9294 -9501
rect 9518 -9499 9552 -9465
rect 9621 -9499 9655 -9465
rect 9724 -9499 9758 -9465
rect 9832 -9535 9866 -9501
rect 9931 -9535 9965 -9501
rect 10030 -9535 10064 -9501
rect 10380 -9499 10414 -9465
rect 10640 -9535 10674 -9501
rect 10815 -9509 10849 -9475
rect 11015 -9509 11049 -9475
rect 11236 -9509 11270 -9475
rect 11356 -9509 11390 -9475
rect 11668 -9499 11702 -9465
rect 11928 -9535 11962 -9501
rect 13692 -9509 13726 -9475
rect 14119 -9509 14153 -9475
rect 14187 -9509 14221 -9475
rect 14255 -9509 14289 -9475
rect 14323 -9509 14357 -9475
rect 14391 -9509 14425 -9475
rect 14459 -9509 14493 -9475
rect 14527 -9509 14561 -9475
rect 14595 -9509 14629 -9475
rect 14663 -9509 14697 -9475
rect 14731 -9509 14765 -9475
rect 14799 -9509 14833 -9475
rect 14867 -9509 14901 -9475
rect 14935 -9509 14969 -9475
rect 15003 -9509 15037 -9475
rect 15071 -9509 15105 -9475
rect 15139 -9509 15173 -9475
rect 15686 -9499 15720 -9465
rect 15814 -9499 15848 -9465
rect 15942 -9499 15976 -9465
rect 16070 -9499 16104 -9465
rect 16178 -9535 16212 -9501
rect 16306 -9535 16340 -9501
rect 16434 -9535 16468 -9501
rect 16562 -9535 16596 -9501
rect -2902 -10107 -2868 -10073
rect -2803 -10107 -2769 -10073
rect -2704 -10107 -2670 -10073
rect -2596 -10143 -2562 -10109
rect -2493 -10143 -2459 -10109
rect -2390 -10143 -2356 -10109
rect -1522 -10107 -1488 -10073
rect -1423 -10107 -1389 -10073
rect -1324 -10107 -1290 -10073
rect -1216 -10143 -1182 -10109
rect -1113 -10143 -1079 -10109
rect -1010 -10143 -976 -10109
rect -786 -10107 -752 -10073
rect -687 -10107 -653 -10073
rect -588 -10107 -554 -10073
rect -480 -10143 -446 -10109
rect -377 -10143 -343 -10109
rect -274 -10143 -240 -10109
rect -16 -10143 18 -10109
rect 244 -10107 278 -10073
rect 464 -10133 498 -10099
rect 584 -10133 618 -10099
rect 805 -10133 839 -10099
rect 1005 -10133 1039 -10099
rect 1272 -10143 1306 -10109
rect 1532 -10107 1566 -10073
rect 1790 -10107 1824 -10073
rect 1889 -10107 1923 -10073
rect 1988 -10107 2022 -10073
rect 2096 -10143 2130 -10109
rect 2199 -10143 2233 -10109
rect 2302 -10143 2336 -10109
rect 2560 -10143 2594 -10109
rect 2820 -10107 2854 -10073
rect 3040 -10133 3074 -10099
rect 3160 -10133 3194 -10099
rect 3381 -10133 3415 -10099
rect 3581 -10133 3615 -10099
rect 3848 -10143 3882 -10109
rect 4108 -10107 4142 -10073
rect 4366 -10107 4400 -10073
rect 4465 -10107 4499 -10073
rect 4564 -10107 4598 -10073
rect 4672 -10143 4706 -10109
rect 4775 -10143 4809 -10109
rect 4878 -10143 4912 -10109
rect 5136 -10143 5170 -10109
rect 5396 -10107 5430 -10073
rect 5616 -10133 5650 -10099
rect 5736 -10133 5770 -10099
rect 5957 -10133 5991 -10099
rect 6157 -10133 6191 -10099
rect 6424 -10143 6458 -10109
rect 6684 -10107 6718 -10073
rect 6942 -10107 6976 -10073
rect 7041 -10107 7075 -10073
rect 7140 -10107 7174 -10073
rect 7248 -10143 7282 -10109
rect 7351 -10143 7385 -10109
rect 7454 -10143 7488 -10109
rect 7712 -10143 7746 -10109
rect 7972 -10107 8006 -10073
rect 8192 -10133 8226 -10099
rect 8312 -10133 8346 -10099
rect 8533 -10133 8567 -10099
rect 8733 -10133 8767 -10099
rect 9000 -10143 9034 -10109
rect 9260 -10107 9294 -10073
rect 9518 -10107 9552 -10073
rect 9617 -10107 9651 -10073
rect 9716 -10107 9750 -10073
rect 9824 -10143 9858 -10109
rect 9927 -10143 9961 -10109
rect 10030 -10143 10064 -10109
rect 10380 -10143 10414 -10109
rect 10640 -10107 10674 -10073
rect 10768 -10133 10802 -10099
rect 10888 -10133 10922 -10099
rect 11109 -10133 11143 -10099
rect 11309 -10133 11343 -10099
rect 11668 -10143 11702 -10109
rect 11928 -10107 11962 -10073
rect 12574 -10133 12608 -10099
rect 12642 -10133 12676 -10099
rect 12710 -10133 12744 -10099
rect 12778 -10133 12812 -10099
rect 12846 -10133 12880 -10099
rect 12914 -10133 12948 -10099
rect 13232 -10107 13266 -10073
rect 13492 -10143 13526 -10109
rect 13692 -10133 13726 -10099
rect 14119 -10133 14153 -10099
rect 14187 -10133 14221 -10099
rect 14255 -10133 14289 -10099
rect 14323 -10133 14357 -10099
rect 14391 -10133 14425 -10099
rect 14459 -10133 14493 -10099
rect 14527 -10133 14561 -10099
rect 14595 -10133 14629 -10099
rect 14663 -10133 14697 -10099
rect 14731 -10133 14765 -10099
rect 14799 -10133 14833 -10099
rect 14867 -10133 14901 -10099
rect 14935 -10133 14969 -10099
rect 15003 -10133 15037 -10099
rect 15071 -10133 15105 -10099
rect 15139 -10133 15173 -10099
rect 15682 -10107 15716 -10073
rect 15810 -10107 15844 -10073
rect 15938 -10107 15972 -10073
rect 16066 -10107 16100 -10073
rect 16174 -10143 16208 -10109
rect 16302 -10143 16336 -10109
rect 16430 -10143 16464 -10109
rect 16558 -10143 16592 -10109
rect -2902 -10587 -2868 -10553
rect -2799 -10587 -2765 -10553
rect -2696 -10587 -2662 -10553
rect -2588 -10623 -2554 -10589
rect -2489 -10623 -2455 -10589
rect -2390 -10623 -2356 -10589
rect -1954 -10597 -1920 -10563
rect -1522 -10587 -1488 -10553
rect -1419 -10587 -1385 -10553
rect -1316 -10587 -1282 -10553
rect -1208 -10623 -1174 -10589
rect -1109 -10623 -1075 -10589
rect -1010 -10623 -976 -10589
rect -786 -10587 -752 -10553
rect -683 -10587 -649 -10553
rect -580 -10587 -546 -10553
rect -472 -10623 -438 -10589
rect -373 -10623 -339 -10589
rect -274 -10623 -240 -10589
rect -16 -10587 18 -10553
rect 244 -10623 278 -10589
rect 511 -10597 545 -10563
rect 711 -10597 745 -10563
rect 932 -10597 966 -10563
rect 1052 -10597 1086 -10563
rect 1272 -10587 1306 -10553
rect 1532 -10623 1566 -10589
rect 1790 -10587 1824 -10553
rect 1893 -10587 1927 -10553
rect 1996 -10587 2030 -10553
rect 2104 -10623 2138 -10589
rect 2203 -10623 2237 -10589
rect 2302 -10623 2336 -10589
rect 2560 -10587 2594 -10553
rect 2820 -10623 2854 -10589
rect 3087 -10597 3121 -10563
rect 3287 -10597 3321 -10563
rect 3508 -10597 3542 -10563
rect 3628 -10597 3662 -10563
rect 3848 -10587 3882 -10553
rect 4108 -10623 4142 -10589
rect 4366 -10587 4400 -10553
rect 4469 -10587 4503 -10553
rect 4572 -10587 4606 -10553
rect 4680 -10623 4714 -10589
rect 4779 -10623 4813 -10589
rect 4878 -10623 4912 -10589
rect 5136 -10587 5170 -10553
rect 5396 -10623 5430 -10589
rect 5663 -10597 5697 -10563
rect 5863 -10597 5897 -10563
rect 6084 -10597 6118 -10563
rect 6204 -10597 6238 -10563
rect 6424 -10587 6458 -10553
rect 6684 -10623 6718 -10589
rect 6942 -10587 6976 -10553
rect 7045 -10587 7079 -10553
rect 7148 -10587 7182 -10553
rect 7256 -10623 7290 -10589
rect 7355 -10623 7389 -10589
rect 7454 -10623 7488 -10589
rect 7712 -10587 7746 -10553
rect 7972 -10623 8006 -10589
rect 8239 -10597 8273 -10563
rect 8439 -10597 8473 -10563
rect 8660 -10597 8694 -10563
rect 8780 -10597 8814 -10563
rect 9000 -10587 9034 -10553
rect 9260 -10623 9294 -10589
rect 9518 -10587 9552 -10553
rect 9621 -10587 9655 -10553
rect 9724 -10587 9758 -10553
rect 9832 -10623 9866 -10589
rect 9931 -10623 9965 -10589
rect 10030 -10623 10064 -10589
rect 10380 -10587 10414 -10553
rect 10640 -10623 10674 -10589
rect 10815 -10597 10849 -10563
rect 11015 -10597 11049 -10563
rect 11236 -10597 11270 -10563
rect 11356 -10597 11390 -10563
rect 11668 -10587 11702 -10553
rect 11928 -10623 11962 -10589
rect 13662 -10587 13696 -10553
rect 13790 -10587 13824 -10553
rect 13918 -10587 13952 -10553
rect 14046 -10587 14080 -10553
rect 14154 -10623 14188 -10589
rect 14282 -10623 14316 -10589
rect 14410 -10623 14444 -10589
rect 14538 -10623 14572 -10589
rect 14858 -10587 14892 -10553
rect 14986 -10587 15020 -10553
rect 15114 -10587 15148 -10553
rect 15242 -10587 15276 -10553
rect 15350 -10623 15384 -10589
rect 15478 -10623 15512 -10589
rect 15606 -10623 15640 -10589
rect 15734 -10623 15768 -10589
rect 16050 -10587 16084 -10553
rect 16153 -10587 16187 -10553
rect 16256 -10587 16290 -10553
rect 16364 -10623 16398 -10589
rect 16463 -10623 16497 -10589
rect 16562 -10623 16596 -10589
rect -2902 -11195 -2868 -11161
rect -2803 -11195 -2769 -11161
rect -2704 -11195 -2670 -11161
rect -2596 -11231 -2562 -11197
rect -2493 -11231 -2459 -11197
rect -2390 -11231 -2356 -11197
rect -1522 -11231 -1488 -11197
rect -1419 -11231 -1385 -11197
rect -1316 -11231 -1282 -11197
rect -1208 -11195 -1174 -11161
rect -1109 -11195 -1075 -11161
rect -1010 -11195 -976 -11161
rect -786 -11231 -752 -11197
rect -683 -11231 -649 -11197
rect -580 -11231 -546 -11197
rect -472 -11195 -438 -11161
rect -373 -11195 -339 -11161
rect -274 -11195 -240 -11161
rect -16 -11231 18 -11197
rect 244 -11195 278 -11161
rect 511 -11221 545 -11187
rect 711 -11221 745 -11187
rect 932 -11221 966 -11187
rect 1052 -11221 1086 -11187
rect 1272 -11231 1306 -11197
rect 1532 -11195 1566 -11161
rect 1790 -11195 1824 -11161
rect 1889 -11195 1923 -11161
rect 1988 -11195 2022 -11161
rect 2096 -11231 2130 -11197
rect 2199 -11231 2233 -11197
rect 2302 -11231 2336 -11197
rect 2560 -11231 2594 -11197
rect 2820 -11195 2854 -11161
rect 3087 -11221 3121 -11187
rect 3287 -11221 3321 -11187
rect 3508 -11221 3542 -11187
rect 3628 -11221 3662 -11187
rect 3848 -11231 3882 -11197
rect 4108 -11195 4142 -11161
rect 4366 -11195 4400 -11161
rect 4465 -11195 4499 -11161
rect 4564 -11195 4598 -11161
rect 4672 -11231 4706 -11197
rect 4775 -11231 4809 -11197
rect 4878 -11231 4912 -11197
rect 5136 -11231 5170 -11197
rect 5396 -11195 5430 -11161
rect 5663 -11221 5697 -11187
rect 5863 -11221 5897 -11187
rect 6084 -11221 6118 -11187
rect 6204 -11221 6238 -11187
rect 6424 -11231 6458 -11197
rect 6684 -11195 6718 -11161
rect 6942 -11195 6976 -11161
rect 7041 -11195 7075 -11161
rect 7140 -11195 7174 -11161
rect 7248 -11231 7282 -11197
rect 7351 -11231 7385 -11197
rect 7454 -11231 7488 -11197
rect 7712 -11231 7746 -11197
rect 7972 -11195 8006 -11161
rect 8239 -11221 8273 -11187
rect 8439 -11221 8473 -11187
rect 8660 -11221 8694 -11187
rect 8780 -11221 8814 -11187
rect 9000 -11231 9034 -11197
rect 9260 -11195 9294 -11161
rect 9518 -11195 9552 -11161
rect 9617 -11195 9651 -11161
rect 9716 -11195 9750 -11161
rect 9824 -11231 9858 -11197
rect 9927 -11231 9961 -11197
rect 10030 -11231 10064 -11197
rect 10380 -11231 10414 -11197
rect 10640 -11195 10674 -11161
rect 10815 -11221 10849 -11187
rect 11015 -11221 11049 -11187
rect 11236 -11221 11270 -11187
rect 11356 -11221 11390 -11187
rect 11668 -11231 11702 -11197
rect 11928 -11195 11962 -11161
rect 13662 -11231 13696 -11197
rect 13790 -11231 13824 -11197
rect 13918 -11231 13952 -11197
rect 14046 -11231 14080 -11197
rect 14154 -11195 14188 -11161
rect 14282 -11195 14316 -11161
rect 14410 -11195 14444 -11161
rect 14538 -11195 14572 -11161
rect 14858 -11231 14892 -11197
rect 14986 -11231 15020 -11197
rect 15114 -11231 15148 -11197
rect 15242 -11231 15276 -11197
rect 15350 -11195 15384 -11161
rect 15478 -11195 15512 -11161
rect 15606 -11195 15640 -11161
rect 15734 -11195 15768 -11161
rect 16050 -11231 16084 -11197
rect 16153 -11231 16187 -11197
rect 16256 -11231 16290 -11197
rect 16364 -11195 16398 -11161
rect 16463 -11195 16497 -11161
rect 16562 -11195 16596 -11161
rect -2902 -11675 -2868 -11641
rect -2799 -11675 -2765 -11641
rect -2696 -11675 -2662 -11641
rect -2588 -11711 -2554 -11677
rect -2489 -11711 -2455 -11677
rect -2390 -11711 -2356 -11677
rect -1522 -11711 -1488 -11677
rect -1423 -11711 -1389 -11677
rect -1324 -11711 -1290 -11677
rect -1216 -11675 -1182 -11641
rect -1113 -11675 -1079 -11641
rect -1010 -11675 -976 -11641
rect -786 -11711 -752 -11677
rect -687 -11711 -653 -11677
rect -588 -11711 -554 -11677
rect -480 -11675 -446 -11641
rect -377 -11675 -343 -11641
rect -274 -11675 -240 -11641
rect -16 -11675 18 -11641
rect 244 -11711 278 -11677
rect 464 -11685 498 -11651
rect 584 -11685 618 -11651
rect 805 -11685 839 -11651
rect 1005 -11685 1039 -11651
rect 1272 -11675 1306 -11641
rect 1532 -11711 1566 -11677
rect 1790 -11675 1824 -11641
rect 1893 -11675 1927 -11641
rect 1996 -11675 2030 -11641
rect 2104 -11711 2138 -11677
rect 2203 -11711 2237 -11677
rect 2302 -11711 2336 -11677
rect 2560 -11675 2594 -11641
rect 2820 -11711 2854 -11677
rect 3040 -11685 3074 -11651
rect 3160 -11685 3194 -11651
rect 3381 -11685 3415 -11651
rect 3581 -11685 3615 -11651
rect 3848 -11675 3882 -11641
rect 4108 -11711 4142 -11677
rect 4366 -11675 4400 -11641
rect 4469 -11675 4503 -11641
rect 4572 -11675 4606 -11641
rect 4680 -11711 4714 -11677
rect 4779 -11711 4813 -11677
rect 4878 -11711 4912 -11677
rect 5136 -11675 5170 -11641
rect 5396 -11711 5430 -11677
rect 5616 -11685 5650 -11651
rect 5736 -11685 5770 -11651
rect 5957 -11685 5991 -11651
rect 6157 -11685 6191 -11651
rect 6424 -11675 6458 -11641
rect 6684 -11711 6718 -11677
rect 6942 -11675 6976 -11641
rect 7045 -11675 7079 -11641
rect 7148 -11675 7182 -11641
rect 7256 -11711 7290 -11677
rect 7355 -11711 7389 -11677
rect 7454 -11711 7488 -11677
rect 7712 -11675 7746 -11641
rect 7972 -11711 8006 -11677
rect 8192 -11685 8226 -11651
rect 8312 -11685 8346 -11651
rect 8533 -11685 8567 -11651
rect 8733 -11685 8767 -11651
rect 9000 -11675 9034 -11641
rect 9260 -11711 9294 -11677
rect 9518 -11675 9552 -11641
rect 9621 -11675 9655 -11641
rect 9724 -11675 9758 -11641
rect 9832 -11711 9866 -11677
rect 9931 -11711 9965 -11677
rect 10030 -11711 10064 -11677
rect 10380 -11675 10414 -11641
rect 10640 -11711 10674 -11677
rect 10768 -11685 10802 -11651
rect 10888 -11685 10922 -11651
rect 11109 -11685 11143 -11651
rect 11309 -11685 11343 -11651
rect 11668 -11675 11702 -11641
rect 11928 -11711 11962 -11677
rect 12574 -11685 12608 -11651
rect 12642 -11685 12676 -11651
rect 12710 -11685 12744 -11651
rect 12778 -11685 12812 -11651
rect 12846 -11685 12880 -11651
rect 12914 -11685 12948 -11651
rect 13232 -11711 13266 -11677
rect 13492 -11675 13526 -11641
rect 13692 -11685 13726 -11651
rect 14119 -11685 14153 -11651
rect 14187 -11685 14221 -11651
rect 14255 -11685 14289 -11651
rect 14323 -11685 14357 -11651
rect 14391 -11685 14425 -11651
rect 14459 -11685 14493 -11651
rect 14527 -11685 14561 -11651
rect 14595 -11685 14629 -11651
rect 14663 -11685 14697 -11651
rect 14731 -11685 14765 -11651
rect 14799 -11685 14833 -11651
rect 14867 -11685 14901 -11651
rect 14935 -11685 14969 -11651
rect 15003 -11685 15037 -11651
rect 15071 -11685 15105 -11651
rect 15139 -11685 15173 -11651
rect 15682 -11711 15716 -11677
rect 15810 -11711 15844 -11677
rect 15938 -11711 15972 -11677
rect 16066 -11711 16100 -11677
rect 16174 -11675 16208 -11641
rect 16302 -11675 16336 -11641
rect 16430 -11675 16464 -11641
rect 16558 -11675 16592 -11641
rect -2902 -12283 -2868 -12249
rect -2803 -12283 -2769 -12249
rect -2704 -12283 -2670 -12249
rect -2596 -12319 -2562 -12285
rect -2493 -12319 -2459 -12285
rect -2390 -12319 -2356 -12285
rect -1522 -12319 -1488 -12285
rect -1419 -12319 -1385 -12285
rect -1316 -12319 -1282 -12285
rect -1208 -12283 -1174 -12249
rect -1109 -12283 -1075 -12249
rect -1010 -12283 -976 -12249
rect -777 -12309 -743 -12275
rect -577 -12309 -543 -12275
rect -356 -12309 -322 -12275
rect -236 -12309 -202 -12275
rect -16 -12319 18 -12285
rect 244 -12283 278 -12249
rect 511 -12309 545 -12275
rect 711 -12309 745 -12275
rect 932 -12309 966 -12275
rect 1052 -12309 1086 -12275
rect 1272 -12319 1306 -12285
rect 1532 -12283 1566 -12249
rect 1790 -12283 1824 -12249
rect 1889 -12283 1923 -12249
rect 1988 -12283 2022 -12249
rect 2096 -12319 2130 -12285
rect 2199 -12319 2233 -12285
rect 2302 -12319 2336 -12285
rect 2560 -12319 2594 -12285
rect 2820 -12283 2854 -12249
rect 3087 -12309 3121 -12275
rect 3287 -12309 3321 -12275
rect 3508 -12309 3542 -12275
rect 3628 -12309 3662 -12275
rect 3848 -12319 3882 -12285
rect 4108 -12283 4142 -12249
rect 4366 -12283 4400 -12249
rect 4465 -12283 4499 -12249
rect 4564 -12283 4598 -12249
rect 4672 -12319 4706 -12285
rect 4775 -12319 4809 -12285
rect 4878 -12319 4912 -12285
rect 5136 -12319 5170 -12285
rect 5396 -12283 5430 -12249
rect 5663 -12309 5697 -12275
rect 5863 -12309 5897 -12275
rect 6084 -12309 6118 -12275
rect 6204 -12309 6238 -12275
rect 6424 -12319 6458 -12285
rect 6684 -12283 6718 -12249
rect 6942 -12283 6976 -12249
rect 7041 -12283 7075 -12249
rect 7140 -12283 7174 -12249
rect 7248 -12319 7282 -12285
rect 7351 -12319 7385 -12285
rect 7454 -12319 7488 -12285
rect 7712 -12319 7746 -12285
rect 7972 -12283 8006 -12249
rect 8239 -12309 8273 -12275
rect 8439 -12309 8473 -12275
rect 8660 -12309 8694 -12275
rect 8780 -12309 8814 -12275
rect 9000 -12319 9034 -12285
rect 9260 -12283 9294 -12249
rect 9518 -12283 9552 -12249
rect 9617 -12283 9651 -12249
rect 9716 -12283 9750 -12249
rect 9824 -12319 9858 -12285
rect 9927 -12319 9961 -12285
rect 10030 -12319 10064 -12285
rect 10380 -12319 10414 -12285
rect 10640 -12283 10674 -12249
rect 10815 -12309 10849 -12275
rect 11015 -12309 11049 -12275
rect 11236 -12309 11270 -12275
rect 11356 -12309 11390 -12275
rect 11668 -12319 11702 -12285
rect 11928 -12283 11962 -12249
rect 13692 -12309 13726 -12275
rect 14119 -12309 14153 -12275
rect 14187 -12309 14221 -12275
rect 14255 -12309 14289 -12275
rect 14323 -12309 14357 -12275
rect 14391 -12309 14425 -12275
rect 14459 -12309 14493 -12275
rect 14527 -12309 14561 -12275
rect 14595 -12309 14629 -12275
rect 14663 -12309 14697 -12275
rect 14731 -12309 14765 -12275
rect 14799 -12309 14833 -12275
rect 14867 -12309 14901 -12275
rect 14935 -12309 14969 -12275
rect 15003 -12309 15037 -12275
rect 15071 -12309 15105 -12275
rect 15139 -12309 15173 -12275
rect 15686 -12319 15720 -12285
rect 15814 -12319 15848 -12285
rect 15942 -12319 15976 -12285
rect 16070 -12319 16104 -12285
rect 16178 -12283 16212 -12249
rect 16306 -12283 16340 -12249
rect 16434 -12283 16468 -12249
rect 16562 -12283 16596 -12249
rect -2902 -12763 -2868 -12729
rect -2799 -12763 -2765 -12729
rect -2696 -12763 -2662 -12729
rect -2588 -12799 -2554 -12765
rect -2489 -12799 -2455 -12765
rect -2390 -12799 -2356 -12765
rect -1522 -12799 -1488 -12765
rect -1423 -12799 -1389 -12765
rect -1324 -12799 -1290 -12765
rect -1216 -12763 -1182 -12729
rect -1113 -12763 -1079 -12729
rect -1010 -12763 -976 -12729
rect -786 -12799 -752 -12765
rect -687 -12799 -653 -12765
rect -588 -12799 -554 -12765
rect -480 -12763 -446 -12729
rect -377 -12763 -343 -12729
rect -274 -12763 -240 -12729
rect -16 -12763 18 -12729
rect 244 -12799 278 -12765
rect 464 -12773 498 -12739
rect 584 -12773 618 -12739
rect 805 -12773 839 -12739
rect 1005 -12773 1039 -12739
rect 1272 -12763 1306 -12729
rect 1532 -12799 1566 -12765
rect 1790 -12763 1824 -12729
rect 1893 -12763 1927 -12729
rect 1996 -12763 2030 -12729
rect 2104 -12799 2138 -12765
rect 2203 -12799 2237 -12765
rect 2302 -12799 2336 -12765
rect 2560 -12763 2594 -12729
rect 2820 -12799 2854 -12765
rect 3040 -12773 3074 -12739
rect 3160 -12773 3194 -12739
rect 3381 -12773 3415 -12739
rect 3581 -12773 3615 -12739
rect 3848 -12763 3882 -12729
rect 4108 -12799 4142 -12765
rect 4366 -12763 4400 -12729
rect 4469 -12763 4503 -12729
rect 4572 -12763 4606 -12729
rect 4680 -12799 4714 -12765
rect 4779 -12799 4813 -12765
rect 4878 -12799 4912 -12765
rect 5136 -12763 5170 -12729
rect 5396 -12799 5430 -12765
rect 5616 -12773 5650 -12739
rect 5736 -12773 5770 -12739
rect 5957 -12773 5991 -12739
rect 6157 -12773 6191 -12739
rect 6424 -12763 6458 -12729
rect 6684 -12799 6718 -12765
rect 6942 -12763 6976 -12729
rect 7045 -12763 7079 -12729
rect 7148 -12763 7182 -12729
rect 7256 -12799 7290 -12765
rect 7355 -12799 7389 -12765
rect 7454 -12799 7488 -12765
rect 7712 -12763 7746 -12729
rect 7972 -12799 8006 -12765
rect 8192 -12773 8226 -12739
rect 8312 -12773 8346 -12739
rect 8533 -12773 8567 -12739
rect 8733 -12773 8767 -12739
rect 9000 -12763 9034 -12729
rect 9260 -12799 9294 -12765
rect 9518 -12763 9552 -12729
rect 9621 -12763 9655 -12729
rect 9724 -12763 9758 -12729
rect 9832 -12799 9866 -12765
rect 9931 -12799 9965 -12765
rect 10030 -12799 10064 -12765
rect 10380 -12763 10414 -12729
rect 10640 -12799 10674 -12765
rect 10768 -12773 10802 -12739
rect 10888 -12773 10922 -12739
rect 11109 -12773 11143 -12739
rect 11309 -12773 11343 -12739
rect 11668 -12763 11702 -12729
rect 11928 -12799 11962 -12765
rect 12574 -12773 12608 -12739
rect 12642 -12773 12676 -12739
rect 12710 -12773 12744 -12739
rect 12778 -12773 12812 -12739
rect 12846 -12773 12880 -12739
rect 12914 -12773 12948 -12739
rect 13232 -12799 13266 -12765
rect 13492 -12763 13526 -12729
rect 13692 -12773 13726 -12739
rect 14119 -12773 14153 -12739
rect 14187 -12773 14221 -12739
rect 14255 -12773 14289 -12739
rect 14323 -12773 14357 -12739
rect 14391 -12773 14425 -12739
rect 14459 -12773 14493 -12739
rect 14527 -12773 14561 -12739
rect 14595 -12773 14629 -12739
rect 14663 -12773 14697 -12739
rect 14731 -12773 14765 -12739
rect 14799 -12773 14833 -12739
rect 14867 -12773 14901 -12739
rect 14935 -12773 14969 -12739
rect 15003 -12773 15037 -12739
rect 15071 -12773 15105 -12739
rect 15139 -12773 15173 -12739
rect 15682 -12799 15716 -12765
rect 15810 -12799 15844 -12765
rect 15938 -12799 15972 -12765
rect 16066 -12799 16100 -12765
rect 16174 -12763 16208 -12729
rect 16302 -12763 16336 -12729
rect 16430 -12763 16464 -12729
rect 16558 -12763 16592 -12729
rect -2902 -13371 -2868 -13337
rect -2803 -13371 -2769 -13337
rect -2704 -13371 -2670 -13337
rect -2596 -13407 -2562 -13373
rect -2493 -13407 -2459 -13373
rect -2390 -13407 -2356 -13373
rect -1522 -13407 -1488 -13373
rect -1419 -13407 -1385 -13373
rect -1316 -13407 -1282 -13373
rect -1208 -13371 -1174 -13337
rect -1109 -13371 -1075 -13337
rect -1010 -13371 -976 -13337
rect -786 -13407 -752 -13373
rect -683 -13407 -649 -13373
rect -580 -13407 -546 -13373
rect -472 -13371 -438 -13337
rect -373 -13371 -339 -13337
rect -274 -13371 -240 -13337
rect -16 -13407 18 -13373
rect 244 -13371 278 -13337
rect 511 -13397 545 -13363
rect 711 -13397 745 -13363
rect 932 -13397 966 -13363
rect 1052 -13397 1086 -13363
rect 1272 -13407 1306 -13373
rect 1532 -13371 1566 -13337
rect 1790 -13371 1824 -13337
rect 1889 -13371 1923 -13337
rect 1988 -13371 2022 -13337
rect 2096 -13407 2130 -13373
rect 2199 -13407 2233 -13373
rect 2302 -13407 2336 -13373
rect 2560 -13407 2594 -13373
rect 2820 -13371 2854 -13337
rect 3087 -13397 3121 -13363
rect 3287 -13397 3321 -13363
rect 3508 -13397 3542 -13363
rect 3628 -13397 3662 -13363
rect 3848 -13407 3882 -13373
rect 4108 -13371 4142 -13337
rect 4366 -13371 4400 -13337
rect 4465 -13371 4499 -13337
rect 4564 -13371 4598 -13337
rect 4672 -13407 4706 -13373
rect 4775 -13407 4809 -13373
rect 4878 -13407 4912 -13373
rect 5136 -13407 5170 -13373
rect 5396 -13371 5430 -13337
rect 5663 -13397 5697 -13363
rect 5863 -13397 5897 -13363
rect 6084 -13397 6118 -13363
rect 6204 -13397 6238 -13363
rect 6424 -13407 6458 -13373
rect 6684 -13371 6718 -13337
rect 6942 -13371 6976 -13337
rect 7041 -13371 7075 -13337
rect 7140 -13371 7174 -13337
rect 7248 -13407 7282 -13373
rect 7351 -13407 7385 -13373
rect 7454 -13407 7488 -13373
rect 7712 -13407 7746 -13373
rect 7972 -13371 8006 -13337
rect 8239 -13397 8273 -13363
rect 8439 -13397 8473 -13363
rect 8660 -13397 8694 -13363
rect 8780 -13397 8814 -13363
rect 9000 -13407 9034 -13373
rect 9260 -13371 9294 -13337
rect 9518 -13371 9552 -13337
rect 9617 -13371 9651 -13337
rect 9716 -13371 9750 -13337
rect 9824 -13407 9858 -13373
rect 9927 -13407 9961 -13373
rect 10030 -13407 10064 -13373
rect 10380 -13407 10414 -13373
rect 10640 -13371 10674 -13337
rect 10815 -13397 10849 -13363
rect 11015 -13397 11049 -13363
rect 11236 -13397 11270 -13363
rect 11356 -13397 11390 -13363
rect 11668 -13407 11702 -13373
rect 11928 -13371 11962 -13337
rect 13692 -13397 13726 -13363
rect 14119 -13397 14153 -13363
rect 14187 -13397 14221 -13363
rect 14255 -13397 14289 -13363
rect 14323 -13397 14357 -13363
rect 14391 -13397 14425 -13363
rect 14459 -13397 14493 -13363
rect 14527 -13397 14561 -13363
rect 14595 -13397 14629 -13363
rect 14663 -13397 14697 -13363
rect 14731 -13397 14765 -13363
rect 14799 -13397 14833 -13363
rect 14867 -13397 14901 -13363
rect 14935 -13397 14969 -13363
rect 15003 -13397 15037 -13363
rect 15071 -13397 15105 -13363
rect 15139 -13397 15173 -13363
rect 15686 -13407 15720 -13373
rect 15814 -13407 15848 -13373
rect 15942 -13407 15976 -13373
rect 16070 -13407 16104 -13373
rect 16178 -13371 16212 -13337
rect 16306 -13371 16340 -13337
rect 16434 -13371 16468 -13337
rect 16562 -13371 16596 -13337
rect -2902 -13851 -2868 -13817
rect -2799 -13851 -2765 -13817
rect -2696 -13851 -2662 -13817
rect -2588 -13887 -2554 -13853
rect -2489 -13887 -2455 -13853
rect -2390 -13887 -2356 -13853
rect -1396 -13887 -1362 -13853
rect -1136 -13851 -1102 -13817
rect -937 -13861 -903 -13827
rect -769 -13861 -735 -13827
rect -568 -13887 -534 -13853
rect -308 -13851 -274 -13817
rect -30 -13861 4 -13827
rect 38 -13861 72 -13827
rect 106 -13861 140 -13827
rect 174 -13861 208 -13827
rect 242 -13861 276 -13827
rect 310 -13861 344 -13827
rect 628 -13887 662 -13853
rect 888 -13851 922 -13817
rect 1082 -13861 1116 -13827
rect 1456 -13887 1490 -13853
rect 1716 -13851 1750 -13817
rect 1916 -13887 1950 -13853
rect 2176 -13851 2210 -13817
rect 2396 -13861 2430 -13827
rect 2516 -13861 2550 -13827
rect 2737 -13861 2771 -13827
rect 2937 -13861 2971 -13827
rect 3204 -13887 3238 -13853
rect 3464 -13851 3498 -13817
rect 4458 -13887 4492 -13853
rect 4586 -13887 4620 -13853
rect 4714 -13887 4748 -13853
rect 4842 -13887 4876 -13853
rect 4950 -13851 4984 -13817
rect 5078 -13851 5112 -13817
rect 5206 -13851 5240 -13817
rect 5334 -13851 5368 -13817
rect 6424 -13887 6458 -13853
rect 6684 -13851 6718 -13817
rect 6904 -13861 6938 -13827
rect 7024 -13861 7058 -13827
rect 7245 -13861 7279 -13827
rect 7445 -13861 7479 -13827
rect 7712 -13887 7746 -13853
rect 7972 -13851 8006 -13817
rect 8192 -13861 8226 -13827
rect 8312 -13861 8346 -13827
rect 8533 -13861 8567 -13827
rect 8733 -13861 8767 -13827
rect 9000 -13887 9034 -13853
rect 9260 -13851 9294 -13817
rect 9480 -13861 9514 -13827
rect 9600 -13861 9634 -13827
rect 9821 -13861 9855 -13827
rect 10021 -13861 10055 -13827
rect 10288 -13887 10322 -13853
rect 10548 -13851 10582 -13817
rect 10749 -13861 10783 -13827
rect 10830 -13861 10864 -13827
rect 10914 -13861 10948 -13827
rect 10998 -13861 11032 -13827
rect 11250 -13861 11284 -13827
rect 11334 -13861 11368 -13827
rect 11668 -13887 11702 -13853
rect 11928 -13851 11962 -13817
rect 13658 -13887 13692 -13853
rect 13786 -13887 13820 -13853
rect 13914 -13887 13948 -13853
rect 14042 -13887 14076 -13853
rect 14150 -13851 14184 -13817
rect 14278 -13851 14312 -13817
rect 14406 -13851 14440 -13817
rect 14534 -13851 14568 -13817
rect 14854 -13887 14888 -13853
rect 14982 -13887 15016 -13853
rect 15110 -13887 15144 -13853
rect 15238 -13887 15272 -13853
rect 15346 -13851 15380 -13817
rect 15474 -13851 15508 -13817
rect 15602 -13851 15636 -13817
rect 15730 -13851 15764 -13817
rect 16050 -13887 16084 -13853
rect 16149 -13887 16183 -13853
rect 16248 -13887 16282 -13853
rect 16356 -13851 16390 -13817
rect 16459 -13851 16493 -13817
rect 16562 -13851 16596 -13817
<< locali >>
rect -2997 -29 -2968 5
rect -2934 -29 -2876 5
rect -2842 -29 -2784 5
rect -2750 -29 -2692 5
rect -2658 -29 -2600 5
rect -2566 -29 -2508 5
rect -2474 -29 -2416 5
rect -2382 -29 -2324 5
rect -2290 -29 -2232 5
rect -2198 -29 -2140 5
rect -2106 -29 -2048 5
rect -2014 -29 -1956 5
rect -1922 -29 -1864 5
rect -1830 -29 -1772 5
rect -1738 -29 -1680 5
rect -1646 -29 -1588 5
rect -1554 -29 -1496 5
rect -1462 -29 -1404 5
rect -1370 -29 -1312 5
rect -1278 -29 -1220 5
rect -1186 -29 -1128 5
rect -1094 -29 -1036 5
rect -1002 -29 -944 5
rect -910 -29 -852 5
rect -818 -29 -760 5
rect -726 -29 -668 5
rect -634 -29 -576 5
rect -542 -29 -484 5
rect -450 -29 -392 5
rect -358 -29 -300 5
rect -266 -29 -208 5
rect -174 -29 -116 5
rect -82 -29 -24 5
rect 10 -29 68 5
rect 102 -29 160 5
rect 194 -29 252 5
rect 286 -29 344 5
rect 378 -29 436 5
rect 470 -29 528 5
rect 562 -29 620 5
rect 654 -29 712 5
rect 746 -29 804 5
rect 838 -29 896 5
rect 930 -29 988 5
rect 1022 -29 1080 5
rect 1114 -29 1172 5
rect 1206 -29 1264 5
rect 1298 -29 1356 5
rect 1390 -29 1448 5
rect 1482 -29 1540 5
rect 1574 -29 1632 5
rect 1666 -29 1724 5
rect 1758 -29 1816 5
rect 1850 -29 1908 5
rect 1942 -29 2000 5
rect 2034 -29 2092 5
rect 2126 -29 2184 5
rect 2218 -29 2276 5
rect 2310 -29 2368 5
rect 2402 -29 2460 5
rect 2494 -29 2552 5
rect 2586 -29 2644 5
rect 2678 -29 2736 5
rect 2770 -29 2828 5
rect 2862 -29 2920 5
rect 2954 -29 3012 5
rect 3046 -29 3104 5
rect 3138 -29 3196 5
rect 3230 -29 3288 5
rect 3322 -29 3380 5
rect 3414 -29 3472 5
rect 3506 -29 3564 5
rect 3598 -29 3656 5
rect 3690 -29 3748 5
rect 3782 -29 3840 5
rect 3874 -29 3932 5
rect 3966 -29 4024 5
rect 4058 -29 4116 5
rect 4150 -29 4208 5
rect 4242 -29 4300 5
rect 4334 -29 4392 5
rect 4426 -29 4484 5
rect 4518 -29 4576 5
rect 4610 -29 4668 5
rect 4702 -29 4760 5
rect 4794 -29 4852 5
rect 4886 -29 4944 5
rect 4978 -29 5036 5
rect 5070 -29 5128 5
rect 5162 -29 5220 5
rect 5254 -29 5312 5
rect 5346 -29 5404 5
rect 5438 -29 5496 5
rect 5530 -29 5588 5
rect 5622 -29 5680 5
rect 5714 -29 5772 5
rect 5806 -29 5864 5
rect 5898 -29 5956 5
rect 5990 -29 6048 5
rect 6082 -29 6140 5
rect 6174 -29 6232 5
rect 6266 -29 6324 5
rect 6358 -29 6416 5
rect 6450 -29 6508 5
rect 6542 -29 6600 5
rect 6634 -29 6692 5
rect 6726 -29 6784 5
rect 6818 -29 6876 5
rect 6910 -29 6968 5
rect 7002 -29 7060 5
rect 7094 -29 7152 5
rect 7186 -29 7244 5
rect 7278 -29 7336 5
rect 7370 -29 7428 5
rect 7462 -29 7520 5
rect 7554 -29 7612 5
rect 7646 -29 7704 5
rect 7738 -29 7796 5
rect 7830 -29 7888 5
rect 7922 -29 7980 5
rect 8014 -29 8072 5
rect 8106 -29 8164 5
rect 8198 -29 8256 5
rect 8290 -29 8348 5
rect 8382 -29 8440 5
rect 8474 -29 8532 5
rect 8566 -29 8624 5
rect 8658 -29 8716 5
rect 8750 -29 8808 5
rect 8842 -29 8900 5
rect 8934 -29 8992 5
rect 9026 -29 9084 5
rect 9118 -29 9176 5
rect 9210 -29 9268 5
rect 9302 -29 9360 5
rect 9394 -29 9452 5
rect 9486 -29 9544 5
rect 9578 -29 9636 5
rect 9670 -29 9728 5
rect 9762 -29 9820 5
rect 9854 -29 9912 5
rect 9946 -29 10004 5
rect 10038 -29 10096 5
rect 10130 -29 10188 5
rect 10222 -29 10280 5
rect 10314 -29 10372 5
rect 10406 -29 10464 5
rect 10498 -29 10556 5
rect 10590 -29 10648 5
rect 10682 -29 10740 5
rect 10774 -29 10832 5
rect 10866 -29 10924 5
rect 10958 -29 11016 5
rect 11050 -29 11108 5
rect 11142 -29 11200 5
rect 11234 -29 11292 5
rect 11326 -29 11384 5
rect 11418 -29 11476 5
rect 11510 -29 11568 5
rect 11602 -29 11660 5
rect 11694 -29 11752 5
rect 11786 -29 11844 5
rect 11878 -29 11936 5
rect 11970 -29 12028 5
rect 12062 -29 12120 5
rect 12154 -29 12212 5
rect 12246 -29 12304 5
rect 12338 -29 12396 5
rect 12430 -29 12488 5
rect 12522 -29 12580 5
rect 12614 -29 12672 5
rect 12706 -29 12764 5
rect 12798 -29 12856 5
rect 12890 -29 12948 5
rect 12982 -29 13040 5
rect 13074 -29 13132 5
rect 13166 -29 13224 5
rect 13258 -29 13316 5
rect 13350 -29 13408 5
rect 13442 -29 13500 5
rect 13534 -29 13592 5
rect 13626 -29 13684 5
rect 13718 -29 13776 5
rect 13810 -29 13868 5
rect 13902 -29 13960 5
rect 13994 -29 14052 5
rect 14086 -29 14144 5
rect 14178 -29 14236 5
rect 14270 -29 14328 5
rect 14362 -29 14420 5
rect 14454 -29 14512 5
rect 14546 -29 14604 5
rect 14638 -29 14696 5
rect 14730 -29 14788 5
rect 14822 -29 14880 5
rect 14914 -29 14972 5
rect 15006 -29 15064 5
rect 15098 -29 15156 5
rect 15190 -29 15248 5
rect 15282 -29 15340 5
rect 15374 -29 15432 5
rect 15466 -29 15524 5
rect 15558 -29 15616 5
rect 15650 -29 15708 5
rect 15742 -29 15800 5
rect 15834 -29 15892 5
rect 15926 -29 15984 5
rect 16018 -29 16076 5
rect 16110 -29 16168 5
rect 16202 -29 16260 5
rect 16294 -29 16352 5
rect 16386 -29 16444 5
rect 16478 -29 16536 5
rect 16570 -29 16628 5
rect 16662 -29 16691 5
rect -2980 -71 -2278 -29
rect -2980 -105 -2962 -71
rect -2928 -105 -2330 -71
rect -2296 -105 -2278 -71
rect -2980 -173 -2278 -105
rect -2980 -207 -2962 -173
rect -2928 -207 -2330 -173
rect -2296 -207 -2278 -173
rect -2980 -247 -2278 -207
rect -2980 -315 -2902 -281
rect -2868 -315 -2803 -281
rect -2769 -315 -2704 -281
rect -2670 -315 -2650 -281
rect -2980 -385 -2650 -315
rect -2616 -317 -2278 -247
rect -2244 -100 -2186 -29
rect -2244 -134 -2232 -100
rect -2198 -134 -2186 -100
rect -2244 -193 -2186 -134
rect -2244 -227 -2232 -193
rect -2198 -227 -2186 -193
rect -2244 -262 -2186 -227
rect -1416 -71 -1082 -29
rect -1416 -105 -1398 -71
rect -1364 -105 -1134 -71
rect -1100 -105 -1082 -71
rect -1416 -173 -1082 -105
rect -1416 -207 -1398 -173
rect -1364 -207 -1134 -173
rect -1100 -207 -1082 -173
rect -1416 -247 -1082 -207
rect -2616 -351 -2596 -317
rect -2562 -351 -2493 -317
rect -2459 -351 -2390 -317
rect -2356 -351 -2278 -317
rect -1416 -315 -1396 -281
rect -1362 -315 -1266 -281
rect -1416 -385 -1266 -315
rect -1232 -317 -1082 -247
rect -1048 -100 -990 -29
rect -1048 -134 -1036 -100
rect -1002 -134 -990 -100
rect -1048 -193 -990 -134
rect -1048 -227 -1036 -193
rect -1002 -227 -990 -193
rect -1048 -262 -990 -227
rect -956 -71 -900 -29
rect -956 -105 -934 -71
rect -956 -139 -900 -105
rect -956 -173 -934 -139
rect -956 -207 -900 -173
rect -956 -241 -934 -207
rect -956 -257 -900 -241
rect -866 -71 -800 -63
rect -866 -105 -850 -71
rect -816 -105 -800 -71
rect -866 -139 -800 -105
rect -866 -173 -850 -139
rect -816 -173 -800 -139
rect -866 -207 -800 -173
rect -866 -241 -850 -207
rect -816 -241 -800 -207
rect -866 -259 -800 -241
rect -766 -71 -714 -29
rect -732 -105 -714 -71
rect -766 -139 -714 -105
rect -732 -173 -714 -139
rect -766 -207 -714 -173
rect -732 -241 -714 -207
rect -766 -257 -714 -241
rect -680 -100 -622 -29
rect -680 -134 -668 -100
rect -634 -134 -622 -100
rect -680 -193 -622 -134
rect -680 -227 -668 -193
rect -634 -227 -622 -193
rect -1232 -351 -1136 -317
rect -1102 -351 -1082 -317
rect -954 -301 -887 -291
rect -954 -335 -943 -301
rect -909 -307 -887 -301
rect -954 -341 -937 -335
rect -903 -341 -887 -307
rect -954 -345 -887 -341
rect -853 -379 -819 -259
rect -680 -262 -622 -227
rect -588 -71 -254 -29
rect -588 -105 -570 -71
rect -536 -105 -306 -71
rect -272 -105 -254 -71
rect -588 -173 -254 -105
rect -588 -207 -570 -173
rect -536 -207 -306 -173
rect -272 -207 -254 -173
rect -588 -247 -254 -207
rect -785 -301 -718 -291
rect -785 -307 -762 -301
rect -785 -341 -769 -307
rect -728 -335 -718 -301
rect -735 -341 -718 -335
rect -588 -315 -568 -281
rect -534 -315 -438 -281
rect -2980 -444 -2278 -385
rect -2980 -478 -2962 -444
rect -2928 -478 -2330 -444
rect -2296 -478 -2278 -444
rect -2980 -539 -2278 -478
rect -2244 -411 -2186 -394
rect -2244 -445 -2232 -411
rect -2198 -445 -2186 -411
rect -2244 -539 -2186 -445
rect -1416 -437 -1082 -385
rect -1416 -471 -1398 -437
rect -1364 -471 -1134 -437
rect -1100 -471 -1082 -437
rect -1416 -539 -1082 -471
rect -1048 -411 -990 -394
rect -1048 -445 -1036 -411
rect -1002 -445 -990 -411
rect -1048 -539 -990 -445
rect -956 -395 -894 -379
rect -956 -429 -934 -395
rect -900 -429 -894 -395
rect -956 -463 -894 -429
rect -956 -497 -934 -463
rect -900 -497 -894 -463
rect -956 -539 -894 -497
rect -853 -395 -714 -379
rect -588 -385 -438 -315
rect -404 -317 -254 -247
rect -220 -100 -162 -29
rect -220 -134 -208 -100
rect -174 -134 -162 -100
rect -220 -193 -162 -134
rect -220 -227 -208 -193
rect -174 -227 -162 -193
rect -128 -78 -59 -29
rect -128 -112 -102 -78
rect -68 -112 -59 -78
rect -128 -146 -59 -112
rect -128 -180 -102 -146
rect -68 -180 -59 -146
rect -128 -196 -59 -180
rect -24 -85 27 -69
rect -24 -119 -16 -85
rect 18 -119 27 -85
rect -24 -173 27 -119
rect -220 -262 -162 -227
rect -24 -207 -16 -173
rect 18 -207 27 -173
rect 61 -78 113 -29
rect 61 -112 70 -78
rect 104 -112 113 -78
rect 61 -146 113 -112
rect 61 -180 70 -146
rect 104 -180 113 -146
rect 61 -196 113 -180
rect 148 -85 199 -69
rect 148 -119 156 -85
rect 190 -119 199 -85
rect 148 -173 199 -119
rect -24 -230 27 -207
rect 148 -207 156 -173
rect 190 -207 199 -173
rect 233 -78 285 -29
rect 233 -112 242 -78
rect 276 -112 285 -78
rect 233 -146 285 -112
rect 233 -180 242 -146
rect 276 -180 285 -146
rect 233 -196 285 -180
rect 319 -85 371 -69
rect 319 -119 328 -85
rect 362 -119 371 -85
rect 319 -173 371 -119
rect 148 -230 199 -207
rect 319 -207 328 -173
rect 362 -207 371 -173
rect 405 -78 482 -29
rect 405 -112 414 -78
rect 448 -112 482 -78
rect 405 -146 482 -112
rect 405 -180 414 -146
rect 448 -180 482 -146
rect 405 -196 482 -180
rect 516 -100 574 -29
rect 516 -134 528 -100
rect 562 -134 574 -100
rect 516 -193 574 -134
rect 319 -230 371 -207
rect 516 -227 528 -193
rect 562 -227 574 -193
rect -404 -351 -308 -317
rect -274 -351 -254 -317
rect -124 -264 482 -230
rect 516 -262 574 -227
rect 608 -71 942 -29
rect 608 -105 626 -71
rect 660 -105 890 -71
rect 924 -105 942 -71
rect 608 -173 942 -105
rect 608 -207 626 -173
rect 660 -207 890 -173
rect 924 -207 942 -173
rect 608 -247 942 -207
rect -124 -377 -90 -264
rect -56 -307 387 -298
rect -56 -341 -30 -307
rect 4 -341 38 -307
rect 72 -341 106 -307
rect 140 -341 174 -307
rect 208 -341 242 -307
rect 276 -341 310 -307
rect 344 -341 387 -307
rect -56 -343 387 -341
rect 422 -345 482 -264
rect 422 -377 434 -345
rect -124 -379 434 -377
rect 468 -379 482 -345
rect -853 -412 -766 -395
rect -853 -446 -848 -412
rect -814 -446 -769 -412
rect -732 -429 -714 -395
rect -735 -446 -714 -429
rect -853 -463 -714 -446
rect -853 -497 -766 -463
rect -732 -497 -714 -463
rect -853 -505 -714 -497
rect -680 -411 -622 -394
rect -680 -445 -668 -411
rect -634 -445 -622 -411
rect -680 -539 -622 -445
rect -588 -437 -254 -385
rect -588 -471 -570 -437
rect -536 -471 -306 -437
rect -272 -471 -254 -437
rect -588 -539 -254 -471
rect -220 -411 -162 -394
rect -124 -411 482 -379
rect 608 -315 628 -281
rect 662 -315 758 -281
rect 608 -385 758 -315
rect 792 -317 942 -247
rect 976 -100 1034 -29
rect 976 -134 988 -100
rect 1022 -134 1034 -100
rect 976 -193 1034 -134
rect 976 -227 988 -193
rect 1022 -227 1034 -193
rect 1068 -71 1120 -29
rect 1068 -105 1086 -71
rect 1068 -173 1120 -105
rect 1068 -207 1086 -173
rect 1068 -223 1120 -207
rect 1154 -71 1220 -63
rect 1154 -105 1170 -71
rect 1204 -105 1220 -71
rect 1154 -173 1220 -105
rect 1154 -207 1170 -173
rect 1204 -207 1220 -173
rect 976 -262 1034 -227
rect 792 -351 888 -317
rect 922 -351 942 -317
rect 1068 -307 1116 -291
rect 1068 -312 1082 -307
rect 1068 -346 1076 -312
rect 1110 -346 1116 -341
rect 1068 -385 1116 -346
rect 516 -411 574 -394
rect -220 -445 -208 -411
rect -174 -445 -162 -411
rect -220 -539 -162 -445
rect -32 -461 27 -445
rect -32 -495 -16 -461
rect 18 -495 27 -461
rect -32 -539 27 -495
rect 61 -450 113 -411
rect 61 -484 70 -450
rect 104 -484 113 -450
rect 61 -500 113 -484
rect 147 -461 199 -445
rect 147 -495 156 -461
rect 190 -495 199 -461
rect 147 -539 199 -495
rect 233 -450 284 -411
rect 516 -445 528 -411
rect 562 -445 574 -411
rect 233 -484 242 -450
rect 276 -484 284 -450
rect 233 -500 284 -484
rect 318 -461 378 -445
rect 318 -495 328 -461
rect 362 -495 378 -461
rect 318 -539 378 -495
rect 516 -539 574 -445
rect 608 -437 942 -385
rect 608 -471 626 -437
rect 660 -471 890 -437
rect 924 -471 942 -437
rect 608 -539 942 -471
rect 976 -411 1034 -394
rect 976 -445 988 -411
rect 1022 -445 1034 -411
rect 976 -539 1034 -445
rect 1068 -419 1076 -385
rect 1110 -419 1116 -385
rect 1068 -481 1116 -419
rect 1154 -298 1220 -207
rect 1254 -71 1310 -29
rect 1288 -105 1310 -71
rect 1254 -173 1310 -105
rect 1288 -207 1310 -173
rect 1254 -223 1310 -207
rect 1344 -100 1402 -29
rect 1344 -134 1356 -100
rect 1390 -134 1402 -100
rect 1344 -193 1402 -134
rect 1344 -227 1356 -193
rect 1390 -227 1402 -193
rect 1344 -262 1402 -227
rect 1436 -71 1770 -29
rect 1436 -105 1454 -71
rect 1488 -105 1718 -71
rect 1752 -105 1770 -71
rect 1436 -173 1770 -105
rect 1436 -207 1454 -173
rect 1488 -207 1718 -173
rect 1752 -207 1770 -173
rect 1436 -247 1770 -207
rect 1154 -306 1310 -298
rect 1154 -340 1171 -306
rect 1205 -340 1263 -306
rect 1297 -340 1310 -306
rect 1154 -404 1310 -340
rect 1436 -315 1456 -281
rect 1490 -315 1586 -281
rect 1436 -385 1586 -315
rect 1620 -317 1770 -247
rect 1804 -100 1862 -29
rect 1804 -134 1816 -100
rect 1850 -134 1862 -100
rect 1804 -193 1862 -134
rect 1804 -227 1816 -193
rect 1850 -227 1862 -193
rect 1804 -262 1862 -227
rect 1896 -71 2230 -29
rect 1896 -105 1914 -71
rect 1948 -105 2178 -71
rect 2212 -105 2230 -71
rect 1896 -173 2230 -105
rect 1896 -207 1914 -173
rect 1948 -207 2178 -173
rect 2212 -207 2230 -173
rect 1896 -247 2230 -207
rect 1620 -351 1716 -317
rect 1750 -351 1770 -317
rect 1896 -315 1916 -281
rect 1950 -315 2046 -281
rect 1896 -385 2046 -315
rect 2080 -317 2230 -247
rect 2264 -100 2322 -29
rect 2264 -134 2276 -100
rect 2310 -134 2322 -100
rect 2264 -193 2322 -134
rect 2264 -227 2276 -193
rect 2310 -227 2322 -193
rect 2264 -262 2322 -227
rect 2356 -78 2425 -63
rect 2356 -112 2375 -78
rect 2409 -112 2425 -78
rect 2356 -146 2425 -112
rect 2356 -180 2375 -146
rect 2409 -180 2425 -146
rect 2356 -230 2425 -180
rect 2459 -78 2525 -29
rect 2459 -112 2475 -78
rect 2509 -112 2525 -78
rect 2459 -146 2525 -112
rect 2459 -180 2475 -146
rect 2509 -180 2525 -146
rect 2459 -196 2525 -180
rect 2615 -78 2685 -63
rect 2615 -112 2633 -78
rect 2667 -112 2685 -78
rect 2615 -146 2685 -112
rect 2615 -180 2633 -146
rect 2667 -180 2685 -146
rect 2356 -264 2550 -230
rect 2480 -293 2550 -264
rect 2615 -292 2685 -180
rect 2737 -79 2787 -63
rect 2771 -113 2787 -79
rect 2737 -147 2787 -113
rect 2771 -181 2787 -147
rect 2737 -223 2787 -181
rect 2877 -78 2943 -29
rect 2877 -112 2893 -78
rect 2927 -112 2943 -78
rect 2877 -146 2943 -112
rect 2877 -180 2893 -146
rect 2927 -180 2943 -146
rect 2877 -189 2943 -180
rect 2977 -79 3058 -63
rect 2977 -113 2991 -79
rect 3025 -113 3058 -79
rect 2977 -147 3058 -113
rect 2977 -181 2991 -147
rect 3025 -181 3058 -147
rect 2977 -218 3058 -181
rect 2737 -257 2855 -223
rect 2821 -291 2855 -257
rect 2080 -351 2176 -317
rect 2210 -351 2230 -317
rect 2356 -301 2446 -298
rect 2356 -335 2369 -301
rect 2403 -307 2446 -301
rect 2356 -341 2396 -335
rect 2430 -341 2446 -307
rect 2480 -307 2566 -293
rect 2480 -341 2516 -307
rect 2550 -341 2566 -307
rect 2480 -351 2566 -341
rect 2615 -307 2787 -292
rect 2615 -341 2737 -307
rect 2771 -341 2787 -307
rect 2615 -342 2787 -341
rect 2821 -307 2974 -291
rect 2821 -341 2937 -307
rect 2971 -341 2974 -307
rect 2480 -375 2550 -351
rect 1154 -452 1219 -404
rect 1344 -411 1402 -394
rect 1154 -486 1169 -452
rect 1203 -486 1219 -452
rect 1154 -505 1219 -486
rect 1253 -454 1310 -438
rect 1287 -488 1310 -454
rect 1253 -539 1310 -488
rect 1344 -445 1356 -411
rect 1390 -445 1402 -411
rect 1344 -539 1402 -445
rect 1436 -437 1770 -385
rect 1436 -471 1454 -437
rect 1488 -471 1718 -437
rect 1752 -471 1770 -437
rect 1436 -539 1770 -471
rect 1804 -411 1862 -394
rect 1804 -445 1816 -411
rect 1850 -445 1862 -411
rect 1804 -539 1862 -445
rect 1896 -437 2230 -385
rect 1896 -471 1914 -437
rect 1948 -471 2178 -437
rect 2212 -471 2230 -437
rect 1896 -539 2230 -471
rect 2264 -411 2322 -394
rect 2264 -445 2276 -411
rect 2310 -445 2322 -411
rect 2264 -539 2322 -445
rect 2356 -409 2550 -375
rect 2356 -452 2422 -409
rect 2356 -486 2375 -452
rect 2409 -486 2422 -452
rect 2356 -505 2422 -486
rect 2456 -452 2522 -443
rect 2456 -486 2472 -452
rect 2506 -486 2522 -452
rect 2456 -539 2522 -486
rect 2615 -452 2685 -342
rect 2821 -357 2974 -341
rect 3008 -302 3058 -218
rect 3092 -100 3150 -29
rect 3092 -134 3104 -100
rect 3138 -134 3150 -100
rect 3092 -193 3150 -134
rect 3092 -227 3104 -193
rect 3138 -227 3150 -193
rect 3092 -262 3150 -227
rect 3184 -71 3518 -29
rect 3184 -105 3202 -71
rect 3236 -105 3466 -71
rect 3500 -105 3518 -71
rect 3184 -173 3518 -105
rect 3184 -207 3202 -173
rect 3236 -207 3466 -173
rect 3500 -207 3518 -173
rect 3184 -247 3518 -207
rect 3008 -336 3015 -302
rect 3049 -336 3058 -302
rect 2821 -376 2855 -357
rect 2615 -486 2632 -452
rect 2666 -486 2685 -452
rect 2615 -505 2685 -486
rect 2737 -410 2855 -376
rect 2737 -452 2787 -410
rect 3008 -428 3058 -336
rect 3184 -315 3204 -281
rect 3238 -315 3334 -281
rect 3184 -385 3334 -315
rect 3368 -317 3518 -247
rect 3552 -100 3610 -29
rect 3552 -134 3564 -100
rect 3598 -134 3610 -100
rect 3552 -193 3610 -134
rect 3552 -227 3564 -193
rect 3598 -227 3610 -193
rect 3552 -262 3610 -227
rect 4380 -71 5449 -29
rect 4380 -105 4398 -71
rect 4432 -105 5398 -71
rect 5432 -105 5449 -71
rect 4380 -173 5449 -105
rect 4380 -207 4398 -173
rect 4432 -207 5398 -173
rect 5432 -207 5449 -173
rect 4380 -247 5449 -207
rect 3368 -351 3464 -317
rect 3498 -351 3518 -317
rect 4380 -315 4458 -281
rect 4492 -315 4586 -281
rect 4620 -315 4714 -281
rect 4748 -315 4842 -281
rect 4876 -315 4896 -281
rect 4380 -385 4896 -315
rect 4930 -317 5449 -247
rect 6312 -100 6370 -29
rect 6312 -134 6324 -100
rect 6358 -134 6370 -100
rect 6312 -193 6370 -134
rect 6312 -227 6324 -193
rect 6358 -227 6370 -193
rect 6312 -262 6370 -227
rect 6404 -71 6738 -29
rect 6404 -105 6422 -71
rect 6456 -105 6686 -71
rect 6720 -105 6738 -71
rect 6404 -173 6738 -105
rect 6404 -207 6422 -173
rect 6456 -207 6686 -173
rect 6720 -207 6738 -173
rect 6404 -247 6738 -207
rect 4930 -351 4950 -317
rect 4984 -351 5078 -317
rect 5112 -351 5206 -317
rect 5240 -351 5334 -317
rect 5368 -351 5449 -317
rect 6404 -315 6424 -281
rect 6458 -315 6554 -281
rect 6404 -385 6554 -315
rect 6588 -317 6738 -247
rect 6772 -100 6830 -29
rect 6772 -134 6784 -100
rect 6818 -134 6830 -100
rect 6772 -193 6830 -134
rect 6772 -227 6784 -193
rect 6818 -227 6830 -193
rect 6772 -262 6830 -227
rect 6864 -78 6933 -63
rect 6864 -112 6883 -78
rect 6917 -112 6933 -78
rect 6864 -146 6933 -112
rect 6864 -180 6883 -146
rect 6917 -180 6933 -146
rect 6864 -230 6933 -180
rect 6967 -78 7033 -29
rect 6967 -112 6983 -78
rect 7017 -112 7033 -78
rect 6967 -146 7033 -112
rect 6967 -180 6983 -146
rect 7017 -180 7033 -146
rect 6967 -196 7033 -180
rect 7123 -78 7193 -63
rect 7123 -112 7141 -78
rect 7175 -112 7193 -78
rect 7123 -146 7193 -112
rect 7123 -180 7141 -146
rect 7175 -180 7193 -146
rect 6864 -264 7058 -230
rect 6988 -293 7058 -264
rect 7123 -292 7193 -180
rect 7245 -79 7295 -63
rect 7279 -113 7295 -79
rect 7245 -147 7295 -113
rect 7279 -181 7295 -147
rect 7245 -223 7295 -181
rect 7385 -78 7451 -29
rect 7385 -112 7401 -78
rect 7435 -112 7451 -78
rect 7385 -146 7451 -112
rect 7385 -180 7401 -146
rect 7435 -180 7451 -146
rect 7385 -189 7451 -180
rect 7485 -79 7566 -63
rect 7485 -113 7499 -79
rect 7533 -113 7566 -79
rect 7485 -147 7566 -113
rect 7485 -181 7499 -147
rect 7533 -181 7566 -147
rect 7485 -218 7566 -181
rect 7245 -257 7363 -223
rect 7329 -291 7363 -257
rect 6588 -351 6684 -317
rect 6718 -351 6738 -317
rect 6864 -302 6954 -298
rect 6864 -336 6876 -302
rect 6910 -307 6954 -302
rect 6864 -341 6904 -336
rect 6938 -341 6954 -307
rect 6988 -307 7074 -293
rect 6988 -341 7024 -307
rect 7058 -341 7074 -307
rect 6988 -351 7074 -341
rect 7123 -307 7295 -292
rect 7123 -341 7245 -307
rect 7279 -341 7295 -307
rect 7123 -342 7295 -341
rect 7329 -307 7482 -291
rect 7329 -341 7445 -307
rect 7479 -341 7482 -307
rect 6988 -375 7058 -351
rect 2771 -486 2787 -452
rect 2737 -505 2787 -486
rect 2877 -452 2943 -436
rect 2877 -486 2893 -452
rect 2927 -486 2943 -452
rect 2877 -539 2943 -486
rect 2977 -452 3058 -428
rect 2977 -486 2991 -452
rect 3025 -486 3058 -452
rect 2977 -505 3058 -486
rect 3092 -411 3150 -394
rect 3092 -445 3104 -411
rect 3138 -445 3150 -411
rect 3092 -539 3150 -445
rect 3184 -437 3518 -385
rect 3184 -471 3202 -437
rect 3236 -471 3466 -437
rect 3500 -471 3518 -437
rect 3184 -539 3518 -471
rect 3552 -411 3610 -394
rect 3552 -445 3564 -411
rect 3598 -445 3610 -411
rect 3552 -539 3610 -445
rect 4380 -444 5449 -385
rect 4380 -478 4398 -444
rect 4432 -478 5398 -444
rect 5432 -478 5449 -444
rect 4380 -539 5449 -478
rect 6312 -411 6370 -394
rect 6312 -445 6324 -411
rect 6358 -445 6370 -411
rect 6312 -539 6370 -445
rect 6404 -437 6738 -385
rect 6404 -471 6422 -437
rect 6456 -471 6686 -437
rect 6720 -471 6738 -437
rect 6404 -539 6738 -471
rect 6772 -411 6830 -394
rect 6772 -445 6784 -411
rect 6818 -445 6830 -411
rect 6772 -539 6830 -445
rect 6864 -409 7058 -375
rect 6864 -452 6930 -409
rect 6864 -486 6883 -452
rect 6917 -486 6930 -452
rect 6864 -505 6930 -486
rect 6964 -452 7030 -443
rect 6964 -486 6980 -452
rect 7014 -486 7030 -452
rect 6964 -539 7030 -486
rect 7123 -452 7193 -342
rect 7329 -357 7482 -341
rect 7516 -302 7566 -218
rect 7600 -100 7658 -29
rect 7600 -134 7612 -100
rect 7646 -134 7658 -100
rect 7600 -193 7658 -134
rect 7600 -227 7612 -193
rect 7646 -227 7658 -193
rect 7600 -262 7658 -227
rect 7692 -71 8026 -29
rect 7692 -105 7710 -71
rect 7744 -105 7974 -71
rect 8008 -105 8026 -71
rect 7692 -173 8026 -105
rect 7692 -207 7710 -173
rect 7744 -207 7974 -173
rect 8008 -207 8026 -173
rect 7692 -247 8026 -207
rect 7516 -336 7522 -302
rect 7556 -336 7566 -302
rect 7329 -376 7363 -357
rect 7123 -486 7140 -452
rect 7174 -486 7193 -452
rect 7123 -505 7193 -486
rect 7245 -410 7363 -376
rect 7245 -452 7295 -410
rect 7516 -428 7566 -336
rect 7692 -315 7712 -281
rect 7746 -315 7842 -281
rect 7692 -385 7842 -315
rect 7876 -317 8026 -247
rect 8060 -100 8118 -29
rect 8060 -134 8072 -100
rect 8106 -134 8118 -100
rect 8060 -193 8118 -134
rect 8060 -227 8072 -193
rect 8106 -227 8118 -193
rect 8060 -262 8118 -227
rect 8152 -78 8221 -63
rect 8152 -112 8171 -78
rect 8205 -112 8221 -78
rect 8152 -146 8221 -112
rect 8152 -180 8171 -146
rect 8205 -180 8221 -146
rect 8152 -230 8221 -180
rect 8255 -78 8321 -29
rect 8255 -112 8271 -78
rect 8305 -112 8321 -78
rect 8255 -146 8321 -112
rect 8255 -180 8271 -146
rect 8305 -180 8321 -146
rect 8255 -196 8321 -180
rect 8411 -78 8481 -63
rect 8411 -112 8429 -78
rect 8463 -112 8481 -78
rect 8411 -146 8481 -112
rect 8411 -180 8429 -146
rect 8463 -180 8481 -146
rect 8152 -264 8346 -230
rect 8276 -293 8346 -264
rect 8411 -292 8481 -180
rect 8533 -79 8583 -63
rect 8567 -113 8583 -79
rect 8533 -147 8583 -113
rect 8567 -181 8583 -147
rect 8533 -223 8583 -181
rect 8673 -78 8739 -29
rect 8673 -112 8689 -78
rect 8723 -112 8739 -78
rect 8673 -146 8739 -112
rect 8673 -180 8689 -146
rect 8723 -180 8739 -146
rect 8673 -189 8739 -180
rect 8773 -79 8854 -63
rect 8773 -113 8787 -79
rect 8821 -113 8854 -79
rect 8773 -147 8854 -113
rect 8773 -181 8787 -147
rect 8821 -181 8854 -147
rect 8773 -218 8854 -181
rect 8533 -257 8651 -223
rect 8617 -291 8651 -257
rect 7876 -351 7972 -317
rect 8006 -351 8026 -317
rect 8152 -303 8242 -298
rect 8152 -337 8164 -303
rect 8198 -307 8242 -303
rect 8152 -341 8192 -337
rect 8226 -341 8242 -307
rect 8276 -307 8362 -293
rect 8276 -341 8312 -307
rect 8346 -341 8362 -307
rect 8276 -351 8362 -341
rect 8411 -307 8583 -292
rect 8411 -341 8533 -307
rect 8567 -341 8583 -307
rect 8411 -342 8583 -341
rect 8617 -307 8770 -291
rect 8617 -341 8733 -307
rect 8767 -341 8770 -307
rect 8276 -375 8346 -351
rect 7279 -486 7295 -452
rect 7245 -505 7295 -486
rect 7385 -452 7451 -436
rect 7385 -486 7401 -452
rect 7435 -486 7451 -452
rect 7385 -539 7451 -486
rect 7485 -452 7566 -428
rect 7485 -486 7499 -452
rect 7533 -486 7566 -452
rect 7485 -505 7566 -486
rect 7600 -411 7658 -394
rect 7600 -445 7612 -411
rect 7646 -445 7658 -411
rect 7600 -539 7658 -445
rect 7692 -437 8026 -385
rect 7692 -471 7710 -437
rect 7744 -471 7974 -437
rect 8008 -471 8026 -437
rect 7692 -539 8026 -471
rect 8060 -411 8118 -394
rect 8060 -445 8072 -411
rect 8106 -445 8118 -411
rect 8060 -539 8118 -445
rect 8152 -409 8346 -375
rect 8152 -452 8218 -409
rect 8152 -486 8171 -452
rect 8205 -486 8218 -452
rect 8152 -505 8218 -486
rect 8252 -452 8318 -443
rect 8252 -486 8268 -452
rect 8302 -486 8318 -452
rect 8252 -539 8318 -486
rect 8411 -452 8481 -342
rect 8617 -357 8770 -341
rect 8804 -301 8854 -218
rect 8888 -100 8946 -29
rect 8888 -134 8900 -100
rect 8934 -134 8946 -100
rect 8888 -193 8946 -134
rect 8888 -227 8900 -193
rect 8934 -227 8946 -193
rect 8888 -262 8946 -227
rect 8980 -71 9314 -29
rect 8980 -105 8998 -71
rect 9032 -105 9262 -71
rect 9296 -105 9314 -71
rect 8980 -173 9314 -105
rect 8980 -207 8998 -173
rect 9032 -207 9262 -173
rect 9296 -207 9314 -173
rect 8980 -247 9314 -207
rect 8804 -335 8811 -301
rect 8845 -335 8854 -301
rect 8617 -376 8651 -357
rect 8411 -486 8428 -452
rect 8462 -486 8481 -452
rect 8411 -505 8481 -486
rect 8533 -410 8651 -376
rect 8533 -452 8583 -410
rect 8804 -428 8854 -335
rect 8980 -315 9000 -281
rect 9034 -315 9130 -281
rect 8980 -385 9130 -315
rect 9164 -317 9314 -247
rect 9348 -100 9406 -29
rect 9348 -134 9360 -100
rect 9394 -134 9406 -100
rect 9348 -193 9406 -134
rect 9348 -227 9360 -193
rect 9394 -227 9406 -193
rect 9348 -262 9406 -227
rect 9440 -78 9509 -63
rect 9440 -112 9459 -78
rect 9493 -112 9509 -78
rect 9440 -146 9509 -112
rect 9440 -180 9459 -146
rect 9493 -180 9509 -146
rect 9440 -230 9509 -180
rect 9543 -78 9609 -29
rect 9543 -112 9559 -78
rect 9593 -112 9609 -78
rect 9543 -146 9609 -112
rect 9543 -180 9559 -146
rect 9593 -180 9609 -146
rect 9543 -196 9609 -180
rect 9699 -78 9769 -63
rect 9699 -112 9717 -78
rect 9751 -112 9769 -78
rect 9699 -146 9769 -112
rect 9699 -180 9717 -146
rect 9751 -180 9769 -146
rect 9440 -264 9634 -230
rect 9564 -293 9634 -264
rect 9699 -292 9769 -180
rect 9821 -79 9871 -63
rect 9855 -113 9871 -79
rect 9821 -147 9871 -113
rect 9855 -181 9871 -147
rect 9821 -223 9871 -181
rect 9961 -78 10027 -29
rect 9961 -112 9977 -78
rect 10011 -112 10027 -78
rect 9961 -146 10027 -112
rect 9961 -180 9977 -146
rect 10011 -180 10027 -146
rect 9961 -189 10027 -180
rect 10061 -79 10142 -63
rect 10061 -113 10075 -79
rect 10109 -113 10142 -79
rect 10061 -147 10142 -113
rect 10061 -181 10075 -147
rect 10109 -181 10142 -147
rect 10061 -218 10142 -181
rect 9821 -257 9939 -223
rect 9905 -291 9939 -257
rect 9164 -351 9260 -317
rect 9294 -351 9314 -317
rect 9440 -301 9530 -298
rect 9440 -335 9453 -301
rect 9487 -307 9530 -301
rect 9440 -341 9480 -335
rect 9514 -341 9530 -307
rect 9564 -307 9650 -293
rect 9564 -341 9600 -307
rect 9634 -341 9650 -307
rect 9564 -351 9650 -341
rect 9699 -307 9871 -292
rect 9699 -341 9821 -307
rect 9855 -341 9871 -307
rect 9699 -342 9871 -341
rect 9905 -307 10058 -291
rect 9905 -341 10021 -307
rect 10055 -341 10058 -307
rect 9564 -375 9634 -351
rect 8567 -486 8583 -452
rect 8533 -505 8583 -486
rect 8673 -452 8739 -436
rect 8673 -486 8689 -452
rect 8723 -486 8739 -452
rect 8673 -539 8739 -486
rect 8773 -452 8854 -428
rect 8773 -486 8787 -452
rect 8821 -486 8854 -452
rect 8773 -505 8854 -486
rect 8888 -411 8946 -394
rect 8888 -445 8900 -411
rect 8934 -445 8946 -411
rect 8888 -539 8946 -445
rect 8980 -437 9314 -385
rect 8980 -471 8998 -437
rect 9032 -471 9262 -437
rect 9296 -471 9314 -437
rect 8980 -539 9314 -471
rect 9348 -411 9406 -394
rect 9348 -445 9360 -411
rect 9394 -445 9406 -411
rect 9348 -539 9406 -445
rect 9440 -409 9634 -375
rect 9440 -452 9506 -409
rect 9440 -486 9459 -452
rect 9493 -486 9506 -452
rect 9440 -505 9506 -486
rect 9540 -452 9606 -443
rect 9540 -486 9556 -452
rect 9590 -486 9606 -452
rect 9540 -539 9606 -486
rect 9699 -452 9769 -342
rect 9905 -357 10058 -341
rect 10092 -300 10142 -218
rect 10176 -100 10234 -29
rect 10176 -134 10188 -100
rect 10222 -134 10234 -100
rect 10176 -193 10234 -134
rect 10176 -227 10188 -193
rect 10222 -227 10234 -193
rect 10176 -262 10234 -227
rect 10268 -71 10602 -29
rect 10268 -105 10286 -71
rect 10320 -105 10550 -71
rect 10584 -105 10602 -71
rect 10268 -173 10602 -105
rect 10268 -207 10286 -173
rect 10320 -207 10550 -173
rect 10584 -207 10602 -173
rect 10268 -247 10602 -207
rect 10092 -334 10099 -300
rect 10133 -334 10142 -300
rect 9905 -376 9939 -357
rect 9699 -486 9716 -452
rect 9750 -486 9769 -452
rect 9699 -505 9769 -486
rect 9821 -410 9939 -376
rect 9821 -452 9871 -410
rect 10092 -428 10142 -334
rect 10268 -315 10288 -281
rect 10322 -315 10418 -281
rect 10268 -385 10418 -315
rect 10452 -317 10602 -247
rect 10636 -100 10694 -29
rect 10636 -134 10648 -100
rect 10682 -134 10694 -100
rect 10636 -193 10694 -134
rect 10636 -227 10648 -193
rect 10682 -227 10694 -193
rect 10636 -262 10694 -227
rect 10729 -71 10780 -29
rect 10729 -105 10746 -71
rect 10729 -139 10780 -105
rect 10729 -173 10746 -139
rect 10729 -207 10780 -173
rect 10729 -241 10746 -207
rect 10729 -257 10780 -241
rect 10814 -71 10880 -63
rect 10814 -105 10830 -71
rect 10864 -105 10880 -71
rect 10814 -139 10880 -105
rect 10814 -173 10830 -139
rect 10864 -173 10880 -139
rect 10814 -207 10880 -173
rect 10914 -71 10948 -29
rect 10914 -139 10948 -105
rect 10914 -189 10948 -173
rect 10982 -71 11048 -63
rect 10982 -105 10998 -71
rect 11032 -105 11048 -71
rect 10982 -139 11048 -105
rect 10982 -173 10998 -139
rect 11032 -173 11048 -139
rect 10814 -241 10830 -207
rect 10864 -223 10880 -207
rect 10982 -207 11048 -173
rect 11082 -71 11116 -29
rect 11082 -139 11116 -105
rect 11082 -189 11116 -173
rect 11150 -71 11216 -63
rect 11150 -105 11166 -71
rect 11200 -105 11216 -71
rect 11150 -139 11216 -105
rect 11150 -173 11166 -139
rect 11200 -173 11216 -139
rect 10982 -223 10998 -207
rect 10864 -241 10998 -223
rect 11032 -223 11048 -207
rect 11150 -207 11216 -173
rect 11250 -71 11284 -29
rect 11250 -139 11284 -105
rect 11250 -189 11284 -173
rect 11318 -71 11384 -63
rect 11318 -105 11334 -71
rect 11368 -105 11384 -71
rect 11318 -139 11384 -105
rect 11318 -173 11334 -139
rect 11368 -173 11384 -139
rect 11150 -223 11166 -207
rect 11032 -241 11166 -223
rect 11200 -223 11216 -207
rect 11318 -207 11384 -173
rect 11418 -71 11468 -29
rect 11452 -105 11468 -71
rect 11418 -139 11468 -105
rect 11452 -173 11468 -139
rect 11418 -189 11468 -173
rect 11556 -100 11614 -29
rect 11556 -134 11568 -100
rect 11602 -134 11614 -100
rect 11318 -223 11334 -207
rect 11200 -241 11334 -223
rect 11368 -241 11384 -207
rect 10814 -257 11384 -241
rect 11556 -193 11614 -134
rect 11556 -227 11568 -193
rect 11602 -227 11614 -193
rect 11093 -268 11200 -257
rect 11556 -262 11614 -227
rect 11648 -71 11982 -29
rect 11648 -105 11666 -71
rect 11700 -105 11930 -71
rect 11964 -105 11982 -71
rect 11648 -173 11982 -105
rect 11648 -207 11666 -173
rect 11700 -207 11930 -173
rect 11964 -207 11982 -173
rect 11648 -247 11982 -207
rect 10452 -351 10548 -317
rect 10582 -351 10602 -317
rect 10733 -301 11057 -291
rect 10733 -335 10741 -301
rect 10775 -307 10832 -301
rect 10866 -302 11057 -301
rect 10866 -307 10925 -302
rect 10959 -307 11017 -302
rect 10733 -341 10749 -335
rect 10783 -341 10830 -307
rect 10866 -335 10914 -307
rect 10864 -341 10914 -335
rect 10959 -336 10998 -307
rect 11051 -336 11057 -302
rect 10948 -341 10998 -336
rect 11032 -341 11057 -336
rect 11093 -302 11129 -268
rect 11163 -302 11200 -268
rect 11093 -341 11200 -302
rect 11234 -299 11522 -291
rect 11234 -341 11250 -299
rect 11284 -307 11344 -299
rect 11284 -341 11334 -307
rect 11378 -333 11522 -299
rect 11368 -341 11522 -333
rect 11648 -315 11668 -281
rect 11702 -315 11798 -281
rect 9855 -486 9871 -452
rect 9821 -505 9871 -486
rect 9961 -452 10027 -436
rect 9961 -486 9977 -452
rect 10011 -486 10027 -452
rect 9961 -539 10027 -486
rect 10061 -452 10142 -428
rect 10061 -486 10075 -452
rect 10109 -486 10142 -452
rect 10061 -505 10142 -486
rect 10176 -411 10234 -394
rect 10176 -445 10188 -411
rect 10222 -445 10234 -411
rect 10176 -539 10234 -445
rect 10268 -437 10602 -385
rect 10268 -471 10286 -437
rect 10320 -471 10550 -437
rect 10584 -471 10602 -437
rect 10268 -539 10602 -471
rect 10636 -411 10694 -394
rect 10636 -445 10648 -411
rect 10682 -445 10694 -411
rect 10636 -539 10694 -445
rect 10729 -395 11116 -375
rect 10729 -429 10746 -395
rect 10780 -413 10914 -395
rect 10780 -429 10796 -413
rect 10729 -463 10796 -429
rect 10898 -429 10914 -413
rect 10948 -413 11082 -395
rect 10948 -429 10964 -413
rect 10729 -497 10746 -463
rect 10780 -497 10796 -463
rect 10729 -505 10796 -497
rect 10830 -463 10864 -447
rect 10830 -539 10864 -497
rect 10898 -463 10964 -429
rect 11066 -429 11082 -413
rect 11150 -395 11200 -341
rect 11418 -395 11468 -379
rect 11648 -385 11798 -315
rect 11832 -317 11982 -247
rect 13488 -100 13546 -29
rect 13488 -134 13500 -100
rect 13534 -134 13546 -100
rect 13488 -193 13546 -134
rect 13488 -227 13500 -193
rect 13534 -227 13546 -193
rect 13488 -262 13546 -227
rect 13580 -71 14649 -29
rect 13580 -105 13598 -71
rect 13632 -105 14598 -71
rect 14632 -105 14649 -71
rect 13580 -173 14649 -105
rect 13580 -207 13598 -173
rect 13632 -207 14598 -173
rect 14632 -207 14649 -173
rect 13580 -247 14649 -207
rect 11832 -351 11928 -317
rect 11962 -351 11982 -317
rect 13580 -315 13658 -281
rect 13692 -315 13786 -281
rect 13820 -315 13914 -281
rect 13948 -315 14042 -281
rect 14076 -315 14096 -281
rect 13580 -385 14096 -315
rect 14130 -317 14649 -247
rect 14684 -100 14742 -29
rect 14684 -134 14696 -100
rect 14730 -134 14742 -100
rect 14684 -193 14742 -134
rect 14684 -227 14696 -193
rect 14730 -227 14742 -193
rect 14684 -262 14742 -227
rect 14776 -71 15845 -29
rect 14776 -105 14794 -71
rect 14828 -105 15794 -71
rect 15828 -105 15845 -71
rect 14776 -173 15845 -105
rect 14776 -207 14794 -173
rect 14828 -207 15794 -173
rect 15828 -207 15845 -173
rect 14776 -247 15845 -207
rect 14130 -351 14150 -317
rect 14184 -351 14278 -317
rect 14312 -351 14406 -317
rect 14440 -351 14534 -317
rect 14568 -351 14649 -317
rect 14776 -315 14854 -281
rect 14888 -315 14982 -281
rect 15016 -315 15110 -281
rect 15144 -315 15238 -281
rect 15272 -315 15292 -281
rect 14776 -385 15292 -315
rect 15326 -317 15845 -247
rect 15880 -100 15938 -29
rect 15880 -134 15892 -100
rect 15926 -134 15938 -100
rect 15880 -193 15938 -134
rect 15880 -227 15892 -193
rect 15926 -227 15938 -193
rect 15880 -262 15938 -227
rect 15972 -71 16674 -29
rect 15972 -105 15990 -71
rect 16024 -105 16622 -71
rect 16656 -105 16674 -71
rect 15972 -173 16674 -105
rect 15972 -207 15990 -173
rect 16024 -207 16622 -173
rect 16656 -207 16674 -173
rect 15972 -247 16674 -207
rect 15326 -351 15346 -317
rect 15380 -351 15474 -317
rect 15508 -351 15602 -317
rect 15636 -351 15730 -317
rect 15764 -351 15845 -317
rect 15972 -315 16050 -281
rect 16084 -315 16149 -281
rect 16183 -315 16248 -281
rect 16282 -315 16302 -281
rect 15972 -385 16302 -315
rect 16336 -317 16674 -247
rect 16336 -351 16356 -317
rect 16390 -351 16459 -317
rect 16493 -351 16562 -317
rect 16596 -351 16674 -317
rect 11150 -429 11166 -395
rect 11200 -429 11334 -395
rect 11368 -429 11384 -395
rect 11452 -429 11468 -395
rect 10898 -497 10914 -463
rect 10948 -497 10964 -463
rect 10898 -505 10964 -497
rect 10998 -463 11032 -447
rect 10998 -539 11032 -497
rect 11066 -463 11116 -429
rect 11418 -463 11468 -429
rect 11066 -497 11082 -463
rect 11116 -497 11250 -463
rect 11284 -497 11418 -463
rect 11452 -497 11468 -463
rect 11066 -505 11468 -497
rect 11556 -411 11614 -394
rect 11556 -445 11568 -411
rect 11602 -445 11614 -411
rect 11556 -539 11614 -445
rect 11648 -437 11982 -385
rect 11648 -471 11666 -437
rect 11700 -471 11930 -437
rect 11964 -471 11982 -437
rect 11648 -539 11982 -471
rect 13488 -411 13546 -394
rect 13488 -445 13500 -411
rect 13534 -445 13546 -411
rect 13488 -539 13546 -445
rect 13580 -444 14649 -385
rect 13580 -478 13598 -444
rect 13632 -478 14598 -444
rect 14632 -478 14649 -444
rect 13580 -539 14649 -478
rect 14684 -411 14742 -394
rect 14684 -445 14696 -411
rect 14730 -445 14742 -411
rect 14684 -539 14742 -445
rect 14776 -444 15845 -385
rect 14776 -478 14794 -444
rect 14828 -478 15794 -444
rect 15828 -478 15845 -444
rect 14776 -539 15845 -478
rect 15880 -411 15938 -394
rect 15880 -445 15892 -411
rect 15926 -445 15938 -411
rect 15880 -539 15938 -445
rect 15972 -444 16674 -385
rect 15972 -478 15990 -444
rect 16024 -478 16622 -444
rect 16656 -478 16674 -444
rect 15972 -539 16674 -478
rect -2997 -573 -2968 -539
rect -2934 -573 -2876 -539
rect -2842 -573 -2784 -539
rect -2750 -573 -2692 -539
rect -2658 -573 -2600 -539
rect -2566 -573 -2508 -539
rect -2474 -573 -2416 -539
rect -2382 -573 -2324 -539
rect -2290 -573 -2232 -539
rect -2198 -573 -2140 -539
rect -2106 -573 -2048 -539
rect -2014 -573 -1956 -539
rect -1922 -573 -1864 -539
rect -1830 -573 -1772 -539
rect -1738 -573 -1680 -539
rect -1646 -573 -1588 -539
rect -1554 -573 -1496 -539
rect -1462 -573 -1404 -539
rect -1370 -573 -1312 -539
rect -1278 -573 -1220 -539
rect -1186 -573 -1128 -539
rect -1094 -573 -1036 -539
rect -1002 -573 -944 -539
rect -910 -573 -852 -539
rect -818 -573 -760 -539
rect -726 -573 -668 -539
rect -634 -573 -576 -539
rect -542 -573 -484 -539
rect -450 -573 -392 -539
rect -358 -573 -300 -539
rect -266 -573 -208 -539
rect -174 -573 -116 -539
rect -82 -573 -24 -539
rect 10 -573 68 -539
rect 102 -573 160 -539
rect 194 -573 252 -539
rect 286 -573 344 -539
rect 378 -573 436 -539
rect 470 -573 528 -539
rect 562 -573 620 -539
rect 654 -573 712 -539
rect 746 -573 804 -539
rect 838 -573 896 -539
rect 930 -573 988 -539
rect 1022 -573 1080 -539
rect 1114 -573 1172 -539
rect 1206 -573 1264 -539
rect 1298 -573 1356 -539
rect 1390 -573 1448 -539
rect 1482 -573 1540 -539
rect 1574 -573 1632 -539
rect 1666 -573 1724 -539
rect 1758 -573 1816 -539
rect 1850 -573 1908 -539
rect 1942 -573 2000 -539
rect 2034 -573 2092 -539
rect 2126 -573 2184 -539
rect 2218 -573 2276 -539
rect 2310 -573 2368 -539
rect 2402 -573 2460 -539
rect 2494 -573 2552 -539
rect 2586 -573 2644 -539
rect 2678 -573 2736 -539
rect 2770 -573 2828 -539
rect 2862 -573 2920 -539
rect 2954 -573 3012 -539
rect 3046 -573 3104 -539
rect 3138 -573 3196 -539
rect 3230 -573 3288 -539
rect 3322 -573 3380 -539
rect 3414 -573 3472 -539
rect 3506 -573 3564 -539
rect 3598 -573 3656 -539
rect 3690 -573 3748 -539
rect 3782 -573 3840 -539
rect 3874 -573 3932 -539
rect 3966 -573 4024 -539
rect 4058 -573 4116 -539
rect 4150 -573 4208 -539
rect 4242 -573 4300 -539
rect 4334 -573 4392 -539
rect 4426 -573 4484 -539
rect 4518 -573 4576 -539
rect 4610 -573 4668 -539
rect 4702 -573 4760 -539
rect 4794 -573 4852 -539
rect 4886 -573 4944 -539
rect 4978 -573 5036 -539
rect 5070 -573 5128 -539
rect 5162 -573 5220 -539
rect 5254 -573 5312 -539
rect 5346 -573 5404 -539
rect 5438 -573 5496 -539
rect 5530 -573 5588 -539
rect 5622 -573 5680 -539
rect 5714 -573 5772 -539
rect 5806 -573 5864 -539
rect 5898 -573 5956 -539
rect 5990 -573 6048 -539
rect 6082 -573 6140 -539
rect 6174 -573 6232 -539
rect 6266 -573 6324 -539
rect 6358 -573 6416 -539
rect 6450 -573 6508 -539
rect 6542 -573 6600 -539
rect 6634 -573 6692 -539
rect 6726 -573 6784 -539
rect 6818 -573 6876 -539
rect 6910 -573 6968 -539
rect 7002 -573 7060 -539
rect 7094 -573 7152 -539
rect 7186 -573 7244 -539
rect 7278 -573 7336 -539
rect 7370 -573 7428 -539
rect 7462 -573 7520 -539
rect 7554 -573 7612 -539
rect 7646 -573 7704 -539
rect 7738 -573 7796 -539
rect 7830 -573 7888 -539
rect 7922 -573 7980 -539
rect 8014 -573 8072 -539
rect 8106 -573 8164 -539
rect 8198 -573 8256 -539
rect 8290 -573 8348 -539
rect 8382 -573 8440 -539
rect 8474 -573 8532 -539
rect 8566 -573 8624 -539
rect 8658 -573 8716 -539
rect 8750 -573 8808 -539
rect 8842 -573 8900 -539
rect 8934 -573 8992 -539
rect 9026 -573 9084 -539
rect 9118 -573 9176 -539
rect 9210 -573 9268 -539
rect 9302 -573 9360 -539
rect 9394 -573 9452 -539
rect 9486 -573 9544 -539
rect 9578 -573 9636 -539
rect 9670 -573 9728 -539
rect 9762 -573 9820 -539
rect 9854 -573 9912 -539
rect 9946 -573 10004 -539
rect 10038 -573 10096 -539
rect 10130 -573 10188 -539
rect 10222 -573 10280 -539
rect 10314 -573 10372 -539
rect 10406 -573 10464 -539
rect 10498 -573 10556 -539
rect 10590 -573 10648 -539
rect 10682 -573 10740 -539
rect 10774 -573 10832 -539
rect 10866 -573 10924 -539
rect 10958 -573 11016 -539
rect 11050 -573 11108 -539
rect 11142 -573 11200 -539
rect 11234 -573 11292 -539
rect 11326 -573 11384 -539
rect 11418 -573 11476 -539
rect 11510 -573 11568 -539
rect 11602 -573 11660 -539
rect 11694 -573 11752 -539
rect 11786 -573 11844 -539
rect 11878 -573 11936 -539
rect 11970 -573 12028 -539
rect 12062 -573 12120 -539
rect 12154 -573 12212 -539
rect 12246 -573 12304 -539
rect 12338 -573 12396 -539
rect 12430 -573 12488 -539
rect 12522 -573 12580 -539
rect 12614 -573 12672 -539
rect 12706 -573 12764 -539
rect 12798 -573 12856 -539
rect 12890 -573 12948 -539
rect 12982 -573 13040 -539
rect 13074 -573 13132 -539
rect 13166 -573 13224 -539
rect 13258 -573 13316 -539
rect 13350 -573 13408 -539
rect 13442 -573 13500 -539
rect 13534 -573 13592 -539
rect 13626 -573 13684 -539
rect 13718 -573 13776 -539
rect 13810 -573 13868 -539
rect 13902 -573 13960 -539
rect 13994 -573 14052 -539
rect 14086 -573 14144 -539
rect 14178 -573 14236 -539
rect 14270 -573 14328 -539
rect 14362 -573 14420 -539
rect 14454 -573 14512 -539
rect 14546 -573 14604 -539
rect 14638 -573 14696 -539
rect 14730 -573 14788 -539
rect 14822 -573 14880 -539
rect 14914 -573 14972 -539
rect 15006 -573 15064 -539
rect 15098 -573 15156 -539
rect 15190 -573 15248 -539
rect 15282 -573 15340 -539
rect 15374 -573 15432 -539
rect 15466 -573 15524 -539
rect 15558 -573 15616 -539
rect 15650 -573 15708 -539
rect 15742 -573 15800 -539
rect 15834 -573 15892 -539
rect 15926 -573 15984 -539
rect 16018 -573 16076 -539
rect 16110 -573 16168 -539
rect 16202 -573 16260 -539
rect 16294 -573 16352 -539
rect 16386 -573 16444 -539
rect 16478 -573 16536 -539
rect 16570 -573 16628 -539
rect 16662 -573 16691 -539
rect -2980 -634 -2278 -573
rect -2980 -668 -2962 -634
rect -2928 -668 -2330 -634
rect -2296 -668 -2278 -634
rect -2980 -727 -2278 -668
rect -2244 -667 -2186 -573
rect -2244 -701 -2232 -667
rect -2198 -701 -2186 -667
rect -2244 -718 -2186 -701
rect -1600 -634 -898 -573
rect -1600 -668 -1582 -634
rect -1548 -668 -950 -634
rect -916 -668 -898 -634
rect -1600 -727 -898 -668
rect -864 -634 -162 -573
rect -864 -668 -846 -634
rect -812 -668 -214 -634
rect -180 -668 -162 -634
rect -864 -727 -162 -668
rect -128 -667 -70 -573
rect -128 -701 -116 -667
rect -82 -701 -70 -667
rect -128 -718 -70 -701
rect -36 -641 298 -573
rect -36 -675 -18 -641
rect 16 -675 246 -641
rect 280 -675 298 -641
rect -36 -727 298 -675
rect 332 -667 390 -573
rect 332 -701 344 -667
rect 378 -701 390 -667
rect 332 -718 390 -701
rect 424 -626 505 -607
rect 424 -660 457 -626
rect 491 -660 505 -626
rect 424 -684 505 -660
rect 539 -626 605 -573
rect 539 -660 555 -626
rect 589 -660 605 -626
rect 539 -676 605 -660
rect 695 -626 745 -607
rect 695 -660 711 -626
rect -2980 -795 -2902 -761
rect -2868 -795 -2799 -761
rect -2765 -795 -2696 -761
rect -2662 -795 -2642 -761
rect -2980 -865 -2642 -795
rect -2608 -797 -2278 -727
rect -2608 -831 -2588 -797
rect -2554 -831 -2489 -797
rect -2455 -831 -2390 -797
rect -2356 -831 -2278 -797
rect -1600 -795 -1522 -761
rect -1488 -795 -1419 -761
rect -1385 -795 -1316 -761
rect -1282 -795 -1262 -761
rect -2980 -905 -2278 -865
rect -2980 -939 -2962 -905
rect -2928 -939 -2330 -905
rect -2296 -939 -2278 -905
rect -2980 -1007 -2278 -939
rect -2980 -1041 -2962 -1007
rect -2928 -1041 -2330 -1007
rect -2296 -1041 -2278 -1007
rect -2980 -1083 -2278 -1041
rect -2244 -885 -2186 -850
rect -2244 -919 -2232 -885
rect -2198 -919 -2186 -885
rect -2244 -978 -2186 -919
rect -2244 -1012 -2232 -978
rect -2198 -1012 -2186 -978
rect -2244 -1083 -2186 -1012
rect -1600 -865 -1262 -795
rect -1228 -797 -898 -727
rect -1228 -831 -1208 -797
rect -1174 -831 -1109 -797
rect -1075 -831 -1010 -797
rect -976 -831 -898 -797
rect -864 -795 -786 -761
rect -752 -795 -683 -761
rect -649 -795 -580 -761
rect -546 -795 -526 -761
rect -864 -865 -526 -795
rect -492 -797 -162 -727
rect -492 -831 -472 -797
rect -438 -831 -373 -797
rect -339 -831 -274 -797
rect -240 -831 -162 -797
rect -36 -795 -16 -761
rect 18 -795 114 -761
rect -1600 -905 -898 -865
rect -1600 -939 -1582 -905
rect -1548 -939 -950 -905
rect -916 -939 -898 -905
rect -1600 -1007 -898 -939
rect -1600 -1041 -1582 -1007
rect -1548 -1041 -950 -1007
rect -916 -1041 -898 -1007
rect -1600 -1083 -898 -1041
rect -864 -905 -162 -865
rect -864 -939 -846 -905
rect -812 -939 -214 -905
rect -180 -939 -162 -905
rect -864 -1007 -162 -939
rect -864 -1041 -846 -1007
rect -812 -1041 -214 -1007
rect -180 -1041 -162 -1007
rect -864 -1083 -162 -1041
rect -128 -885 -70 -850
rect -128 -919 -116 -885
rect -82 -919 -70 -885
rect -128 -978 -70 -919
rect -128 -1012 -116 -978
rect -82 -1012 -70 -978
rect -128 -1083 -70 -1012
rect -36 -865 114 -795
rect 148 -797 298 -727
rect 148 -831 244 -797
rect 278 -831 298 -797
rect 424 -812 474 -684
rect 695 -702 745 -660
rect 627 -736 745 -702
rect 797 -626 867 -607
rect 797 -660 816 -626
rect 850 -660 867 -626
rect 627 -755 661 -736
rect 424 -846 433 -812
rect 467 -846 474 -812
rect 508 -771 661 -755
rect 797 -770 867 -660
rect 960 -626 1026 -573
rect 960 -660 976 -626
rect 1010 -660 1026 -626
rect 960 -669 1026 -660
rect 1060 -626 1126 -607
rect 1060 -660 1073 -626
rect 1107 -660 1126 -626
rect 1060 -703 1126 -660
rect 932 -737 1126 -703
rect 1160 -667 1218 -573
rect 1160 -701 1172 -667
rect 1206 -701 1218 -667
rect 1160 -718 1218 -701
rect 1252 -641 1586 -573
rect 1252 -675 1270 -641
rect 1304 -675 1534 -641
rect 1568 -675 1586 -641
rect 1252 -727 1586 -675
rect 1620 -667 1678 -573
rect 1620 -701 1632 -667
rect 1666 -701 1678 -667
rect 1620 -718 1678 -701
rect 1712 -634 2414 -573
rect 1712 -668 1730 -634
rect 1764 -668 2362 -634
rect 2396 -668 2414 -634
rect 1712 -727 2414 -668
rect 2448 -667 2506 -573
rect 2448 -701 2460 -667
rect 2494 -701 2506 -667
rect 2448 -718 2506 -701
rect 2540 -641 2874 -573
rect 2540 -675 2558 -641
rect 2592 -675 2822 -641
rect 2856 -675 2874 -641
rect 2540 -727 2874 -675
rect 2908 -667 2966 -573
rect 2908 -701 2920 -667
rect 2954 -701 2966 -667
rect 2908 -718 2966 -701
rect 3000 -626 3081 -607
rect 3000 -660 3033 -626
rect 3067 -660 3081 -626
rect 3000 -684 3081 -660
rect 3115 -626 3181 -573
rect 3115 -660 3131 -626
rect 3165 -660 3181 -626
rect 3115 -676 3181 -660
rect 3271 -626 3321 -607
rect 3271 -660 3287 -626
rect 932 -761 1002 -737
rect 508 -805 511 -771
rect 545 -805 661 -771
rect 508 -821 661 -805
rect 695 -771 867 -770
rect 695 -805 711 -771
rect 745 -805 867 -771
rect 695 -820 867 -805
rect 916 -771 1002 -761
rect 916 -805 932 -771
rect 966 -805 1002 -771
rect 916 -819 1002 -805
rect 1036 -809 1052 -771
rect 1086 -809 1126 -771
rect 1036 -814 1126 -809
rect 1252 -795 1272 -761
rect 1306 -795 1402 -761
rect -36 -905 298 -865
rect -36 -939 -18 -905
rect 16 -939 246 -905
rect 280 -939 298 -905
rect -36 -1007 298 -939
rect -36 -1041 -18 -1007
rect 16 -1041 246 -1007
rect 280 -1041 298 -1007
rect -36 -1083 298 -1041
rect 332 -885 390 -850
rect 332 -919 344 -885
rect 378 -919 390 -885
rect 332 -978 390 -919
rect 332 -1012 344 -978
rect 378 -1012 390 -978
rect 332 -1083 390 -1012
rect 424 -894 474 -846
rect 627 -855 661 -821
rect 627 -889 745 -855
rect 424 -931 505 -894
rect 424 -965 457 -931
rect 491 -965 505 -931
rect 424 -999 505 -965
rect 424 -1033 457 -999
rect 491 -1033 505 -999
rect 424 -1049 505 -1033
rect 539 -932 605 -923
rect 539 -966 555 -932
rect 589 -966 605 -932
rect 539 -1000 605 -966
rect 539 -1034 555 -1000
rect 589 -1034 605 -1000
rect 539 -1083 605 -1034
rect 695 -931 745 -889
rect 695 -965 711 -931
rect 695 -999 745 -965
rect 695 -1033 711 -999
rect 695 -1049 745 -1033
rect 797 -932 867 -820
rect 932 -848 1002 -819
rect 932 -882 1126 -848
rect 797 -966 815 -932
rect 849 -966 867 -932
rect 797 -1000 867 -966
rect 797 -1034 815 -1000
rect 849 -1034 867 -1000
rect 797 -1049 867 -1034
rect 957 -932 1023 -916
rect 957 -966 973 -932
rect 1007 -966 1023 -932
rect 957 -1000 1023 -966
rect 957 -1034 973 -1000
rect 1007 -1034 1023 -1000
rect 957 -1083 1023 -1034
rect 1057 -932 1126 -882
rect 1057 -966 1073 -932
rect 1107 -966 1126 -932
rect 1057 -1000 1126 -966
rect 1057 -1034 1073 -1000
rect 1107 -1034 1126 -1000
rect 1057 -1049 1126 -1034
rect 1160 -885 1218 -850
rect 1160 -919 1172 -885
rect 1206 -919 1218 -885
rect 1160 -978 1218 -919
rect 1160 -1012 1172 -978
rect 1206 -1012 1218 -978
rect 1160 -1083 1218 -1012
rect 1252 -865 1402 -795
rect 1436 -797 1586 -727
rect 1436 -831 1532 -797
rect 1566 -831 1586 -797
rect 1712 -795 1790 -761
rect 1824 -795 1893 -761
rect 1927 -795 1996 -761
rect 2030 -795 2050 -761
rect 1252 -905 1586 -865
rect 1252 -939 1270 -905
rect 1304 -939 1534 -905
rect 1568 -939 1586 -905
rect 1252 -1007 1586 -939
rect 1252 -1041 1270 -1007
rect 1304 -1041 1534 -1007
rect 1568 -1041 1586 -1007
rect 1252 -1083 1586 -1041
rect 1620 -885 1678 -850
rect 1620 -919 1632 -885
rect 1666 -919 1678 -885
rect 1620 -978 1678 -919
rect 1620 -1012 1632 -978
rect 1666 -1012 1678 -978
rect 1620 -1083 1678 -1012
rect 1712 -865 2050 -795
rect 2084 -797 2414 -727
rect 2084 -831 2104 -797
rect 2138 -831 2203 -797
rect 2237 -831 2302 -797
rect 2336 -831 2414 -797
rect 2540 -795 2560 -761
rect 2594 -795 2690 -761
rect 1712 -905 2414 -865
rect 1712 -939 1730 -905
rect 1764 -939 2362 -905
rect 2396 -939 2414 -905
rect 1712 -1007 2414 -939
rect 1712 -1041 1730 -1007
rect 1764 -1041 2362 -1007
rect 2396 -1041 2414 -1007
rect 1712 -1083 2414 -1041
rect 2448 -885 2506 -850
rect 2448 -919 2460 -885
rect 2494 -919 2506 -885
rect 2448 -978 2506 -919
rect 2448 -1012 2460 -978
rect 2494 -1012 2506 -978
rect 2448 -1083 2506 -1012
rect 2540 -865 2690 -795
rect 2724 -797 2874 -727
rect 2724 -831 2820 -797
rect 2854 -831 2874 -797
rect 3000 -775 3050 -684
rect 3271 -702 3321 -660
rect 3203 -736 3321 -702
rect 3373 -626 3443 -607
rect 3373 -660 3392 -626
rect 3426 -660 3443 -626
rect 3203 -755 3237 -736
rect 3000 -809 3012 -775
rect 3046 -809 3050 -775
rect 2540 -905 2874 -865
rect 2540 -939 2558 -905
rect 2592 -939 2822 -905
rect 2856 -939 2874 -905
rect 2540 -1007 2874 -939
rect 2540 -1041 2558 -1007
rect 2592 -1041 2822 -1007
rect 2856 -1041 2874 -1007
rect 2540 -1083 2874 -1041
rect 2908 -885 2966 -850
rect 2908 -919 2920 -885
rect 2954 -919 2966 -885
rect 2908 -978 2966 -919
rect 2908 -1012 2920 -978
rect 2954 -1012 2966 -978
rect 2908 -1083 2966 -1012
rect 3000 -894 3050 -809
rect 3084 -771 3237 -755
rect 3373 -770 3443 -660
rect 3536 -626 3602 -573
rect 3536 -660 3552 -626
rect 3586 -660 3602 -626
rect 3536 -669 3602 -660
rect 3636 -626 3702 -607
rect 3636 -660 3649 -626
rect 3683 -660 3702 -626
rect 3636 -703 3702 -660
rect 3508 -737 3702 -703
rect 3736 -667 3794 -573
rect 3736 -701 3748 -667
rect 3782 -701 3794 -667
rect 3736 -718 3794 -701
rect 3828 -641 4162 -573
rect 3828 -675 3846 -641
rect 3880 -675 4110 -641
rect 4144 -675 4162 -641
rect 3828 -727 4162 -675
rect 4196 -667 4254 -573
rect 4196 -701 4208 -667
rect 4242 -701 4254 -667
rect 4196 -718 4254 -701
rect 4288 -634 4990 -573
rect 4288 -668 4306 -634
rect 4340 -668 4938 -634
rect 4972 -668 4990 -634
rect 4288 -727 4990 -668
rect 5024 -667 5082 -573
rect 5024 -701 5036 -667
rect 5070 -701 5082 -667
rect 5024 -718 5082 -701
rect 5116 -641 5450 -573
rect 5116 -675 5134 -641
rect 5168 -675 5398 -641
rect 5432 -675 5450 -641
rect 5116 -727 5450 -675
rect 5484 -667 5542 -573
rect 5484 -701 5496 -667
rect 5530 -701 5542 -667
rect 5484 -718 5542 -701
rect 5576 -626 5657 -607
rect 5576 -660 5609 -626
rect 5643 -660 5657 -626
rect 5576 -684 5657 -660
rect 5691 -626 5757 -573
rect 5691 -660 5707 -626
rect 5741 -660 5757 -626
rect 5691 -676 5757 -660
rect 5847 -626 5897 -607
rect 5847 -660 5863 -626
rect 3508 -761 3578 -737
rect 3084 -805 3087 -771
rect 3121 -805 3237 -771
rect 3084 -821 3237 -805
rect 3271 -771 3443 -770
rect 3271 -805 3287 -771
rect 3321 -805 3443 -771
rect 3271 -820 3443 -805
rect 3492 -771 3578 -761
rect 3492 -805 3508 -771
rect 3542 -805 3578 -771
rect 3492 -819 3578 -805
rect 3612 -775 3628 -771
rect 3612 -809 3626 -775
rect 3662 -805 3702 -771
rect 3660 -809 3702 -805
rect 3612 -814 3702 -809
rect 3828 -795 3848 -761
rect 3882 -795 3978 -761
rect 3203 -855 3237 -821
rect 3203 -889 3321 -855
rect 3000 -931 3081 -894
rect 3000 -965 3033 -931
rect 3067 -965 3081 -931
rect 3000 -999 3081 -965
rect 3000 -1033 3033 -999
rect 3067 -1033 3081 -999
rect 3000 -1049 3081 -1033
rect 3115 -932 3181 -923
rect 3115 -966 3131 -932
rect 3165 -966 3181 -932
rect 3115 -1000 3181 -966
rect 3115 -1034 3131 -1000
rect 3165 -1034 3181 -1000
rect 3115 -1083 3181 -1034
rect 3271 -931 3321 -889
rect 3271 -965 3287 -931
rect 3271 -999 3321 -965
rect 3271 -1033 3287 -999
rect 3271 -1049 3321 -1033
rect 3373 -932 3443 -820
rect 3508 -848 3578 -819
rect 3508 -882 3702 -848
rect 3373 -966 3391 -932
rect 3425 -966 3443 -932
rect 3373 -1000 3443 -966
rect 3373 -1034 3391 -1000
rect 3425 -1034 3443 -1000
rect 3373 -1049 3443 -1034
rect 3533 -932 3599 -916
rect 3533 -966 3549 -932
rect 3583 -966 3599 -932
rect 3533 -1000 3599 -966
rect 3533 -1034 3549 -1000
rect 3583 -1034 3599 -1000
rect 3533 -1083 3599 -1034
rect 3633 -932 3702 -882
rect 3633 -966 3649 -932
rect 3683 -966 3702 -932
rect 3633 -1000 3702 -966
rect 3633 -1034 3649 -1000
rect 3683 -1034 3702 -1000
rect 3633 -1049 3702 -1034
rect 3736 -885 3794 -850
rect 3736 -919 3748 -885
rect 3782 -919 3794 -885
rect 3736 -978 3794 -919
rect 3736 -1012 3748 -978
rect 3782 -1012 3794 -978
rect 3736 -1083 3794 -1012
rect 3828 -865 3978 -795
rect 4012 -797 4162 -727
rect 4012 -831 4108 -797
rect 4142 -831 4162 -797
rect 4288 -795 4366 -761
rect 4400 -795 4469 -761
rect 4503 -795 4572 -761
rect 4606 -795 4626 -761
rect 3828 -905 4162 -865
rect 3828 -939 3846 -905
rect 3880 -939 4110 -905
rect 4144 -939 4162 -905
rect 3828 -1007 4162 -939
rect 3828 -1041 3846 -1007
rect 3880 -1041 4110 -1007
rect 4144 -1041 4162 -1007
rect 3828 -1083 4162 -1041
rect 4196 -885 4254 -850
rect 4196 -919 4208 -885
rect 4242 -919 4254 -885
rect 4196 -978 4254 -919
rect 4196 -1012 4208 -978
rect 4242 -1012 4254 -978
rect 4196 -1083 4254 -1012
rect 4288 -865 4626 -795
rect 4660 -797 4990 -727
rect 4660 -831 4680 -797
rect 4714 -831 4779 -797
rect 4813 -831 4878 -797
rect 4912 -831 4990 -797
rect 5116 -795 5136 -761
rect 5170 -795 5266 -761
rect 4288 -905 4990 -865
rect 4288 -939 4306 -905
rect 4340 -939 4938 -905
rect 4972 -939 4990 -905
rect 4288 -1007 4990 -939
rect 4288 -1041 4306 -1007
rect 4340 -1041 4938 -1007
rect 4972 -1041 4990 -1007
rect 4288 -1083 4990 -1041
rect 5024 -885 5082 -850
rect 5024 -919 5036 -885
rect 5070 -919 5082 -885
rect 5024 -978 5082 -919
rect 5024 -1012 5036 -978
rect 5070 -1012 5082 -978
rect 5024 -1083 5082 -1012
rect 5116 -865 5266 -795
rect 5300 -797 5450 -727
rect 5300 -831 5396 -797
rect 5430 -831 5450 -797
rect 5576 -775 5626 -684
rect 5847 -702 5897 -660
rect 5779 -736 5897 -702
rect 5949 -626 6019 -607
rect 5949 -660 5968 -626
rect 6002 -660 6019 -626
rect 5779 -755 5813 -736
rect 5576 -809 5586 -775
rect 5620 -809 5626 -775
rect 5116 -905 5450 -865
rect 5116 -939 5134 -905
rect 5168 -939 5398 -905
rect 5432 -939 5450 -905
rect 5116 -1007 5450 -939
rect 5116 -1041 5134 -1007
rect 5168 -1041 5398 -1007
rect 5432 -1041 5450 -1007
rect 5116 -1083 5450 -1041
rect 5484 -885 5542 -850
rect 5484 -919 5496 -885
rect 5530 -919 5542 -885
rect 5484 -978 5542 -919
rect 5484 -1012 5496 -978
rect 5530 -1012 5542 -978
rect 5484 -1083 5542 -1012
rect 5576 -894 5626 -809
rect 5660 -771 5813 -755
rect 5949 -770 6019 -660
rect 6112 -626 6178 -573
rect 6112 -660 6128 -626
rect 6162 -660 6178 -626
rect 6112 -669 6178 -660
rect 6212 -626 6278 -607
rect 6212 -660 6225 -626
rect 6259 -660 6278 -626
rect 6212 -703 6278 -660
rect 6084 -737 6278 -703
rect 6312 -667 6370 -573
rect 6312 -701 6324 -667
rect 6358 -701 6370 -667
rect 6312 -718 6370 -701
rect 6404 -641 6738 -573
rect 6404 -675 6422 -641
rect 6456 -675 6686 -641
rect 6720 -675 6738 -641
rect 6404 -727 6738 -675
rect 6772 -667 6830 -573
rect 6772 -701 6784 -667
rect 6818 -701 6830 -667
rect 6772 -718 6830 -701
rect 6864 -634 7566 -573
rect 6864 -668 6882 -634
rect 6916 -668 7514 -634
rect 7548 -668 7566 -634
rect 6864 -727 7566 -668
rect 7600 -667 7658 -573
rect 7600 -701 7612 -667
rect 7646 -701 7658 -667
rect 7600 -718 7658 -701
rect 7692 -641 8026 -573
rect 7692 -675 7710 -641
rect 7744 -675 7974 -641
rect 8008 -675 8026 -641
rect 7692 -727 8026 -675
rect 8060 -667 8118 -573
rect 8060 -701 8072 -667
rect 8106 -701 8118 -667
rect 8060 -718 8118 -701
rect 8152 -626 8233 -607
rect 8152 -660 8185 -626
rect 8219 -660 8233 -626
rect 8152 -684 8233 -660
rect 8267 -626 8333 -573
rect 8267 -660 8283 -626
rect 8317 -660 8333 -626
rect 8267 -676 8333 -660
rect 8423 -626 8473 -607
rect 8423 -660 8439 -626
rect 6084 -761 6154 -737
rect 5660 -805 5663 -771
rect 5697 -805 5813 -771
rect 5660 -821 5813 -805
rect 5847 -771 6019 -770
rect 5847 -805 5863 -771
rect 5897 -805 6019 -771
rect 5847 -820 6019 -805
rect 6068 -771 6154 -761
rect 6068 -805 6084 -771
rect 6118 -805 6154 -771
rect 6068 -819 6154 -805
rect 6188 -775 6204 -771
rect 6188 -809 6200 -775
rect 6238 -805 6278 -771
rect 6234 -809 6278 -805
rect 6188 -814 6278 -809
rect 6404 -795 6424 -761
rect 6458 -795 6554 -761
rect 5779 -855 5813 -821
rect 5779 -889 5897 -855
rect 5576 -931 5657 -894
rect 5576 -965 5609 -931
rect 5643 -965 5657 -931
rect 5576 -999 5657 -965
rect 5576 -1033 5609 -999
rect 5643 -1033 5657 -999
rect 5576 -1049 5657 -1033
rect 5691 -932 5757 -923
rect 5691 -966 5707 -932
rect 5741 -966 5757 -932
rect 5691 -1000 5757 -966
rect 5691 -1034 5707 -1000
rect 5741 -1034 5757 -1000
rect 5691 -1083 5757 -1034
rect 5847 -931 5897 -889
rect 5847 -965 5863 -931
rect 5847 -999 5897 -965
rect 5847 -1033 5863 -999
rect 5847 -1049 5897 -1033
rect 5949 -932 6019 -820
rect 6084 -848 6154 -819
rect 6084 -882 6278 -848
rect 5949 -966 5967 -932
rect 6001 -966 6019 -932
rect 5949 -1000 6019 -966
rect 5949 -1034 5967 -1000
rect 6001 -1034 6019 -1000
rect 5949 -1049 6019 -1034
rect 6109 -932 6175 -916
rect 6109 -966 6125 -932
rect 6159 -966 6175 -932
rect 6109 -1000 6175 -966
rect 6109 -1034 6125 -1000
rect 6159 -1034 6175 -1000
rect 6109 -1083 6175 -1034
rect 6209 -932 6278 -882
rect 6209 -966 6225 -932
rect 6259 -966 6278 -932
rect 6209 -1000 6278 -966
rect 6209 -1034 6225 -1000
rect 6259 -1034 6278 -1000
rect 6209 -1049 6278 -1034
rect 6312 -885 6370 -850
rect 6312 -919 6324 -885
rect 6358 -919 6370 -885
rect 6312 -978 6370 -919
rect 6312 -1012 6324 -978
rect 6358 -1012 6370 -978
rect 6312 -1083 6370 -1012
rect 6404 -865 6554 -795
rect 6588 -797 6738 -727
rect 6588 -831 6684 -797
rect 6718 -831 6738 -797
rect 6864 -795 6942 -761
rect 6976 -795 7045 -761
rect 7079 -795 7148 -761
rect 7182 -795 7202 -761
rect 6404 -905 6738 -865
rect 6404 -939 6422 -905
rect 6456 -939 6686 -905
rect 6720 -939 6738 -905
rect 6404 -1007 6738 -939
rect 6404 -1041 6422 -1007
rect 6456 -1041 6686 -1007
rect 6720 -1041 6738 -1007
rect 6404 -1083 6738 -1041
rect 6772 -885 6830 -850
rect 6772 -919 6784 -885
rect 6818 -919 6830 -885
rect 6772 -978 6830 -919
rect 6772 -1012 6784 -978
rect 6818 -1012 6830 -978
rect 6772 -1083 6830 -1012
rect 6864 -865 7202 -795
rect 7236 -797 7566 -727
rect 7236 -831 7256 -797
rect 7290 -831 7355 -797
rect 7389 -831 7454 -797
rect 7488 -831 7566 -797
rect 7692 -795 7712 -761
rect 7746 -795 7842 -761
rect 6864 -905 7566 -865
rect 6864 -939 6882 -905
rect 6916 -939 7514 -905
rect 7548 -939 7566 -905
rect 6864 -1007 7566 -939
rect 6864 -1041 6882 -1007
rect 6916 -1041 7514 -1007
rect 7548 -1041 7566 -1007
rect 6864 -1083 7566 -1041
rect 7600 -885 7658 -850
rect 7600 -919 7612 -885
rect 7646 -919 7658 -885
rect 7600 -978 7658 -919
rect 7600 -1012 7612 -978
rect 7646 -1012 7658 -978
rect 7600 -1083 7658 -1012
rect 7692 -865 7842 -795
rect 7876 -797 8026 -727
rect 7876 -831 7972 -797
rect 8006 -831 8026 -797
rect 8152 -775 8202 -684
rect 8423 -702 8473 -660
rect 8355 -736 8473 -702
rect 8525 -626 8595 -607
rect 8525 -660 8544 -626
rect 8578 -660 8595 -626
rect 8355 -755 8389 -736
rect 8152 -809 8160 -775
rect 8194 -809 8202 -775
rect 7692 -905 8026 -865
rect 7692 -939 7710 -905
rect 7744 -939 7974 -905
rect 8008 -939 8026 -905
rect 7692 -1007 8026 -939
rect 7692 -1041 7710 -1007
rect 7744 -1041 7974 -1007
rect 8008 -1041 8026 -1007
rect 7692 -1083 8026 -1041
rect 8060 -885 8118 -850
rect 8060 -919 8072 -885
rect 8106 -919 8118 -885
rect 8060 -978 8118 -919
rect 8060 -1012 8072 -978
rect 8106 -1012 8118 -978
rect 8060 -1083 8118 -1012
rect 8152 -894 8202 -809
rect 8236 -771 8389 -755
rect 8525 -770 8595 -660
rect 8688 -626 8754 -573
rect 8688 -660 8704 -626
rect 8738 -660 8754 -626
rect 8688 -669 8754 -660
rect 8788 -626 8854 -607
rect 8788 -660 8801 -626
rect 8835 -660 8854 -626
rect 8788 -703 8854 -660
rect 8660 -737 8854 -703
rect 8888 -667 8946 -573
rect 8888 -701 8900 -667
rect 8934 -701 8946 -667
rect 8888 -718 8946 -701
rect 8980 -641 9314 -573
rect 8980 -675 8998 -641
rect 9032 -675 9262 -641
rect 9296 -675 9314 -641
rect 8980 -727 9314 -675
rect 9348 -667 9406 -573
rect 9348 -701 9360 -667
rect 9394 -701 9406 -667
rect 9348 -718 9406 -701
rect 9440 -634 10142 -573
rect 9440 -668 9458 -634
rect 9492 -668 10090 -634
rect 10124 -668 10142 -634
rect 9440 -727 10142 -668
rect 10176 -667 10234 -573
rect 10176 -701 10188 -667
rect 10222 -701 10234 -667
rect 10176 -718 10234 -701
rect 10360 -641 10694 -573
rect 10360 -675 10378 -641
rect 10412 -675 10642 -641
rect 10676 -675 10694 -641
rect 10360 -727 10694 -675
rect 8660 -761 8730 -737
rect 8236 -805 8239 -771
rect 8273 -805 8389 -771
rect 8236 -821 8389 -805
rect 8423 -771 8595 -770
rect 8423 -805 8439 -771
rect 8473 -805 8595 -771
rect 8423 -820 8595 -805
rect 8644 -771 8730 -761
rect 8644 -805 8660 -771
rect 8694 -805 8730 -771
rect 8644 -819 8730 -805
rect 8764 -775 8780 -771
rect 8764 -809 8774 -775
rect 8814 -805 8854 -771
rect 8808 -809 8854 -805
rect 8764 -814 8854 -809
rect 8980 -795 9000 -761
rect 9034 -795 9130 -761
rect 8355 -855 8389 -821
rect 8355 -889 8473 -855
rect 8152 -931 8233 -894
rect 8152 -965 8185 -931
rect 8219 -965 8233 -931
rect 8152 -999 8233 -965
rect 8152 -1033 8185 -999
rect 8219 -1033 8233 -999
rect 8152 -1049 8233 -1033
rect 8267 -932 8333 -923
rect 8267 -966 8283 -932
rect 8317 -966 8333 -932
rect 8267 -1000 8333 -966
rect 8267 -1034 8283 -1000
rect 8317 -1034 8333 -1000
rect 8267 -1083 8333 -1034
rect 8423 -931 8473 -889
rect 8423 -965 8439 -931
rect 8423 -999 8473 -965
rect 8423 -1033 8439 -999
rect 8423 -1049 8473 -1033
rect 8525 -932 8595 -820
rect 8660 -848 8730 -819
rect 8660 -882 8854 -848
rect 8525 -966 8543 -932
rect 8577 -966 8595 -932
rect 8525 -1000 8595 -966
rect 8525 -1034 8543 -1000
rect 8577 -1034 8595 -1000
rect 8525 -1049 8595 -1034
rect 8685 -932 8751 -916
rect 8685 -966 8701 -932
rect 8735 -966 8751 -932
rect 8685 -1000 8751 -966
rect 8685 -1034 8701 -1000
rect 8735 -1034 8751 -1000
rect 8685 -1083 8751 -1034
rect 8785 -932 8854 -882
rect 8785 -966 8801 -932
rect 8835 -966 8854 -932
rect 8785 -1000 8854 -966
rect 8785 -1034 8801 -1000
rect 8835 -1034 8854 -1000
rect 8785 -1049 8854 -1034
rect 8888 -885 8946 -850
rect 8888 -919 8900 -885
rect 8934 -919 8946 -885
rect 8888 -978 8946 -919
rect 8888 -1012 8900 -978
rect 8934 -1012 8946 -978
rect 8888 -1083 8946 -1012
rect 8980 -865 9130 -795
rect 9164 -797 9314 -727
rect 9164 -831 9260 -797
rect 9294 -831 9314 -797
rect 9440 -795 9518 -761
rect 9552 -795 9621 -761
rect 9655 -795 9724 -761
rect 9758 -795 9778 -761
rect 8980 -905 9314 -865
rect 8980 -939 8998 -905
rect 9032 -939 9262 -905
rect 9296 -939 9314 -905
rect 8980 -1007 9314 -939
rect 8980 -1041 8998 -1007
rect 9032 -1041 9262 -1007
rect 9296 -1041 9314 -1007
rect 8980 -1083 9314 -1041
rect 9348 -885 9406 -850
rect 9348 -919 9360 -885
rect 9394 -919 9406 -885
rect 9348 -978 9406 -919
rect 9348 -1012 9360 -978
rect 9394 -1012 9406 -978
rect 9348 -1083 9406 -1012
rect 9440 -865 9778 -795
rect 9812 -797 10142 -727
rect 9812 -831 9832 -797
rect 9866 -831 9931 -797
rect 9965 -831 10030 -797
rect 10064 -831 10142 -797
rect 10360 -795 10380 -761
rect 10414 -795 10510 -761
rect 9440 -905 10142 -865
rect 9440 -939 9458 -905
rect 9492 -939 10090 -905
rect 10124 -939 10142 -905
rect 9440 -1007 10142 -939
rect 9440 -1041 9458 -1007
rect 9492 -1041 10090 -1007
rect 10124 -1041 10142 -1007
rect 9440 -1083 10142 -1041
rect 10176 -885 10234 -850
rect 10176 -919 10188 -885
rect 10222 -919 10234 -885
rect 10176 -978 10234 -919
rect 10176 -1012 10188 -978
rect 10222 -1012 10234 -978
rect 10176 -1083 10234 -1012
rect 10360 -865 10510 -795
rect 10544 -797 10694 -727
rect 10544 -831 10640 -797
rect 10674 -831 10694 -797
rect 10728 -626 10809 -607
rect 10728 -660 10761 -626
rect 10795 -660 10809 -626
rect 10728 -684 10809 -660
rect 10843 -626 10909 -573
rect 10843 -660 10859 -626
rect 10893 -660 10909 -626
rect 10843 -676 10909 -660
rect 10999 -626 11049 -607
rect 10999 -660 11015 -626
rect 10728 -777 10778 -684
rect 10999 -702 11049 -660
rect 10931 -736 11049 -702
rect 11101 -626 11171 -607
rect 11101 -660 11120 -626
rect 11154 -660 11171 -626
rect 10931 -755 10965 -736
rect 10728 -811 10737 -777
rect 10771 -811 10778 -777
rect 10360 -905 10694 -865
rect 10360 -939 10378 -905
rect 10412 -939 10642 -905
rect 10676 -939 10694 -905
rect 10360 -1007 10694 -939
rect 10360 -1041 10378 -1007
rect 10412 -1041 10642 -1007
rect 10676 -1041 10694 -1007
rect 10360 -1083 10694 -1041
rect 10728 -894 10778 -811
rect 10812 -771 10965 -755
rect 11101 -770 11171 -660
rect 11264 -626 11330 -573
rect 11264 -660 11280 -626
rect 11314 -660 11330 -626
rect 11264 -669 11330 -660
rect 11364 -626 11430 -607
rect 11364 -660 11377 -626
rect 11411 -660 11430 -626
rect 11364 -703 11430 -660
rect 11236 -737 11430 -703
rect 11464 -667 11522 -573
rect 11464 -701 11476 -667
rect 11510 -701 11522 -667
rect 11464 -718 11522 -701
rect 11648 -641 11982 -573
rect 11648 -675 11666 -641
rect 11700 -675 11930 -641
rect 11964 -675 11982 -641
rect 11648 -727 11982 -675
rect 13580 -667 13638 -573
rect 13580 -701 13592 -667
rect 13626 -701 13638 -667
rect 13672 -615 13733 -573
rect 13672 -649 13690 -615
rect 13724 -649 13733 -615
rect 13672 -675 13733 -649
rect 13769 -628 13819 -609
rect 13769 -662 13776 -628
rect 13810 -662 13819 -628
rect 13580 -718 13638 -701
rect 11236 -761 11306 -737
rect 10812 -805 10815 -771
rect 10849 -805 10965 -771
rect 10812 -821 10965 -805
rect 10999 -771 11171 -770
rect 10999 -805 11015 -771
rect 11049 -805 11171 -771
rect 10999 -820 11171 -805
rect 11220 -771 11306 -761
rect 11220 -805 11236 -771
rect 11270 -805 11306 -771
rect 11220 -819 11306 -805
rect 11340 -805 11356 -771
rect 11390 -778 11430 -771
rect 11340 -812 11369 -805
rect 11403 -812 11430 -778
rect 11340 -814 11430 -812
rect 11648 -795 11668 -761
rect 11702 -795 11798 -761
rect 10931 -855 10965 -821
rect 10931 -889 11049 -855
rect 10728 -931 10809 -894
rect 10728 -965 10761 -931
rect 10795 -965 10809 -931
rect 10728 -999 10809 -965
rect 10728 -1033 10761 -999
rect 10795 -1033 10809 -999
rect 10728 -1049 10809 -1033
rect 10843 -932 10909 -923
rect 10843 -966 10859 -932
rect 10893 -966 10909 -932
rect 10843 -1000 10909 -966
rect 10843 -1034 10859 -1000
rect 10893 -1034 10909 -1000
rect 10843 -1083 10909 -1034
rect 10999 -931 11049 -889
rect 10999 -965 11015 -931
rect 10999 -999 11049 -965
rect 10999 -1033 11015 -999
rect 10999 -1049 11049 -1033
rect 11101 -932 11171 -820
rect 11236 -848 11306 -819
rect 11236 -882 11430 -848
rect 11101 -966 11119 -932
rect 11153 -966 11171 -932
rect 11101 -1000 11171 -966
rect 11101 -1034 11119 -1000
rect 11153 -1034 11171 -1000
rect 11101 -1049 11171 -1034
rect 11261 -932 11327 -916
rect 11261 -966 11277 -932
rect 11311 -966 11327 -932
rect 11261 -1000 11327 -966
rect 11261 -1034 11277 -1000
rect 11311 -1034 11327 -1000
rect 11261 -1083 11327 -1034
rect 11361 -932 11430 -882
rect 11361 -966 11377 -932
rect 11411 -966 11430 -932
rect 11361 -1000 11430 -966
rect 11361 -1034 11377 -1000
rect 11411 -1034 11430 -1000
rect 11361 -1049 11430 -1034
rect 11464 -885 11522 -850
rect 11464 -919 11476 -885
rect 11510 -919 11522 -885
rect 11464 -978 11522 -919
rect 11464 -1012 11476 -978
rect 11510 -1012 11522 -978
rect 11464 -1083 11522 -1012
rect 11648 -865 11798 -795
rect 11832 -797 11982 -727
rect 11832 -831 11928 -797
rect 11962 -831 11982 -797
rect 13672 -746 13735 -709
rect 13672 -780 13685 -746
rect 13719 -771 13735 -746
rect 13672 -805 13692 -780
rect 13726 -805 13735 -771
rect 13672 -821 13735 -805
rect 13769 -771 13819 -662
rect 13853 -628 13905 -573
rect 13853 -662 13862 -628
rect 13896 -662 13905 -628
rect 13853 -678 13905 -662
rect 13941 -628 13991 -609
rect 13941 -662 13948 -628
rect 13982 -662 13991 -628
rect 13941 -771 13991 -662
rect 14025 -628 14077 -573
rect 14025 -662 14034 -628
rect 14068 -662 14077 -628
rect 14025 -685 14077 -662
rect 14111 -628 14163 -612
rect 14111 -662 14120 -628
rect 14154 -662 14163 -628
rect 14111 -703 14163 -662
rect 14197 -619 14249 -573
rect 14197 -653 14206 -619
rect 14240 -653 14249 -619
rect 14197 -669 14249 -653
rect 14283 -628 14335 -612
rect 14283 -662 14292 -628
rect 14326 -662 14335 -628
rect 14283 -703 14335 -662
rect 14369 -619 14421 -573
rect 14369 -653 14378 -619
rect 14412 -653 14421 -619
rect 14369 -669 14421 -653
rect 14455 -628 14507 -612
rect 14455 -662 14464 -628
rect 14498 -662 14507 -628
rect 14455 -703 14507 -662
rect 14541 -619 14590 -573
rect 14541 -653 14550 -619
rect 14584 -653 14590 -619
rect 14541 -669 14590 -653
rect 14624 -628 14679 -612
rect 14624 -662 14636 -628
rect 14670 -662 14679 -628
rect 14624 -703 14679 -662
rect 14713 -619 14762 -573
rect 14713 -653 14722 -619
rect 14756 -653 14762 -619
rect 14713 -669 14762 -653
rect 14796 -628 14848 -612
rect 14796 -662 14807 -628
rect 14841 -662 14848 -628
rect 14796 -703 14848 -662
rect 14884 -619 14934 -573
rect 14884 -653 14893 -619
rect 14927 -653 14934 -619
rect 14884 -669 14934 -653
rect 14968 -628 15020 -612
rect 14968 -662 14979 -628
rect 15013 -662 15020 -628
rect 14968 -703 15020 -662
rect 15056 -619 15106 -573
rect 15056 -653 15065 -619
rect 15099 -653 15106 -619
rect 15056 -669 15106 -653
rect 15140 -628 15192 -612
rect 15140 -662 15151 -628
rect 15185 -662 15192 -628
rect 15140 -703 15192 -662
rect 15228 -619 15280 -573
rect 15228 -653 15237 -619
rect 15271 -653 15280 -619
rect 15228 -669 15280 -653
rect 15314 -628 15366 -612
rect 15314 -662 15323 -628
rect 15357 -662 15366 -628
rect 15314 -703 15366 -662
rect 15400 -619 15460 -573
rect 15400 -653 15409 -619
rect 15443 -653 15460 -619
rect 15400 -669 15460 -653
rect 15512 -667 15570 -573
rect 15512 -701 15524 -667
rect 15558 -701 15570 -667
rect 14111 -728 15460 -703
rect 15512 -718 15570 -701
rect 15605 -634 16674 -573
rect 15605 -668 15622 -634
rect 15656 -668 16622 -634
rect 16656 -668 16674 -634
rect 15605 -727 16674 -668
rect 14111 -737 15248 -728
rect 15227 -762 15248 -737
rect 15282 -729 15460 -728
rect 15282 -762 15340 -729
rect 15227 -763 15340 -762
rect 15374 -763 15460 -729
rect 13769 -805 14119 -771
rect 14153 -805 14187 -771
rect 14221 -805 14255 -771
rect 14289 -805 14323 -771
rect 14357 -805 14391 -771
rect 14425 -805 14459 -771
rect 14493 -805 14527 -771
rect 14561 -805 14595 -771
rect 14629 -805 14663 -771
rect 14697 -805 14731 -771
rect 14765 -805 14799 -771
rect 14833 -805 14867 -771
rect 14901 -805 14935 -771
rect 14969 -805 15003 -771
rect 15037 -805 15071 -771
rect 15105 -805 15139 -771
rect 15173 -805 15193 -771
rect 13769 -821 15193 -805
rect 11648 -905 11982 -865
rect 11648 -939 11666 -905
rect 11700 -939 11930 -905
rect 11964 -939 11982 -905
rect 11648 -1007 11982 -939
rect 11648 -1041 11666 -1007
rect 11700 -1041 11930 -1007
rect 11964 -1041 11982 -1007
rect 11648 -1083 11982 -1041
rect 13580 -885 13638 -850
rect 13580 -919 13592 -885
rect 13626 -919 13638 -885
rect 13580 -978 13638 -919
rect 13580 -1012 13592 -978
rect 13626 -1012 13638 -978
rect 13580 -1083 13638 -1012
rect 13674 -939 13733 -921
rect 13674 -973 13690 -939
rect 13724 -973 13733 -939
rect 13674 -1007 13733 -973
rect 13674 -1041 13690 -1007
rect 13724 -1041 13733 -1007
rect 13674 -1083 13733 -1041
rect 13769 -931 13818 -821
rect 13769 -965 13776 -931
rect 13810 -965 13818 -931
rect 13769 -999 13818 -965
rect 13769 -1033 13776 -999
rect 13810 -1033 13818 -999
rect 13769 -1049 13818 -1033
rect 13853 -939 13905 -921
rect 13853 -973 13862 -939
rect 13896 -973 13905 -939
rect 13853 -1007 13905 -973
rect 13853 -1041 13862 -1007
rect 13896 -1041 13905 -1007
rect 13853 -1083 13905 -1041
rect 13941 -923 13991 -821
rect 15227 -824 15460 -763
rect 15227 -855 15248 -824
rect 14111 -858 15248 -855
rect 15282 -858 15341 -824
rect 15375 -858 15460 -824
rect 15605 -795 15686 -761
rect 15720 -795 15814 -761
rect 15848 -795 15942 -761
rect 15976 -795 16070 -761
rect 16104 -795 16124 -761
rect 14111 -877 15460 -858
rect 14111 -911 14120 -877
rect 14154 -903 14292 -877
rect 14154 -911 14163 -903
rect 13941 -957 13948 -923
rect 13982 -957 13991 -923
rect 13941 -991 13991 -957
rect 13941 -1025 13948 -991
rect 13982 -1025 13991 -991
rect 13941 -1048 13991 -1025
rect 14025 -939 14077 -923
rect 14025 -973 14034 -939
rect 14068 -973 14077 -939
rect 14025 -1007 14077 -973
rect 14025 -1041 14034 -1007
rect 14068 -1041 14077 -1007
rect 14025 -1082 14077 -1041
rect 14111 -963 14163 -911
rect 14283 -911 14292 -903
rect 14326 -903 14464 -877
rect 14326 -911 14335 -903
rect 14111 -997 14120 -963
rect 14154 -997 14163 -963
rect 14111 -1048 14163 -997
rect 14197 -983 14249 -937
rect 14197 -1017 14206 -983
rect 14240 -1017 14249 -983
rect 14197 -1082 14249 -1017
rect 14283 -963 14335 -911
rect 14455 -911 14464 -903
rect 14498 -903 14636 -877
rect 14498 -911 14507 -903
rect 14283 -997 14292 -963
rect 14326 -997 14335 -963
rect 14283 -1048 14335 -997
rect 14369 -983 14421 -937
rect 14369 -1017 14378 -983
rect 14412 -1017 14421 -983
rect 14369 -1082 14421 -1017
rect 14455 -963 14507 -911
rect 14627 -911 14636 -903
rect 14670 -903 14807 -877
rect 14670 -911 14679 -903
rect 14455 -997 14464 -963
rect 14498 -997 14507 -963
rect 14455 -1048 14507 -997
rect 14541 -983 14593 -937
rect 14541 -1017 14550 -983
rect 14584 -1017 14593 -983
rect 14541 -1082 14593 -1017
rect 14627 -963 14679 -911
rect 14796 -911 14807 -903
rect 14841 -903 14979 -877
rect 14841 -911 14848 -903
rect 14627 -997 14636 -963
rect 14670 -997 14679 -963
rect 14627 -1048 14679 -997
rect 14713 -983 14762 -937
rect 14713 -1017 14722 -983
rect 14756 -1017 14762 -983
rect 14713 -1082 14762 -1017
rect 14796 -963 14848 -911
rect 14968 -911 14979 -903
rect 15013 -903 15151 -877
rect 15013 -911 15020 -903
rect 14796 -997 14807 -963
rect 14841 -997 14848 -963
rect 14796 -1048 14848 -997
rect 14885 -983 14934 -937
rect 14885 -1017 14893 -983
rect 14927 -1017 14934 -983
rect 14885 -1082 14934 -1017
rect 14968 -963 15020 -911
rect 15140 -911 15151 -903
rect 15185 -900 15323 -877
rect 15185 -911 15192 -900
rect 14968 -997 14979 -963
rect 15013 -997 15020 -963
rect 14968 -1048 15020 -997
rect 15057 -983 15106 -937
rect 15057 -1017 15065 -983
rect 15099 -1017 15106 -983
rect 15057 -1082 15106 -1017
rect 15140 -963 15192 -911
rect 15314 -911 15323 -900
rect 15357 -900 15460 -877
rect 15512 -885 15570 -850
rect 15357 -911 15372 -900
rect 15140 -997 15151 -963
rect 15185 -997 15192 -963
rect 15140 -1048 15192 -997
rect 15229 -983 15280 -937
rect 15229 -1017 15237 -983
rect 15271 -1017 15280 -983
rect 15229 -1082 15280 -1017
rect 15314 -963 15372 -911
rect 15512 -919 15524 -885
rect 15558 -919 15570 -885
rect 15314 -997 15323 -963
rect 15357 -997 15372 -963
rect 15314 -1048 15372 -997
rect 15406 -983 15460 -934
rect 15406 -1017 15409 -983
rect 15443 -1017 15460 -983
rect 14025 -1083 15280 -1082
rect 15406 -1083 15460 -1017
rect 15512 -978 15570 -919
rect 15512 -1012 15524 -978
rect 15558 -1012 15570 -978
rect 15512 -1083 15570 -1012
rect 15605 -865 16124 -795
rect 16158 -797 16674 -727
rect 16158 -831 16178 -797
rect 16212 -831 16306 -797
rect 16340 -831 16434 -797
rect 16468 -831 16562 -797
rect 16596 -831 16674 -797
rect 15605 -905 16674 -865
rect 15605 -939 15622 -905
rect 15656 -939 16622 -905
rect 16656 -939 16674 -905
rect 15605 -1007 16674 -939
rect 15605 -1041 15622 -1007
rect 15656 -1041 16622 -1007
rect 16656 -1041 16674 -1007
rect 15605 -1083 16674 -1041
rect -2997 -1117 -2968 -1083
rect -2934 -1117 -2876 -1083
rect -2842 -1117 -2784 -1083
rect -2750 -1117 -2692 -1083
rect -2658 -1117 -2600 -1083
rect -2566 -1117 -2508 -1083
rect -2474 -1117 -2416 -1083
rect -2382 -1117 -2324 -1083
rect -2290 -1117 -2232 -1083
rect -2198 -1117 -2140 -1083
rect -2106 -1117 -2048 -1083
rect -2014 -1117 -1956 -1083
rect -1922 -1117 -1864 -1083
rect -1830 -1117 -1772 -1083
rect -1738 -1117 -1680 -1083
rect -1646 -1117 -1588 -1083
rect -1554 -1117 -1496 -1083
rect -1462 -1117 -1404 -1083
rect -1370 -1117 -1312 -1083
rect -1278 -1117 -1220 -1083
rect -1186 -1117 -1128 -1083
rect -1094 -1117 -1036 -1083
rect -1002 -1117 -944 -1083
rect -910 -1117 -852 -1083
rect -818 -1117 -760 -1083
rect -726 -1117 -668 -1083
rect -634 -1117 -576 -1083
rect -542 -1117 -484 -1083
rect -450 -1117 -392 -1083
rect -358 -1117 -300 -1083
rect -266 -1117 -208 -1083
rect -174 -1117 -116 -1083
rect -82 -1117 -24 -1083
rect 10 -1117 68 -1083
rect 102 -1117 160 -1083
rect 194 -1117 252 -1083
rect 286 -1117 344 -1083
rect 378 -1117 436 -1083
rect 470 -1117 528 -1083
rect 562 -1117 620 -1083
rect 654 -1117 712 -1083
rect 746 -1117 804 -1083
rect 838 -1117 896 -1083
rect 930 -1117 988 -1083
rect 1022 -1117 1080 -1083
rect 1114 -1117 1172 -1083
rect 1206 -1117 1264 -1083
rect 1298 -1117 1356 -1083
rect 1390 -1117 1448 -1083
rect 1482 -1117 1540 -1083
rect 1574 -1117 1632 -1083
rect 1666 -1117 1724 -1083
rect 1758 -1117 1816 -1083
rect 1850 -1117 1908 -1083
rect 1942 -1117 2000 -1083
rect 2034 -1117 2092 -1083
rect 2126 -1117 2184 -1083
rect 2218 -1117 2276 -1083
rect 2310 -1117 2368 -1083
rect 2402 -1117 2460 -1083
rect 2494 -1117 2552 -1083
rect 2586 -1117 2644 -1083
rect 2678 -1117 2736 -1083
rect 2770 -1117 2828 -1083
rect 2862 -1117 2920 -1083
rect 2954 -1117 3012 -1083
rect 3046 -1117 3104 -1083
rect 3138 -1117 3196 -1083
rect 3230 -1117 3288 -1083
rect 3322 -1117 3380 -1083
rect 3414 -1117 3472 -1083
rect 3506 -1117 3564 -1083
rect 3598 -1117 3656 -1083
rect 3690 -1117 3748 -1083
rect 3782 -1117 3840 -1083
rect 3874 -1117 3932 -1083
rect 3966 -1117 4024 -1083
rect 4058 -1117 4116 -1083
rect 4150 -1117 4208 -1083
rect 4242 -1117 4300 -1083
rect 4334 -1117 4392 -1083
rect 4426 -1117 4484 -1083
rect 4518 -1117 4576 -1083
rect 4610 -1117 4668 -1083
rect 4702 -1117 4760 -1083
rect 4794 -1117 4852 -1083
rect 4886 -1117 4944 -1083
rect 4978 -1117 5036 -1083
rect 5070 -1117 5128 -1083
rect 5162 -1117 5220 -1083
rect 5254 -1117 5312 -1083
rect 5346 -1117 5404 -1083
rect 5438 -1117 5496 -1083
rect 5530 -1117 5588 -1083
rect 5622 -1117 5680 -1083
rect 5714 -1117 5772 -1083
rect 5806 -1117 5864 -1083
rect 5898 -1117 5956 -1083
rect 5990 -1117 6048 -1083
rect 6082 -1117 6140 -1083
rect 6174 -1117 6232 -1083
rect 6266 -1117 6324 -1083
rect 6358 -1117 6416 -1083
rect 6450 -1117 6508 -1083
rect 6542 -1117 6600 -1083
rect 6634 -1117 6692 -1083
rect 6726 -1117 6784 -1083
rect 6818 -1117 6876 -1083
rect 6910 -1117 6968 -1083
rect 7002 -1117 7060 -1083
rect 7094 -1117 7152 -1083
rect 7186 -1117 7244 -1083
rect 7278 -1117 7336 -1083
rect 7370 -1117 7428 -1083
rect 7462 -1117 7520 -1083
rect 7554 -1117 7612 -1083
rect 7646 -1117 7704 -1083
rect 7738 -1117 7796 -1083
rect 7830 -1117 7888 -1083
rect 7922 -1117 7980 -1083
rect 8014 -1117 8072 -1083
rect 8106 -1117 8164 -1083
rect 8198 -1117 8256 -1083
rect 8290 -1117 8348 -1083
rect 8382 -1117 8440 -1083
rect 8474 -1117 8532 -1083
rect 8566 -1117 8624 -1083
rect 8658 -1117 8716 -1083
rect 8750 -1117 8808 -1083
rect 8842 -1117 8900 -1083
rect 8934 -1117 8992 -1083
rect 9026 -1117 9084 -1083
rect 9118 -1117 9176 -1083
rect 9210 -1117 9268 -1083
rect 9302 -1117 9360 -1083
rect 9394 -1117 9452 -1083
rect 9486 -1117 9544 -1083
rect 9578 -1117 9636 -1083
rect 9670 -1117 9728 -1083
rect 9762 -1117 9820 -1083
rect 9854 -1117 9912 -1083
rect 9946 -1117 10004 -1083
rect 10038 -1117 10096 -1083
rect 10130 -1117 10188 -1083
rect 10222 -1117 10280 -1083
rect 10314 -1117 10372 -1083
rect 10406 -1117 10464 -1083
rect 10498 -1117 10556 -1083
rect 10590 -1117 10648 -1083
rect 10682 -1117 10740 -1083
rect 10774 -1117 10832 -1083
rect 10866 -1117 10924 -1083
rect 10958 -1117 11016 -1083
rect 11050 -1117 11108 -1083
rect 11142 -1117 11200 -1083
rect 11234 -1117 11292 -1083
rect 11326 -1117 11384 -1083
rect 11418 -1117 11476 -1083
rect 11510 -1117 11568 -1083
rect 11602 -1117 11660 -1083
rect 11694 -1117 11752 -1083
rect 11786 -1117 11844 -1083
rect 11878 -1117 11936 -1083
rect 11970 -1117 12028 -1083
rect 12062 -1117 12120 -1083
rect 12154 -1117 12212 -1083
rect 12246 -1117 12304 -1083
rect 12338 -1117 12396 -1083
rect 12430 -1117 12488 -1083
rect 12522 -1117 12580 -1083
rect 12614 -1117 12672 -1083
rect 12706 -1117 12764 -1083
rect 12798 -1117 12856 -1083
rect 12890 -1117 12948 -1083
rect 12982 -1117 13040 -1083
rect 13074 -1117 13132 -1083
rect 13166 -1117 13224 -1083
rect 13258 -1117 13316 -1083
rect 13350 -1117 13408 -1083
rect 13442 -1117 13500 -1083
rect 13534 -1117 13592 -1083
rect 13626 -1117 13684 -1083
rect 13718 -1117 13776 -1083
rect 13810 -1117 13868 -1083
rect 13902 -1117 13960 -1083
rect 13994 -1117 14052 -1083
rect 14086 -1117 14144 -1083
rect 14178 -1117 14236 -1083
rect 14270 -1117 14328 -1083
rect 14362 -1117 14420 -1083
rect 14454 -1117 14512 -1083
rect 14546 -1117 14604 -1083
rect 14638 -1117 14696 -1083
rect 14730 -1117 14788 -1083
rect 14822 -1117 14880 -1083
rect 14914 -1117 14972 -1083
rect 15006 -1117 15064 -1083
rect 15098 -1117 15156 -1083
rect 15190 -1117 15248 -1083
rect 15282 -1117 15340 -1083
rect 15374 -1117 15432 -1083
rect 15466 -1117 15524 -1083
rect 15558 -1117 15616 -1083
rect 15650 -1117 15708 -1083
rect 15742 -1117 15800 -1083
rect 15834 -1117 15892 -1083
rect 15926 -1117 15984 -1083
rect 16018 -1117 16076 -1083
rect 16110 -1117 16168 -1083
rect 16202 -1117 16260 -1083
rect 16294 -1117 16352 -1083
rect 16386 -1117 16444 -1083
rect 16478 -1117 16536 -1083
rect 16570 -1117 16628 -1083
rect 16662 -1117 16691 -1083
rect -2980 -1159 -2278 -1117
rect -2980 -1193 -2962 -1159
rect -2928 -1193 -2330 -1159
rect -2296 -1193 -2278 -1159
rect -2980 -1261 -2278 -1193
rect -2980 -1295 -2962 -1261
rect -2928 -1295 -2330 -1261
rect -2296 -1295 -2278 -1261
rect -2980 -1335 -2278 -1295
rect -2980 -1403 -2902 -1369
rect -2868 -1403 -2803 -1369
rect -2769 -1403 -2704 -1369
rect -2670 -1403 -2650 -1369
rect -2980 -1473 -2650 -1403
rect -2616 -1405 -2278 -1335
rect -2244 -1188 -2186 -1117
rect -2244 -1222 -2232 -1188
rect -2198 -1222 -2186 -1188
rect -2244 -1281 -2186 -1222
rect -2244 -1315 -2232 -1281
rect -2198 -1315 -2186 -1281
rect -2244 -1350 -2186 -1315
rect -1600 -1159 -898 -1117
rect -1600 -1193 -1582 -1159
rect -1548 -1193 -950 -1159
rect -916 -1193 -898 -1159
rect -1600 -1261 -898 -1193
rect -1600 -1295 -1582 -1261
rect -1548 -1295 -950 -1261
rect -916 -1295 -898 -1261
rect -1600 -1335 -898 -1295
rect -864 -1159 -162 -1117
rect -864 -1193 -846 -1159
rect -812 -1193 -214 -1159
rect -180 -1193 -162 -1159
rect -864 -1261 -162 -1193
rect -864 -1295 -846 -1261
rect -812 -1295 -214 -1261
rect -180 -1295 -162 -1261
rect -864 -1335 -162 -1295
rect -2616 -1439 -2596 -1405
rect -2562 -1439 -2493 -1405
rect -2459 -1439 -2390 -1405
rect -2356 -1439 -2278 -1405
rect -1600 -1403 -1522 -1369
rect -1488 -1403 -1423 -1369
rect -1389 -1403 -1324 -1369
rect -1290 -1403 -1270 -1369
rect -1600 -1473 -1270 -1403
rect -1236 -1405 -898 -1335
rect -1236 -1439 -1216 -1405
rect -1182 -1439 -1113 -1405
rect -1079 -1439 -1010 -1405
rect -976 -1439 -898 -1405
rect -864 -1403 -786 -1369
rect -752 -1403 -687 -1369
rect -653 -1403 -588 -1369
rect -554 -1403 -534 -1369
rect -864 -1473 -534 -1403
rect -500 -1405 -162 -1335
rect -128 -1188 -70 -1117
rect -128 -1222 -116 -1188
rect -82 -1222 -70 -1188
rect -128 -1281 -70 -1222
rect -128 -1315 -116 -1281
rect -82 -1315 -70 -1281
rect -128 -1350 -70 -1315
rect -36 -1159 298 -1117
rect -36 -1193 -18 -1159
rect 16 -1193 246 -1159
rect 280 -1193 298 -1159
rect -36 -1261 298 -1193
rect -36 -1295 -18 -1261
rect 16 -1295 246 -1261
rect 280 -1295 298 -1261
rect -36 -1335 298 -1295
rect 332 -1188 390 -1117
rect 332 -1222 344 -1188
rect 378 -1222 390 -1188
rect 332 -1281 390 -1222
rect 332 -1315 344 -1281
rect 378 -1315 390 -1281
rect -500 -1439 -480 -1405
rect -446 -1439 -377 -1405
rect -343 -1439 -274 -1405
rect -240 -1439 -162 -1405
rect -36 -1405 114 -1335
rect 332 -1350 390 -1315
rect 424 -1166 493 -1151
rect 424 -1200 443 -1166
rect 477 -1200 493 -1166
rect 424 -1234 493 -1200
rect 424 -1268 443 -1234
rect 477 -1268 493 -1234
rect 424 -1318 493 -1268
rect 527 -1166 593 -1117
rect 527 -1200 543 -1166
rect 577 -1200 593 -1166
rect 527 -1234 593 -1200
rect 527 -1268 543 -1234
rect 577 -1268 593 -1234
rect 527 -1284 593 -1268
rect 683 -1166 753 -1151
rect 683 -1200 701 -1166
rect 735 -1200 753 -1166
rect 683 -1234 753 -1200
rect 683 -1268 701 -1234
rect 735 -1268 753 -1234
rect 424 -1352 618 -1318
rect -36 -1439 -16 -1405
rect 18 -1439 114 -1405
rect 148 -1403 244 -1369
rect 278 -1403 298 -1369
rect 548 -1381 618 -1352
rect 683 -1380 753 -1268
rect 805 -1167 855 -1151
rect 839 -1201 855 -1167
rect 805 -1235 855 -1201
rect 839 -1269 855 -1235
rect 805 -1311 855 -1269
rect 945 -1166 1011 -1117
rect 945 -1200 961 -1166
rect 995 -1200 1011 -1166
rect 945 -1234 1011 -1200
rect 945 -1268 961 -1234
rect 995 -1268 1011 -1234
rect 945 -1277 1011 -1268
rect 1045 -1167 1126 -1151
rect 1045 -1201 1059 -1167
rect 1093 -1201 1126 -1167
rect 1045 -1235 1126 -1201
rect 1045 -1269 1059 -1235
rect 1093 -1269 1126 -1235
rect 1045 -1306 1126 -1269
rect 805 -1345 923 -1311
rect 889 -1379 923 -1345
rect 148 -1473 298 -1403
rect 424 -1392 514 -1386
rect 424 -1426 432 -1392
rect 466 -1395 514 -1392
rect 424 -1429 464 -1426
rect 498 -1429 514 -1395
rect 548 -1395 634 -1381
rect 548 -1429 584 -1395
rect 618 -1429 634 -1395
rect 548 -1439 634 -1429
rect 683 -1395 855 -1380
rect 683 -1429 805 -1395
rect 839 -1429 855 -1395
rect 683 -1430 855 -1429
rect 889 -1395 1042 -1379
rect 889 -1429 1005 -1395
rect 1039 -1429 1042 -1395
rect 548 -1463 618 -1439
rect -2980 -1532 -2278 -1473
rect -2980 -1566 -2962 -1532
rect -2928 -1566 -2330 -1532
rect -2296 -1566 -2278 -1532
rect -2980 -1627 -2278 -1566
rect -2244 -1499 -2186 -1482
rect -2244 -1533 -2232 -1499
rect -2198 -1533 -2186 -1499
rect -2244 -1627 -2186 -1533
rect -1600 -1532 -898 -1473
rect -1600 -1566 -1582 -1532
rect -1548 -1566 -950 -1532
rect -916 -1566 -898 -1532
rect -1600 -1627 -898 -1566
rect -864 -1532 -162 -1473
rect -864 -1566 -846 -1532
rect -812 -1566 -214 -1532
rect -180 -1566 -162 -1532
rect -864 -1627 -162 -1566
rect -128 -1499 -70 -1482
rect -128 -1533 -116 -1499
rect -82 -1533 -70 -1499
rect -128 -1627 -70 -1533
rect -36 -1525 298 -1473
rect -36 -1559 -18 -1525
rect 16 -1559 246 -1525
rect 280 -1559 298 -1525
rect -36 -1627 298 -1559
rect 332 -1499 390 -1482
rect 332 -1533 344 -1499
rect 378 -1533 390 -1499
rect 332 -1627 390 -1533
rect 424 -1497 618 -1463
rect 424 -1540 490 -1497
rect 424 -1574 443 -1540
rect 477 -1574 490 -1540
rect 424 -1593 490 -1574
rect 524 -1540 590 -1531
rect 524 -1574 540 -1540
rect 574 -1574 590 -1540
rect 524 -1627 590 -1574
rect 683 -1540 753 -1430
rect 889 -1445 1042 -1429
rect 1076 -1389 1126 -1306
rect 1160 -1188 1218 -1117
rect 1160 -1222 1172 -1188
rect 1206 -1222 1218 -1188
rect 1160 -1281 1218 -1222
rect 1160 -1315 1172 -1281
rect 1206 -1315 1218 -1281
rect 1160 -1350 1218 -1315
rect 1252 -1159 1586 -1117
rect 1252 -1193 1270 -1159
rect 1304 -1193 1534 -1159
rect 1568 -1193 1586 -1159
rect 1252 -1261 1586 -1193
rect 1252 -1295 1270 -1261
rect 1304 -1295 1534 -1261
rect 1568 -1295 1586 -1261
rect 1252 -1335 1586 -1295
rect 1620 -1188 1678 -1117
rect 1620 -1222 1632 -1188
rect 1666 -1222 1678 -1188
rect 1620 -1281 1678 -1222
rect 1620 -1315 1632 -1281
rect 1666 -1315 1678 -1281
rect 1076 -1423 1082 -1389
rect 1116 -1423 1126 -1389
rect 889 -1464 923 -1445
rect 683 -1574 700 -1540
rect 734 -1574 753 -1540
rect 683 -1593 753 -1574
rect 805 -1498 923 -1464
rect 805 -1540 855 -1498
rect 1076 -1516 1126 -1423
rect 1252 -1405 1402 -1335
rect 1620 -1350 1678 -1315
rect 1712 -1159 2414 -1117
rect 1712 -1193 1730 -1159
rect 1764 -1193 2362 -1159
rect 2396 -1193 2414 -1159
rect 1712 -1261 2414 -1193
rect 1712 -1295 1730 -1261
rect 1764 -1295 2362 -1261
rect 2396 -1295 2414 -1261
rect 1712 -1335 2414 -1295
rect 1252 -1439 1272 -1405
rect 1306 -1439 1402 -1405
rect 1436 -1403 1532 -1369
rect 1566 -1403 1586 -1369
rect 1436 -1473 1586 -1403
rect 839 -1574 855 -1540
rect 805 -1593 855 -1574
rect 945 -1540 1011 -1524
rect 945 -1574 961 -1540
rect 995 -1574 1011 -1540
rect 945 -1627 1011 -1574
rect 1045 -1540 1126 -1516
rect 1045 -1574 1059 -1540
rect 1093 -1574 1126 -1540
rect 1045 -1593 1126 -1574
rect 1160 -1499 1218 -1482
rect 1160 -1533 1172 -1499
rect 1206 -1533 1218 -1499
rect 1160 -1627 1218 -1533
rect 1252 -1525 1586 -1473
rect 1712 -1403 1790 -1369
rect 1824 -1403 1889 -1369
rect 1923 -1403 1988 -1369
rect 2022 -1403 2042 -1369
rect 1712 -1473 2042 -1403
rect 2076 -1405 2414 -1335
rect 2448 -1188 2506 -1117
rect 2448 -1222 2460 -1188
rect 2494 -1222 2506 -1188
rect 2448 -1281 2506 -1222
rect 2448 -1315 2460 -1281
rect 2494 -1315 2506 -1281
rect 2448 -1350 2506 -1315
rect 2540 -1159 2874 -1117
rect 2540 -1193 2558 -1159
rect 2592 -1193 2822 -1159
rect 2856 -1193 2874 -1159
rect 2540 -1261 2874 -1193
rect 2540 -1295 2558 -1261
rect 2592 -1295 2822 -1261
rect 2856 -1295 2874 -1261
rect 2540 -1335 2874 -1295
rect 2908 -1188 2966 -1117
rect 2908 -1222 2920 -1188
rect 2954 -1222 2966 -1188
rect 2908 -1281 2966 -1222
rect 2908 -1315 2920 -1281
rect 2954 -1315 2966 -1281
rect 2076 -1439 2096 -1405
rect 2130 -1439 2199 -1405
rect 2233 -1439 2302 -1405
rect 2336 -1439 2414 -1405
rect 2540 -1405 2690 -1335
rect 2908 -1350 2966 -1315
rect 3000 -1166 3069 -1151
rect 3000 -1200 3019 -1166
rect 3053 -1200 3069 -1166
rect 3000 -1234 3069 -1200
rect 3000 -1268 3019 -1234
rect 3053 -1268 3069 -1234
rect 3000 -1318 3069 -1268
rect 3103 -1166 3169 -1117
rect 3103 -1200 3119 -1166
rect 3153 -1200 3169 -1166
rect 3103 -1234 3169 -1200
rect 3103 -1268 3119 -1234
rect 3153 -1268 3169 -1234
rect 3103 -1284 3169 -1268
rect 3259 -1166 3329 -1151
rect 3259 -1200 3277 -1166
rect 3311 -1200 3329 -1166
rect 3259 -1234 3329 -1200
rect 3259 -1268 3277 -1234
rect 3311 -1268 3329 -1234
rect 3000 -1352 3194 -1318
rect 2540 -1439 2560 -1405
rect 2594 -1439 2690 -1405
rect 2724 -1403 2820 -1369
rect 2854 -1403 2874 -1369
rect 3124 -1381 3194 -1352
rect 3259 -1380 3329 -1268
rect 3381 -1167 3431 -1151
rect 3415 -1201 3431 -1167
rect 3381 -1235 3431 -1201
rect 3415 -1269 3431 -1235
rect 3381 -1311 3431 -1269
rect 3521 -1166 3587 -1117
rect 3521 -1200 3537 -1166
rect 3571 -1200 3587 -1166
rect 3521 -1234 3587 -1200
rect 3521 -1268 3537 -1234
rect 3571 -1268 3587 -1234
rect 3521 -1277 3587 -1268
rect 3621 -1167 3702 -1151
rect 3621 -1201 3635 -1167
rect 3669 -1201 3702 -1167
rect 3621 -1235 3702 -1201
rect 3621 -1269 3635 -1235
rect 3669 -1269 3702 -1235
rect 3621 -1306 3702 -1269
rect 3381 -1345 3499 -1311
rect 3465 -1379 3499 -1345
rect 2724 -1473 2874 -1403
rect 3000 -1389 3090 -1386
rect 3000 -1395 3042 -1389
rect 3000 -1429 3040 -1395
rect 3076 -1423 3090 -1389
rect 3074 -1429 3090 -1423
rect 3124 -1395 3210 -1381
rect 3124 -1429 3160 -1395
rect 3194 -1429 3210 -1395
rect 3124 -1439 3210 -1429
rect 3259 -1395 3431 -1380
rect 3259 -1429 3381 -1395
rect 3415 -1429 3431 -1395
rect 3259 -1430 3431 -1429
rect 3465 -1395 3618 -1379
rect 3465 -1429 3581 -1395
rect 3615 -1429 3618 -1395
rect 3124 -1463 3194 -1439
rect 1252 -1559 1270 -1525
rect 1304 -1559 1534 -1525
rect 1568 -1559 1586 -1525
rect 1252 -1627 1586 -1559
rect 1620 -1499 1678 -1482
rect 1620 -1533 1632 -1499
rect 1666 -1533 1678 -1499
rect 1620 -1627 1678 -1533
rect 1712 -1532 2414 -1473
rect 1712 -1566 1730 -1532
rect 1764 -1566 2362 -1532
rect 2396 -1566 2414 -1532
rect 1712 -1627 2414 -1566
rect 2448 -1499 2506 -1482
rect 2448 -1533 2460 -1499
rect 2494 -1533 2506 -1499
rect 2448 -1627 2506 -1533
rect 2540 -1525 2874 -1473
rect 2540 -1559 2558 -1525
rect 2592 -1559 2822 -1525
rect 2856 -1559 2874 -1525
rect 2540 -1627 2874 -1559
rect 2908 -1499 2966 -1482
rect 2908 -1533 2920 -1499
rect 2954 -1533 2966 -1499
rect 2908 -1627 2966 -1533
rect 3000 -1497 3194 -1463
rect 3000 -1540 3066 -1497
rect 3000 -1574 3019 -1540
rect 3053 -1574 3066 -1540
rect 3000 -1593 3066 -1574
rect 3100 -1540 3166 -1531
rect 3100 -1574 3116 -1540
rect 3150 -1574 3166 -1540
rect 3100 -1627 3166 -1574
rect 3259 -1540 3329 -1430
rect 3465 -1445 3618 -1429
rect 3652 -1389 3702 -1306
rect 3736 -1188 3794 -1117
rect 3736 -1222 3748 -1188
rect 3782 -1222 3794 -1188
rect 3736 -1281 3794 -1222
rect 3736 -1315 3748 -1281
rect 3782 -1315 3794 -1281
rect 3736 -1350 3794 -1315
rect 3828 -1159 4162 -1117
rect 3828 -1193 3846 -1159
rect 3880 -1193 4110 -1159
rect 4144 -1193 4162 -1159
rect 3828 -1261 4162 -1193
rect 3828 -1295 3846 -1261
rect 3880 -1295 4110 -1261
rect 4144 -1295 4162 -1261
rect 3828 -1335 4162 -1295
rect 4196 -1188 4254 -1117
rect 4196 -1222 4208 -1188
rect 4242 -1222 4254 -1188
rect 4196 -1281 4254 -1222
rect 4196 -1315 4208 -1281
rect 4242 -1315 4254 -1281
rect 3652 -1423 3656 -1389
rect 3690 -1423 3702 -1389
rect 3465 -1464 3499 -1445
rect 3259 -1574 3276 -1540
rect 3310 -1574 3329 -1540
rect 3259 -1593 3329 -1574
rect 3381 -1498 3499 -1464
rect 3381 -1540 3431 -1498
rect 3652 -1516 3702 -1423
rect 3828 -1405 3978 -1335
rect 4196 -1350 4254 -1315
rect 4288 -1159 4990 -1117
rect 4288 -1193 4306 -1159
rect 4340 -1193 4938 -1159
rect 4972 -1193 4990 -1159
rect 4288 -1261 4990 -1193
rect 4288 -1295 4306 -1261
rect 4340 -1295 4938 -1261
rect 4972 -1295 4990 -1261
rect 4288 -1335 4990 -1295
rect 3828 -1439 3848 -1405
rect 3882 -1439 3978 -1405
rect 4012 -1403 4108 -1369
rect 4142 -1403 4162 -1369
rect 4012 -1473 4162 -1403
rect 3415 -1574 3431 -1540
rect 3381 -1593 3431 -1574
rect 3521 -1540 3587 -1524
rect 3521 -1574 3537 -1540
rect 3571 -1574 3587 -1540
rect 3521 -1627 3587 -1574
rect 3621 -1540 3702 -1516
rect 3621 -1574 3635 -1540
rect 3669 -1574 3702 -1540
rect 3621 -1593 3702 -1574
rect 3736 -1499 3794 -1482
rect 3736 -1533 3748 -1499
rect 3782 -1533 3794 -1499
rect 3736 -1627 3794 -1533
rect 3828 -1525 4162 -1473
rect 4288 -1403 4366 -1369
rect 4400 -1403 4465 -1369
rect 4499 -1403 4564 -1369
rect 4598 -1403 4618 -1369
rect 4288 -1473 4618 -1403
rect 4652 -1405 4990 -1335
rect 5024 -1188 5082 -1117
rect 5024 -1222 5036 -1188
rect 5070 -1222 5082 -1188
rect 5024 -1281 5082 -1222
rect 5024 -1315 5036 -1281
rect 5070 -1315 5082 -1281
rect 5024 -1350 5082 -1315
rect 5116 -1159 5450 -1117
rect 5116 -1193 5134 -1159
rect 5168 -1193 5398 -1159
rect 5432 -1193 5450 -1159
rect 5116 -1261 5450 -1193
rect 5116 -1295 5134 -1261
rect 5168 -1295 5398 -1261
rect 5432 -1295 5450 -1261
rect 5116 -1335 5450 -1295
rect 5484 -1188 5542 -1117
rect 5484 -1222 5496 -1188
rect 5530 -1222 5542 -1188
rect 5484 -1281 5542 -1222
rect 5484 -1315 5496 -1281
rect 5530 -1315 5542 -1281
rect 4652 -1439 4672 -1405
rect 4706 -1439 4775 -1405
rect 4809 -1439 4878 -1405
rect 4912 -1439 4990 -1405
rect 5116 -1405 5266 -1335
rect 5484 -1350 5542 -1315
rect 5576 -1166 5645 -1151
rect 5576 -1200 5595 -1166
rect 5629 -1200 5645 -1166
rect 5576 -1234 5645 -1200
rect 5576 -1268 5595 -1234
rect 5629 -1268 5645 -1234
rect 5576 -1318 5645 -1268
rect 5679 -1166 5745 -1117
rect 5679 -1200 5695 -1166
rect 5729 -1200 5745 -1166
rect 5679 -1234 5745 -1200
rect 5679 -1268 5695 -1234
rect 5729 -1268 5745 -1234
rect 5679 -1284 5745 -1268
rect 5835 -1166 5905 -1151
rect 5835 -1200 5853 -1166
rect 5887 -1200 5905 -1166
rect 5835 -1234 5905 -1200
rect 5835 -1268 5853 -1234
rect 5887 -1268 5905 -1234
rect 5576 -1352 5770 -1318
rect 5116 -1439 5136 -1405
rect 5170 -1439 5266 -1405
rect 5300 -1403 5396 -1369
rect 5430 -1403 5450 -1369
rect 5700 -1381 5770 -1352
rect 5835 -1380 5905 -1268
rect 5957 -1167 6007 -1151
rect 5991 -1201 6007 -1167
rect 5957 -1235 6007 -1201
rect 5991 -1269 6007 -1235
rect 5957 -1311 6007 -1269
rect 6097 -1166 6163 -1117
rect 6097 -1200 6113 -1166
rect 6147 -1200 6163 -1166
rect 6097 -1234 6163 -1200
rect 6097 -1268 6113 -1234
rect 6147 -1268 6163 -1234
rect 6097 -1277 6163 -1268
rect 6197 -1167 6278 -1151
rect 6197 -1201 6211 -1167
rect 6245 -1201 6278 -1167
rect 6197 -1235 6278 -1201
rect 6197 -1269 6211 -1235
rect 6245 -1269 6278 -1235
rect 6197 -1306 6278 -1269
rect 5957 -1345 6075 -1311
rect 6041 -1379 6075 -1345
rect 5300 -1473 5450 -1403
rect 5576 -1389 5666 -1386
rect 5576 -1429 5616 -1389
rect 5650 -1429 5666 -1389
rect 5700 -1395 5786 -1381
rect 5700 -1429 5736 -1395
rect 5770 -1429 5786 -1395
rect 5700 -1439 5786 -1429
rect 5835 -1395 6007 -1380
rect 5835 -1429 5957 -1395
rect 5991 -1429 6007 -1395
rect 5835 -1430 6007 -1429
rect 6041 -1395 6194 -1379
rect 6041 -1429 6157 -1395
rect 6191 -1429 6194 -1395
rect 5700 -1463 5770 -1439
rect 3828 -1559 3846 -1525
rect 3880 -1559 4110 -1525
rect 4144 -1559 4162 -1525
rect 3828 -1627 4162 -1559
rect 4196 -1499 4254 -1482
rect 4196 -1533 4208 -1499
rect 4242 -1533 4254 -1499
rect 4196 -1627 4254 -1533
rect 4288 -1532 4990 -1473
rect 4288 -1566 4306 -1532
rect 4340 -1566 4938 -1532
rect 4972 -1566 4990 -1532
rect 4288 -1627 4990 -1566
rect 5024 -1499 5082 -1482
rect 5024 -1533 5036 -1499
rect 5070 -1533 5082 -1499
rect 5024 -1627 5082 -1533
rect 5116 -1525 5450 -1473
rect 5116 -1559 5134 -1525
rect 5168 -1559 5398 -1525
rect 5432 -1559 5450 -1525
rect 5116 -1627 5450 -1559
rect 5484 -1499 5542 -1482
rect 5484 -1533 5496 -1499
rect 5530 -1533 5542 -1499
rect 5484 -1627 5542 -1533
rect 5576 -1497 5770 -1463
rect 5576 -1540 5642 -1497
rect 5576 -1574 5595 -1540
rect 5629 -1574 5642 -1540
rect 5576 -1593 5642 -1574
rect 5676 -1540 5742 -1531
rect 5676 -1574 5692 -1540
rect 5726 -1574 5742 -1540
rect 5676 -1627 5742 -1574
rect 5835 -1540 5905 -1430
rect 6041 -1445 6194 -1429
rect 6228 -1389 6278 -1306
rect 6312 -1188 6370 -1117
rect 6312 -1222 6324 -1188
rect 6358 -1222 6370 -1188
rect 6312 -1281 6370 -1222
rect 6312 -1315 6324 -1281
rect 6358 -1315 6370 -1281
rect 6312 -1350 6370 -1315
rect 6404 -1159 6738 -1117
rect 6404 -1193 6422 -1159
rect 6456 -1193 6686 -1159
rect 6720 -1193 6738 -1159
rect 6404 -1261 6738 -1193
rect 6404 -1295 6422 -1261
rect 6456 -1295 6686 -1261
rect 6720 -1295 6738 -1261
rect 6404 -1335 6738 -1295
rect 6772 -1188 6830 -1117
rect 6772 -1222 6784 -1188
rect 6818 -1222 6830 -1188
rect 6772 -1281 6830 -1222
rect 6772 -1315 6784 -1281
rect 6818 -1315 6830 -1281
rect 6228 -1423 6230 -1389
rect 6264 -1423 6278 -1389
rect 6041 -1464 6075 -1445
rect 5835 -1574 5852 -1540
rect 5886 -1574 5905 -1540
rect 5835 -1593 5905 -1574
rect 5957 -1498 6075 -1464
rect 5957 -1540 6007 -1498
rect 6228 -1516 6278 -1423
rect 6404 -1405 6554 -1335
rect 6772 -1350 6830 -1315
rect 6864 -1159 7566 -1117
rect 6864 -1193 6882 -1159
rect 6916 -1193 7514 -1159
rect 7548 -1193 7566 -1159
rect 6864 -1261 7566 -1193
rect 6864 -1295 6882 -1261
rect 6916 -1295 7514 -1261
rect 7548 -1295 7566 -1261
rect 6864 -1335 7566 -1295
rect 6404 -1439 6424 -1405
rect 6458 -1439 6554 -1405
rect 6588 -1403 6684 -1369
rect 6718 -1403 6738 -1369
rect 6588 -1473 6738 -1403
rect 5991 -1574 6007 -1540
rect 5957 -1593 6007 -1574
rect 6097 -1540 6163 -1524
rect 6097 -1574 6113 -1540
rect 6147 -1574 6163 -1540
rect 6097 -1627 6163 -1574
rect 6197 -1540 6278 -1516
rect 6197 -1574 6211 -1540
rect 6245 -1574 6278 -1540
rect 6197 -1593 6278 -1574
rect 6312 -1499 6370 -1482
rect 6312 -1533 6324 -1499
rect 6358 -1533 6370 -1499
rect 6312 -1627 6370 -1533
rect 6404 -1525 6738 -1473
rect 6864 -1403 6942 -1369
rect 6976 -1403 7041 -1369
rect 7075 -1403 7140 -1369
rect 7174 -1403 7194 -1369
rect 6864 -1473 7194 -1403
rect 7228 -1405 7566 -1335
rect 7600 -1188 7658 -1117
rect 7600 -1222 7612 -1188
rect 7646 -1222 7658 -1188
rect 7600 -1281 7658 -1222
rect 7600 -1315 7612 -1281
rect 7646 -1315 7658 -1281
rect 7600 -1350 7658 -1315
rect 7692 -1159 8026 -1117
rect 7692 -1193 7710 -1159
rect 7744 -1193 7974 -1159
rect 8008 -1193 8026 -1159
rect 7692 -1261 8026 -1193
rect 7692 -1295 7710 -1261
rect 7744 -1295 7974 -1261
rect 8008 -1295 8026 -1261
rect 7692 -1335 8026 -1295
rect 8060 -1188 8118 -1117
rect 8060 -1222 8072 -1188
rect 8106 -1222 8118 -1188
rect 8060 -1281 8118 -1222
rect 8060 -1315 8072 -1281
rect 8106 -1315 8118 -1281
rect 7228 -1439 7248 -1405
rect 7282 -1439 7351 -1405
rect 7385 -1439 7454 -1405
rect 7488 -1439 7566 -1405
rect 7692 -1405 7842 -1335
rect 8060 -1350 8118 -1315
rect 8152 -1166 8221 -1151
rect 8152 -1200 8171 -1166
rect 8205 -1200 8221 -1166
rect 8152 -1234 8221 -1200
rect 8152 -1268 8171 -1234
rect 8205 -1268 8221 -1234
rect 8152 -1318 8221 -1268
rect 8255 -1166 8321 -1117
rect 8255 -1200 8271 -1166
rect 8305 -1200 8321 -1166
rect 8255 -1234 8321 -1200
rect 8255 -1268 8271 -1234
rect 8305 -1268 8321 -1234
rect 8255 -1284 8321 -1268
rect 8411 -1166 8481 -1151
rect 8411 -1200 8429 -1166
rect 8463 -1200 8481 -1166
rect 8411 -1234 8481 -1200
rect 8411 -1268 8429 -1234
rect 8463 -1268 8481 -1234
rect 8152 -1352 8346 -1318
rect 7692 -1439 7712 -1405
rect 7746 -1439 7842 -1405
rect 7876 -1403 7972 -1369
rect 8006 -1403 8026 -1369
rect 8276 -1381 8346 -1352
rect 8411 -1380 8481 -1268
rect 8533 -1167 8583 -1151
rect 8567 -1201 8583 -1167
rect 8533 -1235 8583 -1201
rect 8567 -1269 8583 -1235
rect 8533 -1311 8583 -1269
rect 8673 -1166 8739 -1117
rect 8673 -1200 8689 -1166
rect 8723 -1200 8739 -1166
rect 8673 -1234 8739 -1200
rect 8673 -1268 8689 -1234
rect 8723 -1268 8739 -1234
rect 8673 -1277 8739 -1268
rect 8773 -1167 8854 -1151
rect 8773 -1201 8787 -1167
rect 8821 -1201 8854 -1167
rect 8773 -1235 8854 -1201
rect 8773 -1269 8787 -1235
rect 8821 -1269 8854 -1235
rect 8773 -1306 8854 -1269
rect 8533 -1345 8651 -1311
rect 8617 -1379 8651 -1345
rect 7876 -1473 8026 -1403
rect 8152 -1389 8242 -1386
rect 8152 -1423 8190 -1389
rect 8224 -1395 8242 -1389
rect 8152 -1429 8192 -1423
rect 8226 -1429 8242 -1395
rect 8276 -1395 8362 -1381
rect 8276 -1429 8312 -1395
rect 8346 -1429 8362 -1395
rect 8276 -1439 8362 -1429
rect 8411 -1395 8583 -1380
rect 8411 -1429 8533 -1395
rect 8567 -1429 8583 -1395
rect 8411 -1430 8583 -1429
rect 8617 -1395 8770 -1379
rect 8617 -1429 8733 -1395
rect 8767 -1429 8770 -1395
rect 8276 -1463 8346 -1439
rect 6404 -1559 6422 -1525
rect 6456 -1559 6686 -1525
rect 6720 -1559 6738 -1525
rect 6404 -1627 6738 -1559
rect 6772 -1499 6830 -1482
rect 6772 -1533 6784 -1499
rect 6818 -1533 6830 -1499
rect 6772 -1627 6830 -1533
rect 6864 -1532 7566 -1473
rect 6864 -1566 6882 -1532
rect 6916 -1566 7514 -1532
rect 7548 -1566 7566 -1532
rect 6864 -1627 7566 -1566
rect 7600 -1499 7658 -1482
rect 7600 -1533 7612 -1499
rect 7646 -1533 7658 -1499
rect 7600 -1627 7658 -1533
rect 7692 -1525 8026 -1473
rect 7692 -1559 7710 -1525
rect 7744 -1559 7974 -1525
rect 8008 -1559 8026 -1525
rect 7692 -1627 8026 -1559
rect 8060 -1499 8118 -1482
rect 8060 -1533 8072 -1499
rect 8106 -1533 8118 -1499
rect 8060 -1627 8118 -1533
rect 8152 -1497 8346 -1463
rect 8152 -1540 8218 -1497
rect 8152 -1574 8171 -1540
rect 8205 -1574 8218 -1540
rect 8152 -1593 8218 -1574
rect 8252 -1540 8318 -1531
rect 8252 -1574 8268 -1540
rect 8302 -1574 8318 -1540
rect 8252 -1627 8318 -1574
rect 8411 -1540 8481 -1430
rect 8617 -1445 8770 -1429
rect 8804 -1389 8854 -1306
rect 8888 -1188 8946 -1117
rect 8888 -1222 8900 -1188
rect 8934 -1222 8946 -1188
rect 8888 -1281 8946 -1222
rect 8888 -1315 8900 -1281
rect 8934 -1315 8946 -1281
rect 8888 -1350 8946 -1315
rect 8980 -1159 9314 -1117
rect 8980 -1193 8998 -1159
rect 9032 -1193 9262 -1159
rect 9296 -1193 9314 -1159
rect 8980 -1261 9314 -1193
rect 8980 -1295 8998 -1261
rect 9032 -1295 9262 -1261
rect 9296 -1295 9314 -1261
rect 8980 -1335 9314 -1295
rect 9348 -1188 9406 -1117
rect 9348 -1222 9360 -1188
rect 9394 -1222 9406 -1188
rect 9348 -1281 9406 -1222
rect 9348 -1315 9360 -1281
rect 9394 -1315 9406 -1281
rect 8838 -1423 8854 -1389
rect 8617 -1464 8651 -1445
rect 8411 -1574 8428 -1540
rect 8462 -1574 8481 -1540
rect 8411 -1593 8481 -1574
rect 8533 -1498 8651 -1464
rect 8533 -1540 8583 -1498
rect 8804 -1516 8854 -1423
rect 8980 -1405 9130 -1335
rect 9348 -1350 9406 -1315
rect 9440 -1159 10142 -1117
rect 9440 -1193 9458 -1159
rect 9492 -1193 10090 -1159
rect 10124 -1193 10142 -1159
rect 9440 -1261 10142 -1193
rect 9440 -1295 9458 -1261
rect 9492 -1295 10090 -1261
rect 10124 -1295 10142 -1261
rect 9440 -1335 10142 -1295
rect 8980 -1439 9000 -1405
rect 9034 -1439 9130 -1405
rect 9164 -1403 9260 -1369
rect 9294 -1403 9314 -1369
rect 9164 -1473 9314 -1403
rect 8567 -1574 8583 -1540
rect 8533 -1593 8583 -1574
rect 8673 -1540 8739 -1524
rect 8673 -1574 8689 -1540
rect 8723 -1574 8739 -1540
rect 8673 -1627 8739 -1574
rect 8773 -1540 8854 -1516
rect 8773 -1574 8787 -1540
rect 8821 -1574 8854 -1540
rect 8773 -1593 8854 -1574
rect 8888 -1499 8946 -1482
rect 8888 -1533 8900 -1499
rect 8934 -1533 8946 -1499
rect 8888 -1627 8946 -1533
rect 8980 -1525 9314 -1473
rect 9440 -1403 9518 -1369
rect 9552 -1403 9617 -1369
rect 9651 -1403 9716 -1369
rect 9750 -1403 9770 -1369
rect 9440 -1473 9770 -1403
rect 9804 -1405 10142 -1335
rect 10176 -1188 10234 -1117
rect 10176 -1222 10188 -1188
rect 10222 -1222 10234 -1188
rect 10176 -1281 10234 -1222
rect 10176 -1315 10188 -1281
rect 10222 -1315 10234 -1281
rect 10176 -1350 10234 -1315
rect 10360 -1159 10694 -1117
rect 10360 -1193 10378 -1159
rect 10412 -1193 10642 -1159
rect 10676 -1193 10694 -1159
rect 10360 -1261 10694 -1193
rect 10360 -1295 10378 -1261
rect 10412 -1295 10642 -1261
rect 10676 -1295 10694 -1261
rect 10360 -1335 10694 -1295
rect 10728 -1166 10797 -1151
rect 10728 -1200 10747 -1166
rect 10781 -1200 10797 -1166
rect 10728 -1234 10797 -1200
rect 10728 -1268 10747 -1234
rect 10781 -1268 10797 -1234
rect 10728 -1318 10797 -1268
rect 10831 -1166 10897 -1117
rect 10831 -1200 10847 -1166
rect 10881 -1200 10897 -1166
rect 10831 -1234 10897 -1200
rect 10831 -1268 10847 -1234
rect 10881 -1268 10897 -1234
rect 10831 -1284 10897 -1268
rect 10987 -1166 11057 -1151
rect 10987 -1200 11005 -1166
rect 11039 -1200 11057 -1166
rect 10987 -1234 11057 -1200
rect 10987 -1268 11005 -1234
rect 11039 -1268 11057 -1234
rect 9804 -1439 9824 -1405
rect 9858 -1439 9927 -1405
rect 9961 -1439 10030 -1405
rect 10064 -1439 10142 -1405
rect 10360 -1405 10510 -1335
rect 10728 -1352 10922 -1318
rect 10360 -1439 10380 -1405
rect 10414 -1439 10510 -1405
rect 10544 -1403 10640 -1369
rect 10674 -1403 10694 -1369
rect 10852 -1381 10922 -1352
rect 10987 -1380 11057 -1268
rect 11109 -1167 11159 -1151
rect 11143 -1201 11159 -1167
rect 11109 -1235 11159 -1201
rect 11143 -1269 11159 -1235
rect 11109 -1311 11159 -1269
rect 11249 -1166 11315 -1117
rect 11249 -1200 11265 -1166
rect 11299 -1200 11315 -1166
rect 11249 -1234 11315 -1200
rect 11249 -1268 11265 -1234
rect 11299 -1268 11315 -1234
rect 11249 -1277 11315 -1268
rect 11349 -1167 11430 -1151
rect 11349 -1201 11363 -1167
rect 11397 -1201 11430 -1167
rect 11349 -1235 11430 -1201
rect 11349 -1269 11363 -1235
rect 11397 -1269 11430 -1235
rect 11349 -1306 11430 -1269
rect 11109 -1345 11227 -1311
rect 11193 -1379 11227 -1345
rect 11380 -1355 11430 -1306
rect 11464 -1188 11522 -1117
rect 11464 -1222 11476 -1188
rect 11510 -1222 11522 -1188
rect 11464 -1281 11522 -1222
rect 11464 -1315 11476 -1281
rect 11510 -1315 11522 -1281
rect 11464 -1350 11522 -1315
rect 11648 -1159 11982 -1117
rect 11648 -1193 11666 -1159
rect 11700 -1193 11930 -1159
rect 11964 -1193 11982 -1159
rect 11648 -1261 11982 -1193
rect 11648 -1295 11666 -1261
rect 11700 -1295 11930 -1261
rect 11964 -1295 11982 -1261
rect 11648 -1335 11982 -1295
rect 12384 -1188 12442 -1117
rect 12384 -1222 12396 -1188
rect 12430 -1222 12442 -1188
rect 12384 -1281 12442 -1222
rect 12384 -1315 12396 -1281
rect 12430 -1315 12442 -1281
rect 12476 -1166 12545 -1117
rect 12476 -1200 12502 -1166
rect 12536 -1200 12545 -1166
rect 12476 -1234 12545 -1200
rect 12476 -1268 12502 -1234
rect 12536 -1268 12545 -1234
rect 12476 -1284 12545 -1268
rect 12580 -1173 12631 -1157
rect 12580 -1207 12588 -1173
rect 12622 -1207 12631 -1173
rect 12580 -1261 12631 -1207
rect 10544 -1473 10694 -1403
rect 10728 -1389 10818 -1386
rect 10728 -1423 10764 -1389
rect 10798 -1395 10818 -1389
rect 10728 -1429 10768 -1423
rect 10802 -1429 10818 -1395
rect 10852 -1395 10938 -1381
rect 10852 -1429 10888 -1395
rect 10922 -1429 10938 -1395
rect 10852 -1439 10938 -1429
rect 10987 -1395 11159 -1380
rect 10987 -1429 11109 -1395
rect 11143 -1429 11159 -1395
rect 10987 -1430 11159 -1429
rect 11193 -1395 11346 -1379
rect 11193 -1429 11309 -1395
rect 11343 -1429 11346 -1395
rect 10852 -1463 10922 -1439
rect 8980 -1559 8998 -1525
rect 9032 -1559 9262 -1525
rect 9296 -1559 9314 -1525
rect 8980 -1627 9314 -1559
rect 9348 -1499 9406 -1482
rect 9348 -1533 9360 -1499
rect 9394 -1533 9406 -1499
rect 9348 -1627 9406 -1533
rect 9440 -1532 10142 -1473
rect 9440 -1566 9458 -1532
rect 9492 -1566 10090 -1532
rect 10124 -1566 10142 -1532
rect 9440 -1627 10142 -1566
rect 10176 -1499 10234 -1482
rect 10176 -1533 10188 -1499
rect 10222 -1533 10234 -1499
rect 10176 -1627 10234 -1533
rect 10360 -1525 10694 -1473
rect 10360 -1559 10378 -1525
rect 10412 -1559 10642 -1525
rect 10676 -1559 10694 -1525
rect 10360 -1627 10694 -1559
rect 10728 -1497 10922 -1463
rect 10728 -1540 10794 -1497
rect 10728 -1574 10747 -1540
rect 10781 -1574 10794 -1540
rect 10728 -1593 10794 -1574
rect 10828 -1540 10894 -1531
rect 10828 -1574 10844 -1540
rect 10878 -1574 10894 -1540
rect 10828 -1627 10894 -1574
rect 10987 -1540 11057 -1430
rect 11193 -1445 11346 -1429
rect 11380 -1389 11387 -1355
rect 11421 -1389 11430 -1355
rect 11193 -1464 11227 -1445
rect 10987 -1574 11004 -1540
rect 11038 -1574 11057 -1540
rect 10987 -1593 11057 -1574
rect 11109 -1498 11227 -1464
rect 11109 -1540 11159 -1498
rect 11380 -1516 11430 -1389
rect 11648 -1405 11798 -1335
rect 12384 -1350 12442 -1315
rect 12580 -1295 12588 -1261
rect 12622 -1295 12631 -1261
rect 12665 -1166 12717 -1117
rect 12665 -1200 12674 -1166
rect 12708 -1200 12717 -1166
rect 12665 -1234 12717 -1200
rect 12665 -1268 12674 -1234
rect 12708 -1268 12717 -1234
rect 12665 -1284 12717 -1268
rect 12752 -1173 12803 -1157
rect 12752 -1207 12760 -1173
rect 12794 -1207 12803 -1173
rect 12752 -1261 12803 -1207
rect 12580 -1318 12631 -1295
rect 12752 -1295 12760 -1261
rect 12794 -1295 12803 -1261
rect 12837 -1166 12889 -1117
rect 12837 -1200 12846 -1166
rect 12880 -1200 12889 -1166
rect 12837 -1234 12889 -1200
rect 12837 -1268 12846 -1234
rect 12880 -1268 12889 -1234
rect 12837 -1284 12889 -1268
rect 12923 -1173 12975 -1157
rect 12923 -1207 12932 -1173
rect 12966 -1207 12975 -1173
rect 12923 -1261 12975 -1207
rect 12752 -1318 12803 -1295
rect 12923 -1295 12932 -1261
rect 12966 -1295 12975 -1261
rect 13009 -1166 13086 -1117
rect 13009 -1200 13018 -1166
rect 13052 -1200 13086 -1166
rect 13009 -1234 13086 -1200
rect 13009 -1268 13018 -1234
rect 13052 -1268 13086 -1234
rect 13009 -1284 13086 -1268
rect 13120 -1188 13178 -1117
rect 13120 -1222 13132 -1188
rect 13166 -1222 13178 -1188
rect 13120 -1281 13178 -1222
rect 12923 -1318 12975 -1295
rect 13120 -1315 13132 -1281
rect 13166 -1315 13178 -1281
rect 12480 -1352 13086 -1318
rect 13120 -1350 13178 -1315
rect 13212 -1159 13546 -1117
rect 13212 -1193 13230 -1159
rect 13264 -1193 13494 -1159
rect 13528 -1193 13546 -1159
rect 13212 -1261 13546 -1193
rect 13212 -1295 13230 -1261
rect 13264 -1295 13494 -1261
rect 13528 -1295 13546 -1261
rect 13212 -1335 13546 -1295
rect 11648 -1439 11668 -1405
rect 11702 -1439 11798 -1405
rect 11832 -1403 11928 -1369
rect 11962 -1403 11982 -1369
rect 11832 -1473 11982 -1403
rect 11143 -1574 11159 -1540
rect 11109 -1593 11159 -1574
rect 11249 -1540 11315 -1524
rect 11249 -1574 11265 -1540
rect 11299 -1574 11315 -1540
rect 11249 -1627 11315 -1574
rect 11349 -1540 11430 -1516
rect 11349 -1574 11363 -1540
rect 11397 -1574 11430 -1540
rect 11349 -1593 11430 -1574
rect 11464 -1499 11522 -1482
rect 11464 -1533 11476 -1499
rect 11510 -1533 11522 -1499
rect 11464 -1627 11522 -1533
rect 11648 -1525 11982 -1473
rect 12480 -1465 12514 -1352
rect 13026 -1385 13086 -1352
rect 12548 -1392 12991 -1386
rect 12548 -1426 12558 -1392
rect 12592 -1395 12642 -1392
rect 12676 -1395 12739 -1392
rect 12773 -1395 12836 -1392
rect 12870 -1395 12942 -1392
rect 12548 -1429 12574 -1426
rect 12608 -1429 12642 -1395
rect 12676 -1429 12710 -1395
rect 12773 -1426 12778 -1395
rect 12744 -1429 12778 -1426
rect 12812 -1426 12836 -1395
rect 12812 -1429 12846 -1426
rect 12880 -1429 12914 -1395
rect 12976 -1426 12991 -1392
rect 12948 -1429 12991 -1426
rect 12548 -1431 12991 -1429
rect 13026 -1419 13038 -1385
rect 13072 -1419 13086 -1385
rect 13026 -1457 13086 -1419
rect 13026 -1465 13038 -1457
rect 11648 -1559 11666 -1525
rect 11700 -1559 11930 -1525
rect 11964 -1559 11982 -1525
rect 11648 -1627 11982 -1559
rect 12384 -1499 12442 -1482
rect 12480 -1491 13038 -1465
rect 13072 -1491 13086 -1457
rect 13212 -1403 13232 -1369
rect 13266 -1403 13362 -1369
rect 13212 -1473 13362 -1403
rect 13396 -1405 13546 -1335
rect 13580 -1188 13638 -1117
rect 13580 -1222 13592 -1188
rect 13626 -1222 13638 -1188
rect 13580 -1281 13638 -1222
rect 13674 -1159 13733 -1117
rect 13674 -1193 13690 -1159
rect 13724 -1193 13733 -1159
rect 13674 -1227 13733 -1193
rect 13674 -1261 13690 -1227
rect 13724 -1261 13733 -1227
rect 13674 -1279 13733 -1261
rect 13769 -1167 13818 -1151
rect 13769 -1201 13776 -1167
rect 13810 -1201 13818 -1167
rect 13769 -1235 13818 -1201
rect 13769 -1269 13776 -1235
rect 13810 -1269 13818 -1235
rect 13580 -1315 13592 -1281
rect 13626 -1315 13638 -1281
rect 13580 -1350 13638 -1315
rect 13769 -1379 13818 -1269
rect 13853 -1159 13905 -1117
rect 14025 -1118 15280 -1117
rect 13853 -1193 13862 -1159
rect 13896 -1193 13905 -1159
rect 13853 -1227 13905 -1193
rect 13853 -1261 13862 -1227
rect 13896 -1261 13905 -1227
rect 13853 -1279 13905 -1261
rect 13941 -1175 13991 -1152
rect 13941 -1209 13948 -1175
rect 13982 -1209 13991 -1175
rect 13941 -1243 13991 -1209
rect 13941 -1277 13948 -1243
rect 13982 -1277 13991 -1243
rect 14025 -1159 14077 -1118
rect 14025 -1193 14034 -1159
rect 14068 -1193 14077 -1159
rect 14025 -1227 14077 -1193
rect 14025 -1261 14034 -1227
rect 14068 -1261 14077 -1227
rect 14025 -1277 14077 -1261
rect 14111 -1203 14163 -1152
rect 14111 -1237 14120 -1203
rect 14154 -1237 14163 -1203
rect 13941 -1379 13991 -1277
rect 14111 -1289 14163 -1237
rect 14197 -1183 14249 -1118
rect 14197 -1217 14206 -1183
rect 14240 -1217 14249 -1183
rect 14197 -1263 14249 -1217
rect 14283 -1203 14335 -1152
rect 14283 -1237 14292 -1203
rect 14326 -1237 14335 -1203
rect 14111 -1323 14120 -1289
rect 14154 -1297 14163 -1289
rect 14283 -1289 14335 -1237
rect 14369 -1183 14421 -1118
rect 14369 -1217 14378 -1183
rect 14412 -1217 14421 -1183
rect 14369 -1263 14421 -1217
rect 14455 -1203 14507 -1152
rect 14455 -1237 14464 -1203
rect 14498 -1237 14507 -1203
rect 14283 -1297 14292 -1289
rect 14154 -1323 14292 -1297
rect 14326 -1297 14335 -1289
rect 14455 -1289 14507 -1237
rect 14541 -1183 14593 -1118
rect 14541 -1217 14550 -1183
rect 14584 -1217 14593 -1183
rect 14541 -1263 14593 -1217
rect 14627 -1203 14679 -1152
rect 14627 -1237 14636 -1203
rect 14670 -1237 14679 -1203
rect 14455 -1297 14464 -1289
rect 14326 -1323 14464 -1297
rect 14498 -1297 14507 -1289
rect 14627 -1289 14679 -1237
rect 14713 -1183 14762 -1118
rect 14713 -1217 14722 -1183
rect 14756 -1217 14762 -1183
rect 14713 -1263 14762 -1217
rect 14796 -1203 14848 -1152
rect 14796 -1237 14807 -1203
rect 14841 -1237 14848 -1203
rect 14627 -1297 14636 -1289
rect 14498 -1323 14636 -1297
rect 14670 -1297 14679 -1289
rect 14796 -1289 14848 -1237
rect 14885 -1183 14934 -1118
rect 14885 -1217 14893 -1183
rect 14927 -1217 14934 -1183
rect 14885 -1263 14934 -1217
rect 14968 -1203 15020 -1152
rect 14968 -1237 14979 -1203
rect 15013 -1237 15020 -1203
rect 14796 -1297 14807 -1289
rect 14670 -1323 14807 -1297
rect 14841 -1297 14848 -1289
rect 14968 -1289 15020 -1237
rect 15057 -1183 15106 -1118
rect 15057 -1217 15065 -1183
rect 15099 -1217 15106 -1183
rect 15057 -1263 15106 -1217
rect 15140 -1203 15192 -1152
rect 15140 -1237 15151 -1203
rect 15185 -1237 15192 -1203
rect 14968 -1297 14979 -1289
rect 14841 -1323 14979 -1297
rect 15013 -1297 15020 -1289
rect 15140 -1289 15192 -1237
rect 15229 -1183 15280 -1118
rect 15229 -1217 15237 -1183
rect 15271 -1217 15280 -1183
rect 15229 -1263 15280 -1217
rect 15314 -1203 15372 -1152
rect 15314 -1237 15323 -1203
rect 15357 -1237 15372 -1203
rect 15140 -1297 15151 -1289
rect 15013 -1323 15151 -1297
rect 15185 -1300 15192 -1289
rect 15314 -1289 15372 -1237
rect 15406 -1183 15460 -1117
rect 15406 -1217 15409 -1183
rect 15443 -1217 15460 -1183
rect 15406 -1266 15460 -1217
rect 15512 -1188 15570 -1117
rect 15512 -1222 15524 -1188
rect 15558 -1222 15570 -1188
rect 15314 -1300 15323 -1289
rect 15185 -1323 15323 -1300
rect 15357 -1300 15372 -1289
rect 15512 -1281 15570 -1222
rect 15357 -1323 15460 -1300
rect 14111 -1338 15460 -1323
rect 14111 -1345 15248 -1338
rect 15227 -1372 15248 -1345
rect 15282 -1339 15460 -1338
rect 15282 -1372 15340 -1339
rect 15227 -1373 15340 -1372
rect 15374 -1373 15460 -1339
rect 15512 -1315 15524 -1281
rect 15558 -1315 15570 -1281
rect 15512 -1350 15570 -1315
rect 15604 -1159 16673 -1117
rect 15604 -1193 15622 -1159
rect 15656 -1193 16622 -1159
rect 16656 -1193 16673 -1159
rect 15604 -1261 16673 -1193
rect 15604 -1295 15622 -1261
rect 15656 -1295 16622 -1261
rect 16656 -1295 16673 -1261
rect 15604 -1335 16673 -1295
rect 13396 -1439 13492 -1405
rect 13526 -1439 13546 -1405
rect 13672 -1395 13735 -1379
rect 13672 -1422 13692 -1395
rect 13672 -1456 13684 -1422
rect 13726 -1429 13735 -1395
rect 13718 -1456 13735 -1429
rect 12480 -1499 13086 -1491
rect 13120 -1499 13178 -1482
rect 12384 -1533 12396 -1499
rect 12430 -1533 12442 -1499
rect 12384 -1627 12442 -1533
rect 12572 -1549 12631 -1533
rect 12572 -1583 12588 -1549
rect 12622 -1583 12631 -1549
rect 12572 -1627 12631 -1583
rect 12665 -1538 12717 -1499
rect 12665 -1572 12674 -1538
rect 12708 -1572 12717 -1538
rect 12665 -1588 12717 -1572
rect 12751 -1549 12803 -1533
rect 12751 -1583 12760 -1549
rect 12794 -1583 12803 -1549
rect 12751 -1627 12803 -1583
rect 12837 -1538 12888 -1499
rect 13120 -1533 13132 -1499
rect 13166 -1533 13178 -1499
rect 12837 -1572 12846 -1538
rect 12880 -1572 12888 -1538
rect 12837 -1588 12888 -1572
rect 12922 -1549 12982 -1533
rect 12922 -1583 12932 -1549
rect 12966 -1583 12982 -1549
rect 12922 -1627 12982 -1583
rect 13120 -1627 13178 -1533
rect 13212 -1525 13546 -1473
rect 13212 -1559 13230 -1525
rect 13264 -1559 13494 -1525
rect 13528 -1559 13546 -1525
rect 13212 -1627 13546 -1559
rect 13580 -1499 13638 -1482
rect 13672 -1491 13735 -1456
rect 13769 -1395 15193 -1379
rect 13769 -1429 14119 -1395
rect 14153 -1429 14187 -1395
rect 14221 -1429 14255 -1395
rect 14289 -1429 14323 -1395
rect 14357 -1429 14391 -1395
rect 14425 -1429 14459 -1395
rect 14493 -1429 14527 -1395
rect 14561 -1429 14595 -1395
rect 14629 -1429 14663 -1395
rect 14697 -1429 14731 -1395
rect 14765 -1429 14799 -1395
rect 14833 -1429 14867 -1395
rect 14901 -1429 14935 -1395
rect 14969 -1429 15003 -1395
rect 15037 -1429 15071 -1395
rect 15105 -1429 15139 -1395
rect 15173 -1429 15193 -1395
rect 13580 -1533 13592 -1499
rect 13626 -1533 13638 -1499
rect 13580 -1627 13638 -1533
rect 13672 -1551 13733 -1525
rect 13672 -1585 13690 -1551
rect 13724 -1585 13733 -1551
rect 13672 -1627 13733 -1585
rect 13769 -1538 13819 -1429
rect 13769 -1572 13776 -1538
rect 13810 -1572 13819 -1538
rect 13769 -1591 13819 -1572
rect 13853 -1538 13905 -1522
rect 13853 -1572 13862 -1538
rect 13896 -1572 13905 -1538
rect 13853 -1627 13905 -1572
rect 13941 -1538 13991 -1429
rect 15227 -1434 15460 -1373
rect 15227 -1463 15248 -1434
rect 14111 -1468 15248 -1463
rect 15282 -1468 15341 -1434
rect 15375 -1468 15460 -1434
rect 14111 -1497 15460 -1468
rect 15604 -1403 15682 -1369
rect 15716 -1403 15810 -1369
rect 15844 -1403 15938 -1369
rect 15972 -1403 16066 -1369
rect 16100 -1403 16120 -1369
rect 15604 -1473 16120 -1403
rect 16154 -1405 16673 -1335
rect 16154 -1439 16174 -1405
rect 16208 -1439 16302 -1405
rect 16336 -1439 16430 -1405
rect 16464 -1439 16558 -1405
rect 16592 -1439 16673 -1405
rect 13941 -1572 13948 -1538
rect 13982 -1572 13991 -1538
rect 13941 -1591 13991 -1572
rect 14025 -1538 14077 -1515
rect 14025 -1572 14034 -1538
rect 14068 -1572 14077 -1538
rect 14025 -1627 14077 -1572
rect 14111 -1538 14163 -1497
rect 14111 -1572 14120 -1538
rect 14154 -1572 14163 -1538
rect 14111 -1588 14163 -1572
rect 14197 -1547 14249 -1531
rect 14197 -1581 14206 -1547
rect 14240 -1581 14249 -1547
rect 14197 -1627 14249 -1581
rect 14283 -1538 14335 -1497
rect 14283 -1572 14292 -1538
rect 14326 -1572 14335 -1538
rect 14283 -1588 14335 -1572
rect 14369 -1547 14421 -1531
rect 14369 -1581 14378 -1547
rect 14412 -1581 14421 -1547
rect 14369 -1627 14421 -1581
rect 14455 -1538 14507 -1497
rect 14455 -1572 14464 -1538
rect 14498 -1572 14507 -1538
rect 14455 -1588 14507 -1572
rect 14541 -1547 14590 -1531
rect 14541 -1581 14550 -1547
rect 14584 -1581 14590 -1547
rect 14541 -1627 14590 -1581
rect 14624 -1538 14679 -1497
rect 14624 -1572 14636 -1538
rect 14670 -1572 14679 -1538
rect 14624 -1588 14679 -1572
rect 14713 -1547 14762 -1531
rect 14713 -1581 14722 -1547
rect 14756 -1581 14762 -1547
rect 14713 -1627 14762 -1581
rect 14796 -1538 14848 -1497
rect 14796 -1572 14807 -1538
rect 14841 -1572 14848 -1538
rect 14796 -1588 14848 -1572
rect 14884 -1547 14934 -1531
rect 14884 -1581 14893 -1547
rect 14927 -1581 14934 -1547
rect 14884 -1627 14934 -1581
rect 14968 -1538 15020 -1497
rect 14968 -1572 14979 -1538
rect 15013 -1572 15020 -1538
rect 14968 -1588 15020 -1572
rect 15056 -1547 15106 -1531
rect 15056 -1581 15065 -1547
rect 15099 -1581 15106 -1547
rect 15056 -1627 15106 -1581
rect 15140 -1538 15192 -1497
rect 15140 -1572 15151 -1538
rect 15185 -1572 15192 -1538
rect 15140 -1588 15192 -1572
rect 15228 -1547 15280 -1531
rect 15228 -1581 15237 -1547
rect 15271 -1581 15280 -1547
rect 15228 -1627 15280 -1581
rect 15314 -1538 15366 -1497
rect 15512 -1499 15570 -1482
rect 15314 -1572 15323 -1538
rect 15357 -1572 15366 -1538
rect 15314 -1588 15366 -1572
rect 15400 -1547 15460 -1531
rect 15400 -1581 15409 -1547
rect 15443 -1581 15460 -1547
rect 15400 -1627 15460 -1581
rect 15512 -1533 15524 -1499
rect 15558 -1533 15570 -1499
rect 15512 -1627 15570 -1533
rect 15604 -1532 16673 -1473
rect 15604 -1566 15622 -1532
rect 15656 -1566 16622 -1532
rect 16656 -1566 16673 -1532
rect 15604 -1627 16673 -1566
rect -2997 -1661 -2968 -1627
rect -2934 -1661 -2876 -1627
rect -2842 -1661 -2784 -1627
rect -2750 -1661 -2692 -1627
rect -2658 -1661 -2600 -1627
rect -2566 -1661 -2508 -1627
rect -2474 -1661 -2416 -1627
rect -2382 -1661 -2324 -1627
rect -2290 -1661 -2232 -1627
rect -2198 -1661 -2140 -1627
rect -2106 -1661 -2048 -1627
rect -2014 -1661 -1956 -1627
rect -1922 -1661 -1864 -1627
rect -1830 -1661 -1772 -1627
rect -1738 -1661 -1680 -1627
rect -1646 -1661 -1588 -1627
rect -1554 -1661 -1496 -1627
rect -1462 -1661 -1404 -1627
rect -1370 -1661 -1312 -1627
rect -1278 -1661 -1220 -1627
rect -1186 -1661 -1128 -1627
rect -1094 -1661 -1036 -1627
rect -1002 -1661 -944 -1627
rect -910 -1661 -852 -1627
rect -818 -1661 -760 -1627
rect -726 -1661 -668 -1627
rect -634 -1661 -576 -1627
rect -542 -1661 -484 -1627
rect -450 -1661 -392 -1627
rect -358 -1661 -300 -1627
rect -266 -1661 -208 -1627
rect -174 -1661 -116 -1627
rect -82 -1661 -24 -1627
rect 10 -1661 68 -1627
rect 102 -1661 160 -1627
rect 194 -1661 252 -1627
rect 286 -1661 344 -1627
rect 378 -1661 436 -1627
rect 470 -1661 528 -1627
rect 562 -1661 620 -1627
rect 654 -1661 712 -1627
rect 746 -1661 804 -1627
rect 838 -1661 896 -1627
rect 930 -1661 988 -1627
rect 1022 -1661 1080 -1627
rect 1114 -1661 1172 -1627
rect 1206 -1661 1264 -1627
rect 1298 -1661 1356 -1627
rect 1390 -1661 1448 -1627
rect 1482 -1661 1540 -1627
rect 1574 -1661 1632 -1627
rect 1666 -1661 1724 -1627
rect 1758 -1661 1816 -1627
rect 1850 -1661 1908 -1627
rect 1942 -1661 2000 -1627
rect 2034 -1661 2092 -1627
rect 2126 -1661 2184 -1627
rect 2218 -1661 2276 -1627
rect 2310 -1661 2368 -1627
rect 2402 -1661 2460 -1627
rect 2494 -1661 2552 -1627
rect 2586 -1661 2644 -1627
rect 2678 -1661 2736 -1627
rect 2770 -1661 2828 -1627
rect 2862 -1661 2920 -1627
rect 2954 -1661 3012 -1627
rect 3046 -1661 3104 -1627
rect 3138 -1661 3196 -1627
rect 3230 -1661 3288 -1627
rect 3322 -1661 3380 -1627
rect 3414 -1661 3472 -1627
rect 3506 -1661 3564 -1627
rect 3598 -1661 3656 -1627
rect 3690 -1661 3748 -1627
rect 3782 -1661 3840 -1627
rect 3874 -1661 3932 -1627
rect 3966 -1661 4024 -1627
rect 4058 -1661 4116 -1627
rect 4150 -1661 4208 -1627
rect 4242 -1661 4300 -1627
rect 4334 -1661 4392 -1627
rect 4426 -1661 4484 -1627
rect 4518 -1661 4576 -1627
rect 4610 -1661 4668 -1627
rect 4702 -1661 4760 -1627
rect 4794 -1661 4852 -1627
rect 4886 -1661 4944 -1627
rect 4978 -1661 5036 -1627
rect 5070 -1661 5128 -1627
rect 5162 -1661 5220 -1627
rect 5254 -1661 5312 -1627
rect 5346 -1661 5404 -1627
rect 5438 -1661 5496 -1627
rect 5530 -1661 5588 -1627
rect 5622 -1661 5680 -1627
rect 5714 -1661 5772 -1627
rect 5806 -1661 5864 -1627
rect 5898 -1661 5956 -1627
rect 5990 -1661 6048 -1627
rect 6082 -1661 6140 -1627
rect 6174 -1661 6232 -1627
rect 6266 -1661 6324 -1627
rect 6358 -1661 6416 -1627
rect 6450 -1661 6508 -1627
rect 6542 -1661 6600 -1627
rect 6634 -1661 6692 -1627
rect 6726 -1661 6784 -1627
rect 6818 -1661 6876 -1627
rect 6910 -1661 6968 -1627
rect 7002 -1661 7060 -1627
rect 7094 -1661 7152 -1627
rect 7186 -1661 7244 -1627
rect 7278 -1661 7336 -1627
rect 7370 -1661 7428 -1627
rect 7462 -1661 7520 -1627
rect 7554 -1661 7612 -1627
rect 7646 -1661 7704 -1627
rect 7738 -1661 7796 -1627
rect 7830 -1661 7888 -1627
rect 7922 -1661 7980 -1627
rect 8014 -1661 8072 -1627
rect 8106 -1661 8164 -1627
rect 8198 -1661 8256 -1627
rect 8290 -1661 8348 -1627
rect 8382 -1661 8440 -1627
rect 8474 -1661 8532 -1627
rect 8566 -1661 8624 -1627
rect 8658 -1661 8716 -1627
rect 8750 -1661 8808 -1627
rect 8842 -1661 8900 -1627
rect 8934 -1661 8992 -1627
rect 9026 -1661 9084 -1627
rect 9118 -1661 9176 -1627
rect 9210 -1661 9268 -1627
rect 9302 -1661 9360 -1627
rect 9394 -1661 9452 -1627
rect 9486 -1661 9544 -1627
rect 9578 -1661 9636 -1627
rect 9670 -1661 9728 -1627
rect 9762 -1661 9820 -1627
rect 9854 -1661 9912 -1627
rect 9946 -1661 10004 -1627
rect 10038 -1661 10096 -1627
rect 10130 -1661 10188 -1627
rect 10222 -1661 10280 -1627
rect 10314 -1661 10372 -1627
rect 10406 -1661 10464 -1627
rect 10498 -1661 10556 -1627
rect 10590 -1661 10648 -1627
rect 10682 -1661 10740 -1627
rect 10774 -1661 10832 -1627
rect 10866 -1661 10924 -1627
rect 10958 -1661 11016 -1627
rect 11050 -1661 11108 -1627
rect 11142 -1661 11200 -1627
rect 11234 -1661 11292 -1627
rect 11326 -1661 11384 -1627
rect 11418 -1661 11476 -1627
rect 11510 -1661 11568 -1627
rect 11602 -1661 11660 -1627
rect 11694 -1661 11752 -1627
rect 11786 -1661 11844 -1627
rect 11878 -1661 11936 -1627
rect 11970 -1661 12028 -1627
rect 12062 -1661 12120 -1627
rect 12154 -1661 12212 -1627
rect 12246 -1661 12304 -1627
rect 12338 -1661 12396 -1627
rect 12430 -1661 12488 -1627
rect 12522 -1661 12580 -1627
rect 12614 -1661 12672 -1627
rect 12706 -1661 12764 -1627
rect 12798 -1661 12856 -1627
rect 12890 -1661 12948 -1627
rect 12982 -1661 13040 -1627
rect 13074 -1661 13132 -1627
rect 13166 -1661 13224 -1627
rect 13258 -1661 13316 -1627
rect 13350 -1661 13408 -1627
rect 13442 -1661 13500 -1627
rect 13534 -1661 13592 -1627
rect 13626 -1661 13684 -1627
rect 13718 -1661 13776 -1627
rect 13810 -1661 13868 -1627
rect 13902 -1661 13960 -1627
rect 13994 -1661 14052 -1627
rect 14086 -1661 14144 -1627
rect 14178 -1661 14236 -1627
rect 14270 -1661 14328 -1627
rect 14362 -1661 14420 -1627
rect 14454 -1661 14512 -1627
rect 14546 -1661 14604 -1627
rect 14638 -1661 14696 -1627
rect 14730 -1661 14788 -1627
rect 14822 -1661 14880 -1627
rect 14914 -1661 14972 -1627
rect 15006 -1661 15064 -1627
rect 15098 -1661 15156 -1627
rect 15190 -1661 15248 -1627
rect 15282 -1661 15340 -1627
rect 15374 -1661 15432 -1627
rect 15466 -1661 15524 -1627
rect 15558 -1661 15616 -1627
rect 15650 -1661 15708 -1627
rect 15742 -1661 15800 -1627
rect 15834 -1661 15892 -1627
rect 15926 -1661 15984 -1627
rect 16018 -1661 16076 -1627
rect 16110 -1661 16168 -1627
rect 16202 -1661 16260 -1627
rect 16294 -1661 16352 -1627
rect 16386 -1661 16444 -1627
rect 16478 -1661 16536 -1627
rect 16570 -1661 16628 -1627
rect 16662 -1661 16691 -1627
rect -2980 -1722 -2278 -1661
rect -2980 -1756 -2962 -1722
rect -2928 -1756 -2330 -1722
rect -2296 -1756 -2278 -1722
rect -2980 -1815 -2278 -1756
rect -2244 -1755 -2186 -1661
rect -2244 -1789 -2232 -1755
rect -2198 -1789 -2186 -1755
rect -2244 -1806 -2186 -1789
rect -1600 -1722 -898 -1661
rect -1600 -1756 -1582 -1722
rect -1548 -1756 -950 -1722
rect -916 -1756 -898 -1722
rect -1600 -1815 -898 -1756
rect -2980 -1883 -2902 -1849
rect -2868 -1883 -2799 -1849
rect -2765 -1883 -2696 -1849
rect -2662 -1883 -2642 -1849
rect -2980 -1953 -2642 -1883
rect -2608 -1885 -2278 -1815
rect -2608 -1919 -2588 -1885
rect -2554 -1919 -2489 -1885
rect -2455 -1919 -2390 -1885
rect -2356 -1919 -2278 -1885
rect -1600 -1883 -1522 -1849
rect -1488 -1883 -1419 -1849
rect -1385 -1883 -1316 -1849
rect -1282 -1883 -1262 -1849
rect -2980 -1993 -2278 -1953
rect -2980 -2027 -2962 -1993
rect -2928 -2027 -2330 -1993
rect -2296 -2027 -2278 -1993
rect -2980 -2095 -2278 -2027
rect -2980 -2129 -2962 -2095
rect -2928 -2129 -2330 -2095
rect -2296 -2129 -2278 -2095
rect -2980 -2171 -2278 -2129
rect -2244 -1973 -2186 -1938
rect -2244 -2007 -2232 -1973
rect -2198 -2007 -2186 -1973
rect -2244 -2066 -2186 -2007
rect -2244 -2100 -2232 -2066
rect -2198 -2100 -2186 -2066
rect -2244 -2171 -2186 -2100
rect -1600 -1953 -1262 -1883
rect -1228 -1885 -898 -1815
rect -1228 -1919 -1208 -1885
rect -1174 -1919 -1109 -1885
rect -1075 -1919 -1010 -1885
rect -976 -1919 -898 -1885
rect -864 -1714 -783 -1695
rect -864 -1748 -831 -1714
rect -797 -1748 -783 -1714
rect -864 -1772 -783 -1748
rect -749 -1714 -683 -1661
rect -749 -1748 -733 -1714
rect -699 -1748 -683 -1714
rect -749 -1764 -683 -1748
rect -593 -1714 -543 -1695
rect -593 -1748 -577 -1714
rect -864 -1900 -814 -1772
rect -593 -1790 -543 -1748
rect -661 -1824 -543 -1790
rect -491 -1714 -421 -1695
rect -491 -1748 -472 -1714
rect -438 -1748 -421 -1714
rect -661 -1843 -627 -1824
rect -864 -1934 -856 -1900
rect -822 -1934 -814 -1900
rect -780 -1859 -627 -1843
rect -491 -1858 -421 -1748
rect -328 -1714 -262 -1661
rect -328 -1748 -312 -1714
rect -278 -1748 -262 -1714
rect -328 -1757 -262 -1748
rect -228 -1714 -162 -1695
rect -228 -1748 -215 -1714
rect -181 -1748 -162 -1714
rect -228 -1791 -162 -1748
rect -356 -1825 -162 -1791
rect -128 -1755 -70 -1661
rect -128 -1789 -116 -1755
rect -82 -1789 -70 -1755
rect -128 -1806 -70 -1789
rect -36 -1729 298 -1661
rect -36 -1763 -18 -1729
rect 16 -1763 246 -1729
rect 280 -1763 298 -1729
rect -36 -1815 298 -1763
rect 332 -1755 390 -1661
rect 332 -1789 344 -1755
rect 378 -1789 390 -1755
rect 332 -1806 390 -1789
rect 424 -1714 505 -1695
rect 424 -1748 457 -1714
rect 491 -1748 505 -1714
rect 424 -1772 505 -1748
rect 539 -1714 605 -1661
rect 539 -1748 555 -1714
rect 589 -1748 605 -1714
rect 539 -1764 605 -1748
rect 695 -1714 745 -1695
rect 695 -1748 711 -1714
rect -356 -1849 -286 -1825
rect -780 -1893 -777 -1859
rect -743 -1893 -627 -1859
rect -780 -1909 -627 -1893
rect -593 -1859 -421 -1858
rect -593 -1893 -577 -1859
rect -543 -1893 -421 -1859
rect -593 -1908 -421 -1893
rect -372 -1859 -286 -1849
rect -372 -1893 -356 -1859
rect -322 -1893 -286 -1859
rect -372 -1907 -286 -1893
rect -252 -1893 -236 -1859
rect -202 -1865 -162 -1859
rect -252 -1899 -210 -1893
rect -176 -1899 -162 -1865
rect -252 -1902 -162 -1899
rect -36 -1883 -16 -1849
rect 18 -1883 114 -1849
rect -1600 -1993 -898 -1953
rect -1600 -2027 -1582 -1993
rect -1548 -2027 -950 -1993
rect -916 -2027 -898 -1993
rect -1600 -2095 -898 -2027
rect -1600 -2129 -1582 -2095
rect -1548 -2129 -950 -2095
rect -916 -2129 -898 -2095
rect -1600 -2171 -898 -2129
rect -864 -1982 -814 -1934
rect -661 -1943 -627 -1909
rect -661 -1977 -543 -1943
rect -864 -2019 -783 -1982
rect -864 -2053 -831 -2019
rect -797 -2053 -783 -2019
rect -864 -2087 -783 -2053
rect -864 -2121 -831 -2087
rect -797 -2121 -783 -2087
rect -864 -2137 -783 -2121
rect -749 -2020 -683 -2011
rect -749 -2054 -733 -2020
rect -699 -2054 -683 -2020
rect -749 -2088 -683 -2054
rect -749 -2122 -733 -2088
rect -699 -2122 -683 -2088
rect -749 -2171 -683 -2122
rect -593 -2019 -543 -1977
rect -593 -2053 -577 -2019
rect -593 -2087 -543 -2053
rect -593 -2121 -577 -2087
rect -593 -2137 -543 -2121
rect -491 -2020 -421 -1908
rect -356 -1936 -286 -1907
rect -356 -1970 -162 -1936
rect -491 -2054 -473 -2020
rect -439 -2054 -421 -2020
rect -491 -2088 -421 -2054
rect -491 -2122 -473 -2088
rect -439 -2122 -421 -2088
rect -491 -2137 -421 -2122
rect -331 -2020 -265 -2004
rect -331 -2054 -315 -2020
rect -281 -2054 -265 -2020
rect -331 -2088 -265 -2054
rect -331 -2122 -315 -2088
rect -281 -2122 -265 -2088
rect -331 -2171 -265 -2122
rect -231 -2020 -162 -1970
rect -231 -2054 -215 -2020
rect -181 -2054 -162 -2020
rect -231 -2088 -162 -2054
rect -231 -2122 -215 -2088
rect -181 -2122 -162 -2088
rect -231 -2137 -162 -2122
rect -128 -1973 -70 -1938
rect -128 -2007 -116 -1973
rect -82 -2007 -70 -1973
rect -128 -2066 -70 -2007
rect -128 -2100 -116 -2066
rect -82 -2100 -70 -2066
rect -128 -2171 -70 -2100
rect -36 -1953 114 -1883
rect 148 -1885 298 -1815
rect 148 -1919 244 -1885
rect 278 -1919 298 -1885
rect 424 -1900 474 -1772
rect 695 -1790 745 -1748
rect 627 -1824 745 -1790
rect 797 -1714 867 -1695
rect 797 -1748 816 -1714
rect 850 -1748 867 -1714
rect 627 -1843 661 -1824
rect 424 -1934 432 -1900
rect 466 -1934 474 -1900
rect 508 -1859 661 -1843
rect 797 -1858 867 -1748
rect 960 -1714 1026 -1661
rect 960 -1748 976 -1714
rect 1010 -1748 1026 -1714
rect 960 -1757 1026 -1748
rect 1060 -1714 1126 -1695
rect 1060 -1748 1073 -1714
rect 1107 -1748 1126 -1714
rect 1060 -1791 1126 -1748
rect 932 -1825 1126 -1791
rect 1160 -1755 1218 -1661
rect 1160 -1789 1172 -1755
rect 1206 -1789 1218 -1755
rect 1160 -1806 1218 -1789
rect 1252 -1729 1586 -1661
rect 1252 -1763 1270 -1729
rect 1304 -1763 1534 -1729
rect 1568 -1763 1586 -1729
rect 1252 -1815 1586 -1763
rect 1620 -1755 1678 -1661
rect 1620 -1789 1632 -1755
rect 1666 -1789 1678 -1755
rect 1620 -1806 1678 -1789
rect 1712 -1722 2414 -1661
rect 1712 -1756 1730 -1722
rect 1764 -1756 2362 -1722
rect 2396 -1756 2414 -1722
rect 1712 -1815 2414 -1756
rect 2448 -1755 2506 -1661
rect 2448 -1789 2460 -1755
rect 2494 -1789 2506 -1755
rect 2448 -1806 2506 -1789
rect 2540 -1729 2874 -1661
rect 2540 -1763 2558 -1729
rect 2592 -1763 2822 -1729
rect 2856 -1763 2874 -1729
rect 2540 -1815 2874 -1763
rect 2908 -1755 2966 -1661
rect 2908 -1789 2920 -1755
rect 2954 -1789 2966 -1755
rect 2908 -1806 2966 -1789
rect 3000 -1714 3081 -1695
rect 3000 -1748 3033 -1714
rect 3067 -1748 3081 -1714
rect 3000 -1772 3081 -1748
rect 3115 -1714 3181 -1661
rect 3115 -1748 3131 -1714
rect 3165 -1748 3181 -1714
rect 3115 -1764 3181 -1748
rect 3271 -1714 3321 -1695
rect 3271 -1748 3287 -1714
rect 932 -1849 1002 -1825
rect 508 -1893 511 -1859
rect 545 -1893 661 -1859
rect 508 -1909 661 -1893
rect 695 -1859 867 -1858
rect 695 -1893 711 -1859
rect 745 -1893 867 -1859
rect 695 -1908 867 -1893
rect 916 -1859 1002 -1849
rect 916 -1893 932 -1859
rect 966 -1893 1002 -1859
rect 916 -1907 1002 -1893
rect 1036 -1893 1052 -1859
rect 1086 -1866 1126 -1859
rect 1036 -1900 1054 -1893
rect 1088 -1900 1126 -1866
rect 1036 -1902 1126 -1900
rect 1252 -1883 1272 -1849
rect 1306 -1883 1402 -1849
rect -36 -1993 298 -1953
rect -36 -2027 -18 -1993
rect 16 -2027 246 -1993
rect 280 -2027 298 -1993
rect -36 -2095 298 -2027
rect -36 -2129 -18 -2095
rect 16 -2129 246 -2095
rect 280 -2129 298 -2095
rect -36 -2171 298 -2129
rect 332 -1973 390 -1938
rect 332 -2007 344 -1973
rect 378 -2007 390 -1973
rect 332 -2066 390 -2007
rect 332 -2100 344 -2066
rect 378 -2100 390 -2066
rect 332 -2171 390 -2100
rect 424 -1982 474 -1934
rect 627 -1943 661 -1909
rect 627 -1977 745 -1943
rect 424 -2019 505 -1982
rect 424 -2053 457 -2019
rect 491 -2053 505 -2019
rect 424 -2087 505 -2053
rect 424 -2121 457 -2087
rect 491 -2121 505 -2087
rect 424 -2137 505 -2121
rect 539 -2020 605 -2011
rect 539 -2054 555 -2020
rect 589 -2054 605 -2020
rect 539 -2088 605 -2054
rect 539 -2122 555 -2088
rect 589 -2122 605 -2088
rect 539 -2171 605 -2122
rect 695 -2019 745 -1977
rect 695 -2053 711 -2019
rect 695 -2087 745 -2053
rect 695 -2121 711 -2087
rect 695 -2137 745 -2121
rect 797 -2020 867 -1908
rect 932 -1936 1002 -1907
rect 932 -1970 1126 -1936
rect 797 -2054 815 -2020
rect 849 -2054 867 -2020
rect 797 -2088 867 -2054
rect 797 -2122 815 -2088
rect 849 -2122 867 -2088
rect 797 -2137 867 -2122
rect 957 -2020 1023 -2004
rect 957 -2054 973 -2020
rect 1007 -2054 1023 -2020
rect 957 -2088 1023 -2054
rect 957 -2122 973 -2088
rect 1007 -2122 1023 -2088
rect 957 -2171 1023 -2122
rect 1057 -2020 1126 -1970
rect 1057 -2054 1073 -2020
rect 1107 -2054 1126 -2020
rect 1057 -2088 1126 -2054
rect 1057 -2122 1073 -2088
rect 1107 -2122 1126 -2088
rect 1057 -2137 1126 -2122
rect 1160 -1973 1218 -1938
rect 1160 -2007 1172 -1973
rect 1206 -2007 1218 -1973
rect 1160 -2066 1218 -2007
rect 1160 -2100 1172 -2066
rect 1206 -2100 1218 -2066
rect 1160 -2171 1218 -2100
rect 1252 -1953 1402 -1883
rect 1436 -1885 1586 -1815
rect 1436 -1919 1532 -1885
rect 1566 -1919 1586 -1885
rect 1712 -1883 1790 -1849
rect 1824 -1883 1893 -1849
rect 1927 -1883 1996 -1849
rect 2030 -1883 2050 -1849
rect 1252 -1993 1586 -1953
rect 1252 -2027 1270 -1993
rect 1304 -2027 1534 -1993
rect 1568 -2027 1586 -1993
rect 1252 -2095 1586 -2027
rect 1252 -2129 1270 -2095
rect 1304 -2129 1534 -2095
rect 1568 -2129 1586 -2095
rect 1252 -2171 1586 -2129
rect 1620 -1973 1678 -1938
rect 1620 -2007 1632 -1973
rect 1666 -2007 1678 -1973
rect 1620 -2066 1678 -2007
rect 1620 -2100 1632 -2066
rect 1666 -2100 1678 -2066
rect 1620 -2171 1678 -2100
rect 1712 -1953 2050 -1883
rect 2084 -1885 2414 -1815
rect 2084 -1919 2104 -1885
rect 2138 -1919 2203 -1885
rect 2237 -1919 2302 -1885
rect 2336 -1919 2414 -1885
rect 2540 -1883 2560 -1849
rect 2594 -1883 2690 -1849
rect 1712 -1993 2414 -1953
rect 1712 -2027 1730 -1993
rect 1764 -2027 2362 -1993
rect 2396 -2027 2414 -1993
rect 1712 -2095 2414 -2027
rect 1712 -2129 1730 -2095
rect 1764 -2129 2362 -2095
rect 2396 -2129 2414 -2095
rect 1712 -2171 2414 -2129
rect 2448 -1973 2506 -1938
rect 2448 -2007 2460 -1973
rect 2494 -2007 2506 -1973
rect 2448 -2066 2506 -2007
rect 2448 -2100 2460 -2066
rect 2494 -2100 2506 -2066
rect 2448 -2171 2506 -2100
rect 2540 -1953 2690 -1883
rect 2724 -1885 2874 -1815
rect 2724 -1919 2820 -1885
rect 2854 -1919 2874 -1885
rect 3000 -1866 3050 -1772
rect 3271 -1790 3321 -1748
rect 3203 -1824 3321 -1790
rect 3373 -1714 3443 -1695
rect 3373 -1748 3392 -1714
rect 3426 -1748 3443 -1714
rect 3203 -1843 3237 -1824
rect 3000 -1900 3014 -1866
rect 3048 -1900 3050 -1866
rect 2540 -1993 2874 -1953
rect 2540 -2027 2558 -1993
rect 2592 -2027 2822 -1993
rect 2856 -2027 2874 -1993
rect 2540 -2095 2874 -2027
rect 2540 -2129 2558 -2095
rect 2592 -2129 2822 -2095
rect 2856 -2129 2874 -2095
rect 2540 -2171 2874 -2129
rect 2908 -1973 2966 -1938
rect 2908 -2007 2920 -1973
rect 2954 -2007 2966 -1973
rect 2908 -2066 2966 -2007
rect 2908 -2100 2920 -2066
rect 2954 -2100 2966 -2066
rect 2908 -2171 2966 -2100
rect 3000 -1982 3050 -1900
rect 3084 -1859 3237 -1843
rect 3373 -1858 3443 -1748
rect 3536 -1714 3602 -1661
rect 3536 -1748 3552 -1714
rect 3586 -1748 3602 -1714
rect 3536 -1757 3602 -1748
rect 3636 -1714 3702 -1695
rect 3636 -1748 3649 -1714
rect 3683 -1748 3702 -1714
rect 3636 -1791 3702 -1748
rect 3508 -1825 3702 -1791
rect 3736 -1755 3794 -1661
rect 3736 -1789 3748 -1755
rect 3782 -1789 3794 -1755
rect 3736 -1806 3794 -1789
rect 3828 -1729 4162 -1661
rect 3828 -1763 3846 -1729
rect 3880 -1763 4110 -1729
rect 4144 -1763 4162 -1729
rect 3828 -1815 4162 -1763
rect 4196 -1755 4254 -1661
rect 4196 -1789 4208 -1755
rect 4242 -1789 4254 -1755
rect 4196 -1806 4254 -1789
rect 4288 -1722 4990 -1661
rect 4288 -1756 4306 -1722
rect 4340 -1756 4938 -1722
rect 4972 -1756 4990 -1722
rect 4288 -1815 4990 -1756
rect 5024 -1755 5082 -1661
rect 5024 -1789 5036 -1755
rect 5070 -1789 5082 -1755
rect 5024 -1806 5082 -1789
rect 5116 -1729 5450 -1661
rect 5116 -1763 5134 -1729
rect 5168 -1763 5398 -1729
rect 5432 -1763 5450 -1729
rect 5116 -1815 5450 -1763
rect 5484 -1755 5542 -1661
rect 5484 -1789 5496 -1755
rect 5530 -1789 5542 -1755
rect 5484 -1806 5542 -1789
rect 5576 -1714 5657 -1695
rect 5576 -1748 5609 -1714
rect 5643 -1748 5657 -1714
rect 5576 -1772 5657 -1748
rect 5691 -1714 5757 -1661
rect 5691 -1748 5707 -1714
rect 5741 -1748 5757 -1714
rect 5691 -1764 5757 -1748
rect 5847 -1714 5897 -1695
rect 5847 -1748 5863 -1714
rect 3508 -1849 3578 -1825
rect 3084 -1893 3087 -1859
rect 3121 -1893 3237 -1859
rect 3084 -1909 3237 -1893
rect 3271 -1859 3443 -1858
rect 3271 -1893 3287 -1859
rect 3321 -1893 3443 -1859
rect 3271 -1908 3443 -1893
rect 3492 -1859 3578 -1849
rect 3492 -1893 3508 -1859
rect 3542 -1893 3578 -1859
rect 3492 -1907 3578 -1893
rect 3612 -1900 3628 -1859
rect 3662 -1900 3702 -1859
rect 3612 -1902 3702 -1900
rect 3828 -1883 3848 -1849
rect 3882 -1883 3978 -1849
rect 3203 -1943 3237 -1909
rect 3203 -1977 3321 -1943
rect 3000 -2019 3081 -1982
rect 3000 -2053 3033 -2019
rect 3067 -2053 3081 -2019
rect 3000 -2087 3081 -2053
rect 3000 -2121 3033 -2087
rect 3067 -2121 3081 -2087
rect 3000 -2137 3081 -2121
rect 3115 -2020 3181 -2011
rect 3115 -2054 3131 -2020
rect 3165 -2054 3181 -2020
rect 3115 -2088 3181 -2054
rect 3115 -2122 3131 -2088
rect 3165 -2122 3181 -2088
rect 3115 -2171 3181 -2122
rect 3271 -2019 3321 -1977
rect 3271 -2053 3287 -2019
rect 3271 -2087 3321 -2053
rect 3271 -2121 3287 -2087
rect 3271 -2137 3321 -2121
rect 3373 -2020 3443 -1908
rect 3508 -1936 3578 -1907
rect 3508 -1970 3702 -1936
rect 3373 -2054 3391 -2020
rect 3425 -2054 3443 -2020
rect 3373 -2088 3443 -2054
rect 3373 -2122 3391 -2088
rect 3425 -2122 3443 -2088
rect 3373 -2137 3443 -2122
rect 3533 -2020 3599 -2004
rect 3533 -2054 3549 -2020
rect 3583 -2054 3599 -2020
rect 3533 -2088 3599 -2054
rect 3533 -2122 3549 -2088
rect 3583 -2122 3599 -2088
rect 3533 -2171 3599 -2122
rect 3633 -2020 3702 -1970
rect 3633 -2054 3649 -2020
rect 3683 -2054 3702 -2020
rect 3633 -2088 3702 -2054
rect 3633 -2122 3649 -2088
rect 3683 -2122 3702 -2088
rect 3633 -2137 3702 -2122
rect 3736 -1973 3794 -1938
rect 3736 -2007 3748 -1973
rect 3782 -2007 3794 -1973
rect 3736 -2066 3794 -2007
rect 3736 -2100 3748 -2066
rect 3782 -2100 3794 -2066
rect 3736 -2171 3794 -2100
rect 3828 -1953 3978 -1883
rect 4012 -1885 4162 -1815
rect 4012 -1919 4108 -1885
rect 4142 -1919 4162 -1885
rect 4288 -1883 4366 -1849
rect 4400 -1883 4469 -1849
rect 4503 -1883 4572 -1849
rect 4606 -1883 4626 -1849
rect 3828 -1993 4162 -1953
rect 3828 -2027 3846 -1993
rect 3880 -2027 4110 -1993
rect 4144 -2027 4162 -1993
rect 3828 -2095 4162 -2027
rect 3828 -2129 3846 -2095
rect 3880 -2129 4110 -2095
rect 4144 -2129 4162 -2095
rect 3828 -2171 4162 -2129
rect 4196 -1973 4254 -1938
rect 4196 -2007 4208 -1973
rect 4242 -2007 4254 -1973
rect 4196 -2066 4254 -2007
rect 4196 -2100 4208 -2066
rect 4242 -2100 4254 -2066
rect 4196 -2171 4254 -2100
rect 4288 -1953 4626 -1883
rect 4660 -1885 4990 -1815
rect 4660 -1919 4680 -1885
rect 4714 -1919 4779 -1885
rect 4813 -1919 4878 -1885
rect 4912 -1919 4990 -1885
rect 5116 -1883 5136 -1849
rect 5170 -1883 5266 -1849
rect 4288 -1993 4990 -1953
rect 4288 -2027 4306 -1993
rect 4340 -2027 4938 -1993
rect 4972 -2027 4990 -1993
rect 4288 -2095 4990 -2027
rect 4288 -2129 4306 -2095
rect 4340 -2129 4938 -2095
rect 4972 -2129 4990 -2095
rect 4288 -2171 4990 -2129
rect 5024 -1973 5082 -1938
rect 5024 -2007 5036 -1973
rect 5070 -2007 5082 -1973
rect 5024 -2066 5082 -2007
rect 5024 -2100 5036 -2066
rect 5070 -2100 5082 -2066
rect 5024 -2171 5082 -2100
rect 5116 -1953 5266 -1883
rect 5300 -1885 5450 -1815
rect 5300 -1919 5396 -1885
rect 5430 -1919 5450 -1885
rect 5576 -1866 5626 -1772
rect 5847 -1790 5897 -1748
rect 5779 -1824 5897 -1790
rect 5949 -1714 6019 -1695
rect 5949 -1748 5968 -1714
rect 6002 -1748 6019 -1714
rect 5779 -1843 5813 -1824
rect 5576 -1900 5588 -1866
rect 5622 -1900 5626 -1866
rect 5116 -1993 5450 -1953
rect 5116 -2027 5134 -1993
rect 5168 -2027 5398 -1993
rect 5432 -2027 5450 -1993
rect 5116 -2095 5450 -2027
rect 5116 -2129 5134 -2095
rect 5168 -2129 5398 -2095
rect 5432 -2129 5450 -2095
rect 5116 -2171 5450 -2129
rect 5484 -1973 5542 -1938
rect 5484 -2007 5496 -1973
rect 5530 -2007 5542 -1973
rect 5484 -2066 5542 -2007
rect 5484 -2100 5496 -2066
rect 5530 -2100 5542 -2066
rect 5484 -2171 5542 -2100
rect 5576 -1982 5626 -1900
rect 5660 -1859 5813 -1843
rect 5949 -1858 6019 -1748
rect 6112 -1714 6178 -1661
rect 6112 -1748 6128 -1714
rect 6162 -1748 6178 -1714
rect 6112 -1757 6178 -1748
rect 6212 -1714 6278 -1695
rect 6212 -1748 6225 -1714
rect 6259 -1748 6278 -1714
rect 6212 -1791 6278 -1748
rect 6084 -1825 6278 -1791
rect 6312 -1755 6370 -1661
rect 6312 -1789 6324 -1755
rect 6358 -1789 6370 -1755
rect 6312 -1806 6370 -1789
rect 6404 -1729 6738 -1661
rect 6404 -1763 6422 -1729
rect 6456 -1763 6686 -1729
rect 6720 -1763 6738 -1729
rect 6404 -1815 6738 -1763
rect 6772 -1755 6830 -1661
rect 6772 -1789 6784 -1755
rect 6818 -1789 6830 -1755
rect 6772 -1806 6830 -1789
rect 6864 -1722 7566 -1661
rect 6864 -1756 6882 -1722
rect 6916 -1756 7514 -1722
rect 7548 -1756 7566 -1722
rect 6864 -1815 7566 -1756
rect 7600 -1755 7658 -1661
rect 7600 -1789 7612 -1755
rect 7646 -1789 7658 -1755
rect 7600 -1806 7658 -1789
rect 7692 -1729 8026 -1661
rect 7692 -1763 7710 -1729
rect 7744 -1763 7974 -1729
rect 8008 -1763 8026 -1729
rect 7692 -1815 8026 -1763
rect 8060 -1755 8118 -1661
rect 8060 -1789 8072 -1755
rect 8106 -1789 8118 -1755
rect 8060 -1806 8118 -1789
rect 8152 -1714 8233 -1695
rect 8152 -1748 8185 -1714
rect 8219 -1748 8233 -1714
rect 8152 -1772 8233 -1748
rect 8267 -1714 8333 -1661
rect 8267 -1748 8283 -1714
rect 8317 -1748 8333 -1714
rect 8267 -1764 8333 -1748
rect 8423 -1714 8473 -1695
rect 8423 -1748 8439 -1714
rect 6084 -1849 6154 -1825
rect 5660 -1893 5663 -1859
rect 5697 -1893 5813 -1859
rect 5660 -1909 5813 -1893
rect 5847 -1859 6019 -1858
rect 5847 -1893 5863 -1859
rect 5897 -1893 6019 -1859
rect 5847 -1908 6019 -1893
rect 6068 -1859 6154 -1849
rect 6068 -1893 6084 -1859
rect 6118 -1893 6154 -1859
rect 6068 -1907 6154 -1893
rect 6188 -1866 6204 -1859
rect 6188 -1900 6202 -1866
rect 6238 -1893 6278 -1859
rect 6236 -1900 6278 -1893
rect 6188 -1902 6278 -1900
rect 6404 -1883 6424 -1849
rect 6458 -1883 6554 -1849
rect 5779 -1943 5813 -1909
rect 5779 -1977 5897 -1943
rect 5576 -2019 5657 -1982
rect 5576 -2053 5609 -2019
rect 5643 -2053 5657 -2019
rect 5576 -2087 5657 -2053
rect 5576 -2121 5609 -2087
rect 5643 -2121 5657 -2087
rect 5576 -2137 5657 -2121
rect 5691 -2020 5757 -2011
rect 5691 -2054 5707 -2020
rect 5741 -2054 5757 -2020
rect 5691 -2088 5757 -2054
rect 5691 -2122 5707 -2088
rect 5741 -2122 5757 -2088
rect 5691 -2171 5757 -2122
rect 5847 -2019 5897 -1977
rect 5847 -2053 5863 -2019
rect 5847 -2087 5897 -2053
rect 5847 -2121 5863 -2087
rect 5847 -2137 5897 -2121
rect 5949 -2020 6019 -1908
rect 6084 -1936 6154 -1907
rect 6084 -1970 6278 -1936
rect 5949 -2054 5967 -2020
rect 6001 -2054 6019 -2020
rect 5949 -2088 6019 -2054
rect 5949 -2122 5967 -2088
rect 6001 -2122 6019 -2088
rect 5949 -2137 6019 -2122
rect 6109 -2020 6175 -2004
rect 6109 -2054 6125 -2020
rect 6159 -2054 6175 -2020
rect 6109 -2088 6175 -2054
rect 6109 -2122 6125 -2088
rect 6159 -2122 6175 -2088
rect 6109 -2171 6175 -2122
rect 6209 -2020 6278 -1970
rect 6209 -2054 6225 -2020
rect 6259 -2054 6278 -2020
rect 6209 -2088 6278 -2054
rect 6209 -2122 6225 -2088
rect 6259 -2122 6278 -2088
rect 6209 -2137 6278 -2122
rect 6312 -1973 6370 -1938
rect 6312 -2007 6324 -1973
rect 6358 -2007 6370 -1973
rect 6312 -2066 6370 -2007
rect 6312 -2100 6324 -2066
rect 6358 -2100 6370 -2066
rect 6312 -2171 6370 -2100
rect 6404 -1953 6554 -1883
rect 6588 -1885 6738 -1815
rect 6588 -1919 6684 -1885
rect 6718 -1919 6738 -1885
rect 6864 -1883 6942 -1849
rect 6976 -1883 7045 -1849
rect 7079 -1883 7148 -1849
rect 7182 -1883 7202 -1849
rect 6404 -1993 6738 -1953
rect 6404 -2027 6422 -1993
rect 6456 -2027 6686 -1993
rect 6720 -2027 6738 -1993
rect 6404 -2095 6738 -2027
rect 6404 -2129 6422 -2095
rect 6456 -2129 6686 -2095
rect 6720 -2129 6738 -2095
rect 6404 -2171 6738 -2129
rect 6772 -1973 6830 -1938
rect 6772 -2007 6784 -1973
rect 6818 -2007 6830 -1973
rect 6772 -2066 6830 -2007
rect 6772 -2100 6784 -2066
rect 6818 -2100 6830 -2066
rect 6772 -2171 6830 -2100
rect 6864 -1953 7202 -1883
rect 7236 -1885 7566 -1815
rect 7236 -1919 7256 -1885
rect 7290 -1919 7355 -1885
rect 7389 -1919 7454 -1885
rect 7488 -1919 7566 -1885
rect 7692 -1883 7712 -1849
rect 7746 -1883 7842 -1849
rect 6864 -1993 7566 -1953
rect 6864 -2027 6882 -1993
rect 6916 -2027 7514 -1993
rect 7548 -2027 7566 -1993
rect 6864 -2095 7566 -2027
rect 6864 -2129 6882 -2095
rect 6916 -2129 7514 -2095
rect 7548 -2129 7566 -2095
rect 6864 -2171 7566 -2129
rect 7600 -1973 7658 -1938
rect 7600 -2007 7612 -1973
rect 7646 -2007 7658 -1973
rect 7600 -2066 7658 -2007
rect 7600 -2100 7612 -2066
rect 7646 -2100 7658 -2066
rect 7600 -2171 7658 -2100
rect 7692 -1953 7842 -1883
rect 7876 -1885 8026 -1815
rect 7876 -1919 7972 -1885
rect 8006 -1919 8026 -1885
rect 8152 -1866 8202 -1772
rect 8423 -1790 8473 -1748
rect 8355 -1824 8473 -1790
rect 8525 -1714 8595 -1695
rect 8525 -1748 8544 -1714
rect 8578 -1748 8595 -1714
rect 8355 -1843 8389 -1824
rect 8152 -1900 8162 -1866
rect 8196 -1900 8202 -1866
rect 7692 -1993 8026 -1953
rect 7692 -2027 7710 -1993
rect 7744 -2027 7974 -1993
rect 8008 -2027 8026 -1993
rect 7692 -2095 8026 -2027
rect 7692 -2129 7710 -2095
rect 7744 -2129 7974 -2095
rect 8008 -2129 8026 -2095
rect 7692 -2171 8026 -2129
rect 8060 -1973 8118 -1938
rect 8060 -2007 8072 -1973
rect 8106 -2007 8118 -1973
rect 8060 -2066 8118 -2007
rect 8060 -2100 8072 -2066
rect 8106 -2100 8118 -2066
rect 8060 -2171 8118 -2100
rect 8152 -1982 8202 -1900
rect 8236 -1859 8389 -1843
rect 8525 -1858 8595 -1748
rect 8688 -1714 8754 -1661
rect 8688 -1748 8704 -1714
rect 8738 -1748 8754 -1714
rect 8688 -1757 8754 -1748
rect 8788 -1714 8854 -1695
rect 8788 -1748 8801 -1714
rect 8835 -1748 8854 -1714
rect 8788 -1791 8854 -1748
rect 8660 -1825 8854 -1791
rect 8888 -1755 8946 -1661
rect 8888 -1789 8900 -1755
rect 8934 -1789 8946 -1755
rect 8888 -1806 8946 -1789
rect 8980 -1729 9314 -1661
rect 8980 -1763 8998 -1729
rect 9032 -1763 9262 -1729
rect 9296 -1763 9314 -1729
rect 8980 -1815 9314 -1763
rect 9348 -1755 9406 -1661
rect 9348 -1789 9360 -1755
rect 9394 -1789 9406 -1755
rect 9348 -1806 9406 -1789
rect 9440 -1722 10142 -1661
rect 9440 -1756 9458 -1722
rect 9492 -1756 10090 -1722
rect 10124 -1756 10142 -1722
rect 9440 -1815 10142 -1756
rect 10176 -1755 10234 -1661
rect 10176 -1789 10188 -1755
rect 10222 -1789 10234 -1755
rect 10176 -1806 10234 -1789
rect 10360 -1729 10694 -1661
rect 10360 -1763 10378 -1729
rect 10412 -1763 10642 -1729
rect 10676 -1763 10694 -1729
rect 10360 -1815 10694 -1763
rect 8660 -1849 8730 -1825
rect 8236 -1893 8239 -1859
rect 8273 -1893 8389 -1859
rect 8236 -1909 8389 -1893
rect 8423 -1859 8595 -1858
rect 8423 -1893 8439 -1859
rect 8473 -1893 8595 -1859
rect 8423 -1908 8595 -1893
rect 8644 -1859 8730 -1849
rect 8644 -1893 8660 -1859
rect 8694 -1893 8730 -1859
rect 8644 -1907 8730 -1893
rect 8764 -1866 8780 -1859
rect 8764 -1900 8776 -1866
rect 8814 -1893 8854 -1859
rect 8810 -1900 8854 -1893
rect 8764 -1902 8854 -1900
rect 8980 -1883 9000 -1849
rect 9034 -1883 9130 -1849
rect 8355 -1943 8389 -1909
rect 8355 -1977 8473 -1943
rect 8152 -2019 8233 -1982
rect 8152 -2053 8185 -2019
rect 8219 -2053 8233 -2019
rect 8152 -2087 8233 -2053
rect 8152 -2121 8185 -2087
rect 8219 -2121 8233 -2087
rect 8152 -2137 8233 -2121
rect 8267 -2020 8333 -2011
rect 8267 -2054 8283 -2020
rect 8317 -2054 8333 -2020
rect 8267 -2088 8333 -2054
rect 8267 -2122 8283 -2088
rect 8317 -2122 8333 -2088
rect 8267 -2171 8333 -2122
rect 8423 -2019 8473 -1977
rect 8423 -2053 8439 -2019
rect 8423 -2087 8473 -2053
rect 8423 -2121 8439 -2087
rect 8423 -2137 8473 -2121
rect 8525 -2020 8595 -1908
rect 8660 -1936 8730 -1907
rect 8660 -1970 8854 -1936
rect 8525 -2054 8543 -2020
rect 8577 -2054 8595 -2020
rect 8525 -2088 8595 -2054
rect 8525 -2122 8543 -2088
rect 8577 -2122 8595 -2088
rect 8525 -2137 8595 -2122
rect 8685 -2020 8751 -2004
rect 8685 -2054 8701 -2020
rect 8735 -2054 8751 -2020
rect 8685 -2088 8751 -2054
rect 8685 -2122 8701 -2088
rect 8735 -2122 8751 -2088
rect 8685 -2171 8751 -2122
rect 8785 -2020 8854 -1970
rect 8785 -2054 8801 -2020
rect 8835 -2054 8854 -2020
rect 8785 -2088 8854 -2054
rect 8785 -2122 8801 -2088
rect 8835 -2122 8854 -2088
rect 8785 -2137 8854 -2122
rect 8888 -1973 8946 -1938
rect 8888 -2007 8900 -1973
rect 8934 -2007 8946 -1973
rect 8888 -2066 8946 -2007
rect 8888 -2100 8900 -2066
rect 8934 -2100 8946 -2066
rect 8888 -2171 8946 -2100
rect 8980 -1953 9130 -1883
rect 9164 -1885 9314 -1815
rect 9164 -1919 9260 -1885
rect 9294 -1919 9314 -1885
rect 9440 -1883 9518 -1849
rect 9552 -1883 9621 -1849
rect 9655 -1883 9724 -1849
rect 9758 -1883 9778 -1849
rect 8980 -1993 9314 -1953
rect 8980 -2027 8998 -1993
rect 9032 -2027 9262 -1993
rect 9296 -2027 9314 -1993
rect 8980 -2095 9314 -2027
rect 8980 -2129 8998 -2095
rect 9032 -2129 9262 -2095
rect 9296 -2129 9314 -2095
rect 8980 -2171 9314 -2129
rect 9348 -1973 9406 -1938
rect 9348 -2007 9360 -1973
rect 9394 -2007 9406 -1973
rect 9348 -2066 9406 -2007
rect 9348 -2100 9360 -2066
rect 9394 -2100 9406 -2066
rect 9348 -2171 9406 -2100
rect 9440 -1953 9778 -1883
rect 9812 -1885 10142 -1815
rect 9812 -1919 9832 -1885
rect 9866 -1919 9931 -1885
rect 9965 -1919 10030 -1885
rect 10064 -1919 10142 -1885
rect 10360 -1883 10380 -1849
rect 10414 -1883 10510 -1849
rect 9440 -1993 10142 -1953
rect 9440 -2027 9458 -1993
rect 9492 -2027 10090 -1993
rect 10124 -2027 10142 -1993
rect 9440 -2095 10142 -2027
rect 9440 -2129 9458 -2095
rect 9492 -2129 10090 -2095
rect 10124 -2129 10142 -2095
rect 9440 -2171 10142 -2129
rect 10176 -1973 10234 -1938
rect 10176 -2007 10188 -1973
rect 10222 -2007 10234 -1973
rect 10176 -2066 10234 -2007
rect 10176 -2100 10188 -2066
rect 10222 -2100 10234 -2066
rect 10176 -2171 10234 -2100
rect 10360 -1953 10510 -1883
rect 10544 -1885 10694 -1815
rect 10544 -1919 10640 -1885
rect 10674 -1919 10694 -1885
rect 10728 -1714 10809 -1695
rect 10728 -1748 10761 -1714
rect 10795 -1748 10809 -1714
rect 10728 -1772 10809 -1748
rect 10843 -1714 10909 -1661
rect 10843 -1748 10859 -1714
rect 10893 -1748 10909 -1714
rect 10843 -1764 10909 -1748
rect 10999 -1714 11049 -1695
rect 10999 -1748 11015 -1714
rect 10728 -1866 10778 -1772
rect 10999 -1790 11049 -1748
rect 10931 -1824 11049 -1790
rect 11101 -1714 11171 -1695
rect 11101 -1748 11120 -1714
rect 11154 -1748 11171 -1714
rect 10931 -1843 10965 -1824
rect 10728 -1900 10736 -1866
rect 10770 -1900 10778 -1866
rect 10360 -1993 10694 -1953
rect 10360 -2027 10378 -1993
rect 10412 -2027 10642 -1993
rect 10676 -2027 10694 -1993
rect 10360 -2095 10694 -2027
rect 10360 -2129 10378 -2095
rect 10412 -2129 10642 -2095
rect 10676 -2129 10694 -2095
rect 10360 -2171 10694 -2129
rect 10728 -1982 10778 -1900
rect 10812 -1859 10965 -1843
rect 11101 -1858 11171 -1748
rect 11264 -1714 11330 -1661
rect 11264 -1748 11280 -1714
rect 11314 -1748 11330 -1714
rect 11264 -1757 11330 -1748
rect 11364 -1714 11430 -1695
rect 11364 -1748 11377 -1714
rect 11411 -1748 11430 -1714
rect 11364 -1791 11430 -1748
rect 11236 -1825 11430 -1791
rect 11464 -1755 11522 -1661
rect 11464 -1789 11476 -1755
rect 11510 -1789 11522 -1755
rect 11464 -1806 11522 -1789
rect 11648 -1729 11982 -1661
rect 11648 -1763 11666 -1729
rect 11700 -1763 11930 -1729
rect 11964 -1763 11982 -1729
rect 11648 -1815 11982 -1763
rect 13580 -1755 13638 -1661
rect 13580 -1789 13592 -1755
rect 13626 -1789 13638 -1755
rect 13672 -1703 13733 -1661
rect 13672 -1737 13690 -1703
rect 13724 -1737 13733 -1703
rect 13672 -1763 13733 -1737
rect 13769 -1716 13819 -1697
rect 13769 -1750 13776 -1716
rect 13810 -1750 13819 -1716
rect 13580 -1806 13638 -1789
rect 11236 -1849 11306 -1825
rect 10812 -1893 10815 -1859
rect 10849 -1893 10965 -1859
rect 10812 -1909 10965 -1893
rect 10999 -1859 11171 -1858
rect 10999 -1893 11015 -1859
rect 11049 -1893 11171 -1859
rect 10999 -1908 11171 -1893
rect 11220 -1859 11306 -1849
rect 11220 -1893 11236 -1859
rect 11270 -1893 11306 -1859
rect 11220 -1907 11306 -1893
rect 11340 -1893 11356 -1859
rect 11390 -1863 11430 -1859
rect 11340 -1897 11386 -1893
rect 11420 -1897 11430 -1863
rect 11340 -1902 11430 -1897
rect 11648 -1883 11668 -1849
rect 11702 -1883 11798 -1849
rect 10931 -1943 10965 -1909
rect 10931 -1977 11049 -1943
rect 10728 -2019 10809 -1982
rect 10728 -2053 10761 -2019
rect 10795 -2053 10809 -2019
rect 10728 -2087 10809 -2053
rect 10728 -2121 10761 -2087
rect 10795 -2121 10809 -2087
rect 10728 -2137 10809 -2121
rect 10843 -2020 10909 -2011
rect 10843 -2054 10859 -2020
rect 10893 -2054 10909 -2020
rect 10843 -2088 10909 -2054
rect 10843 -2122 10859 -2088
rect 10893 -2122 10909 -2088
rect 10843 -2171 10909 -2122
rect 10999 -2019 11049 -1977
rect 10999 -2053 11015 -2019
rect 10999 -2087 11049 -2053
rect 10999 -2121 11015 -2087
rect 10999 -2137 11049 -2121
rect 11101 -2020 11171 -1908
rect 11236 -1936 11306 -1907
rect 11236 -1970 11430 -1936
rect 11101 -2054 11119 -2020
rect 11153 -2054 11171 -2020
rect 11101 -2088 11171 -2054
rect 11101 -2122 11119 -2088
rect 11153 -2122 11171 -2088
rect 11101 -2137 11171 -2122
rect 11261 -2020 11327 -2004
rect 11261 -2054 11277 -2020
rect 11311 -2054 11327 -2020
rect 11261 -2088 11327 -2054
rect 11261 -2122 11277 -2088
rect 11311 -2122 11327 -2088
rect 11261 -2171 11327 -2122
rect 11361 -2020 11430 -1970
rect 11361 -2054 11377 -2020
rect 11411 -2054 11430 -2020
rect 11361 -2088 11430 -2054
rect 11361 -2122 11377 -2088
rect 11411 -2122 11430 -2088
rect 11361 -2137 11430 -2122
rect 11464 -1973 11522 -1938
rect 11464 -2007 11476 -1973
rect 11510 -2007 11522 -1973
rect 11464 -2066 11522 -2007
rect 11464 -2100 11476 -2066
rect 11510 -2100 11522 -2066
rect 11464 -2171 11522 -2100
rect 11648 -1953 11798 -1883
rect 11832 -1885 11982 -1815
rect 11832 -1919 11928 -1885
rect 11962 -1919 11982 -1885
rect 13672 -1832 13735 -1797
rect 13672 -1866 13685 -1832
rect 13719 -1859 13735 -1832
rect 13672 -1893 13692 -1866
rect 13726 -1893 13735 -1859
rect 13672 -1909 13735 -1893
rect 13769 -1859 13819 -1750
rect 13853 -1716 13905 -1661
rect 13853 -1750 13862 -1716
rect 13896 -1750 13905 -1716
rect 13853 -1766 13905 -1750
rect 13941 -1716 13991 -1697
rect 13941 -1750 13948 -1716
rect 13982 -1750 13991 -1716
rect 13941 -1859 13991 -1750
rect 14025 -1716 14077 -1661
rect 14025 -1750 14034 -1716
rect 14068 -1750 14077 -1716
rect 14025 -1773 14077 -1750
rect 14111 -1716 14163 -1700
rect 14111 -1750 14120 -1716
rect 14154 -1750 14163 -1716
rect 14111 -1791 14163 -1750
rect 14197 -1707 14249 -1661
rect 14197 -1741 14206 -1707
rect 14240 -1741 14249 -1707
rect 14197 -1757 14249 -1741
rect 14283 -1716 14335 -1700
rect 14283 -1750 14292 -1716
rect 14326 -1750 14335 -1716
rect 14283 -1791 14335 -1750
rect 14369 -1707 14421 -1661
rect 14369 -1741 14378 -1707
rect 14412 -1741 14421 -1707
rect 14369 -1757 14421 -1741
rect 14455 -1716 14507 -1700
rect 14455 -1750 14464 -1716
rect 14498 -1750 14507 -1716
rect 14455 -1791 14507 -1750
rect 14541 -1707 14590 -1661
rect 14541 -1741 14550 -1707
rect 14584 -1741 14590 -1707
rect 14541 -1757 14590 -1741
rect 14624 -1716 14679 -1700
rect 14624 -1750 14636 -1716
rect 14670 -1750 14679 -1716
rect 14624 -1791 14679 -1750
rect 14713 -1707 14762 -1661
rect 14713 -1741 14722 -1707
rect 14756 -1741 14762 -1707
rect 14713 -1757 14762 -1741
rect 14796 -1716 14848 -1700
rect 14796 -1750 14807 -1716
rect 14841 -1750 14848 -1716
rect 14796 -1791 14848 -1750
rect 14884 -1707 14934 -1661
rect 14884 -1741 14893 -1707
rect 14927 -1741 14934 -1707
rect 14884 -1757 14934 -1741
rect 14968 -1716 15020 -1700
rect 14968 -1750 14979 -1716
rect 15013 -1750 15020 -1716
rect 14968 -1791 15020 -1750
rect 15056 -1707 15106 -1661
rect 15056 -1741 15065 -1707
rect 15099 -1741 15106 -1707
rect 15056 -1757 15106 -1741
rect 15140 -1716 15192 -1700
rect 15140 -1750 15151 -1716
rect 15185 -1750 15192 -1716
rect 15140 -1791 15192 -1750
rect 15228 -1707 15280 -1661
rect 15228 -1741 15237 -1707
rect 15271 -1741 15280 -1707
rect 15228 -1757 15280 -1741
rect 15314 -1716 15366 -1700
rect 15314 -1750 15323 -1716
rect 15357 -1750 15366 -1716
rect 15314 -1791 15366 -1750
rect 15400 -1707 15460 -1661
rect 15400 -1741 15409 -1707
rect 15443 -1741 15460 -1707
rect 15400 -1757 15460 -1741
rect 15512 -1755 15570 -1661
rect 15512 -1789 15524 -1755
rect 15558 -1789 15570 -1755
rect 14111 -1816 15460 -1791
rect 15512 -1806 15570 -1789
rect 15605 -1722 16674 -1661
rect 15605 -1756 15622 -1722
rect 15656 -1756 16622 -1722
rect 16656 -1756 16674 -1722
rect 15605 -1815 16674 -1756
rect 14111 -1825 15248 -1816
rect 15227 -1850 15248 -1825
rect 15282 -1817 15460 -1816
rect 15282 -1850 15340 -1817
rect 15227 -1851 15340 -1850
rect 15374 -1851 15460 -1817
rect 13769 -1893 14119 -1859
rect 14153 -1893 14187 -1859
rect 14221 -1893 14255 -1859
rect 14289 -1893 14323 -1859
rect 14357 -1893 14391 -1859
rect 14425 -1893 14459 -1859
rect 14493 -1893 14527 -1859
rect 14561 -1893 14595 -1859
rect 14629 -1893 14663 -1859
rect 14697 -1893 14731 -1859
rect 14765 -1893 14799 -1859
rect 14833 -1893 14867 -1859
rect 14901 -1893 14935 -1859
rect 14969 -1893 15003 -1859
rect 15037 -1893 15071 -1859
rect 15105 -1893 15139 -1859
rect 15173 -1893 15193 -1859
rect 13769 -1909 15193 -1893
rect 11648 -1993 11982 -1953
rect 11648 -2027 11666 -1993
rect 11700 -2027 11930 -1993
rect 11964 -2027 11982 -1993
rect 11648 -2095 11982 -2027
rect 11648 -2129 11666 -2095
rect 11700 -2129 11930 -2095
rect 11964 -2129 11982 -2095
rect 11648 -2171 11982 -2129
rect 13580 -1973 13638 -1938
rect 13580 -2007 13592 -1973
rect 13626 -2007 13638 -1973
rect 13580 -2066 13638 -2007
rect 13580 -2100 13592 -2066
rect 13626 -2100 13638 -2066
rect 13580 -2171 13638 -2100
rect 13674 -2027 13733 -2009
rect 13674 -2061 13690 -2027
rect 13724 -2061 13733 -2027
rect 13674 -2095 13733 -2061
rect 13674 -2129 13690 -2095
rect 13724 -2129 13733 -2095
rect 13674 -2171 13733 -2129
rect 13769 -2019 13818 -1909
rect 13769 -2053 13776 -2019
rect 13810 -2053 13818 -2019
rect 13769 -2087 13818 -2053
rect 13769 -2121 13776 -2087
rect 13810 -2121 13818 -2087
rect 13769 -2137 13818 -2121
rect 13853 -2027 13905 -2009
rect 13853 -2061 13862 -2027
rect 13896 -2061 13905 -2027
rect 13853 -2095 13905 -2061
rect 13853 -2129 13862 -2095
rect 13896 -2129 13905 -2095
rect 13853 -2171 13905 -2129
rect 13941 -2011 13991 -1909
rect 15227 -1912 15460 -1851
rect 15227 -1943 15248 -1912
rect 14111 -1946 15248 -1943
rect 15282 -1946 15341 -1912
rect 15375 -1946 15460 -1912
rect 15605 -1883 15686 -1849
rect 15720 -1883 15814 -1849
rect 15848 -1883 15942 -1849
rect 15976 -1883 16070 -1849
rect 16104 -1883 16124 -1849
rect 14111 -1965 15460 -1946
rect 14111 -1999 14120 -1965
rect 14154 -1991 14292 -1965
rect 14154 -1999 14163 -1991
rect 13941 -2045 13948 -2011
rect 13982 -2045 13991 -2011
rect 13941 -2079 13991 -2045
rect 13941 -2113 13948 -2079
rect 13982 -2113 13991 -2079
rect 13941 -2136 13991 -2113
rect 14025 -2027 14077 -2011
rect 14025 -2061 14034 -2027
rect 14068 -2061 14077 -2027
rect 14025 -2095 14077 -2061
rect 14025 -2129 14034 -2095
rect 14068 -2129 14077 -2095
rect 14025 -2170 14077 -2129
rect 14111 -2051 14163 -1999
rect 14283 -1999 14292 -1991
rect 14326 -1991 14464 -1965
rect 14326 -1999 14335 -1991
rect 14111 -2085 14120 -2051
rect 14154 -2085 14163 -2051
rect 14111 -2136 14163 -2085
rect 14197 -2071 14249 -2025
rect 14197 -2105 14206 -2071
rect 14240 -2105 14249 -2071
rect 14197 -2170 14249 -2105
rect 14283 -2051 14335 -1999
rect 14455 -1999 14464 -1991
rect 14498 -1991 14636 -1965
rect 14498 -1999 14507 -1991
rect 14283 -2085 14292 -2051
rect 14326 -2085 14335 -2051
rect 14283 -2136 14335 -2085
rect 14369 -2071 14421 -2025
rect 14369 -2105 14378 -2071
rect 14412 -2105 14421 -2071
rect 14369 -2170 14421 -2105
rect 14455 -2051 14507 -1999
rect 14627 -1999 14636 -1991
rect 14670 -1991 14807 -1965
rect 14670 -1999 14679 -1991
rect 14455 -2085 14464 -2051
rect 14498 -2085 14507 -2051
rect 14455 -2136 14507 -2085
rect 14541 -2071 14593 -2025
rect 14541 -2105 14550 -2071
rect 14584 -2105 14593 -2071
rect 14541 -2170 14593 -2105
rect 14627 -2051 14679 -1999
rect 14796 -1999 14807 -1991
rect 14841 -1991 14979 -1965
rect 14841 -1999 14848 -1991
rect 14627 -2085 14636 -2051
rect 14670 -2085 14679 -2051
rect 14627 -2136 14679 -2085
rect 14713 -2071 14762 -2025
rect 14713 -2105 14722 -2071
rect 14756 -2105 14762 -2071
rect 14713 -2170 14762 -2105
rect 14796 -2051 14848 -1999
rect 14968 -1999 14979 -1991
rect 15013 -1991 15151 -1965
rect 15013 -1999 15020 -1991
rect 14796 -2085 14807 -2051
rect 14841 -2085 14848 -2051
rect 14796 -2136 14848 -2085
rect 14885 -2071 14934 -2025
rect 14885 -2105 14893 -2071
rect 14927 -2105 14934 -2071
rect 14885 -2170 14934 -2105
rect 14968 -2051 15020 -1999
rect 15140 -1999 15151 -1991
rect 15185 -1988 15323 -1965
rect 15185 -1999 15192 -1988
rect 14968 -2085 14979 -2051
rect 15013 -2085 15020 -2051
rect 14968 -2136 15020 -2085
rect 15057 -2071 15106 -2025
rect 15057 -2105 15065 -2071
rect 15099 -2105 15106 -2071
rect 15057 -2170 15106 -2105
rect 15140 -2051 15192 -1999
rect 15314 -1999 15323 -1988
rect 15357 -1988 15460 -1965
rect 15512 -1973 15570 -1938
rect 15357 -1999 15372 -1988
rect 15140 -2085 15151 -2051
rect 15185 -2085 15192 -2051
rect 15140 -2136 15192 -2085
rect 15229 -2071 15280 -2025
rect 15229 -2105 15237 -2071
rect 15271 -2105 15280 -2071
rect 15229 -2170 15280 -2105
rect 15314 -2051 15372 -1999
rect 15512 -2007 15524 -1973
rect 15558 -2007 15570 -1973
rect 15314 -2085 15323 -2051
rect 15357 -2085 15372 -2051
rect 15314 -2136 15372 -2085
rect 15406 -2071 15460 -2022
rect 15406 -2105 15409 -2071
rect 15443 -2105 15460 -2071
rect 14025 -2171 15280 -2170
rect 15406 -2171 15460 -2105
rect 15512 -2066 15570 -2007
rect 15512 -2100 15524 -2066
rect 15558 -2100 15570 -2066
rect 15512 -2171 15570 -2100
rect 15605 -1953 16124 -1883
rect 16158 -1885 16674 -1815
rect 16158 -1919 16178 -1885
rect 16212 -1919 16306 -1885
rect 16340 -1919 16434 -1885
rect 16468 -1919 16562 -1885
rect 16596 -1919 16674 -1885
rect 15605 -1993 16674 -1953
rect 15605 -2027 15622 -1993
rect 15656 -2027 16622 -1993
rect 16656 -2027 16674 -1993
rect 15605 -2095 16674 -2027
rect 15605 -2129 15622 -2095
rect 15656 -2129 16622 -2095
rect 16656 -2129 16674 -2095
rect 15605 -2171 16674 -2129
rect -2997 -2205 -2968 -2171
rect -2934 -2205 -2876 -2171
rect -2842 -2205 -2784 -2171
rect -2750 -2205 -2692 -2171
rect -2658 -2205 -2600 -2171
rect -2566 -2205 -2508 -2171
rect -2474 -2205 -2416 -2171
rect -2382 -2205 -2324 -2171
rect -2290 -2205 -2232 -2171
rect -2198 -2205 -2140 -2171
rect -2106 -2205 -2048 -2171
rect -2014 -2205 -1956 -2171
rect -1922 -2205 -1864 -2171
rect -1830 -2205 -1772 -2171
rect -1738 -2205 -1680 -2171
rect -1646 -2205 -1588 -2171
rect -1554 -2205 -1496 -2171
rect -1462 -2205 -1404 -2171
rect -1370 -2205 -1312 -2171
rect -1278 -2205 -1220 -2171
rect -1186 -2205 -1128 -2171
rect -1094 -2205 -1036 -2171
rect -1002 -2205 -944 -2171
rect -910 -2205 -852 -2171
rect -818 -2205 -760 -2171
rect -726 -2205 -668 -2171
rect -634 -2205 -576 -2171
rect -542 -2205 -484 -2171
rect -450 -2205 -392 -2171
rect -358 -2205 -300 -2171
rect -266 -2205 -208 -2171
rect -174 -2205 -116 -2171
rect -82 -2205 -24 -2171
rect 10 -2205 68 -2171
rect 102 -2205 160 -2171
rect 194 -2205 252 -2171
rect 286 -2205 344 -2171
rect 378 -2205 436 -2171
rect 470 -2205 528 -2171
rect 562 -2205 620 -2171
rect 654 -2205 712 -2171
rect 746 -2205 804 -2171
rect 838 -2205 896 -2171
rect 930 -2205 988 -2171
rect 1022 -2205 1080 -2171
rect 1114 -2205 1172 -2171
rect 1206 -2205 1264 -2171
rect 1298 -2205 1356 -2171
rect 1390 -2205 1448 -2171
rect 1482 -2205 1540 -2171
rect 1574 -2205 1632 -2171
rect 1666 -2205 1724 -2171
rect 1758 -2205 1816 -2171
rect 1850 -2205 1908 -2171
rect 1942 -2205 2000 -2171
rect 2034 -2205 2092 -2171
rect 2126 -2205 2184 -2171
rect 2218 -2205 2276 -2171
rect 2310 -2205 2368 -2171
rect 2402 -2205 2460 -2171
rect 2494 -2205 2552 -2171
rect 2586 -2205 2644 -2171
rect 2678 -2205 2736 -2171
rect 2770 -2205 2828 -2171
rect 2862 -2205 2920 -2171
rect 2954 -2205 3012 -2171
rect 3046 -2205 3104 -2171
rect 3138 -2205 3196 -2171
rect 3230 -2205 3288 -2171
rect 3322 -2205 3380 -2171
rect 3414 -2205 3472 -2171
rect 3506 -2205 3564 -2171
rect 3598 -2205 3656 -2171
rect 3690 -2205 3748 -2171
rect 3782 -2205 3840 -2171
rect 3874 -2205 3932 -2171
rect 3966 -2205 4024 -2171
rect 4058 -2205 4116 -2171
rect 4150 -2205 4208 -2171
rect 4242 -2205 4300 -2171
rect 4334 -2205 4392 -2171
rect 4426 -2205 4484 -2171
rect 4518 -2205 4576 -2171
rect 4610 -2205 4668 -2171
rect 4702 -2205 4760 -2171
rect 4794 -2205 4852 -2171
rect 4886 -2205 4944 -2171
rect 4978 -2205 5036 -2171
rect 5070 -2205 5128 -2171
rect 5162 -2205 5220 -2171
rect 5254 -2205 5312 -2171
rect 5346 -2205 5404 -2171
rect 5438 -2205 5496 -2171
rect 5530 -2205 5588 -2171
rect 5622 -2205 5680 -2171
rect 5714 -2205 5772 -2171
rect 5806 -2205 5864 -2171
rect 5898 -2205 5956 -2171
rect 5990 -2205 6048 -2171
rect 6082 -2205 6140 -2171
rect 6174 -2205 6232 -2171
rect 6266 -2205 6324 -2171
rect 6358 -2205 6416 -2171
rect 6450 -2205 6508 -2171
rect 6542 -2205 6600 -2171
rect 6634 -2205 6692 -2171
rect 6726 -2205 6784 -2171
rect 6818 -2205 6876 -2171
rect 6910 -2205 6968 -2171
rect 7002 -2205 7060 -2171
rect 7094 -2205 7152 -2171
rect 7186 -2205 7244 -2171
rect 7278 -2205 7336 -2171
rect 7370 -2205 7428 -2171
rect 7462 -2205 7520 -2171
rect 7554 -2205 7612 -2171
rect 7646 -2205 7704 -2171
rect 7738 -2205 7796 -2171
rect 7830 -2205 7888 -2171
rect 7922 -2205 7980 -2171
rect 8014 -2205 8072 -2171
rect 8106 -2205 8164 -2171
rect 8198 -2205 8256 -2171
rect 8290 -2205 8348 -2171
rect 8382 -2205 8440 -2171
rect 8474 -2205 8532 -2171
rect 8566 -2205 8624 -2171
rect 8658 -2205 8716 -2171
rect 8750 -2205 8808 -2171
rect 8842 -2205 8900 -2171
rect 8934 -2205 8992 -2171
rect 9026 -2205 9084 -2171
rect 9118 -2205 9176 -2171
rect 9210 -2205 9268 -2171
rect 9302 -2205 9360 -2171
rect 9394 -2205 9452 -2171
rect 9486 -2205 9544 -2171
rect 9578 -2205 9636 -2171
rect 9670 -2205 9728 -2171
rect 9762 -2205 9820 -2171
rect 9854 -2205 9912 -2171
rect 9946 -2205 10004 -2171
rect 10038 -2205 10096 -2171
rect 10130 -2205 10188 -2171
rect 10222 -2205 10280 -2171
rect 10314 -2205 10372 -2171
rect 10406 -2205 10464 -2171
rect 10498 -2205 10556 -2171
rect 10590 -2205 10648 -2171
rect 10682 -2205 10740 -2171
rect 10774 -2205 10832 -2171
rect 10866 -2205 10924 -2171
rect 10958 -2205 11016 -2171
rect 11050 -2205 11108 -2171
rect 11142 -2205 11200 -2171
rect 11234 -2205 11292 -2171
rect 11326 -2205 11384 -2171
rect 11418 -2205 11476 -2171
rect 11510 -2205 11568 -2171
rect 11602 -2205 11660 -2171
rect 11694 -2205 11752 -2171
rect 11786 -2205 11844 -2171
rect 11878 -2205 11936 -2171
rect 11970 -2205 12028 -2171
rect 12062 -2205 12120 -2171
rect 12154 -2205 12212 -2171
rect 12246 -2205 12304 -2171
rect 12338 -2205 12396 -2171
rect 12430 -2205 12488 -2171
rect 12522 -2205 12580 -2171
rect 12614 -2205 12672 -2171
rect 12706 -2205 12764 -2171
rect 12798 -2205 12856 -2171
rect 12890 -2205 12948 -2171
rect 12982 -2205 13040 -2171
rect 13074 -2205 13132 -2171
rect 13166 -2205 13224 -2171
rect 13258 -2205 13316 -2171
rect 13350 -2205 13408 -2171
rect 13442 -2205 13500 -2171
rect 13534 -2205 13592 -2171
rect 13626 -2205 13684 -2171
rect 13718 -2205 13776 -2171
rect 13810 -2205 13868 -2171
rect 13902 -2205 13960 -2171
rect 13994 -2205 14052 -2171
rect 14086 -2205 14144 -2171
rect 14178 -2205 14236 -2171
rect 14270 -2205 14328 -2171
rect 14362 -2205 14420 -2171
rect 14454 -2205 14512 -2171
rect 14546 -2205 14604 -2171
rect 14638 -2205 14696 -2171
rect 14730 -2205 14788 -2171
rect 14822 -2205 14880 -2171
rect 14914 -2205 14972 -2171
rect 15006 -2205 15064 -2171
rect 15098 -2205 15156 -2171
rect 15190 -2205 15248 -2171
rect 15282 -2205 15340 -2171
rect 15374 -2205 15432 -2171
rect 15466 -2205 15524 -2171
rect 15558 -2205 15616 -2171
rect 15650 -2205 15708 -2171
rect 15742 -2205 15800 -2171
rect 15834 -2205 15892 -2171
rect 15926 -2205 15984 -2171
rect 16018 -2205 16076 -2171
rect 16110 -2205 16168 -2171
rect 16202 -2205 16260 -2171
rect 16294 -2205 16352 -2171
rect 16386 -2205 16444 -2171
rect 16478 -2205 16536 -2171
rect 16570 -2205 16628 -2171
rect 16662 -2205 16691 -2171
rect -2980 -2247 -2278 -2205
rect -2980 -2281 -2962 -2247
rect -2928 -2281 -2330 -2247
rect -2296 -2281 -2278 -2247
rect -2980 -2349 -2278 -2281
rect -2980 -2383 -2962 -2349
rect -2928 -2383 -2330 -2349
rect -2296 -2383 -2278 -2349
rect -2980 -2423 -2278 -2383
rect -2980 -2491 -2902 -2457
rect -2868 -2491 -2803 -2457
rect -2769 -2491 -2704 -2457
rect -2670 -2491 -2650 -2457
rect -2980 -2561 -2650 -2491
rect -2616 -2493 -2278 -2423
rect -2244 -2276 -2186 -2205
rect -2244 -2310 -2232 -2276
rect -2198 -2310 -2186 -2276
rect -2244 -2369 -2186 -2310
rect -2244 -2403 -2232 -2369
rect -2198 -2403 -2186 -2369
rect -2244 -2438 -2186 -2403
rect -1600 -2247 -898 -2205
rect -1600 -2281 -1582 -2247
rect -1548 -2281 -950 -2247
rect -916 -2281 -898 -2247
rect -1600 -2349 -898 -2281
rect -1600 -2383 -1582 -2349
rect -1548 -2383 -950 -2349
rect -916 -2383 -898 -2349
rect -1600 -2423 -898 -2383
rect -864 -2247 -162 -2205
rect -864 -2281 -846 -2247
rect -812 -2281 -214 -2247
rect -180 -2281 -162 -2247
rect -864 -2349 -162 -2281
rect -864 -2383 -846 -2349
rect -812 -2383 -214 -2349
rect -180 -2383 -162 -2349
rect -864 -2423 -162 -2383
rect -2616 -2527 -2596 -2493
rect -2562 -2527 -2493 -2493
rect -2459 -2527 -2390 -2493
rect -2356 -2527 -2278 -2493
rect -1600 -2491 -1522 -2457
rect -1488 -2491 -1423 -2457
rect -1389 -2491 -1324 -2457
rect -1290 -2491 -1270 -2457
rect -1600 -2561 -1270 -2491
rect -1236 -2493 -898 -2423
rect -1236 -2527 -1216 -2493
rect -1182 -2527 -1113 -2493
rect -1079 -2527 -1010 -2493
rect -976 -2527 -898 -2493
rect -864 -2491 -786 -2457
rect -752 -2491 -687 -2457
rect -653 -2491 -588 -2457
rect -554 -2491 -534 -2457
rect -864 -2561 -534 -2491
rect -500 -2493 -162 -2423
rect -128 -2276 -70 -2205
rect -128 -2310 -116 -2276
rect -82 -2310 -70 -2276
rect -128 -2369 -70 -2310
rect -128 -2403 -116 -2369
rect -82 -2403 -70 -2369
rect -128 -2438 -70 -2403
rect -36 -2247 298 -2205
rect -36 -2281 -18 -2247
rect 16 -2281 246 -2247
rect 280 -2281 298 -2247
rect -36 -2349 298 -2281
rect -36 -2383 -18 -2349
rect 16 -2383 246 -2349
rect 280 -2383 298 -2349
rect -36 -2423 298 -2383
rect 332 -2276 390 -2205
rect 332 -2310 344 -2276
rect 378 -2310 390 -2276
rect 332 -2369 390 -2310
rect 332 -2403 344 -2369
rect 378 -2403 390 -2369
rect -500 -2527 -480 -2493
rect -446 -2527 -377 -2493
rect -343 -2527 -274 -2493
rect -240 -2527 -162 -2493
rect -36 -2493 114 -2423
rect 332 -2438 390 -2403
rect 424 -2254 493 -2239
rect 424 -2288 443 -2254
rect 477 -2288 493 -2254
rect 424 -2322 493 -2288
rect 424 -2356 443 -2322
rect 477 -2356 493 -2322
rect 424 -2406 493 -2356
rect 527 -2254 593 -2205
rect 527 -2288 543 -2254
rect 577 -2288 593 -2254
rect 527 -2322 593 -2288
rect 527 -2356 543 -2322
rect 577 -2356 593 -2322
rect 527 -2372 593 -2356
rect 683 -2254 753 -2239
rect 683 -2288 701 -2254
rect 735 -2288 753 -2254
rect 683 -2322 753 -2288
rect 683 -2356 701 -2322
rect 735 -2356 753 -2322
rect 424 -2440 618 -2406
rect -36 -2527 -16 -2493
rect 18 -2527 114 -2493
rect 148 -2491 244 -2457
rect 278 -2491 298 -2457
rect 548 -2469 618 -2440
rect 683 -2468 753 -2356
rect 805 -2255 855 -2239
rect 839 -2289 855 -2255
rect 805 -2323 855 -2289
rect 839 -2357 855 -2323
rect 805 -2399 855 -2357
rect 945 -2254 1011 -2205
rect 945 -2288 961 -2254
rect 995 -2288 1011 -2254
rect 945 -2322 1011 -2288
rect 945 -2356 961 -2322
rect 995 -2356 1011 -2322
rect 945 -2365 1011 -2356
rect 1045 -2255 1126 -2239
rect 1045 -2289 1059 -2255
rect 1093 -2289 1126 -2255
rect 1045 -2323 1126 -2289
rect 1045 -2357 1059 -2323
rect 1093 -2357 1126 -2323
rect 1045 -2394 1126 -2357
rect 805 -2433 923 -2399
rect 889 -2467 923 -2433
rect 148 -2561 298 -2491
rect 424 -2480 514 -2474
rect 424 -2514 436 -2480
rect 470 -2483 514 -2480
rect 424 -2517 464 -2514
rect 498 -2517 514 -2483
rect 548 -2483 634 -2469
rect 548 -2517 584 -2483
rect 618 -2517 634 -2483
rect 548 -2527 634 -2517
rect 683 -2483 855 -2468
rect 683 -2517 805 -2483
rect 839 -2517 855 -2483
rect 683 -2518 855 -2517
rect 889 -2483 1042 -2467
rect 889 -2517 1005 -2483
rect 1039 -2517 1042 -2483
rect 548 -2551 618 -2527
rect -2980 -2620 -2278 -2561
rect -2980 -2654 -2962 -2620
rect -2928 -2654 -2330 -2620
rect -2296 -2654 -2278 -2620
rect -2980 -2715 -2278 -2654
rect -2244 -2587 -2186 -2570
rect -2244 -2621 -2232 -2587
rect -2198 -2621 -2186 -2587
rect -2244 -2715 -2186 -2621
rect -1600 -2620 -898 -2561
rect -1600 -2654 -1582 -2620
rect -1548 -2654 -950 -2620
rect -916 -2654 -898 -2620
rect -1600 -2715 -898 -2654
rect -864 -2620 -162 -2561
rect -864 -2654 -846 -2620
rect -812 -2654 -214 -2620
rect -180 -2654 -162 -2620
rect -864 -2715 -162 -2654
rect -128 -2587 -70 -2570
rect -128 -2621 -116 -2587
rect -82 -2621 -70 -2587
rect -128 -2715 -70 -2621
rect -36 -2613 298 -2561
rect -36 -2647 -18 -2613
rect 16 -2647 246 -2613
rect 280 -2647 298 -2613
rect -36 -2715 298 -2647
rect 332 -2587 390 -2570
rect 332 -2621 344 -2587
rect 378 -2621 390 -2587
rect 332 -2715 390 -2621
rect 424 -2585 618 -2551
rect 424 -2628 490 -2585
rect 424 -2662 443 -2628
rect 477 -2662 490 -2628
rect 424 -2681 490 -2662
rect 524 -2628 590 -2619
rect 524 -2662 540 -2628
rect 574 -2662 590 -2628
rect 524 -2715 590 -2662
rect 683 -2628 753 -2518
rect 889 -2533 1042 -2517
rect 1076 -2478 1126 -2394
rect 1160 -2276 1218 -2205
rect 1160 -2310 1172 -2276
rect 1206 -2310 1218 -2276
rect 1160 -2369 1218 -2310
rect 1160 -2403 1172 -2369
rect 1206 -2403 1218 -2369
rect 1160 -2438 1218 -2403
rect 1252 -2247 1586 -2205
rect 1252 -2281 1270 -2247
rect 1304 -2281 1534 -2247
rect 1568 -2281 1586 -2247
rect 1252 -2349 1586 -2281
rect 1252 -2383 1270 -2349
rect 1304 -2383 1534 -2349
rect 1568 -2383 1586 -2349
rect 1252 -2423 1586 -2383
rect 1620 -2276 1678 -2205
rect 1620 -2310 1632 -2276
rect 1666 -2310 1678 -2276
rect 1620 -2369 1678 -2310
rect 1620 -2403 1632 -2369
rect 1666 -2403 1678 -2369
rect 1076 -2512 1081 -2478
rect 1115 -2512 1126 -2478
rect 889 -2552 923 -2533
rect 683 -2662 700 -2628
rect 734 -2662 753 -2628
rect 683 -2681 753 -2662
rect 805 -2586 923 -2552
rect 805 -2628 855 -2586
rect 1076 -2604 1126 -2512
rect 1252 -2493 1402 -2423
rect 1620 -2438 1678 -2403
rect 1712 -2247 2414 -2205
rect 1712 -2281 1730 -2247
rect 1764 -2281 2362 -2247
rect 2396 -2281 2414 -2247
rect 1712 -2349 2414 -2281
rect 1712 -2383 1730 -2349
rect 1764 -2383 2362 -2349
rect 2396 -2383 2414 -2349
rect 1712 -2423 2414 -2383
rect 1252 -2527 1272 -2493
rect 1306 -2527 1402 -2493
rect 1436 -2491 1532 -2457
rect 1566 -2491 1586 -2457
rect 1436 -2561 1586 -2491
rect 839 -2662 855 -2628
rect 805 -2681 855 -2662
rect 945 -2628 1011 -2612
rect 945 -2662 961 -2628
rect 995 -2662 1011 -2628
rect 945 -2715 1011 -2662
rect 1045 -2628 1126 -2604
rect 1045 -2662 1059 -2628
rect 1093 -2662 1126 -2628
rect 1045 -2681 1126 -2662
rect 1160 -2587 1218 -2570
rect 1160 -2621 1172 -2587
rect 1206 -2621 1218 -2587
rect 1160 -2715 1218 -2621
rect 1252 -2613 1586 -2561
rect 1712 -2491 1790 -2457
rect 1824 -2491 1889 -2457
rect 1923 -2491 1988 -2457
rect 2022 -2491 2042 -2457
rect 1712 -2561 2042 -2491
rect 2076 -2493 2414 -2423
rect 2448 -2276 2506 -2205
rect 2448 -2310 2460 -2276
rect 2494 -2310 2506 -2276
rect 2448 -2369 2506 -2310
rect 2448 -2403 2460 -2369
rect 2494 -2403 2506 -2369
rect 2448 -2438 2506 -2403
rect 2540 -2247 2874 -2205
rect 2540 -2281 2558 -2247
rect 2592 -2281 2822 -2247
rect 2856 -2281 2874 -2247
rect 2540 -2349 2874 -2281
rect 2540 -2383 2558 -2349
rect 2592 -2383 2822 -2349
rect 2856 -2383 2874 -2349
rect 2540 -2423 2874 -2383
rect 2908 -2276 2966 -2205
rect 2908 -2310 2920 -2276
rect 2954 -2310 2966 -2276
rect 2908 -2369 2966 -2310
rect 2908 -2403 2920 -2369
rect 2954 -2403 2966 -2369
rect 2076 -2527 2096 -2493
rect 2130 -2527 2199 -2493
rect 2233 -2527 2302 -2493
rect 2336 -2527 2414 -2493
rect 2540 -2493 2690 -2423
rect 2908 -2438 2966 -2403
rect 3000 -2254 3069 -2239
rect 3000 -2288 3019 -2254
rect 3053 -2288 3069 -2254
rect 3000 -2322 3069 -2288
rect 3000 -2356 3019 -2322
rect 3053 -2356 3069 -2322
rect 3000 -2406 3069 -2356
rect 3103 -2254 3169 -2205
rect 3103 -2288 3119 -2254
rect 3153 -2288 3169 -2254
rect 3103 -2322 3169 -2288
rect 3103 -2356 3119 -2322
rect 3153 -2356 3169 -2322
rect 3103 -2372 3169 -2356
rect 3259 -2254 3329 -2239
rect 3259 -2288 3277 -2254
rect 3311 -2288 3329 -2254
rect 3259 -2322 3329 -2288
rect 3259 -2356 3277 -2322
rect 3311 -2356 3329 -2322
rect 3000 -2440 3194 -2406
rect 2540 -2527 2560 -2493
rect 2594 -2527 2690 -2493
rect 2724 -2491 2820 -2457
rect 2854 -2491 2874 -2457
rect 3124 -2469 3194 -2440
rect 3259 -2468 3329 -2356
rect 3381 -2255 3431 -2239
rect 3415 -2289 3431 -2255
rect 3381 -2323 3431 -2289
rect 3415 -2357 3431 -2323
rect 3381 -2399 3431 -2357
rect 3521 -2254 3587 -2205
rect 3521 -2288 3537 -2254
rect 3571 -2288 3587 -2254
rect 3521 -2322 3587 -2288
rect 3521 -2356 3537 -2322
rect 3571 -2356 3587 -2322
rect 3521 -2365 3587 -2356
rect 3621 -2255 3702 -2239
rect 3621 -2289 3635 -2255
rect 3669 -2289 3702 -2255
rect 3621 -2323 3702 -2289
rect 3621 -2357 3635 -2323
rect 3669 -2357 3702 -2323
rect 3621 -2394 3702 -2357
rect 3381 -2433 3499 -2399
rect 3465 -2467 3499 -2433
rect 2724 -2561 2874 -2491
rect 3000 -2478 3090 -2474
rect 3000 -2483 3041 -2478
rect 3000 -2517 3040 -2483
rect 3075 -2512 3090 -2478
rect 3074 -2517 3090 -2512
rect 3124 -2483 3210 -2469
rect 3124 -2517 3160 -2483
rect 3194 -2517 3210 -2483
rect 3124 -2527 3210 -2517
rect 3259 -2483 3431 -2468
rect 3259 -2517 3381 -2483
rect 3415 -2517 3431 -2483
rect 3259 -2518 3431 -2517
rect 3465 -2483 3618 -2467
rect 3465 -2517 3581 -2483
rect 3615 -2517 3618 -2483
rect 3124 -2551 3194 -2527
rect 1252 -2647 1270 -2613
rect 1304 -2647 1534 -2613
rect 1568 -2647 1586 -2613
rect 1252 -2715 1586 -2647
rect 1620 -2587 1678 -2570
rect 1620 -2621 1632 -2587
rect 1666 -2621 1678 -2587
rect 1620 -2715 1678 -2621
rect 1712 -2620 2414 -2561
rect 1712 -2654 1730 -2620
rect 1764 -2654 2362 -2620
rect 2396 -2654 2414 -2620
rect 1712 -2715 2414 -2654
rect 2448 -2587 2506 -2570
rect 2448 -2621 2460 -2587
rect 2494 -2621 2506 -2587
rect 2448 -2715 2506 -2621
rect 2540 -2613 2874 -2561
rect 2540 -2647 2558 -2613
rect 2592 -2647 2822 -2613
rect 2856 -2647 2874 -2613
rect 2540 -2715 2874 -2647
rect 2908 -2587 2966 -2570
rect 2908 -2621 2920 -2587
rect 2954 -2621 2966 -2587
rect 2908 -2715 2966 -2621
rect 3000 -2585 3194 -2551
rect 3000 -2628 3066 -2585
rect 3000 -2662 3019 -2628
rect 3053 -2662 3066 -2628
rect 3000 -2681 3066 -2662
rect 3100 -2628 3166 -2619
rect 3100 -2662 3116 -2628
rect 3150 -2662 3166 -2628
rect 3100 -2715 3166 -2662
rect 3259 -2628 3329 -2518
rect 3465 -2533 3618 -2517
rect 3652 -2478 3702 -2394
rect 3736 -2276 3794 -2205
rect 3736 -2310 3748 -2276
rect 3782 -2310 3794 -2276
rect 3736 -2369 3794 -2310
rect 3736 -2403 3748 -2369
rect 3782 -2403 3794 -2369
rect 3736 -2438 3794 -2403
rect 3828 -2247 4162 -2205
rect 3828 -2281 3846 -2247
rect 3880 -2281 4110 -2247
rect 4144 -2281 4162 -2247
rect 3828 -2349 4162 -2281
rect 3828 -2383 3846 -2349
rect 3880 -2383 4110 -2349
rect 4144 -2383 4162 -2349
rect 3828 -2423 4162 -2383
rect 4196 -2276 4254 -2205
rect 4196 -2310 4208 -2276
rect 4242 -2310 4254 -2276
rect 4196 -2369 4254 -2310
rect 4196 -2403 4208 -2369
rect 4242 -2403 4254 -2369
rect 3652 -2512 3655 -2478
rect 3689 -2512 3702 -2478
rect 3465 -2552 3499 -2533
rect 3259 -2662 3276 -2628
rect 3310 -2662 3329 -2628
rect 3259 -2681 3329 -2662
rect 3381 -2586 3499 -2552
rect 3381 -2628 3431 -2586
rect 3652 -2604 3702 -2512
rect 3828 -2493 3978 -2423
rect 4196 -2438 4254 -2403
rect 4288 -2247 4990 -2205
rect 4288 -2281 4306 -2247
rect 4340 -2281 4938 -2247
rect 4972 -2281 4990 -2247
rect 4288 -2349 4990 -2281
rect 4288 -2383 4306 -2349
rect 4340 -2383 4938 -2349
rect 4972 -2383 4990 -2349
rect 4288 -2423 4990 -2383
rect 3828 -2527 3848 -2493
rect 3882 -2527 3978 -2493
rect 4012 -2491 4108 -2457
rect 4142 -2491 4162 -2457
rect 4012 -2561 4162 -2491
rect 3415 -2662 3431 -2628
rect 3381 -2681 3431 -2662
rect 3521 -2628 3587 -2612
rect 3521 -2662 3537 -2628
rect 3571 -2662 3587 -2628
rect 3521 -2715 3587 -2662
rect 3621 -2628 3702 -2604
rect 3621 -2662 3635 -2628
rect 3669 -2662 3702 -2628
rect 3621 -2681 3702 -2662
rect 3736 -2587 3794 -2570
rect 3736 -2621 3748 -2587
rect 3782 -2621 3794 -2587
rect 3736 -2715 3794 -2621
rect 3828 -2613 4162 -2561
rect 4288 -2491 4366 -2457
rect 4400 -2491 4465 -2457
rect 4499 -2491 4564 -2457
rect 4598 -2491 4618 -2457
rect 4288 -2561 4618 -2491
rect 4652 -2493 4990 -2423
rect 5024 -2276 5082 -2205
rect 5024 -2310 5036 -2276
rect 5070 -2310 5082 -2276
rect 5024 -2369 5082 -2310
rect 5024 -2403 5036 -2369
rect 5070 -2403 5082 -2369
rect 5024 -2438 5082 -2403
rect 5116 -2247 5450 -2205
rect 5116 -2281 5134 -2247
rect 5168 -2281 5398 -2247
rect 5432 -2281 5450 -2247
rect 5116 -2349 5450 -2281
rect 5116 -2383 5134 -2349
rect 5168 -2383 5398 -2349
rect 5432 -2383 5450 -2349
rect 5116 -2423 5450 -2383
rect 5484 -2276 5542 -2205
rect 5484 -2310 5496 -2276
rect 5530 -2310 5542 -2276
rect 5484 -2369 5542 -2310
rect 5484 -2403 5496 -2369
rect 5530 -2403 5542 -2369
rect 4652 -2527 4672 -2493
rect 4706 -2527 4775 -2493
rect 4809 -2527 4878 -2493
rect 4912 -2527 4990 -2493
rect 5116 -2493 5266 -2423
rect 5484 -2438 5542 -2403
rect 5576 -2254 5645 -2239
rect 5576 -2288 5595 -2254
rect 5629 -2288 5645 -2254
rect 5576 -2322 5645 -2288
rect 5576 -2356 5595 -2322
rect 5629 -2356 5645 -2322
rect 5576 -2406 5645 -2356
rect 5679 -2254 5745 -2205
rect 5679 -2288 5695 -2254
rect 5729 -2288 5745 -2254
rect 5679 -2322 5745 -2288
rect 5679 -2356 5695 -2322
rect 5729 -2356 5745 -2322
rect 5679 -2372 5745 -2356
rect 5835 -2254 5905 -2239
rect 5835 -2288 5853 -2254
rect 5887 -2288 5905 -2254
rect 5835 -2322 5905 -2288
rect 5835 -2356 5853 -2322
rect 5887 -2356 5905 -2322
rect 5576 -2440 5770 -2406
rect 5116 -2527 5136 -2493
rect 5170 -2527 5266 -2493
rect 5300 -2491 5396 -2457
rect 5430 -2491 5450 -2457
rect 5700 -2469 5770 -2440
rect 5835 -2468 5905 -2356
rect 5957 -2255 6007 -2239
rect 5991 -2289 6007 -2255
rect 5957 -2323 6007 -2289
rect 5991 -2357 6007 -2323
rect 5957 -2399 6007 -2357
rect 6097 -2254 6163 -2205
rect 6097 -2288 6113 -2254
rect 6147 -2288 6163 -2254
rect 6097 -2322 6163 -2288
rect 6097 -2356 6113 -2322
rect 6147 -2356 6163 -2322
rect 6097 -2365 6163 -2356
rect 6197 -2255 6278 -2239
rect 6197 -2289 6211 -2255
rect 6245 -2289 6278 -2255
rect 6197 -2323 6278 -2289
rect 6197 -2357 6211 -2323
rect 6245 -2357 6278 -2323
rect 6197 -2394 6278 -2357
rect 5957 -2433 6075 -2399
rect 6041 -2467 6075 -2433
rect 5300 -2561 5450 -2491
rect 5576 -2478 5666 -2474
rect 5576 -2512 5615 -2478
rect 5649 -2483 5666 -2478
rect 5576 -2517 5616 -2512
rect 5650 -2517 5666 -2483
rect 5700 -2483 5786 -2469
rect 5700 -2517 5736 -2483
rect 5770 -2517 5786 -2483
rect 5700 -2527 5786 -2517
rect 5835 -2483 6007 -2468
rect 5835 -2517 5957 -2483
rect 5991 -2517 6007 -2483
rect 5835 -2518 6007 -2517
rect 6041 -2483 6194 -2467
rect 6041 -2517 6157 -2483
rect 6191 -2517 6194 -2483
rect 5700 -2551 5770 -2527
rect 3828 -2647 3846 -2613
rect 3880 -2647 4110 -2613
rect 4144 -2647 4162 -2613
rect 3828 -2715 4162 -2647
rect 4196 -2587 4254 -2570
rect 4196 -2621 4208 -2587
rect 4242 -2621 4254 -2587
rect 4196 -2715 4254 -2621
rect 4288 -2620 4990 -2561
rect 4288 -2654 4306 -2620
rect 4340 -2654 4938 -2620
rect 4972 -2654 4990 -2620
rect 4288 -2715 4990 -2654
rect 5024 -2587 5082 -2570
rect 5024 -2621 5036 -2587
rect 5070 -2621 5082 -2587
rect 5024 -2715 5082 -2621
rect 5116 -2613 5450 -2561
rect 5116 -2647 5134 -2613
rect 5168 -2647 5398 -2613
rect 5432 -2647 5450 -2613
rect 5116 -2715 5450 -2647
rect 5484 -2587 5542 -2570
rect 5484 -2621 5496 -2587
rect 5530 -2621 5542 -2587
rect 5484 -2715 5542 -2621
rect 5576 -2585 5770 -2551
rect 5576 -2628 5642 -2585
rect 5576 -2662 5595 -2628
rect 5629 -2662 5642 -2628
rect 5576 -2681 5642 -2662
rect 5676 -2628 5742 -2619
rect 5676 -2662 5692 -2628
rect 5726 -2662 5742 -2628
rect 5676 -2715 5742 -2662
rect 5835 -2628 5905 -2518
rect 6041 -2533 6194 -2517
rect 6228 -2478 6278 -2394
rect 6312 -2276 6370 -2205
rect 6312 -2310 6324 -2276
rect 6358 -2310 6370 -2276
rect 6312 -2369 6370 -2310
rect 6312 -2403 6324 -2369
rect 6358 -2403 6370 -2369
rect 6312 -2438 6370 -2403
rect 6404 -2247 6738 -2205
rect 6404 -2281 6422 -2247
rect 6456 -2281 6686 -2247
rect 6720 -2281 6738 -2247
rect 6404 -2349 6738 -2281
rect 6404 -2383 6422 -2349
rect 6456 -2383 6686 -2349
rect 6720 -2383 6738 -2349
rect 6404 -2423 6738 -2383
rect 6772 -2276 6830 -2205
rect 6772 -2310 6784 -2276
rect 6818 -2310 6830 -2276
rect 6772 -2369 6830 -2310
rect 6772 -2403 6784 -2369
rect 6818 -2403 6830 -2369
rect 6228 -2512 6229 -2478
rect 6263 -2512 6278 -2478
rect 6041 -2552 6075 -2533
rect 5835 -2662 5852 -2628
rect 5886 -2662 5905 -2628
rect 5835 -2681 5905 -2662
rect 5957 -2586 6075 -2552
rect 5957 -2628 6007 -2586
rect 6228 -2604 6278 -2512
rect 6404 -2493 6554 -2423
rect 6772 -2438 6830 -2403
rect 6864 -2247 7566 -2205
rect 6864 -2281 6882 -2247
rect 6916 -2281 7514 -2247
rect 7548 -2281 7566 -2247
rect 6864 -2349 7566 -2281
rect 6864 -2383 6882 -2349
rect 6916 -2383 7514 -2349
rect 7548 -2383 7566 -2349
rect 6864 -2423 7566 -2383
rect 6404 -2527 6424 -2493
rect 6458 -2527 6554 -2493
rect 6588 -2491 6684 -2457
rect 6718 -2491 6738 -2457
rect 6588 -2561 6738 -2491
rect 5991 -2662 6007 -2628
rect 5957 -2681 6007 -2662
rect 6097 -2628 6163 -2612
rect 6097 -2662 6113 -2628
rect 6147 -2662 6163 -2628
rect 6097 -2715 6163 -2662
rect 6197 -2628 6278 -2604
rect 6197 -2662 6211 -2628
rect 6245 -2662 6278 -2628
rect 6197 -2681 6278 -2662
rect 6312 -2587 6370 -2570
rect 6312 -2621 6324 -2587
rect 6358 -2621 6370 -2587
rect 6312 -2715 6370 -2621
rect 6404 -2613 6738 -2561
rect 6864 -2491 6942 -2457
rect 6976 -2491 7041 -2457
rect 7075 -2491 7140 -2457
rect 7174 -2491 7194 -2457
rect 6864 -2561 7194 -2491
rect 7228 -2493 7566 -2423
rect 7600 -2276 7658 -2205
rect 7600 -2310 7612 -2276
rect 7646 -2310 7658 -2276
rect 7600 -2369 7658 -2310
rect 7600 -2403 7612 -2369
rect 7646 -2403 7658 -2369
rect 7600 -2438 7658 -2403
rect 7692 -2247 8026 -2205
rect 7692 -2281 7710 -2247
rect 7744 -2281 7974 -2247
rect 8008 -2281 8026 -2247
rect 7692 -2349 8026 -2281
rect 7692 -2383 7710 -2349
rect 7744 -2383 7974 -2349
rect 8008 -2383 8026 -2349
rect 7692 -2423 8026 -2383
rect 8060 -2276 8118 -2205
rect 8060 -2310 8072 -2276
rect 8106 -2310 8118 -2276
rect 8060 -2369 8118 -2310
rect 8060 -2403 8072 -2369
rect 8106 -2403 8118 -2369
rect 7228 -2527 7248 -2493
rect 7282 -2527 7351 -2493
rect 7385 -2527 7454 -2493
rect 7488 -2527 7566 -2493
rect 7692 -2493 7842 -2423
rect 8060 -2438 8118 -2403
rect 8152 -2254 8221 -2239
rect 8152 -2288 8171 -2254
rect 8205 -2288 8221 -2254
rect 8152 -2322 8221 -2288
rect 8152 -2356 8171 -2322
rect 8205 -2356 8221 -2322
rect 8152 -2406 8221 -2356
rect 8255 -2254 8321 -2205
rect 8255 -2288 8271 -2254
rect 8305 -2288 8321 -2254
rect 8255 -2322 8321 -2288
rect 8255 -2356 8271 -2322
rect 8305 -2356 8321 -2322
rect 8255 -2372 8321 -2356
rect 8411 -2254 8481 -2239
rect 8411 -2288 8429 -2254
rect 8463 -2288 8481 -2254
rect 8411 -2322 8481 -2288
rect 8411 -2356 8429 -2322
rect 8463 -2356 8481 -2322
rect 8152 -2440 8346 -2406
rect 7692 -2527 7712 -2493
rect 7746 -2527 7842 -2493
rect 7876 -2491 7972 -2457
rect 8006 -2491 8026 -2457
rect 8276 -2469 8346 -2440
rect 8411 -2468 8481 -2356
rect 8533 -2255 8583 -2239
rect 8567 -2289 8583 -2255
rect 8533 -2323 8583 -2289
rect 8567 -2357 8583 -2323
rect 8533 -2399 8583 -2357
rect 8673 -2254 8739 -2205
rect 8673 -2288 8689 -2254
rect 8723 -2288 8739 -2254
rect 8673 -2322 8739 -2288
rect 8673 -2356 8689 -2322
rect 8723 -2356 8739 -2322
rect 8673 -2365 8739 -2356
rect 8773 -2255 8854 -2239
rect 8773 -2289 8787 -2255
rect 8821 -2289 8854 -2255
rect 8773 -2323 8854 -2289
rect 8773 -2357 8787 -2323
rect 8821 -2357 8854 -2323
rect 8773 -2394 8854 -2357
rect 8533 -2433 8651 -2399
rect 8617 -2467 8651 -2433
rect 7876 -2561 8026 -2491
rect 8152 -2478 8242 -2474
rect 8152 -2512 8189 -2478
rect 8223 -2483 8242 -2478
rect 8152 -2517 8192 -2512
rect 8226 -2517 8242 -2483
rect 8276 -2483 8362 -2469
rect 8276 -2517 8312 -2483
rect 8346 -2517 8362 -2483
rect 8276 -2527 8362 -2517
rect 8411 -2483 8583 -2468
rect 8411 -2517 8533 -2483
rect 8567 -2517 8583 -2483
rect 8411 -2518 8583 -2517
rect 8617 -2483 8770 -2467
rect 8617 -2517 8733 -2483
rect 8767 -2517 8770 -2483
rect 8276 -2551 8346 -2527
rect 6404 -2647 6422 -2613
rect 6456 -2647 6686 -2613
rect 6720 -2647 6738 -2613
rect 6404 -2715 6738 -2647
rect 6772 -2587 6830 -2570
rect 6772 -2621 6784 -2587
rect 6818 -2621 6830 -2587
rect 6772 -2715 6830 -2621
rect 6864 -2620 7566 -2561
rect 6864 -2654 6882 -2620
rect 6916 -2654 7514 -2620
rect 7548 -2654 7566 -2620
rect 6864 -2715 7566 -2654
rect 7600 -2587 7658 -2570
rect 7600 -2621 7612 -2587
rect 7646 -2621 7658 -2587
rect 7600 -2715 7658 -2621
rect 7692 -2613 8026 -2561
rect 7692 -2647 7710 -2613
rect 7744 -2647 7974 -2613
rect 8008 -2647 8026 -2613
rect 7692 -2715 8026 -2647
rect 8060 -2587 8118 -2570
rect 8060 -2621 8072 -2587
rect 8106 -2621 8118 -2587
rect 8060 -2715 8118 -2621
rect 8152 -2585 8346 -2551
rect 8152 -2628 8218 -2585
rect 8152 -2662 8171 -2628
rect 8205 -2662 8218 -2628
rect 8152 -2681 8218 -2662
rect 8252 -2628 8318 -2619
rect 8252 -2662 8268 -2628
rect 8302 -2662 8318 -2628
rect 8252 -2715 8318 -2662
rect 8411 -2628 8481 -2518
rect 8617 -2533 8770 -2517
rect 8804 -2478 8854 -2394
rect 8888 -2276 8946 -2205
rect 8888 -2310 8900 -2276
rect 8934 -2310 8946 -2276
rect 8888 -2369 8946 -2310
rect 8888 -2403 8900 -2369
rect 8934 -2403 8946 -2369
rect 8888 -2438 8946 -2403
rect 8980 -2247 9314 -2205
rect 8980 -2281 8998 -2247
rect 9032 -2281 9262 -2247
rect 9296 -2281 9314 -2247
rect 8980 -2349 9314 -2281
rect 8980 -2383 8998 -2349
rect 9032 -2383 9262 -2349
rect 9296 -2383 9314 -2349
rect 8980 -2423 9314 -2383
rect 9348 -2276 9406 -2205
rect 9348 -2310 9360 -2276
rect 9394 -2310 9406 -2276
rect 9348 -2369 9406 -2310
rect 9348 -2403 9360 -2369
rect 9394 -2403 9406 -2369
rect 8804 -2512 8806 -2478
rect 8840 -2512 8854 -2478
rect 8617 -2552 8651 -2533
rect 8411 -2662 8428 -2628
rect 8462 -2662 8481 -2628
rect 8411 -2681 8481 -2662
rect 8533 -2586 8651 -2552
rect 8533 -2628 8583 -2586
rect 8804 -2604 8854 -2512
rect 8980 -2493 9130 -2423
rect 9348 -2438 9406 -2403
rect 9440 -2247 10142 -2205
rect 9440 -2281 9458 -2247
rect 9492 -2281 10090 -2247
rect 10124 -2281 10142 -2247
rect 9440 -2349 10142 -2281
rect 9440 -2383 9458 -2349
rect 9492 -2383 10090 -2349
rect 10124 -2383 10142 -2349
rect 9440 -2423 10142 -2383
rect 8980 -2527 9000 -2493
rect 9034 -2527 9130 -2493
rect 9164 -2491 9260 -2457
rect 9294 -2491 9314 -2457
rect 9164 -2561 9314 -2491
rect 8567 -2662 8583 -2628
rect 8533 -2681 8583 -2662
rect 8673 -2628 8739 -2612
rect 8673 -2662 8689 -2628
rect 8723 -2662 8739 -2628
rect 8673 -2715 8739 -2662
rect 8773 -2628 8854 -2604
rect 8773 -2662 8787 -2628
rect 8821 -2662 8854 -2628
rect 8773 -2681 8854 -2662
rect 8888 -2587 8946 -2570
rect 8888 -2621 8900 -2587
rect 8934 -2621 8946 -2587
rect 8888 -2715 8946 -2621
rect 8980 -2613 9314 -2561
rect 9440 -2491 9518 -2457
rect 9552 -2491 9617 -2457
rect 9651 -2491 9716 -2457
rect 9750 -2491 9770 -2457
rect 9440 -2561 9770 -2491
rect 9804 -2493 10142 -2423
rect 10176 -2276 10234 -2205
rect 10176 -2310 10188 -2276
rect 10222 -2310 10234 -2276
rect 10176 -2369 10234 -2310
rect 10176 -2403 10188 -2369
rect 10222 -2403 10234 -2369
rect 10176 -2438 10234 -2403
rect 10360 -2247 10694 -2205
rect 10360 -2281 10378 -2247
rect 10412 -2281 10642 -2247
rect 10676 -2281 10694 -2247
rect 10360 -2349 10694 -2281
rect 10360 -2383 10378 -2349
rect 10412 -2383 10642 -2349
rect 10676 -2383 10694 -2349
rect 10360 -2423 10694 -2383
rect 10728 -2254 10797 -2239
rect 10728 -2288 10747 -2254
rect 10781 -2288 10797 -2254
rect 10728 -2322 10797 -2288
rect 10728 -2356 10747 -2322
rect 10781 -2356 10797 -2322
rect 10728 -2406 10797 -2356
rect 10831 -2254 10897 -2205
rect 10831 -2288 10847 -2254
rect 10881 -2288 10897 -2254
rect 10831 -2322 10897 -2288
rect 10831 -2356 10847 -2322
rect 10881 -2356 10897 -2322
rect 10831 -2372 10897 -2356
rect 10987 -2254 11057 -2239
rect 10987 -2288 11005 -2254
rect 11039 -2288 11057 -2254
rect 10987 -2322 11057 -2288
rect 10987 -2356 11005 -2322
rect 11039 -2356 11057 -2322
rect 9804 -2527 9824 -2493
rect 9858 -2527 9927 -2493
rect 9961 -2527 10030 -2493
rect 10064 -2527 10142 -2493
rect 10360 -2493 10510 -2423
rect 10728 -2440 10922 -2406
rect 10360 -2527 10380 -2493
rect 10414 -2527 10510 -2493
rect 10544 -2491 10640 -2457
rect 10674 -2491 10694 -2457
rect 10852 -2469 10922 -2440
rect 10987 -2468 11057 -2356
rect 11109 -2255 11159 -2239
rect 11143 -2289 11159 -2255
rect 11109 -2323 11159 -2289
rect 11143 -2357 11159 -2323
rect 11109 -2399 11159 -2357
rect 11249 -2254 11315 -2205
rect 11249 -2288 11265 -2254
rect 11299 -2288 11315 -2254
rect 11249 -2322 11315 -2288
rect 11249 -2356 11265 -2322
rect 11299 -2356 11315 -2322
rect 11249 -2365 11315 -2356
rect 11349 -2255 11430 -2239
rect 11349 -2289 11363 -2255
rect 11397 -2289 11430 -2255
rect 11349 -2323 11430 -2289
rect 11349 -2357 11363 -2323
rect 11397 -2357 11430 -2323
rect 11349 -2394 11430 -2357
rect 11109 -2433 11227 -2399
rect 11193 -2467 11227 -2433
rect 11380 -2445 11430 -2394
rect 11464 -2276 11522 -2205
rect 11464 -2310 11476 -2276
rect 11510 -2310 11522 -2276
rect 11464 -2369 11522 -2310
rect 11464 -2403 11476 -2369
rect 11510 -2403 11522 -2369
rect 11464 -2438 11522 -2403
rect 11648 -2247 11982 -2205
rect 11648 -2281 11666 -2247
rect 11700 -2281 11930 -2247
rect 11964 -2281 11982 -2247
rect 11648 -2349 11982 -2281
rect 11648 -2383 11666 -2349
rect 11700 -2383 11930 -2349
rect 11964 -2383 11982 -2349
rect 11648 -2423 11982 -2383
rect 12384 -2276 12442 -2205
rect 12384 -2310 12396 -2276
rect 12430 -2310 12442 -2276
rect 12384 -2369 12442 -2310
rect 12384 -2403 12396 -2369
rect 12430 -2403 12442 -2369
rect 12476 -2254 12545 -2205
rect 12476 -2288 12502 -2254
rect 12536 -2288 12545 -2254
rect 12476 -2322 12545 -2288
rect 12476 -2356 12502 -2322
rect 12536 -2356 12545 -2322
rect 12476 -2372 12545 -2356
rect 12580 -2261 12631 -2245
rect 12580 -2295 12588 -2261
rect 12622 -2295 12631 -2261
rect 12580 -2349 12631 -2295
rect 10544 -2561 10694 -2491
rect 10728 -2478 10818 -2474
rect 10728 -2512 10763 -2478
rect 10797 -2483 10818 -2478
rect 10728 -2517 10768 -2512
rect 10802 -2517 10818 -2483
rect 10852 -2483 10938 -2469
rect 10852 -2517 10888 -2483
rect 10922 -2517 10938 -2483
rect 10852 -2527 10938 -2517
rect 10987 -2483 11159 -2468
rect 10987 -2517 11109 -2483
rect 11143 -2517 11159 -2483
rect 10987 -2518 11159 -2517
rect 11193 -2483 11346 -2467
rect 11193 -2517 11309 -2483
rect 11343 -2517 11346 -2483
rect 10852 -2551 10922 -2527
rect 8980 -2647 8998 -2613
rect 9032 -2647 9262 -2613
rect 9296 -2647 9314 -2613
rect 8980 -2715 9314 -2647
rect 9348 -2587 9406 -2570
rect 9348 -2621 9360 -2587
rect 9394 -2621 9406 -2587
rect 9348 -2715 9406 -2621
rect 9440 -2620 10142 -2561
rect 9440 -2654 9458 -2620
rect 9492 -2654 10090 -2620
rect 10124 -2654 10142 -2620
rect 9440 -2715 10142 -2654
rect 10176 -2587 10234 -2570
rect 10176 -2621 10188 -2587
rect 10222 -2621 10234 -2587
rect 10176 -2715 10234 -2621
rect 10360 -2613 10694 -2561
rect 10360 -2647 10378 -2613
rect 10412 -2647 10642 -2613
rect 10676 -2647 10694 -2613
rect 10360 -2715 10694 -2647
rect 10728 -2585 10922 -2551
rect 10728 -2628 10794 -2585
rect 10728 -2662 10747 -2628
rect 10781 -2662 10794 -2628
rect 10728 -2681 10794 -2662
rect 10828 -2628 10894 -2619
rect 10828 -2662 10844 -2628
rect 10878 -2662 10894 -2628
rect 10828 -2715 10894 -2662
rect 10987 -2628 11057 -2518
rect 11193 -2533 11346 -2517
rect 11380 -2479 11386 -2445
rect 11420 -2479 11430 -2445
rect 11193 -2552 11227 -2533
rect 10987 -2662 11004 -2628
rect 11038 -2662 11057 -2628
rect 10987 -2681 11057 -2662
rect 11109 -2586 11227 -2552
rect 11109 -2628 11159 -2586
rect 11380 -2604 11430 -2479
rect 11648 -2493 11798 -2423
rect 12384 -2438 12442 -2403
rect 12580 -2383 12588 -2349
rect 12622 -2383 12631 -2349
rect 12665 -2254 12717 -2205
rect 12665 -2288 12674 -2254
rect 12708 -2288 12717 -2254
rect 12665 -2322 12717 -2288
rect 12665 -2356 12674 -2322
rect 12708 -2356 12717 -2322
rect 12665 -2372 12717 -2356
rect 12752 -2261 12803 -2245
rect 12752 -2295 12760 -2261
rect 12794 -2295 12803 -2261
rect 12752 -2349 12803 -2295
rect 12580 -2406 12631 -2383
rect 12752 -2383 12760 -2349
rect 12794 -2383 12803 -2349
rect 12837 -2254 12889 -2205
rect 12837 -2288 12846 -2254
rect 12880 -2288 12889 -2254
rect 12837 -2322 12889 -2288
rect 12837 -2356 12846 -2322
rect 12880 -2356 12889 -2322
rect 12837 -2372 12889 -2356
rect 12923 -2261 12975 -2245
rect 12923 -2295 12932 -2261
rect 12966 -2295 12975 -2261
rect 12923 -2349 12975 -2295
rect 12752 -2406 12803 -2383
rect 12923 -2383 12932 -2349
rect 12966 -2383 12975 -2349
rect 13009 -2254 13086 -2205
rect 13009 -2288 13018 -2254
rect 13052 -2288 13086 -2254
rect 13009 -2322 13086 -2288
rect 13009 -2356 13018 -2322
rect 13052 -2356 13086 -2322
rect 13009 -2372 13086 -2356
rect 13120 -2276 13178 -2205
rect 13120 -2310 13132 -2276
rect 13166 -2310 13178 -2276
rect 13120 -2369 13178 -2310
rect 12923 -2406 12975 -2383
rect 13120 -2403 13132 -2369
rect 13166 -2403 13178 -2369
rect 12480 -2407 13086 -2406
rect 12514 -2440 13086 -2407
rect 13120 -2438 13178 -2403
rect 13212 -2247 13546 -2205
rect 13212 -2281 13230 -2247
rect 13264 -2281 13494 -2247
rect 13528 -2281 13546 -2247
rect 13212 -2349 13546 -2281
rect 13212 -2383 13230 -2349
rect 13264 -2383 13494 -2349
rect 13528 -2383 13546 -2349
rect 13212 -2423 13546 -2383
rect 11648 -2527 11668 -2493
rect 11702 -2527 11798 -2493
rect 11832 -2491 11928 -2457
rect 11962 -2491 11982 -2457
rect 11832 -2561 11982 -2491
rect 11143 -2662 11159 -2628
rect 11109 -2681 11159 -2662
rect 11249 -2628 11315 -2612
rect 11249 -2662 11265 -2628
rect 11299 -2662 11315 -2628
rect 11249 -2715 11315 -2662
rect 11349 -2628 11430 -2604
rect 11349 -2662 11363 -2628
rect 11397 -2662 11430 -2628
rect 11349 -2681 11430 -2662
rect 11464 -2587 11522 -2570
rect 11464 -2621 11476 -2587
rect 11510 -2621 11522 -2587
rect 11464 -2715 11522 -2621
rect 11648 -2613 11982 -2561
rect 12480 -2481 12514 -2441
rect 13026 -2466 13086 -2440
rect 12480 -2553 12514 -2515
rect 12548 -2477 12991 -2474
rect 12548 -2479 12858 -2477
rect 12548 -2513 12568 -2479
rect 12602 -2483 12659 -2479
rect 12693 -2483 12765 -2479
rect 12799 -2483 12858 -2479
rect 12892 -2483 12942 -2477
rect 12548 -2517 12574 -2513
rect 12608 -2517 12642 -2483
rect 12693 -2513 12710 -2483
rect 12676 -2517 12710 -2513
rect 12744 -2513 12765 -2483
rect 12744 -2517 12778 -2513
rect 12812 -2517 12846 -2483
rect 12892 -2511 12914 -2483
rect 12976 -2511 12991 -2477
rect 12880 -2517 12914 -2511
rect 12948 -2517 12991 -2511
rect 12548 -2519 12991 -2517
rect 13026 -2500 13039 -2466
rect 13073 -2500 13086 -2466
rect 13026 -2543 13086 -2500
rect 13026 -2553 13042 -2543
rect 11648 -2647 11666 -2613
rect 11700 -2647 11930 -2613
rect 11964 -2647 11982 -2613
rect 11648 -2715 11982 -2647
rect 12384 -2587 12442 -2570
rect 12514 -2577 13042 -2553
rect 13076 -2577 13086 -2543
rect 13212 -2491 13232 -2457
rect 13266 -2491 13362 -2457
rect 13212 -2561 13362 -2491
rect 13396 -2493 13546 -2423
rect 13580 -2276 13638 -2205
rect 13580 -2310 13592 -2276
rect 13626 -2310 13638 -2276
rect 13580 -2369 13638 -2310
rect 13674 -2247 13733 -2205
rect 13674 -2281 13690 -2247
rect 13724 -2281 13733 -2247
rect 13674 -2315 13733 -2281
rect 13674 -2349 13690 -2315
rect 13724 -2349 13733 -2315
rect 13674 -2367 13733 -2349
rect 13769 -2255 13818 -2239
rect 13769 -2289 13776 -2255
rect 13810 -2289 13818 -2255
rect 13769 -2323 13818 -2289
rect 13769 -2357 13776 -2323
rect 13810 -2357 13818 -2323
rect 13580 -2403 13592 -2369
rect 13626 -2403 13638 -2369
rect 13580 -2438 13638 -2403
rect 13769 -2467 13818 -2357
rect 13853 -2247 13905 -2205
rect 14025 -2206 15280 -2205
rect 13853 -2281 13862 -2247
rect 13896 -2281 13905 -2247
rect 13853 -2315 13905 -2281
rect 13853 -2349 13862 -2315
rect 13896 -2349 13905 -2315
rect 13853 -2367 13905 -2349
rect 13941 -2263 13991 -2240
rect 13941 -2297 13948 -2263
rect 13982 -2297 13991 -2263
rect 13941 -2331 13991 -2297
rect 13941 -2365 13948 -2331
rect 13982 -2365 13991 -2331
rect 14025 -2247 14077 -2206
rect 14025 -2281 14034 -2247
rect 14068 -2281 14077 -2247
rect 14025 -2315 14077 -2281
rect 14025 -2349 14034 -2315
rect 14068 -2349 14077 -2315
rect 14025 -2365 14077 -2349
rect 14111 -2291 14163 -2240
rect 14111 -2325 14120 -2291
rect 14154 -2325 14163 -2291
rect 13941 -2467 13991 -2365
rect 14111 -2377 14163 -2325
rect 14197 -2271 14249 -2206
rect 14197 -2305 14206 -2271
rect 14240 -2305 14249 -2271
rect 14197 -2351 14249 -2305
rect 14283 -2291 14335 -2240
rect 14283 -2325 14292 -2291
rect 14326 -2325 14335 -2291
rect 14111 -2411 14120 -2377
rect 14154 -2385 14163 -2377
rect 14283 -2377 14335 -2325
rect 14369 -2271 14421 -2206
rect 14369 -2305 14378 -2271
rect 14412 -2305 14421 -2271
rect 14369 -2351 14421 -2305
rect 14455 -2291 14507 -2240
rect 14455 -2325 14464 -2291
rect 14498 -2325 14507 -2291
rect 14283 -2385 14292 -2377
rect 14154 -2411 14292 -2385
rect 14326 -2385 14335 -2377
rect 14455 -2377 14507 -2325
rect 14541 -2271 14593 -2206
rect 14541 -2305 14550 -2271
rect 14584 -2305 14593 -2271
rect 14541 -2351 14593 -2305
rect 14627 -2291 14679 -2240
rect 14627 -2325 14636 -2291
rect 14670 -2325 14679 -2291
rect 14455 -2385 14464 -2377
rect 14326 -2411 14464 -2385
rect 14498 -2385 14507 -2377
rect 14627 -2377 14679 -2325
rect 14713 -2271 14762 -2206
rect 14713 -2305 14722 -2271
rect 14756 -2305 14762 -2271
rect 14713 -2351 14762 -2305
rect 14796 -2291 14848 -2240
rect 14796 -2325 14807 -2291
rect 14841 -2325 14848 -2291
rect 14627 -2385 14636 -2377
rect 14498 -2411 14636 -2385
rect 14670 -2385 14679 -2377
rect 14796 -2377 14848 -2325
rect 14885 -2271 14934 -2206
rect 14885 -2305 14893 -2271
rect 14927 -2305 14934 -2271
rect 14885 -2351 14934 -2305
rect 14968 -2291 15020 -2240
rect 14968 -2325 14979 -2291
rect 15013 -2325 15020 -2291
rect 14796 -2385 14807 -2377
rect 14670 -2411 14807 -2385
rect 14841 -2385 14848 -2377
rect 14968 -2377 15020 -2325
rect 15057 -2271 15106 -2206
rect 15057 -2305 15065 -2271
rect 15099 -2305 15106 -2271
rect 15057 -2351 15106 -2305
rect 15140 -2291 15192 -2240
rect 15140 -2325 15151 -2291
rect 15185 -2325 15192 -2291
rect 14968 -2385 14979 -2377
rect 14841 -2411 14979 -2385
rect 15013 -2385 15020 -2377
rect 15140 -2377 15192 -2325
rect 15229 -2271 15280 -2206
rect 15229 -2305 15237 -2271
rect 15271 -2305 15280 -2271
rect 15229 -2351 15280 -2305
rect 15314 -2291 15372 -2240
rect 15314 -2325 15323 -2291
rect 15357 -2325 15372 -2291
rect 15140 -2385 15151 -2377
rect 15013 -2411 15151 -2385
rect 15185 -2388 15192 -2377
rect 15314 -2377 15372 -2325
rect 15406 -2271 15460 -2205
rect 15406 -2305 15409 -2271
rect 15443 -2305 15460 -2271
rect 15406 -2354 15460 -2305
rect 15512 -2276 15570 -2205
rect 15512 -2310 15524 -2276
rect 15558 -2310 15570 -2276
rect 15314 -2388 15323 -2377
rect 15185 -2411 15323 -2388
rect 15357 -2388 15372 -2377
rect 15512 -2369 15570 -2310
rect 15357 -2411 15460 -2388
rect 14111 -2426 15460 -2411
rect 14111 -2433 15248 -2426
rect 15227 -2460 15248 -2433
rect 15282 -2460 15340 -2426
rect 15374 -2460 15460 -2426
rect 15512 -2403 15524 -2369
rect 15558 -2403 15570 -2369
rect 15512 -2438 15570 -2403
rect 15604 -2247 16673 -2205
rect 15604 -2281 15622 -2247
rect 15656 -2281 16622 -2247
rect 16656 -2281 16673 -2247
rect 15604 -2349 16673 -2281
rect 15604 -2383 15622 -2349
rect 15656 -2383 16622 -2349
rect 16656 -2383 16673 -2349
rect 15604 -2423 16673 -2383
rect 13396 -2527 13492 -2493
rect 13526 -2527 13546 -2493
rect 13672 -2483 13735 -2467
rect 13672 -2510 13692 -2483
rect 13672 -2544 13685 -2510
rect 13726 -2517 13735 -2483
rect 13719 -2544 13735 -2517
rect 12514 -2587 13086 -2577
rect 13120 -2587 13178 -2570
rect 12384 -2621 12396 -2587
rect 12430 -2621 12442 -2587
rect 12384 -2715 12442 -2621
rect 12572 -2637 12631 -2621
rect 12572 -2671 12588 -2637
rect 12622 -2671 12631 -2637
rect 12572 -2715 12631 -2671
rect 12665 -2626 12717 -2587
rect 12665 -2660 12674 -2626
rect 12708 -2660 12717 -2626
rect 12665 -2676 12717 -2660
rect 12751 -2637 12803 -2621
rect 12751 -2671 12760 -2637
rect 12794 -2671 12803 -2637
rect 12751 -2715 12803 -2671
rect 12837 -2626 12888 -2587
rect 13120 -2621 13132 -2587
rect 13166 -2621 13178 -2587
rect 12837 -2660 12846 -2626
rect 12880 -2660 12888 -2626
rect 12837 -2676 12888 -2660
rect 12922 -2637 12982 -2621
rect 12922 -2671 12932 -2637
rect 12966 -2671 12982 -2637
rect 12922 -2715 12982 -2671
rect 13120 -2715 13178 -2621
rect 13212 -2613 13546 -2561
rect 13212 -2647 13230 -2613
rect 13264 -2647 13494 -2613
rect 13528 -2647 13546 -2613
rect 13212 -2715 13546 -2647
rect 13580 -2587 13638 -2570
rect 13672 -2579 13735 -2544
rect 13769 -2483 15193 -2467
rect 13769 -2517 14119 -2483
rect 14153 -2517 14187 -2483
rect 14221 -2517 14255 -2483
rect 14289 -2517 14323 -2483
rect 14357 -2517 14391 -2483
rect 14425 -2517 14459 -2483
rect 14493 -2517 14527 -2483
rect 14561 -2517 14595 -2483
rect 14629 -2517 14663 -2483
rect 14697 -2517 14731 -2483
rect 14765 -2517 14799 -2483
rect 14833 -2517 14867 -2483
rect 14901 -2517 14935 -2483
rect 14969 -2517 15003 -2483
rect 15037 -2517 15071 -2483
rect 15105 -2517 15139 -2483
rect 15173 -2517 15193 -2483
rect 13580 -2621 13592 -2587
rect 13626 -2621 13638 -2587
rect 13580 -2715 13638 -2621
rect 13672 -2639 13733 -2613
rect 13672 -2673 13690 -2639
rect 13724 -2673 13733 -2639
rect 13672 -2715 13733 -2673
rect 13769 -2626 13819 -2517
rect 13769 -2660 13776 -2626
rect 13810 -2660 13819 -2626
rect 13769 -2679 13819 -2660
rect 13853 -2626 13905 -2610
rect 13853 -2660 13862 -2626
rect 13896 -2660 13905 -2626
rect 13853 -2715 13905 -2660
rect 13941 -2626 13991 -2517
rect 15227 -2522 15460 -2460
rect 15227 -2551 15248 -2522
rect 14111 -2556 15248 -2551
rect 15282 -2556 15341 -2522
rect 15375 -2556 15460 -2522
rect 14111 -2585 15460 -2556
rect 15604 -2491 15682 -2457
rect 15716 -2491 15810 -2457
rect 15844 -2491 15938 -2457
rect 15972 -2491 16066 -2457
rect 16100 -2491 16120 -2457
rect 15604 -2561 16120 -2491
rect 16154 -2493 16673 -2423
rect 16154 -2527 16174 -2493
rect 16208 -2527 16302 -2493
rect 16336 -2527 16430 -2493
rect 16464 -2527 16558 -2493
rect 16592 -2527 16673 -2493
rect 13941 -2660 13948 -2626
rect 13982 -2660 13991 -2626
rect 13941 -2679 13991 -2660
rect 14025 -2626 14077 -2603
rect 14025 -2660 14034 -2626
rect 14068 -2660 14077 -2626
rect 14025 -2715 14077 -2660
rect 14111 -2626 14163 -2585
rect 14111 -2660 14120 -2626
rect 14154 -2660 14163 -2626
rect 14111 -2676 14163 -2660
rect 14197 -2635 14249 -2619
rect 14197 -2669 14206 -2635
rect 14240 -2669 14249 -2635
rect 14197 -2715 14249 -2669
rect 14283 -2626 14335 -2585
rect 14283 -2660 14292 -2626
rect 14326 -2660 14335 -2626
rect 14283 -2676 14335 -2660
rect 14369 -2635 14421 -2619
rect 14369 -2669 14378 -2635
rect 14412 -2669 14421 -2635
rect 14369 -2715 14421 -2669
rect 14455 -2626 14507 -2585
rect 14455 -2660 14464 -2626
rect 14498 -2660 14507 -2626
rect 14455 -2676 14507 -2660
rect 14541 -2635 14590 -2619
rect 14541 -2669 14550 -2635
rect 14584 -2669 14590 -2635
rect 14541 -2715 14590 -2669
rect 14624 -2626 14679 -2585
rect 14624 -2660 14636 -2626
rect 14670 -2660 14679 -2626
rect 14624 -2676 14679 -2660
rect 14713 -2635 14762 -2619
rect 14713 -2669 14722 -2635
rect 14756 -2669 14762 -2635
rect 14713 -2715 14762 -2669
rect 14796 -2626 14848 -2585
rect 14796 -2660 14807 -2626
rect 14841 -2660 14848 -2626
rect 14796 -2676 14848 -2660
rect 14884 -2635 14934 -2619
rect 14884 -2669 14893 -2635
rect 14927 -2669 14934 -2635
rect 14884 -2715 14934 -2669
rect 14968 -2626 15020 -2585
rect 14968 -2660 14979 -2626
rect 15013 -2660 15020 -2626
rect 14968 -2676 15020 -2660
rect 15056 -2635 15106 -2619
rect 15056 -2669 15065 -2635
rect 15099 -2669 15106 -2635
rect 15056 -2715 15106 -2669
rect 15140 -2626 15192 -2585
rect 15140 -2660 15151 -2626
rect 15185 -2660 15192 -2626
rect 15140 -2676 15192 -2660
rect 15228 -2635 15280 -2619
rect 15228 -2669 15237 -2635
rect 15271 -2669 15280 -2635
rect 15228 -2715 15280 -2669
rect 15314 -2626 15366 -2585
rect 15512 -2587 15570 -2570
rect 15314 -2660 15323 -2626
rect 15357 -2660 15366 -2626
rect 15314 -2676 15366 -2660
rect 15400 -2635 15460 -2619
rect 15400 -2669 15409 -2635
rect 15443 -2669 15460 -2635
rect 15400 -2715 15460 -2669
rect 15512 -2621 15524 -2587
rect 15558 -2621 15570 -2587
rect 15512 -2715 15570 -2621
rect 15604 -2620 16673 -2561
rect 15604 -2654 15622 -2620
rect 15656 -2654 16622 -2620
rect 16656 -2654 16673 -2620
rect 15604 -2715 16673 -2654
rect -2997 -2749 -2968 -2715
rect -2934 -2749 -2876 -2715
rect -2842 -2749 -2784 -2715
rect -2750 -2749 -2692 -2715
rect -2658 -2749 -2600 -2715
rect -2566 -2749 -2508 -2715
rect -2474 -2749 -2416 -2715
rect -2382 -2749 -2324 -2715
rect -2290 -2749 -2232 -2715
rect -2198 -2749 -2140 -2715
rect -2106 -2749 -2048 -2715
rect -2014 -2749 -1956 -2715
rect -1922 -2749 -1864 -2715
rect -1830 -2749 -1772 -2715
rect -1738 -2749 -1680 -2715
rect -1646 -2749 -1588 -2715
rect -1554 -2749 -1496 -2715
rect -1462 -2749 -1404 -2715
rect -1370 -2749 -1312 -2715
rect -1278 -2749 -1220 -2715
rect -1186 -2749 -1128 -2715
rect -1094 -2749 -1036 -2715
rect -1002 -2749 -944 -2715
rect -910 -2749 -852 -2715
rect -818 -2749 -760 -2715
rect -726 -2749 -668 -2715
rect -634 -2749 -576 -2715
rect -542 -2749 -484 -2715
rect -450 -2749 -392 -2715
rect -358 -2749 -300 -2715
rect -266 -2749 -208 -2715
rect -174 -2749 -116 -2715
rect -82 -2749 -24 -2715
rect 10 -2749 68 -2715
rect 102 -2749 160 -2715
rect 194 -2749 252 -2715
rect 286 -2749 344 -2715
rect 378 -2749 436 -2715
rect 470 -2749 528 -2715
rect 562 -2749 620 -2715
rect 654 -2749 712 -2715
rect 746 -2749 804 -2715
rect 838 -2749 896 -2715
rect 930 -2749 988 -2715
rect 1022 -2749 1080 -2715
rect 1114 -2749 1172 -2715
rect 1206 -2749 1264 -2715
rect 1298 -2749 1356 -2715
rect 1390 -2749 1448 -2715
rect 1482 -2749 1540 -2715
rect 1574 -2749 1632 -2715
rect 1666 -2749 1724 -2715
rect 1758 -2749 1816 -2715
rect 1850 -2749 1908 -2715
rect 1942 -2749 2000 -2715
rect 2034 -2749 2092 -2715
rect 2126 -2749 2184 -2715
rect 2218 -2749 2276 -2715
rect 2310 -2749 2368 -2715
rect 2402 -2749 2460 -2715
rect 2494 -2749 2552 -2715
rect 2586 -2749 2644 -2715
rect 2678 -2749 2736 -2715
rect 2770 -2749 2828 -2715
rect 2862 -2749 2920 -2715
rect 2954 -2749 3012 -2715
rect 3046 -2749 3104 -2715
rect 3138 -2749 3196 -2715
rect 3230 -2749 3288 -2715
rect 3322 -2749 3380 -2715
rect 3414 -2749 3472 -2715
rect 3506 -2749 3564 -2715
rect 3598 -2749 3656 -2715
rect 3690 -2749 3748 -2715
rect 3782 -2749 3840 -2715
rect 3874 -2749 3932 -2715
rect 3966 -2749 4024 -2715
rect 4058 -2749 4116 -2715
rect 4150 -2749 4208 -2715
rect 4242 -2749 4300 -2715
rect 4334 -2749 4392 -2715
rect 4426 -2749 4484 -2715
rect 4518 -2749 4576 -2715
rect 4610 -2749 4668 -2715
rect 4702 -2749 4760 -2715
rect 4794 -2749 4852 -2715
rect 4886 -2749 4944 -2715
rect 4978 -2749 5036 -2715
rect 5070 -2749 5128 -2715
rect 5162 -2749 5220 -2715
rect 5254 -2749 5312 -2715
rect 5346 -2749 5404 -2715
rect 5438 -2749 5496 -2715
rect 5530 -2749 5588 -2715
rect 5622 -2749 5680 -2715
rect 5714 -2749 5772 -2715
rect 5806 -2749 5864 -2715
rect 5898 -2749 5956 -2715
rect 5990 -2749 6048 -2715
rect 6082 -2749 6140 -2715
rect 6174 -2749 6232 -2715
rect 6266 -2749 6324 -2715
rect 6358 -2749 6416 -2715
rect 6450 -2749 6508 -2715
rect 6542 -2749 6600 -2715
rect 6634 -2749 6692 -2715
rect 6726 -2749 6784 -2715
rect 6818 -2749 6876 -2715
rect 6910 -2749 6968 -2715
rect 7002 -2749 7060 -2715
rect 7094 -2749 7152 -2715
rect 7186 -2749 7244 -2715
rect 7278 -2749 7336 -2715
rect 7370 -2749 7428 -2715
rect 7462 -2749 7520 -2715
rect 7554 -2749 7612 -2715
rect 7646 -2749 7704 -2715
rect 7738 -2749 7796 -2715
rect 7830 -2749 7888 -2715
rect 7922 -2749 7980 -2715
rect 8014 -2749 8072 -2715
rect 8106 -2749 8164 -2715
rect 8198 -2749 8256 -2715
rect 8290 -2749 8348 -2715
rect 8382 -2749 8440 -2715
rect 8474 -2749 8532 -2715
rect 8566 -2749 8624 -2715
rect 8658 -2749 8716 -2715
rect 8750 -2749 8808 -2715
rect 8842 -2749 8900 -2715
rect 8934 -2749 8992 -2715
rect 9026 -2749 9084 -2715
rect 9118 -2749 9176 -2715
rect 9210 -2749 9268 -2715
rect 9302 -2749 9360 -2715
rect 9394 -2749 9452 -2715
rect 9486 -2749 9544 -2715
rect 9578 -2749 9636 -2715
rect 9670 -2749 9728 -2715
rect 9762 -2749 9820 -2715
rect 9854 -2749 9912 -2715
rect 9946 -2749 10004 -2715
rect 10038 -2749 10096 -2715
rect 10130 -2749 10188 -2715
rect 10222 -2749 10280 -2715
rect 10314 -2749 10372 -2715
rect 10406 -2749 10464 -2715
rect 10498 -2749 10556 -2715
rect 10590 -2749 10648 -2715
rect 10682 -2749 10740 -2715
rect 10774 -2749 10832 -2715
rect 10866 -2749 10924 -2715
rect 10958 -2749 11016 -2715
rect 11050 -2749 11108 -2715
rect 11142 -2749 11200 -2715
rect 11234 -2749 11292 -2715
rect 11326 -2749 11384 -2715
rect 11418 -2749 11476 -2715
rect 11510 -2749 11568 -2715
rect 11602 -2749 11660 -2715
rect 11694 -2749 11752 -2715
rect 11786 -2749 11844 -2715
rect 11878 -2749 11936 -2715
rect 11970 -2749 12028 -2715
rect 12062 -2749 12120 -2715
rect 12154 -2749 12212 -2715
rect 12246 -2749 12304 -2715
rect 12338 -2749 12396 -2715
rect 12430 -2749 12488 -2715
rect 12522 -2749 12580 -2715
rect 12614 -2749 12672 -2715
rect 12706 -2749 12764 -2715
rect 12798 -2749 12856 -2715
rect 12890 -2749 12948 -2715
rect 12982 -2749 13040 -2715
rect 13074 -2749 13132 -2715
rect 13166 -2749 13224 -2715
rect 13258 -2749 13316 -2715
rect 13350 -2749 13408 -2715
rect 13442 -2749 13500 -2715
rect 13534 -2749 13592 -2715
rect 13626 -2749 13684 -2715
rect 13718 -2749 13776 -2715
rect 13810 -2749 13868 -2715
rect 13902 -2749 13960 -2715
rect 13994 -2749 14052 -2715
rect 14086 -2749 14144 -2715
rect 14178 -2749 14236 -2715
rect 14270 -2749 14328 -2715
rect 14362 -2749 14420 -2715
rect 14454 -2749 14512 -2715
rect 14546 -2749 14604 -2715
rect 14638 -2749 14696 -2715
rect 14730 -2749 14788 -2715
rect 14822 -2749 14880 -2715
rect 14914 -2749 14972 -2715
rect 15006 -2749 15064 -2715
rect 15098 -2749 15156 -2715
rect 15190 -2749 15248 -2715
rect 15282 -2749 15340 -2715
rect 15374 -2749 15432 -2715
rect 15466 -2749 15524 -2715
rect 15558 -2749 15616 -2715
rect 15650 -2749 15708 -2715
rect 15742 -2749 15800 -2715
rect 15834 -2749 15892 -2715
rect 15926 -2749 15984 -2715
rect 16018 -2749 16076 -2715
rect 16110 -2749 16168 -2715
rect 16202 -2749 16260 -2715
rect 16294 -2749 16352 -2715
rect 16386 -2749 16444 -2715
rect 16478 -2749 16536 -2715
rect 16570 -2749 16628 -2715
rect 16662 -2749 16691 -2715
rect -2980 -2810 -2278 -2749
rect -2980 -2844 -2962 -2810
rect -2928 -2844 -2330 -2810
rect -2296 -2844 -2278 -2810
rect -2980 -2903 -2278 -2844
rect -2244 -2843 -2186 -2749
rect -1882 -2802 -1817 -2783
rect -2244 -2877 -2232 -2843
rect -2198 -2877 -2186 -2843
rect -2244 -2894 -2186 -2877
rect -2980 -2971 -2902 -2937
rect -2868 -2971 -2799 -2937
rect -2765 -2971 -2696 -2937
rect -2662 -2971 -2642 -2937
rect -2980 -3041 -2642 -2971
rect -2608 -2973 -2278 -2903
rect -2608 -3007 -2588 -2973
rect -2554 -3007 -2489 -2973
rect -2455 -3007 -2390 -2973
rect -2356 -3007 -2278 -2973
rect -1968 -2947 -1920 -2807
rect -1968 -2952 -1954 -2947
rect -1968 -2986 -1960 -2952
rect -1926 -2986 -1920 -2981
rect -1968 -2997 -1920 -2986
rect -1882 -2836 -1867 -2802
rect -1833 -2836 -1817 -2802
rect -1882 -2884 -1817 -2836
rect -1783 -2800 -1726 -2749
rect -1749 -2834 -1726 -2800
rect -1783 -2850 -1726 -2834
rect -1692 -2843 -1634 -2749
rect -1692 -2877 -1680 -2843
rect -1646 -2877 -1634 -2843
rect -1882 -2915 -1726 -2884
rect -1692 -2894 -1634 -2877
rect -1600 -2810 -898 -2749
rect -1600 -2844 -1582 -2810
rect -1548 -2844 -950 -2810
rect -916 -2844 -898 -2810
rect -1600 -2903 -898 -2844
rect -864 -2810 -162 -2749
rect -864 -2844 -846 -2810
rect -812 -2844 -214 -2810
rect -180 -2844 -162 -2810
rect -864 -2903 -162 -2844
rect -128 -2843 -70 -2749
rect -128 -2877 -116 -2843
rect -82 -2877 -70 -2843
rect -128 -2894 -70 -2877
rect -36 -2817 298 -2749
rect -36 -2851 -18 -2817
rect 16 -2851 246 -2817
rect 280 -2851 298 -2817
rect -36 -2903 298 -2851
rect 332 -2843 390 -2749
rect 332 -2877 344 -2843
rect 378 -2877 390 -2843
rect 332 -2894 390 -2877
rect 424 -2802 505 -2783
rect 424 -2836 457 -2802
rect 491 -2836 505 -2802
rect 424 -2860 505 -2836
rect 539 -2802 605 -2749
rect 539 -2836 555 -2802
rect 589 -2836 605 -2802
rect 539 -2852 605 -2836
rect 695 -2802 745 -2783
rect 695 -2836 711 -2802
rect -1882 -2949 -1783 -2915
rect -1749 -2949 -1726 -2915
rect -1882 -2990 -1726 -2949
rect -1600 -2971 -1522 -2937
rect -1488 -2971 -1419 -2937
rect -1385 -2971 -1316 -2937
rect -1282 -2971 -1262 -2937
rect -2980 -3081 -2278 -3041
rect -2980 -3115 -2962 -3081
rect -2928 -3115 -2330 -3081
rect -2296 -3115 -2278 -3081
rect -2980 -3183 -2278 -3115
rect -2980 -3217 -2962 -3183
rect -2928 -3217 -2330 -3183
rect -2296 -3217 -2278 -3183
rect -2980 -3259 -2278 -3217
rect -2244 -3061 -2186 -3026
rect -2244 -3095 -2232 -3061
rect -2198 -3095 -2186 -3061
rect -2244 -3154 -2186 -3095
rect -2244 -3188 -2232 -3154
rect -2198 -3188 -2186 -3154
rect -2244 -3259 -2186 -3188
rect -1968 -3081 -1916 -3065
rect -1968 -3115 -1950 -3081
rect -1968 -3183 -1916 -3115
rect -1968 -3217 -1950 -3183
rect -1968 -3259 -1916 -3217
rect -1882 -3081 -1816 -2990
rect -1692 -3061 -1634 -3026
rect -1882 -3115 -1866 -3081
rect -1832 -3115 -1816 -3081
rect -1882 -3183 -1816 -3115
rect -1882 -3217 -1866 -3183
rect -1832 -3217 -1816 -3183
rect -1882 -3225 -1816 -3217
rect -1782 -3081 -1726 -3065
rect -1748 -3115 -1726 -3081
rect -1782 -3183 -1726 -3115
rect -1748 -3217 -1726 -3183
rect -1782 -3259 -1726 -3217
rect -1692 -3095 -1680 -3061
rect -1646 -3095 -1634 -3061
rect -1692 -3154 -1634 -3095
rect -1692 -3188 -1680 -3154
rect -1646 -3188 -1634 -3154
rect -1692 -3259 -1634 -3188
rect -1600 -3041 -1262 -2971
rect -1228 -2973 -898 -2903
rect -1228 -3007 -1208 -2973
rect -1174 -3007 -1109 -2973
rect -1075 -3007 -1010 -2973
rect -976 -3007 -898 -2973
rect -864 -2971 -786 -2937
rect -752 -2971 -683 -2937
rect -649 -2971 -580 -2937
rect -546 -2971 -526 -2937
rect -864 -3041 -526 -2971
rect -492 -2973 -162 -2903
rect -492 -3007 -472 -2973
rect -438 -3007 -373 -2973
rect -339 -3007 -274 -2973
rect -240 -3007 -162 -2973
rect -36 -2971 -16 -2937
rect 18 -2971 114 -2937
rect -1600 -3081 -898 -3041
rect -1600 -3115 -1582 -3081
rect -1548 -3115 -950 -3081
rect -916 -3115 -898 -3081
rect -1600 -3183 -898 -3115
rect -1600 -3217 -1582 -3183
rect -1548 -3217 -950 -3183
rect -916 -3217 -898 -3183
rect -1600 -3259 -898 -3217
rect -864 -3081 -162 -3041
rect -864 -3115 -846 -3081
rect -812 -3115 -214 -3081
rect -180 -3115 -162 -3081
rect -864 -3183 -162 -3115
rect -864 -3217 -846 -3183
rect -812 -3217 -214 -3183
rect -180 -3217 -162 -3183
rect -864 -3259 -162 -3217
rect -128 -3061 -70 -3026
rect -128 -3095 -116 -3061
rect -82 -3095 -70 -3061
rect -128 -3154 -70 -3095
rect -128 -3188 -116 -3154
rect -82 -3188 -70 -3154
rect -128 -3259 -70 -3188
rect -36 -3041 114 -2971
rect 148 -2973 298 -2903
rect 148 -3007 244 -2973
rect 278 -3007 298 -2973
rect 424 -2987 474 -2860
rect 695 -2878 745 -2836
rect 627 -2912 745 -2878
rect 797 -2802 867 -2783
rect 797 -2836 816 -2802
rect 850 -2836 867 -2802
rect 627 -2931 661 -2912
rect 424 -3021 429 -2987
rect 463 -3021 474 -2987
rect 508 -2947 661 -2931
rect 797 -2946 867 -2836
rect 960 -2802 1026 -2749
rect 960 -2836 976 -2802
rect 1010 -2836 1026 -2802
rect 960 -2845 1026 -2836
rect 1060 -2802 1126 -2783
rect 1060 -2836 1073 -2802
rect 1107 -2836 1126 -2802
rect 1060 -2879 1126 -2836
rect 932 -2913 1126 -2879
rect 1160 -2843 1218 -2749
rect 1160 -2877 1172 -2843
rect 1206 -2877 1218 -2843
rect 1160 -2894 1218 -2877
rect 1252 -2817 1586 -2749
rect 1252 -2851 1270 -2817
rect 1304 -2851 1534 -2817
rect 1568 -2851 1586 -2817
rect 1252 -2903 1586 -2851
rect 1620 -2843 1678 -2749
rect 1620 -2877 1632 -2843
rect 1666 -2877 1678 -2843
rect 1620 -2894 1678 -2877
rect 1712 -2810 2414 -2749
rect 1712 -2844 1730 -2810
rect 1764 -2844 2362 -2810
rect 2396 -2844 2414 -2810
rect 1712 -2903 2414 -2844
rect 2448 -2843 2506 -2749
rect 2448 -2877 2460 -2843
rect 2494 -2877 2506 -2843
rect 2448 -2894 2506 -2877
rect 2540 -2817 2874 -2749
rect 2540 -2851 2558 -2817
rect 2592 -2851 2822 -2817
rect 2856 -2851 2874 -2817
rect 2540 -2903 2874 -2851
rect 2908 -2843 2966 -2749
rect 2908 -2877 2920 -2843
rect 2954 -2877 2966 -2843
rect 2908 -2894 2966 -2877
rect 3000 -2802 3081 -2783
rect 3000 -2836 3033 -2802
rect 3067 -2836 3081 -2802
rect 3000 -2860 3081 -2836
rect 3115 -2802 3181 -2749
rect 3115 -2836 3131 -2802
rect 3165 -2836 3181 -2802
rect 3115 -2852 3181 -2836
rect 3271 -2802 3321 -2783
rect 3271 -2836 3287 -2802
rect 932 -2937 1002 -2913
rect 508 -2981 511 -2947
rect 545 -2981 661 -2947
rect 508 -2997 661 -2981
rect 695 -2947 867 -2946
rect 695 -2981 711 -2947
rect 745 -2981 867 -2947
rect 695 -2996 867 -2981
rect 916 -2947 1002 -2937
rect 916 -2981 932 -2947
rect 966 -2981 1002 -2947
rect 916 -2995 1002 -2981
rect 1036 -2981 1052 -2947
rect 1086 -2952 1126 -2947
rect 1036 -2986 1072 -2981
rect 1106 -2986 1126 -2952
rect 1036 -2990 1126 -2986
rect 1252 -2971 1272 -2937
rect 1306 -2971 1402 -2937
rect -36 -3081 298 -3041
rect -36 -3115 -18 -3081
rect 16 -3115 246 -3081
rect 280 -3115 298 -3081
rect -36 -3183 298 -3115
rect -36 -3217 -18 -3183
rect 16 -3217 246 -3183
rect 280 -3217 298 -3183
rect -36 -3259 298 -3217
rect 332 -3061 390 -3026
rect 332 -3095 344 -3061
rect 378 -3095 390 -3061
rect 332 -3154 390 -3095
rect 332 -3188 344 -3154
rect 378 -3188 390 -3154
rect 332 -3259 390 -3188
rect 424 -3070 474 -3021
rect 627 -3031 661 -2997
rect 627 -3065 745 -3031
rect 424 -3107 505 -3070
rect 424 -3141 457 -3107
rect 491 -3141 505 -3107
rect 424 -3175 505 -3141
rect 424 -3209 457 -3175
rect 491 -3209 505 -3175
rect 424 -3225 505 -3209
rect 539 -3108 605 -3099
rect 539 -3142 555 -3108
rect 589 -3142 605 -3108
rect 539 -3176 605 -3142
rect 539 -3210 555 -3176
rect 589 -3210 605 -3176
rect 539 -3259 605 -3210
rect 695 -3107 745 -3065
rect 695 -3141 711 -3107
rect 695 -3175 745 -3141
rect 695 -3209 711 -3175
rect 695 -3225 745 -3209
rect 797 -3108 867 -2996
rect 932 -3024 1002 -2995
rect 932 -3058 1126 -3024
rect 797 -3142 815 -3108
rect 849 -3142 867 -3108
rect 797 -3176 867 -3142
rect 797 -3210 815 -3176
rect 849 -3210 867 -3176
rect 797 -3225 867 -3210
rect 957 -3108 1023 -3092
rect 957 -3142 973 -3108
rect 1007 -3142 1023 -3108
rect 957 -3176 1023 -3142
rect 957 -3210 973 -3176
rect 1007 -3210 1023 -3176
rect 957 -3259 1023 -3210
rect 1057 -3108 1126 -3058
rect 1057 -3142 1073 -3108
rect 1107 -3142 1126 -3108
rect 1057 -3176 1126 -3142
rect 1057 -3210 1073 -3176
rect 1107 -3210 1126 -3176
rect 1057 -3225 1126 -3210
rect 1160 -3061 1218 -3026
rect 1160 -3095 1172 -3061
rect 1206 -3095 1218 -3061
rect 1160 -3154 1218 -3095
rect 1160 -3188 1172 -3154
rect 1206 -3188 1218 -3154
rect 1160 -3259 1218 -3188
rect 1252 -3041 1402 -2971
rect 1436 -2973 1586 -2903
rect 1436 -3007 1532 -2973
rect 1566 -3007 1586 -2973
rect 1712 -2971 1790 -2937
rect 1824 -2971 1893 -2937
rect 1927 -2971 1996 -2937
rect 2030 -2971 2050 -2937
rect 1252 -3081 1586 -3041
rect 1252 -3115 1270 -3081
rect 1304 -3115 1534 -3081
rect 1568 -3115 1586 -3081
rect 1252 -3183 1586 -3115
rect 1252 -3217 1270 -3183
rect 1304 -3217 1534 -3183
rect 1568 -3217 1586 -3183
rect 1252 -3259 1586 -3217
rect 1620 -3061 1678 -3026
rect 1620 -3095 1632 -3061
rect 1666 -3095 1678 -3061
rect 1620 -3154 1678 -3095
rect 1620 -3188 1632 -3154
rect 1666 -3188 1678 -3154
rect 1620 -3259 1678 -3188
rect 1712 -3041 2050 -2971
rect 2084 -2973 2414 -2903
rect 2084 -3007 2104 -2973
rect 2138 -3007 2203 -2973
rect 2237 -3007 2302 -2973
rect 2336 -3007 2414 -2973
rect 2540 -2971 2560 -2937
rect 2594 -2971 2690 -2937
rect 1712 -3081 2414 -3041
rect 1712 -3115 1730 -3081
rect 1764 -3115 2362 -3081
rect 2396 -3115 2414 -3081
rect 1712 -3183 2414 -3115
rect 1712 -3217 1730 -3183
rect 1764 -3217 2362 -3183
rect 2396 -3217 2414 -3183
rect 1712 -3259 2414 -3217
rect 2448 -3061 2506 -3026
rect 2448 -3095 2460 -3061
rect 2494 -3095 2506 -3061
rect 2448 -3154 2506 -3095
rect 2448 -3188 2460 -3154
rect 2494 -3188 2506 -3154
rect 2448 -3259 2506 -3188
rect 2540 -3041 2690 -2971
rect 2724 -2973 2874 -2903
rect 2724 -3007 2820 -2973
rect 2854 -3007 2874 -2973
rect 3000 -2953 3050 -2860
rect 3271 -2878 3321 -2836
rect 3203 -2912 3321 -2878
rect 3373 -2802 3443 -2783
rect 3373 -2836 3392 -2802
rect 3426 -2836 3443 -2802
rect 3203 -2931 3237 -2912
rect 3000 -2987 3016 -2953
rect 2540 -3081 2874 -3041
rect 2540 -3115 2558 -3081
rect 2592 -3115 2822 -3081
rect 2856 -3115 2874 -3081
rect 2540 -3183 2874 -3115
rect 2540 -3217 2558 -3183
rect 2592 -3217 2822 -3183
rect 2856 -3217 2874 -3183
rect 2540 -3259 2874 -3217
rect 2908 -3061 2966 -3026
rect 2908 -3095 2920 -3061
rect 2954 -3095 2966 -3061
rect 2908 -3154 2966 -3095
rect 2908 -3188 2920 -3154
rect 2954 -3188 2966 -3154
rect 2908 -3259 2966 -3188
rect 3000 -3070 3050 -2987
rect 3084 -2947 3237 -2931
rect 3373 -2946 3443 -2836
rect 3536 -2802 3602 -2749
rect 3536 -2836 3552 -2802
rect 3586 -2836 3602 -2802
rect 3536 -2845 3602 -2836
rect 3636 -2802 3702 -2783
rect 3636 -2836 3649 -2802
rect 3683 -2836 3702 -2802
rect 3636 -2879 3702 -2836
rect 3508 -2913 3702 -2879
rect 3736 -2843 3794 -2749
rect 3736 -2877 3748 -2843
rect 3782 -2877 3794 -2843
rect 3736 -2894 3794 -2877
rect 3828 -2817 4162 -2749
rect 3828 -2851 3846 -2817
rect 3880 -2851 4110 -2817
rect 4144 -2851 4162 -2817
rect 3828 -2903 4162 -2851
rect 4196 -2843 4254 -2749
rect 4196 -2877 4208 -2843
rect 4242 -2877 4254 -2843
rect 4196 -2894 4254 -2877
rect 4288 -2810 4990 -2749
rect 4288 -2844 4306 -2810
rect 4340 -2844 4938 -2810
rect 4972 -2844 4990 -2810
rect 4288 -2903 4990 -2844
rect 5024 -2843 5082 -2749
rect 5024 -2877 5036 -2843
rect 5070 -2877 5082 -2843
rect 5024 -2894 5082 -2877
rect 5116 -2817 5450 -2749
rect 5116 -2851 5134 -2817
rect 5168 -2851 5398 -2817
rect 5432 -2851 5450 -2817
rect 5116 -2903 5450 -2851
rect 5484 -2843 5542 -2749
rect 5484 -2877 5496 -2843
rect 5530 -2877 5542 -2843
rect 5484 -2894 5542 -2877
rect 5576 -2802 5657 -2783
rect 5576 -2836 5609 -2802
rect 5643 -2836 5657 -2802
rect 5576 -2860 5657 -2836
rect 5691 -2802 5757 -2749
rect 5691 -2836 5707 -2802
rect 5741 -2836 5757 -2802
rect 5691 -2852 5757 -2836
rect 5847 -2802 5897 -2783
rect 5847 -2836 5863 -2802
rect 3508 -2937 3578 -2913
rect 3084 -2981 3087 -2947
rect 3121 -2981 3237 -2947
rect 3084 -2997 3237 -2981
rect 3271 -2947 3443 -2946
rect 3271 -2981 3287 -2947
rect 3321 -2981 3443 -2947
rect 3271 -2996 3443 -2981
rect 3492 -2947 3578 -2937
rect 3492 -2981 3508 -2947
rect 3542 -2981 3578 -2947
rect 3492 -2995 3578 -2981
rect 3612 -2981 3628 -2947
rect 3662 -2953 3702 -2947
rect 3612 -2987 3630 -2981
rect 3664 -2987 3702 -2953
rect 3612 -2990 3702 -2987
rect 3828 -2971 3848 -2937
rect 3882 -2971 3978 -2937
rect 3203 -3031 3237 -2997
rect 3203 -3065 3321 -3031
rect 3000 -3107 3081 -3070
rect 3000 -3141 3033 -3107
rect 3067 -3141 3081 -3107
rect 3000 -3175 3081 -3141
rect 3000 -3209 3033 -3175
rect 3067 -3209 3081 -3175
rect 3000 -3225 3081 -3209
rect 3115 -3108 3181 -3099
rect 3115 -3142 3131 -3108
rect 3165 -3142 3181 -3108
rect 3115 -3176 3181 -3142
rect 3115 -3210 3131 -3176
rect 3165 -3210 3181 -3176
rect 3115 -3259 3181 -3210
rect 3271 -3107 3321 -3065
rect 3271 -3141 3287 -3107
rect 3271 -3175 3321 -3141
rect 3271 -3209 3287 -3175
rect 3271 -3225 3321 -3209
rect 3373 -3108 3443 -2996
rect 3508 -3024 3578 -2995
rect 3508 -3058 3702 -3024
rect 3373 -3142 3391 -3108
rect 3425 -3142 3443 -3108
rect 3373 -3176 3443 -3142
rect 3373 -3210 3391 -3176
rect 3425 -3210 3443 -3176
rect 3373 -3225 3443 -3210
rect 3533 -3108 3599 -3092
rect 3533 -3142 3549 -3108
rect 3583 -3142 3599 -3108
rect 3533 -3176 3599 -3142
rect 3533 -3210 3549 -3176
rect 3583 -3210 3599 -3176
rect 3533 -3259 3599 -3210
rect 3633 -3108 3702 -3058
rect 3633 -3142 3649 -3108
rect 3683 -3142 3702 -3108
rect 3633 -3176 3702 -3142
rect 3633 -3210 3649 -3176
rect 3683 -3210 3702 -3176
rect 3633 -3225 3702 -3210
rect 3736 -3061 3794 -3026
rect 3736 -3095 3748 -3061
rect 3782 -3095 3794 -3061
rect 3736 -3154 3794 -3095
rect 3736 -3188 3748 -3154
rect 3782 -3188 3794 -3154
rect 3736 -3259 3794 -3188
rect 3828 -3041 3978 -2971
rect 4012 -2973 4162 -2903
rect 4012 -3007 4108 -2973
rect 4142 -3007 4162 -2973
rect 4288 -2971 4366 -2937
rect 4400 -2971 4469 -2937
rect 4503 -2971 4572 -2937
rect 4606 -2971 4626 -2937
rect 3828 -3081 4162 -3041
rect 3828 -3115 3846 -3081
rect 3880 -3115 4110 -3081
rect 4144 -3115 4162 -3081
rect 3828 -3183 4162 -3115
rect 3828 -3217 3846 -3183
rect 3880 -3217 4110 -3183
rect 4144 -3217 4162 -3183
rect 3828 -3259 4162 -3217
rect 4196 -3061 4254 -3026
rect 4196 -3095 4208 -3061
rect 4242 -3095 4254 -3061
rect 4196 -3154 4254 -3095
rect 4196 -3188 4208 -3154
rect 4242 -3188 4254 -3154
rect 4196 -3259 4254 -3188
rect 4288 -3041 4626 -2971
rect 4660 -2973 4990 -2903
rect 4660 -3007 4680 -2973
rect 4714 -3007 4779 -2973
rect 4813 -3007 4878 -2973
rect 4912 -3007 4990 -2973
rect 5116 -2971 5136 -2937
rect 5170 -2971 5266 -2937
rect 4288 -3081 4990 -3041
rect 4288 -3115 4306 -3081
rect 4340 -3115 4938 -3081
rect 4972 -3115 4990 -3081
rect 4288 -3183 4990 -3115
rect 4288 -3217 4306 -3183
rect 4340 -3217 4938 -3183
rect 4972 -3217 4990 -3183
rect 4288 -3259 4990 -3217
rect 5024 -3061 5082 -3026
rect 5024 -3095 5036 -3061
rect 5070 -3095 5082 -3061
rect 5024 -3154 5082 -3095
rect 5024 -3188 5036 -3154
rect 5070 -3188 5082 -3154
rect 5024 -3259 5082 -3188
rect 5116 -3041 5266 -2971
rect 5300 -2973 5450 -2903
rect 5300 -3007 5396 -2973
rect 5430 -3007 5450 -2973
rect 5576 -2953 5626 -2860
rect 5847 -2878 5897 -2836
rect 5779 -2912 5897 -2878
rect 5949 -2802 6019 -2783
rect 5949 -2836 5968 -2802
rect 6002 -2836 6019 -2802
rect 5779 -2931 5813 -2912
rect 5576 -2987 5590 -2953
rect 5624 -2987 5626 -2953
rect 5116 -3081 5450 -3041
rect 5116 -3115 5134 -3081
rect 5168 -3115 5398 -3081
rect 5432 -3115 5450 -3081
rect 5116 -3183 5450 -3115
rect 5116 -3217 5134 -3183
rect 5168 -3217 5398 -3183
rect 5432 -3217 5450 -3183
rect 5116 -3259 5450 -3217
rect 5484 -3061 5542 -3026
rect 5484 -3095 5496 -3061
rect 5530 -3095 5542 -3061
rect 5484 -3154 5542 -3095
rect 5484 -3188 5496 -3154
rect 5530 -3188 5542 -3154
rect 5484 -3259 5542 -3188
rect 5576 -3070 5626 -2987
rect 5660 -2947 5813 -2931
rect 5949 -2946 6019 -2836
rect 6112 -2802 6178 -2749
rect 6112 -2836 6128 -2802
rect 6162 -2836 6178 -2802
rect 6112 -2845 6178 -2836
rect 6212 -2802 6278 -2783
rect 6212 -2836 6225 -2802
rect 6259 -2836 6278 -2802
rect 6212 -2879 6278 -2836
rect 6084 -2913 6278 -2879
rect 6312 -2843 6370 -2749
rect 6312 -2877 6324 -2843
rect 6358 -2877 6370 -2843
rect 6312 -2894 6370 -2877
rect 6404 -2817 6738 -2749
rect 6404 -2851 6422 -2817
rect 6456 -2851 6686 -2817
rect 6720 -2851 6738 -2817
rect 6404 -2903 6738 -2851
rect 6772 -2843 6830 -2749
rect 6772 -2877 6784 -2843
rect 6818 -2877 6830 -2843
rect 6772 -2894 6830 -2877
rect 6864 -2810 7566 -2749
rect 6864 -2844 6882 -2810
rect 6916 -2844 7514 -2810
rect 7548 -2844 7566 -2810
rect 6864 -2903 7566 -2844
rect 7600 -2843 7658 -2749
rect 7600 -2877 7612 -2843
rect 7646 -2877 7658 -2843
rect 7600 -2894 7658 -2877
rect 7692 -2817 8026 -2749
rect 7692 -2851 7710 -2817
rect 7744 -2851 7974 -2817
rect 8008 -2851 8026 -2817
rect 7692 -2903 8026 -2851
rect 8060 -2843 8118 -2749
rect 8060 -2877 8072 -2843
rect 8106 -2877 8118 -2843
rect 8060 -2894 8118 -2877
rect 8152 -2802 8233 -2783
rect 8152 -2836 8185 -2802
rect 8219 -2836 8233 -2802
rect 8152 -2860 8233 -2836
rect 8267 -2802 8333 -2749
rect 8267 -2836 8283 -2802
rect 8317 -2836 8333 -2802
rect 8267 -2852 8333 -2836
rect 8423 -2802 8473 -2783
rect 8423 -2836 8439 -2802
rect 6084 -2937 6154 -2913
rect 5660 -2981 5663 -2947
rect 5697 -2981 5813 -2947
rect 5660 -2997 5813 -2981
rect 5847 -2947 6019 -2946
rect 5847 -2981 5863 -2947
rect 5897 -2981 6019 -2947
rect 5847 -2996 6019 -2981
rect 6068 -2947 6154 -2937
rect 6068 -2981 6084 -2947
rect 6118 -2981 6154 -2947
rect 6068 -2995 6154 -2981
rect 6188 -2987 6204 -2947
rect 6238 -2987 6278 -2947
rect 6188 -2990 6278 -2987
rect 6404 -2971 6424 -2937
rect 6458 -2971 6554 -2937
rect 5779 -3031 5813 -2997
rect 5779 -3065 5897 -3031
rect 5576 -3107 5657 -3070
rect 5576 -3141 5609 -3107
rect 5643 -3141 5657 -3107
rect 5576 -3175 5657 -3141
rect 5576 -3209 5609 -3175
rect 5643 -3209 5657 -3175
rect 5576 -3225 5657 -3209
rect 5691 -3108 5757 -3099
rect 5691 -3142 5707 -3108
rect 5741 -3142 5757 -3108
rect 5691 -3176 5757 -3142
rect 5691 -3210 5707 -3176
rect 5741 -3210 5757 -3176
rect 5691 -3259 5757 -3210
rect 5847 -3107 5897 -3065
rect 5847 -3141 5863 -3107
rect 5847 -3175 5897 -3141
rect 5847 -3209 5863 -3175
rect 5847 -3225 5897 -3209
rect 5949 -3108 6019 -2996
rect 6084 -3024 6154 -2995
rect 6084 -3058 6278 -3024
rect 5949 -3142 5967 -3108
rect 6001 -3142 6019 -3108
rect 5949 -3176 6019 -3142
rect 5949 -3210 5967 -3176
rect 6001 -3210 6019 -3176
rect 5949 -3225 6019 -3210
rect 6109 -3108 6175 -3092
rect 6109 -3142 6125 -3108
rect 6159 -3142 6175 -3108
rect 6109 -3176 6175 -3142
rect 6109 -3210 6125 -3176
rect 6159 -3210 6175 -3176
rect 6109 -3259 6175 -3210
rect 6209 -3108 6278 -3058
rect 6209 -3142 6225 -3108
rect 6259 -3142 6278 -3108
rect 6209 -3176 6278 -3142
rect 6209 -3210 6225 -3176
rect 6259 -3210 6278 -3176
rect 6209 -3225 6278 -3210
rect 6312 -3061 6370 -3026
rect 6312 -3095 6324 -3061
rect 6358 -3095 6370 -3061
rect 6312 -3154 6370 -3095
rect 6312 -3188 6324 -3154
rect 6358 -3188 6370 -3154
rect 6312 -3259 6370 -3188
rect 6404 -3041 6554 -2971
rect 6588 -2973 6738 -2903
rect 6588 -3007 6684 -2973
rect 6718 -3007 6738 -2973
rect 6864 -2971 6942 -2937
rect 6976 -2971 7045 -2937
rect 7079 -2971 7148 -2937
rect 7182 -2971 7202 -2937
rect 6404 -3081 6738 -3041
rect 6404 -3115 6422 -3081
rect 6456 -3115 6686 -3081
rect 6720 -3115 6738 -3081
rect 6404 -3183 6738 -3115
rect 6404 -3217 6422 -3183
rect 6456 -3217 6686 -3183
rect 6720 -3217 6738 -3183
rect 6404 -3259 6738 -3217
rect 6772 -3061 6830 -3026
rect 6772 -3095 6784 -3061
rect 6818 -3095 6830 -3061
rect 6772 -3154 6830 -3095
rect 6772 -3188 6784 -3154
rect 6818 -3188 6830 -3154
rect 6772 -3259 6830 -3188
rect 6864 -3041 7202 -2971
rect 7236 -2973 7566 -2903
rect 7236 -3007 7256 -2973
rect 7290 -3007 7355 -2973
rect 7389 -3007 7454 -2973
rect 7488 -3007 7566 -2973
rect 7692 -2971 7712 -2937
rect 7746 -2971 7842 -2937
rect 6864 -3081 7566 -3041
rect 6864 -3115 6882 -3081
rect 6916 -3115 7514 -3081
rect 7548 -3115 7566 -3081
rect 6864 -3183 7566 -3115
rect 6864 -3217 6882 -3183
rect 6916 -3217 7514 -3183
rect 7548 -3217 7566 -3183
rect 6864 -3259 7566 -3217
rect 7600 -3061 7658 -3026
rect 7600 -3095 7612 -3061
rect 7646 -3095 7658 -3061
rect 7600 -3154 7658 -3095
rect 7600 -3188 7612 -3154
rect 7646 -3188 7658 -3154
rect 7600 -3259 7658 -3188
rect 7692 -3041 7842 -2971
rect 7876 -2973 8026 -2903
rect 7876 -3007 7972 -2973
rect 8006 -3007 8026 -2973
rect 8152 -2953 8202 -2860
rect 8423 -2878 8473 -2836
rect 8355 -2912 8473 -2878
rect 8525 -2802 8595 -2783
rect 8525 -2836 8544 -2802
rect 8578 -2836 8595 -2802
rect 8355 -2931 8389 -2912
rect 8152 -2987 8164 -2953
rect 8198 -2987 8202 -2953
rect 7692 -3081 8026 -3041
rect 7692 -3115 7710 -3081
rect 7744 -3115 7974 -3081
rect 8008 -3115 8026 -3081
rect 7692 -3183 8026 -3115
rect 7692 -3217 7710 -3183
rect 7744 -3217 7974 -3183
rect 8008 -3217 8026 -3183
rect 7692 -3259 8026 -3217
rect 8060 -3061 8118 -3026
rect 8060 -3095 8072 -3061
rect 8106 -3095 8118 -3061
rect 8060 -3154 8118 -3095
rect 8060 -3188 8072 -3154
rect 8106 -3188 8118 -3154
rect 8060 -3259 8118 -3188
rect 8152 -3070 8202 -2987
rect 8236 -2947 8389 -2931
rect 8525 -2946 8595 -2836
rect 8688 -2802 8754 -2749
rect 8688 -2836 8704 -2802
rect 8738 -2836 8754 -2802
rect 8688 -2845 8754 -2836
rect 8788 -2802 8854 -2783
rect 8788 -2836 8801 -2802
rect 8835 -2836 8854 -2802
rect 8788 -2879 8854 -2836
rect 8660 -2913 8854 -2879
rect 8888 -2843 8946 -2749
rect 8888 -2877 8900 -2843
rect 8934 -2877 8946 -2843
rect 8888 -2894 8946 -2877
rect 8980 -2817 9314 -2749
rect 8980 -2851 8998 -2817
rect 9032 -2851 9262 -2817
rect 9296 -2851 9314 -2817
rect 8980 -2903 9314 -2851
rect 9348 -2843 9406 -2749
rect 9348 -2877 9360 -2843
rect 9394 -2877 9406 -2843
rect 9348 -2894 9406 -2877
rect 9440 -2810 10142 -2749
rect 9440 -2844 9458 -2810
rect 9492 -2844 10090 -2810
rect 10124 -2844 10142 -2810
rect 9440 -2903 10142 -2844
rect 10176 -2843 10234 -2749
rect 10176 -2877 10188 -2843
rect 10222 -2877 10234 -2843
rect 10176 -2894 10234 -2877
rect 10360 -2817 10694 -2749
rect 10360 -2851 10378 -2817
rect 10412 -2851 10642 -2817
rect 10676 -2851 10694 -2817
rect 10360 -2903 10694 -2851
rect 8660 -2937 8730 -2913
rect 8236 -2981 8239 -2947
rect 8273 -2981 8389 -2947
rect 8236 -2997 8389 -2981
rect 8423 -2947 8595 -2946
rect 8423 -2981 8439 -2947
rect 8473 -2981 8595 -2947
rect 8423 -2996 8595 -2981
rect 8644 -2947 8730 -2937
rect 8644 -2981 8660 -2947
rect 8694 -2981 8730 -2947
rect 8644 -2995 8730 -2981
rect 8764 -2953 8780 -2947
rect 8764 -2987 8778 -2953
rect 8814 -2981 8854 -2947
rect 8812 -2987 8854 -2981
rect 8764 -2990 8854 -2987
rect 8980 -2971 9000 -2937
rect 9034 -2971 9130 -2937
rect 8355 -3031 8389 -2997
rect 8355 -3065 8473 -3031
rect 8152 -3107 8233 -3070
rect 8152 -3141 8185 -3107
rect 8219 -3141 8233 -3107
rect 8152 -3175 8233 -3141
rect 8152 -3209 8185 -3175
rect 8219 -3209 8233 -3175
rect 8152 -3225 8233 -3209
rect 8267 -3108 8333 -3099
rect 8267 -3142 8283 -3108
rect 8317 -3142 8333 -3108
rect 8267 -3176 8333 -3142
rect 8267 -3210 8283 -3176
rect 8317 -3210 8333 -3176
rect 8267 -3259 8333 -3210
rect 8423 -3107 8473 -3065
rect 8423 -3141 8439 -3107
rect 8423 -3175 8473 -3141
rect 8423 -3209 8439 -3175
rect 8423 -3225 8473 -3209
rect 8525 -3108 8595 -2996
rect 8660 -3024 8730 -2995
rect 8660 -3058 8854 -3024
rect 8525 -3142 8543 -3108
rect 8577 -3142 8595 -3108
rect 8525 -3176 8595 -3142
rect 8525 -3210 8543 -3176
rect 8577 -3210 8595 -3176
rect 8525 -3225 8595 -3210
rect 8685 -3108 8751 -3092
rect 8685 -3142 8701 -3108
rect 8735 -3142 8751 -3108
rect 8685 -3176 8751 -3142
rect 8685 -3210 8701 -3176
rect 8735 -3210 8751 -3176
rect 8685 -3259 8751 -3210
rect 8785 -3108 8854 -3058
rect 8785 -3142 8801 -3108
rect 8835 -3142 8854 -3108
rect 8785 -3176 8854 -3142
rect 8785 -3210 8801 -3176
rect 8835 -3210 8854 -3176
rect 8785 -3225 8854 -3210
rect 8888 -3061 8946 -3026
rect 8888 -3095 8900 -3061
rect 8934 -3095 8946 -3061
rect 8888 -3154 8946 -3095
rect 8888 -3188 8900 -3154
rect 8934 -3188 8946 -3154
rect 8888 -3259 8946 -3188
rect 8980 -3041 9130 -2971
rect 9164 -2973 9314 -2903
rect 9164 -3007 9260 -2973
rect 9294 -3007 9314 -2973
rect 9440 -2971 9518 -2937
rect 9552 -2971 9621 -2937
rect 9655 -2971 9724 -2937
rect 9758 -2971 9778 -2937
rect 8980 -3081 9314 -3041
rect 8980 -3115 8998 -3081
rect 9032 -3115 9262 -3081
rect 9296 -3115 9314 -3081
rect 8980 -3183 9314 -3115
rect 8980 -3217 8998 -3183
rect 9032 -3217 9262 -3183
rect 9296 -3217 9314 -3183
rect 8980 -3259 9314 -3217
rect 9348 -3061 9406 -3026
rect 9348 -3095 9360 -3061
rect 9394 -3095 9406 -3061
rect 9348 -3154 9406 -3095
rect 9348 -3188 9360 -3154
rect 9394 -3188 9406 -3154
rect 9348 -3259 9406 -3188
rect 9440 -3041 9778 -2971
rect 9812 -2973 10142 -2903
rect 9812 -3007 9832 -2973
rect 9866 -3007 9931 -2973
rect 9965 -3007 10030 -2973
rect 10064 -3007 10142 -2973
rect 10360 -2971 10380 -2937
rect 10414 -2971 10510 -2937
rect 9440 -3081 10142 -3041
rect 9440 -3115 9458 -3081
rect 9492 -3115 10090 -3081
rect 10124 -3115 10142 -3081
rect 9440 -3183 10142 -3115
rect 9440 -3217 9458 -3183
rect 9492 -3217 10090 -3183
rect 10124 -3217 10142 -3183
rect 9440 -3259 10142 -3217
rect 10176 -3061 10234 -3026
rect 10176 -3095 10188 -3061
rect 10222 -3095 10234 -3061
rect 10176 -3154 10234 -3095
rect 10176 -3188 10188 -3154
rect 10222 -3188 10234 -3154
rect 10176 -3259 10234 -3188
rect 10360 -3041 10510 -2971
rect 10544 -2973 10694 -2903
rect 10544 -3007 10640 -2973
rect 10674 -3007 10694 -2973
rect 10728 -2802 10809 -2783
rect 10728 -2836 10761 -2802
rect 10795 -2836 10809 -2802
rect 10728 -2860 10809 -2836
rect 10843 -2802 10909 -2749
rect 10843 -2836 10859 -2802
rect 10893 -2836 10909 -2802
rect 10843 -2852 10909 -2836
rect 10999 -2802 11049 -2783
rect 10999 -2836 11015 -2802
rect 10728 -2954 10778 -2860
rect 10999 -2878 11049 -2836
rect 10931 -2912 11049 -2878
rect 11101 -2802 11171 -2783
rect 11101 -2836 11120 -2802
rect 11154 -2836 11171 -2802
rect 10931 -2931 10965 -2912
rect 10728 -2988 10738 -2954
rect 10772 -2988 10778 -2954
rect 10360 -3081 10694 -3041
rect 10360 -3115 10378 -3081
rect 10412 -3115 10642 -3081
rect 10676 -3115 10694 -3081
rect 10360 -3183 10694 -3115
rect 10360 -3217 10378 -3183
rect 10412 -3217 10642 -3183
rect 10676 -3217 10694 -3183
rect 10360 -3259 10694 -3217
rect 10728 -3070 10778 -2988
rect 10812 -2947 10965 -2931
rect 11101 -2946 11171 -2836
rect 11264 -2802 11330 -2749
rect 11264 -2836 11280 -2802
rect 11314 -2836 11330 -2802
rect 11264 -2845 11330 -2836
rect 11364 -2802 11430 -2783
rect 11364 -2836 11377 -2802
rect 11411 -2836 11430 -2802
rect 11364 -2879 11430 -2836
rect 11236 -2913 11430 -2879
rect 11464 -2843 11522 -2749
rect 11464 -2877 11476 -2843
rect 11510 -2877 11522 -2843
rect 11464 -2894 11522 -2877
rect 11648 -2817 11982 -2749
rect 11648 -2851 11666 -2817
rect 11700 -2851 11930 -2817
rect 11964 -2851 11982 -2817
rect 11648 -2903 11982 -2851
rect 13488 -2843 13546 -2749
rect 13488 -2877 13500 -2843
rect 13534 -2877 13546 -2843
rect 13488 -2894 13546 -2877
rect 13581 -2810 14650 -2749
rect 13581 -2844 13598 -2810
rect 13632 -2844 14598 -2810
rect 14632 -2844 14650 -2810
rect 13581 -2903 14650 -2844
rect 14684 -2843 14742 -2749
rect 14684 -2877 14696 -2843
rect 14730 -2877 14742 -2843
rect 14684 -2894 14742 -2877
rect 14777 -2810 15846 -2749
rect 14777 -2844 14794 -2810
rect 14828 -2844 15794 -2810
rect 15828 -2844 15846 -2810
rect 14777 -2903 15846 -2844
rect 15880 -2843 15938 -2749
rect 15880 -2877 15892 -2843
rect 15926 -2877 15938 -2843
rect 15880 -2894 15938 -2877
rect 15972 -2810 16674 -2749
rect 15972 -2844 15990 -2810
rect 16024 -2844 16622 -2810
rect 16656 -2844 16674 -2810
rect 15972 -2903 16674 -2844
rect 11236 -2937 11306 -2913
rect 10812 -2981 10815 -2947
rect 10849 -2981 10965 -2947
rect 10812 -2997 10965 -2981
rect 10999 -2947 11171 -2946
rect 10999 -2981 11015 -2947
rect 11049 -2981 11171 -2947
rect 10999 -2996 11171 -2981
rect 11220 -2947 11306 -2937
rect 11220 -2981 11236 -2947
rect 11270 -2981 11306 -2947
rect 11220 -2995 11306 -2981
rect 11340 -2981 11356 -2947
rect 11390 -2952 11430 -2947
rect 11340 -2986 11384 -2981
rect 11418 -2986 11430 -2952
rect 11340 -2990 11430 -2986
rect 11648 -2971 11668 -2937
rect 11702 -2971 11798 -2937
rect 10931 -3031 10965 -2997
rect 10931 -3065 11049 -3031
rect 10728 -3107 10809 -3070
rect 10728 -3141 10761 -3107
rect 10795 -3141 10809 -3107
rect 10728 -3175 10809 -3141
rect 10728 -3209 10761 -3175
rect 10795 -3209 10809 -3175
rect 10728 -3225 10809 -3209
rect 10843 -3108 10909 -3099
rect 10843 -3142 10859 -3108
rect 10893 -3142 10909 -3108
rect 10843 -3176 10909 -3142
rect 10843 -3210 10859 -3176
rect 10893 -3210 10909 -3176
rect 10843 -3259 10909 -3210
rect 10999 -3107 11049 -3065
rect 10999 -3141 11015 -3107
rect 10999 -3175 11049 -3141
rect 10999 -3209 11015 -3175
rect 10999 -3225 11049 -3209
rect 11101 -3108 11171 -2996
rect 11236 -3024 11306 -2995
rect 11236 -3058 11430 -3024
rect 11101 -3142 11119 -3108
rect 11153 -3142 11171 -3108
rect 11101 -3176 11171 -3142
rect 11101 -3210 11119 -3176
rect 11153 -3210 11171 -3176
rect 11101 -3225 11171 -3210
rect 11261 -3108 11327 -3092
rect 11261 -3142 11277 -3108
rect 11311 -3142 11327 -3108
rect 11261 -3176 11327 -3142
rect 11261 -3210 11277 -3176
rect 11311 -3210 11327 -3176
rect 11261 -3259 11327 -3210
rect 11361 -3108 11430 -3058
rect 11361 -3142 11377 -3108
rect 11411 -3142 11430 -3108
rect 11361 -3176 11430 -3142
rect 11361 -3210 11377 -3176
rect 11411 -3210 11430 -3176
rect 11361 -3225 11430 -3210
rect 11464 -3061 11522 -3026
rect 11464 -3095 11476 -3061
rect 11510 -3095 11522 -3061
rect 11464 -3154 11522 -3095
rect 11464 -3188 11476 -3154
rect 11510 -3188 11522 -3154
rect 11464 -3259 11522 -3188
rect 11648 -3041 11798 -2971
rect 11832 -2973 11982 -2903
rect 11832 -3007 11928 -2973
rect 11962 -3007 11982 -2973
rect 13581 -2971 13662 -2937
rect 13696 -2971 13790 -2937
rect 13824 -2971 13918 -2937
rect 13952 -2971 14046 -2937
rect 14080 -2971 14100 -2937
rect 11648 -3081 11982 -3041
rect 11648 -3115 11666 -3081
rect 11700 -3115 11930 -3081
rect 11964 -3115 11982 -3081
rect 11648 -3183 11982 -3115
rect 11648 -3217 11666 -3183
rect 11700 -3217 11930 -3183
rect 11964 -3217 11982 -3183
rect 11648 -3259 11982 -3217
rect 13488 -3061 13546 -3026
rect 13488 -3095 13500 -3061
rect 13534 -3095 13546 -3061
rect 13488 -3154 13546 -3095
rect 13488 -3188 13500 -3154
rect 13534 -3188 13546 -3154
rect 13488 -3259 13546 -3188
rect 13581 -3041 14100 -2971
rect 14134 -2973 14650 -2903
rect 14134 -3007 14154 -2973
rect 14188 -3007 14282 -2973
rect 14316 -3007 14410 -2973
rect 14444 -3007 14538 -2973
rect 14572 -3007 14650 -2973
rect 14777 -2971 14858 -2937
rect 14892 -2971 14986 -2937
rect 15020 -2971 15114 -2937
rect 15148 -2971 15242 -2937
rect 15276 -2971 15296 -2937
rect 13581 -3081 14650 -3041
rect 13581 -3115 13598 -3081
rect 13632 -3115 14598 -3081
rect 14632 -3115 14650 -3081
rect 13581 -3183 14650 -3115
rect 13581 -3217 13598 -3183
rect 13632 -3217 14598 -3183
rect 14632 -3217 14650 -3183
rect 13581 -3259 14650 -3217
rect 14684 -3061 14742 -3026
rect 14684 -3095 14696 -3061
rect 14730 -3095 14742 -3061
rect 14684 -3154 14742 -3095
rect 14684 -3188 14696 -3154
rect 14730 -3188 14742 -3154
rect 14684 -3259 14742 -3188
rect 14777 -3041 15296 -2971
rect 15330 -2973 15846 -2903
rect 15330 -3007 15350 -2973
rect 15384 -3007 15478 -2973
rect 15512 -3007 15606 -2973
rect 15640 -3007 15734 -2973
rect 15768 -3007 15846 -2973
rect 15972 -2971 16050 -2937
rect 16084 -2971 16153 -2937
rect 16187 -2971 16256 -2937
rect 16290 -2971 16310 -2937
rect 14777 -3081 15846 -3041
rect 14777 -3115 14794 -3081
rect 14828 -3115 15794 -3081
rect 15828 -3115 15846 -3081
rect 14777 -3183 15846 -3115
rect 14777 -3217 14794 -3183
rect 14828 -3217 15794 -3183
rect 15828 -3217 15846 -3183
rect 14777 -3259 15846 -3217
rect 15880 -3061 15938 -3026
rect 15880 -3095 15892 -3061
rect 15926 -3095 15938 -3061
rect 15880 -3154 15938 -3095
rect 15880 -3188 15892 -3154
rect 15926 -3188 15938 -3154
rect 15880 -3259 15938 -3188
rect 15972 -3041 16310 -2971
rect 16344 -2973 16674 -2903
rect 16344 -3007 16364 -2973
rect 16398 -3007 16463 -2973
rect 16497 -3007 16562 -2973
rect 16596 -3007 16674 -2973
rect 15972 -3081 16674 -3041
rect 15972 -3115 15990 -3081
rect 16024 -3115 16622 -3081
rect 16656 -3115 16674 -3081
rect 15972 -3183 16674 -3115
rect 15972 -3217 15990 -3183
rect 16024 -3217 16622 -3183
rect 16656 -3217 16674 -3183
rect 15972 -3259 16674 -3217
rect -2997 -3293 -2968 -3259
rect -2934 -3293 -2876 -3259
rect -2842 -3293 -2784 -3259
rect -2750 -3293 -2692 -3259
rect -2658 -3293 -2600 -3259
rect -2566 -3293 -2508 -3259
rect -2474 -3293 -2416 -3259
rect -2382 -3293 -2324 -3259
rect -2290 -3293 -2232 -3259
rect -2198 -3293 -2140 -3259
rect -2106 -3293 -2048 -3259
rect -2014 -3293 -1956 -3259
rect -1922 -3293 -1864 -3259
rect -1830 -3293 -1772 -3259
rect -1738 -3293 -1680 -3259
rect -1646 -3293 -1588 -3259
rect -1554 -3293 -1496 -3259
rect -1462 -3293 -1404 -3259
rect -1370 -3293 -1312 -3259
rect -1278 -3293 -1220 -3259
rect -1186 -3293 -1128 -3259
rect -1094 -3293 -1036 -3259
rect -1002 -3293 -944 -3259
rect -910 -3293 -852 -3259
rect -818 -3293 -760 -3259
rect -726 -3293 -668 -3259
rect -634 -3293 -576 -3259
rect -542 -3293 -484 -3259
rect -450 -3293 -392 -3259
rect -358 -3293 -300 -3259
rect -266 -3293 -208 -3259
rect -174 -3293 -116 -3259
rect -82 -3293 -24 -3259
rect 10 -3293 68 -3259
rect 102 -3293 160 -3259
rect 194 -3293 252 -3259
rect 286 -3293 344 -3259
rect 378 -3293 436 -3259
rect 470 -3293 528 -3259
rect 562 -3293 620 -3259
rect 654 -3293 712 -3259
rect 746 -3293 804 -3259
rect 838 -3293 896 -3259
rect 930 -3293 988 -3259
rect 1022 -3293 1080 -3259
rect 1114 -3293 1172 -3259
rect 1206 -3293 1264 -3259
rect 1298 -3293 1356 -3259
rect 1390 -3293 1448 -3259
rect 1482 -3293 1540 -3259
rect 1574 -3293 1632 -3259
rect 1666 -3293 1724 -3259
rect 1758 -3293 1816 -3259
rect 1850 -3293 1908 -3259
rect 1942 -3293 2000 -3259
rect 2034 -3293 2092 -3259
rect 2126 -3293 2184 -3259
rect 2218 -3293 2276 -3259
rect 2310 -3293 2368 -3259
rect 2402 -3293 2460 -3259
rect 2494 -3293 2552 -3259
rect 2586 -3293 2644 -3259
rect 2678 -3293 2736 -3259
rect 2770 -3293 2828 -3259
rect 2862 -3293 2920 -3259
rect 2954 -3293 3012 -3259
rect 3046 -3293 3104 -3259
rect 3138 -3293 3196 -3259
rect 3230 -3293 3288 -3259
rect 3322 -3293 3380 -3259
rect 3414 -3293 3472 -3259
rect 3506 -3293 3564 -3259
rect 3598 -3293 3656 -3259
rect 3690 -3293 3748 -3259
rect 3782 -3293 3840 -3259
rect 3874 -3293 3932 -3259
rect 3966 -3293 4024 -3259
rect 4058 -3293 4116 -3259
rect 4150 -3293 4208 -3259
rect 4242 -3293 4300 -3259
rect 4334 -3293 4392 -3259
rect 4426 -3293 4484 -3259
rect 4518 -3293 4576 -3259
rect 4610 -3293 4668 -3259
rect 4702 -3293 4760 -3259
rect 4794 -3293 4852 -3259
rect 4886 -3293 4944 -3259
rect 4978 -3293 5036 -3259
rect 5070 -3293 5128 -3259
rect 5162 -3293 5220 -3259
rect 5254 -3293 5312 -3259
rect 5346 -3293 5404 -3259
rect 5438 -3293 5496 -3259
rect 5530 -3293 5588 -3259
rect 5622 -3293 5680 -3259
rect 5714 -3293 5772 -3259
rect 5806 -3293 5864 -3259
rect 5898 -3293 5956 -3259
rect 5990 -3293 6048 -3259
rect 6082 -3293 6140 -3259
rect 6174 -3293 6232 -3259
rect 6266 -3293 6324 -3259
rect 6358 -3293 6416 -3259
rect 6450 -3293 6508 -3259
rect 6542 -3293 6600 -3259
rect 6634 -3293 6692 -3259
rect 6726 -3293 6784 -3259
rect 6818 -3293 6876 -3259
rect 6910 -3293 6968 -3259
rect 7002 -3293 7060 -3259
rect 7094 -3293 7152 -3259
rect 7186 -3293 7244 -3259
rect 7278 -3293 7336 -3259
rect 7370 -3293 7428 -3259
rect 7462 -3293 7520 -3259
rect 7554 -3293 7612 -3259
rect 7646 -3293 7704 -3259
rect 7738 -3293 7796 -3259
rect 7830 -3293 7888 -3259
rect 7922 -3293 7980 -3259
rect 8014 -3293 8072 -3259
rect 8106 -3293 8164 -3259
rect 8198 -3293 8256 -3259
rect 8290 -3293 8348 -3259
rect 8382 -3293 8440 -3259
rect 8474 -3293 8532 -3259
rect 8566 -3293 8624 -3259
rect 8658 -3293 8716 -3259
rect 8750 -3293 8808 -3259
rect 8842 -3293 8900 -3259
rect 8934 -3293 8992 -3259
rect 9026 -3293 9084 -3259
rect 9118 -3293 9176 -3259
rect 9210 -3293 9268 -3259
rect 9302 -3293 9360 -3259
rect 9394 -3293 9452 -3259
rect 9486 -3293 9544 -3259
rect 9578 -3293 9636 -3259
rect 9670 -3293 9728 -3259
rect 9762 -3293 9820 -3259
rect 9854 -3293 9912 -3259
rect 9946 -3293 10004 -3259
rect 10038 -3293 10096 -3259
rect 10130 -3293 10188 -3259
rect 10222 -3293 10280 -3259
rect 10314 -3293 10372 -3259
rect 10406 -3293 10464 -3259
rect 10498 -3293 10556 -3259
rect 10590 -3293 10648 -3259
rect 10682 -3293 10740 -3259
rect 10774 -3293 10832 -3259
rect 10866 -3293 10924 -3259
rect 10958 -3293 11016 -3259
rect 11050 -3293 11108 -3259
rect 11142 -3293 11200 -3259
rect 11234 -3293 11292 -3259
rect 11326 -3293 11384 -3259
rect 11418 -3293 11476 -3259
rect 11510 -3293 11568 -3259
rect 11602 -3293 11660 -3259
rect 11694 -3293 11752 -3259
rect 11786 -3293 11844 -3259
rect 11878 -3293 11936 -3259
rect 11970 -3293 12028 -3259
rect 12062 -3293 12120 -3259
rect 12154 -3293 12212 -3259
rect 12246 -3293 12304 -3259
rect 12338 -3293 12396 -3259
rect 12430 -3293 12488 -3259
rect 12522 -3293 12580 -3259
rect 12614 -3293 12672 -3259
rect 12706 -3293 12764 -3259
rect 12798 -3293 12856 -3259
rect 12890 -3293 12948 -3259
rect 12982 -3293 13040 -3259
rect 13074 -3293 13132 -3259
rect 13166 -3293 13224 -3259
rect 13258 -3293 13316 -3259
rect 13350 -3293 13408 -3259
rect 13442 -3293 13500 -3259
rect 13534 -3293 13592 -3259
rect 13626 -3293 13684 -3259
rect 13718 -3293 13776 -3259
rect 13810 -3293 13868 -3259
rect 13902 -3293 13960 -3259
rect 13994 -3293 14052 -3259
rect 14086 -3293 14144 -3259
rect 14178 -3293 14236 -3259
rect 14270 -3293 14328 -3259
rect 14362 -3293 14420 -3259
rect 14454 -3293 14512 -3259
rect 14546 -3293 14604 -3259
rect 14638 -3293 14696 -3259
rect 14730 -3293 14788 -3259
rect 14822 -3293 14880 -3259
rect 14914 -3293 14972 -3259
rect 15006 -3293 15064 -3259
rect 15098 -3293 15156 -3259
rect 15190 -3293 15248 -3259
rect 15282 -3293 15340 -3259
rect 15374 -3293 15432 -3259
rect 15466 -3293 15524 -3259
rect 15558 -3293 15616 -3259
rect 15650 -3293 15708 -3259
rect 15742 -3293 15800 -3259
rect 15834 -3293 15892 -3259
rect 15926 -3293 15984 -3259
rect 16018 -3293 16076 -3259
rect 16110 -3293 16168 -3259
rect 16202 -3293 16260 -3259
rect 16294 -3293 16352 -3259
rect 16386 -3293 16444 -3259
rect 16478 -3293 16536 -3259
rect 16570 -3293 16628 -3259
rect 16662 -3293 16691 -3259
rect -2980 -3335 -2278 -3293
rect -2980 -3369 -2962 -3335
rect -2928 -3369 -2330 -3335
rect -2296 -3369 -2278 -3335
rect -2980 -3437 -2278 -3369
rect -2980 -3471 -2962 -3437
rect -2928 -3471 -2330 -3437
rect -2296 -3471 -2278 -3437
rect -2980 -3511 -2278 -3471
rect -2980 -3579 -2902 -3545
rect -2868 -3579 -2803 -3545
rect -2769 -3579 -2704 -3545
rect -2670 -3579 -2650 -3545
rect -2980 -3649 -2650 -3579
rect -2616 -3581 -2278 -3511
rect -2244 -3364 -2186 -3293
rect -2244 -3398 -2232 -3364
rect -2198 -3398 -2186 -3364
rect -2244 -3457 -2186 -3398
rect -2244 -3491 -2232 -3457
rect -2198 -3491 -2186 -3457
rect -2244 -3526 -2186 -3491
rect -1600 -3335 -898 -3293
rect -1600 -3369 -1582 -3335
rect -1548 -3369 -950 -3335
rect -916 -3369 -898 -3335
rect -1600 -3437 -898 -3369
rect -1600 -3471 -1582 -3437
rect -1548 -3471 -950 -3437
rect -916 -3471 -898 -3437
rect -1600 -3511 -898 -3471
rect -864 -3335 -162 -3293
rect -864 -3369 -846 -3335
rect -812 -3369 -214 -3335
rect -180 -3369 -162 -3335
rect -864 -3437 -162 -3369
rect -864 -3471 -846 -3437
rect -812 -3471 -214 -3437
rect -180 -3471 -162 -3437
rect -864 -3511 -162 -3471
rect -128 -3364 -70 -3293
rect -128 -3398 -116 -3364
rect -82 -3398 -70 -3364
rect -128 -3457 -70 -3398
rect -128 -3491 -116 -3457
rect -82 -3491 -70 -3457
rect -2616 -3615 -2596 -3581
rect -2562 -3615 -2493 -3581
rect -2459 -3615 -2390 -3581
rect -2356 -3615 -2278 -3581
rect -1600 -3581 -1262 -3511
rect -1600 -3615 -1522 -3581
rect -1488 -3615 -1419 -3581
rect -1385 -3615 -1316 -3581
rect -1282 -3615 -1262 -3581
rect -1228 -3579 -1208 -3545
rect -1174 -3579 -1109 -3545
rect -1075 -3579 -1010 -3545
rect -976 -3579 -898 -3545
rect -1228 -3649 -898 -3579
rect -864 -3581 -526 -3511
rect -128 -3526 -70 -3491
rect -36 -3335 298 -3293
rect -36 -3369 -18 -3335
rect 16 -3369 246 -3335
rect 280 -3369 298 -3335
rect -36 -3437 298 -3369
rect -36 -3471 -18 -3437
rect 16 -3471 246 -3437
rect 280 -3471 298 -3437
rect -36 -3511 298 -3471
rect 332 -3364 390 -3293
rect 332 -3398 344 -3364
rect 378 -3398 390 -3364
rect 332 -3457 390 -3398
rect 332 -3491 344 -3457
rect 378 -3491 390 -3457
rect -864 -3615 -786 -3581
rect -752 -3615 -683 -3581
rect -649 -3615 -580 -3581
rect -546 -3615 -526 -3581
rect -492 -3579 -472 -3545
rect -438 -3579 -373 -3545
rect -339 -3579 -274 -3545
rect -240 -3579 -162 -3545
rect -492 -3649 -162 -3579
rect -36 -3581 114 -3511
rect 332 -3526 390 -3491
rect 424 -3343 505 -3327
rect 424 -3377 457 -3343
rect 491 -3377 505 -3343
rect 424 -3411 505 -3377
rect 424 -3445 457 -3411
rect 491 -3445 505 -3411
rect 424 -3482 505 -3445
rect 539 -3342 605 -3293
rect 539 -3376 555 -3342
rect 589 -3376 605 -3342
rect 539 -3410 605 -3376
rect 539 -3444 555 -3410
rect 589 -3444 605 -3410
rect 539 -3453 605 -3444
rect 695 -3343 745 -3327
rect 695 -3377 711 -3343
rect 695 -3411 745 -3377
rect 695 -3445 711 -3411
rect 424 -3531 474 -3482
rect 695 -3487 745 -3445
rect -36 -3615 -16 -3581
rect 18 -3615 114 -3581
rect 148 -3579 244 -3545
rect 278 -3579 298 -3545
rect 148 -3649 298 -3579
rect -2980 -3708 -2278 -3649
rect -2980 -3742 -2962 -3708
rect -2928 -3742 -2330 -3708
rect -2296 -3742 -2278 -3708
rect -2980 -3803 -2278 -3742
rect -2244 -3675 -2186 -3658
rect -2244 -3709 -2232 -3675
rect -2198 -3709 -2186 -3675
rect -2244 -3803 -2186 -3709
rect -1600 -3708 -898 -3649
rect -1600 -3742 -1582 -3708
rect -1548 -3742 -950 -3708
rect -916 -3742 -898 -3708
rect -1600 -3803 -898 -3742
rect -864 -3708 -162 -3649
rect -864 -3742 -846 -3708
rect -812 -3742 -214 -3708
rect -180 -3742 -162 -3708
rect -864 -3803 -162 -3742
rect -128 -3675 -70 -3658
rect -128 -3709 -116 -3675
rect -82 -3709 -70 -3675
rect -128 -3803 -70 -3709
rect -36 -3701 298 -3649
rect 424 -3565 432 -3531
rect 466 -3565 474 -3531
rect 627 -3521 745 -3487
rect 797 -3342 867 -3327
rect 797 -3376 815 -3342
rect 849 -3376 867 -3342
rect 797 -3410 867 -3376
rect 797 -3444 815 -3410
rect 849 -3444 867 -3410
rect 627 -3555 661 -3521
rect -36 -3735 -18 -3701
rect 16 -3735 246 -3701
rect 280 -3735 298 -3701
rect -36 -3803 298 -3735
rect 332 -3675 390 -3658
rect 332 -3709 344 -3675
rect 378 -3709 390 -3675
rect 332 -3803 390 -3709
rect 424 -3692 474 -3565
rect 508 -3571 661 -3555
rect 797 -3556 867 -3444
rect 957 -3342 1023 -3293
rect 957 -3376 973 -3342
rect 1007 -3376 1023 -3342
rect 957 -3410 1023 -3376
rect 957 -3444 973 -3410
rect 1007 -3444 1023 -3410
rect 957 -3460 1023 -3444
rect 1057 -3342 1126 -3327
rect 1057 -3376 1073 -3342
rect 1107 -3376 1126 -3342
rect 1057 -3410 1126 -3376
rect 1057 -3444 1073 -3410
rect 1107 -3444 1126 -3410
rect 1057 -3494 1126 -3444
rect 508 -3605 511 -3571
rect 545 -3605 661 -3571
rect 508 -3621 661 -3605
rect 695 -3571 867 -3556
rect 932 -3528 1126 -3494
rect 1160 -3364 1218 -3293
rect 1160 -3398 1172 -3364
rect 1206 -3398 1218 -3364
rect 1160 -3457 1218 -3398
rect 1160 -3491 1172 -3457
rect 1206 -3491 1218 -3457
rect 1160 -3526 1218 -3491
rect 1252 -3335 1586 -3293
rect 1252 -3369 1270 -3335
rect 1304 -3369 1534 -3335
rect 1568 -3369 1586 -3335
rect 1252 -3437 1586 -3369
rect 1252 -3471 1270 -3437
rect 1304 -3471 1534 -3437
rect 1568 -3471 1586 -3437
rect 1252 -3511 1586 -3471
rect 1620 -3364 1678 -3293
rect 1620 -3398 1632 -3364
rect 1666 -3398 1678 -3364
rect 1620 -3457 1678 -3398
rect 1620 -3491 1632 -3457
rect 1666 -3491 1678 -3457
rect 932 -3557 1002 -3528
rect 695 -3605 711 -3571
rect 745 -3605 867 -3571
rect 695 -3606 867 -3605
rect 627 -3640 661 -3621
rect 627 -3674 745 -3640
rect 424 -3716 505 -3692
rect 424 -3750 457 -3716
rect 491 -3750 505 -3716
rect 424 -3769 505 -3750
rect 539 -3716 605 -3700
rect 539 -3750 555 -3716
rect 589 -3750 605 -3716
rect 539 -3803 605 -3750
rect 695 -3716 745 -3674
rect 695 -3750 711 -3716
rect 695 -3769 745 -3750
rect 797 -3716 867 -3606
rect 916 -3571 1002 -3557
rect 916 -3605 932 -3571
rect 966 -3605 1002 -3571
rect 1036 -3568 1126 -3562
rect 1036 -3571 1070 -3568
rect 1036 -3605 1052 -3571
rect 1104 -3602 1126 -3568
rect 1086 -3605 1126 -3602
rect 1252 -3581 1402 -3511
rect 1620 -3526 1678 -3491
rect 1712 -3335 2414 -3293
rect 1712 -3369 1730 -3335
rect 1764 -3369 2362 -3335
rect 2396 -3369 2414 -3335
rect 1712 -3437 2414 -3369
rect 1712 -3471 1730 -3437
rect 1764 -3471 2362 -3437
rect 2396 -3471 2414 -3437
rect 1712 -3511 2414 -3471
rect 916 -3615 1002 -3605
rect 1252 -3615 1272 -3581
rect 1306 -3615 1402 -3581
rect 1436 -3579 1532 -3545
rect 1566 -3579 1586 -3545
rect 932 -3639 1002 -3615
rect 932 -3673 1126 -3639
rect 1436 -3649 1586 -3579
rect 797 -3750 816 -3716
rect 850 -3750 867 -3716
rect 797 -3769 867 -3750
rect 960 -3716 1026 -3707
rect 960 -3750 976 -3716
rect 1010 -3750 1026 -3716
rect 960 -3803 1026 -3750
rect 1060 -3716 1126 -3673
rect 1060 -3750 1073 -3716
rect 1107 -3750 1126 -3716
rect 1060 -3769 1126 -3750
rect 1160 -3675 1218 -3658
rect 1160 -3709 1172 -3675
rect 1206 -3709 1218 -3675
rect 1160 -3803 1218 -3709
rect 1252 -3701 1586 -3649
rect 1712 -3579 1790 -3545
rect 1824 -3579 1889 -3545
rect 1923 -3579 1988 -3545
rect 2022 -3579 2042 -3545
rect 1712 -3649 2042 -3579
rect 2076 -3581 2414 -3511
rect 2448 -3364 2506 -3293
rect 2448 -3398 2460 -3364
rect 2494 -3398 2506 -3364
rect 2448 -3457 2506 -3398
rect 2448 -3491 2460 -3457
rect 2494 -3491 2506 -3457
rect 2448 -3526 2506 -3491
rect 2540 -3335 2874 -3293
rect 2540 -3369 2558 -3335
rect 2592 -3369 2822 -3335
rect 2856 -3369 2874 -3335
rect 2540 -3437 2874 -3369
rect 2540 -3471 2558 -3437
rect 2592 -3471 2822 -3437
rect 2856 -3471 2874 -3437
rect 2540 -3511 2874 -3471
rect 2908 -3364 2966 -3293
rect 2908 -3398 2920 -3364
rect 2954 -3398 2966 -3364
rect 2908 -3457 2966 -3398
rect 2908 -3491 2920 -3457
rect 2954 -3491 2966 -3457
rect 2076 -3615 2096 -3581
rect 2130 -3615 2199 -3581
rect 2233 -3615 2302 -3581
rect 2336 -3615 2414 -3581
rect 2540 -3581 2690 -3511
rect 2908 -3526 2966 -3491
rect 3000 -3343 3081 -3327
rect 3000 -3377 3033 -3343
rect 3067 -3377 3081 -3343
rect 3000 -3411 3081 -3377
rect 3000 -3445 3033 -3411
rect 3067 -3445 3081 -3411
rect 3000 -3482 3081 -3445
rect 3115 -3342 3181 -3293
rect 3115 -3376 3131 -3342
rect 3165 -3376 3181 -3342
rect 3115 -3410 3181 -3376
rect 3115 -3444 3131 -3410
rect 3165 -3444 3181 -3410
rect 3115 -3453 3181 -3444
rect 3271 -3343 3321 -3327
rect 3271 -3377 3287 -3343
rect 3271 -3411 3321 -3377
rect 3271 -3445 3287 -3411
rect 2540 -3615 2560 -3581
rect 2594 -3615 2690 -3581
rect 2724 -3579 2820 -3545
rect 2854 -3579 2874 -3545
rect 2724 -3649 2874 -3579
rect 1252 -3735 1270 -3701
rect 1304 -3735 1534 -3701
rect 1568 -3735 1586 -3701
rect 1252 -3803 1586 -3735
rect 1620 -3675 1678 -3658
rect 1620 -3709 1632 -3675
rect 1666 -3709 1678 -3675
rect 1620 -3803 1678 -3709
rect 1712 -3708 2414 -3649
rect 1712 -3742 1730 -3708
rect 1764 -3742 2362 -3708
rect 2396 -3742 2414 -3708
rect 1712 -3803 2414 -3742
rect 2448 -3675 2506 -3658
rect 2448 -3709 2460 -3675
rect 2494 -3709 2506 -3675
rect 2448 -3803 2506 -3709
rect 2540 -3701 2874 -3649
rect 3000 -3565 3050 -3482
rect 3271 -3487 3321 -3445
rect 3203 -3521 3321 -3487
rect 3373 -3342 3443 -3327
rect 3373 -3376 3391 -3342
rect 3425 -3376 3443 -3342
rect 3373 -3410 3443 -3376
rect 3373 -3444 3391 -3410
rect 3425 -3444 3443 -3410
rect 3203 -3555 3237 -3521
rect 3000 -3599 3016 -3565
rect 2540 -3735 2558 -3701
rect 2592 -3735 2822 -3701
rect 2856 -3735 2874 -3701
rect 2540 -3803 2874 -3735
rect 2908 -3675 2966 -3658
rect 2908 -3709 2920 -3675
rect 2954 -3709 2966 -3675
rect 2908 -3803 2966 -3709
rect 3000 -3692 3050 -3599
rect 3084 -3571 3237 -3555
rect 3373 -3556 3443 -3444
rect 3533 -3342 3599 -3293
rect 3533 -3376 3549 -3342
rect 3583 -3376 3599 -3342
rect 3533 -3410 3599 -3376
rect 3533 -3444 3549 -3410
rect 3583 -3444 3599 -3410
rect 3533 -3460 3599 -3444
rect 3633 -3342 3702 -3327
rect 3633 -3376 3649 -3342
rect 3683 -3376 3702 -3342
rect 3633 -3410 3702 -3376
rect 3633 -3444 3649 -3410
rect 3683 -3444 3702 -3410
rect 3633 -3494 3702 -3444
rect 3084 -3605 3087 -3571
rect 3121 -3605 3237 -3571
rect 3084 -3621 3237 -3605
rect 3271 -3571 3443 -3556
rect 3508 -3528 3702 -3494
rect 3736 -3364 3794 -3293
rect 3736 -3398 3748 -3364
rect 3782 -3398 3794 -3364
rect 3736 -3457 3794 -3398
rect 3736 -3491 3748 -3457
rect 3782 -3491 3794 -3457
rect 3736 -3526 3794 -3491
rect 3828 -3335 4162 -3293
rect 3828 -3369 3846 -3335
rect 3880 -3369 4110 -3335
rect 4144 -3369 4162 -3335
rect 3828 -3437 4162 -3369
rect 3828 -3471 3846 -3437
rect 3880 -3471 4110 -3437
rect 4144 -3471 4162 -3437
rect 3828 -3511 4162 -3471
rect 4196 -3364 4254 -3293
rect 4196 -3398 4208 -3364
rect 4242 -3398 4254 -3364
rect 4196 -3457 4254 -3398
rect 4196 -3491 4208 -3457
rect 4242 -3491 4254 -3457
rect 3508 -3557 3578 -3528
rect 3271 -3605 3287 -3571
rect 3321 -3605 3443 -3571
rect 3271 -3606 3443 -3605
rect 3203 -3640 3237 -3621
rect 3203 -3674 3321 -3640
rect 3000 -3716 3081 -3692
rect 3000 -3750 3033 -3716
rect 3067 -3750 3081 -3716
rect 3000 -3769 3081 -3750
rect 3115 -3716 3181 -3700
rect 3115 -3750 3131 -3716
rect 3165 -3750 3181 -3716
rect 3115 -3803 3181 -3750
rect 3271 -3716 3321 -3674
rect 3271 -3750 3287 -3716
rect 3271 -3769 3321 -3750
rect 3373 -3716 3443 -3606
rect 3492 -3571 3578 -3557
rect 3492 -3605 3508 -3571
rect 3542 -3605 3578 -3571
rect 3612 -3565 3702 -3562
rect 3612 -3571 3630 -3565
rect 3612 -3605 3628 -3571
rect 3664 -3599 3702 -3565
rect 3662 -3605 3702 -3599
rect 3828 -3581 3978 -3511
rect 4196 -3526 4254 -3491
rect 4288 -3335 4990 -3293
rect 4288 -3369 4306 -3335
rect 4340 -3369 4938 -3335
rect 4972 -3369 4990 -3335
rect 4288 -3437 4990 -3369
rect 4288 -3471 4306 -3437
rect 4340 -3471 4938 -3437
rect 4972 -3471 4990 -3437
rect 4288 -3511 4990 -3471
rect 3492 -3615 3578 -3605
rect 3828 -3615 3848 -3581
rect 3882 -3615 3978 -3581
rect 4012 -3579 4108 -3545
rect 4142 -3579 4162 -3545
rect 3508 -3639 3578 -3615
rect 3508 -3673 3702 -3639
rect 4012 -3649 4162 -3579
rect 3373 -3750 3392 -3716
rect 3426 -3750 3443 -3716
rect 3373 -3769 3443 -3750
rect 3536 -3716 3602 -3707
rect 3536 -3750 3552 -3716
rect 3586 -3750 3602 -3716
rect 3536 -3803 3602 -3750
rect 3636 -3716 3702 -3673
rect 3636 -3750 3649 -3716
rect 3683 -3750 3702 -3716
rect 3636 -3769 3702 -3750
rect 3736 -3675 3794 -3658
rect 3736 -3709 3748 -3675
rect 3782 -3709 3794 -3675
rect 3736 -3803 3794 -3709
rect 3828 -3701 4162 -3649
rect 4288 -3579 4366 -3545
rect 4400 -3579 4465 -3545
rect 4499 -3579 4564 -3545
rect 4598 -3579 4618 -3545
rect 4288 -3649 4618 -3579
rect 4652 -3581 4990 -3511
rect 5024 -3364 5082 -3293
rect 5024 -3398 5036 -3364
rect 5070 -3398 5082 -3364
rect 5024 -3457 5082 -3398
rect 5024 -3491 5036 -3457
rect 5070 -3491 5082 -3457
rect 5024 -3526 5082 -3491
rect 5116 -3335 5450 -3293
rect 5116 -3369 5134 -3335
rect 5168 -3369 5398 -3335
rect 5432 -3369 5450 -3335
rect 5116 -3437 5450 -3369
rect 5116 -3471 5134 -3437
rect 5168 -3471 5398 -3437
rect 5432 -3471 5450 -3437
rect 5116 -3511 5450 -3471
rect 5484 -3364 5542 -3293
rect 5484 -3398 5496 -3364
rect 5530 -3398 5542 -3364
rect 5484 -3457 5542 -3398
rect 5484 -3491 5496 -3457
rect 5530 -3491 5542 -3457
rect 4652 -3615 4672 -3581
rect 4706 -3615 4775 -3581
rect 4809 -3615 4878 -3581
rect 4912 -3615 4990 -3581
rect 5116 -3581 5266 -3511
rect 5484 -3526 5542 -3491
rect 5576 -3343 5657 -3327
rect 5576 -3377 5609 -3343
rect 5643 -3377 5657 -3343
rect 5576 -3411 5657 -3377
rect 5576 -3445 5609 -3411
rect 5643 -3445 5657 -3411
rect 5576 -3482 5657 -3445
rect 5691 -3342 5757 -3293
rect 5691 -3376 5707 -3342
rect 5741 -3376 5757 -3342
rect 5691 -3410 5757 -3376
rect 5691 -3444 5707 -3410
rect 5741 -3444 5757 -3410
rect 5691 -3453 5757 -3444
rect 5847 -3343 5897 -3327
rect 5847 -3377 5863 -3343
rect 5847 -3411 5897 -3377
rect 5847 -3445 5863 -3411
rect 5116 -3615 5136 -3581
rect 5170 -3615 5266 -3581
rect 5300 -3579 5396 -3545
rect 5430 -3579 5450 -3545
rect 5300 -3649 5450 -3579
rect 3828 -3735 3846 -3701
rect 3880 -3735 4110 -3701
rect 4144 -3735 4162 -3701
rect 3828 -3803 4162 -3735
rect 4196 -3675 4254 -3658
rect 4196 -3709 4208 -3675
rect 4242 -3709 4254 -3675
rect 4196 -3803 4254 -3709
rect 4288 -3708 4990 -3649
rect 4288 -3742 4306 -3708
rect 4340 -3742 4938 -3708
rect 4972 -3742 4990 -3708
rect 4288 -3803 4990 -3742
rect 5024 -3675 5082 -3658
rect 5024 -3709 5036 -3675
rect 5070 -3709 5082 -3675
rect 5024 -3803 5082 -3709
rect 5116 -3701 5450 -3649
rect 5576 -3565 5626 -3482
rect 5847 -3487 5897 -3445
rect 5779 -3521 5897 -3487
rect 5949 -3342 6019 -3327
rect 5949 -3376 5967 -3342
rect 6001 -3376 6019 -3342
rect 5949 -3410 6019 -3376
rect 5949 -3444 5967 -3410
rect 6001 -3444 6019 -3410
rect 5779 -3555 5813 -3521
rect 5576 -3599 5590 -3565
rect 5624 -3599 5626 -3565
rect 5116 -3735 5134 -3701
rect 5168 -3735 5398 -3701
rect 5432 -3735 5450 -3701
rect 5116 -3803 5450 -3735
rect 5484 -3675 5542 -3658
rect 5484 -3709 5496 -3675
rect 5530 -3709 5542 -3675
rect 5484 -3803 5542 -3709
rect 5576 -3692 5626 -3599
rect 5660 -3571 5813 -3555
rect 5949 -3556 6019 -3444
rect 6109 -3342 6175 -3293
rect 6109 -3376 6125 -3342
rect 6159 -3376 6175 -3342
rect 6109 -3410 6175 -3376
rect 6109 -3444 6125 -3410
rect 6159 -3444 6175 -3410
rect 6109 -3460 6175 -3444
rect 6209 -3342 6278 -3327
rect 6209 -3376 6225 -3342
rect 6259 -3376 6278 -3342
rect 6209 -3410 6278 -3376
rect 6209 -3444 6225 -3410
rect 6259 -3444 6278 -3410
rect 6209 -3494 6278 -3444
rect 5660 -3605 5663 -3571
rect 5697 -3605 5813 -3571
rect 5660 -3621 5813 -3605
rect 5847 -3571 6019 -3556
rect 6084 -3528 6278 -3494
rect 6312 -3364 6370 -3293
rect 6312 -3398 6324 -3364
rect 6358 -3398 6370 -3364
rect 6312 -3457 6370 -3398
rect 6312 -3491 6324 -3457
rect 6358 -3491 6370 -3457
rect 6312 -3526 6370 -3491
rect 6404 -3335 6738 -3293
rect 6404 -3369 6422 -3335
rect 6456 -3369 6686 -3335
rect 6720 -3369 6738 -3335
rect 6404 -3437 6738 -3369
rect 6404 -3471 6422 -3437
rect 6456 -3471 6686 -3437
rect 6720 -3471 6738 -3437
rect 6404 -3511 6738 -3471
rect 6772 -3364 6830 -3293
rect 6772 -3398 6784 -3364
rect 6818 -3398 6830 -3364
rect 6772 -3457 6830 -3398
rect 6772 -3491 6784 -3457
rect 6818 -3491 6830 -3457
rect 6084 -3557 6154 -3528
rect 5847 -3605 5863 -3571
rect 5897 -3605 6019 -3571
rect 5847 -3606 6019 -3605
rect 5779 -3640 5813 -3621
rect 5779 -3674 5897 -3640
rect 5576 -3716 5657 -3692
rect 5576 -3750 5609 -3716
rect 5643 -3750 5657 -3716
rect 5576 -3769 5657 -3750
rect 5691 -3716 5757 -3700
rect 5691 -3750 5707 -3716
rect 5741 -3750 5757 -3716
rect 5691 -3803 5757 -3750
rect 5847 -3716 5897 -3674
rect 5847 -3750 5863 -3716
rect 5847 -3769 5897 -3750
rect 5949 -3716 6019 -3606
rect 6068 -3571 6154 -3557
rect 6068 -3605 6084 -3571
rect 6118 -3605 6154 -3571
rect 6188 -3565 6278 -3562
rect 6188 -3605 6204 -3565
rect 6238 -3605 6278 -3565
rect 6404 -3581 6554 -3511
rect 6772 -3526 6830 -3491
rect 6864 -3335 7566 -3293
rect 6864 -3369 6882 -3335
rect 6916 -3369 7514 -3335
rect 7548 -3369 7566 -3335
rect 6864 -3437 7566 -3369
rect 6864 -3471 6882 -3437
rect 6916 -3471 7514 -3437
rect 7548 -3471 7566 -3437
rect 6864 -3511 7566 -3471
rect 6068 -3615 6154 -3605
rect 6404 -3615 6424 -3581
rect 6458 -3615 6554 -3581
rect 6588 -3579 6684 -3545
rect 6718 -3579 6738 -3545
rect 6084 -3639 6154 -3615
rect 6084 -3673 6278 -3639
rect 6588 -3649 6738 -3579
rect 5949 -3750 5968 -3716
rect 6002 -3750 6019 -3716
rect 5949 -3769 6019 -3750
rect 6112 -3716 6178 -3707
rect 6112 -3750 6128 -3716
rect 6162 -3750 6178 -3716
rect 6112 -3803 6178 -3750
rect 6212 -3716 6278 -3673
rect 6212 -3750 6225 -3716
rect 6259 -3750 6278 -3716
rect 6212 -3769 6278 -3750
rect 6312 -3675 6370 -3658
rect 6312 -3709 6324 -3675
rect 6358 -3709 6370 -3675
rect 6312 -3803 6370 -3709
rect 6404 -3701 6738 -3649
rect 6864 -3579 6942 -3545
rect 6976 -3579 7041 -3545
rect 7075 -3579 7140 -3545
rect 7174 -3579 7194 -3545
rect 6864 -3649 7194 -3579
rect 7228 -3581 7566 -3511
rect 7600 -3364 7658 -3293
rect 7600 -3398 7612 -3364
rect 7646 -3398 7658 -3364
rect 7600 -3457 7658 -3398
rect 7600 -3491 7612 -3457
rect 7646 -3491 7658 -3457
rect 7600 -3526 7658 -3491
rect 7692 -3335 8026 -3293
rect 7692 -3369 7710 -3335
rect 7744 -3369 7974 -3335
rect 8008 -3369 8026 -3335
rect 7692 -3437 8026 -3369
rect 7692 -3471 7710 -3437
rect 7744 -3471 7974 -3437
rect 8008 -3471 8026 -3437
rect 7692 -3511 8026 -3471
rect 8060 -3364 8118 -3293
rect 8060 -3398 8072 -3364
rect 8106 -3398 8118 -3364
rect 8060 -3457 8118 -3398
rect 8060 -3491 8072 -3457
rect 8106 -3491 8118 -3457
rect 7228 -3615 7248 -3581
rect 7282 -3615 7351 -3581
rect 7385 -3615 7454 -3581
rect 7488 -3615 7566 -3581
rect 7692 -3581 7842 -3511
rect 8060 -3526 8118 -3491
rect 8152 -3343 8233 -3327
rect 8152 -3377 8185 -3343
rect 8219 -3377 8233 -3343
rect 8152 -3411 8233 -3377
rect 8152 -3445 8185 -3411
rect 8219 -3445 8233 -3411
rect 8152 -3482 8233 -3445
rect 8267 -3342 8333 -3293
rect 8267 -3376 8283 -3342
rect 8317 -3376 8333 -3342
rect 8267 -3410 8333 -3376
rect 8267 -3444 8283 -3410
rect 8317 -3444 8333 -3410
rect 8267 -3453 8333 -3444
rect 8423 -3343 8473 -3327
rect 8423 -3377 8439 -3343
rect 8423 -3411 8473 -3377
rect 8423 -3445 8439 -3411
rect 7692 -3615 7712 -3581
rect 7746 -3615 7842 -3581
rect 7876 -3579 7972 -3545
rect 8006 -3579 8026 -3545
rect 7876 -3649 8026 -3579
rect 6404 -3735 6422 -3701
rect 6456 -3735 6686 -3701
rect 6720 -3735 6738 -3701
rect 6404 -3803 6738 -3735
rect 6772 -3675 6830 -3658
rect 6772 -3709 6784 -3675
rect 6818 -3709 6830 -3675
rect 6772 -3803 6830 -3709
rect 6864 -3708 7566 -3649
rect 6864 -3742 6882 -3708
rect 6916 -3742 7514 -3708
rect 7548 -3742 7566 -3708
rect 6864 -3803 7566 -3742
rect 7600 -3675 7658 -3658
rect 7600 -3709 7612 -3675
rect 7646 -3709 7658 -3675
rect 7600 -3803 7658 -3709
rect 7692 -3701 8026 -3649
rect 8152 -3565 8202 -3482
rect 8423 -3487 8473 -3445
rect 8355 -3521 8473 -3487
rect 8525 -3342 8595 -3327
rect 8525 -3376 8543 -3342
rect 8577 -3376 8595 -3342
rect 8525 -3410 8595 -3376
rect 8525 -3444 8543 -3410
rect 8577 -3444 8595 -3410
rect 8355 -3555 8389 -3521
rect 8152 -3599 8164 -3565
rect 8198 -3599 8202 -3565
rect 7692 -3735 7710 -3701
rect 7744 -3735 7974 -3701
rect 8008 -3735 8026 -3701
rect 7692 -3803 8026 -3735
rect 8060 -3675 8118 -3658
rect 8060 -3709 8072 -3675
rect 8106 -3709 8118 -3675
rect 8060 -3803 8118 -3709
rect 8152 -3692 8202 -3599
rect 8236 -3571 8389 -3555
rect 8525 -3556 8595 -3444
rect 8685 -3342 8751 -3293
rect 8685 -3376 8701 -3342
rect 8735 -3376 8751 -3342
rect 8685 -3410 8751 -3376
rect 8685 -3444 8701 -3410
rect 8735 -3444 8751 -3410
rect 8685 -3460 8751 -3444
rect 8785 -3342 8854 -3327
rect 8785 -3376 8801 -3342
rect 8835 -3376 8854 -3342
rect 8785 -3410 8854 -3376
rect 8785 -3444 8801 -3410
rect 8835 -3444 8854 -3410
rect 8785 -3494 8854 -3444
rect 8236 -3605 8239 -3571
rect 8273 -3605 8389 -3571
rect 8236 -3621 8389 -3605
rect 8423 -3571 8595 -3556
rect 8660 -3528 8854 -3494
rect 8888 -3364 8946 -3293
rect 8888 -3398 8900 -3364
rect 8934 -3398 8946 -3364
rect 8888 -3457 8946 -3398
rect 8888 -3491 8900 -3457
rect 8934 -3491 8946 -3457
rect 8888 -3526 8946 -3491
rect 8980 -3335 9314 -3293
rect 8980 -3369 8998 -3335
rect 9032 -3369 9262 -3335
rect 9296 -3369 9314 -3335
rect 8980 -3437 9314 -3369
rect 8980 -3471 8998 -3437
rect 9032 -3471 9262 -3437
rect 9296 -3471 9314 -3437
rect 8980 -3511 9314 -3471
rect 9348 -3364 9406 -3293
rect 9348 -3398 9360 -3364
rect 9394 -3398 9406 -3364
rect 9348 -3457 9406 -3398
rect 9348 -3491 9360 -3457
rect 9394 -3491 9406 -3457
rect 8660 -3557 8730 -3528
rect 8423 -3605 8439 -3571
rect 8473 -3605 8595 -3571
rect 8423 -3606 8595 -3605
rect 8355 -3640 8389 -3621
rect 8355 -3674 8473 -3640
rect 8152 -3716 8233 -3692
rect 8152 -3750 8185 -3716
rect 8219 -3750 8233 -3716
rect 8152 -3769 8233 -3750
rect 8267 -3716 8333 -3700
rect 8267 -3750 8283 -3716
rect 8317 -3750 8333 -3716
rect 8267 -3803 8333 -3750
rect 8423 -3716 8473 -3674
rect 8423 -3750 8439 -3716
rect 8423 -3769 8473 -3750
rect 8525 -3716 8595 -3606
rect 8644 -3571 8730 -3557
rect 8644 -3605 8660 -3571
rect 8694 -3605 8730 -3571
rect 8764 -3565 8854 -3562
rect 8764 -3599 8778 -3565
rect 8812 -3571 8854 -3565
rect 8764 -3605 8780 -3599
rect 8814 -3605 8854 -3571
rect 8980 -3581 9130 -3511
rect 9348 -3526 9406 -3491
rect 9440 -3335 10142 -3293
rect 9440 -3369 9458 -3335
rect 9492 -3369 10090 -3335
rect 10124 -3369 10142 -3335
rect 9440 -3437 10142 -3369
rect 9440 -3471 9458 -3437
rect 9492 -3471 10090 -3437
rect 10124 -3471 10142 -3437
rect 9440 -3511 10142 -3471
rect 8644 -3615 8730 -3605
rect 8980 -3615 9000 -3581
rect 9034 -3615 9130 -3581
rect 9164 -3579 9260 -3545
rect 9294 -3579 9314 -3545
rect 8660 -3639 8730 -3615
rect 8660 -3673 8854 -3639
rect 9164 -3649 9314 -3579
rect 8525 -3750 8544 -3716
rect 8578 -3750 8595 -3716
rect 8525 -3769 8595 -3750
rect 8688 -3716 8754 -3707
rect 8688 -3750 8704 -3716
rect 8738 -3750 8754 -3716
rect 8688 -3803 8754 -3750
rect 8788 -3716 8854 -3673
rect 8788 -3750 8801 -3716
rect 8835 -3750 8854 -3716
rect 8788 -3769 8854 -3750
rect 8888 -3675 8946 -3658
rect 8888 -3709 8900 -3675
rect 8934 -3709 8946 -3675
rect 8888 -3803 8946 -3709
rect 8980 -3701 9314 -3649
rect 9440 -3579 9518 -3545
rect 9552 -3579 9617 -3545
rect 9651 -3579 9716 -3545
rect 9750 -3579 9770 -3545
rect 9440 -3649 9770 -3579
rect 9804 -3581 10142 -3511
rect 10176 -3364 10234 -3293
rect 10176 -3398 10188 -3364
rect 10222 -3398 10234 -3364
rect 10176 -3457 10234 -3398
rect 10176 -3491 10188 -3457
rect 10222 -3491 10234 -3457
rect 10176 -3526 10234 -3491
rect 10360 -3335 10694 -3293
rect 10360 -3369 10378 -3335
rect 10412 -3369 10642 -3335
rect 10676 -3369 10694 -3335
rect 10360 -3437 10694 -3369
rect 10360 -3471 10378 -3437
rect 10412 -3471 10642 -3437
rect 10676 -3471 10694 -3437
rect 10360 -3511 10694 -3471
rect 10728 -3343 10809 -3327
rect 10728 -3377 10761 -3343
rect 10795 -3377 10809 -3343
rect 10728 -3411 10809 -3377
rect 10728 -3445 10761 -3411
rect 10795 -3445 10809 -3411
rect 10728 -3482 10809 -3445
rect 10843 -3342 10909 -3293
rect 10843 -3376 10859 -3342
rect 10893 -3376 10909 -3342
rect 10843 -3410 10909 -3376
rect 10843 -3444 10859 -3410
rect 10893 -3444 10909 -3410
rect 10843 -3453 10909 -3444
rect 10999 -3343 11049 -3327
rect 10999 -3377 11015 -3343
rect 10999 -3411 11049 -3377
rect 10999 -3445 11015 -3411
rect 9804 -3615 9824 -3581
rect 9858 -3615 9927 -3581
rect 9961 -3615 10030 -3581
rect 10064 -3615 10142 -3581
rect 10360 -3581 10510 -3511
rect 10360 -3615 10380 -3581
rect 10414 -3615 10510 -3581
rect 10544 -3579 10640 -3545
rect 10674 -3579 10694 -3545
rect 10544 -3649 10694 -3579
rect 8980 -3735 8998 -3701
rect 9032 -3735 9262 -3701
rect 9296 -3735 9314 -3701
rect 8980 -3803 9314 -3735
rect 9348 -3675 9406 -3658
rect 9348 -3709 9360 -3675
rect 9394 -3709 9406 -3675
rect 9348 -3803 9406 -3709
rect 9440 -3708 10142 -3649
rect 9440 -3742 9458 -3708
rect 9492 -3742 10090 -3708
rect 10124 -3742 10142 -3708
rect 9440 -3803 10142 -3742
rect 10176 -3675 10234 -3658
rect 10176 -3709 10188 -3675
rect 10222 -3709 10234 -3675
rect 10176 -3803 10234 -3709
rect 10360 -3701 10694 -3649
rect 10360 -3735 10378 -3701
rect 10412 -3735 10642 -3701
rect 10676 -3735 10694 -3701
rect 10360 -3803 10694 -3735
rect 10728 -3568 10778 -3482
rect 10999 -3487 11049 -3445
rect 10931 -3521 11049 -3487
rect 11101 -3342 11171 -3327
rect 11101 -3376 11119 -3342
rect 11153 -3376 11171 -3342
rect 11101 -3410 11171 -3376
rect 11101 -3444 11119 -3410
rect 11153 -3444 11171 -3410
rect 10931 -3555 10965 -3521
rect 10728 -3602 10735 -3568
rect 10769 -3602 10778 -3568
rect 10728 -3692 10778 -3602
rect 10812 -3571 10965 -3555
rect 11101 -3556 11171 -3444
rect 11261 -3342 11327 -3293
rect 11261 -3376 11277 -3342
rect 11311 -3376 11327 -3342
rect 11261 -3410 11327 -3376
rect 11261 -3444 11277 -3410
rect 11311 -3444 11327 -3410
rect 11261 -3460 11327 -3444
rect 11361 -3342 11430 -3327
rect 11361 -3376 11377 -3342
rect 11411 -3376 11430 -3342
rect 11361 -3410 11430 -3376
rect 11361 -3444 11377 -3410
rect 11411 -3444 11430 -3410
rect 11361 -3494 11430 -3444
rect 10812 -3605 10815 -3571
rect 10849 -3605 10965 -3571
rect 10812 -3621 10965 -3605
rect 10999 -3571 11171 -3556
rect 11236 -3528 11430 -3494
rect 11464 -3364 11522 -3293
rect 11464 -3398 11476 -3364
rect 11510 -3398 11522 -3364
rect 11464 -3457 11522 -3398
rect 11464 -3491 11476 -3457
rect 11510 -3491 11522 -3457
rect 11464 -3526 11522 -3491
rect 11648 -3335 11982 -3293
rect 11648 -3369 11666 -3335
rect 11700 -3369 11930 -3335
rect 11964 -3369 11982 -3335
rect 11648 -3437 11982 -3369
rect 11648 -3471 11666 -3437
rect 11700 -3471 11930 -3437
rect 11964 -3471 11982 -3437
rect 11648 -3511 11982 -3471
rect 13488 -3364 13546 -3293
rect 13488 -3398 13500 -3364
rect 13534 -3398 13546 -3364
rect 13488 -3457 13546 -3398
rect 13488 -3491 13500 -3457
rect 13534 -3491 13546 -3457
rect 11236 -3557 11306 -3528
rect 10999 -3605 11015 -3571
rect 11049 -3605 11171 -3571
rect 10999 -3606 11171 -3605
rect 10931 -3640 10965 -3621
rect 10931 -3674 11049 -3640
rect 10728 -3716 10809 -3692
rect 10728 -3750 10761 -3716
rect 10795 -3750 10809 -3716
rect 10728 -3769 10809 -3750
rect 10843 -3716 10909 -3700
rect 10843 -3750 10859 -3716
rect 10893 -3750 10909 -3716
rect 10843 -3803 10909 -3750
rect 10999 -3716 11049 -3674
rect 10999 -3750 11015 -3716
rect 10999 -3769 11049 -3750
rect 11101 -3716 11171 -3606
rect 11220 -3571 11306 -3557
rect 11220 -3605 11236 -3571
rect 11270 -3605 11306 -3571
rect 11340 -3567 11430 -3562
rect 11340 -3571 11383 -3567
rect 11340 -3605 11356 -3571
rect 11417 -3601 11430 -3567
rect 11390 -3605 11430 -3601
rect 11648 -3581 11798 -3511
rect 13488 -3526 13546 -3491
rect 13581 -3335 14650 -3293
rect 13581 -3369 13598 -3335
rect 13632 -3369 14598 -3335
rect 14632 -3369 14650 -3335
rect 13581 -3437 14650 -3369
rect 13581 -3471 13598 -3437
rect 13632 -3471 14598 -3437
rect 14632 -3471 14650 -3437
rect 13581 -3511 14650 -3471
rect 14684 -3364 14742 -3293
rect 14684 -3398 14696 -3364
rect 14730 -3398 14742 -3364
rect 14684 -3457 14742 -3398
rect 14684 -3491 14696 -3457
rect 14730 -3491 14742 -3457
rect 11220 -3615 11306 -3605
rect 11648 -3615 11668 -3581
rect 11702 -3615 11798 -3581
rect 11832 -3579 11928 -3545
rect 11962 -3579 11982 -3545
rect 11236 -3639 11306 -3615
rect 11236 -3673 11430 -3639
rect 11832 -3649 11982 -3579
rect 13581 -3581 14100 -3511
rect 14684 -3526 14742 -3491
rect 14777 -3335 15846 -3293
rect 14777 -3369 14794 -3335
rect 14828 -3369 15794 -3335
rect 15828 -3369 15846 -3335
rect 14777 -3437 15846 -3369
rect 14777 -3471 14794 -3437
rect 14828 -3471 15794 -3437
rect 15828 -3471 15846 -3437
rect 14777 -3511 15846 -3471
rect 15880 -3364 15938 -3293
rect 15880 -3398 15892 -3364
rect 15926 -3398 15938 -3364
rect 15880 -3457 15938 -3398
rect 15880 -3491 15892 -3457
rect 15926 -3491 15938 -3457
rect 13581 -3615 13662 -3581
rect 13696 -3615 13790 -3581
rect 13824 -3615 13918 -3581
rect 13952 -3615 14046 -3581
rect 14080 -3615 14100 -3581
rect 14134 -3579 14154 -3545
rect 14188 -3579 14282 -3545
rect 14316 -3579 14410 -3545
rect 14444 -3579 14538 -3545
rect 14572 -3579 14650 -3545
rect 14134 -3649 14650 -3579
rect 14777 -3581 15296 -3511
rect 15880 -3526 15938 -3491
rect 15972 -3335 16674 -3293
rect 15972 -3369 15990 -3335
rect 16024 -3369 16622 -3335
rect 16656 -3369 16674 -3335
rect 15972 -3437 16674 -3369
rect 15972 -3471 15990 -3437
rect 16024 -3471 16622 -3437
rect 16656 -3471 16674 -3437
rect 15972 -3511 16674 -3471
rect 14777 -3615 14858 -3581
rect 14892 -3615 14986 -3581
rect 15020 -3615 15114 -3581
rect 15148 -3615 15242 -3581
rect 15276 -3615 15296 -3581
rect 15330 -3579 15350 -3545
rect 15384 -3579 15478 -3545
rect 15512 -3579 15606 -3545
rect 15640 -3579 15734 -3545
rect 15768 -3579 15846 -3545
rect 15330 -3649 15846 -3579
rect 15972 -3581 16310 -3511
rect 15972 -3615 16050 -3581
rect 16084 -3615 16153 -3581
rect 16187 -3615 16256 -3581
rect 16290 -3615 16310 -3581
rect 16344 -3579 16364 -3545
rect 16398 -3579 16463 -3545
rect 16497 -3579 16562 -3545
rect 16596 -3579 16674 -3545
rect 16344 -3649 16674 -3579
rect 11101 -3750 11120 -3716
rect 11154 -3750 11171 -3716
rect 11101 -3769 11171 -3750
rect 11264 -3716 11330 -3707
rect 11264 -3750 11280 -3716
rect 11314 -3750 11330 -3716
rect 11264 -3803 11330 -3750
rect 11364 -3716 11430 -3673
rect 11364 -3750 11377 -3716
rect 11411 -3750 11430 -3716
rect 11364 -3769 11430 -3750
rect 11464 -3675 11522 -3658
rect 11464 -3709 11476 -3675
rect 11510 -3709 11522 -3675
rect 11464 -3803 11522 -3709
rect 11648 -3701 11982 -3649
rect 11648 -3735 11666 -3701
rect 11700 -3735 11930 -3701
rect 11964 -3735 11982 -3701
rect 11648 -3803 11982 -3735
rect 13488 -3675 13546 -3658
rect 13488 -3709 13500 -3675
rect 13534 -3709 13546 -3675
rect 13488 -3803 13546 -3709
rect 13581 -3708 14650 -3649
rect 13581 -3742 13598 -3708
rect 13632 -3742 14598 -3708
rect 14632 -3742 14650 -3708
rect 13581 -3803 14650 -3742
rect 14684 -3675 14742 -3658
rect 14684 -3709 14696 -3675
rect 14730 -3709 14742 -3675
rect 14684 -3803 14742 -3709
rect 14777 -3708 15846 -3649
rect 14777 -3742 14794 -3708
rect 14828 -3742 15794 -3708
rect 15828 -3742 15846 -3708
rect 14777 -3803 15846 -3742
rect 15880 -3675 15938 -3658
rect 15880 -3709 15892 -3675
rect 15926 -3709 15938 -3675
rect 15880 -3803 15938 -3709
rect 15972 -3708 16674 -3649
rect 15972 -3742 15990 -3708
rect 16024 -3742 16622 -3708
rect 16656 -3742 16674 -3708
rect 15972 -3803 16674 -3742
rect -2997 -3837 -2968 -3803
rect -2934 -3837 -2876 -3803
rect -2842 -3837 -2784 -3803
rect -2750 -3837 -2692 -3803
rect -2658 -3837 -2600 -3803
rect -2566 -3837 -2508 -3803
rect -2474 -3837 -2416 -3803
rect -2382 -3837 -2324 -3803
rect -2290 -3837 -2232 -3803
rect -2198 -3837 -2140 -3803
rect -2106 -3837 -2048 -3803
rect -2014 -3837 -1956 -3803
rect -1922 -3837 -1864 -3803
rect -1830 -3837 -1772 -3803
rect -1738 -3837 -1680 -3803
rect -1646 -3837 -1588 -3803
rect -1554 -3837 -1496 -3803
rect -1462 -3837 -1404 -3803
rect -1370 -3837 -1312 -3803
rect -1278 -3837 -1220 -3803
rect -1186 -3837 -1128 -3803
rect -1094 -3837 -1036 -3803
rect -1002 -3837 -944 -3803
rect -910 -3837 -852 -3803
rect -818 -3837 -760 -3803
rect -726 -3837 -668 -3803
rect -634 -3837 -576 -3803
rect -542 -3837 -484 -3803
rect -450 -3837 -392 -3803
rect -358 -3837 -300 -3803
rect -266 -3837 -208 -3803
rect -174 -3837 -116 -3803
rect -82 -3837 -24 -3803
rect 10 -3837 68 -3803
rect 102 -3837 160 -3803
rect 194 -3837 252 -3803
rect 286 -3837 344 -3803
rect 378 -3837 436 -3803
rect 470 -3837 528 -3803
rect 562 -3837 620 -3803
rect 654 -3837 712 -3803
rect 746 -3837 804 -3803
rect 838 -3837 896 -3803
rect 930 -3837 988 -3803
rect 1022 -3837 1080 -3803
rect 1114 -3837 1172 -3803
rect 1206 -3837 1264 -3803
rect 1298 -3837 1356 -3803
rect 1390 -3837 1448 -3803
rect 1482 -3837 1540 -3803
rect 1574 -3837 1632 -3803
rect 1666 -3837 1724 -3803
rect 1758 -3837 1816 -3803
rect 1850 -3837 1908 -3803
rect 1942 -3837 2000 -3803
rect 2034 -3837 2092 -3803
rect 2126 -3837 2184 -3803
rect 2218 -3837 2276 -3803
rect 2310 -3837 2368 -3803
rect 2402 -3837 2460 -3803
rect 2494 -3837 2552 -3803
rect 2586 -3837 2644 -3803
rect 2678 -3837 2736 -3803
rect 2770 -3837 2828 -3803
rect 2862 -3837 2920 -3803
rect 2954 -3837 3012 -3803
rect 3046 -3837 3104 -3803
rect 3138 -3837 3196 -3803
rect 3230 -3837 3288 -3803
rect 3322 -3837 3380 -3803
rect 3414 -3837 3472 -3803
rect 3506 -3837 3564 -3803
rect 3598 -3837 3656 -3803
rect 3690 -3837 3748 -3803
rect 3782 -3837 3840 -3803
rect 3874 -3837 3932 -3803
rect 3966 -3837 4024 -3803
rect 4058 -3837 4116 -3803
rect 4150 -3837 4208 -3803
rect 4242 -3837 4300 -3803
rect 4334 -3837 4392 -3803
rect 4426 -3837 4484 -3803
rect 4518 -3837 4576 -3803
rect 4610 -3837 4668 -3803
rect 4702 -3837 4760 -3803
rect 4794 -3837 4852 -3803
rect 4886 -3837 4944 -3803
rect 4978 -3837 5036 -3803
rect 5070 -3837 5128 -3803
rect 5162 -3837 5220 -3803
rect 5254 -3837 5312 -3803
rect 5346 -3837 5404 -3803
rect 5438 -3837 5496 -3803
rect 5530 -3837 5588 -3803
rect 5622 -3837 5680 -3803
rect 5714 -3837 5772 -3803
rect 5806 -3837 5864 -3803
rect 5898 -3837 5956 -3803
rect 5990 -3837 6048 -3803
rect 6082 -3837 6140 -3803
rect 6174 -3837 6232 -3803
rect 6266 -3837 6324 -3803
rect 6358 -3837 6416 -3803
rect 6450 -3837 6508 -3803
rect 6542 -3837 6600 -3803
rect 6634 -3837 6692 -3803
rect 6726 -3837 6784 -3803
rect 6818 -3837 6876 -3803
rect 6910 -3837 6968 -3803
rect 7002 -3837 7060 -3803
rect 7094 -3837 7152 -3803
rect 7186 -3837 7244 -3803
rect 7278 -3837 7336 -3803
rect 7370 -3837 7428 -3803
rect 7462 -3837 7520 -3803
rect 7554 -3837 7612 -3803
rect 7646 -3837 7704 -3803
rect 7738 -3837 7796 -3803
rect 7830 -3837 7888 -3803
rect 7922 -3837 7980 -3803
rect 8014 -3837 8072 -3803
rect 8106 -3837 8164 -3803
rect 8198 -3837 8256 -3803
rect 8290 -3837 8348 -3803
rect 8382 -3837 8440 -3803
rect 8474 -3837 8532 -3803
rect 8566 -3837 8624 -3803
rect 8658 -3837 8716 -3803
rect 8750 -3837 8808 -3803
rect 8842 -3837 8900 -3803
rect 8934 -3837 8992 -3803
rect 9026 -3837 9084 -3803
rect 9118 -3837 9176 -3803
rect 9210 -3837 9268 -3803
rect 9302 -3837 9360 -3803
rect 9394 -3837 9452 -3803
rect 9486 -3837 9544 -3803
rect 9578 -3837 9636 -3803
rect 9670 -3837 9728 -3803
rect 9762 -3837 9820 -3803
rect 9854 -3837 9912 -3803
rect 9946 -3837 10004 -3803
rect 10038 -3837 10096 -3803
rect 10130 -3837 10188 -3803
rect 10222 -3837 10280 -3803
rect 10314 -3837 10372 -3803
rect 10406 -3837 10464 -3803
rect 10498 -3837 10556 -3803
rect 10590 -3837 10648 -3803
rect 10682 -3837 10740 -3803
rect 10774 -3837 10832 -3803
rect 10866 -3837 10924 -3803
rect 10958 -3837 11016 -3803
rect 11050 -3837 11108 -3803
rect 11142 -3837 11200 -3803
rect 11234 -3837 11292 -3803
rect 11326 -3837 11384 -3803
rect 11418 -3837 11476 -3803
rect 11510 -3837 11568 -3803
rect 11602 -3837 11660 -3803
rect 11694 -3837 11752 -3803
rect 11786 -3837 11844 -3803
rect 11878 -3837 11936 -3803
rect 11970 -3837 12028 -3803
rect 12062 -3837 12120 -3803
rect 12154 -3837 12212 -3803
rect 12246 -3837 12304 -3803
rect 12338 -3837 12396 -3803
rect 12430 -3837 12488 -3803
rect 12522 -3837 12580 -3803
rect 12614 -3837 12672 -3803
rect 12706 -3837 12764 -3803
rect 12798 -3837 12856 -3803
rect 12890 -3837 12948 -3803
rect 12982 -3837 13040 -3803
rect 13074 -3837 13132 -3803
rect 13166 -3837 13224 -3803
rect 13258 -3837 13316 -3803
rect 13350 -3837 13408 -3803
rect 13442 -3837 13500 -3803
rect 13534 -3837 13592 -3803
rect 13626 -3837 13684 -3803
rect 13718 -3837 13776 -3803
rect 13810 -3837 13868 -3803
rect 13902 -3837 13960 -3803
rect 13994 -3837 14052 -3803
rect 14086 -3837 14144 -3803
rect 14178 -3837 14236 -3803
rect 14270 -3837 14328 -3803
rect 14362 -3837 14420 -3803
rect 14454 -3837 14512 -3803
rect 14546 -3837 14604 -3803
rect 14638 -3837 14696 -3803
rect 14730 -3837 14788 -3803
rect 14822 -3837 14880 -3803
rect 14914 -3837 14972 -3803
rect 15006 -3837 15064 -3803
rect 15098 -3837 15156 -3803
rect 15190 -3837 15248 -3803
rect 15282 -3837 15340 -3803
rect 15374 -3837 15432 -3803
rect 15466 -3837 15524 -3803
rect 15558 -3837 15616 -3803
rect 15650 -3837 15708 -3803
rect 15742 -3837 15800 -3803
rect 15834 -3837 15892 -3803
rect 15926 -3837 15984 -3803
rect 16018 -3837 16076 -3803
rect 16110 -3837 16168 -3803
rect 16202 -3837 16260 -3803
rect 16294 -3837 16352 -3803
rect 16386 -3837 16444 -3803
rect 16478 -3837 16536 -3803
rect 16570 -3837 16628 -3803
rect 16662 -3837 16691 -3803
rect -2980 -3898 -2278 -3837
rect -2980 -3932 -2962 -3898
rect -2928 -3932 -2330 -3898
rect -2296 -3932 -2278 -3898
rect -2980 -3991 -2278 -3932
rect -2244 -3931 -2186 -3837
rect -2244 -3965 -2232 -3931
rect -2198 -3965 -2186 -3931
rect -2244 -3982 -2186 -3965
rect -1600 -3898 -898 -3837
rect -1600 -3932 -1582 -3898
rect -1548 -3932 -950 -3898
rect -916 -3932 -898 -3898
rect -2980 -4059 -2902 -4025
rect -2868 -4059 -2799 -4025
rect -2765 -4059 -2696 -4025
rect -2662 -4059 -2642 -4025
rect -2980 -4129 -2642 -4059
rect -2608 -4061 -2278 -3991
rect -2608 -4095 -2588 -4061
rect -2554 -4095 -2489 -4061
rect -2455 -4095 -2390 -4061
rect -2356 -4095 -2278 -4061
rect -1600 -3991 -898 -3932
rect -864 -3898 -162 -3837
rect -864 -3932 -846 -3898
rect -812 -3932 -214 -3898
rect -180 -3932 -162 -3898
rect -864 -3991 -162 -3932
rect -128 -3931 -70 -3837
rect -128 -3965 -116 -3931
rect -82 -3965 -70 -3931
rect -128 -3982 -70 -3965
rect -36 -3905 298 -3837
rect -36 -3939 -18 -3905
rect 16 -3939 246 -3905
rect 280 -3939 298 -3905
rect -36 -3991 298 -3939
rect 332 -3931 390 -3837
rect 332 -3965 344 -3931
rect 378 -3965 390 -3931
rect 332 -3982 390 -3965
rect 424 -3890 490 -3871
rect 424 -3924 443 -3890
rect 477 -3924 490 -3890
rect 424 -3967 490 -3924
rect 524 -3890 590 -3837
rect 524 -3924 540 -3890
rect 574 -3924 590 -3890
rect 524 -3933 590 -3924
rect 683 -3890 753 -3871
rect 683 -3924 700 -3890
rect 734 -3924 753 -3890
rect -1600 -4061 -1270 -3991
rect -1600 -4095 -1522 -4061
rect -1488 -4095 -1423 -4061
rect -1389 -4095 -1324 -4061
rect -1290 -4095 -1270 -4061
rect -1236 -4059 -1216 -4025
rect -1182 -4059 -1113 -4025
rect -1079 -4059 -1010 -4025
rect -976 -4059 -898 -4025
rect -2980 -4169 -2278 -4129
rect -2980 -4203 -2962 -4169
rect -2928 -4203 -2330 -4169
rect -2296 -4203 -2278 -4169
rect -2980 -4271 -2278 -4203
rect -2980 -4305 -2962 -4271
rect -2928 -4305 -2330 -4271
rect -2296 -4305 -2278 -4271
rect -2980 -4347 -2278 -4305
rect -2244 -4149 -2186 -4114
rect -1236 -4129 -898 -4059
rect -864 -4061 -534 -3991
rect -864 -4095 -786 -4061
rect -752 -4095 -687 -4061
rect -653 -4095 -588 -4061
rect -554 -4095 -534 -4061
rect -500 -4059 -480 -4025
rect -446 -4059 -377 -4025
rect -343 -4059 -274 -4025
rect -240 -4059 -162 -4025
rect -500 -4129 -162 -4059
rect -36 -4059 -16 -4025
rect 18 -4059 114 -4025
rect -2244 -4183 -2232 -4149
rect -2198 -4183 -2186 -4149
rect -2244 -4242 -2186 -4183
rect -2244 -4276 -2232 -4242
rect -2198 -4276 -2186 -4242
rect -2244 -4347 -2186 -4276
rect -1600 -4169 -898 -4129
rect -1600 -4203 -1582 -4169
rect -1548 -4203 -950 -4169
rect -916 -4203 -898 -4169
rect -1600 -4271 -898 -4203
rect -1600 -4305 -1582 -4271
rect -1548 -4305 -950 -4271
rect -916 -4305 -898 -4271
rect -1600 -4347 -898 -4305
rect -864 -4169 -162 -4129
rect -864 -4203 -846 -4169
rect -812 -4203 -214 -4169
rect -180 -4203 -162 -4169
rect -864 -4271 -162 -4203
rect -864 -4305 -846 -4271
rect -812 -4305 -214 -4271
rect -180 -4305 -162 -4271
rect -864 -4347 -162 -4305
rect -128 -4149 -70 -4114
rect -128 -4183 -116 -4149
rect -82 -4183 -70 -4149
rect -128 -4242 -70 -4183
rect -128 -4276 -116 -4242
rect -82 -4276 -70 -4242
rect -128 -4347 -70 -4276
rect -36 -4129 114 -4059
rect 148 -4061 298 -3991
rect 424 -4001 618 -3967
rect 548 -4025 618 -4001
rect 548 -4035 634 -4025
rect 148 -4095 244 -4061
rect 278 -4095 298 -4061
rect 424 -4040 464 -4035
rect 424 -4074 436 -4040
rect 498 -4069 514 -4035
rect 470 -4074 514 -4069
rect 424 -4078 514 -4074
rect 548 -4069 584 -4035
rect 618 -4069 634 -4035
rect 548 -4083 634 -4069
rect 683 -4034 753 -3924
rect 805 -3890 855 -3871
rect 839 -3924 855 -3890
rect 805 -3966 855 -3924
rect 945 -3890 1011 -3837
rect 945 -3924 961 -3890
rect 995 -3924 1011 -3890
rect 945 -3940 1011 -3924
rect 1045 -3890 1126 -3871
rect 1045 -3924 1059 -3890
rect 1093 -3924 1126 -3890
rect 1045 -3948 1126 -3924
rect 805 -4000 923 -3966
rect 889 -4019 923 -4000
rect 683 -4035 855 -4034
rect 683 -4069 805 -4035
rect 839 -4069 855 -4035
rect 548 -4112 618 -4083
rect -36 -4169 298 -4129
rect -36 -4203 -18 -4169
rect 16 -4203 246 -4169
rect 280 -4203 298 -4169
rect -36 -4271 298 -4203
rect -36 -4305 -18 -4271
rect 16 -4305 246 -4271
rect 280 -4305 298 -4271
rect -36 -4347 298 -4305
rect 332 -4149 390 -4114
rect 332 -4183 344 -4149
rect 378 -4183 390 -4149
rect 332 -4242 390 -4183
rect 332 -4276 344 -4242
rect 378 -4276 390 -4242
rect 332 -4347 390 -4276
rect 424 -4146 618 -4112
rect 683 -4084 855 -4069
rect 889 -4035 1042 -4019
rect 889 -4069 1005 -4035
rect 1039 -4069 1042 -4035
rect 424 -4196 493 -4146
rect 424 -4230 443 -4196
rect 477 -4230 493 -4196
rect 424 -4264 493 -4230
rect 424 -4298 443 -4264
rect 477 -4298 493 -4264
rect 424 -4313 493 -4298
rect 527 -4196 593 -4180
rect 527 -4230 543 -4196
rect 577 -4230 593 -4196
rect 527 -4264 593 -4230
rect 527 -4298 543 -4264
rect 577 -4298 593 -4264
rect 527 -4347 593 -4298
rect 683 -4196 753 -4084
rect 889 -4085 1042 -4069
rect 1076 -4040 1126 -3948
rect 1160 -3931 1218 -3837
rect 1160 -3965 1172 -3931
rect 1206 -3965 1218 -3931
rect 1160 -3982 1218 -3965
rect 1252 -3905 1586 -3837
rect 1252 -3939 1270 -3905
rect 1304 -3939 1534 -3905
rect 1568 -3939 1586 -3905
rect 1252 -3991 1586 -3939
rect 1620 -3931 1678 -3837
rect 1620 -3965 1632 -3931
rect 1666 -3965 1678 -3931
rect 1620 -3982 1678 -3965
rect 1712 -3898 2414 -3837
rect 1712 -3932 1730 -3898
rect 1764 -3932 2362 -3898
rect 2396 -3932 2414 -3898
rect 1712 -3991 2414 -3932
rect 2448 -3931 2506 -3837
rect 2448 -3965 2460 -3931
rect 2494 -3965 2506 -3931
rect 2448 -3982 2506 -3965
rect 2540 -3905 2874 -3837
rect 2540 -3939 2558 -3905
rect 2592 -3939 2822 -3905
rect 2856 -3939 2874 -3905
rect 2540 -3991 2874 -3939
rect 2908 -3931 2966 -3837
rect 2908 -3965 2920 -3931
rect 2954 -3965 2966 -3931
rect 2908 -3982 2966 -3965
rect 3000 -3890 3066 -3871
rect 3000 -3924 3019 -3890
rect 3053 -3924 3066 -3890
rect 3000 -3967 3066 -3924
rect 3100 -3890 3166 -3837
rect 3100 -3924 3116 -3890
rect 3150 -3924 3166 -3890
rect 3100 -3933 3166 -3924
rect 3259 -3890 3329 -3871
rect 3259 -3924 3276 -3890
rect 3310 -3924 3329 -3890
rect 1076 -4074 1081 -4040
rect 1115 -4074 1126 -4040
rect 889 -4119 923 -4085
rect 683 -4230 701 -4196
rect 735 -4230 753 -4196
rect 683 -4264 753 -4230
rect 683 -4298 701 -4264
rect 735 -4298 753 -4264
rect 683 -4313 753 -4298
rect 805 -4153 923 -4119
rect 805 -4195 855 -4153
rect 1076 -4158 1126 -4074
rect 1252 -4059 1272 -4025
rect 1306 -4059 1402 -4025
rect 839 -4229 855 -4195
rect 805 -4263 855 -4229
rect 839 -4297 855 -4263
rect 805 -4313 855 -4297
rect 945 -4196 1011 -4187
rect 945 -4230 961 -4196
rect 995 -4230 1011 -4196
rect 945 -4264 1011 -4230
rect 945 -4298 961 -4264
rect 995 -4298 1011 -4264
rect 945 -4347 1011 -4298
rect 1045 -4195 1126 -4158
rect 1045 -4229 1059 -4195
rect 1093 -4229 1126 -4195
rect 1045 -4263 1126 -4229
rect 1045 -4297 1059 -4263
rect 1093 -4297 1126 -4263
rect 1045 -4313 1126 -4297
rect 1160 -4149 1218 -4114
rect 1160 -4183 1172 -4149
rect 1206 -4183 1218 -4149
rect 1160 -4242 1218 -4183
rect 1160 -4276 1172 -4242
rect 1206 -4276 1218 -4242
rect 1160 -4347 1218 -4276
rect 1252 -4129 1402 -4059
rect 1436 -4061 1586 -3991
rect 1436 -4095 1532 -4061
rect 1566 -4095 1586 -4061
rect 1712 -4059 1790 -4025
rect 1824 -4059 1893 -4025
rect 1927 -4059 1996 -4025
rect 2030 -4059 2050 -4025
rect 1252 -4169 1586 -4129
rect 1252 -4203 1270 -4169
rect 1304 -4203 1534 -4169
rect 1568 -4203 1586 -4169
rect 1252 -4271 1586 -4203
rect 1252 -4305 1270 -4271
rect 1304 -4305 1534 -4271
rect 1568 -4305 1586 -4271
rect 1252 -4347 1586 -4305
rect 1620 -4149 1678 -4114
rect 1620 -4183 1632 -4149
rect 1666 -4183 1678 -4149
rect 1620 -4242 1678 -4183
rect 1620 -4276 1632 -4242
rect 1666 -4276 1678 -4242
rect 1620 -4347 1678 -4276
rect 1712 -4129 2050 -4059
rect 2084 -4061 2414 -3991
rect 2084 -4095 2104 -4061
rect 2138 -4095 2203 -4061
rect 2237 -4095 2302 -4061
rect 2336 -4095 2414 -4061
rect 2540 -4059 2560 -4025
rect 2594 -4059 2690 -4025
rect 1712 -4169 2414 -4129
rect 1712 -4203 1730 -4169
rect 1764 -4203 2362 -4169
rect 2396 -4203 2414 -4169
rect 1712 -4271 2414 -4203
rect 1712 -4305 1730 -4271
rect 1764 -4305 2362 -4271
rect 2396 -4305 2414 -4271
rect 1712 -4347 2414 -4305
rect 2448 -4149 2506 -4114
rect 2448 -4183 2460 -4149
rect 2494 -4183 2506 -4149
rect 2448 -4242 2506 -4183
rect 2448 -4276 2460 -4242
rect 2494 -4276 2506 -4242
rect 2448 -4347 2506 -4276
rect 2540 -4129 2690 -4059
rect 2724 -4061 2874 -3991
rect 3000 -4001 3194 -3967
rect 3124 -4025 3194 -4001
rect 3124 -4035 3210 -4025
rect 2724 -4095 2820 -4061
rect 2854 -4095 2874 -4061
rect 3000 -4069 3040 -4035
rect 3074 -4040 3090 -4035
rect 3000 -4074 3041 -4069
rect 3075 -4074 3090 -4040
rect 3000 -4078 3090 -4074
rect 3124 -4069 3160 -4035
rect 3194 -4069 3210 -4035
rect 3124 -4083 3210 -4069
rect 3259 -4034 3329 -3924
rect 3381 -3890 3431 -3871
rect 3415 -3924 3431 -3890
rect 3381 -3966 3431 -3924
rect 3521 -3890 3587 -3837
rect 3521 -3924 3537 -3890
rect 3571 -3924 3587 -3890
rect 3521 -3940 3587 -3924
rect 3621 -3890 3702 -3871
rect 3621 -3924 3635 -3890
rect 3669 -3924 3702 -3890
rect 3621 -3948 3702 -3924
rect 3381 -4000 3499 -3966
rect 3465 -4019 3499 -4000
rect 3259 -4035 3431 -4034
rect 3259 -4069 3381 -4035
rect 3415 -4069 3431 -4035
rect 3124 -4112 3194 -4083
rect 2540 -4169 2874 -4129
rect 2540 -4203 2558 -4169
rect 2592 -4203 2822 -4169
rect 2856 -4203 2874 -4169
rect 2540 -4271 2874 -4203
rect 2540 -4305 2558 -4271
rect 2592 -4305 2822 -4271
rect 2856 -4305 2874 -4271
rect 2540 -4347 2874 -4305
rect 2908 -4149 2966 -4114
rect 2908 -4183 2920 -4149
rect 2954 -4183 2966 -4149
rect 2908 -4242 2966 -4183
rect 2908 -4276 2920 -4242
rect 2954 -4276 2966 -4242
rect 2908 -4347 2966 -4276
rect 3000 -4146 3194 -4112
rect 3259 -4084 3431 -4069
rect 3465 -4035 3618 -4019
rect 3465 -4069 3581 -4035
rect 3615 -4069 3618 -4035
rect 3000 -4196 3069 -4146
rect 3000 -4230 3019 -4196
rect 3053 -4230 3069 -4196
rect 3000 -4264 3069 -4230
rect 3000 -4298 3019 -4264
rect 3053 -4298 3069 -4264
rect 3000 -4313 3069 -4298
rect 3103 -4196 3169 -4180
rect 3103 -4230 3119 -4196
rect 3153 -4230 3169 -4196
rect 3103 -4264 3169 -4230
rect 3103 -4298 3119 -4264
rect 3153 -4298 3169 -4264
rect 3103 -4347 3169 -4298
rect 3259 -4196 3329 -4084
rect 3465 -4085 3618 -4069
rect 3652 -4040 3702 -3948
rect 3736 -3931 3794 -3837
rect 3736 -3965 3748 -3931
rect 3782 -3965 3794 -3931
rect 3736 -3982 3794 -3965
rect 3828 -3905 4162 -3837
rect 3828 -3939 3846 -3905
rect 3880 -3939 4110 -3905
rect 4144 -3939 4162 -3905
rect 3828 -3991 4162 -3939
rect 4196 -3931 4254 -3837
rect 4196 -3965 4208 -3931
rect 4242 -3965 4254 -3931
rect 4196 -3982 4254 -3965
rect 4288 -3898 4990 -3837
rect 4288 -3932 4306 -3898
rect 4340 -3932 4938 -3898
rect 4972 -3932 4990 -3898
rect 4288 -3991 4990 -3932
rect 5024 -3931 5082 -3837
rect 5024 -3965 5036 -3931
rect 5070 -3965 5082 -3931
rect 5024 -3982 5082 -3965
rect 5116 -3905 5450 -3837
rect 5116 -3939 5134 -3905
rect 5168 -3939 5398 -3905
rect 5432 -3939 5450 -3905
rect 5116 -3991 5450 -3939
rect 5484 -3931 5542 -3837
rect 5484 -3965 5496 -3931
rect 5530 -3965 5542 -3931
rect 5484 -3982 5542 -3965
rect 5576 -3890 5642 -3871
rect 5576 -3924 5595 -3890
rect 5629 -3924 5642 -3890
rect 5576 -3967 5642 -3924
rect 5676 -3890 5742 -3837
rect 5676 -3924 5692 -3890
rect 5726 -3924 5742 -3890
rect 5676 -3933 5742 -3924
rect 5835 -3890 5905 -3871
rect 5835 -3924 5852 -3890
rect 5886 -3924 5905 -3890
rect 3652 -4074 3655 -4040
rect 3689 -4074 3702 -4040
rect 3465 -4119 3499 -4085
rect 3259 -4230 3277 -4196
rect 3311 -4230 3329 -4196
rect 3259 -4264 3329 -4230
rect 3259 -4298 3277 -4264
rect 3311 -4298 3329 -4264
rect 3259 -4313 3329 -4298
rect 3381 -4153 3499 -4119
rect 3381 -4195 3431 -4153
rect 3652 -4158 3702 -4074
rect 3828 -4059 3848 -4025
rect 3882 -4059 3978 -4025
rect 3415 -4229 3431 -4195
rect 3381 -4263 3431 -4229
rect 3415 -4297 3431 -4263
rect 3381 -4313 3431 -4297
rect 3521 -4196 3587 -4187
rect 3521 -4230 3537 -4196
rect 3571 -4230 3587 -4196
rect 3521 -4264 3587 -4230
rect 3521 -4298 3537 -4264
rect 3571 -4298 3587 -4264
rect 3521 -4347 3587 -4298
rect 3621 -4195 3702 -4158
rect 3621 -4229 3635 -4195
rect 3669 -4229 3702 -4195
rect 3621 -4263 3702 -4229
rect 3621 -4297 3635 -4263
rect 3669 -4297 3702 -4263
rect 3621 -4313 3702 -4297
rect 3736 -4149 3794 -4114
rect 3736 -4183 3748 -4149
rect 3782 -4183 3794 -4149
rect 3736 -4242 3794 -4183
rect 3736 -4276 3748 -4242
rect 3782 -4276 3794 -4242
rect 3736 -4347 3794 -4276
rect 3828 -4129 3978 -4059
rect 4012 -4061 4162 -3991
rect 4012 -4095 4108 -4061
rect 4142 -4095 4162 -4061
rect 4288 -4059 4366 -4025
rect 4400 -4059 4469 -4025
rect 4503 -4059 4572 -4025
rect 4606 -4059 4626 -4025
rect 3828 -4169 4162 -4129
rect 3828 -4203 3846 -4169
rect 3880 -4203 4110 -4169
rect 4144 -4203 4162 -4169
rect 3828 -4271 4162 -4203
rect 3828 -4305 3846 -4271
rect 3880 -4305 4110 -4271
rect 4144 -4305 4162 -4271
rect 3828 -4347 4162 -4305
rect 4196 -4149 4254 -4114
rect 4196 -4183 4208 -4149
rect 4242 -4183 4254 -4149
rect 4196 -4242 4254 -4183
rect 4196 -4276 4208 -4242
rect 4242 -4276 4254 -4242
rect 4196 -4347 4254 -4276
rect 4288 -4129 4626 -4059
rect 4660 -4061 4990 -3991
rect 4660 -4095 4680 -4061
rect 4714 -4095 4779 -4061
rect 4813 -4095 4878 -4061
rect 4912 -4095 4990 -4061
rect 5116 -4059 5136 -4025
rect 5170 -4059 5266 -4025
rect 4288 -4169 4990 -4129
rect 4288 -4203 4306 -4169
rect 4340 -4203 4938 -4169
rect 4972 -4203 4990 -4169
rect 4288 -4271 4990 -4203
rect 4288 -4305 4306 -4271
rect 4340 -4305 4938 -4271
rect 4972 -4305 4990 -4271
rect 4288 -4347 4990 -4305
rect 5024 -4149 5082 -4114
rect 5024 -4183 5036 -4149
rect 5070 -4183 5082 -4149
rect 5024 -4242 5082 -4183
rect 5024 -4276 5036 -4242
rect 5070 -4276 5082 -4242
rect 5024 -4347 5082 -4276
rect 5116 -4129 5266 -4059
rect 5300 -4061 5450 -3991
rect 5576 -4001 5770 -3967
rect 5700 -4025 5770 -4001
rect 5700 -4035 5786 -4025
rect 5300 -4095 5396 -4061
rect 5430 -4095 5450 -4061
rect 5576 -4040 5616 -4035
rect 5576 -4074 5615 -4040
rect 5650 -4069 5666 -4035
rect 5649 -4074 5666 -4069
rect 5576 -4078 5666 -4074
rect 5700 -4069 5736 -4035
rect 5770 -4069 5786 -4035
rect 5700 -4083 5786 -4069
rect 5835 -4034 5905 -3924
rect 5957 -3890 6007 -3871
rect 5991 -3924 6007 -3890
rect 5957 -3966 6007 -3924
rect 6097 -3890 6163 -3837
rect 6097 -3924 6113 -3890
rect 6147 -3924 6163 -3890
rect 6097 -3940 6163 -3924
rect 6197 -3890 6278 -3871
rect 6197 -3924 6211 -3890
rect 6245 -3924 6278 -3890
rect 6197 -3948 6278 -3924
rect 5957 -4000 6075 -3966
rect 6041 -4019 6075 -4000
rect 5835 -4035 6007 -4034
rect 5835 -4069 5957 -4035
rect 5991 -4069 6007 -4035
rect 5700 -4112 5770 -4083
rect 5116 -4169 5450 -4129
rect 5116 -4203 5134 -4169
rect 5168 -4203 5398 -4169
rect 5432 -4203 5450 -4169
rect 5116 -4271 5450 -4203
rect 5116 -4305 5134 -4271
rect 5168 -4305 5398 -4271
rect 5432 -4305 5450 -4271
rect 5116 -4347 5450 -4305
rect 5484 -4149 5542 -4114
rect 5484 -4183 5496 -4149
rect 5530 -4183 5542 -4149
rect 5484 -4242 5542 -4183
rect 5484 -4276 5496 -4242
rect 5530 -4276 5542 -4242
rect 5484 -4347 5542 -4276
rect 5576 -4146 5770 -4112
rect 5835 -4084 6007 -4069
rect 6041 -4035 6194 -4019
rect 6041 -4069 6157 -4035
rect 6191 -4069 6194 -4035
rect 5576 -4196 5645 -4146
rect 5576 -4230 5595 -4196
rect 5629 -4230 5645 -4196
rect 5576 -4264 5645 -4230
rect 5576 -4298 5595 -4264
rect 5629 -4298 5645 -4264
rect 5576 -4313 5645 -4298
rect 5679 -4196 5745 -4180
rect 5679 -4230 5695 -4196
rect 5729 -4230 5745 -4196
rect 5679 -4264 5745 -4230
rect 5679 -4298 5695 -4264
rect 5729 -4298 5745 -4264
rect 5679 -4347 5745 -4298
rect 5835 -4196 5905 -4084
rect 6041 -4085 6194 -4069
rect 6228 -4040 6278 -3948
rect 6312 -3931 6370 -3837
rect 6312 -3965 6324 -3931
rect 6358 -3965 6370 -3931
rect 6312 -3982 6370 -3965
rect 6404 -3905 6738 -3837
rect 6404 -3939 6422 -3905
rect 6456 -3939 6686 -3905
rect 6720 -3939 6738 -3905
rect 6404 -3991 6738 -3939
rect 6772 -3931 6830 -3837
rect 6772 -3965 6784 -3931
rect 6818 -3965 6830 -3931
rect 6772 -3982 6830 -3965
rect 6864 -3898 7566 -3837
rect 6864 -3932 6882 -3898
rect 6916 -3932 7514 -3898
rect 7548 -3932 7566 -3898
rect 6864 -3991 7566 -3932
rect 7600 -3931 7658 -3837
rect 7600 -3965 7612 -3931
rect 7646 -3965 7658 -3931
rect 7600 -3982 7658 -3965
rect 7692 -3905 8026 -3837
rect 7692 -3939 7710 -3905
rect 7744 -3939 7974 -3905
rect 8008 -3939 8026 -3905
rect 7692 -3991 8026 -3939
rect 8060 -3931 8118 -3837
rect 8060 -3965 8072 -3931
rect 8106 -3965 8118 -3931
rect 8060 -3982 8118 -3965
rect 8152 -3890 8218 -3871
rect 8152 -3924 8171 -3890
rect 8205 -3924 8218 -3890
rect 8152 -3967 8218 -3924
rect 8252 -3890 8318 -3837
rect 8252 -3924 8268 -3890
rect 8302 -3924 8318 -3890
rect 8252 -3933 8318 -3924
rect 8411 -3890 8481 -3871
rect 8411 -3924 8428 -3890
rect 8462 -3924 8481 -3890
rect 6228 -4074 6229 -4040
rect 6263 -4074 6278 -4040
rect 6041 -4119 6075 -4085
rect 5835 -4230 5853 -4196
rect 5887 -4230 5905 -4196
rect 5835 -4264 5905 -4230
rect 5835 -4298 5853 -4264
rect 5887 -4298 5905 -4264
rect 5835 -4313 5905 -4298
rect 5957 -4153 6075 -4119
rect 5957 -4195 6007 -4153
rect 6228 -4158 6278 -4074
rect 6404 -4059 6424 -4025
rect 6458 -4059 6554 -4025
rect 5991 -4229 6007 -4195
rect 5957 -4263 6007 -4229
rect 5991 -4297 6007 -4263
rect 5957 -4313 6007 -4297
rect 6097 -4196 6163 -4187
rect 6097 -4230 6113 -4196
rect 6147 -4230 6163 -4196
rect 6097 -4264 6163 -4230
rect 6097 -4298 6113 -4264
rect 6147 -4298 6163 -4264
rect 6097 -4347 6163 -4298
rect 6197 -4195 6278 -4158
rect 6197 -4229 6211 -4195
rect 6245 -4229 6278 -4195
rect 6197 -4263 6278 -4229
rect 6197 -4297 6211 -4263
rect 6245 -4297 6278 -4263
rect 6197 -4313 6278 -4297
rect 6312 -4149 6370 -4114
rect 6312 -4183 6324 -4149
rect 6358 -4183 6370 -4149
rect 6312 -4242 6370 -4183
rect 6312 -4276 6324 -4242
rect 6358 -4276 6370 -4242
rect 6312 -4347 6370 -4276
rect 6404 -4129 6554 -4059
rect 6588 -4061 6738 -3991
rect 6588 -4095 6684 -4061
rect 6718 -4095 6738 -4061
rect 6864 -4059 6942 -4025
rect 6976 -4059 7045 -4025
rect 7079 -4059 7148 -4025
rect 7182 -4059 7202 -4025
rect 6404 -4169 6738 -4129
rect 6404 -4203 6422 -4169
rect 6456 -4203 6686 -4169
rect 6720 -4203 6738 -4169
rect 6404 -4271 6738 -4203
rect 6404 -4305 6422 -4271
rect 6456 -4305 6686 -4271
rect 6720 -4305 6738 -4271
rect 6404 -4347 6738 -4305
rect 6772 -4149 6830 -4114
rect 6772 -4183 6784 -4149
rect 6818 -4183 6830 -4149
rect 6772 -4242 6830 -4183
rect 6772 -4276 6784 -4242
rect 6818 -4276 6830 -4242
rect 6772 -4347 6830 -4276
rect 6864 -4129 7202 -4059
rect 7236 -4061 7566 -3991
rect 7236 -4095 7256 -4061
rect 7290 -4095 7355 -4061
rect 7389 -4095 7454 -4061
rect 7488 -4095 7566 -4061
rect 7692 -4059 7712 -4025
rect 7746 -4059 7842 -4025
rect 6864 -4169 7566 -4129
rect 6864 -4203 6882 -4169
rect 6916 -4203 7514 -4169
rect 7548 -4203 7566 -4169
rect 6864 -4271 7566 -4203
rect 6864 -4305 6882 -4271
rect 6916 -4305 7514 -4271
rect 7548 -4305 7566 -4271
rect 6864 -4347 7566 -4305
rect 7600 -4149 7658 -4114
rect 7600 -4183 7612 -4149
rect 7646 -4183 7658 -4149
rect 7600 -4242 7658 -4183
rect 7600 -4276 7612 -4242
rect 7646 -4276 7658 -4242
rect 7600 -4347 7658 -4276
rect 7692 -4129 7842 -4059
rect 7876 -4061 8026 -3991
rect 8152 -4001 8346 -3967
rect 8276 -4025 8346 -4001
rect 8276 -4035 8362 -4025
rect 7876 -4095 7972 -4061
rect 8006 -4095 8026 -4061
rect 8152 -4040 8192 -4035
rect 8152 -4074 8189 -4040
rect 8226 -4069 8242 -4035
rect 8223 -4074 8242 -4069
rect 8152 -4078 8242 -4074
rect 8276 -4069 8312 -4035
rect 8346 -4069 8362 -4035
rect 8276 -4083 8362 -4069
rect 8411 -4034 8481 -3924
rect 8533 -3890 8583 -3871
rect 8567 -3924 8583 -3890
rect 8533 -3966 8583 -3924
rect 8673 -3890 8739 -3837
rect 8673 -3924 8689 -3890
rect 8723 -3924 8739 -3890
rect 8673 -3940 8739 -3924
rect 8773 -3890 8854 -3871
rect 8773 -3924 8787 -3890
rect 8821 -3924 8854 -3890
rect 8773 -3948 8854 -3924
rect 8533 -4000 8651 -3966
rect 8617 -4019 8651 -4000
rect 8411 -4035 8583 -4034
rect 8411 -4069 8533 -4035
rect 8567 -4069 8583 -4035
rect 8276 -4112 8346 -4083
rect 7692 -4169 8026 -4129
rect 7692 -4203 7710 -4169
rect 7744 -4203 7974 -4169
rect 8008 -4203 8026 -4169
rect 7692 -4271 8026 -4203
rect 7692 -4305 7710 -4271
rect 7744 -4305 7974 -4271
rect 8008 -4305 8026 -4271
rect 7692 -4347 8026 -4305
rect 8060 -4149 8118 -4114
rect 8060 -4183 8072 -4149
rect 8106 -4183 8118 -4149
rect 8060 -4242 8118 -4183
rect 8060 -4276 8072 -4242
rect 8106 -4276 8118 -4242
rect 8060 -4347 8118 -4276
rect 8152 -4146 8346 -4112
rect 8411 -4084 8583 -4069
rect 8617 -4035 8770 -4019
rect 8617 -4069 8733 -4035
rect 8767 -4069 8770 -4035
rect 8152 -4196 8221 -4146
rect 8152 -4230 8171 -4196
rect 8205 -4230 8221 -4196
rect 8152 -4264 8221 -4230
rect 8152 -4298 8171 -4264
rect 8205 -4298 8221 -4264
rect 8152 -4313 8221 -4298
rect 8255 -4196 8321 -4180
rect 8255 -4230 8271 -4196
rect 8305 -4230 8321 -4196
rect 8255 -4264 8321 -4230
rect 8255 -4298 8271 -4264
rect 8305 -4298 8321 -4264
rect 8255 -4347 8321 -4298
rect 8411 -4196 8481 -4084
rect 8617 -4085 8770 -4069
rect 8804 -4040 8854 -3948
rect 8888 -3931 8946 -3837
rect 8888 -3965 8900 -3931
rect 8934 -3965 8946 -3931
rect 8888 -3982 8946 -3965
rect 8980 -3905 9314 -3837
rect 8980 -3939 8998 -3905
rect 9032 -3939 9262 -3905
rect 9296 -3939 9314 -3905
rect 8980 -3991 9314 -3939
rect 9348 -3931 9406 -3837
rect 9348 -3965 9360 -3931
rect 9394 -3965 9406 -3931
rect 9348 -3982 9406 -3965
rect 9440 -3898 10142 -3837
rect 9440 -3932 9458 -3898
rect 9492 -3932 10090 -3898
rect 10124 -3932 10142 -3898
rect 9440 -3991 10142 -3932
rect 10176 -3931 10234 -3837
rect 10176 -3965 10188 -3931
rect 10222 -3965 10234 -3931
rect 10176 -3982 10234 -3965
rect 10360 -3905 10694 -3837
rect 10360 -3939 10378 -3905
rect 10412 -3939 10642 -3905
rect 10676 -3939 10694 -3905
rect 10360 -3991 10694 -3939
rect 8804 -4074 8806 -4040
rect 8840 -4074 8854 -4040
rect 8617 -4119 8651 -4085
rect 8411 -4230 8429 -4196
rect 8463 -4230 8481 -4196
rect 8411 -4264 8481 -4230
rect 8411 -4298 8429 -4264
rect 8463 -4298 8481 -4264
rect 8411 -4313 8481 -4298
rect 8533 -4153 8651 -4119
rect 8533 -4195 8583 -4153
rect 8804 -4158 8854 -4074
rect 8980 -4059 9000 -4025
rect 9034 -4059 9130 -4025
rect 8567 -4229 8583 -4195
rect 8533 -4263 8583 -4229
rect 8567 -4297 8583 -4263
rect 8533 -4313 8583 -4297
rect 8673 -4196 8739 -4187
rect 8673 -4230 8689 -4196
rect 8723 -4230 8739 -4196
rect 8673 -4264 8739 -4230
rect 8673 -4298 8689 -4264
rect 8723 -4298 8739 -4264
rect 8673 -4347 8739 -4298
rect 8773 -4195 8854 -4158
rect 8773 -4229 8787 -4195
rect 8821 -4229 8854 -4195
rect 8773 -4263 8854 -4229
rect 8773 -4297 8787 -4263
rect 8821 -4297 8854 -4263
rect 8773 -4313 8854 -4297
rect 8888 -4149 8946 -4114
rect 8888 -4183 8900 -4149
rect 8934 -4183 8946 -4149
rect 8888 -4242 8946 -4183
rect 8888 -4276 8900 -4242
rect 8934 -4276 8946 -4242
rect 8888 -4347 8946 -4276
rect 8980 -4129 9130 -4059
rect 9164 -4061 9314 -3991
rect 9164 -4095 9260 -4061
rect 9294 -4095 9314 -4061
rect 9440 -4059 9518 -4025
rect 9552 -4059 9621 -4025
rect 9655 -4059 9724 -4025
rect 9758 -4059 9778 -4025
rect 8980 -4169 9314 -4129
rect 8980 -4203 8998 -4169
rect 9032 -4203 9262 -4169
rect 9296 -4203 9314 -4169
rect 8980 -4271 9314 -4203
rect 8980 -4305 8998 -4271
rect 9032 -4305 9262 -4271
rect 9296 -4305 9314 -4271
rect 8980 -4347 9314 -4305
rect 9348 -4149 9406 -4114
rect 9348 -4183 9360 -4149
rect 9394 -4183 9406 -4149
rect 9348 -4242 9406 -4183
rect 9348 -4276 9360 -4242
rect 9394 -4276 9406 -4242
rect 9348 -4347 9406 -4276
rect 9440 -4129 9778 -4059
rect 9812 -4061 10142 -3991
rect 9812 -4095 9832 -4061
rect 9866 -4095 9931 -4061
rect 9965 -4095 10030 -4061
rect 10064 -4095 10142 -4061
rect 10360 -4059 10380 -4025
rect 10414 -4059 10510 -4025
rect 9440 -4169 10142 -4129
rect 9440 -4203 9458 -4169
rect 9492 -4203 10090 -4169
rect 10124 -4203 10142 -4169
rect 9440 -4271 10142 -4203
rect 9440 -4305 9458 -4271
rect 9492 -4305 10090 -4271
rect 10124 -4305 10142 -4271
rect 9440 -4347 10142 -4305
rect 10176 -4149 10234 -4114
rect 10176 -4183 10188 -4149
rect 10222 -4183 10234 -4149
rect 10176 -4242 10234 -4183
rect 10176 -4276 10188 -4242
rect 10222 -4276 10234 -4242
rect 10176 -4347 10234 -4276
rect 10360 -4129 10510 -4059
rect 10544 -4061 10694 -3991
rect 10728 -3890 10794 -3871
rect 10728 -3924 10747 -3890
rect 10781 -3924 10794 -3890
rect 10728 -3967 10794 -3924
rect 10828 -3890 10894 -3837
rect 10828 -3924 10844 -3890
rect 10878 -3924 10894 -3890
rect 10828 -3933 10894 -3924
rect 10987 -3890 11057 -3871
rect 10987 -3924 11004 -3890
rect 11038 -3924 11057 -3890
rect 10728 -4001 10922 -3967
rect 10852 -4025 10922 -4001
rect 10852 -4035 10938 -4025
rect 10544 -4095 10640 -4061
rect 10674 -4095 10694 -4061
rect 10728 -4040 10768 -4035
rect 10728 -4074 10763 -4040
rect 10802 -4069 10818 -4035
rect 10797 -4074 10818 -4069
rect 10728 -4078 10818 -4074
rect 10852 -4069 10888 -4035
rect 10922 -4069 10938 -4035
rect 10852 -4083 10938 -4069
rect 10987 -4034 11057 -3924
rect 11109 -3890 11159 -3871
rect 11143 -3924 11159 -3890
rect 11109 -3966 11159 -3924
rect 11249 -3890 11315 -3837
rect 11249 -3924 11265 -3890
rect 11299 -3924 11315 -3890
rect 11249 -3940 11315 -3924
rect 11349 -3890 11430 -3871
rect 11349 -3924 11363 -3890
rect 11397 -3924 11430 -3890
rect 11349 -3948 11430 -3924
rect 11109 -4000 11227 -3966
rect 11193 -4019 11227 -4000
rect 10987 -4035 11159 -4034
rect 10987 -4069 11109 -4035
rect 11143 -4069 11159 -4035
rect 10852 -4112 10922 -4083
rect 10360 -4169 10694 -4129
rect 10360 -4203 10378 -4169
rect 10412 -4203 10642 -4169
rect 10676 -4203 10694 -4169
rect 10360 -4271 10694 -4203
rect 10360 -4305 10378 -4271
rect 10412 -4305 10642 -4271
rect 10676 -4305 10694 -4271
rect 10360 -4347 10694 -4305
rect 10728 -4146 10922 -4112
rect 10987 -4084 11159 -4069
rect 11193 -4035 11346 -4019
rect 11193 -4069 11309 -4035
rect 11343 -4069 11346 -4035
rect 10728 -4196 10797 -4146
rect 10728 -4230 10747 -4196
rect 10781 -4230 10797 -4196
rect 10728 -4264 10797 -4230
rect 10728 -4298 10747 -4264
rect 10781 -4298 10797 -4264
rect 10728 -4313 10797 -4298
rect 10831 -4196 10897 -4180
rect 10831 -4230 10847 -4196
rect 10881 -4230 10897 -4196
rect 10831 -4264 10897 -4230
rect 10831 -4298 10847 -4264
rect 10881 -4298 10897 -4264
rect 10831 -4347 10897 -4298
rect 10987 -4196 11057 -4084
rect 11193 -4085 11346 -4069
rect 11380 -4077 11430 -3948
rect 11464 -3931 11522 -3837
rect 11464 -3965 11476 -3931
rect 11510 -3965 11522 -3931
rect 11464 -3982 11522 -3965
rect 11648 -3905 11982 -3837
rect 11648 -3939 11666 -3905
rect 11700 -3939 11930 -3905
rect 11964 -3939 11982 -3905
rect 11648 -3991 11982 -3939
rect 12384 -3931 12442 -3837
rect 12572 -3881 12631 -3837
rect 12572 -3915 12588 -3881
rect 12622 -3915 12631 -3881
rect 12572 -3931 12631 -3915
rect 12665 -3892 12717 -3876
rect 12665 -3926 12674 -3892
rect 12708 -3926 12717 -3892
rect 12384 -3965 12396 -3931
rect 12430 -3965 12442 -3931
rect 12665 -3965 12717 -3926
rect 12751 -3881 12803 -3837
rect 12751 -3915 12760 -3881
rect 12794 -3915 12803 -3881
rect 12751 -3931 12803 -3915
rect 12837 -3892 12888 -3876
rect 12837 -3926 12846 -3892
rect 12880 -3926 12888 -3892
rect 12837 -3965 12888 -3926
rect 12922 -3881 12982 -3837
rect 12922 -3915 12932 -3881
rect 12966 -3915 12982 -3881
rect 12922 -3931 12982 -3915
rect 13120 -3931 13178 -3837
rect 13120 -3965 13132 -3931
rect 13166 -3965 13178 -3931
rect 12384 -3982 12442 -3965
rect 11193 -4119 11227 -4085
rect 10987 -4230 11005 -4196
rect 11039 -4230 11057 -4196
rect 10987 -4264 11057 -4230
rect 10987 -4298 11005 -4264
rect 11039 -4298 11057 -4264
rect 10987 -4313 11057 -4298
rect 11109 -4153 11227 -4119
rect 11380 -4111 11386 -4077
rect 11420 -4111 11430 -4077
rect 11109 -4195 11159 -4153
rect 11380 -4158 11430 -4111
rect 11648 -4059 11668 -4025
rect 11702 -4059 11798 -4025
rect 11143 -4229 11159 -4195
rect 11109 -4263 11159 -4229
rect 11143 -4297 11159 -4263
rect 11109 -4313 11159 -4297
rect 11249 -4196 11315 -4187
rect 11249 -4230 11265 -4196
rect 11299 -4230 11315 -4196
rect 11249 -4264 11315 -4230
rect 11249 -4298 11265 -4264
rect 11299 -4298 11315 -4264
rect 11249 -4347 11315 -4298
rect 11349 -4195 11430 -4158
rect 11349 -4229 11363 -4195
rect 11397 -4229 11430 -4195
rect 11349 -4263 11430 -4229
rect 11349 -4297 11363 -4263
rect 11397 -4297 11430 -4263
rect 11349 -4313 11430 -4297
rect 11464 -4149 11522 -4114
rect 11464 -4183 11476 -4149
rect 11510 -4183 11522 -4149
rect 11464 -4242 11522 -4183
rect 11464 -4276 11476 -4242
rect 11510 -4276 11522 -4242
rect 11464 -4347 11522 -4276
rect 11648 -4129 11798 -4059
rect 11832 -4061 11982 -3991
rect 11832 -4095 11928 -4061
rect 11962 -4095 11982 -4061
rect 12514 -3975 13086 -3965
rect 12514 -3999 13042 -3975
rect 12480 -4037 12514 -3999
rect 13026 -4009 13042 -3999
rect 13076 -4009 13086 -3975
rect 13120 -3982 13178 -3965
rect 13212 -3905 13546 -3837
rect 13212 -3939 13230 -3905
rect 13264 -3939 13494 -3905
rect 13528 -3939 13546 -3905
rect 12480 -4111 12514 -4071
rect 12548 -4035 12991 -4033
rect 12548 -4039 12574 -4035
rect 12548 -4073 12568 -4039
rect 12608 -4069 12642 -4035
rect 12676 -4039 12710 -4035
rect 12693 -4069 12710 -4039
rect 12744 -4039 12778 -4035
rect 12744 -4069 12765 -4039
rect 12812 -4069 12846 -4035
rect 12880 -4041 12914 -4035
rect 12948 -4041 12991 -4035
rect 12892 -4069 12914 -4041
rect 12602 -4073 12659 -4069
rect 12693 -4073 12765 -4069
rect 12799 -4073 12858 -4069
rect 12548 -4075 12858 -4073
rect 12892 -4075 12942 -4069
rect 12976 -4075 12991 -4041
rect 12548 -4078 12991 -4075
rect 13026 -4052 13086 -4009
rect 11648 -4169 11982 -4129
rect 11648 -4203 11666 -4169
rect 11700 -4203 11930 -4169
rect 11964 -4203 11982 -4169
rect 11648 -4271 11982 -4203
rect 11648 -4305 11666 -4271
rect 11700 -4305 11930 -4271
rect 11964 -4305 11982 -4271
rect 11648 -4347 11982 -4305
rect 12384 -4149 12442 -4114
rect 13026 -4086 13039 -4052
rect 13073 -4086 13086 -4052
rect 13026 -4112 13086 -4086
rect 13212 -3991 13546 -3939
rect 13580 -3931 13638 -3837
rect 13580 -3965 13592 -3931
rect 13626 -3965 13638 -3931
rect 13672 -3879 13733 -3837
rect 13672 -3913 13690 -3879
rect 13724 -3913 13733 -3879
rect 13672 -3939 13733 -3913
rect 13769 -3892 13819 -3873
rect 13769 -3926 13776 -3892
rect 13810 -3926 13819 -3892
rect 13580 -3982 13638 -3965
rect 13212 -4061 13362 -3991
rect 13672 -4008 13735 -3973
rect 13212 -4095 13232 -4061
rect 13266 -4095 13362 -4061
rect 13396 -4059 13492 -4025
rect 13526 -4059 13546 -4025
rect 12514 -4145 13086 -4112
rect 12480 -4146 13086 -4145
rect 12384 -4183 12396 -4149
rect 12430 -4183 12442 -4149
rect 12580 -4169 12631 -4146
rect 12384 -4242 12442 -4183
rect 12384 -4276 12396 -4242
rect 12430 -4276 12442 -4242
rect 12384 -4347 12442 -4276
rect 12476 -4196 12545 -4180
rect 12476 -4230 12502 -4196
rect 12536 -4230 12545 -4196
rect 12476 -4264 12545 -4230
rect 12476 -4298 12502 -4264
rect 12536 -4298 12545 -4264
rect 12476 -4347 12545 -4298
rect 12580 -4203 12588 -4169
rect 12622 -4203 12631 -4169
rect 12752 -4169 12803 -4146
rect 12580 -4257 12631 -4203
rect 12580 -4291 12588 -4257
rect 12622 -4291 12631 -4257
rect 12580 -4307 12631 -4291
rect 12665 -4196 12717 -4180
rect 12665 -4230 12674 -4196
rect 12708 -4230 12717 -4196
rect 12665 -4264 12717 -4230
rect 12665 -4298 12674 -4264
rect 12708 -4298 12717 -4264
rect 12665 -4347 12717 -4298
rect 12752 -4203 12760 -4169
rect 12794 -4203 12803 -4169
rect 12923 -4169 12975 -4146
rect 12752 -4257 12803 -4203
rect 12752 -4291 12760 -4257
rect 12794 -4291 12803 -4257
rect 12752 -4307 12803 -4291
rect 12837 -4196 12889 -4180
rect 12837 -4230 12846 -4196
rect 12880 -4230 12889 -4196
rect 12837 -4264 12889 -4230
rect 12837 -4298 12846 -4264
rect 12880 -4298 12889 -4264
rect 12837 -4347 12889 -4298
rect 12923 -4203 12932 -4169
rect 12966 -4203 12975 -4169
rect 13120 -4149 13178 -4114
rect 13396 -4129 13546 -4059
rect 13672 -4042 13685 -4008
rect 13719 -4035 13735 -4008
rect 13672 -4069 13692 -4042
rect 13726 -4069 13735 -4035
rect 13672 -4085 13735 -4069
rect 13769 -4035 13819 -3926
rect 13853 -3892 13905 -3837
rect 13853 -3926 13862 -3892
rect 13896 -3926 13905 -3892
rect 13853 -3942 13905 -3926
rect 13941 -3892 13991 -3873
rect 13941 -3926 13948 -3892
rect 13982 -3926 13991 -3892
rect 13941 -4035 13991 -3926
rect 14025 -3892 14077 -3837
rect 14025 -3926 14034 -3892
rect 14068 -3926 14077 -3892
rect 14025 -3949 14077 -3926
rect 14111 -3892 14163 -3876
rect 14111 -3926 14120 -3892
rect 14154 -3926 14163 -3892
rect 14111 -3967 14163 -3926
rect 14197 -3883 14249 -3837
rect 14197 -3917 14206 -3883
rect 14240 -3917 14249 -3883
rect 14197 -3933 14249 -3917
rect 14283 -3892 14335 -3876
rect 14283 -3926 14292 -3892
rect 14326 -3926 14335 -3892
rect 14283 -3967 14335 -3926
rect 14369 -3883 14421 -3837
rect 14369 -3917 14378 -3883
rect 14412 -3917 14421 -3883
rect 14369 -3933 14421 -3917
rect 14455 -3892 14507 -3876
rect 14455 -3926 14464 -3892
rect 14498 -3926 14507 -3892
rect 14455 -3967 14507 -3926
rect 14541 -3883 14590 -3837
rect 14541 -3917 14550 -3883
rect 14584 -3917 14590 -3883
rect 14541 -3933 14590 -3917
rect 14624 -3892 14679 -3876
rect 14624 -3926 14636 -3892
rect 14670 -3926 14679 -3892
rect 14624 -3967 14679 -3926
rect 14713 -3883 14762 -3837
rect 14713 -3917 14722 -3883
rect 14756 -3917 14762 -3883
rect 14713 -3933 14762 -3917
rect 14796 -3892 14848 -3876
rect 14796 -3926 14807 -3892
rect 14841 -3926 14848 -3892
rect 14796 -3967 14848 -3926
rect 14884 -3883 14934 -3837
rect 14884 -3917 14893 -3883
rect 14927 -3917 14934 -3883
rect 14884 -3933 14934 -3917
rect 14968 -3892 15020 -3876
rect 14968 -3926 14979 -3892
rect 15013 -3926 15020 -3892
rect 14968 -3967 15020 -3926
rect 15056 -3883 15106 -3837
rect 15056 -3917 15065 -3883
rect 15099 -3917 15106 -3883
rect 15056 -3933 15106 -3917
rect 15140 -3892 15192 -3876
rect 15140 -3926 15151 -3892
rect 15185 -3926 15192 -3892
rect 15140 -3967 15192 -3926
rect 15228 -3883 15280 -3837
rect 15228 -3917 15237 -3883
rect 15271 -3917 15280 -3883
rect 15228 -3933 15280 -3917
rect 15314 -3892 15366 -3876
rect 15314 -3926 15323 -3892
rect 15357 -3926 15366 -3892
rect 15314 -3967 15366 -3926
rect 15400 -3883 15460 -3837
rect 15400 -3917 15409 -3883
rect 15443 -3917 15460 -3883
rect 15400 -3933 15460 -3917
rect 15512 -3931 15570 -3837
rect 15512 -3965 15524 -3931
rect 15558 -3965 15570 -3931
rect 14111 -3996 15460 -3967
rect 15512 -3982 15570 -3965
rect 15604 -3898 16673 -3837
rect 15604 -3932 15622 -3898
rect 15656 -3932 16622 -3898
rect 16656 -3932 16673 -3898
rect 14111 -4001 15248 -3996
rect 15227 -4030 15248 -4001
rect 15282 -4030 15341 -3996
rect 15375 -4030 15460 -3996
rect 13769 -4069 14119 -4035
rect 14153 -4069 14187 -4035
rect 14221 -4069 14255 -4035
rect 14289 -4069 14323 -4035
rect 14357 -4069 14391 -4035
rect 14425 -4069 14459 -4035
rect 14493 -4069 14527 -4035
rect 14561 -4069 14595 -4035
rect 14629 -4069 14663 -4035
rect 14697 -4069 14731 -4035
rect 14765 -4069 14799 -4035
rect 14833 -4069 14867 -4035
rect 14901 -4069 14935 -4035
rect 14969 -4069 15003 -4035
rect 15037 -4069 15071 -4035
rect 15105 -4069 15139 -4035
rect 15173 -4069 15193 -4035
rect 13769 -4085 15193 -4069
rect 12923 -4257 12975 -4203
rect 12923 -4291 12932 -4257
rect 12966 -4291 12975 -4257
rect 12923 -4307 12975 -4291
rect 13009 -4196 13086 -4180
rect 13009 -4230 13018 -4196
rect 13052 -4230 13086 -4196
rect 13009 -4264 13086 -4230
rect 13009 -4298 13018 -4264
rect 13052 -4298 13086 -4264
rect 13009 -4347 13086 -4298
rect 13120 -4183 13132 -4149
rect 13166 -4183 13178 -4149
rect 13120 -4242 13178 -4183
rect 13120 -4276 13132 -4242
rect 13166 -4276 13178 -4242
rect 13120 -4347 13178 -4276
rect 13212 -4169 13546 -4129
rect 13212 -4203 13230 -4169
rect 13264 -4203 13494 -4169
rect 13528 -4203 13546 -4169
rect 13212 -4271 13546 -4203
rect 13212 -4305 13230 -4271
rect 13264 -4305 13494 -4271
rect 13528 -4305 13546 -4271
rect 13212 -4347 13546 -4305
rect 13580 -4149 13638 -4114
rect 13580 -4183 13592 -4149
rect 13626 -4183 13638 -4149
rect 13580 -4242 13638 -4183
rect 13580 -4276 13592 -4242
rect 13626 -4276 13638 -4242
rect 13580 -4347 13638 -4276
rect 13674 -4203 13733 -4185
rect 13674 -4237 13690 -4203
rect 13724 -4237 13733 -4203
rect 13674 -4271 13733 -4237
rect 13674 -4305 13690 -4271
rect 13724 -4305 13733 -4271
rect 13674 -4347 13733 -4305
rect 13769 -4195 13818 -4085
rect 13769 -4229 13776 -4195
rect 13810 -4229 13818 -4195
rect 13769 -4263 13818 -4229
rect 13769 -4297 13776 -4263
rect 13810 -4297 13818 -4263
rect 13769 -4313 13818 -4297
rect 13853 -4203 13905 -4185
rect 13853 -4237 13862 -4203
rect 13896 -4237 13905 -4203
rect 13853 -4271 13905 -4237
rect 13853 -4305 13862 -4271
rect 13896 -4305 13905 -4271
rect 13853 -4347 13905 -4305
rect 13941 -4187 13991 -4085
rect 15227 -4092 15460 -4030
rect 15227 -4119 15248 -4092
rect 14111 -4126 15248 -4119
rect 15282 -4126 15340 -4092
rect 15374 -4126 15460 -4092
rect 15604 -3991 16673 -3932
rect 15604 -4061 16120 -3991
rect 15604 -4095 15682 -4061
rect 15716 -4095 15810 -4061
rect 15844 -4095 15938 -4061
rect 15972 -4095 16066 -4061
rect 16100 -4095 16120 -4061
rect 16154 -4059 16174 -4025
rect 16208 -4059 16302 -4025
rect 16336 -4059 16430 -4025
rect 16464 -4059 16558 -4025
rect 16592 -4059 16673 -4025
rect 14111 -4141 15460 -4126
rect 14111 -4175 14120 -4141
rect 14154 -4167 14292 -4141
rect 14154 -4175 14163 -4167
rect 13941 -4221 13948 -4187
rect 13982 -4221 13991 -4187
rect 13941 -4255 13991 -4221
rect 13941 -4289 13948 -4255
rect 13982 -4289 13991 -4255
rect 13941 -4312 13991 -4289
rect 14025 -4203 14077 -4187
rect 14025 -4237 14034 -4203
rect 14068 -4237 14077 -4203
rect 14025 -4271 14077 -4237
rect 14025 -4305 14034 -4271
rect 14068 -4305 14077 -4271
rect 14025 -4346 14077 -4305
rect 14111 -4227 14163 -4175
rect 14283 -4175 14292 -4167
rect 14326 -4167 14464 -4141
rect 14326 -4175 14335 -4167
rect 14111 -4261 14120 -4227
rect 14154 -4261 14163 -4227
rect 14111 -4312 14163 -4261
rect 14197 -4247 14249 -4201
rect 14197 -4281 14206 -4247
rect 14240 -4281 14249 -4247
rect 14197 -4346 14249 -4281
rect 14283 -4227 14335 -4175
rect 14455 -4175 14464 -4167
rect 14498 -4167 14636 -4141
rect 14498 -4175 14507 -4167
rect 14283 -4261 14292 -4227
rect 14326 -4261 14335 -4227
rect 14283 -4312 14335 -4261
rect 14369 -4247 14421 -4201
rect 14369 -4281 14378 -4247
rect 14412 -4281 14421 -4247
rect 14369 -4346 14421 -4281
rect 14455 -4227 14507 -4175
rect 14627 -4175 14636 -4167
rect 14670 -4167 14807 -4141
rect 14670 -4175 14679 -4167
rect 14455 -4261 14464 -4227
rect 14498 -4261 14507 -4227
rect 14455 -4312 14507 -4261
rect 14541 -4247 14593 -4201
rect 14541 -4281 14550 -4247
rect 14584 -4281 14593 -4247
rect 14541 -4346 14593 -4281
rect 14627 -4227 14679 -4175
rect 14796 -4175 14807 -4167
rect 14841 -4167 14979 -4141
rect 14841 -4175 14848 -4167
rect 14627 -4261 14636 -4227
rect 14670 -4261 14679 -4227
rect 14627 -4312 14679 -4261
rect 14713 -4247 14762 -4201
rect 14713 -4281 14722 -4247
rect 14756 -4281 14762 -4247
rect 14713 -4346 14762 -4281
rect 14796 -4227 14848 -4175
rect 14968 -4175 14979 -4167
rect 15013 -4167 15151 -4141
rect 15013 -4175 15020 -4167
rect 14796 -4261 14807 -4227
rect 14841 -4261 14848 -4227
rect 14796 -4312 14848 -4261
rect 14885 -4247 14934 -4201
rect 14885 -4281 14893 -4247
rect 14927 -4281 14934 -4247
rect 14885 -4346 14934 -4281
rect 14968 -4227 15020 -4175
rect 15140 -4175 15151 -4167
rect 15185 -4164 15323 -4141
rect 15185 -4175 15192 -4164
rect 14968 -4261 14979 -4227
rect 15013 -4261 15020 -4227
rect 14968 -4312 15020 -4261
rect 15057 -4247 15106 -4201
rect 15057 -4281 15065 -4247
rect 15099 -4281 15106 -4247
rect 15057 -4346 15106 -4281
rect 15140 -4227 15192 -4175
rect 15314 -4175 15323 -4164
rect 15357 -4164 15460 -4141
rect 15512 -4149 15570 -4114
rect 16154 -4129 16673 -4059
rect 15357 -4175 15372 -4164
rect 15140 -4261 15151 -4227
rect 15185 -4261 15192 -4227
rect 15140 -4312 15192 -4261
rect 15229 -4247 15280 -4201
rect 15229 -4281 15237 -4247
rect 15271 -4281 15280 -4247
rect 15229 -4346 15280 -4281
rect 15314 -4227 15372 -4175
rect 15512 -4183 15524 -4149
rect 15558 -4183 15570 -4149
rect 15314 -4261 15323 -4227
rect 15357 -4261 15372 -4227
rect 15314 -4312 15372 -4261
rect 15406 -4247 15460 -4198
rect 15406 -4281 15409 -4247
rect 15443 -4281 15460 -4247
rect 14025 -4347 15280 -4346
rect 15406 -4347 15460 -4281
rect 15512 -4242 15570 -4183
rect 15512 -4276 15524 -4242
rect 15558 -4276 15570 -4242
rect 15512 -4347 15570 -4276
rect 15604 -4169 16673 -4129
rect 15604 -4203 15622 -4169
rect 15656 -4203 16622 -4169
rect 16656 -4203 16673 -4169
rect 15604 -4271 16673 -4203
rect 15604 -4305 15622 -4271
rect 15656 -4305 16622 -4271
rect 16656 -4305 16673 -4271
rect 15604 -4347 16673 -4305
rect -2997 -4381 -2968 -4347
rect -2934 -4381 -2876 -4347
rect -2842 -4381 -2784 -4347
rect -2750 -4381 -2692 -4347
rect -2658 -4381 -2600 -4347
rect -2566 -4381 -2508 -4347
rect -2474 -4381 -2416 -4347
rect -2382 -4381 -2324 -4347
rect -2290 -4381 -2232 -4347
rect -2198 -4381 -2140 -4347
rect -2106 -4381 -2048 -4347
rect -2014 -4381 -1956 -4347
rect -1922 -4381 -1864 -4347
rect -1830 -4381 -1772 -4347
rect -1738 -4381 -1680 -4347
rect -1646 -4381 -1588 -4347
rect -1554 -4381 -1496 -4347
rect -1462 -4381 -1404 -4347
rect -1370 -4381 -1312 -4347
rect -1278 -4381 -1220 -4347
rect -1186 -4381 -1128 -4347
rect -1094 -4381 -1036 -4347
rect -1002 -4381 -944 -4347
rect -910 -4381 -852 -4347
rect -818 -4381 -760 -4347
rect -726 -4381 -668 -4347
rect -634 -4381 -576 -4347
rect -542 -4381 -484 -4347
rect -450 -4381 -392 -4347
rect -358 -4381 -300 -4347
rect -266 -4381 -208 -4347
rect -174 -4381 -116 -4347
rect -82 -4381 -24 -4347
rect 10 -4381 68 -4347
rect 102 -4381 160 -4347
rect 194 -4381 252 -4347
rect 286 -4381 344 -4347
rect 378 -4381 436 -4347
rect 470 -4381 528 -4347
rect 562 -4381 620 -4347
rect 654 -4381 712 -4347
rect 746 -4381 804 -4347
rect 838 -4381 896 -4347
rect 930 -4381 988 -4347
rect 1022 -4381 1080 -4347
rect 1114 -4381 1172 -4347
rect 1206 -4381 1264 -4347
rect 1298 -4381 1356 -4347
rect 1390 -4381 1448 -4347
rect 1482 -4381 1540 -4347
rect 1574 -4381 1632 -4347
rect 1666 -4381 1724 -4347
rect 1758 -4381 1816 -4347
rect 1850 -4381 1908 -4347
rect 1942 -4381 2000 -4347
rect 2034 -4381 2092 -4347
rect 2126 -4381 2184 -4347
rect 2218 -4381 2276 -4347
rect 2310 -4381 2368 -4347
rect 2402 -4381 2460 -4347
rect 2494 -4381 2552 -4347
rect 2586 -4381 2644 -4347
rect 2678 -4381 2736 -4347
rect 2770 -4381 2828 -4347
rect 2862 -4381 2920 -4347
rect 2954 -4381 3012 -4347
rect 3046 -4381 3104 -4347
rect 3138 -4381 3196 -4347
rect 3230 -4381 3288 -4347
rect 3322 -4381 3380 -4347
rect 3414 -4381 3472 -4347
rect 3506 -4381 3564 -4347
rect 3598 -4381 3656 -4347
rect 3690 -4381 3748 -4347
rect 3782 -4381 3840 -4347
rect 3874 -4381 3932 -4347
rect 3966 -4381 4024 -4347
rect 4058 -4381 4116 -4347
rect 4150 -4381 4208 -4347
rect 4242 -4381 4300 -4347
rect 4334 -4381 4392 -4347
rect 4426 -4381 4484 -4347
rect 4518 -4381 4576 -4347
rect 4610 -4381 4668 -4347
rect 4702 -4381 4760 -4347
rect 4794 -4381 4852 -4347
rect 4886 -4381 4944 -4347
rect 4978 -4381 5036 -4347
rect 5070 -4381 5128 -4347
rect 5162 -4381 5220 -4347
rect 5254 -4381 5312 -4347
rect 5346 -4381 5404 -4347
rect 5438 -4381 5496 -4347
rect 5530 -4381 5588 -4347
rect 5622 -4381 5680 -4347
rect 5714 -4381 5772 -4347
rect 5806 -4381 5864 -4347
rect 5898 -4381 5956 -4347
rect 5990 -4381 6048 -4347
rect 6082 -4381 6140 -4347
rect 6174 -4381 6232 -4347
rect 6266 -4381 6324 -4347
rect 6358 -4381 6416 -4347
rect 6450 -4381 6508 -4347
rect 6542 -4381 6600 -4347
rect 6634 -4381 6692 -4347
rect 6726 -4381 6784 -4347
rect 6818 -4381 6876 -4347
rect 6910 -4381 6968 -4347
rect 7002 -4381 7060 -4347
rect 7094 -4381 7152 -4347
rect 7186 -4381 7244 -4347
rect 7278 -4381 7336 -4347
rect 7370 -4381 7428 -4347
rect 7462 -4381 7520 -4347
rect 7554 -4381 7612 -4347
rect 7646 -4381 7704 -4347
rect 7738 -4381 7796 -4347
rect 7830 -4381 7888 -4347
rect 7922 -4381 7980 -4347
rect 8014 -4381 8072 -4347
rect 8106 -4381 8164 -4347
rect 8198 -4381 8256 -4347
rect 8290 -4381 8348 -4347
rect 8382 -4381 8440 -4347
rect 8474 -4381 8532 -4347
rect 8566 -4381 8624 -4347
rect 8658 -4381 8716 -4347
rect 8750 -4381 8808 -4347
rect 8842 -4381 8900 -4347
rect 8934 -4381 8992 -4347
rect 9026 -4381 9084 -4347
rect 9118 -4381 9176 -4347
rect 9210 -4381 9268 -4347
rect 9302 -4381 9360 -4347
rect 9394 -4381 9452 -4347
rect 9486 -4381 9544 -4347
rect 9578 -4381 9636 -4347
rect 9670 -4381 9728 -4347
rect 9762 -4381 9820 -4347
rect 9854 -4381 9912 -4347
rect 9946 -4381 10004 -4347
rect 10038 -4381 10096 -4347
rect 10130 -4381 10188 -4347
rect 10222 -4381 10280 -4347
rect 10314 -4381 10372 -4347
rect 10406 -4381 10464 -4347
rect 10498 -4381 10556 -4347
rect 10590 -4381 10648 -4347
rect 10682 -4381 10740 -4347
rect 10774 -4381 10832 -4347
rect 10866 -4381 10924 -4347
rect 10958 -4381 11016 -4347
rect 11050 -4381 11108 -4347
rect 11142 -4381 11200 -4347
rect 11234 -4381 11292 -4347
rect 11326 -4381 11384 -4347
rect 11418 -4381 11476 -4347
rect 11510 -4381 11568 -4347
rect 11602 -4381 11660 -4347
rect 11694 -4381 11752 -4347
rect 11786 -4381 11844 -4347
rect 11878 -4381 11936 -4347
rect 11970 -4381 12028 -4347
rect 12062 -4381 12120 -4347
rect 12154 -4381 12212 -4347
rect 12246 -4381 12304 -4347
rect 12338 -4381 12396 -4347
rect 12430 -4381 12488 -4347
rect 12522 -4381 12580 -4347
rect 12614 -4381 12672 -4347
rect 12706 -4381 12764 -4347
rect 12798 -4381 12856 -4347
rect 12890 -4381 12948 -4347
rect 12982 -4381 13040 -4347
rect 13074 -4381 13132 -4347
rect 13166 -4381 13224 -4347
rect 13258 -4381 13316 -4347
rect 13350 -4381 13408 -4347
rect 13442 -4381 13500 -4347
rect 13534 -4381 13592 -4347
rect 13626 -4381 13684 -4347
rect 13718 -4381 13776 -4347
rect 13810 -4381 13868 -4347
rect 13902 -4381 13960 -4347
rect 13994 -4381 14052 -4347
rect 14086 -4381 14144 -4347
rect 14178 -4381 14236 -4347
rect 14270 -4381 14328 -4347
rect 14362 -4381 14420 -4347
rect 14454 -4381 14512 -4347
rect 14546 -4381 14604 -4347
rect 14638 -4381 14696 -4347
rect 14730 -4381 14788 -4347
rect 14822 -4381 14880 -4347
rect 14914 -4381 14972 -4347
rect 15006 -4381 15064 -4347
rect 15098 -4381 15156 -4347
rect 15190 -4381 15248 -4347
rect 15282 -4381 15340 -4347
rect 15374 -4381 15432 -4347
rect 15466 -4381 15524 -4347
rect 15558 -4381 15616 -4347
rect 15650 -4381 15708 -4347
rect 15742 -4381 15800 -4347
rect 15834 -4381 15892 -4347
rect 15926 -4381 15984 -4347
rect 16018 -4381 16076 -4347
rect 16110 -4381 16168 -4347
rect 16202 -4381 16260 -4347
rect 16294 -4381 16352 -4347
rect 16386 -4381 16444 -4347
rect 16478 -4381 16536 -4347
rect 16570 -4381 16628 -4347
rect 16662 -4381 16691 -4347
rect -2980 -4423 -2278 -4381
rect -2980 -4457 -2962 -4423
rect -2928 -4457 -2330 -4423
rect -2296 -4457 -2278 -4423
rect -2980 -4525 -2278 -4457
rect -2980 -4559 -2962 -4525
rect -2928 -4559 -2330 -4525
rect -2296 -4559 -2278 -4525
rect -2980 -4599 -2278 -4559
rect -2980 -4667 -2902 -4633
rect -2868 -4667 -2803 -4633
rect -2769 -4667 -2704 -4633
rect -2670 -4667 -2650 -4633
rect -2980 -4737 -2650 -4667
rect -2616 -4669 -2278 -4599
rect -2244 -4452 -2186 -4381
rect -2244 -4486 -2232 -4452
rect -2198 -4486 -2186 -4452
rect -2244 -4545 -2186 -4486
rect -2244 -4579 -2232 -4545
rect -2198 -4579 -2186 -4545
rect -2244 -4614 -2186 -4579
rect -1600 -4423 -898 -4381
rect -1600 -4457 -1582 -4423
rect -1548 -4457 -950 -4423
rect -916 -4457 -898 -4423
rect -1600 -4525 -898 -4457
rect -1600 -4559 -1582 -4525
rect -1548 -4559 -950 -4525
rect -916 -4559 -898 -4525
rect -1600 -4599 -898 -4559
rect -864 -4431 -783 -4415
rect -864 -4465 -831 -4431
rect -797 -4465 -783 -4431
rect -864 -4499 -783 -4465
rect -864 -4533 -831 -4499
rect -797 -4533 -783 -4499
rect -864 -4570 -783 -4533
rect -749 -4430 -683 -4381
rect -749 -4464 -733 -4430
rect -699 -4464 -683 -4430
rect -749 -4498 -683 -4464
rect -749 -4532 -733 -4498
rect -699 -4532 -683 -4498
rect -749 -4541 -683 -4532
rect -593 -4431 -543 -4415
rect -593 -4465 -577 -4431
rect -593 -4499 -543 -4465
rect -593 -4533 -577 -4499
rect -2616 -4703 -2596 -4669
rect -2562 -4703 -2493 -4669
rect -2459 -4703 -2390 -4669
rect -2356 -4703 -2278 -4669
rect -1600 -4669 -1262 -4599
rect -864 -4619 -814 -4570
rect -593 -4575 -543 -4533
rect -1600 -4703 -1522 -4669
rect -1488 -4703 -1419 -4669
rect -1385 -4703 -1316 -4669
rect -1282 -4703 -1262 -4669
rect -1228 -4667 -1208 -4633
rect -1174 -4667 -1109 -4633
rect -1075 -4667 -1010 -4633
rect -976 -4667 -898 -4633
rect -1228 -4737 -898 -4667
rect -2980 -4796 -2278 -4737
rect -2980 -4830 -2962 -4796
rect -2928 -4830 -2330 -4796
rect -2296 -4830 -2278 -4796
rect -2980 -4891 -2278 -4830
rect -2244 -4763 -2186 -4746
rect -2244 -4797 -2232 -4763
rect -2198 -4797 -2186 -4763
rect -2244 -4891 -2186 -4797
rect -1600 -4796 -898 -4737
rect -1600 -4830 -1582 -4796
rect -1548 -4830 -950 -4796
rect -916 -4830 -898 -4796
rect -1600 -4891 -898 -4830
rect -864 -4653 -855 -4619
rect -821 -4653 -814 -4619
rect -661 -4609 -543 -4575
rect -491 -4430 -421 -4415
rect -491 -4464 -473 -4430
rect -439 -4464 -421 -4430
rect -491 -4498 -421 -4464
rect -491 -4532 -473 -4498
rect -439 -4532 -421 -4498
rect -661 -4643 -627 -4609
rect -864 -4780 -814 -4653
rect -780 -4659 -627 -4643
rect -491 -4644 -421 -4532
rect -331 -4430 -265 -4381
rect -331 -4464 -315 -4430
rect -281 -4464 -265 -4430
rect -331 -4498 -265 -4464
rect -331 -4532 -315 -4498
rect -281 -4532 -265 -4498
rect -331 -4548 -265 -4532
rect -231 -4430 -162 -4415
rect -231 -4464 -215 -4430
rect -181 -4464 -162 -4430
rect -231 -4498 -162 -4464
rect -231 -4532 -215 -4498
rect -181 -4532 -162 -4498
rect -231 -4582 -162 -4532
rect -780 -4693 -777 -4659
rect -743 -4693 -627 -4659
rect -780 -4709 -627 -4693
rect -593 -4659 -421 -4644
rect -356 -4616 -162 -4582
rect -128 -4452 -70 -4381
rect -128 -4486 -116 -4452
rect -82 -4486 -70 -4452
rect -128 -4545 -70 -4486
rect -128 -4579 -116 -4545
rect -82 -4579 -70 -4545
rect -128 -4614 -70 -4579
rect -36 -4423 298 -4381
rect -36 -4457 -18 -4423
rect 16 -4457 246 -4423
rect 280 -4457 298 -4423
rect -36 -4525 298 -4457
rect -36 -4559 -18 -4525
rect 16 -4559 246 -4525
rect 280 -4559 298 -4525
rect -36 -4599 298 -4559
rect 332 -4452 390 -4381
rect 332 -4486 344 -4452
rect 378 -4486 390 -4452
rect 332 -4545 390 -4486
rect 332 -4579 344 -4545
rect 378 -4579 390 -4545
rect -356 -4645 -286 -4616
rect -593 -4693 -577 -4659
rect -543 -4693 -421 -4659
rect -593 -4694 -421 -4693
rect -661 -4728 -627 -4709
rect -661 -4762 -543 -4728
rect -864 -4804 -783 -4780
rect -864 -4838 -831 -4804
rect -797 -4838 -783 -4804
rect -864 -4857 -783 -4838
rect -749 -4804 -683 -4788
rect -749 -4838 -733 -4804
rect -699 -4838 -683 -4804
rect -749 -4891 -683 -4838
rect -593 -4804 -543 -4762
rect -593 -4838 -577 -4804
rect -593 -4857 -543 -4838
rect -491 -4804 -421 -4694
rect -372 -4659 -286 -4645
rect -372 -4693 -356 -4659
rect -322 -4693 -286 -4659
rect -252 -4656 -162 -4650
rect -252 -4659 -210 -4656
rect -252 -4693 -236 -4659
rect -176 -4690 -162 -4656
rect -202 -4693 -162 -4690
rect -36 -4669 114 -4599
rect 332 -4614 390 -4579
rect 424 -4431 505 -4415
rect 424 -4465 457 -4431
rect 491 -4465 505 -4431
rect 424 -4499 505 -4465
rect 424 -4533 457 -4499
rect 491 -4533 505 -4499
rect 424 -4570 505 -4533
rect 539 -4430 605 -4381
rect 539 -4464 555 -4430
rect 589 -4464 605 -4430
rect 539 -4498 605 -4464
rect 539 -4532 555 -4498
rect 589 -4532 605 -4498
rect 539 -4541 605 -4532
rect 695 -4431 745 -4415
rect 695 -4465 711 -4431
rect 695 -4499 745 -4465
rect 695 -4533 711 -4499
rect 424 -4619 474 -4570
rect 695 -4575 745 -4533
rect -372 -4703 -286 -4693
rect -36 -4703 -16 -4669
rect 18 -4703 114 -4669
rect 148 -4667 244 -4633
rect 278 -4667 298 -4633
rect -356 -4727 -286 -4703
rect -356 -4761 -162 -4727
rect 148 -4737 298 -4667
rect -491 -4838 -472 -4804
rect -438 -4838 -421 -4804
rect -491 -4857 -421 -4838
rect -328 -4804 -262 -4795
rect -328 -4838 -312 -4804
rect -278 -4838 -262 -4804
rect -328 -4891 -262 -4838
rect -228 -4804 -162 -4761
rect -228 -4838 -215 -4804
rect -181 -4838 -162 -4804
rect -228 -4857 -162 -4838
rect -128 -4763 -70 -4746
rect -128 -4797 -116 -4763
rect -82 -4797 -70 -4763
rect -128 -4891 -70 -4797
rect -36 -4789 298 -4737
rect 424 -4653 433 -4619
rect 467 -4653 474 -4619
rect 627 -4609 745 -4575
rect 797 -4430 867 -4415
rect 797 -4464 815 -4430
rect 849 -4464 867 -4430
rect 797 -4498 867 -4464
rect 797 -4532 815 -4498
rect 849 -4532 867 -4498
rect 627 -4643 661 -4609
rect -36 -4823 -18 -4789
rect 16 -4823 246 -4789
rect 280 -4823 298 -4789
rect -36 -4891 298 -4823
rect 332 -4763 390 -4746
rect 332 -4797 344 -4763
rect 378 -4797 390 -4763
rect 332 -4891 390 -4797
rect 424 -4780 474 -4653
rect 508 -4659 661 -4643
rect 797 -4644 867 -4532
rect 957 -4430 1023 -4381
rect 957 -4464 973 -4430
rect 1007 -4464 1023 -4430
rect 957 -4498 1023 -4464
rect 957 -4532 973 -4498
rect 1007 -4532 1023 -4498
rect 957 -4548 1023 -4532
rect 1057 -4430 1126 -4415
rect 1057 -4464 1073 -4430
rect 1107 -4464 1126 -4430
rect 1057 -4498 1126 -4464
rect 1057 -4532 1073 -4498
rect 1107 -4532 1126 -4498
rect 1057 -4582 1126 -4532
rect 508 -4693 511 -4659
rect 545 -4693 661 -4659
rect 508 -4709 661 -4693
rect 695 -4659 867 -4644
rect 932 -4616 1126 -4582
rect 1160 -4452 1218 -4381
rect 1160 -4486 1172 -4452
rect 1206 -4486 1218 -4452
rect 1160 -4545 1218 -4486
rect 1160 -4579 1172 -4545
rect 1206 -4579 1218 -4545
rect 1160 -4614 1218 -4579
rect 1252 -4423 1586 -4381
rect 1252 -4457 1270 -4423
rect 1304 -4457 1534 -4423
rect 1568 -4457 1586 -4423
rect 1252 -4525 1586 -4457
rect 1252 -4559 1270 -4525
rect 1304 -4559 1534 -4525
rect 1568 -4559 1586 -4525
rect 1252 -4599 1586 -4559
rect 1620 -4452 1678 -4381
rect 1620 -4486 1632 -4452
rect 1666 -4486 1678 -4452
rect 1620 -4545 1678 -4486
rect 1620 -4579 1632 -4545
rect 1666 -4579 1678 -4545
rect 932 -4645 1002 -4616
rect 695 -4693 711 -4659
rect 745 -4693 867 -4659
rect 695 -4694 867 -4693
rect 627 -4728 661 -4709
rect 627 -4762 745 -4728
rect 424 -4804 505 -4780
rect 424 -4838 457 -4804
rect 491 -4838 505 -4804
rect 424 -4857 505 -4838
rect 539 -4804 605 -4788
rect 539 -4838 555 -4804
rect 589 -4838 605 -4804
rect 539 -4891 605 -4838
rect 695 -4804 745 -4762
rect 695 -4838 711 -4804
rect 695 -4857 745 -4838
rect 797 -4804 867 -4694
rect 916 -4659 1002 -4645
rect 916 -4693 932 -4659
rect 966 -4693 1002 -4659
rect 1036 -4652 1126 -4650
rect 1036 -4659 1054 -4652
rect 1036 -4693 1052 -4659
rect 1088 -4686 1126 -4652
rect 1086 -4693 1126 -4686
rect 1252 -4669 1402 -4599
rect 1620 -4614 1678 -4579
rect 1712 -4423 2414 -4381
rect 1712 -4457 1730 -4423
rect 1764 -4457 2362 -4423
rect 2396 -4457 2414 -4423
rect 1712 -4525 2414 -4457
rect 1712 -4559 1730 -4525
rect 1764 -4559 2362 -4525
rect 2396 -4559 2414 -4525
rect 1712 -4599 2414 -4559
rect 916 -4703 1002 -4693
rect 1252 -4703 1272 -4669
rect 1306 -4703 1402 -4669
rect 1436 -4667 1532 -4633
rect 1566 -4667 1586 -4633
rect 932 -4727 1002 -4703
rect 932 -4761 1126 -4727
rect 1436 -4737 1586 -4667
rect 797 -4838 816 -4804
rect 850 -4838 867 -4804
rect 797 -4857 867 -4838
rect 960 -4804 1026 -4795
rect 960 -4838 976 -4804
rect 1010 -4838 1026 -4804
rect 960 -4891 1026 -4838
rect 1060 -4804 1126 -4761
rect 1060 -4838 1073 -4804
rect 1107 -4838 1126 -4804
rect 1060 -4857 1126 -4838
rect 1160 -4763 1218 -4746
rect 1160 -4797 1172 -4763
rect 1206 -4797 1218 -4763
rect 1160 -4891 1218 -4797
rect 1252 -4789 1586 -4737
rect 1712 -4667 1790 -4633
rect 1824 -4667 1889 -4633
rect 1923 -4667 1988 -4633
rect 2022 -4667 2042 -4633
rect 1712 -4737 2042 -4667
rect 2076 -4669 2414 -4599
rect 2448 -4452 2506 -4381
rect 2448 -4486 2460 -4452
rect 2494 -4486 2506 -4452
rect 2448 -4545 2506 -4486
rect 2448 -4579 2460 -4545
rect 2494 -4579 2506 -4545
rect 2448 -4614 2506 -4579
rect 2540 -4423 2874 -4381
rect 2540 -4457 2558 -4423
rect 2592 -4457 2822 -4423
rect 2856 -4457 2874 -4423
rect 2540 -4525 2874 -4457
rect 2540 -4559 2558 -4525
rect 2592 -4559 2822 -4525
rect 2856 -4559 2874 -4525
rect 2540 -4599 2874 -4559
rect 2908 -4452 2966 -4381
rect 2908 -4486 2920 -4452
rect 2954 -4486 2966 -4452
rect 2908 -4545 2966 -4486
rect 2908 -4579 2920 -4545
rect 2954 -4579 2966 -4545
rect 2076 -4703 2096 -4669
rect 2130 -4703 2199 -4669
rect 2233 -4703 2302 -4669
rect 2336 -4703 2414 -4669
rect 2540 -4669 2690 -4599
rect 2908 -4614 2966 -4579
rect 3000 -4431 3081 -4415
rect 3000 -4465 3033 -4431
rect 3067 -4465 3081 -4431
rect 3000 -4499 3081 -4465
rect 3000 -4533 3033 -4499
rect 3067 -4533 3081 -4499
rect 3000 -4570 3081 -4533
rect 3115 -4430 3181 -4381
rect 3115 -4464 3131 -4430
rect 3165 -4464 3181 -4430
rect 3115 -4498 3181 -4464
rect 3115 -4532 3131 -4498
rect 3165 -4532 3181 -4498
rect 3115 -4541 3181 -4532
rect 3271 -4431 3321 -4415
rect 3271 -4465 3287 -4431
rect 3271 -4499 3321 -4465
rect 3271 -4533 3287 -4499
rect 2540 -4703 2560 -4669
rect 2594 -4703 2690 -4669
rect 2724 -4667 2820 -4633
rect 2854 -4667 2874 -4633
rect 2724 -4737 2874 -4667
rect 1252 -4823 1270 -4789
rect 1304 -4823 1534 -4789
rect 1568 -4823 1586 -4789
rect 1252 -4891 1586 -4823
rect 1620 -4763 1678 -4746
rect 1620 -4797 1632 -4763
rect 1666 -4797 1678 -4763
rect 1620 -4891 1678 -4797
rect 1712 -4796 2414 -4737
rect 1712 -4830 1730 -4796
rect 1764 -4830 2362 -4796
rect 2396 -4830 2414 -4796
rect 1712 -4891 2414 -4830
rect 2448 -4763 2506 -4746
rect 2448 -4797 2460 -4763
rect 2494 -4797 2506 -4763
rect 2448 -4891 2506 -4797
rect 2540 -4789 2874 -4737
rect 3000 -4652 3050 -4570
rect 3271 -4575 3321 -4533
rect 3203 -4609 3321 -4575
rect 3373 -4430 3443 -4415
rect 3373 -4464 3391 -4430
rect 3425 -4464 3443 -4430
rect 3373 -4498 3443 -4464
rect 3373 -4532 3391 -4498
rect 3425 -4532 3443 -4498
rect 3203 -4643 3237 -4609
rect 3000 -4686 3014 -4652
rect 3048 -4686 3050 -4652
rect 2540 -4823 2558 -4789
rect 2592 -4823 2822 -4789
rect 2856 -4823 2874 -4789
rect 2540 -4891 2874 -4823
rect 2908 -4763 2966 -4746
rect 2908 -4797 2920 -4763
rect 2954 -4797 2966 -4763
rect 2908 -4891 2966 -4797
rect 3000 -4780 3050 -4686
rect 3084 -4659 3237 -4643
rect 3373 -4644 3443 -4532
rect 3533 -4430 3599 -4381
rect 3533 -4464 3549 -4430
rect 3583 -4464 3599 -4430
rect 3533 -4498 3599 -4464
rect 3533 -4532 3549 -4498
rect 3583 -4532 3599 -4498
rect 3533 -4548 3599 -4532
rect 3633 -4430 3702 -4415
rect 3633 -4464 3649 -4430
rect 3683 -4464 3702 -4430
rect 3633 -4498 3702 -4464
rect 3633 -4532 3649 -4498
rect 3683 -4532 3702 -4498
rect 3633 -4582 3702 -4532
rect 3084 -4693 3087 -4659
rect 3121 -4693 3237 -4659
rect 3084 -4709 3237 -4693
rect 3271 -4659 3443 -4644
rect 3508 -4616 3702 -4582
rect 3736 -4452 3794 -4381
rect 3736 -4486 3748 -4452
rect 3782 -4486 3794 -4452
rect 3736 -4545 3794 -4486
rect 3736 -4579 3748 -4545
rect 3782 -4579 3794 -4545
rect 3736 -4614 3794 -4579
rect 3828 -4423 4162 -4381
rect 3828 -4457 3846 -4423
rect 3880 -4457 4110 -4423
rect 4144 -4457 4162 -4423
rect 3828 -4525 4162 -4457
rect 3828 -4559 3846 -4525
rect 3880 -4559 4110 -4525
rect 4144 -4559 4162 -4525
rect 3828 -4599 4162 -4559
rect 4196 -4452 4254 -4381
rect 4196 -4486 4208 -4452
rect 4242 -4486 4254 -4452
rect 4196 -4545 4254 -4486
rect 4196 -4579 4208 -4545
rect 4242 -4579 4254 -4545
rect 3508 -4645 3578 -4616
rect 3271 -4693 3287 -4659
rect 3321 -4693 3443 -4659
rect 3271 -4694 3443 -4693
rect 3203 -4728 3237 -4709
rect 3203 -4762 3321 -4728
rect 3000 -4804 3081 -4780
rect 3000 -4838 3033 -4804
rect 3067 -4838 3081 -4804
rect 3000 -4857 3081 -4838
rect 3115 -4804 3181 -4788
rect 3115 -4838 3131 -4804
rect 3165 -4838 3181 -4804
rect 3115 -4891 3181 -4838
rect 3271 -4804 3321 -4762
rect 3271 -4838 3287 -4804
rect 3271 -4857 3321 -4838
rect 3373 -4804 3443 -4694
rect 3492 -4659 3578 -4645
rect 3492 -4693 3508 -4659
rect 3542 -4693 3578 -4659
rect 3612 -4652 3702 -4650
rect 3612 -4693 3628 -4652
rect 3662 -4693 3702 -4652
rect 3828 -4669 3978 -4599
rect 4196 -4614 4254 -4579
rect 4288 -4423 4990 -4381
rect 4288 -4457 4306 -4423
rect 4340 -4457 4938 -4423
rect 4972 -4457 4990 -4423
rect 4288 -4525 4990 -4457
rect 4288 -4559 4306 -4525
rect 4340 -4559 4938 -4525
rect 4972 -4559 4990 -4525
rect 4288 -4599 4990 -4559
rect 3492 -4703 3578 -4693
rect 3828 -4703 3848 -4669
rect 3882 -4703 3978 -4669
rect 4012 -4667 4108 -4633
rect 4142 -4667 4162 -4633
rect 3508 -4727 3578 -4703
rect 3508 -4761 3702 -4727
rect 4012 -4737 4162 -4667
rect 3373 -4838 3392 -4804
rect 3426 -4838 3443 -4804
rect 3373 -4857 3443 -4838
rect 3536 -4804 3602 -4795
rect 3536 -4838 3552 -4804
rect 3586 -4838 3602 -4804
rect 3536 -4891 3602 -4838
rect 3636 -4804 3702 -4761
rect 3636 -4838 3649 -4804
rect 3683 -4838 3702 -4804
rect 3636 -4857 3702 -4838
rect 3736 -4763 3794 -4746
rect 3736 -4797 3748 -4763
rect 3782 -4797 3794 -4763
rect 3736 -4891 3794 -4797
rect 3828 -4789 4162 -4737
rect 4288 -4667 4366 -4633
rect 4400 -4667 4465 -4633
rect 4499 -4667 4564 -4633
rect 4598 -4667 4618 -4633
rect 4288 -4737 4618 -4667
rect 4652 -4669 4990 -4599
rect 5024 -4452 5082 -4381
rect 5024 -4486 5036 -4452
rect 5070 -4486 5082 -4452
rect 5024 -4545 5082 -4486
rect 5024 -4579 5036 -4545
rect 5070 -4579 5082 -4545
rect 5024 -4614 5082 -4579
rect 5116 -4423 5450 -4381
rect 5116 -4457 5134 -4423
rect 5168 -4457 5398 -4423
rect 5432 -4457 5450 -4423
rect 5116 -4525 5450 -4457
rect 5116 -4559 5134 -4525
rect 5168 -4559 5398 -4525
rect 5432 -4559 5450 -4525
rect 5116 -4599 5450 -4559
rect 5484 -4452 5542 -4381
rect 5484 -4486 5496 -4452
rect 5530 -4486 5542 -4452
rect 5484 -4545 5542 -4486
rect 5484 -4579 5496 -4545
rect 5530 -4579 5542 -4545
rect 4652 -4703 4672 -4669
rect 4706 -4703 4775 -4669
rect 4809 -4703 4878 -4669
rect 4912 -4703 4990 -4669
rect 5116 -4669 5266 -4599
rect 5484 -4614 5542 -4579
rect 5576 -4431 5657 -4415
rect 5576 -4465 5609 -4431
rect 5643 -4465 5657 -4431
rect 5576 -4499 5657 -4465
rect 5576 -4533 5609 -4499
rect 5643 -4533 5657 -4499
rect 5576 -4570 5657 -4533
rect 5691 -4430 5757 -4381
rect 5691 -4464 5707 -4430
rect 5741 -4464 5757 -4430
rect 5691 -4498 5757 -4464
rect 5691 -4532 5707 -4498
rect 5741 -4532 5757 -4498
rect 5691 -4541 5757 -4532
rect 5847 -4431 5897 -4415
rect 5847 -4465 5863 -4431
rect 5847 -4499 5897 -4465
rect 5847 -4533 5863 -4499
rect 5116 -4703 5136 -4669
rect 5170 -4703 5266 -4669
rect 5300 -4667 5396 -4633
rect 5430 -4667 5450 -4633
rect 5300 -4737 5450 -4667
rect 3828 -4823 3846 -4789
rect 3880 -4823 4110 -4789
rect 4144 -4823 4162 -4789
rect 3828 -4891 4162 -4823
rect 4196 -4763 4254 -4746
rect 4196 -4797 4208 -4763
rect 4242 -4797 4254 -4763
rect 4196 -4891 4254 -4797
rect 4288 -4796 4990 -4737
rect 4288 -4830 4306 -4796
rect 4340 -4830 4938 -4796
rect 4972 -4830 4990 -4796
rect 4288 -4891 4990 -4830
rect 5024 -4763 5082 -4746
rect 5024 -4797 5036 -4763
rect 5070 -4797 5082 -4763
rect 5024 -4891 5082 -4797
rect 5116 -4789 5450 -4737
rect 5576 -4652 5626 -4570
rect 5847 -4575 5897 -4533
rect 5779 -4609 5897 -4575
rect 5949 -4430 6019 -4415
rect 5949 -4464 5967 -4430
rect 6001 -4464 6019 -4430
rect 5949 -4498 6019 -4464
rect 5949 -4532 5967 -4498
rect 6001 -4532 6019 -4498
rect 5779 -4643 5813 -4609
rect 5576 -4686 5588 -4652
rect 5622 -4686 5626 -4652
rect 5116 -4823 5134 -4789
rect 5168 -4823 5398 -4789
rect 5432 -4823 5450 -4789
rect 5116 -4891 5450 -4823
rect 5484 -4763 5542 -4746
rect 5484 -4797 5496 -4763
rect 5530 -4797 5542 -4763
rect 5484 -4891 5542 -4797
rect 5576 -4780 5626 -4686
rect 5660 -4659 5813 -4643
rect 5949 -4644 6019 -4532
rect 6109 -4430 6175 -4381
rect 6109 -4464 6125 -4430
rect 6159 -4464 6175 -4430
rect 6109 -4498 6175 -4464
rect 6109 -4532 6125 -4498
rect 6159 -4532 6175 -4498
rect 6109 -4548 6175 -4532
rect 6209 -4430 6278 -4415
rect 6209 -4464 6225 -4430
rect 6259 -4464 6278 -4430
rect 6209 -4498 6278 -4464
rect 6209 -4532 6225 -4498
rect 6259 -4532 6278 -4498
rect 6209 -4582 6278 -4532
rect 5660 -4693 5663 -4659
rect 5697 -4693 5813 -4659
rect 5660 -4709 5813 -4693
rect 5847 -4659 6019 -4644
rect 6084 -4616 6278 -4582
rect 6312 -4452 6370 -4381
rect 6312 -4486 6324 -4452
rect 6358 -4486 6370 -4452
rect 6312 -4545 6370 -4486
rect 6312 -4579 6324 -4545
rect 6358 -4579 6370 -4545
rect 6312 -4614 6370 -4579
rect 6404 -4423 6738 -4381
rect 6404 -4457 6422 -4423
rect 6456 -4457 6686 -4423
rect 6720 -4457 6738 -4423
rect 6404 -4525 6738 -4457
rect 6404 -4559 6422 -4525
rect 6456 -4559 6686 -4525
rect 6720 -4559 6738 -4525
rect 6404 -4599 6738 -4559
rect 6772 -4452 6830 -4381
rect 6772 -4486 6784 -4452
rect 6818 -4486 6830 -4452
rect 6772 -4545 6830 -4486
rect 6772 -4579 6784 -4545
rect 6818 -4579 6830 -4545
rect 6084 -4645 6154 -4616
rect 5847 -4693 5863 -4659
rect 5897 -4693 6019 -4659
rect 5847 -4694 6019 -4693
rect 5779 -4728 5813 -4709
rect 5779 -4762 5897 -4728
rect 5576 -4804 5657 -4780
rect 5576 -4838 5609 -4804
rect 5643 -4838 5657 -4804
rect 5576 -4857 5657 -4838
rect 5691 -4804 5757 -4788
rect 5691 -4838 5707 -4804
rect 5741 -4838 5757 -4804
rect 5691 -4891 5757 -4838
rect 5847 -4804 5897 -4762
rect 5847 -4838 5863 -4804
rect 5847 -4857 5897 -4838
rect 5949 -4804 6019 -4694
rect 6068 -4659 6154 -4645
rect 6068 -4693 6084 -4659
rect 6118 -4693 6154 -4659
rect 6188 -4652 6278 -4650
rect 6188 -4686 6202 -4652
rect 6236 -4659 6278 -4652
rect 6188 -4693 6204 -4686
rect 6238 -4693 6278 -4659
rect 6404 -4669 6554 -4599
rect 6772 -4614 6830 -4579
rect 6864 -4423 7566 -4381
rect 6864 -4457 6882 -4423
rect 6916 -4457 7514 -4423
rect 7548 -4457 7566 -4423
rect 6864 -4525 7566 -4457
rect 6864 -4559 6882 -4525
rect 6916 -4559 7514 -4525
rect 7548 -4559 7566 -4525
rect 6864 -4599 7566 -4559
rect 6068 -4703 6154 -4693
rect 6404 -4703 6424 -4669
rect 6458 -4703 6554 -4669
rect 6588 -4667 6684 -4633
rect 6718 -4667 6738 -4633
rect 6084 -4727 6154 -4703
rect 6084 -4761 6278 -4727
rect 6588 -4737 6738 -4667
rect 5949 -4838 5968 -4804
rect 6002 -4838 6019 -4804
rect 5949 -4857 6019 -4838
rect 6112 -4804 6178 -4795
rect 6112 -4838 6128 -4804
rect 6162 -4838 6178 -4804
rect 6112 -4891 6178 -4838
rect 6212 -4804 6278 -4761
rect 6212 -4838 6225 -4804
rect 6259 -4838 6278 -4804
rect 6212 -4857 6278 -4838
rect 6312 -4763 6370 -4746
rect 6312 -4797 6324 -4763
rect 6358 -4797 6370 -4763
rect 6312 -4891 6370 -4797
rect 6404 -4789 6738 -4737
rect 6864 -4667 6942 -4633
rect 6976 -4667 7041 -4633
rect 7075 -4667 7140 -4633
rect 7174 -4667 7194 -4633
rect 6864 -4737 7194 -4667
rect 7228 -4669 7566 -4599
rect 7600 -4452 7658 -4381
rect 7600 -4486 7612 -4452
rect 7646 -4486 7658 -4452
rect 7600 -4545 7658 -4486
rect 7600 -4579 7612 -4545
rect 7646 -4579 7658 -4545
rect 7600 -4614 7658 -4579
rect 7692 -4423 8026 -4381
rect 7692 -4457 7710 -4423
rect 7744 -4457 7974 -4423
rect 8008 -4457 8026 -4423
rect 7692 -4525 8026 -4457
rect 7692 -4559 7710 -4525
rect 7744 -4559 7974 -4525
rect 8008 -4559 8026 -4525
rect 7692 -4599 8026 -4559
rect 8060 -4452 8118 -4381
rect 8060 -4486 8072 -4452
rect 8106 -4486 8118 -4452
rect 8060 -4545 8118 -4486
rect 8060 -4579 8072 -4545
rect 8106 -4579 8118 -4545
rect 7228 -4703 7248 -4669
rect 7282 -4703 7351 -4669
rect 7385 -4703 7454 -4669
rect 7488 -4703 7566 -4669
rect 7692 -4669 7842 -4599
rect 8060 -4614 8118 -4579
rect 8152 -4431 8233 -4415
rect 8152 -4465 8185 -4431
rect 8219 -4465 8233 -4431
rect 8152 -4499 8233 -4465
rect 8152 -4533 8185 -4499
rect 8219 -4533 8233 -4499
rect 8152 -4570 8233 -4533
rect 8267 -4430 8333 -4381
rect 8267 -4464 8283 -4430
rect 8317 -4464 8333 -4430
rect 8267 -4498 8333 -4464
rect 8267 -4532 8283 -4498
rect 8317 -4532 8333 -4498
rect 8267 -4541 8333 -4532
rect 8423 -4431 8473 -4415
rect 8423 -4465 8439 -4431
rect 8423 -4499 8473 -4465
rect 8423 -4533 8439 -4499
rect 7692 -4703 7712 -4669
rect 7746 -4703 7842 -4669
rect 7876 -4667 7972 -4633
rect 8006 -4667 8026 -4633
rect 7876 -4737 8026 -4667
rect 6404 -4823 6422 -4789
rect 6456 -4823 6686 -4789
rect 6720 -4823 6738 -4789
rect 6404 -4891 6738 -4823
rect 6772 -4763 6830 -4746
rect 6772 -4797 6784 -4763
rect 6818 -4797 6830 -4763
rect 6772 -4891 6830 -4797
rect 6864 -4796 7566 -4737
rect 6864 -4830 6882 -4796
rect 6916 -4830 7514 -4796
rect 7548 -4830 7566 -4796
rect 6864 -4891 7566 -4830
rect 7600 -4763 7658 -4746
rect 7600 -4797 7612 -4763
rect 7646 -4797 7658 -4763
rect 7600 -4891 7658 -4797
rect 7692 -4789 8026 -4737
rect 8152 -4652 8202 -4570
rect 8423 -4575 8473 -4533
rect 8355 -4609 8473 -4575
rect 8525 -4430 8595 -4415
rect 8525 -4464 8543 -4430
rect 8577 -4464 8595 -4430
rect 8525 -4498 8595 -4464
rect 8525 -4532 8543 -4498
rect 8577 -4532 8595 -4498
rect 8355 -4643 8389 -4609
rect 8152 -4686 8162 -4652
rect 8196 -4686 8202 -4652
rect 7692 -4823 7710 -4789
rect 7744 -4823 7974 -4789
rect 8008 -4823 8026 -4789
rect 7692 -4891 8026 -4823
rect 8060 -4763 8118 -4746
rect 8060 -4797 8072 -4763
rect 8106 -4797 8118 -4763
rect 8060 -4891 8118 -4797
rect 8152 -4780 8202 -4686
rect 8236 -4659 8389 -4643
rect 8525 -4644 8595 -4532
rect 8685 -4430 8751 -4381
rect 8685 -4464 8701 -4430
rect 8735 -4464 8751 -4430
rect 8685 -4498 8751 -4464
rect 8685 -4532 8701 -4498
rect 8735 -4532 8751 -4498
rect 8685 -4548 8751 -4532
rect 8785 -4430 8854 -4415
rect 8785 -4464 8801 -4430
rect 8835 -4464 8854 -4430
rect 8785 -4498 8854 -4464
rect 8785 -4532 8801 -4498
rect 8835 -4532 8854 -4498
rect 8785 -4582 8854 -4532
rect 8236 -4693 8239 -4659
rect 8273 -4693 8389 -4659
rect 8236 -4709 8389 -4693
rect 8423 -4659 8595 -4644
rect 8660 -4616 8854 -4582
rect 8888 -4452 8946 -4381
rect 8888 -4486 8900 -4452
rect 8934 -4486 8946 -4452
rect 8888 -4545 8946 -4486
rect 8888 -4579 8900 -4545
rect 8934 -4579 8946 -4545
rect 8888 -4614 8946 -4579
rect 8980 -4423 9314 -4381
rect 8980 -4457 8998 -4423
rect 9032 -4457 9262 -4423
rect 9296 -4457 9314 -4423
rect 8980 -4525 9314 -4457
rect 8980 -4559 8998 -4525
rect 9032 -4559 9262 -4525
rect 9296 -4559 9314 -4525
rect 8980 -4599 9314 -4559
rect 9348 -4452 9406 -4381
rect 9348 -4486 9360 -4452
rect 9394 -4486 9406 -4452
rect 9348 -4545 9406 -4486
rect 9348 -4579 9360 -4545
rect 9394 -4579 9406 -4545
rect 8660 -4645 8730 -4616
rect 8423 -4693 8439 -4659
rect 8473 -4693 8595 -4659
rect 8423 -4694 8595 -4693
rect 8355 -4728 8389 -4709
rect 8355 -4762 8473 -4728
rect 8152 -4804 8233 -4780
rect 8152 -4838 8185 -4804
rect 8219 -4838 8233 -4804
rect 8152 -4857 8233 -4838
rect 8267 -4804 8333 -4788
rect 8267 -4838 8283 -4804
rect 8317 -4838 8333 -4804
rect 8267 -4891 8333 -4838
rect 8423 -4804 8473 -4762
rect 8423 -4838 8439 -4804
rect 8423 -4857 8473 -4838
rect 8525 -4804 8595 -4694
rect 8644 -4659 8730 -4645
rect 8644 -4693 8660 -4659
rect 8694 -4693 8730 -4659
rect 8764 -4652 8854 -4650
rect 8764 -4686 8776 -4652
rect 8810 -4659 8854 -4652
rect 8764 -4693 8780 -4686
rect 8814 -4693 8854 -4659
rect 8980 -4669 9130 -4599
rect 9348 -4614 9406 -4579
rect 9440 -4423 10142 -4381
rect 9440 -4457 9458 -4423
rect 9492 -4457 10090 -4423
rect 10124 -4457 10142 -4423
rect 9440 -4525 10142 -4457
rect 9440 -4559 9458 -4525
rect 9492 -4559 10090 -4525
rect 10124 -4559 10142 -4525
rect 9440 -4599 10142 -4559
rect 8644 -4703 8730 -4693
rect 8980 -4703 9000 -4669
rect 9034 -4703 9130 -4669
rect 9164 -4667 9260 -4633
rect 9294 -4667 9314 -4633
rect 8660 -4727 8730 -4703
rect 8660 -4761 8854 -4727
rect 9164 -4737 9314 -4667
rect 8525 -4838 8544 -4804
rect 8578 -4838 8595 -4804
rect 8525 -4857 8595 -4838
rect 8688 -4804 8754 -4795
rect 8688 -4838 8704 -4804
rect 8738 -4838 8754 -4804
rect 8688 -4891 8754 -4838
rect 8788 -4804 8854 -4761
rect 8788 -4838 8801 -4804
rect 8835 -4838 8854 -4804
rect 8788 -4857 8854 -4838
rect 8888 -4763 8946 -4746
rect 8888 -4797 8900 -4763
rect 8934 -4797 8946 -4763
rect 8888 -4891 8946 -4797
rect 8980 -4789 9314 -4737
rect 9440 -4667 9518 -4633
rect 9552 -4667 9617 -4633
rect 9651 -4667 9716 -4633
rect 9750 -4667 9770 -4633
rect 9440 -4737 9770 -4667
rect 9804 -4669 10142 -4599
rect 10176 -4452 10234 -4381
rect 10176 -4486 10188 -4452
rect 10222 -4486 10234 -4452
rect 10176 -4545 10234 -4486
rect 10176 -4579 10188 -4545
rect 10222 -4579 10234 -4545
rect 10176 -4614 10234 -4579
rect 10360 -4423 10694 -4381
rect 10360 -4457 10378 -4423
rect 10412 -4457 10642 -4423
rect 10676 -4457 10694 -4423
rect 10360 -4525 10694 -4457
rect 10360 -4559 10378 -4525
rect 10412 -4559 10642 -4525
rect 10676 -4559 10694 -4525
rect 10360 -4599 10694 -4559
rect 10728 -4431 10809 -4415
rect 10728 -4465 10761 -4431
rect 10795 -4465 10809 -4431
rect 10728 -4499 10809 -4465
rect 10728 -4533 10761 -4499
rect 10795 -4533 10809 -4499
rect 10728 -4570 10809 -4533
rect 10843 -4430 10909 -4381
rect 10843 -4464 10859 -4430
rect 10893 -4464 10909 -4430
rect 10843 -4498 10909 -4464
rect 10843 -4532 10859 -4498
rect 10893 -4532 10909 -4498
rect 10843 -4541 10909 -4532
rect 10999 -4431 11049 -4415
rect 10999 -4465 11015 -4431
rect 10999 -4499 11049 -4465
rect 10999 -4533 11015 -4499
rect 9804 -4703 9824 -4669
rect 9858 -4703 9927 -4669
rect 9961 -4703 10030 -4669
rect 10064 -4703 10142 -4669
rect 10360 -4669 10510 -4599
rect 10360 -4703 10380 -4669
rect 10414 -4703 10510 -4669
rect 10544 -4667 10640 -4633
rect 10674 -4667 10694 -4633
rect 10544 -4737 10694 -4667
rect 8980 -4823 8998 -4789
rect 9032 -4823 9262 -4789
rect 9296 -4823 9314 -4789
rect 8980 -4891 9314 -4823
rect 9348 -4763 9406 -4746
rect 9348 -4797 9360 -4763
rect 9394 -4797 9406 -4763
rect 9348 -4891 9406 -4797
rect 9440 -4796 10142 -4737
rect 9440 -4830 9458 -4796
rect 9492 -4830 10090 -4796
rect 10124 -4830 10142 -4796
rect 9440 -4891 10142 -4830
rect 10176 -4763 10234 -4746
rect 10176 -4797 10188 -4763
rect 10222 -4797 10234 -4763
rect 10176 -4891 10234 -4797
rect 10360 -4789 10694 -4737
rect 10360 -4823 10378 -4789
rect 10412 -4823 10642 -4789
rect 10676 -4823 10694 -4789
rect 10360 -4891 10694 -4823
rect 10728 -4652 10778 -4570
rect 10999 -4575 11049 -4533
rect 10931 -4609 11049 -4575
rect 11101 -4430 11171 -4415
rect 11101 -4464 11119 -4430
rect 11153 -4464 11171 -4430
rect 11101 -4498 11171 -4464
rect 11101 -4532 11119 -4498
rect 11153 -4532 11171 -4498
rect 10931 -4643 10965 -4609
rect 10728 -4686 10736 -4652
rect 10770 -4686 10778 -4652
rect 10728 -4780 10778 -4686
rect 10812 -4659 10965 -4643
rect 11101 -4644 11171 -4532
rect 11261 -4430 11327 -4381
rect 11261 -4464 11277 -4430
rect 11311 -4464 11327 -4430
rect 11261 -4498 11327 -4464
rect 11261 -4532 11277 -4498
rect 11311 -4532 11327 -4498
rect 11261 -4548 11327 -4532
rect 11361 -4430 11430 -4415
rect 11361 -4464 11377 -4430
rect 11411 -4464 11430 -4430
rect 11361 -4498 11430 -4464
rect 11361 -4532 11377 -4498
rect 11411 -4532 11430 -4498
rect 11361 -4582 11430 -4532
rect 10812 -4693 10815 -4659
rect 10849 -4693 10965 -4659
rect 10812 -4709 10965 -4693
rect 10999 -4659 11171 -4644
rect 11236 -4616 11430 -4582
rect 11464 -4452 11522 -4381
rect 11464 -4486 11476 -4452
rect 11510 -4486 11522 -4452
rect 11464 -4545 11522 -4486
rect 11464 -4579 11476 -4545
rect 11510 -4579 11522 -4545
rect 11464 -4614 11522 -4579
rect 11648 -4423 11982 -4381
rect 11648 -4457 11666 -4423
rect 11700 -4457 11930 -4423
rect 11964 -4457 11982 -4423
rect 11648 -4525 11982 -4457
rect 11648 -4559 11666 -4525
rect 11700 -4559 11930 -4525
rect 11964 -4559 11982 -4525
rect 11648 -4599 11982 -4559
rect 13580 -4452 13638 -4381
rect 13580 -4486 13592 -4452
rect 13626 -4486 13638 -4452
rect 13580 -4545 13638 -4486
rect 13674 -4423 13733 -4381
rect 13674 -4457 13690 -4423
rect 13724 -4457 13733 -4423
rect 13674 -4491 13733 -4457
rect 13674 -4525 13690 -4491
rect 13724 -4525 13733 -4491
rect 13674 -4543 13733 -4525
rect 13769 -4431 13818 -4415
rect 13769 -4465 13776 -4431
rect 13810 -4465 13818 -4431
rect 13769 -4499 13818 -4465
rect 13769 -4533 13776 -4499
rect 13810 -4533 13818 -4499
rect 13580 -4579 13592 -4545
rect 13626 -4579 13638 -4545
rect 11236 -4645 11306 -4616
rect 10999 -4693 11015 -4659
rect 11049 -4693 11171 -4659
rect 10999 -4694 11171 -4693
rect 10931 -4728 10965 -4709
rect 10931 -4762 11049 -4728
rect 10728 -4804 10809 -4780
rect 10728 -4838 10761 -4804
rect 10795 -4838 10809 -4804
rect 10728 -4857 10809 -4838
rect 10843 -4804 10909 -4788
rect 10843 -4838 10859 -4804
rect 10893 -4838 10909 -4804
rect 10843 -4891 10909 -4838
rect 10999 -4804 11049 -4762
rect 10999 -4838 11015 -4804
rect 10999 -4857 11049 -4838
rect 11101 -4804 11171 -4694
rect 11220 -4659 11306 -4645
rect 11220 -4693 11236 -4659
rect 11270 -4693 11306 -4659
rect 11340 -4657 11430 -4650
rect 11340 -4659 11384 -4657
rect 11340 -4693 11356 -4659
rect 11418 -4691 11430 -4657
rect 11390 -4693 11430 -4691
rect 11648 -4669 11798 -4599
rect 13580 -4614 13638 -4579
rect 11220 -4703 11306 -4693
rect 11648 -4703 11668 -4669
rect 11702 -4703 11798 -4669
rect 11832 -4667 11928 -4633
rect 11962 -4667 11982 -4633
rect 13769 -4643 13818 -4533
rect 13853 -4423 13905 -4381
rect 14025 -4382 15280 -4381
rect 13853 -4457 13862 -4423
rect 13896 -4457 13905 -4423
rect 13853 -4491 13905 -4457
rect 13853 -4525 13862 -4491
rect 13896 -4525 13905 -4491
rect 13853 -4543 13905 -4525
rect 13941 -4439 13991 -4416
rect 13941 -4473 13948 -4439
rect 13982 -4473 13991 -4439
rect 13941 -4507 13991 -4473
rect 13941 -4541 13948 -4507
rect 13982 -4541 13991 -4507
rect 14025 -4423 14077 -4382
rect 14025 -4457 14034 -4423
rect 14068 -4457 14077 -4423
rect 14025 -4491 14077 -4457
rect 14025 -4525 14034 -4491
rect 14068 -4525 14077 -4491
rect 14025 -4541 14077 -4525
rect 14111 -4467 14163 -4416
rect 14111 -4501 14120 -4467
rect 14154 -4501 14163 -4467
rect 13941 -4643 13991 -4541
rect 14111 -4553 14163 -4501
rect 14197 -4447 14249 -4382
rect 14197 -4481 14206 -4447
rect 14240 -4481 14249 -4447
rect 14197 -4527 14249 -4481
rect 14283 -4467 14335 -4416
rect 14283 -4501 14292 -4467
rect 14326 -4501 14335 -4467
rect 14111 -4587 14120 -4553
rect 14154 -4561 14163 -4553
rect 14283 -4553 14335 -4501
rect 14369 -4447 14421 -4382
rect 14369 -4481 14378 -4447
rect 14412 -4481 14421 -4447
rect 14369 -4527 14421 -4481
rect 14455 -4467 14507 -4416
rect 14455 -4501 14464 -4467
rect 14498 -4501 14507 -4467
rect 14283 -4561 14292 -4553
rect 14154 -4587 14292 -4561
rect 14326 -4561 14335 -4553
rect 14455 -4553 14507 -4501
rect 14541 -4447 14593 -4382
rect 14541 -4481 14550 -4447
rect 14584 -4481 14593 -4447
rect 14541 -4527 14593 -4481
rect 14627 -4467 14679 -4416
rect 14627 -4501 14636 -4467
rect 14670 -4501 14679 -4467
rect 14455 -4561 14464 -4553
rect 14326 -4587 14464 -4561
rect 14498 -4561 14507 -4553
rect 14627 -4553 14679 -4501
rect 14713 -4447 14762 -4382
rect 14713 -4481 14722 -4447
rect 14756 -4481 14762 -4447
rect 14713 -4527 14762 -4481
rect 14796 -4467 14848 -4416
rect 14796 -4501 14807 -4467
rect 14841 -4501 14848 -4467
rect 14627 -4561 14636 -4553
rect 14498 -4587 14636 -4561
rect 14670 -4561 14679 -4553
rect 14796 -4553 14848 -4501
rect 14885 -4447 14934 -4382
rect 14885 -4481 14893 -4447
rect 14927 -4481 14934 -4447
rect 14885 -4527 14934 -4481
rect 14968 -4467 15020 -4416
rect 14968 -4501 14979 -4467
rect 15013 -4501 15020 -4467
rect 14796 -4561 14807 -4553
rect 14670 -4587 14807 -4561
rect 14841 -4561 14848 -4553
rect 14968 -4553 15020 -4501
rect 15057 -4447 15106 -4382
rect 15057 -4481 15065 -4447
rect 15099 -4481 15106 -4447
rect 15057 -4527 15106 -4481
rect 15140 -4467 15192 -4416
rect 15140 -4501 15151 -4467
rect 15185 -4501 15192 -4467
rect 14968 -4561 14979 -4553
rect 14841 -4587 14979 -4561
rect 15013 -4561 15020 -4553
rect 15140 -4553 15192 -4501
rect 15229 -4447 15280 -4382
rect 15229 -4481 15237 -4447
rect 15271 -4481 15280 -4447
rect 15229 -4527 15280 -4481
rect 15314 -4467 15372 -4416
rect 15314 -4501 15323 -4467
rect 15357 -4501 15372 -4467
rect 15140 -4561 15151 -4553
rect 15013 -4587 15151 -4561
rect 15185 -4564 15192 -4553
rect 15314 -4553 15372 -4501
rect 15406 -4447 15460 -4381
rect 15406 -4481 15409 -4447
rect 15443 -4481 15460 -4447
rect 15406 -4530 15460 -4481
rect 15512 -4452 15570 -4381
rect 15512 -4486 15524 -4452
rect 15558 -4486 15570 -4452
rect 15314 -4564 15323 -4553
rect 15185 -4587 15323 -4564
rect 15357 -4564 15372 -4553
rect 15512 -4545 15570 -4486
rect 15357 -4587 15460 -4564
rect 14111 -4606 15460 -4587
rect 14111 -4609 15248 -4606
rect 15227 -4640 15248 -4609
rect 15282 -4640 15341 -4606
rect 15375 -4640 15460 -4606
rect 15512 -4579 15524 -4545
rect 15558 -4579 15570 -4545
rect 15512 -4614 15570 -4579
rect 15605 -4423 16674 -4381
rect 15605 -4457 15622 -4423
rect 15656 -4457 16622 -4423
rect 16656 -4457 16674 -4423
rect 15605 -4525 16674 -4457
rect 15605 -4559 15622 -4525
rect 15656 -4559 16622 -4525
rect 16656 -4559 16674 -4525
rect 15605 -4599 16674 -4559
rect 11236 -4727 11306 -4703
rect 11236 -4761 11430 -4727
rect 11832 -4737 11982 -4667
rect 11101 -4838 11120 -4804
rect 11154 -4838 11171 -4804
rect 11101 -4857 11171 -4838
rect 11264 -4804 11330 -4795
rect 11264 -4838 11280 -4804
rect 11314 -4838 11330 -4804
rect 11264 -4891 11330 -4838
rect 11364 -4804 11430 -4761
rect 11364 -4838 11377 -4804
rect 11411 -4838 11430 -4804
rect 11364 -4857 11430 -4838
rect 11464 -4763 11522 -4746
rect 11464 -4797 11476 -4763
rect 11510 -4797 11522 -4763
rect 11464 -4891 11522 -4797
rect 11648 -4789 11982 -4737
rect 13672 -4659 13735 -4643
rect 13672 -4686 13692 -4659
rect 13672 -4720 13685 -4686
rect 13726 -4693 13735 -4659
rect 13719 -4720 13735 -4693
rect 11648 -4823 11666 -4789
rect 11700 -4823 11930 -4789
rect 11964 -4823 11982 -4789
rect 11648 -4891 11982 -4823
rect 13580 -4763 13638 -4746
rect 13672 -4755 13735 -4720
rect 13769 -4659 15193 -4643
rect 13769 -4693 14119 -4659
rect 14153 -4693 14187 -4659
rect 14221 -4693 14255 -4659
rect 14289 -4693 14323 -4659
rect 14357 -4693 14391 -4659
rect 14425 -4693 14459 -4659
rect 14493 -4693 14527 -4659
rect 14561 -4693 14595 -4659
rect 14629 -4693 14663 -4659
rect 14697 -4693 14731 -4659
rect 14765 -4693 14799 -4659
rect 14833 -4693 14867 -4659
rect 14901 -4693 14935 -4659
rect 14969 -4693 15003 -4659
rect 15037 -4693 15071 -4659
rect 15105 -4693 15139 -4659
rect 15173 -4693 15193 -4659
rect 13580 -4797 13592 -4763
rect 13626 -4797 13638 -4763
rect 13580 -4891 13638 -4797
rect 13672 -4815 13733 -4789
rect 13672 -4849 13690 -4815
rect 13724 -4849 13733 -4815
rect 13672 -4891 13733 -4849
rect 13769 -4802 13819 -4693
rect 13769 -4836 13776 -4802
rect 13810 -4836 13819 -4802
rect 13769 -4855 13819 -4836
rect 13853 -4802 13905 -4786
rect 13853 -4836 13862 -4802
rect 13896 -4836 13905 -4802
rect 13853 -4891 13905 -4836
rect 13941 -4802 13991 -4693
rect 15227 -4701 15460 -4640
rect 15227 -4702 15340 -4701
rect 15227 -4727 15248 -4702
rect 14111 -4736 15248 -4727
rect 15282 -4735 15340 -4702
rect 15374 -4735 15460 -4701
rect 15605 -4669 16124 -4599
rect 15605 -4703 15686 -4669
rect 15720 -4703 15814 -4669
rect 15848 -4703 15942 -4669
rect 15976 -4703 16070 -4669
rect 16104 -4703 16124 -4669
rect 16158 -4667 16178 -4633
rect 16212 -4667 16306 -4633
rect 16340 -4667 16434 -4633
rect 16468 -4667 16562 -4633
rect 16596 -4667 16674 -4633
rect 15282 -4736 15460 -4735
rect 14111 -4761 15460 -4736
rect 16158 -4737 16674 -4667
rect 13941 -4836 13948 -4802
rect 13982 -4836 13991 -4802
rect 13941 -4855 13991 -4836
rect 14025 -4802 14077 -4779
rect 14025 -4836 14034 -4802
rect 14068 -4836 14077 -4802
rect 14025 -4891 14077 -4836
rect 14111 -4802 14163 -4761
rect 14111 -4836 14120 -4802
rect 14154 -4836 14163 -4802
rect 14111 -4852 14163 -4836
rect 14197 -4811 14249 -4795
rect 14197 -4845 14206 -4811
rect 14240 -4845 14249 -4811
rect 14197 -4891 14249 -4845
rect 14283 -4802 14335 -4761
rect 14283 -4836 14292 -4802
rect 14326 -4836 14335 -4802
rect 14283 -4852 14335 -4836
rect 14369 -4811 14421 -4795
rect 14369 -4845 14378 -4811
rect 14412 -4845 14421 -4811
rect 14369 -4891 14421 -4845
rect 14455 -4802 14507 -4761
rect 14455 -4836 14464 -4802
rect 14498 -4836 14507 -4802
rect 14455 -4852 14507 -4836
rect 14541 -4811 14590 -4795
rect 14541 -4845 14550 -4811
rect 14584 -4845 14590 -4811
rect 14541 -4891 14590 -4845
rect 14624 -4802 14679 -4761
rect 14624 -4836 14636 -4802
rect 14670 -4836 14679 -4802
rect 14624 -4852 14679 -4836
rect 14713 -4811 14762 -4795
rect 14713 -4845 14722 -4811
rect 14756 -4845 14762 -4811
rect 14713 -4891 14762 -4845
rect 14796 -4802 14848 -4761
rect 14796 -4836 14807 -4802
rect 14841 -4836 14848 -4802
rect 14796 -4852 14848 -4836
rect 14884 -4811 14934 -4795
rect 14884 -4845 14893 -4811
rect 14927 -4845 14934 -4811
rect 14884 -4891 14934 -4845
rect 14968 -4802 15020 -4761
rect 14968 -4836 14979 -4802
rect 15013 -4836 15020 -4802
rect 14968 -4852 15020 -4836
rect 15056 -4811 15106 -4795
rect 15056 -4845 15065 -4811
rect 15099 -4845 15106 -4811
rect 15056 -4891 15106 -4845
rect 15140 -4802 15192 -4761
rect 15140 -4836 15151 -4802
rect 15185 -4836 15192 -4802
rect 15140 -4852 15192 -4836
rect 15228 -4811 15280 -4795
rect 15228 -4845 15237 -4811
rect 15271 -4845 15280 -4811
rect 15228 -4891 15280 -4845
rect 15314 -4802 15366 -4761
rect 15512 -4763 15570 -4746
rect 15314 -4836 15323 -4802
rect 15357 -4836 15366 -4802
rect 15314 -4852 15366 -4836
rect 15400 -4811 15460 -4795
rect 15400 -4845 15409 -4811
rect 15443 -4845 15460 -4811
rect 15400 -4891 15460 -4845
rect 15512 -4797 15524 -4763
rect 15558 -4797 15570 -4763
rect 15512 -4891 15570 -4797
rect 15605 -4796 16674 -4737
rect 15605 -4830 15622 -4796
rect 15656 -4830 16622 -4796
rect 16656 -4830 16674 -4796
rect 15605 -4891 16674 -4830
rect -2997 -4925 -2968 -4891
rect -2934 -4925 -2876 -4891
rect -2842 -4925 -2784 -4891
rect -2750 -4925 -2692 -4891
rect -2658 -4925 -2600 -4891
rect -2566 -4925 -2508 -4891
rect -2474 -4925 -2416 -4891
rect -2382 -4925 -2324 -4891
rect -2290 -4925 -2232 -4891
rect -2198 -4925 -2140 -4891
rect -2106 -4925 -2048 -4891
rect -2014 -4925 -1956 -4891
rect -1922 -4925 -1864 -4891
rect -1830 -4925 -1772 -4891
rect -1738 -4925 -1680 -4891
rect -1646 -4925 -1588 -4891
rect -1554 -4925 -1496 -4891
rect -1462 -4925 -1404 -4891
rect -1370 -4925 -1312 -4891
rect -1278 -4925 -1220 -4891
rect -1186 -4925 -1128 -4891
rect -1094 -4925 -1036 -4891
rect -1002 -4925 -944 -4891
rect -910 -4925 -852 -4891
rect -818 -4925 -760 -4891
rect -726 -4925 -668 -4891
rect -634 -4925 -576 -4891
rect -542 -4925 -484 -4891
rect -450 -4925 -392 -4891
rect -358 -4925 -300 -4891
rect -266 -4925 -208 -4891
rect -174 -4925 -116 -4891
rect -82 -4925 -24 -4891
rect 10 -4925 68 -4891
rect 102 -4925 160 -4891
rect 194 -4925 252 -4891
rect 286 -4925 344 -4891
rect 378 -4925 436 -4891
rect 470 -4925 528 -4891
rect 562 -4925 620 -4891
rect 654 -4925 712 -4891
rect 746 -4925 804 -4891
rect 838 -4925 896 -4891
rect 930 -4925 988 -4891
rect 1022 -4925 1080 -4891
rect 1114 -4925 1172 -4891
rect 1206 -4925 1264 -4891
rect 1298 -4925 1356 -4891
rect 1390 -4925 1448 -4891
rect 1482 -4925 1540 -4891
rect 1574 -4925 1632 -4891
rect 1666 -4925 1724 -4891
rect 1758 -4925 1816 -4891
rect 1850 -4925 1908 -4891
rect 1942 -4925 2000 -4891
rect 2034 -4925 2092 -4891
rect 2126 -4925 2184 -4891
rect 2218 -4925 2276 -4891
rect 2310 -4925 2368 -4891
rect 2402 -4925 2460 -4891
rect 2494 -4925 2552 -4891
rect 2586 -4925 2644 -4891
rect 2678 -4925 2736 -4891
rect 2770 -4925 2828 -4891
rect 2862 -4925 2920 -4891
rect 2954 -4925 3012 -4891
rect 3046 -4925 3104 -4891
rect 3138 -4925 3196 -4891
rect 3230 -4925 3288 -4891
rect 3322 -4925 3380 -4891
rect 3414 -4925 3472 -4891
rect 3506 -4925 3564 -4891
rect 3598 -4925 3656 -4891
rect 3690 -4925 3748 -4891
rect 3782 -4925 3840 -4891
rect 3874 -4925 3932 -4891
rect 3966 -4925 4024 -4891
rect 4058 -4925 4116 -4891
rect 4150 -4925 4208 -4891
rect 4242 -4925 4300 -4891
rect 4334 -4925 4392 -4891
rect 4426 -4925 4484 -4891
rect 4518 -4925 4576 -4891
rect 4610 -4925 4668 -4891
rect 4702 -4925 4760 -4891
rect 4794 -4925 4852 -4891
rect 4886 -4925 4944 -4891
rect 4978 -4925 5036 -4891
rect 5070 -4925 5128 -4891
rect 5162 -4925 5220 -4891
rect 5254 -4925 5312 -4891
rect 5346 -4925 5404 -4891
rect 5438 -4925 5496 -4891
rect 5530 -4925 5588 -4891
rect 5622 -4925 5680 -4891
rect 5714 -4925 5772 -4891
rect 5806 -4925 5864 -4891
rect 5898 -4925 5956 -4891
rect 5990 -4925 6048 -4891
rect 6082 -4925 6140 -4891
rect 6174 -4925 6232 -4891
rect 6266 -4925 6324 -4891
rect 6358 -4925 6416 -4891
rect 6450 -4925 6508 -4891
rect 6542 -4925 6600 -4891
rect 6634 -4925 6692 -4891
rect 6726 -4925 6784 -4891
rect 6818 -4925 6876 -4891
rect 6910 -4925 6968 -4891
rect 7002 -4925 7060 -4891
rect 7094 -4925 7152 -4891
rect 7186 -4925 7244 -4891
rect 7278 -4925 7336 -4891
rect 7370 -4925 7428 -4891
rect 7462 -4925 7520 -4891
rect 7554 -4925 7612 -4891
rect 7646 -4925 7704 -4891
rect 7738 -4925 7796 -4891
rect 7830 -4925 7888 -4891
rect 7922 -4925 7980 -4891
rect 8014 -4925 8072 -4891
rect 8106 -4925 8164 -4891
rect 8198 -4925 8256 -4891
rect 8290 -4925 8348 -4891
rect 8382 -4925 8440 -4891
rect 8474 -4925 8532 -4891
rect 8566 -4925 8624 -4891
rect 8658 -4925 8716 -4891
rect 8750 -4925 8808 -4891
rect 8842 -4925 8900 -4891
rect 8934 -4925 8992 -4891
rect 9026 -4925 9084 -4891
rect 9118 -4925 9176 -4891
rect 9210 -4925 9268 -4891
rect 9302 -4925 9360 -4891
rect 9394 -4925 9452 -4891
rect 9486 -4925 9544 -4891
rect 9578 -4925 9636 -4891
rect 9670 -4925 9728 -4891
rect 9762 -4925 9820 -4891
rect 9854 -4925 9912 -4891
rect 9946 -4925 10004 -4891
rect 10038 -4925 10096 -4891
rect 10130 -4925 10188 -4891
rect 10222 -4925 10280 -4891
rect 10314 -4925 10372 -4891
rect 10406 -4925 10464 -4891
rect 10498 -4925 10556 -4891
rect 10590 -4925 10648 -4891
rect 10682 -4925 10740 -4891
rect 10774 -4925 10832 -4891
rect 10866 -4925 10924 -4891
rect 10958 -4925 11016 -4891
rect 11050 -4925 11108 -4891
rect 11142 -4925 11200 -4891
rect 11234 -4925 11292 -4891
rect 11326 -4925 11384 -4891
rect 11418 -4925 11476 -4891
rect 11510 -4925 11568 -4891
rect 11602 -4925 11660 -4891
rect 11694 -4925 11752 -4891
rect 11786 -4925 11844 -4891
rect 11878 -4925 11936 -4891
rect 11970 -4925 12028 -4891
rect 12062 -4925 12120 -4891
rect 12154 -4925 12212 -4891
rect 12246 -4925 12304 -4891
rect 12338 -4925 12396 -4891
rect 12430 -4925 12488 -4891
rect 12522 -4925 12580 -4891
rect 12614 -4925 12672 -4891
rect 12706 -4925 12764 -4891
rect 12798 -4925 12856 -4891
rect 12890 -4925 12948 -4891
rect 12982 -4925 13040 -4891
rect 13074 -4925 13132 -4891
rect 13166 -4925 13224 -4891
rect 13258 -4925 13316 -4891
rect 13350 -4925 13408 -4891
rect 13442 -4925 13500 -4891
rect 13534 -4925 13592 -4891
rect 13626 -4925 13684 -4891
rect 13718 -4925 13776 -4891
rect 13810 -4925 13868 -4891
rect 13902 -4925 13960 -4891
rect 13994 -4925 14052 -4891
rect 14086 -4925 14144 -4891
rect 14178 -4925 14236 -4891
rect 14270 -4925 14328 -4891
rect 14362 -4925 14420 -4891
rect 14454 -4925 14512 -4891
rect 14546 -4925 14604 -4891
rect 14638 -4925 14696 -4891
rect 14730 -4925 14788 -4891
rect 14822 -4925 14880 -4891
rect 14914 -4925 14972 -4891
rect 15006 -4925 15064 -4891
rect 15098 -4925 15156 -4891
rect 15190 -4925 15248 -4891
rect 15282 -4925 15340 -4891
rect 15374 -4925 15432 -4891
rect 15466 -4925 15524 -4891
rect 15558 -4925 15616 -4891
rect 15650 -4925 15708 -4891
rect 15742 -4925 15800 -4891
rect 15834 -4925 15892 -4891
rect 15926 -4925 15984 -4891
rect 16018 -4925 16076 -4891
rect 16110 -4925 16168 -4891
rect 16202 -4925 16260 -4891
rect 16294 -4925 16352 -4891
rect 16386 -4925 16444 -4891
rect 16478 -4925 16536 -4891
rect 16570 -4925 16628 -4891
rect 16662 -4925 16691 -4891
rect -2980 -4986 -2278 -4925
rect -2980 -5020 -2962 -4986
rect -2928 -5020 -2330 -4986
rect -2296 -5020 -2278 -4986
rect -2980 -5079 -2278 -5020
rect -2244 -5019 -2186 -4925
rect -2244 -5053 -2232 -5019
rect -2198 -5053 -2186 -5019
rect -2244 -5070 -2186 -5053
rect -1600 -4986 -898 -4925
rect -1600 -5020 -1582 -4986
rect -1548 -5020 -950 -4986
rect -916 -5020 -898 -4986
rect -2980 -5147 -2902 -5113
rect -2868 -5147 -2799 -5113
rect -2765 -5147 -2696 -5113
rect -2662 -5147 -2642 -5113
rect -2980 -5217 -2642 -5147
rect -2608 -5149 -2278 -5079
rect -2608 -5183 -2588 -5149
rect -2554 -5183 -2489 -5149
rect -2455 -5183 -2390 -5149
rect -2356 -5183 -2278 -5149
rect -1600 -5079 -898 -5020
rect -864 -4986 -162 -4925
rect -864 -5020 -846 -4986
rect -812 -5020 -214 -4986
rect -180 -5020 -162 -4986
rect -864 -5079 -162 -5020
rect -128 -5019 -70 -4925
rect -128 -5053 -116 -5019
rect -82 -5053 -70 -5019
rect -128 -5070 -70 -5053
rect -36 -4993 298 -4925
rect -36 -5027 -18 -4993
rect 16 -5027 246 -4993
rect 280 -5027 298 -4993
rect -36 -5079 298 -5027
rect 332 -5019 390 -4925
rect 332 -5053 344 -5019
rect 378 -5053 390 -5019
rect 332 -5070 390 -5053
rect 424 -4978 490 -4959
rect 424 -5012 443 -4978
rect 477 -5012 490 -4978
rect 424 -5055 490 -5012
rect 524 -4978 590 -4925
rect 524 -5012 540 -4978
rect 574 -5012 590 -4978
rect 524 -5021 590 -5012
rect 683 -4978 753 -4959
rect 683 -5012 700 -4978
rect 734 -5012 753 -4978
rect -1600 -5149 -1270 -5079
rect -1600 -5183 -1522 -5149
rect -1488 -5183 -1423 -5149
rect -1389 -5183 -1324 -5149
rect -1290 -5183 -1270 -5149
rect -1236 -5147 -1216 -5113
rect -1182 -5147 -1113 -5113
rect -1079 -5147 -1010 -5113
rect -976 -5147 -898 -5113
rect -2980 -5257 -2278 -5217
rect -2980 -5291 -2962 -5257
rect -2928 -5291 -2330 -5257
rect -2296 -5291 -2278 -5257
rect -2980 -5359 -2278 -5291
rect -2980 -5393 -2962 -5359
rect -2928 -5393 -2330 -5359
rect -2296 -5393 -2278 -5359
rect -2980 -5435 -2278 -5393
rect -2244 -5237 -2186 -5202
rect -1236 -5217 -898 -5147
rect -864 -5149 -534 -5079
rect -864 -5183 -786 -5149
rect -752 -5183 -687 -5149
rect -653 -5183 -588 -5149
rect -554 -5183 -534 -5149
rect -500 -5147 -480 -5113
rect -446 -5147 -377 -5113
rect -343 -5147 -274 -5113
rect -240 -5147 -162 -5113
rect -500 -5217 -162 -5147
rect -36 -5147 -16 -5113
rect 18 -5147 114 -5113
rect -2244 -5271 -2232 -5237
rect -2198 -5271 -2186 -5237
rect -2244 -5330 -2186 -5271
rect -2244 -5364 -2232 -5330
rect -2198 -5364 -2186 -5330
rect -2244 -5435 -2186 -5364
rect -1600 -5257 -898 -5217
rect -1600 -5291 -1582 -5257
rect -1548 -5291 -950 -5257
rect -916 -5291 -898 -5257
rect -1600 -5359 -898 -5291
rect -1600 -5393 -1582 -5359
rect -1548 -5393 -950 -5359
rect -916 -5393 -898 -5359
rect -1600 -5435 -898 -5393
rect -864 -5257 -162 -5217
rect -864 -5291 -846 -5257
rect -812 -5291 -214 -5257
rect -180 -5291 -162 -5257
rect -864 -5359 -162 -5291
rect -864 -5393 -846 -5359
rect -812 -5393 -214 -5359
rect -180 -5393 -162 -5359
rect -864 -5435 -162 -5393
rect -128 -5237 -70 -5202
rect -128 -5271 -116 -5237
rect -82 -5271 -70 -5237
rect -128 -5330 -70 -5271
rect -128 -5364 -116 -5330
rect -82 -5364 -70 -5330
rect -128 -5435 -70 -5364
rect -36 -5217 114 -5147
rect 148 -5149 298 -5079
rect 424 -5089 618 -5055
rect 548 -5113 618 -5089
rect 548 -5123 634 -5113
rect 148 -5183 244 -5149
rect 278 -5183 298 -5149
rect 424 -5128 464 -5123
rect 424 -5162 436 -5128
rect 498 -5157 514 -5123
rect 470 -5162 514 -5157
rect 424 -5166 514 -5162
rect 548 -5157 584 -5123
rect 618 -5157 634 -5123
rect 548 -5171 634 -5157
rect 683 -5122 753 -5012
rect 805 -4978 855 -4959
rect 839 -5012 855 -4978
rect 805 -5054 855 -5012
rect 945 -4978 1011 -4925
rect 945 -5012 961 -4978
rect 995 -5012 1011 -4978
rect 945 -5028 1011 -5012
rect 1045 -4978 1126 -4959
rect 1045 -5012 1059 -4978
rect 1093 -5012 1126 -4978
rect 1045 -5036 1126 -5012
rect 805 -5088 923 -5054
rect 889 -5107 923 -5088
rect 683 -5123 855 -5122
rect 683 -5157 805 -5123
rect 839 -5157 855 -5123
rect 548 -5200 618 -5171
rect -36 -5257 298 -5217
rect -36 -5291 -18 -5257
rect 16 -5291 246 -5257
rect 280 -5291 298 -5257
rect -36 -5359 298 -5291
rect -36 -5393 -18 -5359
rect 16 -5393 246 -5359
rect 280 -5393 298 -5359
rect -36 -5435 298 -5393
rect 332 -5237 390 -5202
rect 332 -5271 344 -5237
rect 378 -5271 390 -5237
rect 332 -5330 390 -5271
rect 332 -5364 344 -5330
rect 378 -5364 390 -5330
rect 332 -5435 390 -5364
rect 424 -5234 618 -5200
rect 683 -5172 855 -5157
rect 889 -5123 1042 -5107
rect 889 -5157 1005 -5123
rect 1039 -5157 1042 -5123
rect 424 -5284 493 -5234
rect 424 -5318 443 -5284
rect 477 -5318 493 -5284
rect 424 -5352 493 -5318
rect 424 -5386 443 -5352
rect 477 -5386 493 -5352
rect 424 -5401 493 -5386
rect 527 -5284 593 -5268
rect 527 -5318 543 -5284
rect 577 -5318 593 -5284
rect 527 -5352 593 -5318
rect 527 -5386 543 -5352
rect 577 -5386 593 -5352
rect 527 -5435 593 -5386
rect 683 -5284 753 -5172
rect 889 -5173 1042 -5157
rect 1076 -5129 1126 -5036
rect 1160 -5019 1218 -4925
rect 1160 -5053 1172 -5019
rect 1206 -5053 1218 -5019
rect 1160 -5070 1218 -5053
rect 1252 -4993 1586 -4925
rect 1252 -5027 1270 -4993
rect 1304 -5027 1534 -4993
rect 1568 -5027 1586 -4993
rect 1252 -5079 1586 -5027
rect 1620 -5019 1678 -4925
rect 1620 -5053 1632 -5019
rect 1666 -5053 1678 -5019
rect 1620 -5070 1678 -5053
rect 1712 -4986 2414 -4925
rect 1712 -5020 1730 -4986
rect 1764 -5020 2362 -4986
rect 2396 -5020 2414 -4986
rect 1712 -5079 2414 -5020
rect 2448 -5019 2506 -4925
rect 2448 -5053 2460 -5019
rect 2494 -5053 2506 -5019
rect 2448 -5070 2506 -5053
rect 2540 -4993 2874 -4925
rect 2540 -5027 2558 -4993
rect 2592 -5027 2822 -4993
rect 2856 -5027 2874 -4993
rect 2540 -5079 2874 -5027
rect 2908 -5019 2966 -4925
rect 2908 -5053 2920 -5019
rect 2954 -5053 2966 -5019
rect 2908 -5070 2966 -5053
rect 3000 -4978 3066 -4959
rect 3000 -5012 3019 -4978
rect 3053 -5012 3066 -4978
rect 3000 -5055 3066 -5012
rect 3100 -4978 3166 -4925
rect 3100 -5012 3116 -4978
rect 3150 -5012 3166 -4978
rect 3100 -5021 3166 -5012
rect 3259 -4978 3329 -4959
rect 3259 -5012 3276 -4978
rect 3310 -5012 3329 -4978
rect 1076 -5163 1082 -5129
rect 1116 -5163 1126 -5129
rect 889 -5207 923 -5173
rect 683 -5318 701 -5284
rect 735 -5318 753 -5284
rect 683 -5352 753 -5318
rect 683 -5386 701 -5352
rect 735 -5386 753 -5352
rect 683 -5401 753 -5386
rect 805 -5241 923 -5207
rect 805 -5283 855 -5241
rect 1076 -5246 1126 -5163
rect 1252 -5147 1272 -5113
rect 1306 -5147 1402 -5113
rect 839 -5317 855 -5283
rect 805 -5351 855 -5317
rect 839 -5385 855 -5351
rect 805 -5401 855 -5385
rect 945 -5284 1011 -5275
rect 945 -5318 961 -5284
rect 995 -5318 1011 -5284
rect 945 -5352 1011 -5318
rect 945 -5386 961 -5352
rect 995 -5386 1011 -5352
rect 945 -5435 1011 -5386
rect 1045 -5283 1126 -5246
rect 1045 -5317 1059 -5283
rect 1093 -5317 1126 -5283
rect 1045 -5351 1126 -5317
rect 1045 -5385 1059 -5351
rect 1093 -5385 1126 -5351
rect 1045 -5401 1126 -5385
rect 1160 -5237 1218 -5202
rect 1160 -5271 1172 -5237
rect 1206 -5271 1218 -5237
rect 1160 -5330 1218 -5271
rect 1160 -5364 1172 -5330
rect 1206 -5364 1218 -5330
rect 1160 -5435 1218 -5364
rect 1252 -5217 1402 -5147
rect 1436 -5149 1586 -5079
rect 1436 -5183 1532 -5149
rect 1566 -5183 1586 -5149
rect 1712 -5147 1790 -5113
rect 1824 -5147 1893 -5113
rect 1927 -5147 1996 -5113
rect 2030 -5147 2050 -5113
rect 1252 -5257 1586 -5217
rect 1252 -5291 1270 -5257
rect 1304 -5291 1534 -5257
rect 1568 -5291 1586 -5257
rect 1252 -5359 1586 -5291
rect 1252 -5393 1270 -5359
rect 1304 -5393 1534 -5359
rect 1568 -5393 1586 -5359
rect 1252 -5435 1586 -5393
rect 1620 -5237 1678 -5202
rect 1620 -5271 1632 -5237
rect 1666 -5271 1678 -5237
rect 1620 -5330 1678 -5271
rect 1620 -5364 1632 -5330
rect 1666 -5364 1678 -5330
rect 1620 -5435 1678 -5364
rect 1712 -5217 2050 -5147
rect 2084 -5149 2414 -5079
rect 2084 -5183 2104 -5149
rect 2138 -5183 2203 -5149
rect 2237 -5183 2302 -5149
rect 2336 -5183 2414 -5149
rect 2540 -5147 2560 -5113
rect 2594 -5147 2690 -5113
rect 1712 -5257 2414 -5217
rect 1712 -5291 1730 -5257
rect 1764 -5291 2362 -5257
rect 2396 -5291 2414 -5257
rect 1712 -5359 2414 -5291
rect 1712 -5393 1730 -5359
rect 1764 -5393 2362 -5359
rect 2396 -5393 2414 -5359
rect 1712 -5435 2414 -5393
rect 2448 -5237 2506 -5202
rect 2448 -5271 2460 -5237
rect 2494 -5271 2506 -5237
rect 2448 -5330 2506 -5271
rect 2448 -5364 2460 -5330
rect 2494 -5364 2506 -5330
rect 2448 -5435 2506 -5364
rect 2540 -5217 2690 -5147
rect 2724 -5149 2874 -5079
rect 3000 -5089 3194 -5055
rect 3124 -5113 3194 -5089
rect 3124 -5123 3210 -5113
rect 2724 -5183 2820 -5149
rect 2854 -5183 2874 -5149
rect 3000 -5157 3040 -5123
rect 3074 -5129 3090 -5123
rect 3000 -5163 3042 -5157
rect 3076 -5163 3090 -5129
rect 3000 -5166 3090 -5163
rect 3124 -5157 3160 -5123
rect 3194 -5157 3210 -5123
rect 3124 -5171 3210 -5157
rect 3259 -5122 3329 -5012
rect 3381 -4978 3431 -4959
rect 3415 -5012 3431 -4978
rect 3381 -5054 3431 -5012
rect 3521 -4978 3587 -4925
rect 3521 -5012 3537 -4978
rect 3571 -5012 3587 -4978
rect 3521 -5028 3587 -5012
rect 3621 -4978 3702 -4959
rect 3621 -5012 3635 -4978
rect 3669 -5012 3702 -4978
rect 3621 -5036 3702 -5012
rect 3381 -5088 3499 -5054
rect 3465 -5107 3499 -5088
rect 3259 -5123 3431 -5122
rect 3259 -5157 3381 -5123
rect 3415 -5157 3431 -5123
rect 3124 -5200 3194 -5171
rect 2540 -5257 2874 -5217
rect 2540 -5291 2558 -5257
rect 2592 -5291 2822 -5257
rect 2856 -5291 2874 -5257
rect 2540 -5359 2874 -5291
rect 2540 -5393 2558 -5359
rect 2592 -5393 2822 -5359
rect 2856 -5393 2874 -5359
rect 2540 -5435 2874 -5393
rect 2908 -5237 2966 -5202
rect 2908 -5271 2920 -5237
rect 2954 -5271 2966 -5237
rect 2908 -5330 2966 -5271
rect 2908 -5364 2920 -5330
rect 2954 -5364 2966 -5330
rect 2908 -5435 2966 -5364
rect 3000 -5234 3194 -5200
rect 3259 -5172 3431 -5157
rect 3465 -5123 3618 -5107
rect 3465 -5157 3581 -5123
rect 3615 -5157 3618 -5123
rect 3000 -5284 3069 -5234
rect 3000 -5318 3019 -5284
rect 3053 -5318 3069 -5284
rect 3000 -5352 3069 -5318
rect 3000 -5386 3019 -5352
rect 3053 -5386 3069 -5352
rect 3000 -5401 3069 -5386
rect 3103 -5284 3169 -5268
rect 3103 -5318 3119 -5284
rect 3153 -5318 3169 -5284
rect 3103 -5352 3169 -5318
rect 3103 -5386 3119 -5352
rect 3153 -5386 3169 -5352
rect 3103 -5435 3169 -5386
rect 3259 -5284 3329 -5172
rect 3465 -5173 3618 -5157
rect 3652 -5129 3702 -5036
rect 3736 -5019 3794 -4925
rect 3736 -5053 3748 -5019
rect 3782 -5053 3794 -5019
rect 3736 -5070 3794 -5053
rect 3828 -4993 4162 -4925
rect 3828 -5027 3846 -4993
rect 3880 -5027 4110 -4993
rect 4144 -5027 4162 -4993
rect 3828 -5079 4162 -5027
rect 4196 -5019 4254 -4925
rect 4196 -5053 4208 -5019
rect 4242 -5053 4254 -5019
rect 4196 -5070 4254 -5053
rect 4288 -4986 4990 -4925
rect 4288 -5020 4306 -4986
rect 4340 -5020 4938 -4986
rect 4972 -5020 4990 -4986
rect 4288 -5079 4990 -5020
rect 5024 -5019 5082 -4925
rect 5024 -5053 5036 -5019
rect 5070 -5053 5082 -5019
rect 5024 -5070 5082 -5053
rect 5116 -4993 5450 -4925
rect 5116 -5027 5134 -4993
rect 5168 -5027 5398 -4993
rect 5432 -5027 5450 -4993
rect 5116 -5079 5450 -5027
rect 5484 -5019 5542 -4925
rect 5484 -5053 5496 -5019
rect 5530 -5053 5542 -5019
rect 5484 -5070 5542 -5053
rect 5576 -4978 5642 -4959
rect 5576 -5012 5595 -4978
rect 5629 -5012 5642 -4978
rect 5576 -5055 5642 -5012
rect 5676 -4978 5742 -4925
rect 5676 -5012 5692 -4978
rect 5726 -5012 5742 -4978
rect 5676 -5021 5742 -5012
rect 5835 -4978 5905 -4959
rect 5835 -5012 5852 -4978
rect 5886 -5012 5905 -4978
rect 3652 -5163 3656 -5129
rect 3690 -5163 3702 -5129
rect 3465 -5207 3499 -5173
rect 3259 -5318 3277 -5284
rect 3311 -5318 3329 -5284
rect 3259 -5352 3329 -5318
rect 3259 -5386 3277 -5352
rect 3311 -5386 3329 -5352
rect 3259 -5401 3329 -5386
rect 3381 -5241 3499 -5207
rect 3381 -5283 3431 -5241
rect 3652 -5246 3702 -5163
rect 3828 -5147 3848 -5113
rect 3882 -5147 3978 -5113
rect 3415 -5317 3431 -5283
rect 3381 -5351 3431 -5317
rect 3415 -5385 3431 -5351
rect 3381 -5401 3431 -5385
rect 3521 -5284 3587 -5275
rect 3521 -5318 3537 -5284
rect 3571 -5318 3587 -5284
rect 3521 -5352 3587 -5318
rect 3521 -5386 3537 -5352
rect 3571 -5386 3587 -5352
rect 3521 -5435 3587 -5386
rect 3621 -5283 3702 -5246
rect 3621 -5317 3635 -5283
rect 3669 -5317 3702 -5283
rect 3621 -5351 3702 -5317
rect 3621 -5385 3635 -5351
rect 3669 -5385 3702 -5351
rect 3621 -5401 3702 -5385
rect 3736 -5237 3794 -5202
rect 3736 -5271 3748 -5237
rect 3782 -5271 3794 -5237
rect 3736 -5330 3794 -5271
rect 3736 -5364 3748 -5330
rect 3782 -5364 3794 -5330
rect 3736 -5435 3794 -5364
rect 3828 -5217 3978 -5147
rect 4012 -5149 4162 -5079
rect 4012 -5183 4108 -5149
rect 4142 -5183 4162 -5149
rect 4288 -5147 4366 -5113
rect 4400 -5147 4469 -5113
rect 4503 -5147 4572 -5113
rect 4606 -5147 4626 -5113
rect 3828 -5257 4162 -5217
rect 3828 -5291 3846 -5257
rect 3880 -5291 4110 -5257
rect 4144 -5291 4162 -5257
rect 3828 -5359 4162 -5291
rect 3828 -5393 3846 -5359
rect 3880 -5393 4110 -5359
rect 4144 -5393 4162 -5359
rect 3828 -5435 4162 -5393
rect 4196 -5237 4254 -5202
rect 4196 -5271 4208 -5237
rect 4242 -5271 4254 -5237
rect 4196 -5330 4254 -5271
rect 4196 -5364 4208 -5330
rect 4242 -5364 4254 -5330
rect 4196 -5435 4254 -5364
rect 4288 -5217 4626 -5147
rect 4660 -5149 4990 -5079
rect 4660 -5183 4680 -5149
rect 4714 -5183 4779 -5149
rect 4813 -5183 4878 -5149
rect 4912 -5183 4990 -5149
rect 5116 -5147 5136 -5113
rect 5170 -5147 5266 -5113
rect 4288 -5257 4990 -5217
rect 4288 -5291 4306 -5257
rect 4340 -5291 4938 -5257
rect 4972 -5291 4990 -5257
rect 4288 -5359 4990 -5291
rect 4288 -5393 4306 -5359
rect 4340 -5393 4938 -5359
rect 4972 -5393 4990 -5359
rect 4288 -5435 4990 -5393
rect 5024 -5237 5082 -5202
rect 5024 -5271 5036 -5237
rect 5070 -5271 5082 -5237
rect 5024 -5330 5082 -5271
rect 5024 -5364 5036 -5330
rect 5070 -5364 5082 -5330
rect 5024 -5435 5082 -5364
rect 5116 -5217 5266 -5147
rect 5300 -5149 5450 -5079
rect 5576 -5089 5770 -5055
rect 5700 -5113 5770 -5089
rect 5700 -5123 5786 -5113
rect 5300 -5183 5396 -5149
rect 5430 -5183 5450 -5149
rect 5576 -5163 5616 -5123
rect 5650 -5163 5666 -5123
rect 5576 -5166 5666 -5163
rect 5700 -5157 5736 -5123
rect 5770 -5157 5786 -5123
rect 5700 -5171 5786 -5157
rect 5835 -5122 5905 -5012
rect 5957 -4978 6007 -4959
rect 5991 -5012 6007 -4978
rect 5957 -5054 6007 -5012
rect 6097 -4978 6163 -4925
rect 6097 -5012 6113 -4978
rect 6147 -5012 6163 -4978
rect 6097 -5028 6163 -5012
rect 6197 -4978 6278 -4959
rect 6197 -5012 6211 -4978
rect 6245 -5012 6278 -4978
rect 6197 -5036 6278 -5012
rect 5957 -5088 6075 -5054
rect 6041 -5107 6075 -5088
rect 5835 -5123 6007 -5122
rect 5835 -5157 5957 -5123
rect 5991 -5157 6007 -5123
rect 5700 -5200 5770 -5171
rect 5116 -5257 5450 -5217
rect 5116 -5291 5134 -5257
rect 5168 -5291 5398 -5257
rect 5432 -5291 5450 -5257
rect 5116 -5359 5450 -5291
rect 5116 -5393 5134 -5359
rect 5168 -5393 5398 -5359
rect 5432 -5393 5450 -5359
rect 5116 -5435 5450 -5393
rect 5484 -5237 5542 -5202
rect 5484 -5271 5496 -5237
rect 5530 -5271 5542 -5237
rect 5484 -5330 5542 -5271
rect 5484 -5364 5496 -5330
rect 5530 -5364 5542 -5330
rect 5484 -5435 5542 -5364
rect 5576 -5234 5770 -5200
rect 5835 -5172 6007 -5157
rect 6041 -5123 6194 -5107
rect 6041 -5157 6157 -5123
rect 6191 -5157 6194 -5123
rect 5576 -5284 5645 -5234
rect 5576 -5318 5595 -5284
rect 5629 -5318 5645 -5284
rect 5576 -5352 5645 -5318
rect 5576 -5386 5595 -5352
rect 5629 -5386 5645 -5352
rect 5576 -5401 5645 -5386
rect 5679 -5284 5745 -5268
rect 5679 -5318 5695 -5284
rect 5729 -5318 5745 -5284
rect 5679 -5352 5745 -5318
rect 5679 -5386 5695 -5352
rect 5729 -5386 5745 -5352
rect 5679 -5435 5745 -5386
rect 5835 -5284 5905 -5172
rect 6041 -5173 6194 -5157
rect 6228 -5129 6278 -5036
rect 6312 -5019 6370 -4925
rect 6312 -5053 6324 -5019
rect 6358 -5053 6370 -5019
rect 6312 -5070 6370 -5053
rect 6404 -4993 6738 -4925
rect 6404 -5027 6422 -4993
rect 6456 -5027 6686 -4993
rect 6720 -5027 6738 -4993
rect 6404 -5079 6738 -5027
rect 6772 -5019 6830 -4925
rect 6772 -5053 6784 -5019
rect 6818 -5053 6830 -5019
rect 6772 -5070 6830 -5053
rect 6864 -4986 7566 -4925
rect 6864 -5020 6882 -4986
rect 6916 -5020 7514 -4986
rect 7548 -5020 7566 -4986
rect 6864 -5079 7566 -5020
rect 7600 -5019 7658 -4925
rect 7600 -5053 7612 -5019
rect 7646 -5053 7658 -5019
rect 7600 -5070 7658 -5053
rect 7692 -4993 8026 -4925
rect 7692 -5027 7710 -4993
rect 7744 -5027 7974 -4993
rect 8008 -5027 8026 -4993
rect 7692 -5079 8026 -5027
rect 8060 -5019 8118 -4925
rect 8060 -5053 8072 -5019
rect 8106 -5053 8118 -5019
rect 8060 -5070 8118 -5053
rect 8152 -4978 8218 -4959
rect 8152 -5012 8171 -4978
rect 8205 -5012 8218 -4978
rect 8152 -5055 8218 -5012
rect 8252 -4978 8318 -4925
rect 8252 -5012 8268 -4978
rect 8302 -5012 8318 -4978
rect 8252 -5021 8318 -5012
rect 8411 -4978 8481 -4959
rect 8411 -5012 8428 -4978
rect 8462 -5012 8481 -4978
rect 6228 -5163 6230 -5129
rect 6264 -5163 6278 -5129
rect 6041 -5207 6075 -5173
rect 5835 -5318 5853 -5284
rect 5887 -5318 5905 -5284
rect 5835 -5352 5905 -5318
rect 5835 -5386 5853 -5352
rect 5887 -5386 5905 -5352
rect 5835 -5401 5905 -5386
rect 5957 -5241 6075 -5207
rect 5957 -5283 6007 -5241
rect 6228 -5246 6278 -5163
rect 6404 -5147 6424 -5113
rect 6458 -5147 6554 -5113
rect 5991 -5317 6007 -5283
rect 5957 -5351 6007 -5317
rect 5991 -5385 6007 -5351
rect 5957 -5401 6007 -5385
rect 6097 -5284 6163 -5275
rect 6097 -5318 6113 -5284
rect 6147 -5318 6163 -5284
rect 6097 -5352 6163 -5318
rect 6097 -5386 6113 -5352
rect 6147 -5386 6163 -5352
rect 6097 -5435 6163 -5386
rect 6197 -5283 6278 -5246
rect 6197 -5317 6211 -5283
rect 6245 -5317 6278 -5283
rect 6197 -5351 6278 -5317
rect 6197 -5385 6211 -5351
rect 6245 -5385 6278 -5351
rect 6197 -5401 6278 -5385
rect 6312 -5237 6370 -5202
rect 6312 -5271 6324 -5237
rect 6358 -5271 6370 -5237
rect 6312 -5330 6370 -5271
rect 6312 -5364 6324 -5330
rect 6358 -5364 6370 -5330
rect 6312 -5435 6370 -5364
rect 6404 -5217 6554 -5147
rect 6588 -5149 6738 -5079
rect 6588 -5183 6684 -5149
rect 6718 -5183 6738 -5149
rect 6864 -5147 6942 -5113
rect 6976 -5147 7045 -5113
rect 7079 -5147 7148 -5113
rect 7182 -5147 7202 -5113
rect 6404 -5257 6738 -5217
rect 6404 -5291 6422 -5257
rect 6456 -5291 6686 -5257
rect 6720 -5291 6738 -5257
rect 6404 -5359 6738 -5291
rect 6404 -5393 6422 -5359
rect 6456 -5393 6686 -5359
rect 6720 -5393 6738 -5359
rect 6404 -5435 6738 -5393
rect 6772 -5237 6830 -5202
rect 6772 -5271 6784 -5237
rect 6818 -5271 6830 -5237
rect 6772 -5330 6830 -5271
rect 6772 -5364 6784 -5330
rect 6818 -5364 6830 -5330
rect 6772 -5435 6830 -5364
rect 6864 -5217 7202 -5147
rect 7236 -5149 7566 -5079
rect 7236 -5183 7256 -5149
rect 7290 -5183 7355 -5149
rect 7389 -5183 7454 -5149
rect 7488 -5183 7566 -5149
rect 7692 -5147 7712 -5113
rect 7746 -5147 7842 -5113
rect 6864 -5257 7566 -5217
rect 6864 -5291 6882 -5257
rect 6916 -5291 7514 -5257
rect 7548 -5291 7566 -5257
rect 6864 -5359 7566 -5291
rect 6864 -5393 6882 -5359
rect 6916 -5393 7514 -5359
rect 7548 -5393 7566 -5359
rect 6864 -5435 7566 -5393
rect 7600 -5237 7658 -5202
rect 7600 -5271 7612 -5237
rect 7646 -5271 7658 -5237
rect 7600 -5330 7658 -5271
rect 7600 -5364 7612 -5330
rect 7646 -5364 7658 -5330
rect 7600 -5435 7658 -5364
rect 7692 -5217 7842 -5147
rect 7876 -5149 8026 -5079
rect 8152 -5089 8346 -5055
rect 8276 -5113 8346 -5089
rect 8276 -5123 8362 -5113
rect 7876 -5183 7972 -5149
rect 8006 -5183 8026 -5149
rect 8152 -5129 8192 -5123
rect 8152 -5163 8190 -5129
rect 8226 -5157 8242 -5123
rect 8224 -5163 8242 -5157
rect 8152 -5166 8242 -5163
rect 8276 -5157 8312 -5123
rect 8346 -5157 8362 -5123
rect 8276 -5171 8362 -5157
rect 8411 -5122 8481 -5012
rect 8533 -4978 8583 -4959
rect 8567 -5012 8583 -4978
rect 8533 -5054 8583 -5012
rect 8673 -4978 8739 -4925
rect 8673 -5012 8689 -4978
rect 8723 -5012 8739 -4978
rect 8673 -5028 8739 -5012
rect 8773 -4978 8854 -4959
rect 8773 -5012 8787 -4978
rect 8821 -5012 8854 -4978
rect 8773 -5036 8854 -5012
rect 8533 -5088 8651 -5054
rect 8617 -5107 8651 -5088
rect 8411 -5123 8583 -5122
rect 8411 -5157 8533 -5123
rect 8567 -5157 8583 -5123
rect 8276 -5200 8346 -5171
rect 7692 -5257 8026 -5217
rect 7692 -5291 7710 -5257
rect 7744 -5291 7974 -5257
rect 8008 -5291 8026 -5257
rect 7692 -5359 8026 -5291
rect 7692 -5393 7710 -5359
rect 7744 -5393 7974 -5359
rect 8008 -5393 8026 -5359
rect 7692 -5435 8026 -5393
rect 8060 -5237 8118 -5202
rect 8060 -5271 8072 -5237
rect 8106 -5271 8118 -5237
rect 8060 -5330 8118 -5271
rect 8060 -5364 8072 -5330
rect 8106 -5364 8118 -5330
rect 8060 -5435 8118 -5364
rect 8152 -5234 8346 -5200
rect 8411 -5172 8583 -5157
rect 8617 -5123 8770 -5107
rect 8617 -5157 8733 -5123
rect 8767 -5157 8770 -5123
rect 8152 -5284 8221 -5234
rect 8152 -5318 8171 -5284
rect 8205 -5318 8221 -5284
rect 8152 -5352 8221 -5318
rect 8152 -5386 8171 -5352
rect 8205 -5386 8221 -5352
rect 8152 -5401 8221 -5386
rect 8255 -5284 8321 -5268
rect 8255 -5318 8271 -5284
rect 8305 -5318 8321 -5284
rect 8255 -5352 8321 -5318
rect 8255 -5386 8271 -5352
rect 8305 -5386 8321 -5352
rect 8255 -5435 8321 -5386
rect 8411 -5284 8481 -5172
rect 8617 -5173 8770 -5157
rect 8804 -5129 8854 -5036
rect 8888 -5019 8946 -4925
rect 8888 -5053 8900 -5019
rect 8934 -5053 8946 -5019
rect 8888 -5070 8946 -5053
rect 8980 -4993 9314 -4925
rect 8980 -5027 8998 -4993
rect 9032 -5027 9262 -4993
rect 9296 -5027 9314 -4993
rect 8980 -5079 9314 -5027
rect 9348 -5019 9406 -4925
rect 9348 -5053 9360 -5019
rect 9394 -5053 9406 -5019
rect 9348 -5070 9406 -5053
rect 9440 -4986 10142 -4925
rect 9440 -5020 9458 -4986
rect 9492 -5020 10090 -4986
rect 10124 -5020 10142 -4986
rect 9440 -5079 10142 -5020
rect 10176 -5019 10234 -4925
rect 10176 -5053 10188 -5019
rect 10222 -5053 10234 -5019
rect 10176 -5070 10234 -5053
rect 10360 -4993 10694 -4925
rect 10360 -5027 10378 -4993
rect 10412 -5027 10642 -4993
rect 10676 -5027 10694 -4993
rect 10360 -5079 10694 -5027
rect 8838 -5163 8854 -5129
rect 8617 -5207 8651 -5173
rect 8411 -5318 8429 -5284
rect 8463 -5318 8481 -5284
rect 8411 -5352 8481 -5318
rect 8411 -5386 8429 -5352
rect 8463 -5386 8481 -5352
rect 8411 -5401 8481 -5386
rect 8533 -5241 8651 -5207
rect 8533 -5283 8583 -5241
rect 8804 -5246 8854 -5163
rect 8980 -5147 9000 -5113
rect 9034 -5147 9130 -5113
rect 8567 -5317 8583 -5283
rect 8533 -5351 8583 -5317
rect 8567 -5385 8583 -5351
rect 8533 -5401 8583 -5385
rect 8673 -5284 8739 -5275
rect 8673 -5318 8689 -5284
rect 8723 -5318 8739 -5284
rect 8673 -5352 8739 -5318
rect 8673 -5386 8689 -5352
rect 8723 -5386 8739 -5352
rect 8673 -5435 8739 -5386
rect 8773 -5283 8854 -5246
rect 8773 -5317 8787 -5283
rect 8821 -5317 8854 -5283
rect 8773 -5351 8854 -5317
rect 8773 -5385 8787 -5351
rect 8821 -5385 8854 -5351
rect 8773 -5401 8854 -5385
rect 8888 -5237 8946 -5202
rect 8888 -5271 8900 -5237
rect 8934 -5271 8946 -5237
rect 8888 -5330 8946 -5271
rect 8888 -5364 8900 -5330
rect 8934 -5364 8946 -5330
rect 8888 -5435 8946 -5364
rect 8980 -5217 9130 -5147
rect 9164 -5149 9314 -5079
rect 9164 -5183 9260 -5149
rect 9294 -5183 9314 -5149
rect 9440 -5147 9518 -5113
rect 9552 -5147 9621 -5113
rect 9655 -5147 9724 -5113
rect 9758 -5147 9778 -5113
rect 8980 -5257 9314 -5217
rect 8980 -5291 8998 -5257
rect 9032 -5291 9262 -5257
rect 9296 -5291 9314 -5257
rect 8980 -5359 9314 -5291
rect 8980 -5393 8998 -5359
rect 9032 -5393 9262 -5359
rect 9296 -5393 9314 -5359
rect 8980 -5435 9314 -5393
rect 9348 -5237 9406 -5202
rect 9348 -5271 9360 -5237
rect 9394 -5271 9406 -5237
rect 9348 -5330 9406 -5271
rect 9348 -5364 9360 -5330
rect 9394 -5364 9406 -5330
rect 9348 -5435 9406 -5364
rect 9440 -5217 9778 -5147
rect 9812 -5149 10142 -5079
rect 9812 -5183 9832 -5149
rect 9866 -5183 9931 -5149
rect 9965 -5183 10030 -5149
rect 10064 -5183 10142 -5149
rect 10360 -5147 10380 -5113
rect 10414 -5147 10510 -5113
rect 9440 -5257 10142 -5217
rect 9440 -5291 9458 -5257
rect 9492 -5291 10090 -5257
rect 10124 -5291 10142 -5257
rect 9440 -5359 10142 -5291
rect 9440 -5393 9458 -5359
rect 9492 -5393 10090 -5359
rect 10124 -5393 10142 -5359
rect 9440 -5435 10142 -5393
rect 10176 -5237 10234 -5202
rect 10176 -5271 10188 -5237
rect 10222 -5271 10234 -5237
rect 10176 -5330 10234 -5271
rect 10176 -5364 10188 -5330
rect 10222 -5364 10234 -5330
rect 10176 -5435 10234 -5364
rect 10360 -5217 10510 -5147
rect 10544 -5149 10694 -5079
rect 10728 -4978 10794 -4959
rect 10728 -5012 10747 -4978
rect 10781 -5012 10794 -4978
rect 10728 -5055 10794 -5012
rect 10828 -4978 10894 -4925
rect 10828 -5012 10844 -4978
rect 10878 -5012 10894 -4978
rect 10828 -5021 10894 -5012
rect 10987 -4978 11057 -4959
rect 10987 -5012 11004 -4978
rect 11038 -5012 11057 -4978
rect 10728 -5089 10922 -5055
rect 10852 -5113 10922 -5089
rect 10852 -5123 10938 -5113
rect 10544 -5183 10640 -5149
rect 10674 -5183 10694 -5149
rect 10728 -5129 10768 -5123
rect 10728 -5163 10764 -5129
rect 10802 -5157 10818 -5123
rect 10798 -5163 10818 -5157
rect 10728 -5166 10818 -5163
rect 10852 -5157 10888 -5123
rect 10922 -5157 10938 -5123
rect 10852 -5171 10938 -5157
rect 10987 -5122 11057 -5012
rect 11109 -4978 11159 -4959
rect 11143 -5012 11159 -4978
rect 11109 -5054 11159 -5012
rect 11249 -4978 11315 -4925
rect 11249 -5012 11265 -4978
rect 11299 -5012 11315 -4978
rect 11249 -5028 11315 -5012
rect 11349 -4978 11430 -4959
rect 11349 -5012 11363 -4978
rect 11397 -5012 11430 -4978
rect 11349 -5036 11430 -5012
rect 11109 -5088 11227 -5054
rect 11193 -5107 11227 -5088
rect 10987 -5123 11159 -5122
rect 10987 -5157 11109 -5123
rect 11143 -5157 11159 -5123
rect 10852 -5200 10922 -5171
rect 10360 -5257 10694 -5217
rect 10360 -5291 10378 -5257
rect 10412 -5291 10642 -5257
rect 10676 -5291 10694 -5257
rect 10360 -5359 10694 -5291
rect 10360 -5393 10378 -5359
rect 10412 -5393 10642 -5359
rect 10676 -5393 10694 -5359
rect 10360 -5435 10694 -5393
rect 10728 -5234 10922 -5200
rect 10987 -5172 11159 -5157
rect 11193 -5123 11346 -5107
rect 11193 -5157 11309 -5123
rect 11343 -5157 11346 -5123
rect 10728 -5284 10797 -5234
rect 10728 -5318 10747 -5284
rect 10781 -5318 10797 -5284
rect 10728 -5352 10797 -5318
rect 10728 -5386 10747 -5352
rect 10781 -5386 10797 -5352
rect 10728 -5401 10797 -5386
rect 10831 -5284 10897 -5268
rect 10831 -5318 10847 -5284
rect 10881 -5318 10897 -5284
rect 10831 -5352 10897 -5318
rect 10831 -5386 10847 -5352
rect 10881 -5386 10897 -5352
rect 10831 -5435 10897 -5386
rect 10987 -5284 11057 -5172
rect 11193 -5173 11346 -5157
rect 11380 -5162 11430 -5036
rect 11464 -5019 11522 -4925
rect 11464 -5053 11476 -5019
rect 11510 -5053 11522 -5019
rect 11464 -5070 11522 -5053
rect 11648 -4993 11982 -4925
rect 11648 -5027 11666 -4993
rect 11700 -5027 11930 -4993
rect 11964 -5027 11982 -4993
rect 11648 -5079 11982 -5027
rect 12384 -5019 12442 -4925
rect 12572 -4969 12631 -4925
rect 12572 -5003 12588 -4969
rect 12622 -5003 12631 -4969
rect 12572 -5019 12631 -5003
rect 12665 -4980 12717 -4964
rect 12665 -5014 12674 -4980
rect 12708 -5014 12717 -4980
rect 12384 -5053 12396 -5019
rect 12430 -5053 12442 -5019
rect 12665 -5053 12717 -5014
rect 12751 -4969 12803 -4925
rect 12751 -5003 12760 -4969
rect 12794 -5003 12803 -4969
rect 12751 -5019 12803 -5003
rect 12837 -4980 12888 -4964
rect 12837 -5014 12846 -4980
rect 12880 -5014 12888 -4980
rect 12837 -5053 12888 -5014
rect 12922 -4969 12982 -4925
rect 12922 -5003 12932 -4969
rect 12966 -5003 12982 -4969
rect 12922 -5019 12982 -5003
rect 13120 -5019 13178 -4925
rect 13120 -5053 13132 -5019
rect 13166 -5053 13178 -5019
rect 12384 -5070 12442 -5053
rect 12480 -5061 13086 -5053
rect 11193 -5207 11227 -5173
rect 10987 -5318 11005 -5284
rect 11039 -5318 11057 -5284
rect 10987 -5352 11057 -5318
rect 10987 -5386 11005 -5352
rect 11039 -5386 11057 -5352
rect 10987 -5401 11057 -5386
rect 11109 -5241 11227 -5207
rect 11380 -5196 11389 -5162
rect 11423 -5196 11430 -5162
rect 11109 -5283 11159 -5241
rect 11380 -5246 11430 -5196
rect 11648 -5147 11668 -5113
rect 11702 -5147 11798 -5113
rect 11143 -5317 11159 -5283
rect 11109 -5351 11159 -5317
rect 11143 -5385 11159 -5351
rect 11109 -5401 11159 -5385
rect 11249 -5284 11315 -5275
rect 11249 -5318 11265 -5284
rect 11299 -5318 11315 -5284
rect 11249 -5352 11315 -5318
rect 11249 -5386 11265 -5352
rect 11299 -5386 11315 -5352
rect 11249 -5435 11315 -5386
rect 11349 -5283 11430 -5246
rect 11349 -5317 11363 -5283
rect 11397 -5317 11430 -5283
rect 11349 -5351 11430 -5317
rect 11349 -5385 11363 -5351
rect 11397 -5385 11430 -5351
rect 11349 -5401 11430 -5385
rect 11464 -5237 11522 -5202
rect 11464 -5271 11476 -5237
rect 11510 -5271 11522 -5237
rect 11464 -5330 11522 -5271
rect 11464 -5364 11476 -5330
rect 11510 -5364 11522 -5330
rect 11464 -5435 11522 -5364
rect 11648 -5217 11798 -5147
rect 11832 -5149 11982 -5079
rect 11832 -5183 11928 -5149
rect 11962 -5183 11982 -5149
rect 12480 -5087 13038 -5061
rect 12480 -5200 12514 -5087
rect 13026 -5095 13038 -5087
rect 13072 -5095 13086 -5061
rect 13120 -5070 13178 -5053
rect 13212 -4993 13546 -4925
rect 13212 -5027 13230 -4993
rect 13264 -5027 13494 -4993
rect 13528 -5027 13546 -4993
rect 12548 -5123 12991 -5121
rect 12548 -5126 12574 -5123
rect 12548 -5160 12558 -5126
rect 12608 -5157 12642 -5123
rect 12676 -5157 12710 -5123
rect 12744 -5126 12778 -5123
rect 12773 -5157 12778 -5126
rect 12812 -5126 12846 -5123
rect 12812 -5157 12836 -5126
rect 12880 -5157 12914 -5123
rect 12948 -5126 12991 -5123
rect 12592 -5160 12642 -5157
rect 12676 -5160 12739 -5157
rect 12773 -5160 12836 -5157
rect 12870 -5160 12942 -5157
rect 12976 -5160 12991 -5126
rect 12548 -5166 12991 -5160
rect 13026 -5133 13086 -5095
rect 13026 -5167 13038 -5133
rect 13072 -5167 13086 -5133
rect 13026 -5200 13086 -5167
rect 13212 -5079 13546 -5027
rect 13580 -5019 13638 -4925
rect 13580 -5053 13592 -5019
rect 13626 -5053 13638 -5019
rect 13672 -4967 13733 -4925
rect 13672 -5001 13690 -4967
rect 13724 -5001 13733 -4967
rect 13672 -5027 13733 -5001
rect 13769 -4980 13819 -4961
rect 13769 -5014 13776 -4980
rect 13810 -5014 13819 -4980
rect 13580 -5070 13638 -5053
rect 13212 -5149 13362 -5079
rect 13672 -5096 13735 -5061
rect 13212 -5183 13232 -5149
rect 13266 -5183 13362 -5149
rect 13396 -5147 13492 -5113
rect 13526 -5147 13546 -5113
rect 11648 -5257 11982 -5217
rect 11648 -5291 11666 -5257
rect 11700 -5291 11930 -5257
rect 11964 -5291 11982 -5257
rect 11648 -5359 11982 -5291
rect 11648 -5393 11666 -5359
rect 11700 -5393 11930 -5359
rect 11964 -5393 11982 -5359
rect 11648 -5435 11982 -5393
rect 12384 -5237 12442 -5202
rect 12480 -5234 13086 -5200
rect 12384 -5271 12396 -5237
rect 12430 -5271 12442 -5237
rect 12580 -5257 12631 -5234
rect 12384 -5330 12442 -5271
rect 12384 -5364 12396 -5330
rect 12430 -5364 12442 -5330
rect 12384 -5435 12442 -5364
rect 12476 -5284 12545 -5268
rect 12476 -5318 12502 -5284
rect 12536 -5318 12545 -5284
rect 12476 -5352 12545 -5318
rect 12476 -5386 12502 -5352
rect 12536 -5386 12545 -5352
rect 12476 -5435 12545 -5386
rect 12580 -5291 12588 -5257
rect 12622 -5291 12631 -5257
rect 12752 -5257 12803 -5234
rect 12580 -5345 12631 -5291
rect 12580 -5379 12588 -5345
rect 12622 -5379 12631 -5345
rect 12580 -5395 12631 -5379
rect 12665 -5284 12717 -5268
rect 12665 -5318 12674 -5284
rect 12708 -5318 12717 -5284
rect 12665 -5352 12717 -5318
rect 12665 -5386 12674 -5352
rect 12708 -5386 12717 -5352
rect 12665 -5435 12717 -5386
rect 12752 -5291 12760 -5257
rect 12794 -5291 12803 -5257
rect 12923 -5257 12975 -5234
rect 12752 -5345 12803 -5291
rect 12752 -5379 12760 -5345
rect 12794 -5379 12803 -5345
rect 12752 -5395 12803 -5379
rect 12837 -5284 12889 -5268
rect 12837 -5318 12846 -5284
rect 12880 -5318 12889 -5284
rect 12837 -5352 12889 -5318
rect 12837 -5386 12846 -5352
rect 12880 -5386 12889 -5352
rect 12837 -5435 12889 -5386
rect 12923 -5291 12932 -5257
rect 12966 -5291 12975 -5257
rect 13120 -5237 13178 -5202
rect 13396 -5217 13546 -5147
rect 13672 -5130 13684 -5096
rect 13718 -5123 13735 -5096
rect 13672 -5157 13692 -5130
rect 13726 -5157 13735 -5123
rect 13672 -5173 13735 -5157
rect 13769 -5123 13819 -5014
rect 13853 -4980 13905 -4925
rect 13853 -5014 13862 -4980
rect 13896 -5014 13905 -4980
rect 13853 -5030 13905 -5014
rect 13941 -4980 13991 -4961
rect 13941 -5014 13948 -4980
rect 13982 -5014 13991 -4980
rect 13941 -5123 13991 -5014
rect 14025 -4980 14077 -4925
rect 14025 -5014 14034 -4980
rect 14068 -5014 14077 -4980
rect 14025 -5037 14077 -5014
rect 14111 -4980 14163 -4964
rect 14111 -5014 14120 -4980
rect 14154 -5014 14163 -4980
rect 14111 -5055 14163 -5014
rect 14197 -4971 14249 -4925
rect 14197 -5005 14206 -4971
rect 14240 -5005 14249 -4971
rect 14197 -5021 14249 -5005
rect 14283 -4980 14335 -4964
rect 14283 -5014 14292 -4980
rect 14326 -5014 14335 -4980
rect 14283 -5055 14335 -5014
rect 14369 -4971 14421 -4925
rect 14369 -5005 14378 -4971
rect 14412 -5005 14421 -4971
rect 14369 -5021 14421 -5005
rect 14455 -4980 14507 -4964
rect 14455 -5014 14464 -4980
rect 14498 -5014 14507 -4980
rect 14455 -5055 14507 -5014
rect 14541 -4971 14590 -4925
rect 14541 -5005 14550 -4971
rect 14584 -5005 14590 -4971
rect 14541 -5021 14590 -5005
rect 14624 -4980 14679 -4964
rect 14624 -5014 14636 -4980
rect 14670 -5014 14679 -4980
rect 14624 -5055 14679 -5014
rect 14713 -4971 14762 -4925
rect 14713 -5005 14722 -4971
rect 14756 -5005 14762 -4971
rect 14713 -5021 14762 -5005
rect 14796 -4980 14848 -4964
rect 14796 -5014 14807 -4980
rect 14841 -5014 14848 -4980
rect 14796 -5055 14848 -5014
rect 14884 -4971 14934 -4925
rect 14884 -5005 14893 -4971
rect 14927 -5005 14934 -4971
rect 14884 -5021 14934 -5005
rect 14968 -4980 15020 -4964
rect 14968 -5014 14979 -4980
rect 15013 -5014 15020 -4980
rect 14968 -5055 15020 -5014
rect 15056 -4971 15106 -4925
rect 15056 -5005 15065 -4971
rect 15099 -5005 15106 -4971
rect 15056 -5021 15106 -5005
rect 15140 -4980 15192 -4964
rect 15140 -5014 15151 -4980
rect 15185 -5014 15192 -4980
rect 15140 -5055 15192 -5014
rect 15228 -4971 15280 -4925
rect 15228 -5005 15237 -4971
rect 15271 -5005 15280 -4971
rect 15228 -5021 15280 -5005
rect 15314 -4980 15366 -4964
rect 15314 -5014 15323 -4980
rect 15357 -5014 15366 -4980
rect 15314 -5055 15366 -5014
rect 15400 -4971 15460 -4925
rect 15400 -5005 15409 -4971
rect 15443 -5005 15460 -4971
rect 15400 -5021 15460 -5005
rect 15512 -5019 15570 -4925
rect 15512 -5053 15524 -5019
rect 15558 -5053 15570 -5019
rect 14111 -5084 15460 -5055
rect 15512 -5070 15570 -5053
rect 15604 -4986 16673 -4925
rect 15604 -5020 15622 -4986
rect 15656 -5020 16622 -4986
rect 16656 -5020 16673 -4986
rect 14111 -5089 15248 -5084
rect 15227 -5118 15248 -5089
rect 15282 -5118 15341 -5084
rect 15375 -5118 15460 -5084
rect 13769 -5157 14119 -5123
rect 14153 -5157 14187 -5123
rect 14221 -5157 14255 -5123
rect 14289 -5157 14323 -5123
rect 14357 -5157 14391 -5123
rect 14425 -5157 14459 -5123
rect 14493 -5157 14527 -5123
rect 14561 -5157 14595 -5123
rect 14629 -5157 14663 -5123
rect 14697 -5157 14731 -5123
rect 14765 -5157 14799 -5123
rect 14833 -5157 14867 -5123
rect 14901 -5157 14935 -5123
rect 14969 -5157 15003 -5123
rect 15037 -5157 15071 -5123
rect 15105 -5157 15139 -5123
rect 15173 -5157 15193 -5123
rect 13769 -5173 15193 -5157
rect 12923 -5345 12975 -5291
rect 12923 -5379 12932 -5345
rect 12966 -5379 12975 -5345
rect 12923 -5395 12975 -5379
rect 13009 -5284 13086 -5268
rect 13009 -5318 13018 -5284
rect 13052 -5318 13086 -5284
rect 13009 -5352 13086 -5318
rect 13009 -5386 13018 -5352
rect 13052 -5386 13086 -5352
rect 13009 -5435 13086 -5386
rect 13120 -5271 13132 -5237
rect 13166 -5271 13178 -5237
rect 13120 -5330 13178 -5271
rect 13120 -5364 13132 -5330
rect 13166 -5364 13178 -5330
rect 13120 -5435 13178 -5364
rect 13212 -5257 13546 -5217
rect 13212 -5291 13230 -5257
rect 13264 -5291 13494 -5257
rect 13528 -5291 13546 -5257
rect 13212 -5359 13546 -5291
rect 13212 -5393 13230 -5359
rect 13264 -5393 13494 -5359
rect 13528 -5393 13546 -5359
rect 13212 -5435 13546 -5393
rect 13580 -5237 13638 -5202
rect 13580 -5271 13592 -5237
rect 13626 -5271 13638 -5237
rect 13580 -5330 13638 -5271
rect 13580 -5364 13592 -5330
rect 13626 -5364 13638 -5330
rect 13580 -5435 13638 -5364
rect 13674 -5291 13733 -5273
rect 13674 -5325 13690 -5291
rect 13724 -5325 13733 -5291
rect 13674 -5359 13733 -5325
rect 13674 -5393 13690 -5359
rect 13724 -5393 13733 -5359
rect 13674 -5435 13733 -5393
rect 13769 -5283 13818 -5173
rect 13769 -5317 13776 -5283
rect 13810 -5317 13818 -5283
rect 13769 -5351 13818 -5317
rect 13769 -5385 13776 -5351
rect 13810 -5385 13818 -5351
rect 13769 -5401 13818 -5385
rect 13853 -5291 13905 -5273
rect 13853 -5325 13862 -5291
rect 13896 -5325 13905 -5291
rect 13853 -5359 13905 -5325
rect 13853 -5393 13862 -5359
rect 13896 -5393 13905 -5359
rect 13853 -5435 13905 -5393
rect 13941 -5275 13991 -5173
rect 15227 -5179 15460 -5118
rect 15227 -5180 15340 -5179
rect 15227 -5207 15248 -5180
rect 14111 -5214 15248 -5207
rect 15282 -5213 15340 -5180
rect 15374 -5213 15460 -5179
rect 15604 -5079 16673 -5020
rect 15604 -5149 16120 -5079
rect 15604 -5183 15682 -5149
rect 15716 -5183 15810 -5149
rect 15844 -5183 15938 -5149
rect 15972 -5183 16066 -5149
rect 16100 -5183 16120 -5149
rect 16154 -5147 16174 -5113
rect 16208 -5147 16302 -5113
rect 16336 -5147 16430 -5113
rect 16464 -5147 16558 -5113
rect 16592 -5147 16673 -5113
rect 15282 -5214 15460 -5213
rect 14111 -5229 15460 -5214
rect 14111 -5263 14120 -5229
rect 14154 -5255 14292 -5229
rect 14154 -5263 14163 -5255
rect 13941 -5309 13948 -5275
rect 13982 -5309 13991 -5275
rect 13941 -5343 13991 -5309
rect 13941 -5377 13948 -5343
rect 13982 -5377 13991 -5343
rect 13941 -5400 13991 -5377
rect 14025 -5291 14077 -5275
rect 14025 -5325 14034 -5291
rect 14068 -5325 14077 -5291
rect 14025 -5359 14077 -5325
rect 14025 -5393 14034 -5359
rect 14068 -5393 14077 -5359
rect 14025 -5434 14077 -5393
rect 14111 -5315 14163 -5263
rect 14283 -5263 14292 -5255
rect 14326 -5255 14464 -5229
rect 14326 -5263 14335 -5255
rect 14111 -5349 14120 -5315
rect 14154 -5349 14163 -5315
rect 14111 -5400 14163 -5349
rect 14197 -5335 14249 -5289
rect 14197 -5369 14206 -5335
rect 14240 -5369 14249 -5335
rect 14197 -5434 14249 -5369
rect 14283 -5315 14335 -5263
rect 14455 -5263 14464 -5255
rect 14498 -5255 14636 -5229
rect 14498 -5263 14507 -5255
rect 14283 -5349 14292 -5315
rect 14326 -5349 14335 -5315
rect 14283 -5400 14335 -5349
rect 14369 -5335 14421 -5289
rect 14369 -5369 14378 -5335
rect 14412 -5369 14421 -5335
rect 14369 -5434 14421 -5369
rect 14455 -5315 14507 -5263
rect 14627 -5263 14636 -5255
rect 14670 -5255 14807 -5229
rect 14670 -5263 14679 -5255
rect 14455 -5349 14464 -5315
rect 14498 -5349 14507 -5315
rect 14455 -5400 14507 -5349
rect 14541 -5335 14593 -5289
rect 14541 -5369 14550 -5335
rect 14584 -5369 14593 -5335
rect 14541 -5434 14593 -5369
rect 14627 -5315 14679 -5263
rect 14796 -5263 14807 -5255
rect 14841 -5255 14979 -5229
rect 14841 -5263 14848 -5255
rect 14627 -5349 14636 -5315
rect 14670 -5349 14679 -5315
rect 14627 -5400 14679 -5349
rect 14713 -5335 14762 -5289
rect 14713 -5369 14722 -5335
rect 14756 -5369 14762 -5335
rect 14713 -5434 14762 -5369
rect 14796 -5315 14848 -5263
rect 14968 -5263 14979 -5255
rect 15013 -5255 15151 -5229
rect 15013 -5263 15020 -5255
rect 14796 -5349 14807 -5315
rect 14841 -5349 14848 -5315
rect 14796 -5400 14848 -5349
rect 14885 -5335 14934 -5289
rect 14885 -5369 14893 -5335
rect 14927 -5369 14934 -5335
rect 14885 -5434 14934 -5369
rect 14968 -5315 15020 -5263
rect 15140 -5263 15151 -5255
rect 15185 -5252 15323 -5229
rect 15185 -5263 15192 -5252
rect 14968 -5349 14979 -5315
rect 15013 -5349 15020 -5315
rect 14968 -5400 15020 -5349
rect 15057 -5335 15106 -5289
rect 15057 -5369 15065 -5335
rect 15099 -5369 15106 -5335
rect 15057 -5434 15106 -5369
rect 15140 -5315 15192 -5263
rect 15314 -5263 15323 -5252
rect 15357 -5252 15460 -5229
rect 15512 -5237 15570 -5202
rect 16154 -5217 16673 -5147
rect 15357 -5263 15372 -5252
rect 15140 -5349 15151 -5315
rect 15185 -5349 15192 -5315
rect 15140 -5400 15192 -5349
rect 15229 -5335 15280 -5289
rect 15229 -5369 15237 -5335
rect 15271 -5369 15280 -5335
rect 15229 -5434 15280 -5369
rect 15314 -5315 15372 -5263
rect 15512 -5271 15524 -5237
rect 15558 -5271 15570 -5237
rect 15314 -5349 15323 -5315
rect 15357 -5349 15372 -5315
rect 15314 -5400 15372 -5349
rect 15406 -5335 15460 -5286
rect 15406 -5369 15409 -5335
rect 15443 -5369 15460 -5335
rect 14025 -5435 15280 -5434
rect 15406 -5435 15460 -5369
rect 15512 -5330 15570 -5271
rect 15512 -5364 15524 -5330
rect 15558 -5364 15570 -5330
rect 15512 -5435 15570 -5364
rect 15604 -5257 16673 -5217
rect 15604 -5291 15622 -5257
rect 15656 -5291 16622 -5257
rect 16656 -5291 16673 -5257
rect 15604 -5359 16673 -5291
rect 15604 -5393 15622 -5359
rect 15656 -5393 16622 -5359
rect 16656 -5393 16673 -5359
rect 15604 -5435 16673 -5393
rect -2997 -5469 -2968 -5435
rect -2934 -5469 -2876 -5435
rect -2842 -5469 -2784 -5435
rect -2750 -5469 -2692 -5435
rect -2658 -5469 -2600 -5435
rect -2566 -5469 -2508 -5435
rect -2474 -5469 -2416 -5435
rect -2382 -5469 -2324 -5435
rect -2290 -5469 -2232 -5435
rect -2198 -5469 -2140 -5435
rect -2106 -5469 -2048 -5435
rect -2014 -5469 -1956 -5435
rect -1922 -5469 -1864 -5435
rect -1830 -5469 -1772 -5435
rect -1738 -5469 -1680 -5435
rect -1646 -5469 -1588 -5435
rect -1554 -5469 -1496 -5435
rect -1462 -5469 -1404 -5435
rect -1370 -5469 -1312 -5435
rect -1278 -5469 -1220 -5435
rect -1186 -5469 -1128 -5435
rect -1094 -5469 -1036 -5435
rect -1002 -5469 -944 -5435
rect -910 -5469 -852 -5435
rect -818 -5469 -760 -5435
rect -726 -5469 -668 -5435
rect -634 -5469 -576 -5435
rect -542 -5469 -484 -5435
rect -450 -5469 -392 -5435
rect -358 -5469 -300 -5435
rect -266 -5469 -208 -5435
rect -174 -5469 -116 -5435
rect -82 -5469 -24 -5435
rect 10 -5469 68 -5435
rect 102 -5469 160 -5435
rect 194 -5469 252 -5435
rect 286 -5469 344 -5435
rect 378 -5469 436 -5435
rect 470 -5469 528 -5435
rect 562 -5469 620 -5435
rect 654 -5469 712 -5435
rect 746 -5469 804 -5435
rect 838 -5469 896 -5435
rect 930 -5469 988 -5435
rect 1022 -5469 1080 -5435
rect 1114 -5469 1172 -5435
rect 1206 -5469 1264 -5435
rect 1298 -5469 1356 -5435
rect 1390 -5469 1448 -5435
rect 1482 -5469 1540 -5435
rect 1574 -5469 1632 -5435
rect 1666 -5469 1724 -5435
rect 1758 -5469 1816 -5435
rect 1850 -5469 1908 -5435
rect 1942 -5469 2000 -5435
rect 2034 -5469 2092 -5435
rect 2126 -5469 2184 -5435
rect 2218 -5469 2276 -5435
rect 2310 -5469 2368 -5435
rect 2402 -5469 2460 -5435
rect 2494 -5469 2552 -5435
rect 2586 -5469 2644 -5435
rect 2678 -5469 2736 -5435
rect 2770 -5469 2828 -5435
rect 2862 -5469 2920 -5435
rect 2954 -5469 3012 -5435
rect 3046 -5469 3104 -5435
rect 3138 -5469 3196 -5435
rect 3230 -5469 3288 -5435
rect 3322 -5469 3380 -5435
rect 3414 -5469 3472 -5435
rect 3506 -5469 3564 -5435
rect 3598 -5469 3656 -5435
rect 3690 -5469 3748 -5435
rect 3782 -5469 3840 -5435
rect 3874 -5469 3932 -5435
rect 3966 -5469 4024 -5435
rect 4058 -5469 4116 -5435
rect 4150 -5469 4208 -5435
rect 4242 -5469 4300 -5435
rect 4334 -5469 4392 -5435
rect 4426 -5469 4484 -5435
rect 4518 -5469 4576 -5435
rect 4610 -5469 4668 -5435
rect 4702 -5469 4760 -5435
rect 4794 -5469 4852 -5435
rect 4886 -5469 4944 -5435
rect 4978 -5469 5036 -5435
rect 5070 -5469 5128 -5435
rect 5162 -5469 5220 -5435
rect 5254 -5469 5312 -5435
rect 5346 -5469 5404 -5435
rect 5438 -5469 5496 -5435
rect 5530 -5469 5588 -5435
rect 5622 -5469 5680 -5435
rect 5714 -5469 5772 -5435
rect 5806 -5469 5864 -5435
rect 5898 -5469 5956 -5435
rect 5990 -5469 6048 -5435
rect 6082 -5469 6140 -5435
rect 6174 -5469 6232 -5435
rect 6266 -5469 6324 -5435
rect 6358 -5469 6416 -5435
rect 6450 -5469 6508 -5435
rect 6542 -5469 6600 -5435
rect 6634 -5469 6692 -5435
rect 6726 -5469 6784 -5435
rect 6818 -5469 6876 -5435
rect 6910 -5469 6968 -5435
rect 7002 -5469 7060 -5435
rect 7094 -5469 7152 -5435
rect 7186 -5469 7244 -5435
rect 7278 -5469 7336 -5435
rect 7370 -5469 7428 -5435
rect 7462 -5469 7520 -5435
rect 7554 -5469 7612 -5435
rect 7646 -5469 7704 -5435
rect 7738 -5469 7796 -5435
rect 7830 -5469 7888 -5435
rect 7922 -5469 7980 -5435
rect 8014 -5469 8072 -5435
rect 8106 -5469 8164 -5435
rect 8198 -5469 8256 -5435
rect 8290 -5469 8348 -5435
rect 8382 -5469 8440 -5435
rect 8474 -5469 8532 -5435
rect 8566 -5469 8624 -5435
rect 8658 -5469 8716 -5435
rect 8750 -5469 8808 -5435
rect 8842 -5469 8900 -5435
rect 8934 -5469 8992 -5435
rect 9026 -5469 9084 -5435
rect 9118 -5469 9176 -5435
rect 9210 -5469 9268 -5435
rect 9302 -5469 9360 -5435
rect 9394 -5469 9452 -5435
rect 9486 -5469 9544 -5435
rect 9578 -5469 9636 -5435
rect 9670 -5469 9728 -5435
rect 9762 -5469 9820 -5435
rect 9854 -5469 9912 -5435
rect 9946 -5469 10004 -5435
rect 10038 -5469 10096 -5435
rect 10130 -5469 10188 -5435
rect 10222 -5469 10280 -5435
rect 10314 -5469 10372 -5435
rect 10406 -5469 10464 -5435
rect 10498 -5469 10556 -5435
rect 10590 -5469 10648 -5435
rect 10682 -5469 10740 -5435
rect 10774 -5469 10832 -5435
rect 10866 -5469 10924 -5435
rect 10958 -5469 11016 -5435
rect 11050 -5469 11108 -5435
rect 11142 -5469 11200 -5435
rect 11234 -5469 11292 -5435
rect 11326 -5469 11384 -5435
rect 11418 -5469 11476 -5435
rect 11510 -5469 11568 -5435
rect 11602 -5469 11660 -5435
rect 11694 -5469 11752 -5435
rect 11786 -5469 11844 -5435
rect 11878 -5469 11936 -5435
rect 11970 -5469 12028 -5435
rect 12062 -5469 12120 -5435
rect 12154 -5469 12212 -5435
rect 12246 -5469 12304 -5435
rect 12338 -5469 12396 -5435
rect 12430 -5469 12488 -5435
rect 12522 -5469 12580 -5435
rect 12614 -5469 12672 -5435
rect 12706 -5469 12764 -5435
rect 12798 -5469 12856 -5435
rect 12890 -5469 12948 -5435
rect 12982 -5469 13040 -5435
rect 13074 -5469 13132 -5435
rect 13166 -5469 13224 -5435
rect 13258 -5469 13316 -5435
rect 13350 -5469 13408 -5435
rect 13442 -5469 13500 -5435
rect 13534 -5469 13592 -5435
rect 13626 -5469 13684 -5435
rect 13718 -5469 13776 -5435
rect 13810 -5469 13868 -5435
rect 13902 -5469 13960 -5435
rect 13994 -5469 14052 -5435
rect 14086 -5469 14144 -5435
rect 14178 -5469 14236 -5435
rect 14270 -5469 14328 -5435
rect 14362 -5469 14420 -5435
rect 14454 -5469 14512 -5435
rect 14546 -5469 14604 -5435
rect 14638 -5469 14696 -5435
rect 14730 -5469 14788 -5435
rect 14822 -5469 14880 -5435
rect 14914 -5469 14972 -5435
rect 15006 -5469 15064 -5435
rect 15098 -5469 15156 -5435
rect 15190 -5469 15248 -5435
rect 15282 -5469 15340 -5435
rect 15374 -5469 15432 -5435
rect 15466 -5469 15524 -5435
rect 15558 -5469 15616 -5435
rect 15650 -5469 15708 -5435
rect 15742 -5469 15800 -5435
rect 15834 -5469 15892 -5435
rect 15926 -5469 15984 -5435
rect 16018 -5469 16076 -5435
rect 16110 -5469 16168 -5435
rect 16202 -5469 16260 -5435
rect 16294 -5469 16352 -5435
rect 16386 -5469 16444 -5435
rect 16478 -5469 16536 -5435
rect 16570 -5469 16628 -5435
rect 16662 -5469 16691 -5435
rect -2980 -5511 -2278 -5469
rect -2980 -5545 -2962 -5511
rect -2928 -5545 -2330 -5511
rect -2296 -5545 -2278 -5511
rect -2980 -5613 -2278 -5545
rect -2980 -5647 -2962 -5613
rect -2928 -5647 -2330 -5613
rect -2296 -5647 -2278 -5613
rect -2980 -5687 -2278 -5647
rect -2980 -5755 -2902 -5721
rect -2868 -5755 -2803 -5721
rect -2769 -5755 -2704 -5721
rect -2670 -5755 -2650 -5721
rect -2980 -5825 -2650 -5755
rect -2616 -5757 -2278 -5687
rect -2244 -5540 -2186 -5469
rect -2244 -5574 -2232 -5540
rect -2198 -5574 -2186 -5540
rect -2244 -5633 -2186 -5574
rect -2244 -5667 -2232 -5633
rect -2198 -5667 -2186 -5633
rect -2244 -5702 -2186 -5667
rect -1600 -5511 -898 -5469
rect -1600 -5545 -1582 -5511
rect -1548 -5545 -950 -5511
rect -916 -5545 -898 -5511
rect -1600 -5613 -898 -5545
rect -1600 -5647 -1582 -5613
rect -1548 -5647 -950 -5613
rect -916 -5647 -898 -5613
rect -1600 -5687 -898 -5647
rect -864 -5511 -162 -5469
rect -864 -5545 -846 -5511
rect -812 -5545 -214 -5511
rect -180 -5545 -162 -5511
rect -864 -5613 -162 -5545
rect -864 -5647 -846 -5613
rect -812 -5647 -214 -5613
rect -180 -5647 -162 -5613
rect -864 -5687 -162 -5647
rect -128 -5540 -70 -5469
rect -128 -5574 -116 -5540
rect -82 -5574 -70 -5540
rect -128 -5633 -70 -5574
rect -128 -5667 -116 -5633
rect -82 -5667 -70 -5633
rect -2616 -5791 -2596 -5757
rect -2562 -5791 -2493 -5757
rect -2459 -5791 -2390 -5757
rect -2356 -5791 -2278 -5757
rect -1600 -5757 -1262 -5687
rect -1600 -5791 -1522 -5757
rect -1488 -5791 -1419 -5757
rect -1385 -5791 -1316 -5757
rect -1282 -5791 -1262 -5757
rect -1228 -5755 -1208 -5721
rect -1174 -5755 -1109 -5721
rect -1075 -5755 -1010 -5721
rect -976 -5755 -898 -5721
rect -1228 -5825 -898 -5755
rect -864 -5757 -526 -5687
rect -128 -5702 -70 -5667
rect -36 -5511 298 -5469
rect -36 -5545 -18 -5511
rect 16 -5545 246 -5511
rect 280 -5545 298 -5511
rect -36 -5613 298 -5545
rect -36 -5647 -18 -5613
rect 16 -5647 246 -5613
rect 280 -5647 298 -5613
rect -36 -5687 298 -5647
rect 332 -5540 390 -5469
rect 332 -5574 344 -5540
rect 378 -5574 390 -5540
rect 332 -5633 390 -5574
rect 332 -5667 344 -5633
rect 378 -5667 390 -5633
rect -864 -5791 -786 -5757
rect -752 -5791 -683 -5757
rect -649 -5791 -580 -5757
rect -546 -5791 -526 -5757
rect -492 -5755 -472 -5721
rect -438 -5755 -373 -5721
rect -339 -5755 -274 -5721
rect -240 -5755 -162 -5721
rect -492 -5825 -162 -5755
rect -36 -5757 114 -5687
rect 332 -5702 390 -5667
rect 424 -5519 505 -5503
rect 424 -5553 457 -5519
rect 491 -5553 505 -5519
rect 424 -5587 505 -5553
rect 424 -5621 457 -5587
rect 491 -5621 505 -5587
rect 424 -5658 505 -5621
rect 539 -5518 605 -5469
rect 539 -5552 555 -5518
rect 589 -5552 605 -5518
rect 539 -5586 605 -5552
rect 539 -5620 555 -5586
rect 589 -5620 605 -5586
rect 539 -5629 605 -5620
rect 695 -5519 745 -5503
rect 695 -5553 711 -5519
rect 695 -5587 745 -5553
rect 695 -5621 711 -5587
rect 424 -5708 474 -5658
rect 695 -5663 745 -5621
rect -36 -5791 -16 -5757
rect 18 -5791 114 -5757
rect 148 -5755 244 -5721
rect 278 -5755 298 -5721
rect 148 -5825 298 -5755
rect -2980 -5884 -2278 -5825
rect -2980 -5918 -2962 -5884
rect -2928 -5918 -2330 -5884
rect -2296 -5918 -2278 -5884
rect -2980 -5979 -2278 -5918
rect -2244 -5851 -2186 -5834
rect -2244 -5885 -2232 -5851
rect -2198 -5885 -2186 -5851
rect -2244 -5979 -2186 -5885
rect -1600 -5884 -898 -5825
rect -1600 -5918 -1582 -5884
rect -1548 -5918 -950 -5884
rect -916 -5918 -898 -5884
rect -1600 -5979 -898 -5918
rect -864 -5884 -162 -5825
rect -864 -5918 -846 -5884
rect -812 -5918 -214 -5884
rect -180 -5918 -162 -5884
rect -864 -5979 -162 -5918
rect -128 -5851 -70 -5834
rect -128 -5885 -116 -5851
rect -82 -5885 -70 -5851
rect -128 -5979 -70 -5885
rect -36 -5877 298 -5825
rect 424 -5742 432 -5708
rect 466 -5742 474 -5708
rect 627 -5697 745 -5663
rect 797 -5518 867 -5503
rect 797 -5552 815 -5518
rect 849 -5552 867 -5518
rect 797 -5586 867 -5552
rect 797 -5620 815 -5586
rect 849 -5620 867 -5586
rect 627 -5731 661 -5697
rect -36 -5911 -18 -5877
rect 16 -5911 246 -5877
rect 280 -5911 298 -5877
rect -36 -5979 298 -5911
rect 332 -5851 390 -5834
rect 332 -5885 344 -5851
rect 378 -5885 390 -5851
rect 332 -5979 390 -5885
rect 424 -5868 474 -5742
rect 508 -5747 661 -5731
rect 797 -5732 867 -5620
rect 957 -5518 1023 -5469
rect 957 -5552 973 -5518
rect 1007 -5552 1023 -5518
rect 957 -5586 1023 -5552
rect 957 -5620 973 -5586
rect 1007 -5620 1023 -5586
rect 957 -5636 1023 -5620
rect 1057 -5518 1126 -5503
rect 1057 -5552 1073 -5518
rect 1107 -5552 1126 -5518
rect 1057 -5586 1126 -5552
rect 1057 -5620 1073 -5586
rect 1107 -5620 1126 -5586
rect 1057 -5670 1126 -5620
rect 508 -5781 511 -5747
rect 545 -5781 661 -5747
rect 508 -5797 661 -5781
rect 695 -5747 867 -5732
rect 932 -5704 1126 -5670
rect 1160 -5540 1218 -5469
rect 1160 -5574 1172 -5540
rect 1206 -5574 1218 -5540
rect 1160 -5633 1218 -5574
rect 1160 -5667 1172 -5633
rect 1206 -5667 1218 -5633
rect 1160 -5702 1218 -5667
rect 1252 -5511 1586 -5469
rect 1252 -5545 1270 -5511
rect 1304 -5545 1534 -5511
rect 1568 -5545 1586 -5511
rect 1252 -5613 1586 -5545
rect 1252 -5647 1270 -5613
rect 1304 -5647 1534 -5613
rect 1568 -5647 1586 -5613
rect 1252 -5687 1586 -5647
rect 1620 -5540 1678 -5469
rect 1620 -5574 1632 -5540
rect 1666 -5574 1678 -5540
rect 1620 -5633 1678 -5574
rect 1620 -5667 1632 -5633
rect 1666 -5667 1678 -5633
rect 932 -5733 1002 -5704
rect 695 -5781 711 -5747
rect 745 -5781 867 -5747
rect 695 -5782 867 -5781
rect 627 -5816 661 -5797
rect 627 -5850 745 -5816
rect 424 -5892 505 -5868
rect 424 -5926 457 -5892
rect 491 -5926 505 -5892
rect 424 -5945 505 -5926
rect 539 -5892 605 -5876
rect 539 -5926 555 -5892
rect 589 -5926 605 -5892
rect 539 -5979 605 -5926
rect 695 -5892 745 -5850
rect 695 -5926 711 -5892
rect 695 -5945 745 -5926
rect 797 -5892 867 -5782
rect 916 -5747 1002 -5733
rect 916 -5781 932 -5747
rect 966 -5781 1002 -5747
rect 1036 -5743 1126 -5738
rect 1036 -5781 1052 -5743
rect 1086 -5781 1126 -5743
rect 1252 -5757 1402 -5687
rect 1620 -5702 1678 -5667
rect 1712 -5511 2414 -5469
rect 1712 -5545 1730 -5511
rect 1764 -5545 2362 -5511
rect 2396 -5545 2414 -5511
rect 1712 -5613 2414 -5545
rect 1712 -5647 1730 -5613
rect 1764 -5647 2362 -5613
rect 2396 -5647 2414 -5613
rect 1712 -5687 2414 -5647
rect 916 -5791 1002 -5781
rect 1252 -5791 1272 -5757
rect 1306 -5791 1402 -5757
rect 1436 -5755 1532 -5721
rect 1566 -5755 1586 -5721
rect 932 -5815 1002 -5791
rect 932 -5849 1126 -5815
rect 1436 -5825 1586 -5755
rect 797 -5926 816 -5892
rect 850 -5926 867 -5892
rect 797 -5945 867 -5926
rect 960 -5892 1026 -5883
rect 960 -5926 976 -5892
rect 1010 -5926 1026 -5892
rect 960 -5979 1026 -5926
rect 1060 -5892 1126 -5849
rect 1060 -5926 1073 -5892
rect 1107 -5926 1126 -5892
rect 1060 -5945 1126 -5926
rect 1160 -5851 1218 -5834
rect 1160 -5885 1172 -5851
rect 1206 -5885 1218 -5851
rect 1160 -5979 1218 -5885
rect 1252 -5877 1586 -5825
rect 1712 -5755 1790 -5721
rect 1824 -5755 1889 -5721
rect 1923 -5755 1988 -5721
rect 2022 -5755 2042 -5721
rect 1712 -5825 2042 -5755
rect 2076 -5757 2414 -5687
rect 2448 -5540 2506 -5469
rect 2448 -5574 2460 -5540
rect 2494 -5574 2506 -5540
rect 2448 -5633 2506 -5574
rect 2448 -5667 2460 -5633
rect 2494 -5667 2506 -5633
rect 2448 -5702 2506 -5667
rect 2540 -5511 2874 -5469
rect 2540 -5545 2558 -5511
rect 2592 -5545 2822 -5511
rect 2856 -5545 2874 -5511
rect 2540 -5613 2874 -5545
rect 2540 -5647 2558 -5613
rect 2592 -5647 2822 -5613
rect 2856 -5647 2874 -5613
rect 2540 -5687 2874 -5647
rect 2908 -5540 2966 -5469
rect 2908 -5574 2920 -5540
rect 2954 -5574 2966 -5540
rect 2908 -5633 2966 -5574
rect 2908 -5667 2920 -5633
rect 2954 -5667 2966 -5633
rect 2076 -5791 2096 -5757
rect 2130 -5791 2199 -5757
rect 2233 -5791 2302 -5757
rect 2336 -5791 2414 -5757
rect 2540 -5757 2690 -5687
rect 2908 -5702 2966 -5667
rect 3000 -5519 3081 -5503
rect 3000 -5553 3033 -5519
rect 3067 -5553 3081 -5519
rect 3000 -5587 3081 -5553
rect 3000 -5621 3033 -5587
rect 3067 -5621 3081 -5587
rect 3000 -5658 3081 -5621
rect 3115 -5518 3181 -5469
rect 3115 -5552 3131 -5518
rect 3165 -5552 3181 -5518
rect 3115 -5586 3181 -5552
rect 3115 -5620 3131 -5586
rect 3165 -5620 3181 -5586
rect 3115 -5629 3181 -5620
rect 3271 -5519 3321 -5503
rect 3271 -5553 3287 -5519
rect 3271 -5587 3321 -5553
rect 3271 -5621 3287 -5587
rect 2540 -5791 2560 -5757
rect 2594 -5791 2690 -5757
rect 2724 -5755 2820 -5721
rect 2854 -5755 2874 -5721
rect 2724 -5825 2874 -5755
rect 1252 -5911 1270 -5877
rect 1304 -5911 1534 -5877
rect 1568 -5911 1586 -5877
rect 1252 -5979 1586 -5911
rect 1620 -5851 1678 -5834
rect 1620 -5885 1632 -5851
rect 1666 -5885 1678 -5851
rect 1620 -5979 1678 -5885
rect 1712 -5884 2414 -5825
rect 1712 -5918 1730 -5884
rect 1764 -5918 2362 -5884
rect 2396 -5918 2414 -5884
rect 1712 -5979 2414 -5918
rect 2448 -5851 2506 -5834
rect 2448 -5885 2460 -5851
rect 2494 -5885 2506 -5851
rect 2448 -5979 2506 -5885
rect 2540 -5877 2874 -5825
rect 3000 -5743 3050 -5658
rect 3271 -5663 3321 -5621
rect 3203 -5697 3321 -5663
rect 3373 -5518 3443 -5503
rect 3373 -5552 3391 -5518
rect 3425 -5552 3443 -5518
rect 3373 -5586 3443 -5552
rect 3373 -5620 3391 -5586
rect 3425 -5620 3443 -5586
rect 3203 -5731 3237 -5697
rect 3000 -5777 3012 -5743
rect 3046 -5777 3050 -5743
rect 2540 -5911 2558 -5877
rect 2592 -5911 2822 -5877
rect 2856 -5911 2874 -5877
rect 2540 -5979 2874 -5911
rect 2908 -5851 2966 -5834
rect 2908 -5885 2920 -5851
rect 2954 -5885 2966 -5851
rect 2908 -5979 2966 -5885
rect 3000 -5868 3050 -5777
rect 3084 -5747 3237 -5731
rect 3373 -5732 3443 -5620
rect 3533 -5518 3599 -5469
rect 3533 -5552 3549 -5518
rect 3583 -5552 3599 -5518
rect 3533 -5586 3599 -5552
rect 3533 -5620 3549 -5586
rect 3583 -5620 3599 -5586
rect 3533 -5636 3599 -5620
rect 3633 -5518 3702 -5503
rect 3633 -5552 3649 -5518
rect 3683 -5552 3702 -5518
rect 3633 -5586 3702 -5552
rect 3633 -5620 3649 -5586
rect 3683 -5620 3702 -5586
rect 3633 -5670 3702 -5620
rect 3084 -5781 3087 -5747
rect 3121 -5781 3237 -5747
rect 3084 -5797 3237 -5781
rect 3271 -5747 3443 -5732
rect 3508 -5704 3702 -5670
rect 3736 -5540 3794 -5469
rect 3736 -5574 3748 -5540
rect 3782 -5574 3794 -5540
rect 3736 -5633 3794 -5574
rect 3736 -5667 3748 -5633
rect 3782 -5667 3794 -5633
rect 3736 -5702 3794 -5667
rect 3828 -5511 4162 -5469
rect 3828 -5545 3846 -5511
rect 3880 -5545 4110 -5511
rect 4144 -5545 4162 -5511
rect 3828 -5613 4162 -5545
rect 3828 -5647 3846 -5613
rect 3880 -5647 4110 -5613
rect 4144 -5647 4162 -5613
rect 3828 -5687 4162 -5647
rect 4196 -5540 4254 -5469
rect 4196 -5574 4208 -5540
rect 4242 -5574 4254 -5540
rect 4196 -5633 4254 -5574
rect 4196 -5667 4208 -5633
rect 4242 -5667 4254 -5633
rect 3508 -5733 3578 -5704
rect 3271 -5781 3287 -5747
rect 3321 -5781 3443 -5747
rect 3271 -5782 3443 -5781
rect 3203 -5816 3237 -5797
rect 3203 -5850 3321 -5816
rect 3000 -5892 3081 -5868
rect 3000 -5926 3033 -5892
rect 3067 -5926 3081 -5892
rect 3000 -5945 3081 -5926
rect 3115 -5892 3181 -5876
rect 3115 -5926 3131 -5892
rect 3165 -5926 3181 -5892
rect 3115 -5979 3181 -5926
rect 3271 -5892 3321 -5850
rect 3271 -5926 3287 -5892
rect 3271 -5945 3321 -5926
rect 3373 -5892 3443 -5782
rect 3492 -5747 3578 -5733
rect 3492 -5781 3508 -5747
rect 3542 -5781 3578 -5747
rect 3612 -5743 3702 -5738
rect 3612 -5777 3626 -5743
rect 3660 -5747 3702 -5743
rect 3612 -5781 3628 -5777
rect 3662 -5781 3702 -5747
rect 3828 -5757 3978 -5687
rect 4196 -5702 4254 -5667
rect 4288 -5511 4990 -5469
rect 4288 -5545 4306 -5511
rect 4340 -5545 4938 -5511
rect 4972 -5545 4990 -5511
rect 4288 -5613 4990 -5545
rect 4288 -5647 4306 -5613
rect 4340 -5647 4938 -5613
rect 4972 -5647 4990 -5613
rect 4288 -5687 4990 -5647
rect 3492 -5791 3578 -5781
rect 3828 -5791 3848 -5757
rect 3882 -5791 3978 -5757
rect 4012 -5755 4108 -5721
rect 4142 -5755 4162 -5721
rect 3508 -5815 3578 -5791
rect 3508 -5849 3702 -5815
rect 4012 -5825 4162 -5755
rect 3373 -5926 3392 -5892
rect 3426 -5926 3443 -5892
rect 3373 -5945 3443 -5926
rect 3536 -5892 3602 -5883
rect 3536 -5926 3552 -5892
rect 3586 -5926 3602 -5892
rect 3536 -5979 3602 -5926
rect 3636 -5892 3702 -5849
rect 3636 -5926 3649 -5892
rect 3683 -5926 3702 -5892
rect 3636 -5945 3702 -5926
rect 3736 -5851 3794 -5834
rect 3736 -5885 3748 -5851
rect 3782 -5885 3794 -5851
rect 3736 -5979 3794 -5885
rect 3828 -5877 4162 -5825
rect 4288 -5755 4366 -5721
rect 4400 -5755 4465 -5721
rect 4499 -5755 4564 -5721
rect 4598 -5755 4618 -5721
rect 4288 -5825 4618 -5755
rect 4652 -5757 4990 -5687
rect 5024 -5540 5082 -5469
rect 5024 -5574 5036 -5540
rect 5070 -5574 5082 -5540
rect 5024 -5633 5082 -5574
rect 5024 -5667 5036 -5633
rect 5070 -5667 5082 -5633
rect 5024 -5702 5082 -5667
rect 5116 -5511 5450 -5469
rect 5116 -5545 5134 -5511
rect 5168 -5545 5398 -5511
rect 5432 -5545 5450 -5511
rect 5116 -5613 5450 -5545
rect 5116 -5647 5134 -5613
rect 5168 -5647 5398 -5613
rect 5432 -5647 5450 -5613
rect 5116 -5687 5450 -5647
rect 5484 -5540 5542 -5469
rect 5484 -5574 5496 -5540
rect 5530 -5574 5542 -5540
rect 5484 -5633 5542 -5574
rect 5484 -5667 5496 -5633
rect 5530 -5667 5542 -5633
rect 4652 -5791 4672 -5757
rect 4706 -5791 4775 -5757
rect 4809 -5791 4878 -5757
rect 4912 -5791 4990 -5757
rect 5116 -5757 5266 -5687
rect 5484 -5702 5542 -5667
rect 5576 -5519 5657 -5503
rect 5576 -5553 5609 -5519
rect 5643 -5553 5657 -5519
rect 5576 -5587 5657 -5553
rect 5576 -5621 5609 -5587
rect 5643 -5621 5657 -5587
rect 5576 -5658 5657 -5621
rect 5691 -5518 5757 -5469
rect 5691 -5552 5707 -5518
rect 5741 -5552 5757 -5518
rect 5691 -5586 5757 -5552
rect 5691 -5620 5707 -5586
rect 5741 -5620 5757 -5586
rect 5691 -5629 5757 -5620
rect 5847 -5519 5897 -5503
rect 5847 -5553 5863 -5519
rect 5847 -5587 5897 -5553
rect 5847 -5621 5863 -5587
rect 5116 -5791 5136 -5757
rect 5170 -5791 5266 -5757
rect 5300 -5755 5396 -5721
rect 5430 -5755 5450 -5721
rect 5300 -5825 5450 -5755
rect 3828 -5911 3846 -5877
rect 3880 -5911 4110 -5877
rect 4144 -5911 4162 -5877
rect 3828 -5979 4162 -5911
rect 4196 -5851 4254 -5834
rect 4196 -5885 4208 -5851
rect 4242 -5885 4254 -5851
rect 4196 -5979 4254 -5885
rect 4288 -5884 4990 -5825
rect 4288 -5918 4306 -5884
rect 4340 -5918 4938 -5884
rect 4972 -5918 4990 -5884
rect 4288 -5979 4990 -5918
rect 5024 -5851 5082 -5834
rect 5024 -5885 5036 -5851
rect 5070 -5885 5082 -5851
rect 5024 -5979 5082 -5885
rect 5116 -5877 5450 -5825
rect 5576 -5743 5626 -5658
rect 5847 -5663 5897 -5621
rect 5779 -5697 5897 -5663
rect 5949 -5518 6019 -5503
rect 5949 -5552 5967 -5518
rect 6001 -5552 6019 -5518
rect 5949 -5586 6019 -5552
rect 5949 -5620 5967 -5586
rect 6001 -5620 6019 -5586
rect 5779 -5731 5813 -5697
rect 5576 -5777 5586 -5743
rect 5620 -5777 5626 -5743
rect 5116 -5911 5134 -5877
rect 5168 -5911 5398 -5877
rect 5432 -5911 5450 -5877
rect 5116 -5979 5450 -5911
rect 5484 -5851 5542 -5834
rect 5484 -5885 5496 -5851
rect 5530 -5885 5542 -5851
rect 5484 -5979 5542 -5885
rect 5576 -5868 5626 -5777
rect 5660 -5747 5813 -5731
rect 5949 -5732 6019 -5620
rect 6109 -5518 6175 -5469
rect 6109 -5552 6125 -5518
rect 6159 -5552 6175 -5518
rect 6109 -5586 6175 -5552
rect 6109 -5620 6125 -5586
rect 6159 -5620 6175 -5586
rect 6109 -5636 6175 -5620
rect 6209 -5518 6278 -5503
rect 6209 -5552 6225 -5518
rect 6259 -5552 6278 -5518
rect 6209 -5586 6278 -5552
rect 6209 -5620 6225 -5586
rect 6259 -5620 6278 -5586
rect 6209 -5670 6278 -5620
rect 5660 -5781 5663 -5747
rect 5697 -5781 5813 -5747
rect 5660 -5797 5813 -5781
rect 5847 -5747 6019 -5732
rect 6084 -5704 6278 -5670
rect 6312 -5540 6370 -5469
rect 6312 -5574 6324 -5540
rect 6358 -5574 6370 -5540
rect 6312 -5633 6370 -5574
rect 6312 -5667 6324 -5633
rect 6358 -5667 6370 -5633
rect 6312 -5702 6370 -5667
rect 6404 -5511 6738 -5469
rect 6404 -5545 6422 -5511
rect 6456 -5545 6686 -5511
rect 6720 -5545 6738 -5511
rect 6404 -5613 6738 -5545
rect 6404 -5647 6422 -5613
rect 6456 -5647 6686 -5613
rect 6720 -5647 6738 -5613
rect 6404 -5687 6738 -5647
rect 6772 -5540 6830 -5469
rect 6772 -5574 6784 -5540
rect 6818 -5574 6830 -5540
rect 6772 -5633 6830 -5574
rect 6772 -5667 6784 -5633
rect 6818 -5667 6830 -5633
rect 6084 -5733 6154 -5704
rect 5847 -5781 5863 -5747
rect 5897 -5781 6019 -5747
rect 5847 -5782 6019 -5781
rect 5779 -5816 5813 -5797
rect 5779 -5850 5897 -5816
rect 5576 -5892 5657 -5868
rect 5576 -5926 5609 -5892
rect 5643 -5926 5657 -5892
rect 5576 -5945 5657 -5926
rect 5691 -5892 5757 -5876
rect 5691 -5926 5707 -5892
rect 5741 -5926 5757 -5892
rect 5691 -5979 5757 -5926
rect 5847 -5892 5897 -5850
rect 5847 -5926 5863 -5892
rect 5847 -5945 5897 -5926
rect 5949 -5892 6019 -5782
rect 6068 -5747 6154 -5733
rect 6068 -5781 6084 -5747
rect 6118 -5781 6154 -5747
rect 6188 -5743 6278 -5738
rect 6188 -5777 6200 -5743
rect 6234 -5747 6278 -5743
rect 6188 -5781 6204 -5777
rect 6238 -5781 6278 -5747
rect 6404 -5757 6554 -5687
rect 6772 -5702 6830 -5667
rect 6864 -5511 7566 -5469
rect 6864 -5545 6882 -5511
rect 6916 -5545 7514 -5511
rect 7548 -5545 7566 -5511
rect 6864 -5613 7566 -5545
rect 6864 -5647 6882 -5613
rect 6916 -5647 7514 -5613
rect 7548 -5647 7566 -5613
rect 6864 -5687 7566 -5647
rect 6068 -5791 6154 -5781
rect 6404 -5791 6424 -5757
rect 6458 -5791 6554 -5757
rect 6588 -5755 6684 -5721
rect 6718 -5755 6738 -5721
rect 6084 -5815 6154 -5791
rect 6084 -5849 6278 -5815
rect 6588 -5825 6738 -5755
rect 5949 -5926 5968 -5892
rect 6002 -5926 6019 -5892
rect 5949 -5945 6019 -5926
rect 6112 -5892 6178 -5883
rect 6112 -5926 6128 -5892
rect 6162 -5926 6178 -5892
rect 6112 -5979 6178 -5926
rect 6212 -5892 6278 -5849
rect 6212 -5926 6225 -5892
rect 6259 -5926 6278 -5892
rect 6212 -5945 6278 -5926
rect 6312 -5851 6370 -5834
rect 6312 -5885 6324 -5851
rect 6358 -5885 6370 -5851
rect 6312 -5979 6370 -5885
rect 6404 -5877 6738 -5825
rect 6864 -5755 6942 -5721
rect 6976 -5755 7041 -5721
rect 7075 -5755 7140 -5721
rect 7174 -5755 7194 -5721
rect 6864 -5825 7194 -5755
rect 7228 -5757 7566 -5687
rect 7600 -5540 7658 -5469
rect 7600 -5574 7612 -5540
rect 7646 -5574 7658 -5540
rect 7600 -5633 7658 -5574
rect 7600 -5667 7612 -5633
rect 7646 -5667 7658 -5633
rect 7600 -5702 7658 -5667
rect 7692 -5511 8026 -5469
rect 7692 -5545 7710 -5511
rect 7744 -5545 7974 -5511
rect 8008 -5545 8026 -5511
rect 7692 -5613 8026 -5545
rect 7692 -5647 7710 -5613
rect 7744 -5647 7974 -5613
rect 8008 -5647 8026 -5613
rect 7692 -5687 8026 -5647
rect 8060 -5540 8118 -5469
rect 8060 -5574 8072 -5540
rect 8106 -5574 8118 -5540
rect 8060 -5633 8118 -5574
rect 8060 -5667 8072 -5633
rect 8106 -5667 8118 -5633
rect 7228 -5791 7248 -5757
rect 7282 -5791 7351 -5757
rect 7385 -5791 7454 -5757
rect 7488 -5791 7566 -5757
rect 7692 -5757 7842 -5687
rect 8060 -5702 8118 -5667
rect 8152 -5519 8233 -5503
rect 8152 -5553 8185 -5519
rect 8219 -5553 8233 -5519
rect 8152 -5587 8233 -5553
rect 8152 -5621 8185 -5587
rect 8219 -5621 8233 -5587
rect 8152 -5658 8233 -5621
rect 8267 -5518 8333 -5469
rect 8267 -5552 8283 -5518
rect 8317 -5552 8333 -5518
rect 8267 -5586 8333 -5552
rect 8267 -5620 8283 -5586
rect 8317 -5620 8333 -5586
rect 8267 -5629 8333 -5620
rect 8423 -5519 8473 -5503
rect 8423 -5553 8439 -5519
rect 8423 -5587 8473 -5553
rect 8423 -5621 8439 -5587
rect 7692 -5791 7712 -5757
rect 7746 -5791 7842 -5757
rect 7876 -5755 7972 -5721
rect 8006 -5755 8026 -5721
rect 7876 -5825 8026 -5755
rect 6404 -5911 6422 -5877
rect 6456 -5911 6686 -5877
rect 6720 -5911 6738 -5877
rect 6404 -5979 6738 -5911
rect 6772 -5851 6830 -5834
rect 6772 -5885 6784 -5851
rect 6818 -5885 6830 -5851
rect 6772 -5979 6830 -5885
rect 6864 -5884 7566 -5825
rect 6864 -5918 6882 -5884
rect 6916 -5918 7514 -5884
rect 7548 -5918 7566 -5884
rect 6864 -5979 7566 -5918
rect 7600 -5851 7658 -5834
rect 7600 -5885 7612 -5851
rect 7646 -5885 7658 -5851
rect 7600 -5979 7658 -5885
rect 7692 -5877 8026 -5825
rect 8152 -5743 8202 -5658
rect 8423 -5663 8473 -5621
rect 8355 -5697 8473 -5663
rect 8525 -5518 8595 -5503
rect 8525 -5552 8543 -5518
rect 8577 -5552 8595 -5518
rect 8525 -5586 8595 -5552
rect 8525 -5620 8543 -5586
rect 8577 -5620 8595 -5586
rect 8355 -5731 8389 -5697
rect 8152 -5777 8160 -5743
rect 8194 -5777 8202 -5743
rect 7692 -5911 7710 -5877
rect 7744 -5911 7974 -5877
rect 8008 -5911 8026 -5877
rect 7692 -5979 8026 -5911
rect 8060 -5851 8118 -5834
rect 8060 -5885 8072 -5851
rect 8106 -5885 8118 -5851
rect 8060 -5979 8118 -5885
rect 8152 -5868 8202 -5777
rect 8236 -5747 8389 -5731
rect 8525 -5732 8595 -5620
rect 8685 -5518 8751 -5469
rect 8685 -5552 8701 -5518
rect 8735 -5552 8751 -5518
rect 8685 -5586 8751 -5552
rect 8685 -5620 8701 -5586
rect 8735 -5620 8751 -5586
rect 8685 -5636 8751 -5620
rect 8785 -5518 8854 -5503
rect 8785 -5552 8801 -5518
rect 8835 -5552 8854 -5518
rect 8785 -5586 8854 -5552
rect 8785 -5620 8801 -5586
rect 8835 -5620 8854 -5586
rect 8785 -5670 8854 -5620
rect 8236 -5781 8239 -5747
rect 8273 -5781 8389 -5747
rect 8236 -5797 8389 -5781
rect 8423 -5747 8595 -5732
rect 8660 -5704 8854 -5670
rect 8888 -5540 8946 -5469
rect 8888 -5574 8900 -5540
rect 8934 -5574 8946 -5540
rect 8888 -5633 8946 -5574
rect 8888 -5667 8900 -5633
rect 8934 -5667 8946 -5633
rect 8888 -5702 8946 -5667
rect 8980 -5511 9314 -5469
rect 8980 -5545 8998 -5511
rect 9032 -5545 9262 -5511
rect 9296 -5545 9314 -5511
rect 8980 -5613 9314 -5545
rect 8980 -5647 8998 -5613
rect 9032 -5647 9262 -5613
rect 9296 -5647 9314 -5613
rect 8980 -5687 9314 -5647
rect 9348 -5540 9406 -5469
rect 9348 -5574 9360 -5540
rect 9394 -5574 9406 -5540
rect 9348 -5633 9406 -5574
rect 9348 -5667 9360 -5633
rect 9394 -5667 9406 -5633
rect 8660 -5733 8730 -5704
rect 8423 -5781 8439 -5747
rect 8473 -5781 8595 -5747
rect 8423 -5782 8595 -5781
rect 8355 -5816 8389 -5797
rect 8355 -5850 8473 -5816
rect 8152 -5892 8233 -5868
rect 8152 -5926 8185 -5892
rect 8219 -5926 8233 -5892
rect 8152 -5945 8233 -5926
rect 8267 -5892 8333 -5876
rect 8267 -5926 8283 -5892
rect 8317 -5926 8333 -5892
rect 8267 -5979 8333 -5926
rect 8423 -5892 8473 -5850
rect 8423 -5926 8439 -5892
rect 8423 -5945 8473 -5926
rect 8525 -5892 8595 -5782
rect 8644 -5747 8730 -5733
rect 8644 -5781 8660 -5747
rect 8694 -5781 8730 -5747
rect 8764 -5743 8854 -5738
rect 8764 -5777 8774 -5743
rect 8808 -5747 8854 -5743
rect 8764 -5781 8780 -5777
rect 8814 -5781 8854 -5747
rect 8980 -5757 9130 -5687
rect 9348 -5702 9406 -5667
rect 9440 -5511 10142 -5469
rect 9440 -5545 9458 -5511
rect 9492 -5545 10090 -5511
rect 10124 -5545 10142 -5511
rect 9440 -5613 10142 -5545
rect 9440 -5647 9458 -5613
rect 9492 -5647 10090 -5613
rect 10124 -5647 10142 -5613
rect 9440 -5687 10142 -5647
rect 8644 -5791 8730 -5781
rect 8980 -5791 9000 -5757
rect 9034 -5791 9130 -5757
rect 9164 -5755 9260 -5721
rect 9294 -5755 9314 -5721
rect 8660 -5815 8730 -5791
rect 8660 -5849 8854 -5815
rect 9164 -5825 9314 -5755
rect 8525 -5926 8544 -5892
rect 8578 -5926 8595 -5892
rect 8525 -5945 8595 -5926
rect 8688 -5892 8754 -5883
rect 8688 -5926 8704 -5892
rect 8738 -5926 8754 -5892
rect 8688 -5979 8754 -5926
rect 8788 -5892 8854 -5849
rect 8788 -5926 8801 -5892
rect 8835 -5926 8854 -5892
rect 8788 -5945 8854 -5926
rect 8888 -5851 8946 -5834
rect 8888 -5885 8900 -5851
rect 8934 -5885 8946 -5851
rect 8888 -5979 8946 -5885
rect 8980 -5877 9314 -5825
rect 9440 -5755 9518 -5721
rect 9552 -5755 9617 -5721
rect 9651 -5755 9716 -5721
rect 9750 -5755 9770 -5721
rect 9440 -5825 9770 -5755
rect 9804 -5757 10142 -5687
rect 10176 -5540 10234 -5469
rect 10176 -5574 10188 -5540
rect 10222 -5574 10234 -5540
rect 10176 -5633 10234 -5574
rect 10176 -5667 10188 -5633
rect 10222 -5667 10234 -5633
rect 10176 -5702 10234 -5667
rect 10360 -5511 10694 -5469
rect 10360 -5545 10378 -5511
rect 10412 -5545 10642 -5511
rect 10676 -5545 10694 -5511
rect 10360 -5613 10694 -5545
rect 10360 -5647 10378 -5613
rect 10412 -5647 10642 -5613
rect 10676 -5647 10694 -5613
rect 10360 -5687 10694 -5647
rect 10728 -5519 10809 -5503
rect 10728 -5553 10761 -5519
rect 10795 -5553 10809 -5519
rect 10728 -5587 10809 -5553
rect 10728 -5621 10761 -5587
rect 10795 -5621 10809 -5587
rect 10728 -5658 10809 -5621
rect 10843 -5518 10909 -5469
rect 10843 -5552 10859 -5518
rect 10893 -5552 10909 -5518
rect 10843 -5586 10909 -5552
rect 10843 -5620 10859 -5586
rect 10893 -5620 10909 -5586
rect 10843 -5629 10909 -5620
rect 10999 -5519 11049 -5503
rect 10999 -5553 11015 -5519
rect 10999 -5587 11049 -5553
rect 10999 -5621 11015 -5587
rect 9804 -5791 9824 -5757
rect 9858 -5791 9927 -5757
rect 9961 -5791 10030 -5757
rect 10064 -5791 10142 -5757
rect 10360 -5757 10510 -5687
rect 10360 -5791 10380 -5757
rect 10414 -5791 10510 -5757
rect 10544 -5755 10640 -5721
rect 10674 -5755 10694 -5721
rect 10544 -5825 10694 -5755
rect 8980 -5911 8998 -5877
rect 9032 -5911 9262 -5877
rect 9296 -5911 9314 -5877
rect 8980 -5979 9314 -5911
rect 9348 -5851 9406 -5834
rect 9348 -5885 9360 -5851
rect 9394 -5885 9406 -5851
rect 9348 -5979 9406 -5885
rect 9440 -5884 10142 -5825
rect 9440 -5918 9458 -5884
rect 9492 -5918 10090 -5884
rect 10124 -5918 10142 -5884
rect 9440 -5979 10142 -5918
rect 10176 -5851 10234 -5834
rect 10176 -5885 10188 -5851
rect 10222 -5885 10234 -5851
rect 10176 -5979 10234 -5885
rect 10360 -5877 10694 -5825
rect 10360 -5911 10378 -5877
rect 10412 -5911 10642 -5877
rect 10676 -5911 10694 -5877
rect 10360 -5979 10694 -5911
rect 10728 -5741 10778 -5658
rect 10999 -5663 11049 -5621
rect 10931 -5697 11049 -5663
rect 11101 -5518 11171 -5503
rect 11101 -5552 11119 -5518
rect 11153 -5552 11171 -5518
rect 11101 -5586 11171 -5552
rect 11101 -5620 11119 -5586
rect 11153 -5620 11171 -5586
rect 10931 -5731 10965 -5697
rect 10728 -5775 10737 -5741
rect 10771 -5775 10778 -5741
rect 10728 -5868 10778 -5775
rect 10812 -5747 10965 -5731
rect 11101 -5732 11171 -5620
rect 11261 -5518 11327 -5469
rect 11261 -5552 11277 -5518
rect 11311 -5552 11327 -5518
rect 11261 -5586 11327 -5552
rect 11261 -5620 11277 -5586
rect 11311 -5620 11327 -5586
rect 11261 -5636 11327 -5620
rect 11361 -5518 11430 -5503
rect 11361 -5552 11377 -5518
rect 11411 -5552 11430 -5518
rect 11361 -5586 11430 -5552
rect 11361 -5620 11377 -5586
rect 11411 -5620 11430 -5586
rect 11361 -5670 11430 -5620
rect 10812 -5781 10815 -5747
rect 10849 -5781 10965 -5747
rect 10812 -5797 10965 -5781
rect 10999 -5747 11171 -5732
rect 11236 -5704 11430 -5670
rect 11464 -5540 11522 -5469
rect 11464 -5574 11476 -5540
rect 11510 -5574 11522 -5540
rect 11464 -5633 11522 -5574
rect 11464 -5667 11476 -5633
rect 11510 -5667 11522 -5633
rect 11464 -5702 11522 -5667
rect 11648 -5511 11982 -5469
rect 11648 -5545 11666 -5511
rect 11700 -5545 11930 -5511
rect 11964 -5545 11982 -5511
rect 11648 -5613 11982 -5545
rect 11648 -5647 11666 -5613
rect 11700 -5647 11930 -5613
rect 11964 -5647 11982 -5613
rect 11648 -5687 11982 -5647
rect 13580 -5540 13638 -5469
rect 13580 -5574 13592 -5540
rect 13626 -5574 13638 -5540
rect 13580 -5633 13638 -5574
rect 13674 -5511 13733 -5469
rect 13674 -5545 13690 -5511
rect 13724 -5545 13733 -5511
rect 13674 -5579 13733 -5545
rect 13674 -5613 13690 -5579
rect 13724 -5613 13733 -5579
rect 13674 -5631 13733 -5613
rect 13769 -5519 13818 -5503
rect 13769 -5553 13776 -5519
rect 13810 -5553 13818 -5519
rect 13769 -5587 13818 -5553
rect 13769 -5621 13776 -5587
rect 13810 -5621 13818 -5587
rect 13580 -5667 13592 -5633
rect 13626 -5667 13638 -5633
rect 11236 -5733 11306 -5704
rect 10999 -5781 11015 -5747
rect 11049 -5781 11171 -5747
rect 10999 -5782 11171 -5781
rect 10931 -5816 10965 -5797
rect 10931 -5850 11049 -5816
rect 10728 -5892 10809 -5868
rect 10728 -5926 10761 -5892
rect 10795 -5926 10809 -5892
rect 10728 -5945 10809 -5926
rect 10843 -5892 10909 -5876
rect 10843 -5926 10859 -5892
rect 10893 -5926 10909 -5892
rect 10843 -5979 10909 -5926
rect 10999 -5892 11049 -5850
rect 10999 -5926 11015 -5892
rect 10999 -5945 11049 -5926
rect 11101 -5892 11171 -5782
rect 11220 -5747 11306 -5733
rect 11220 -5781 11236 -5747
rect 11270 -5781 11306 -5747
rect 11340 -5740 11430 -5738
rect 11340 -5747 11369 -5740
rect 11340 -5781 11356 -5747
rect 11403 -5774 11430 -5740
rect 11390 -5781 11430 -5774
rect 11648 -5757 11798 -5687
rect 13580 -5702 13638 -5667
rect 11220 -5791 11306 -5781
rect 11648 -5791 11668 -5757
rect 11702 -5791 11798 -5757
rect 11832 -5755 11928 -5721
rect 11962 -5755 11982 -5721
rect 13769 -5731 13818 -5621
rect 13853 -5511 13905 -5469
rect 14025 -5470 15280 -5469
rect 13853 -5545 13862 -5511
rect 13896 -5545 13905 -5511
rect 13853 -5579 13905 -5545
rect 13853 -5613 13862 -5579
rect 13896 -5613 13905 -5579
rect 13853 -5631 13905 -5613
rect 13941 -5527 13991 -5504
rect 13941 -5561 13948 -5527
rect 13982 -5561 13991 -5527
rect 13941 -5595 13991 -5561
rect 13941 -5629 13948 -5595
rect 13982 -5629 13991 -5595
rect 14025 -5511 14077 -5470
rect 14025 -5545 14034 -5511
rect 14068 -5545 14077 -5511
rect 14025 -5579 14077 -5545
rect 14025 -5613 14034 -5579
rect 14068 -5613 14077 -5579
rect 14025 -5629 14077 -5613
rect 14111 -5555 14163 -5504
rect 14111 -5589 14120 -5555
rect 14154 -5589 14163 -5555
rect 13941 -5731 13991 -5629
rect 14111 -5641 14163 -5589
rect 14197 -5535 14249 -5470
rect 14197 -5569 14206 -5535
rect 14240 -5569 14249 -5535
rect 14197 -5615 14249 -5569
rect 14283 -5555 14335 -5504
rect 14283 -5589 14292 -5555
rect 14326 -5589 14335 -5555
rect 14111 -5675 14120 -5641
rect 14154 -5649 14163 -5641
rect 14283 -5641 14335 -5589
rect 14369 -5535 14421 -5470
rect 14369 -5569 14378 -5535
rect 14412 -5569 14421 -5535
rect 14369 -5615 14421 -5569
rect 14455 -5555 14507 -5504
rect 14455 -5589 14464 -5555
rect 14498 -5589 14507 -5555
rect 14283 -5649 14292 -5641
rect 14154 -5675 14292 -5649
rect 14326 -5649 14335 -5641
rect 14455 -5641 14507 -5589
rect 14541 -5535 14593 -5470
rect 14541 -5569 14550 -5535
rect 14584 -5569 14593 -5535
rect 14541 -5615 14593 -5569
rect 14627 -5555 14679 -5504
rect 14627 -5589 14636 -5555
rect 14670 -5589 14679 -5555
rect 14455 -5649 14464 -5641
rect 14326 -5675 14464 -5649
rect 14498 -5649 14507 -5641
rect 14627 -5641 14679 -5589
rect 14713 -5535 14762 -5470
rect 14713 -5569 14722 -5535
rect 14756 -5569 14762 -5535
rect 14713 -5615 14762 -5569
rect 14796 -5555 14848 -5504
rect 14796 -5589 14807 -5555
rect 14841 -5589 14848 -5555
rect 14627 -5649 14636 -5641
rect 14498 -5675 14636 -5649
rect 14670 -5649 14679 -5641
rect 14796 -5641 14848 -5589
rect 14885 -5535 14934 -5470
rect 14885 -5569 14893 -5535
rect 14927 -5569 14934 -5535
rect 14885 -5615 14934 -5569
rect 14968 -5555 15020 -5504
rect 14968 -5589 14979 -5555
rect 15013 -5589 15020 -5555
rect 14796 -5649 14807 -5641
rect 14670 -5675 14807 -5649
rect 14841 -5649 14848 -5641
rect 14968 -5641 15020 -5589
rect 15057 -5535 15106 -5470
rect 15057 -5569 15065 -5535
rect 15099 -5569 15106 -5535
rect 15057 -5615 15106 -5569
rect 15140 -5555 15192 -5504
rect 15140 -5589 15151 -5555
rect 15185 -5589 15192 -5555
rect 14968 -5649 14979 -5641
rect 14841 -5675 14979 -5649
rect 15013 -5649 15020 -5641
rect 15140 -5641 15192 -5589
rect 15229 -5535 15280 -5470
rect 15229 -5569 15237 -5535
rect 15271 -5569 15280 -5535
rect 15229 -5615 15280 -5569
rect 15314 -5555 15372 -5504
rect 15314 -5589 15323 -5555
rect 15357 -5589 15372 -5555
rect 15140 -5649 15151 -5641
rect 15013 -5675 15151 -5649
rect 15185 -5652 15192 -5641
rect 15314 -5641 15372 -5589
rect 15406 -5535 15460 -5469
rect 15406 -5569 15409 -5535
rect 15443 -5569 15460 -5535
rect 15406 -5618 15460 -5569
rect 15512 -5540 15570 -5469
rect 15512 -5574 15524 -5540
rect 15558 -5574 15570 -5540
rect 15314 -5652 15323 -5641
rect 15185 -5675 15323 -5652
rect 15357 -5652 15372 -5641
rect 15512 -5633 15570 -5574
rect 15357 -5675 15460 -5652
rect 14111 -5694 15460 -5675
rect 14111 -5697 15248 -5694
rect 15227 -5728 15248 -5697
rect 15282 -5728 15341 -5694
rect 15375 -5728 15460 -5694
rect 15512 -5667 15524 -5633
rect 15558 -5667 15570 -5633
rect 15512 -5702 15570 -5667
rect 15605 -5511 16674 -5469
rect 15605 -5545 15622 -5511
rect 15656 -5545 16622 -5511
rect 16656 -5545 16674 -5511
rect 15605 -5613 16674 -5545
rect 15605 -5647 15622 -5613
rect 15656 -5647 16622 -5613
rect 16656 -5647 16674 -5613
rect 15605 -5687 16674 -5647
rect 11236 -5815 11306 -5791
rect 11236 -5849 11430 -5815
rect 11832 -5825 11982 -5755
rect 11101 -5926 11120 -5892
rect 11154 -5926 11171 -5892
rect 11101 -5945 11171 -5926
rect 11264 -5892 11330 -5883
rect 11264 -5926 11280 -5892
rect 11314 -5926 11330 -5892
rect 11264 -5979 11330 -5926
rect 11364 -5892 11430 -5849
rect 11364 -5926 11377 -5892
rect 11411 -5926 11430 -5892
rect 11364 -5945 11430 -5926
rect 11464 -5851 11522 -5834
rect 11464 -5885 11476 -5851
rect 11510 -5885 11522 -5851
rect 11464 -5979 11522 -5885
rect 11648 -5877 11982 -5825
rect 13672 -5747 13735 -5731
rect 13672 -5772 13692 -5747
rect 13672 -5806 13685 -5772
rect 13726 -5781 13735 -5747
rect 13719 -5806 13735 -5781
rect 11648 -5911 11666 -5877
rect 11700 -5911 11930 -5877
rect 11964 -5911 11982 -5877
rect 11648 -5979 11982 -5911
rect 13580 -5851 13638 -5834
rect 13672 -5843 13735 -5806
rect 13769 -5747 15193 -5731
rect 13769 -5781 14119 -5747
rect 14153 -5781 14187 -5747
rect 14221 -5781 14255 -5747
rect 14289 -5781 14323 -5747
rect 14357 -5781 14391 -5747
rect 14425 -5781 14459 -5747
rect 14493 -5781 14527 -5747
rect 14561 -5781 14595 -5747
rect 14629 -5781 14663 -5747
rect 14697 -5781 14731 -5747
rect 14765 -5781 14799 -5747
rect 14833 -5781 14867 -5747
rect 14901 -5781 14935 -5747
rect 14969 -5781 15003 -5747
rect 15037 -5781 15071 -5747
rect 15105 -5781 15139 -5747
rect 15173 -5781 15193 -5747
rect 13580 -5885 13592 -5851
rect 13626 -5885 13638 -5851
rect 13580 -5979 13638 -5885
rect 13672 -5903 13733 -5877
rect 13672 -5937 13690 -5903
rect 13724 -5937 13733 -5903
rect 13672 -5979 13733 -5937
rect 13769 -5890 13819 -5781
rect 13769 -5924 13776 -5890
rect 13810 -5924 13819 -5890
rect 13769 -5943 13819 -5924
rect 13853 -5890 13905 -5874
rect 13853 -5924 13862 -5890
rect 13896 -5924 13905 -5890
rect 13853 -5979 13905 -5924
rect 13941 -5890 13991 -5781
rect 15227 -5789 15460 -5728
rect 15227 -5790 15340 -5789
rect 15227 -5815 15248 -5790
rect 14111 -5824 15248 -5815
rect 15282 -5823 15340 -5790
rect 15374 -5823 15460 -5789
rect 15605 -5757 16124 -5687
rect 15605 -5791 15686 -5757
rect 15720 -5791 15814 -5757
rect 15848 -5791 15942 -5757
rect 15976 -5791 16070 -5757
rect 16104 -5791 16124 -5757
rect 16158 -5755 16178 -5721
rect 16212 -5755 16306 -5721
rect 16340 -5755 16434 -5721
rect 16468 -5755 16562 -5721
rect 16596 -5755 16674 -5721
rect 15282 -5824 15460 -5823
rect 14111 -5849 15460 -5824
rect 16158 -5825 16674 -5755
rect 13941 -5924 13948 -5890
rect 13982 -5924 13991 -5890
rect 13941 -5943 13991 -5924
rect 14025 -5890 14077 -5867
rect 14025 -5924 14034 -5890
rect 14068 -5924 14077 -5890
rect 14025 -5979 14077 -5924
rect 14111 -5890 14163 -5849
rect 14111 -5924 14120 -5890
rect 14154 -5924 14163 -5890
rect 14111 -5940 14163 -5924
rect 14197 -5899 14249 -5883
rect 14197 -5933 14206 -5899
rect 14240 -5933 14249 -5899
rect 14197 -5979 14249 -5933
rect 14283 -5890 14335 -5849
rect 14283 -5924 14292 -5890
rect 14326 -5924 14335 -5890
rect 14283 -5940 14335 -5924
rect 14369 -5899 14421 -5883
rect 14369 -5933 14378 -5899
rect 14412 -5933 14421 -5899
rect 14369 -5979 14421 -5933
rect 14455 -5890 14507 -5849
rect 14455 -5924 14464 -5890
rect 14498 -5924 14507 -5890
rect 14455 -5940 14507 -5924
rect 14541 -5899 14590 -5883
rect 14541 -5933 14550 -5899
rect 14584 -5933 14590 -5899
rect 14541 -5979 14590 -5933
rect 14624 -5890 14679 -5849
rect 14624 -5924 14636 -5890
rect 14670 -5924 14679 -5890
rect 14624 -5940 14679 -5924
rect 14713 -5899 14762 -5883
rect 14713 -5933 14722 -5899
rect 14756 -5933 14762 -5899
rect 14713 -5979 14762 -5933
rect 14796 -5890 14848 -5849
rect 14796 -5924 14807 -5890
rect 14841 -5924 14848 -5890
rect 14796 -5940 14848 -5924
rect 14884 -5899 14934 -5883
rect 14884 -5933 14893 -5899
rect 14927 -5933 14934 -5899
rect 14884 -5979 14934 -5933
rect 14968 -5890 15020 -5849
rect 14968 -5924 14979 -5890
rect 15013 -5924 15020 -5890
rect 14968 -5940 15020 -5924
rect 15056 -5899 15106 -5883
rect 15056 -5933 15065 -5899
rect 15099 -5933 15106 -5899
rect 15056 -5979 15106 -5933
rect 15140 -5890 15192 -5849
rect 15140 -5924 15151 -5890
rect 15185 -5924 15192 -5890
rect 15140 -5940 15192 -5924
rect 15228 -5899 15280 -5883
rect 15228 -5933 15237 -5899
rect 15271 -5933 15280 -5899
rect 15228 -5979 15280 -5933
rect 15314 -5890 15366 -5849
rect 15512 -5851 15570 -5834
rect 15314 -5924 15323 -5890
rect 15357 -5924 15366 -5890
rect 15314 -5940 15366 -5924
rect 15400 -5899 15460 -5883
rect 15400 -5933 15409 -5899
rect 15443 -5933 15460 -5899
rect 15400 -5979 15460 -5933
rect 15512 -5885 15524 -5851
rect 15558 -5885 15570 -5851
rect 15512 -5979 15570 -5885
rect 15605 -5884 16674 -5825
rect 15605 -5918 15622 -5884
rect 15656 -5918 16622 -5884
rect 16656 -5918 16674 -5884
rect 15605 -5979 16674 -5918
rect -2997 -6013 -2968 -5979
rect -2934 -6013 -2876 -5979
rect -2842 -6013 -2784 -5979
rect -2750 -6013 -2692 -5979
rect -2658 -6013 -2600 -5979
rect -2566 -6013 -2508 -5979
rect -2474 -6013 -2416 -5979
rect -2382 -6013 -2324 -5979
rect -2290 -6013 -2232 -5979
rect -2198 -6013 -2140 -5979
rect -2106 -6013 -2048 -5979
rect -2014 -6013 -1956 -5979
rect -1922 -6013 -1864 -5979
rect -1830 -6013 -1772 -5979
rect -1738 -6013 -1680 -5979
rect -1646 -6013 -1588 -5979
rect -1554 -6013 -1496 -5979
rect -1462 -6013 -1404 -5979
rect -1370 -6013 -1312 -5979
rect -1278 -6013 -1220 -5979
rect -1186 -6013 -1128 -5979
rect -1094 -6013 -1036 -5979
rect -1002 -6013 -944 -5979
rect -910 -6013 -852 -5979
rect -818 -6013 -760 -5979
rect -726 -6013 -668 -5979
rect -634 -6013 -576 -5979
rect -542 -6013 -484 -5979
rect -450 -6013 -392 -5979
rect -358 -6013 -300 -5979
rect -266 -6013 -208 -5979
rect -174 -6013 -116 -5979
rect -82 -6013 -24 -5979
rect 10 -6013 68 -5979
rect 102 -6013 160 -5979
rect 194 -6013 252 -5979
rect 286 -6013 344 -5979
rect 378 -6013 436 -5979
rect 470 -6013 528 -5979
rect 562 -6013 620 -5979
rect 654 -6013 712 -5979
rect 746 -6013 804 -5979
rect 838 -6013 896 -5979
rect 930 -6013 988 -5979
rect 1022 -6013 1080 -5979
rect 1114 -6013 1172 -5979
rect 1206 -6013 1264 -5979
rect 1298 -6013 1356 -5979
rect 1390 -6013 1448 -5979
rect 1482 -6013 1540 -5979
rect 1574 -6013 1632 -5979
rect 1666 -6013 1724 -5979
rect 1758 -6013 1816 -5979
rect 1850 -6013 1908 -5979
rect 1942 -6013 2000 -5979
rect 2034 -6013 2092 -5979
rect 2126 -6013 2184 -5979
rect 2218 -6013 2276 -5979
rect 2310 -6013 2368 -5979
rect 2402 -6013 2460 -5979
rect 2494 -6013 2552 -5979
rect 2586 -6013 2644 -5979
rect 2678 -6013 2736 -5979
rect 2770 -6013 2828 -5979
rect 2862 -6013 2920 -5979
rect 2954 -6013 3012 -5979
rect 3046 -6013 3104 -5979
rect 3138 -6013 3196 -5979
rect 3230 -6013 3288 -5979
rect 3322 -6013 3380 -5979
rect 3414 -6013 3472 -5979
rect 3506 -6013 3564 -5979
rect 3598 -6013 3656 -5979
rect 3690 -6013 3748 -5979
rect 3782 -6013 3840 -5979
rect 3874 -6013 3932 -5979
rect 3966 -6013 4024 -5979
rect 4058 -6013 4116 -5979
rect 4150 -6013 4208 -5979
rect 4242 -6013 4300 -5979
rect 4334 -6013 4392 -5979
rect 4426 -6013 4484 -5979
rect 4518 -6013 4576 -5979
rect 4610 -6013 4668 -5979
rect 4702 -6013 4760 -5979
rect 4794 -6013 4852 -5979
rect 4886 -6013 4944 -5979
rect 4978 -6013 5036 -5979
rect 5070 -6013 5128 -5979
rect 5162 -6013 5220 -5979
rect 5254 -6013 5312 -5979
rect 5346 -6013 5404 -5979
rect 5438 -6013 5496 -5979
rect 5530 -6013 5588 -5979
rect 5622 -6013 5680 -5979
rect 5714 -6013 5772 -5979
rect 5806 -6013 5864 -5979
rect 5898 -6013 5956 -5979
rect 5990 -6013 6048 -5979
rect 6082 -6013 6140 -5979
rect 6174 -6013 6232 -5979
rect 6266 -6013 6324 -5979
rect 6358 -6013 6416 -5979
rect 6450 -6013 6508 -5979
rect 6542 -6013 6600 -5979
rect 6634 -6013 6692 -5979
rect 6726 -6013 6784 -5979
rect 6818 -6013 6876 -5979
rect 6910 -6013 6968 -5979
rect 7002 -6013 7060 -5979
rect 7094 -6013 7152 -5979
rect 7186 -6013 7244 -5979
rect 7278 -6013 7336 -5979
rect 7370 -6013 7428 -5979
rect 7462 -6013 7520 -5979
rect 7554 -6013 7612 -5979
rect 7646 -6013 7704 -5979
rect 7738 -6013 7796 -5979
rect 7830 -6013 7888 -5979
rect 7922 -6013 7980 -5979
rect 8014 -6013 8072 -5979
rect 8106 -6013 8164 -5979
rect 8198 -6013 8256 -5979
rect 8290 -6013 8348 -5979
rect 8382 -6013 8440 -5979
rect 8474 -6013 8532 -5979
rect 8566 -6013 8624 -5979
rect 8658 -6013 8716 -5979
rect 8750 -6013 8808 -5979
rect 8842 -6013 8900 -5979
rect 8934 -6013 8992 -5979
rect 9026 -6013 9084 -5979
rect 9118 -6013 9176 -5979
rect 9210 -6013 9268 -5979
rect 9302 -6013 9360 -5979
rect 9394 -6013 9452 -5979
rect 9486 -6013 9544 -5979
rect 9578 -6013 9636 -5979
rect 9670 -6013 9728 -5979
rect 9762 -6013 9820 -5979
rect 9854 -6013 9912 -5979
rect 9946 -6013 10004 -5979
rect 10038 -6013 10096 -5979
rect 10130 -6013 10188 -5979
rect 10222 -6013 10280 -5979
rect 10314 -6013 10372 -5979
rect 10406 -6013 10464 -5979
rect 10498 -6013 10556 -5979
rect 10590 -6013 10648 -5979
rect 10682 -6013 10740 -5979
rect 10774 -6013 10832 -5979
rect 10866 -6013 10924 -5979
rect 10958 -6013 11016 -5979
rect 11050 -6013 11108 -5979
rect 11142 -6013 11200 -5979
rect 11234 -6013 11292 -5979
rect 11326 -6013 11384 -5979
rect 11418 -6013 11476 -5979
rect 11510 -6013 11568 -5979
rect 11602 -6013 11660 -5979
rect 11694 -6013 11752 -5979
rect 11786 -6013 11844 -5979
rect 11878 -6013 11936 -5979
rect 11970 -6013 12028 -5979
rect 12062 -6013 12120 -5979
rect 12154 -6013 12212 -5979
rect 12246 -6013 12304 -5979
rect 12338 -6013 12396 -5979
rect 12430 -6013 12488 -5979
rect 12522 -6013 12580 -5979
rect 12614 -6013 12672 -5979
rect 12706 -6013 12764 -5979
rect 12798 -6013 12856 -5979
rect 12890 -6013 12948 -5979
rect 12982 -6013 13040 -5979
rect 13074 -6013 13132 -5979
rect 13166 -6013 13224 -5979
rect 13258 -6013 13316 -5979
rect 13350 -6013 13408 -5979
rect 13442 -6013 13500 -5979
rect 13534 -6013 13592 -5979
rect 13626 -6013 13684 -5979
rect 13718 -6013 13776 -5979
rect 13810 -6013 13868 -5979
rect 13902 -6013 13960 -5979
rect 13994 -6013 14052 -5979
rect 14086 -6013 14144 -5979
rect 14178 -6013 14236 -5979
rect 14270 -6013 14328 -5979
rect 14362 -6013 14420 -5979
rect 14454 -6013 14512 -5979
rect 14546 -6013 14604 -5979
rect 14638 -6013 14696 -5979
rect 14730 -6013 14788 -5979
rect 14822 -6013 14880 -5979
rect 14914 -6013 14972 -5979
rect 15006 -6013 15064 -5979
rect 15098 -6013 15156 -5979
rect 15190 -6013 15248 -5979
rect 15282 -6013 15340 -5979
rect 15374 -6013 15432 -5979
rect 15466 -6013 15524 -5979
rect 15558 -6013 15616 -5979
rect 15650 -6013 15708 -5979
rect 15742 -6013 15800 -5979
rect 15834 -6013 15892 -5979
rect 15926 -6013 15984 -5979
rect 16018 -6013 16076 -5979
rect 16110 -6013 16168 -5979
rect 16202 -6013 16260 -5979
rect 16294 -6013 16352 -5979
rect 16386 -6013 16444 -5979
rect 16478 -6013 16536 -5979
rect 16570 -6013 16628 -5979
rect 16662 -6013 16691 -5979
rect -2980 -6074 -2278 -6013
rect -2980 -6108 -2962 -6074
rect -2928 -6108 -2330 -6074
rect -2296 -6108 -2278 -6074
rect -2980 -6167 -2278 -6108
rect -2244 -6107 -2186 -6013
rect -2244 -6141 -2232 -6107
rect -2198 -6141 -2186 -6107
rect -2244 -6158 -2186 -6141
rect -1416 -6081 -1082 -6013
rect -1416 -6115 -1398 -6081
rect -1364 -6115 -1134 -6081
rect -1100 -6115 -1082 -6081
rect -2980 -6235 -2902 -6201
rect -2868 -6235 -2799 -6201
rect -2765 -6235 -2696 -6201
rect -2662 -6235 -2642 -6201
rect -2980 -6305 -2642 -6235
rect -2608 -6237 -2278 -6167
rect -2608 -6271 -2588 -6237
rect -2554 -6271 -2489 -6237
rect -2455 -6271 -2390 -6237
rect -2356 -6271 -2278 -6237
rect -1416 -6167 -1082 -6115
rect -1048 -6107 -990 -6013
rect -1048 -6141 -1036 -6107
rect -1002 -6141 -990 -6107
rect -1048 -6158 -990 -6141
rect -956 -6055 -894 -6013
rect -956 -6089 -934 -6055
rect -900 -6089 -894 -6055
rect -956 -6123 -894 -6089
rect -956 -6157 -934 -6123
rect -900 -6157 -894 -6123
rect -1416 -6237 -1266 -6167
rect -956 -6173 -894 -6157
rect -853 -6055 -714 -6047
rect -853 -6089 -766 -6055
rect -732 -6089 -714 -6055
rect -853 -6106 -714 -6089
rect -853 -6140 -848 -6106
rect -814 -6140 -769 -6106
rect -735 -6123 -714 -6106
rect -853 -6157 -766 -6140
rect -732 -6157 -714 -6123
rect -853 -6173 -714 -6157
rect -680 -6107 -622 -6013
rect -680 -6141 -668 -6107
rect -634 -6141 -622 -6107
rect -680 -6158 -622 -6141
rect -588 -6081 -254 -6013
rect -588 -6115 -570 -6081
rect -536 -6115 -306 -6081
rect -272 -6115 -254 -6081
rect -588 -6167 -254 -6115
rect -220 -6107 -162 -6013
rect -32 -6057 27 -6013
rect -32 -6091 -16 -6057
rect 18 -6091 27 -6057
rect -32 -6107 27 -6091
rect 61 -6068 113 -6052
rect 61 -6102 70 -6068
rect 104 -6102 113 -6068
rect -220 -6141 -208 -6107
rect -174 -6141 -162 -6107
rect 61 -6141 113 -6102
rect 147 -6057 199 -6013
rect 147 -6091 156 -6057
rect 190 -6091 199 -6057
rect 147 -6107 199 -6091
rect 233 -6068 284 -6052
rect 233 -6102 242 -6068
rect 276 -6102 284 -6068
rect 233 -6141 284 -6102
rect 318 -6057 378 -6013
rect 318 -6091 328 -6057
rect 362 -6091 378 -6057
rect 318 -6107 378 -6091
rect 516 -6107 574 -6013
rect 516 -6141 528 -6107
rect 562 -6141 574 -6107
rect -220 -6158 -162 -6141
rect -1416 -6271 -1396 -6237
rect -1362 -6271 -1266 -6237
rect -1232 -6235 -1136 -6201
rect -1102 -6235 -1082 -6201
rect -2980 -6345 -2278 -6305
rect -2980 -6379 -2962 -6345
rect -2928 -6379 -2330 -6345
rect -2296 -6379 -2278 -6345
rect -2980 -6447 -2278 -6379
rect -2980 -6481 -2962 -6447
rect -2928 -6481 -2330 -6447
rect -2296 -6481 -2278 -6447
rect -2980 -6523 -2278 -6481
rect -2244 -6325 -2186 -6290
rect -1232 -6305 -1082 -6235
rect -954 -6211 -887 -6207
rect -954 -6245 -937 -6211
rect -903 -6218 -887 -6211
rect -954 -6252 -932 -6245
rect -898 -6252 -887 -6218
rect -954 -6261 -887 -6252
rect -2244 -6359 -2232 -6325
rect -2198 -6359 -2186 -6325
rect -2244 -6418 -2186 -6359
rect -2244 -6452 -2232 -6418
rect -2198 -6452 -2186 -6418
rect -2244 -6523 -2186 -6452
rect -1416 -6345 -1082 -6305
rect -1416 -6379 -1398 -6345
rect -1364 -6379 -1134 -6345
rect -1100 -6379 -1082 -6345
rect -1416 -6447 -1082 -6379
rect -1416 -6481 -1398 -6447
rect -1364 -6481 -1134 -6447
rect -1100 -6481 -1082 -6447
rect -1416 -6523 -1082 -6481
rect -1048 -6325 -990 -6290
rect -853 -6293 -819 -6173
rect -785 -6245 -769 -6211
rect -735 -6217 -718 -6211
rect -785 -6251 -760 -6245
rect -726 -6251 -718 -6217
rect -785 -6261 -718 -6251
rect -588 -6237 -438 -6167
rect -124 -6173 482 -6141
rect 516 -6158 574 -6141
rect 608 -6081 942 -6013
rect 608 -6115 626 -6081
rect 660 -6115 890 -6081
rect 924 -6115 942 -6081
rect -124 -6175 434 -6173
rect -588 -6271 -568 -6237
rect -534 -6271 -438 -6237
rect -404 -6235 -308 -6201
rect -274 -6235 -254 -6201
rect -1048 -6359 -1036 -6325
rect -1002 -6359 -990 -6325
rect -1048 -6418 -990 -6359
rect -1048 -6452 -1036 -6418
rect -1002 -6452 -990 -6418
rect -1048 -6523 -990 -6452
rect -956 -6311 -900 -6295
rect -956 -6345 -934 -6311
rect -956 -6379 -900 -6345
rect -956 -6413 -934 -6379
rect -956 -6447 -900 -6413
rect -956 -6481 -934 -6447
rect -956 -6523 -900 -6481
rect -866 -6311 -800 -6293
rect -866 -6345 -850 -6311
rect -816 -6345 -800 -6311
rect -866 -6379 -800 -6345
rect -866 -6413 -850 -6379
rect -816 -6413 -800 -6379
rect -866 -6447 -800 -6413
rect -866 -6481 -850 -6447
rect -816 -6481 -800 -6447
rect -866 -6489 -800 -6481
rect -766 -6311 -714 -6295
rect -732 -6345 -714 -6311
rect -766 -6379 -714 -6345
rect -732 -6413 -714 -6379
rect -766 -6447 -714 -6413
rect -732 -6481 -714 -6447
rect -766 -6523 -714 -6481
rect -680 -6325 -622 -6290
rect -404 -6305 -254 -6235
rect -124 -6288 -90 -6175
rect 422 -6207 434 -6175
rect 468 -6207 482 -6173
rect -56 -6211 387 -6209
rect -56 -6245 -30 -6211
rect 4 -6245 38 -6211
rect 72 -6245 106 -6211
rect 140 -6245 174 -6211
rect 208 -6245 242 -6211
rect 276 -6245 310 -6211
rect 344 -6245 387 -6211
rect -56 -6254 387 -6245
rect 422 -6288 482 -6207
rect 608 -6167 942 -6115
rect 976 -6107 1034 -6013
rect 1154 -6066 1219 -6047
rect 976 -6141 988 -6107
rect 1022 -6141 1034 -6107
rect 976 -6158 1034 -6141
rect 1068 -6133 1116 -6071
rect 1068 -6167 1076 -6133
rect 1110 -6167 1116 -6133
rect 608 -6237 758 -6167
rect 608 -6271 628 -6237
rect 662 -6271 758 -6237
rect 792 -6235 888 -6201
rect 922 -6235 942 -6201
rect -680 -6359 -668 -6325
rect -634 -6359 -622 -6325
rect -680 -6418 -622 -6359
rect -680 -6452 -668 -6418
rect -634 -6452 -622 -6418
rect -680 -6523 -622 -6452
rect -588 -6345 -254 -6305
rect -588 -6379 -570 -6345
rect -536 -6379 -306 -6345
rect -272 -6379 -254 -6345
rect -588 -6447 -254 -6379
rect -588 -6481 -570 -6447
rect -536 -6481 -306 -6447
rect -272 -6481 -254 -6447
rect -588 -6523 -254 -6481
rect -220 -6325 -162 -6290
rect -124 -6322 482 -6288
rect -220 -6359 -208 -6325
rect -174 -6359 -162 -6325
rect -24 -6345 27 -6322
rect -220 -6418 -162 -6359
rect -220 -6452 -208 -6418
rect -174 -6452 -162 -6418
rect -220 -6523 -162 -6452
rect -128 -6372 -59 -6356
rect -128 -6406 -102 -6372
rect -68 -6406 -59 -6372
rect -128 -6440 -59 -6406
rect -128 -6474 -102 -6440
rect -68 -6474 -59 -6440
rect -128 -6523 -59 -6474
rect -24 -6379 -16 -6345
rect 18 -6379 27 -6345
rect 148 -6345 199 -6322
rect -24 -6433 27 -6379
rect -24 -6467 -16 -6433
rect 18 -6467 27 -6433
rect -24 -6483 27 -6467
rect 61 -6372 113 -6356
rect 61 -6406 70 -6372
rect 104 -6406 113 -6372
rect 61 -6440 113 -6406
rect 61 -6474 70 -6440
rect 104 -6474 113 -6440
rect 61 -6523 113 -6474
rect 148 -6379 156 -6345
rect 190 -6379 199 -6345
rect 319 -6345 371 -6322
rect 148 -6433 199 -6379
rect 148 -6467 156 -6433
rect 190 -6467 199 -6433
rect 148 -6483 199 -6467
rect 233 -6372 285 -6356
rect 233 -6406 242 -6372
rect 276 -6406 285 -6372
rect 233 -6440 285 -6406
rect 233 -6474 242 -6440
rect 276 -6474 285 -6440
rect 233 -6523 285 -6474
rect 319 -6379 328 -6345
rect 362 -6379 371 -6345
rect 516 -6325 574 -6290
rect 792 -6305 942 -6235
rect 1068 -6206 1116 -6167
rect 1068 -6240 1076 -6206
rect 1110 -6211 1116 -6206
rect 1068 -6245 1082 -6240
rect 1068 -6261 1116 -6245
rect 1154 -6100 1169 -6066
rect 1203 -6100 1219 -6066
rect 1154 -6148 1219 -6100
rect 1253 -6064 1310 -6013
rect 1287 -6098 1310 -6064
rect 1253 -6114 1310 -6098
rect 1344 -6107 1402 -6013
rect 1344 -6141 1356 -6107
rect 1390 -6141 1402 -6107
rect 1154 -6212 1310 -6148
rect 1344 -6158 1402 -6141
rect 1436 -6081 1770 -6013
rect 1436 -6115 1454 -6081
rect 1488 -6115 1718 -6081
rect 1752 -6115 1770 -6081
rect 1154 -6246 1171 -6212
rect 1205 -6246 1263 -6212
rect 1297 -6246 1310 -6212
rect 1154 -6254 1310 -6246
rect 1436 -6167 1770 -6115
rect 1804 -6107 1862 -6013
rect 1804 -6141 1816 -6107
rect 1850 -6141 1862 -6107
rect 1804 -6158 1862 -6141
rect 1896 -6081 2230 -6013
rect 1896 -6115 1914 -6081
rect 1948 -6115 2178 -6081
rect 2212 -6115 2230 -6081
rect 1896 -6167 2230 -6115
rect 2264 -6107 2322 -6013
rect 2264 -6141 2276 -6107
rect 2310 -6141 2322 -6107
rect 2264 -6158 2322 -6141
rect 2356 -6066 2422 -6047
rect 2356 -6100 2375 -6066
rect 2409 -6100 2422 -6066
rect 2356 -6143 2422 -6100
rect 2456 -6066 2522 -6013
rect 2456 -6100 2472 -6066
rect 2506 -6100 2522 -6066
rect 2456 -6109 2522 -6100
rect 2615 -6066 2685 -6047
rect 2615 -6100 2632 -6066
rect 2666 -6100 2685 -6066
rect 1436 -6237 1586 -6167
rect 319 -6433 371 -6379
rect 319 -6467 328 -6433
rect 362 -6467 371 -6433
rect 319 -6483 371 -6467
rect 405 -6372 482 -6356
rect 405 -6406 414 -6372
rect 448 -6406 482 -6372
rect 405 -6440 482 -6406
rect 405 -6474 414 -6440
rect 448 -6474 482 -6440
rect 405 -6523 482 -6474
rect 516 -6359 528 -6325
rect 562 -6359 574 -6325
rect 516 -6418 574 -6359
rect 516 -6452 528 -6418
rect 562 -6452 574 -6418
rect 516 -6523 574 -6452
rect 608 -6345 942 -6305
rect 608 -6379 626 -6345
rect 660 -6379 890 -6345
rect 924 -6379 942 -6345
rect 608 -6447 942 -6379
rect 608 -6481 626 -6447
rect 660 -6481 890 -6447
rect 924 -6481 942 -6447
rect 608 -6523 942 -6481
rect 976 -6325 1034 -6290
rect 976 -6359 988 -6325
rect 1022 -6359 1034 -6325
rect 976 -6418 1034 -6359
rect 976 -6452 988 -6418
rect 1022 -6452 1034 -6418
rect 976 -6523 1034 -6452
rect 1068 -6345 1120 -6329
rect 1068 -6379 1086 -6345
rect 1068 -6447 1120 -6379
rect 1068 -6481 1086 -6447
rect 1068 -6523 1120 -6481
rect 1154 -6345 1220 -6254
rect 1436 -6271 1456 -6237
rect 1490 -6271 1586 -6237
rect 1620 -6235 1716 -6201
rect 1750 -6235 1770 -6201
rect 1344 -6325 1402 -6290
rect 1620 -6305 1770 -6235
rect 1896 -6237 2046 -6167
rect 2356 -6177 2550 -6143
rect 2480 -6201 2550 -6177
rect 1896 -6271 1916 -6237
rect 1950 -6271 2046 -6237
rect 2080 -6235 2176 -6201
rect 2210 -6235 2230 -6201
rect 2480 -6211 2566 -6201
rect 1154 -6379 1170 -6345
rect 1204 -6379 1220 -6345
rect 1154 -6447 1220 -6379
rect 1154 -6481 1170 -6447
rect 1204 -6481 1220 -6447
rect 1154 -6489 1220 -6481
rect 1254 -6345 1310 -6329
rect 1288 -6379 1310 -6345
rect 1254 -6447 1310 -6379
rect 1288 -6481 1310 -6447
rect 1254 -6523 1310 -6481
rect 1344 -6359 1356 -6325
rect 1390 -6359 1402 -6325
rect 1344 -6418 1402 -6359
rect 1344 -6452 1356 -6418
rect 1390 -6452 1402 -6418
rect 1344 -6523 1402 -6452
rect 1436 -6345 1770 -6305
rect 1436 -6379 1454 -6345
rect 1488 -6379 1718 -6345
rect 1752 -6379 1770 -6345
rect 1436 -6447 1770 -6379
rect 1436 -6481 1454 -6447
rect 1488 -6481 1718 -6447
rect 1752 -6481 1770 -6447
rect 1436 -6523 1770 -6481
rect 1804 -6325 1862 -6290
rect 2080 -6305 2230 -6235
rect 2356 -6217 2396 -6211
rect 2356 -6251 2369 -6217
rect 2430 -6245 2446 -6211
rect 2403 -6251 2446 -6245
rect 2356 -6254 2446 -6251
rect 2480 -6245 2516 -6211
rect 2550 -6245 2566 -6211
rect 2480 -6259 2566 -6245
rect 2615 -6210 2685 -6100
rect 2737 -6066 2787 -6047
rect 2771 -6100 2787 -6066
rect 2737 -6142 2787 -6100
rect 2877 -6066 2943 -6013
rect 2877 -6100 2893 -6066
rect 2927 -6100 2943 -6066
rect 2877 -6116 2943 -6100
rect 2977 -6066 3058 -6047
rect 2977 -6100 2991 -6066
rect 3025 -6100 3058 -6066
rect 2977 -6124 3058 -6100
rect 2737 -6176 2855 -6142
rect 2821 -6195 2855 -6176
rect 2615 -6211 2787 -6210
rect 2615 -6245 2737 -6211
rect 2771 -6245 2787 -6211
rect 2480 -6288 2550 -6259
rect 1804 -6359 1816 -6325
rect 1850 -6359 1862 -6325
rect 1804 -6418 1862 -6359
rect 1804 -6452 1816 -6418
rect 1850 -6452 1862 -6418
rect 1804 -6523 1862 -6452
rect 1896 -6345 2230 -6305
rect 1896 -6379 1914 -6345
rect 1948 -6379 2178 -6345
rect 2212 -6379 2230 -6345
rect 1896 -6447 2230 -6379
rect 1896 -6481 1914 -6447
rect 1948 -6481 2178 -6447
rect 2212 -6481 2230 -6447
rect 1896 -6523 2230 -6481
rect 2264 -6325 2322 -6290
rect 2264 -6359 2276 -6325
rect 2310 -6359 2322 -6325
rect 2264 -6418 2322 -6359
rect 2264 -6452 2276 -6418
rect 2310 -6452 2322 -6418
rect 2264 -6523 2322 -6452
rect 2356 -6322 2550 -6288
rect 2615 -6260 2787 -6245
rect 2821 -6211 2974 -6195
rect 2821 -6245 2937 -6211
rect 2971 -6245 2974 -6211
rect 2356 -6372 2425 -6322
rect 2356 -6406 2375 -6372
rect 2409 -6406 2425 -6372
rect 2356 -6440 2425 -6406
rect 2356 -6474 2375 -6440
rect 2409 -6474 2425 -6440
rect 2356 -6489 2425 -6474
rect 2459 -6372 2525 -6356
rect 2459 -6406 2475 -6372
rect 2509 -6406 2525 -6372
rect 2459 -6440 2525 -6406
rect 2459 -6474 2475 -6440
rect 2509 -6474 2525 -6440
rect 2459 -6523 2525 -6474
rect 2615 -6372 2685 -6260
rect 2821 -6261 2974 -6245
rect 3008 -6216 3058 -6124
rect 3092 -6107 3150 -6013
rect 3092 -6141 3104 -6107
rect 3138 -6141 3150 -6107
rect 3092 -6158 3150 -6141
rect 3184 -6081 3518 -6013
rect 3184 -6115 3202 -6081
rect 3236 -6115 3466 -6081
rect 3500 -6115 3518 -6081
rect 3008 -6250 3015 -6216
rect 3049 -6250 3058 -6216
rect 2821 -6295 2855 -6261
rect 2615 -6406 2633 -6372
rect 2667 -6406 2685 -6372
rect 2615 -6440 2685 -6406
rect 2615 -6474 2633 -6440
rect 2667 -6474 2685 -6440
rect 2615 -6489 2685 -6474
rect 2737 -6329 2855 -6295
rect 2737 -6371 2787 -6329
rect 3008 -6334 3058 -6250
rect 3184 -6167 3518 -6115
rect 3552 -6107 3610 -6013
rect 3552 -6141 3564 -6107
rect 3598 -6141 3610 -6107
rect 3552 -6158 3610 -6141
rect 4380 -6074 5449 -6013
rect 4380 -6108 4398 -6074
rect 4432 -6108 5398 -6074
rect 5432 -6108 5449 -6074
rect 4380 -6167 5449 -6108
rect 6312 -6107 6370 -6013
rect 6312 -6141 6324 -6107
rect 6358 -6141 6370 -6107
rect 6312 -6158 6370 -6141
rect 6404 -6081 6738 -6013
rect 6404 -6115 6422 -6081
rect 6456 -6115 6686 -6081
rect 6720 -6115 6738 -6081
rect 6404 -6167 6738 -6115
rect 6772 -6107 6830 -6013
rect 6772 -6141 6784 -6107
rect 6818 -6141 6830 -6107
rect 6772 -6158 6830 -6141
rect 6864 -6066 6930 -6047
rect 6864 -6100 6883 -6066
rect 6917 -6100 6930 -6066
rect 6864 -6143 6930 -6100
rect 6964 -6066 7030 -6013
rect 6964 -6100 6980 -6066
rect 7014 -6100 7030 -6066
rect 6964 -6109 7030 -6100
rect 7123 -6066 7193 -6047
rect 7123 -6100 7140 -6066
rect 7174 -6100 7193 -6066
rect 3184 -6237 3334 -6167
rect 3184 -6271 3204 -6237
rect 3238 -6271 3334 -6237
rect 3368 -6235 3464 -6201
rect 3498 -6235 3518 -6201
rect 2771 -6405 2787 -6371
rect 2737 -6439 2787 -6405
rect 2771 -6473 2787 -6439
rect 2737 -6489 2787 -6473
rect 2877 -6372 2943 -6363
rect 2877 -6406 2893 -6372
rect 2927 -6406 2943 -6372
rect 2877 -6440 2943 -6406
rect 2877 -6474 2893 -6440
rect 2927 -6474 2943 -6440
rect 2877 -6523 2943 -6474
rect 2977 -6371 3058 -6334
rect 2977 -6405 2991 -6371
rect 3025 -6405 3058 -6371
rect 2977 -6439 3058 -6405
rect 2977 -6473 2991 -6439
rect 3025 -6473 3058 -6439
rect 2977 -6489 3058 -6473
rect 3092 -6325 3150 -6290
rect 3368 -6305 3518 -6235
rect 4380 -6237 4896 -6167
rect 4380 -6271 4458 -6237
rect 4492 -6271 4586 -6237
rect 4620 -6271 4714 -6237
rect 4748 -6271 4842 -6237
rect 4876 -6271 4896 -6237
rect 4930 -6235 4950 -6201
rect 4984 -6235 5078 -6201
rect 5112 -6235 5206 -6201
rect 5240 -6235 5334 -6201
rect 5368 -6235 5449 -6201
rect 3092 -6359 3104 -6325
rect 3138 -6359 3150 -6325
rect 3092 -6418 3150 -6359
rect 3092 -6452 3104 -6418
rect 3138 -6452 3150 -6418
rect 3092 -6523 3150 -6452
rect 3184 -6345 3518 -6305
rect 3184 -6379 3202 -6345
rect 3236 -6379 3466 -6345
rect 3500 -6379 3518 -6345
rect 3184 -6447 3518 -6379
rect 3184 -6481 3202 -6447
rect 3236 -6481 3466 -6447
rect 3500 -6481 3518 -6447
rect 3184 -6523 3518 -6481
rect 3552 -6325 3610 -6290
rect 4930 -6305 5449 -6235
rect 6404 -6237 6554 -6167
rect 6864 -6177 7058 -6143
rect 6988 -6201 7058 -6177
rect 6404 -6271 6424 -6237
rect 6458 -6271 6554 -6237
rect 6588 -6235 6684 -6201
rect 6718 -6235 6738 -6201
rect 6988 -6211 7074 -6201
rect 3552 -6359 3564 -6325
rect 3598 -6359 3610 -6325
rect 3552 -6418 3610 -6359
rect 3552 -6452 3564 -6418
rect 3598 -6452 3610 -6418
rect 3552 -6523 3610 -6452
rect 4380 -6345 5449 -6305
rect 4380 -6379 4398 -6345
rect 4432 -6379 5398 -6345
rect 5432 -6379 5449 -6345
rect 4380 -6447 5449 -6379
rect 4380 -6481 4398 -6447
rect 4432 -6481 5398 -6447
rect 5432 -6481 5449 -6447
rect 4380 -6523 5449 -6481
rect 6312 -6325 6370 -6290
rect 6588 -6305 6738 -6235
rect 6864 -6216 6904 -6211
rect 6864 -6250 6876 -6216
rect 6938 -6245 6954 -6211
rect 6910 -6250 6954 -6245
rect 6864 -6254 6954 -6250
rect 6988 -6245 7024 -6211
rect 7058 -6245 7074 -6211
rect 6988 -6259 7074 -6245
rect 7123 -6210 7193 -6100
rect 7245 -6066 7295 -6047
rect 7279 -6100 7295 -6066
rect 7245 -6142 7295 -6100
rect 7385 -6066 7451 -6013
rect 7385 -6100 7401 -6066
rect 7435 -6100 7451 -6066
rect 7385 -6116 7451 -6100
rect 7485 -6066 7566 -6047
rect 7485 -6100 7499 -6066
rect 7533 -6100 7566 -6066
rect 7485 -6124 7566 -6100
rect 7245 -6176 7363 -6142
rect 7329 -6195 7363 -6176
rect 7123 -6211 7295 -6210
rect 7123 -6245 7245 -6211
rect 7279 -6245 7295 -6211
rect 6988 -6288 7058 -6259
rect 6312 -6359 6324 -6325
rect 6358 -6359 6370 -6325
rect 6312 -6418 6370 -6359
rect 6312 -6452 6324 -6418
rect 6358 -6452 6370 -6418
rect 6312 -6523 6370 -6452
rect 6404 -6345 6738 -6305
rect 6404 -6379 6422 -6345
rect 6456 -6379 6686 -6345
rect 6720 -6379 6738 -6345
rect 6404 -6447 6738 -6379
rect 6404 -6481 6422 -6447
rect 6456 -6481 6686 -6447
rect 6720 -6481 6738 -6447
rect 6404 -6523 6738 -6481
rect 6772 -6325 6830 -6290
rect 6772 -6359 6784 -6325
rect 6818 -6359 6830 -6325
rect 6772 -6418 6830 -6359
rect 6772 -6452 6784 -6418
rect 6818 -6452 6830 -6418
rect 6772 -6523 6830 -6452
rect 6864 -6322 7058 -6288
rect 7123 -6260 7295 -6245
rect 7329 -6211 7482 -6195
rect 7329 -6245 7445 -6211
rect 7479 -6245 7482 -6211
rect 6864 -6372 6933 -6322
rect 6864 -6406 6883 -6372
rect 6917 -6406 6933 -6372
rect 6864 -6440 6933 -6406
rect 6864 -6474 6883 -6440
rect 6917 -6474 6933 -6440
rect 6864 -6489 6933 -6474
rect 6967 -6372 7033 -6356
rect 6967 -6406 6983 -6372
rect 7017 -6406 7033 -6372
rect 6967 -6440 7033 -6406
rect 6967 -6474 6983 -6440
rect 7017 -6474 7033 -6440
rect 6967 -6523 7033 -6474
rect 7123 -6372 7193 -6260
rect 7329 -6261 7482 -6245
rect 7516 -6216 7566 -6124
rect 7600 -6107 7658 -6013
rect 7600 -6141 7612 -6107
rect 7646 -6141 7658 -6107
rect 7600 -6158 7658 -6141
rect 7692 -6081 8026 -6013
rect 7692 -6115 7710 -6081
rect 7744 -6115 7974 -6081
rect 8008 -6115 8026 -6081
rect 7516 -6250 7522 -6216
rect 7556 -6250 7566 -6216
rect 7329 -6295 7363 -6261
rect 7123 -6406 7141 -6372
rect 7175 -6406 7193 -6372
rect 7123 -6440 7193 -6406
rect 7123 -6474 7141 -6440
rect 7175 -6474 7193 -6440
rect 7123 -6489 7193 -6474
rect 7245 -6329 7363 -6295
rect 7245 -6371 7295 -6329
rect 7516 -6334 7566 -6250
rect 7692 -6167 8026 -6115
rect 8060 -6107 8118 -6013
rect 8060 -6141 8072 -6107
rect 8106 -6141 8118 -6107
rect 8060 -6158 8118 -6141
rect 8152 -6066 8218 -6047
rect 8152 -6100 8171 -6066
rect 8205 -6100 8218 -6066
rect 8152 -6143 8218 -6100
rect 8252 -6066 8318 -6013
rect 8252 -6100 8268 -6066
rect 8302 -6100 8318 -6066
rect 8252 -6109 8318 -6100
rect 8411 -6066 8481 -6047
rect 8411 -6100 8428 -6066
rect 8462 -6100 8481 -6066
rect 7692 -6237 7842 -6167
rect 8152 -6177 8346 -6143
rect 8276 -6201 8346 -6177
rect 7692 -6271 7712 -6237
rect 7746 -6271 7842 -6237
rect 7876 -6235 7972 -6201
rect 8006 -6235 8026 -6201
rect 8276 -6211 8362 -6201
rect 7279 -6405 7295 -6371
rect 7245 -6439 7295 -6405
rect 7279 -6473 7295 -6439
rect 7245 -6489 7295 -6473
rect 7385 -6372 7451 -6363
rect 7385 -6406 7401 -6372
rect 7435 -6406 7451 -6372
rect 7385 -6440 7451 -6406
rect 7385 -6474 7401 -6440
rect 7435 -6474 7451 -6440
rect 7385 -6523 7451 -6474
rect 7485 -6371 7566 -6334
rect 7485 -6405 7499 -6371
rect 7533 -6405 7566 -6371
rect 7485 -6439 7566 -6405
rect 7485 -6473 7499 -6439
rect 7533 -6473 7566 -6439
rect 7485 -6489 7566 -6473
rect 7600 -6325 7658 -6290
rect 7876 -6305 8026 -6235
rect 8152 -6215 8192 -6211
rect 8152 -6249 8164 -6215
rect 8226 -6245 8242 -6211
rect 8198 -6249 8242 -6245
rect 8152 -6254 8242 -6249
rect 8276 -6245 8312 -6211
rect 8346 -6245 8362 -6211
rect 8276 -6259 8362 -6245
rect 8411 -6210 8481 -6100
rect 8533 -6066 8583 -6047
rect 8567 -6100 8583 -6066
rect 8533 -6142 8583 -6100
rect 8673 -6066 8739 -6013
rect 8673 -6100 8689 -6066
rect 8723 -6100 8739 -6066
rect 8673 -6116 8739 -6100
rect 8773 -6066 8854 -6047
rect 8773 -6100 8787 -6066
rect 8821 -6100 8854 -6066
rect 8773 -6124 8854 -6100
rect 8533 -6176 8651 -6142
rect 8617 -6195 8651 -6176
rect 8411 -6211 8583 -6210
rect 8411 -6245 8533 -6211
rect 8567 -6245 8583 -6211
rect 8276 -6288 8346 -6259
rect 7600 -6359 7612 -6325
rect 7646 -6359 7658 -6325
rect 7600 -6418 7658 -6359
rect 7600 -6452 7612 -6418
rect 7646 -6452 7658 -6418
rect 7600 -6523 7658 -6452
rect 7692 -6345 8026 -6305
rect 7692 -6379 7710 -6345
rect 7744 -6379 7974 -6345
rect 8008 -6379 8026 -6345
rect 7692 -6447 8026 -6379
rect 7692 -6481 7710 -6447
rect 7744 -6481 7974 -6447
rect 8008 -6481 8026 -6447
rect 7692 -6523 8026 -6481
rect 8060 -6325 8118 -6290
rect 8060 -6359 8072 -6325
rect 8106 -6359 8118 -6325
rect 8060 -6418 8118 -6359
rect 8060 -6452 8072 -6418
rect 8106 -6452 8118 -6418
rect 8060 -6523 8118 -6452
rect 8152 -6322 8346 -6288
rect 8411 -6260 8583 -6245
rect 8617 -6211 8770 -6195
rect 8617 -6245 8733 -6211
rect 8767 -6245 8770 -6211
rect 8152 -6372 8221 -6322
rect 8152 -6406 8171 -6372
rect 8205 -6406 8221 -6372
rect 8152 -6440 8221 -6406
rect 8152 -6474 8171 -6440
rect 8205 -6474 8221 -6440
rect 8152 -6489 8221 -6474
rect 8255 -6372 8321 -6356
rect 8255 -6406 8271 -6372
rect 8305 -6406 8321 -6372
rect 8255 -6440 8321 -6406
rect 8255 -6474 8271 -6440
rect 8305 -6474 8321 -6440
rect 8255 -6523 8321 -6474
rect 8411 -6372 8481 -6260
rect 8617 -6261 8770 -6245
rect 8804 -6217 8854 -6124
rect 8888 -6107 8946 -6013
rect 8888 -6141 8900 -6107
rect 8934 -6141 8946 -6107
rect 8888 -6158 8946 -6141
rect 8980 -6081 9314 -6013
rect 8980 -6115 8998 -6081
rect 9032 -6115 9262 -6081
rect 9296 -6115 9314 -6081
rect 8804 -6251 8811 -6217
rect 8845 -6251 8854 -6217
rect 8617 -6295 8651 -6261
rect 8411 -6406 8429 -6372
rect 8463 -6406 8481 -6372
rect 8411 -6440 8481 -6406
rect 8411 -6474 8429 -6440
rect 8463 -6474 8481 -6440
rect 8411 -6489 8481 -6474
rect 8533 -6329 8651 -6295
rect 8533 -6371 8583 -6329
rect 8804 -6334 8854 -6251
rect 8980 -6167 9314 -6115
rect 9348 -6107 9406 -6013
rect 9348 -6141 9360 -6107
rect 9394 -6141 9406 -6107
rect 9348 -6158 9406 -6141
rect 9440 -6066 9506 -6047
rect 9440 -6100 9459 -6066
rect 9493 -6100 9506 -6066
rect 9440 -6143 9506 -6100
rect 9540 -6066 9606 -6013
rect 9540 -6100 9556 -6066
rect 9590 -6100 9606 -6066
rect 9540 -6109 9606 -6100
rect 9699 -6066 9769 -6047
rect 9699 -6100 9716 -6066
rect 9750 -6100 9769 -6066
rect 8980 -6237 9130 -6167
rect 9440 -6177 9634 -6143
rect 9564 -6201 9634 -6177
rect 8980 -6271 9000 -6237
rect 9034 -6271 9130 -6237
rect 9164 -6235 9260 -6201
rect 9294 -6235 9314 -6201
rect 9564 -6211 9650 -6201
rect 8567 -6405 8583 -6371
rect 8533 -6439 8583 -6405
rect 8567 -6473 8583 -6439
rect 8533 -6489 8583 -6473
rect 8673 -6372 8739 -6363
rect 8673 -6406 8689 -6372
rect 8723 -6406 8739 -6372
rect 8673 -6440 8739 -6406
rect 8673 -6474 8689 -6440
rect 8723 -6474 8739 -6440
rect 8673 -6523 8739 -6474
rect 8773 -6371 8854 -6334
rect 8773 -6405 8787 -6371
rect 8821 -6405 8854 -6371
rect 8773 -6439 8854 -6405
rect 8773 -6473 8787 -6439
rect 8821 -6473 8854 -6439
rect 8773 -6489 8854 -6473
rect 8888 -6325 8946 -6290
rect 9164 -6305 9314 -6235
rect 9440 -6217 9480 -6211
rect 9440 -6251 9453 -6217
rect 9514 -6245 9530 -6211
rect 9487 -6251 9530 -6245
rect 9440 -6254 9530 -6251
rect 9564 -6245 9600 -6211
rect 9634 -6245 9650 -6211
rect 9564 -6259 9650 -6245
rect 9699 -6210 9769 -6100
rect 9821 -6066 9871 -6047
rect 9855 -6100 9871 -6066
rect 9821 -6142 9871 -6100
rect 9961 -6066 10027 -6013
rect 9961 -6100 9977 -6066
rect 10011 -6100 10027 -6066
rect 9961 -6116 10027 -6100
rect 10061 -6066 10142 -6047
rect 10061 -6100 10075 -6066
rect 10109 -6100 10142 -6066
rect 10061 -6124 10142 -6100
rect 9821 -6176 9939 -6142
rect 9905 -6195 9939 -6176
rect 9699 -6211 9871 -6210
rect 9699 -6245 9821 -6211
rect 9855 -6245 9871 -6211
rect 9564 -6288 9634 -6259
rect 8888 -6359 8900 -6325
rect 8934 -6359 8946 -6325
rect 8888 -6418 8946 -6359
rect 8888 -6452 8900 -6418
rect 8934 -6452 8946 -6418
rect 8888 -6523 8946 -6452
rect 8980 -6345 9314 -6305
rect 8980 -6379 8998 -6345
rect 9032 -6379 9262 -6345
rect 9296 -6379 9314 -6345
rect 8980 -6447 9314 -6379
rect 8980 -6481 8998 -6447
rect 9032 -6481 9262 -6447
rect 9296 -6481 9314 -6447
rect 8980 -6523 9314 -6481
rect 9348 -6325 9406 -6290
rect 9348 -6359 9360 -6325
rect 9394 -6359 9406 -6325
rect 9348 -6418 9406 -6359
rect 9348 -6452 9360 -6418
rect 9394 -6452 9406 -6418
rect 9348 -6523 9406 -6452
rect 9440 -6322 9634 -6288
rect 9699 -6260 9871 -6245
rect 9905 -6211 10058 -6195
rect 9905 -6245 10021 -6211
rect 10055 -6245 10058 -6211
rect 9440 -6372 9509 -6322
rect 9440 -6406 9459 -6372
rect 9493 -6406 9509 -6372
rect 9440 -6440 9509 -6406
rect 9440 -6474 9459 -6440
rect 9493 -6474 9509 -6440
rect 9440 -6489 9509 -6474
rect 9543 -6372 9609 -6356
rect 9543 -6406 9559 -6372
rect 9593 -6406 9609 -6372
rect 9543 -6440 9609 -6406
rect 9543 -6474 9559 -6440
rect 9593 -6474 9609 -6440
rect 9543 -6523 9609 -6474
rect 9699 -6372 9769 -6260
rect 9905 -6261 10058 -6245
rect 10092 -6218 10142 -6124
rect 10176 -6107 10234 -6013
rect 10176 -6141 10188 -6107
rect 10222 -6141 10234 -6107
rect 10176 -6158 10234 -6141
rect 10268 -6081 10602 -6013
rect 10268 -6115 10286 -6081
rect 10320 -6115 10550 -6081
rect 10584 -6115 10602 -6081
rect 10092 -6252 10099 -6218
rect 10133 -6252 10142 -6218
rect 9905 -6295 9939 -6261
rect 9699 -6406 9717 -6372
rect 9751 -6406 9769 -6372
rect 9699 -6440 9769 -6406
rect 9699 -6474 9717 -6440
rect 9751 -6474 9769 -6440
rect 9699 -6489 9769 -6474
rect 9821 -6329 9939 -6295
rect 9821 -6371 9871 -6329
rect 10092 -6334 10142 -6252
rect 10268 -6167 10602 -6115
rect 10636 -6107 10694 -6013
rect 10636 -6141 10648 -6107
rect 10682 -6141 10694 -6107
rect 10636 -6158 10694 -6141
rect 10729 -6055 10796 -6047
rect 10729 -6089 10746 -6055
rect 10780 -6089 10796 -6055
rect 10729 -6123 10796 -6089
rect 10830 -6055 10864 -6013
rect 10830 -6105 10864 -6089
rect 10898 -6055 10964 -6047
rect 10898 -6089 10914 -6055
rect 10948 -6089 10964 -6055
rect 10729 -6157 10746 -6123
rect 10780 -6139 10796 -6123
rect 10898 -6123 10964 -6089
rect 10998 -6055 11032 -6013
rect 10998 -6105 11032 -6089
rect 11066 -6055 11468 -6047
rect 11066 -6089 11082 -6055
rect 11116 -6089 11250 -6055
rect 11284 -6089 11418 -6055
rect 11452 -6089 11468 -6055
rect 10898 -6139 10914 -6123
rect 10780 -6157 10914 -6139
rect 10948 -6139 10964 -6123
rect 11066 -6123 11116 -6089
rect 11418 -6123 11468 -6089
rect 11066 -6139 11082 -6123
rect 10948 -6157 11082 -6139
rect 10268 -6237 10418 -6167
rect 10729 -6177 11116 -6157
rect 11150 -6157 11166 -6123
rect 11200 -6157 11334 -6123
rect 11368 -6157 11384 -6123
rect 11452 -6157 11468 -6123
rect 10268 -6271 10288 -6237
rect 10322 -6271 10418 -6237
rect 10452 -6235 10548 -6201
rect 10582 -6235 10602 -6201
rect 11150 -6211 11200 -6157
rect 11418 -6173 11468 -6157
rect 11556 -6107 11614 -6013
rect 11556 -6141 11568 -6107
rect 11602 -6141 11614 -6107
rect 11556 -6158 11614 -6141
rect 11648 -6081 11982 -6013
rect 11648 -6115 11666 -6081
rect 11700 -6115 11930 -6081
rect 11964 -6115 11982 -6081
rect 11648 -6167 11982 -6115
rect 13488 -6107 13546 -6013
rect 13488 -6141 13500 -6107
rect 13534 -6141 13546 -6107
rect 13488 -6158 13546 -6141
rect 13580 -6074 14649 -6013
rect 13580 -6108 13598 -6074
rect 13632 -6108 14598 -6074
rect 14632 -6108 14649 -6074
rect 13580 -6167 14649 -6108
rect 14684 -6107 14742 -6013
rect 14684 -6141 14696 -6107
rect 14730 -6141 14742 -6107
rect 14684 -6158 14742 -6141
rect 14776 -6074 15845 -6013
rect 14776 -6108 14794 -6074
rect 14828 -6108 15794 -6074
rect 15828 -6108 15845 -6074
rect 14776 -6167 15845 -6108
rect 15880 -6107 15938 -6013
rect 15880 -6141 15892 -6107
rect 15926 -6141 15938 -6107
rect 15880 -6158 15938 -6141
rect 15972 -6074 16674 -6013
rect 15972 -6108 15990 -6074
rect 16024 -6108 16622 -6074
rect 16656 -6108 16674 -6074
rect 15972 -6167 16674 -6108
rect 9855 -6405 9871 -6371
rect 9821 -6439 9871 -6405
rect 9855 -6473 9871 -6439
rect 9821 -6489 9871 -6473
rect 9961 -6372 10027 -6363
rect 9961 -6406 9977 -6372
rect 10011 -6406 10027 -6372
rect 9961 -6440 10027 -6406
rect 9961 -6474 9977 -6440
rect 10011 -6474 10027 -6440
rect 9961 -6523 10027 -6474
rect 10061 -6371 10142 -6334
rect 10061 -6405 10075 -6371
rect 10109 -6405 10142 -6371
rect 10061 -6439 10142 -6405
rect 10061 -6473 10075 -6439
rect 10109 -6473 10142 -6439
rect 10061 -6489 10142 -6473
rect 10176 -6325 10234 -6290
rect 10452 -6305 10602 -6235
rect 10733 -6217 10749 -6211
rect 10733 -6251 10741 -6217
rect 10783 -6245 10830 -6211
rect 10864 -6217 10914 -6211
rect 10948 -6216 10998 -6211
rect 11032 -6216 11057 -6211
rect 10866 -6245 10914 -6217
rect 10959 -6245 10998 -6216
rect 10775 -6251 10832 -6245
rect 10866 -6250 10925 -6245
rect 10959 -6250 11017 -6245
rect 11051 -6250 11057 -6216
rect 10866 -6251 11057 -6250
rect 10733 -6261 11057 -6251
rect 11093 -6250 11200 -6211
rect 11093 -6284 11129 -6250
rect 11163 -6284 11200 -6250
rect 11234 -6253 11250 -6211
rect 11284 -6245 11334 -6211
rect 11368 -6219 11522 -6211
rect 11284 -6253 11344 -6245
rect 11378 -6253 11522 -6219
rect 11234 -6261 11522 -6253
rect 11648 -6237 11798 -6167
rect 11648 -6271 11668 -6237
rect 11702 -6271 11798 -6237
rect 11832 -6235 11928 -6201
rect 11962 -6235 11982 -6201
rect 10176 -6359 10188 -6325
rect 10222 -6359 10234 -6325
rect 10176 -6418 10234 -6359
rect 10176 -6452 10188 -6418
rect 10222 -6452 10234 -6418
rect 10176 -6523 10234 -6452
rect 10268 -6345 10602 -6305
rect 10268 -6379 10286 -6345
rect 10320 -6379 10550 -6345
rect 10584 -6379 10602 -6345
rect 10268 -6447 10602 -6379
rect 10268 -6481 10286 -6447
rect 10320 -6481 10550 -6447
rect 10584 -6481 10602 -6447
rect 10268 -6523 10602 -6481
rect 10636 -6325 10694 -6290
rect 11093 -6295 11200 -6284
rect 10636 -6359 10648 -6325
rect 10682 -6359 10694 -6325
rect 10636 -6418 10694 -6359
rect 10636 -6452 10648 -6418
rect 10682 -6452 10694 -6418
rect 10636 -6523 10694 -6452
rect 10729 -6311 10780 -6295
rect 10729 -6345 10746 -6311
rect 10729 -6379 10780 -6345
rect 10729 -6413 10746 -6379
rect 10729 -6447 10780 -6413
rect 10729 -6481 10746 -6447
rect 10729 -6523 10780 -6481
rect 10814 -6311 11384 -6295
rect 10814 -6345 10830 -6311
rect 10864 -6329 10998 -6311
rect 10864 -6345 10880 -6329
rect 10814 -6379 10880 -6345
rect 10982 -6345 10998 -6329
rect 11032 -6329 11166 -6311
rect 11032 -6345 11048 -6329
rect 10814 -6413 10830 -6379
rect 10864 -6413 10880 -6379
rect 10814 -6447 10880 -6413
rect 10814 -6481 10830 -6447
rect 10864 -6481 10880 -6447
rect 10814 -6489 10880 -6481
rect 10914 -6379 10948 -6363
rect 10914 -6447 10948 -6413
rect 10914 -6523 10948 -6481
rect 10982 -6379 11048 -6345
rect 11150 -6345 11166 -6329
rect 11200 -6329 11334 -6311
rect 11200 -6345 11216 -6329
rect 10982 -6413 10998 -6379
rect 11032 -6413 11048 -6379
rect 10982 -6447 11048 -6413
rect 10982 -6481 10998 -6447
rect 11032 -6481 11048 -6447
rect 10982 -6489 11048 -6481
rect 11082 -6379 11116 -6363
rect 11082 -6447 11116 -6413
rect 11082 -6523 11116 -6481
rect 11150 -6379 11216 -6345
rect 11318 -6345 11334 -6329
rect 11368 -6345 11384 -6311
rect 11150 -6413 11166 -6379
rect 11200 -6413 11216 -6379
rect 11150 -6447 11216 -6413
rect 11150 -6481 11166 -6447
rect 11200 -6481 11216 -6447
rect 11150 -6489 11216 -6481
rect 11250 -6379 11284 -6363
rect 11250 -6447 11284 -6413
rect 11250 -6523 11284 -6481
rect 11318 -6379 11384 -6345
rect 11556 -6325 11614 -6290
rect 11832 -6305 11982 -6235
rect 13580 -6237 14096 -6167
rect 13580 -6271 13658 -6237
rect 13692 -6271 13786 -6237
rect 13820 -6271 13914 -6237
rect 13948 -6271 14042 -6237
rect 14076 -6271 14096 -6237
rect 14130 -6235 14150 -6201
rect 14184 -6235 14278 -6201
rect 14312 -6235 14406 -6201
rect 14440 -6235 14534 -6201
rect 14568 -6235 14649 -6201
rect 11556 -6359 11568 -6325
rect 11602 -6359 11614 -6325
rect 11318 -6413 11334 -6379
rect 11368 -6413 11384 -6379
rect 11318 -6447 11384 -6413
rect 11318 -6481 11334 -6447
rect 11368 -6481 11384 -6447
rect 11318 -6489 11384 -6481
rect 11418 -6379 11468 -6363
rect 11452 -6413 11468 -6379
rect 11418 -6447 11468 -6413
rect 11452 -6481 11468 -6447
rect 11418 -6523 11468 -6481
rect 11556 -6418 11614 -6359
rect 11556 -6452 11568 -6418
rect 11602 -6452 11614 -6418
rect 11556 -6523 11614 -6452
rect 11648 -6345 11982 -6305
rect 11648 -6379 11666 -6345
rect 11700 -6379 11930 -6345
rect 11964 -6379 11982 -6345
rect 11648 -6447 11982 -6379
rect 11648 -6481 11666 -6447
rect 11700 -6481 11930 -6447
rect 11964 -6481 11982 -6447
rect 11648 -6523 11982 -6481
rect 13488 -6325 13546 -6290
rect 14130 -6305 14649 -6235
rect 14776 -6237 15292 -6167
rect 14776 -6271 14854 -6237
rect 14888 -6271 14982 -6237
rect 15016 -6271 15110 -6237
rect 15144 -6271 15238 -6237
rect 15272 -6271 15292 -6237
rect 15326 -6235 15346 -6201
rect 15380 -6235 15474 -6201
rect 15508 -6235 15602 -6201
rect 15636 -6235 15730 -6201
rect 15764 -6235 15845 -6201
rect 13488 -6359 13500 -6325
rect 13534 -6359 13546 -6325
rect 13488 -6418 13546 -6359
rect 13488 -6452 13500 -6418
rect 13534 -6452 13546 -6418
rect 13488 -6523 13546 -6452
rect 13580 -6345 14649 -6305
rect 13580 -6379 13598 -6345
rect 13632 -6379 14598 -6345
rect 14632 -6379 14649 -6345
rect 13580 -6447 14649 -6379
rect 13580 -6481 13598 -6447
rect 13632 -6481 14598 -6447
rect 14632 -6481 14649 -6447
rect 13580 -6523 14649 -6481
rect 14684 -6325 14742 -6290
rect 15326 -6305 15845 -6235
rect 15972 -6237 16302 -6167
rect 15972 -6271 16050 -6237
rect 16084 -6271 16149 -6237
rect 16183 -6271 16248 -6237
rect 16282 -6271 16302 -6237
rect 16336 -6235 16356 -6201
rect 16390 -6235 16459 -6201
rect 16493 -6235 16562 -6201
rect 16596 -6235 16674 -6201
rect 14684 -6359 14696 -6325
rect 14730 -6359 14742 -6325
rect 14684 -6418 14742 -6359
rect 14684 -6452 14696 -6418
rect 14730 -6452 14742 -6418
rect 14684 -6523 14742 -6452
rect 14776 -6345 15845 -6305
rect 14776 -6379 14794 -6345
rect 14828 -6379 15794 -6345
rect 15828 -6379 15845 -6345
rect 14776 -6447 15845 -6379
rect 14776 -6481 14794 -6447
rect 14828 -6481 15794 -6447
rect 15828 -6481 15845 -6447
rect 14776 -6523 15845 -6481
rect 15880 -6325 15938 -6290
rect 16336 -6305 16674 -6235
rect 15880 -6359 15892 -6325
rect 15926 -6359 15938 -6325
rect 15880 -6418 15938 -6359
rect 15880 -6452 15892 -6418
rect 15926 -6452 15938 -6418
rect 15880 -6523 15938 -6452
rect 15972 -6345 16674 -6305
rect 15972 -6379 15990 -6345
rect 16024 -6379 16622 -6345
rect 16656 -6379 16674 -6345
rect 15972 -6447 16674 -6379
rect 15972 -6481 15990 -6447
rect 16024 -6481 16622 -6447
rect 16656 -6481 16674 -6447
rect 15972 -6523 16674 -6481
rect -2997 -6557 -2968 -6523
rect -2934 -6557 -2876 -6523
rect -2842 -6557 -2784 -6523
rect -2750 -6557 -2692 -6523
rect -2658 -6557 -2600 -6523
rect -2566 -6557 -2508 -6523
rect -2474 -6557 -2416 -6523
rect -2382 -6557 -2324 -6523
rect -2290 -6557 -2232 -6523
rect -2198 -6557 -2140 -6523
rect -2106 -6557 -2048 -6523
rect -2014 -6557 -1956 -6523
rect -1922 -6557 -1864 -6523
rect -1830 -6557 -1772 -6523
rect -1738 -6557 -1680 -6523
rect -1646 -6557 -1588 -6523
rect -1554 -6557 -1496 -6523
rect -1462 -6557 -1404 -6523
rect -1370 -6557 -1312 -6523
rect -1278 -6557 -1220 -6523
rect -1186 -6557 -1128 -6523
rect -1094 -6557 -1036 -6523
rect -1002 -6557 -944 -6523
rect -910 -6557 -852 -6523
rect -818 -6557 -760 -6523
rect -726 -6557 -668 -6523
rect -634 -6557 -576 -6523
rect -542 -6557 -484 -6523
rect -450 -6557 -392 -6523
rect -358 -6557 -300 -6523
rect -266 -6557 -208 -6523
rect -174 -6557 -116 -6523
rect -82 -6557 -24 -6523
rect 10 -6557 68 -6523
rect 102 -6557 160 -6523
rect 194 -6557 252 -6523
rect 286 -6557 344 -6523
rect 378 -6557 436 -6523
rect 470 -6557 528 -6523
rect 562 -6557 620 -6523
rect 654 -6557 712 -6523
rect 746 -6557 804 -6523
rect 838 -6557 896 -6523
rect 930 -6557 988 -6523
rect 1022 -6557 1080 -6523
rect 1114 -6557 1172 -6523
rect 1206 -6557 1264 -6523
rect 1298 -6557 1356 -6523
rect 1390 -6557 1448 -6523
rect 1482 -6557 1540 -6523
rect 1574 -6557 1632 -6523
rect 1666 -6557 1724 -6523
rect 1758 -6557 1816 -6523
rect 1850 -6557 1908 -6523
rect 1942 -6557 2000 -6523
rect 2034 -6557 2092 -6523
rect 2126 -6557 2184 -6523
rect 2218 -6557 2276 -6523
rect 2310 -6557 2368 -6523
rect 2402 -6557 2460 -6523
rect 2494 -6557 2552 -6523
rect 2586 -6557 2644 -6523
rect 2678 -6557 2736 -6523
rect 2770 -6557 2828 -6523
rect 2862 -6557 2920 -6523
rect 2954 -6557 3012 -6523
rect 3046 -6557 3104 -6523
rect 3138 -6557 3196 -6523
rect 3230 -6557 3288 -6523
rect 3322 -6557 3380 -6523
rect 3414 -6557 3472 -6523
rect 3506 -6557 3564 -6523
rect 3598 -6557 3656 -6523
rect 3690 -6557 3748 -6523
rect 3782 -6557 3840 -6523
rect 3874 -6557 3932 -6523
rect 3966 -6557 4024 -6523
rect 4058 -6557 4116 -6523
rect 4150 -6557 4208 -6523
rect 4242 -6557 4300 -6523
rect 4334 -6557 4392 -6523
rect 4426 -6557 4484 -6523
rect 4518 -6557 4576 -6523
rect 4610 -6557 4668 -6523
rect 4702 -6557 4760 -6523
rect 4794 -6557 4852 -6523
rect 4886 -6557 4944 -6523
rect 4978 -6557 5036 -6523
rect 5070 -6557 5128 -6523
rect 5162 -6557 5220 -6523
rect 5254 -6557 5312 -6523
rect 5346 -6557 5404 -6523
rect 5438 -6557 5496 -6523
rect 5530 -6557 5588 -6523
rect 5622 -6557 5680 -6523
rect 5714 -6557 5772 -6523
rect 5806 -6557 5864 -6523
rect 5898 -6557 5956 -6523
rect 5990 -6557 6048 -6523
rect 6082 -6557 6140 -6523
rect 6174 -6557 6232 -6523
rect 6266 -6557 6324 -6523
rect 6358 -6557 6416 -6523
rect 6450 -6557 6508 -6523
rect 6542 -6557 6600 -6523
rect 6634 -6557 6692 -6523
rect 6726 -6557 6784 -6523
rect 6818 -6557 6876 -6523
rect 6910 -6557 6968 -6523
rect 7002 -6557 7060 -6523
rect 7094 -6557 7152 -6523
rect 7186 -6557 7244 -6523
rect 7278 -6557 7336 -6523
rect 7370 -6557 7428 -6523
rect 7462 -6557 7520 -6523
rect 7554 -6557 7612 -6523
rect 7646 -6557 7704 -6523
rect 7738 -6557 7796 -6523
rect 7830 -6557 7888 -6523
rect 7922 -6557 7980 -6523
rect 8014 -6557 8072 -6523
rect 8106 -6557 8164 -6523
rect 8198 -6557 8256 -6523
rect 8290 -6557 8348 -6523
rect 8382 -6557 8440 -6523
rect 8474 -6557 8532 -6523
rect 8566 -6557 8624 -6523
rect 8658 -6557 8716 -6523
rect 8750 -6557 8808 -6523
rect 8842 -6557 8900 -6523
rect 8934 -6557 8992 -6523
rect 9026 -6557 9084 -6523
rect 9118 -6557 9176 -6523
rect 9210 -6557 9268 -6523
rect 9302 -6557 9360 -6523
rect 9394 -6557 9452 -6523
rect 9486 -6557 9544 -6523
rect 9578 -6557 9636 -6523
rect 9670 -6557 9728 -6523
rect 9762 -6557 9820 -6523
rect 9854 -6557 9912 -6523
rect 9946 -6557 10004 -6523
rect 10038 -6557 10096 -6523
rect 10130 -6557 10188 -6523
rect 10222 -6557 10280 -6523
rect 10314 -6557 10372 -6523
rect 10406 -6557 10464 -6523
rect 10498 -6557 10556 -6523
rect 10590 -6557 10648 -6523
rect 10682 -6557 10740 -6523
rect 10774 -6557 10832 -6523
rect 10866 -6557 10924 -6523
rect 10958 -6557 11016 -6523
rect 11050 -6557 11108 -6523
rect 11142 -6557 11200 -6523
rect 11234 -6557 11292 -6523
rect 11326 -6557 11384 -6523
rect 11418 -6557 11476 -6523
rect 11510 -6557 11568 -6523
rect 11602 -6557 11660 -6523
rect 11694 -6557 11752 -6523
rect 11786 -6557 11844 -6523
rect 11878 -6557 11936 -6523
rect 11970 -6557 12028 -6523
rect 12062 -6557 12120 -6523
rect 12154 -6557 12212 -6523
rect 12246 -6557 12304 -6523
rect 12338 -6557 12396 -6523
rect 12430 -6557 12488 -6523
rect 12522 -6557 12580 -6523
rect 12614 -6557 12672 -6523
rect 12706 -6557 12764 -6523
rect 12798 -6557 12856 -6523
rect 12890 -6557 12948 -6523
rect 12982 -6557 13040 -6523
rect 13074 -6557 13132 -6523
rect 13166 -6557 13224 -6523
rect 13258 -6557 13316 -6523
rect 13350 -6557 13408 -6523
rect 13442 -6557 13500 -6523
rect 13534 -6557 13592 -6523
rect 13626 -6557 13684 -6523
rect 13718 -6557 13776 -6523
rect 13810 -6557 13868 -6523
rect 13902 -6557 13960 -6523
rect 13994 -6557 14052 -6523
rect 14086 -6557 14144 -6523
rect 14178 -6557 14236 -6523
rect 14270 -6557 14328 -6523
rect 14362 -6557 14420 -6523
rect 14454 -6557 14512 -6523
rect 14546 -6557 14604 -6523
rect 14638 -6557 14696 -6523
rect 14730 -6557 14788 -6523
rect 14822 -6557 14880 -6523
rect 14914 -6557 14972 -6523
rect 15006 -6557 15064 -6523
rect 15098 -6557 15156 -6523
rect 15190 -6557 15248 -6523
rect 15282 -6557 15340 -6523
rect 15374 -6557 15432 -6523
rect 15466 -6557 15524 -6523
rect 15558 -6557 15616 -6523
rect 15650 -6557 15708 -6523
rect 15742 -6557 15800 -6523
rect 15834 -6557 15892 -6523
rect 15926 -6557 15984 -6523
rect 16018 -6557 16076 -6523
rect 16110 -6557 16168 -6523
rect 16202 -6557 16260 -6523
rect 16294 -6557 16352 -6523
rect 16386 -6557 16444 -6523
rect 16478 -6557 16536 -6523
rect 16570 -6557 16628 -6523
rect 16662 -6557 16691 -6523
rect -2980 -6599 -2738 -6557
rect -2980 -6633 -2962 -6599
rect -2928 -6633 -2790 -6599
rect -2756 -6633 -2738 -6599
rect -2980 -6694 -2738 -6633
rect -2980 -6728 -2962 -6694
rect -2928 -6728 -2790 -6694
rect -2756 -6728 -2738 -6694
rect -2980 -6775 -2738 -6728
rect -2980 -6843 -2930 -6809
rect -2896 -6843 -2876 -6809
rect -2980 -6917 -2876 -6843
rect -2842 -6849 -2738 -6775
rect -2704 -6628 -2646 -6557
rect -2704 -6662 -2692 -6628
rect -2658 -6662 -2646 -6628
rect -2704 -6721 -2646 -6662
rect -2704 -6755 -2692 -6721
rect -2658 -6755 -2646 -6721
rect -2594 -6607 -2560 -6591
rect -2594 -6675 -2560 -6641
rect -2526 -6623 -2460 -6557
rect -2526 -6657 -2510 -6623
rect -2476 -6657 -2460 -6623
rect -2426 -6607 -2389 -6591
rect -2392 -6641 -2389 -6607
rect -2426 -6675 -2389 -6641
rect -2341 -6599 -2288 -6557
rect -2341 -6633 -2322 -6599
rect -2341 -6649 -2288 -6633
rect -2254 -6607 -2204 -6591
rect -2254 -6641 -2238 -6607
rect -1907 -6599 -1873 -6557
rect -2560 -6693 -2461 -6691
rect -2560 -6709 -2503 -6693
rect -2594 -6725 -2503 -6709
rect -2704 -6790 -2646 -6755
rect -2507 -6727 -2503 -6725
rect -2469 -6727 -2461 -6693
rect -2842 -6883 -2822 -6849
rect -2788 -6883 -2738 -6849
rect -2611 -6830 -2541 -6759
rect -2611 -6864 -2599 -6830
rect -2565 -6835 -2541 -6830
rect -2611 -6869 -2597 -6864
rect -2563 -6869 -2541 -6835
rect -2611 -6889 -2541 -6869
rect -2507 -6820 -2461 -6727
rect -2507 -6854 -2495 -6820
rect -2980 -6970 -2738 -6917
rect -2980 -7004 -2962 -6970
rect -2928 -7004 -2790 -6970
rect -2756 -7004 -2738 -6970
rect -2980 -7067 -2738 -7004
rect -2704 -6939 -2646 -6922
rect -2507 -6923 -2461 -6854
rect -2704 -6973 -2692 -6939
rect -2658 -6973 -2646 -6939
rect -2704 -7067 -2646 -6973
rect -2594 -6957 -2461 -6923
rect -2392 -6709 -2389 -6675
rect -2254 -6676 -2204 -6641
rect -2162 -6646 -2146 -6612
rect -2112 -6646 -1941 -6612
rect -2426 -6761 -2389 -6709
rect -2265 -6702 -2204 -6676
rect -2115 -6693 -2009 -6680
rect -2426 -6795 -2424 -6761
rect -2390 -6795 -2389 -6761
rect -2594 -6965 -2560 -6957
rect -2426 -6965 -2389 -6795
rect -2355 -6767 -2299 -6751
rect -2355 -6801 -2333 -6767
rect -2355 -6882 -2299 -6801
rect -2355 -6916 -2343 -6882
rect -2309 -6916 -2299 -6882
rect -2355 -6941 -2299 -6916
rect -2265 -6923 -2231 -6702
rect -2115 -6727 -2083 -6693
rect -2049 -6719 -2009 -6693
rect -2197 -6761 -2149 -6740
rect -2197 -6795 -2186 -6761
rect -2152 -6795 -2149 -6761
rect -2197 -6797 -2149 -6795
rect -2197 -6831 -2190 -6797
rect -2156 -6831 -2149 -6797
rect -2197 -6859 -2149 -6831
rect -2115 -6893 -2081 -6727
rect -2047 -6753 -2009 -6719
rect -1975 -6769 -1941 -6646
rect -1907 -6667 -1873 -6633
rect -1907 -6717 -1873 -6701
rect -1839 -6607 -1789 -6591
rect -1839 -6641 -1823 -6607
rect -1531 -6607 -1468 -6557
rect -1839 -6657 -1789 -6641
rect -1744 -6651 -1728 -6617
rect -1694 -6651 -1567 -6617
rect -1975 -6785 -1873 -6769
rect -1975 -6787 -1907 -6785
rect -2265 -6949 -2220 -6923
rect -2186 -6927 -2170 -6893
rect -2136 -6927 -2081 -6893
rect -2186 -6937 -2081 -6927
rect -2047 -6819 -1907 -6787
rect -2047 -6821 -1873 -6819
rect -2594 -7015 -2560 -6999
rect -2526 -7025 -2510 -6991
rect -2476 -7025 -2460 -6991
rect -2392 -6999 -2389 -6965
rect -2426 -7015 -2389 -6999
rect -2338 -6991 -2288 -6975
rect -2526 -7067 -2460 -7025
rect -2338 -7025 -2322 -6991
rect -2254 -6977 -2220 -6949
rect -2047 -6977 -2013 -6821
rect -1907 -6835 -1873 -6821
rect -1971 -6871 -1931 -6865
rect -1839 -6871 -1805 -6657
rect -1771 -6693 -1733 -6691
rect -1771 -6727 -1769 -6693
rect -1735 -6727 -1733 -6693
rect -1771 -6785 -1733 -6727
rect -1737 -6819 -1733 -6785
rect -1771 -6835 -1733 -6819
rect -1699 -6719 -1635 -6685
rect -1699 -6753 -1669 -6719
rect -1699 -6761 -1635 -6753
rect -1699 -6795 -1682 -6761
rect -1648 -6795 -1635 -6761
rect -1971 -6881 -1805 -6871
rect -1699 -6877 -1635 -6795
rect -1937 -6915 -1805 -6881
rect -1971 -6931 -1805 -6915
rect -2254 -7011 -2237 -6977
rect -2203 -7011 -2187 -6977
rect -2148 -7011 -2126 -6977
rect -2092 -7011 -2013 -6977
rect -1949 -6983 -1875 -6967
rect -2338 -7067 -2288 -7025
rect -1949 -7017 -1927 -6983
rect -1893 -7017 -1875 -6983
rect -1839 -6977 -1805 -6931
rect -1728 -6893 -1635 -6877
rect -1694 -6927 -1635 -6893
rect -1728 -6943 -1635 -6927
rect -1601 -6819 -1567 -6651
rect -1531 -6641 -1529 -6607
rect -1495 -6641 -1468 -6607
rect -1531 -6657 -1468 -6641
rect -1421 -6599 -1353 -6591
rect -1421 -6633 -1405 -6599
rect -1371 -6633 -1353 -6599
rect -1421 -6670 -1353 -6633
rect -1421 -6703 -1405 -6670
rect -1533 -6704 -1405 -6703
rect -1371 -6704 -1353 -6670
rect -1533 -6719 -1353 -6704
rect -1499 -6741 -1353 -6719
rect -1499 -6753 -1405 -6741
rect -1533 -6775 -1405 -6753
rect -1371 -6775 -1353 -6741
rect -1319 -6629 -1285 -6557
rect -1147 -6599 -1081 -6595
rect -1319 -6709 -1285 -6663
rect -1319 -6759 -1285 -6743
rect -1251 -6605 -1185 -6600
rect -1251 -6639 -1235 -6605
rect -1201 -6639 -1185 -6605
rect -1251 -6673 -1185 -6639
rect -1251 -6707 -1235 -6673
rect -1201 -6707 -1185 -6673
rect -1251 -6741 -1185 -6707
rect -1147 -6633 -1131 -6599
rect -1097 -6633 -1081 -6599
rect -1147 -6667 -1081 -6633
rect -1147 -6701 -1131 -6667
rect -1097 -6701 -1081 -6667
rect -1147 -6741 -1081 -6701
rect -1533 -6778 -1353 -6775
rect -1391 -6819 -1353 -6778
rect -1251 -6775 -1235 -6741
rect -1201 -6769 -1185 -6741
rect -1201 -6775 -1169 -6769
rect -1251 -6785 -1169 -6775
rect -1216 -6795 -1169 -6785
rect -1601 -6835 -1425 -6819
rect -1601 -6869 -1459 -6835
rect -1601 -6885 -1425 -6869
rect -1391 -6835 -1241 -6819
rect -1391 -6869 -1275 -6835
rect -1391 -6885 -1241 -6869
rect -1601 -6977 -1567 -6885
rect -1391 -6919 -1351 -6885
rect -1207 -6911 -1169 -6795
rect -1218 -6919 -1169 -6911
rect -1417 -6922 -1351 -6919
rect -1417 -6956 -1401 -6922
rect -1367 -6956 -1351 -6922
rect -1249 -6920 -1169 -6919
rect -1839 -7011 -1808 -6977
rect -1774 -7011 -1758 -6977
rect -1724 -7011 -1705 -6977
rect -1671 -7011 -1567 -6977
rect -1512 -6977 -1470 -6961
rect -1512 -7011 -1507 -6977
rect -1473 -7011 -1470 -6977
rect -1949 -7067 -1875 -7017
rect -1512 -7067 -1470 -7011
rect -1417 -6990 -1351 -6956
rect -1417 -7024 -1401 -6990
rect -1367 -7024 -1351 -6990
rect -1317 -6961 -1283 -6945
rect -1317 -7067 -1283 -6995
rect -1249 -6954 -1233 -6920
rect -1199 -6936 -1169 -6920
rect -1135 -6819 -1081 -6741
rect -1043 -6599 -1000 -6557
rect -1043 -6633 -1034 -6599
rect -1043 -6667 -1000 -6633
rect -1043 -6701 -1034 -6667
rect -1043 -6735 -1000 -6701
rect -1043 -6769 -1034 -6735
rect -1043 -6785 -1000 -6769
rect -966 -6599 -899 -6591
rect -966 -6633 -950 -6599
rect -916 -6633 -899 -6599
rect -966 -6670 -899 -6633
rect -966 -6704 -950 -6670
rect -916 -6704 -899 -6670
rect -966 -6741 -899 -6704
rect -966 -6775 -950 -6741
rect -916 -6775 -899 -6741
rect -966 -6788 -899 -6775
rect -1135 -6835 -980 -6819
rect -1135 -6869 -1014 -6835
rect -1135 -6885 -980 -6869
rect -946 -6880 -899 -6788
rect -864 -6599 -162 -6557
rect -864 -6633 -846 -6599
rect -812 -6633 -214 -6599
rect -180 -6633 -162 -6599
rect -864 -6701 -162 -6633
rect -864 -6735 -846 -6701
rect -812 -6735 -214 -6701
rect -180 -6735 -162 -6701
rect -864 -6775 -162 -6735
rect -128 -6628 -70 -6557
rect -128 -6662 -116 -6628
rect -82 -6662 -70 -6628
rect -128 -6721 -70 -6662
rect -128 -6755 -116 -6721
rect -82 -6755 -70 -6721
rect -864 -6845 -526 -6775
rect -128 -6790 -70 -6755
rect -36 -6599 666 -6557
rect -36 -6633 -18 -6599
rect 16 -6633 614 -6599
rect 648 -6633 666 -6599
rect -36 -6701 666 -6633
rect -36 -6735 -18 -6701
rect 16 -6735 614 -6701
rect 648 -6735 666 -6701
rect -36 -6775 666 -6735
rect 700 -6599 1402 -6557
rect 700 -6633 718 -6599
rect 752 -6633 1350 -6599
rect 1384 -6633 1402 -6599
rect 700 -6701 1402 -6633
rect 700 -6735 718 -6701
rect 752 -6735 1350 -6701
rect 1384 -6735 1402 -6701
rect 700 -6775 1402 -6735
rect 1436 -6628 1494 -6557
rect 1436 -6662 1448 -6628
rect 1482 -6662 1494 -6628
rect 1436 -6721 1494 -6662
rect 1436 -6755 1448 -6721
rect 1482 -6755 1494 -6721
rect -864 -6879 -786 -6845
rect -752 -6879 -683 -6845
rect -649 -6879 -580 -6845
rect -546 -6879 -526 -6845
rect -492 -6843 -472 -6809
rect -438 -6843 -373 -6809
rect -339 -6843 -274 -6809
rect -240 -6843 -162 -6809
rect -1199 -6954 -1183 -6936
rect -1249 -6960 -1183 -6954
rect -1249 -7022 -1233 -6960
rect -1199 -7022 -1183 -6960
rect -1135 -6961 -1095 -6885
rect -946 -6902 -940 -6880
rect -1145 -6965 -1095 -6961
rect -1145 -6999 -1129 -6965
rect -950 -6914 -940 -6902
rect -906 -6914 -899 -6880
rect -492 -6913 -162 -6843
rect -36 -6845 302 -6775
rect -36 -6879 42 -6845
rect 76 -6879 145 -6845
rect 179 -6879 248 -6845
rect 282 -6879 302 -6845
rect 336 -6843 356 -6809
rect 390 -6843 455 -6809
rect 489 -6843 554 -6809
rect 588 -6843 666 -6809
rect 336 -6913 666 -6843
rect 700 -6845 1038 -6775
rect 1436 -6790 1494 -6755
rect 1528 -6599 2230 -6557
rect 1528 -6633 1546 -6599
rect 1580 -6633 2178 -6599
rect 2212 -6633 2230 -6599
rect 1528 -6701 2230 -6633
rect 1528 -6735 1546 -6701
rect 1580 -6735 2178 -6701
rect 2212 -6735 2230 -6701
rect 1528 -6775 2230 -6735
rect 2264 -6599 2966 -6557
rect 2264 -6633 2282 -6599
rect 2316 -6633 2914 -6599
rect 2948 -6633 2966 -6599
rect 2264 -6701 2966 -6633
rect 2264 -6735 2282 -6701
rect 2316 -6735 2914 -6701
rect 2948 -6735 2966 -6701
rect 2264 -6775 2966 -6735
rect 3000 -6628 3058 -6557
rect 3000 -6662 3012 -6628
rect 3046 -6662 3058 -6628
rect 3000 -6721 3058 -6662
rect 3000 -6755 3012 -6721
rect 3046 -6755 3058 -6721
rect 700 -6879 778 -6845
rect 812 -6879 881 -6845
rect 915 -6879 984 -6845
rect 1018 -6879 1038 -6845
rect 1072 -6843 1092 -6809
rect 1126 -6843 1191 -6809
rect 1225 -6843 1290 -6809
rect 1324 -6843 1402 -6809
rect 1072 -6913 1402 -6843
rect 1528 -6845 1866 -6775
rect 1528 -6879 1606 -6845
rect 1640 -6879 1709 -6845
rect 1743 -6879 1812 -6845
rect 1846 -6879 1866 -6845
rect 1900 -6843 1920 -6809
rect 1954 -6843 2019 -6809
rect 2053 -6843 2118 -6809
rect 2152 -6843 2230 -6809
rect 1900 -6913 2230 -6843
rect 2264 -6845 2602 -6775
rect 3000 -6790 3058 -6755
rect 3092 -6599 3794 -6557
rect 3092 -6633 3110 -6599
rect 3144 -6633 3742 -6599
rect 3776 -6633 3794 -6599
rect 3092 -6701 3794 -6633
rect 3092 -6735 3110 -6701
rect 3144 -6735 3742 -6701
rect 3776 -6735 3794 -6701
rect 3092 -6775 3794 -6735
rect 3828 -6599 4530 -6557
rect 3828 -6633 3846 -6599
rect 3880 -6633 4478 -6599
rect 4512 -6633 4530 -6599
rect 3828 -6701 4530 -6633
rect 3828 -6735 3846 -6701
rect 3880 -6735 4478 -6701
rect 4512 -6735 4530 -6701
rect 3828 -6775 4530 -6735
rect 4564 -6628 4622 -6557
rect 4564 -6662 4576 -6628
rect 4610 -6662 4622 -6628
rect 4564 -6721 4622 -6662
rect 4564 -6755 4576 -6721
rect 4610 -6755 4622 -6721
rect 2264 -6879 2342 -6845
rect 2376 -6879 2445 -6845
rect 2479 -6879 2548 -6845
rect 2582 -6879 2602 -6845
rect 2636 -6843 2656 -6809
rect 2690 -6843 2755 -6809
rect 2789 -6843 2854 -6809
rect 2888 -6843 2966 -6809
rect 2636 -6913 2966 -6843
rect 3092 -6845 3430 -6775
rect 3092 -6879 3170 -6845
rect 3204 -6879 3273 -6845
rect 3307 -6879 3376 -6845
rect 3410 -6879 3430 -6845
rect 3464 -6843 3484 -6809
rect 3518 -6843 3583 -6809
rect 3617 -6843 3682 -6809
rect 3716 -6843 3794 -6809
rect 3464 -6913 3794 -6843
rect 3828 -6845 4166 -6775
rect 4564 -6790 4622 -6755
rect 4656 -6599 5358 -6557
rect 4656 -6633 4674 -6599
rect 4708 -6633 5306 -6599
rect 5340 -6633 5358 -6599
rect 4656 -6701 5358 -6633
rect 4656 -6735 4674 -6701
rect 4708 -6735 5306 -6701
rect 5340 -6735 5358 -6701
rect 4656 -6775 5358 -6735
rect 5392 -6599 6094 -6557
rect 5392 -6633 5410 -6599
rect 5444 -6633 6042 -6599
rect 6076 -6633 6094 -6599
rect 5392 -6701 6094 -6633
rect 5392 -6735 5410 -6701
rect 5444 -6735 6042 -6701
rect 6076 -6735 6094 -6701
rect 5392 -6775 6094 -6735
rect 6128 -6628 6186 -6557
rect 6128 -6662 6140 -6628
rect 6174 -6662 6186 -6628
rect 6128 -6721 6186 -6662
rect 6128 -6755 6140 -6721
rect 6174 -6755 6186 -6721
rect 3828 -6879 3906 -6845
rect 3940 -6879 4009 -6845
rect 4043 -6879 4112 -6845
rect 4146 -6879 4166 -6845
rect 4200 -6843 4220 -6809
rect 4254 -6843 4319 -6809
rect 4353 -6843 4418 -6809
rect 4452 -6843 4530 -6809
rect 4200 -6913 4530 -6843
rect 4656 -6845 4994 -6775
rect 4656 -6879 4734 -6845
rect 4768 -6879 4837 -6845
rect 4871 -6879 4940 -6845
rect 4974 -6879 4994 -6845
rect 5028 -6843 5048 -6809
rect 5082 -6843 5147 -6809
rect 5181 -6843 5246 -6809
rect 5280 -6843 5358 -6809
rect 5028 -6913 5358 -6843
rect 5392 -6845 5730 -6775
rect 6128 -6790 6186 -6755
rect 6220 -6599 6922 -6557
rect 6220 -6633 6238 -6599
rect 6272 -6633 6870 -6599
rect 6904 -6633 6922 -6599
rect 6220 -6701 6922 -6633
rect 6220 -6735 6238 -6701
rect 6272 -6735 6870 -6701
rect 6904 -6735 6922 -6701
rect 6220 -6775 6922 -6735
rect 6956 -6599 7658 -6557
rect 6956 -6633 6974 -6599
rect 7008 -6633 7606 -6599
rect 7640 -6633 7658 -6599
rect 6956 -6701 7658 -6633
rect 6956 -6735 6974 -6701
rect 7008 -6735 7606 -6701
rect 7640 -6735 7658 -6701
rect 6956 -6775 7658 -6735
rect 7692 -6628 7750 -6557
rect 7692 -6662 7704 -6628
rect 7738 -6662 7750 -6628
rect 7692 -6721 7750 -6662
rect 7692 -6755 7704 -6721
rect 7738 -6755 7750 -6721
rect 5392 -6879 5470 -6845
rect 5504 -6879 5573 -6845
rect 5607 -6879 5676 -6845
rect 5710 -6879 5730 -6845
rect 5764 -6843 5784 -6809
rect 5818 -6843 5883 -6809
rect 5917 -6843 5982 -6809
rect 6016 -6843 6094 -6809
rect 5764 -6913 6094 -6843
rect 6220 -6845 6558 -6775
rect 6220 -6879 6298 -6845
rect 6332 -6879 6401 -6845
rect 6435 -6879 6504 -6845
rect 6538 -6879 6558 -6845
rect 6592 -6843 6612 -6809
rect 6646 -6843 6711 -6809
rect 6745 -6843 6810 -6809
rect 6844 -6843 6922 -6809
rect 6592 -6913 6922 -6843
rect 6956 -6845 7294 -6775
rect 7692 -6790 7750 -6755
rect 7784 -6599 8486 -6557
rect 7784 -6633 7802 -6599
rect 7836 -6633 8434 -6599
rect 8468 -6633 8486 -6599
rect 7784 -6701 8486 -6633
rect 7784 -6735 7802 -6701
rect 7836 -6735 8434 -6701
rect 8468 -6735 8486 -6701
rect 7784 -6775 8486 -6735
rect 8520 -6599 9222 -6557
rect 8520 -6633 8538 -6599
rect 8572 -6633 9170 -6599
rect 9204 -6633 9222 -6599
rect 8520 -6701 9222 -6633
rect 8520 -6735 8538 -6701
rect 8572 -6735 9170 -6701
rect 9204 -6735 9222 -6701
rect 8520 -6775 9222 -6735
rect 9256 -6628 9314 -6557
rect 9256 -6662 9268 -6628
rect 9302 -6662 9314 -6628
rect 9256 -6721 9314 -6662
rect 9256 -6755 9268 -6721
rect 9302 -6755 9314 -6721
rect 6956 -6879 7034 -6845
rect 7068 -6879 7137 -6845
rect 7171 -6879 7240 -6845
rect 7274 -6879 7294 -6845
rect 7328 -6843 7348 -6809
rect 7382 -6843 7447 -6809
rect 7481 -6843 7546 -6809
rect 7580 -6843 7658 -6809
rect 7328 -6913 7658 -6843
rect 7784 -6845 8122 -6775
rect 7784 -6879 7862 -6845
rect 7896 -6879 7965 -6845
rect 7999 -6879 8068 -6845
rect 8102 -6879 8122 -6845
rect 8156 -6843 8176 -6809
rect 8210 -6843 8275 -6809
rect 8309 -6843 8374 -6809
rect 8408 -6843 8486 -6809
rect 8156 -6913 8486 -6843
rect 8520 -6845 8858 -6775
rect 9256 -6790 9314 -6755
rect 15880 -6628 15938 -6557
rect 15880 -6662 15892 -6628
rect 15926 -6662 15938 -6628
rect 15880 -6721 15938 -6662
rect 15880 -6755 15892 -6721
rect 15926 -6755 15938 -6721
rect 15880 -6790 15938 -6755
rect 15972 -6599 16674 -6557
rect 15972 -6633 15990 -6599
rect 16024 -6633 16622 -6599
rect 16656 -6633 16674 -6599
rect 15972 -6701 16674 -6633
rect 15972 -6735 15990 -6701
rect 16024 -6735 16622 -6701
rect 16656 -6735 16674 -6701
rect 15972 -6775 16674 -6735
rect 8520 -6879 8598 -6845
rect 8632 -6879 8701 -6845
rect 8735 -6879 8804 -6845
rect 8838 -6879 8858 -6845
rect 8892 -6843 8912 -6809
rect 8946 -6843 9011 -6809
rect 9045 -6843 9110 -6809
rect 9144 -6843 9222 -6809
rect 8892 -6913 9222 -6843
rect 15972 -6845 16310 -6775
rect 15972 -6879 16050 -6845
rect 16084 -6879 16153 -6845
rect 16187 -6879 16256 -6845
rect 16290 -6879 16310 -6845
rect 16344 -6843 16364 -6809
rect 16398 -6843 16463 -6809
rect 16497 -6843 16562 -6809
rect 16596 -6843 16674 -6809
rect 16344 -6913 16674 -6843
rect -950 -6953 -899 -6914
rect -1145 -7015 -1095 -6999
rect -1048 -6991 -984 -6975
rect -1249 -7023 -1183 -7022
rect -1048 -7025 -1034 -6991
rect -1000 -7025 -984 -6991
rect -1048 -7067 -984 -7025
rect -916 -6987 -899 -6953
rect -950 -7033 -899 -6987
rect -864 -6972 -162 -6913
rect -864 -7006 -846 -6972
rect -812 -7006 -214 -6972
rect -180 -7006 -162 -6972
rect -864 -7067 -162 -7006
rect -128 -6939 -70 -6922
rect -128 -6973 -116 -6939
rect -82 -6973 -70 -6939
rect -128 -7067 -70 -6973
rect -36 -6972 666 -6913
rect -36 -7006 -18 -6972
rect 16 -7006 614 -6972
rect 648 -7006 666 -6972
rect -36 -7067 666 -7006
rect 700 -6972 1402 -6913
rect 700 -7006 718 -6972
rect 752 -7006 1350 -6972
rect 1384 -7006 1402 -6972
rect 700 -7067 1402 -7006
rect 1436 -6939 1494 -6922
rect 1436 -6973 1448 -6939
rect 1482 -6973 1494 -6939
rect 1436 -7067 1494 -6973
rect 1528 -6972 2230 -6913
rect 1528 -7006 1546 -6972
rect 1580 -7006 2178 -6972
rect 2212 -7006 2230 -6972
rect 1528 -7067 2230 -7006
rect 2264 -6972 2966 -6913
rect 2264 -7006 2282 -6972
rect 2316 -7006 2914 -6972
rect 2948 -7006 2966 -6972
rect 2264 -7067 2966 -7006
rect 3000 -6939 3058 -6922
rect 3000 -6973 3012 -6939
rect 3046 -6973 3058 -6939
rect 3000 -7067 3058 -6973
rect 3092 -6972 3794 -6913
rect 3092 -7006 3110 -6972
rect 3144 -7006 3742 -6972
rect 3776 -7006 3794 -6972
rect 3092 -7067 3794 -7006
rect 3828 -6972 4530 -6913
rect 3828 -7006 3846 -6972
rect 3880 -7006 4478 -6972
rect 4512 -7006 4530 -6972
rect 3828 -7067 4530 -7006
rect 4564 -6939 4622 -6922
rect 4564 -6973 4576 -6939
rect 4610 -6973 4622 -6939
rect 4564 -7067 4622 -6973
rect 4656 -6972 5358 -6913
rect 4656 -7006 4674 -6972
rect 4708 -7006 5306 -6972
rect 5340 -7006 5358 -6972
rect 4656 -7067 5358 -7006
rect 5392 -6972 6094 -6913
rect 5392 -7006 5410 -6972
rect 5444 -7006 6042 -6972
rect 6076 -7006 6094 -6972
rect 5392 -7067 6094 -7006
rect 6128 -6939 6186 -6922
rect 6128 -6973 6140 -6939
rect 6174 -6973 6186 -6939
rect 6128 -7067 6186 -6973
rect 6220 -6972 6922 -6913
rect 6220 -7006 6238 -6972
rect 6272 -7006 6870 -6972
rect 6904 -7006 6922 -6972
rect 6220 -7067 6922 -7006
rect 6956 -6972 7658 -6913
rect 6956 -7006 6974 -6972
rect 7008 -7006 7606 -6972
rect 7640 -7006 7658 -6972
rect 6956 -7067 7658 -7006
rect 7692 -6939 7750 -6922
rect 7692 -6973 7704 -6939
rect 7738 -6973 7750 -6939
rect 7692 -7067 7750 -6973
rect 7784 -6972 8486 -6913
rect 7784 -7006 7802 -6972
rect 7836 -7006 8434 -6972
rect 8468 -7006 8486 -6972
rect 7784 -7067 8486 -7006
rect 8520 -6972 9222 -6913
rect 8520 -7006 8538 -6972
rect 8572 -7006 9170 -6972
rect 9204 -7006 9222 -6972
rect 8520 -7067 9222 -7006
rect 9256 -6939 9314 -6922
rect 9256 -6973 9268 -6939
rect 9302 -6973 9314 -6939
rect 9256 -7067 9314 -6973
rect 15880 -6939 15938 -6922
rect 15880 -6973 15892 -6939
rect 15926 -6973 15938 -6939
rect 15880 -7067 15938 -6973
rect 15972 -6972 16674 -6913
rect 15972 -7006 15990 -6972
rect 16024 -7006 16622 -6972
rect 16656 -7006 16674 -6972
rect 15972 -7067 16674 -7006
rect -2997 -7101 -2968 -7067
rect -2934 -7101 -2876 -7067
rect -2842 -7101 -2784 -7067
rect -2750 -7101 -2692 -7067
rect -2658 -7101 -2600 -7067
rect -2566 -7101 -2508 -7067
rect -2474 -7101 -2416 -7067
rect -2382 -7101 -2324 -7067
rect -2290 -7101 -2232 -7067
rect -2198 -7101 -2140 -7067
rect -2106 -7101 -2048 -7067
rect -2014 -7101 -1956 -7067
rect -1922 -7101 -1864 -7067
rect -1830 -7101 -1772 -7067
rect -1738 -7101 -1680 -7067
rect -1646 -7101 -1588 -7067
rect -1554 -7101 -1496 -7067
rect -1462 -7101 -1404 -7067
rect -1370 -7101 -1312 -7067
rect -1278 -7101 -1220 -7067
rect -1186 -7101 -1128 -7067
rect -1094 -7101 -1036 -7067
rect -1002 -7101 -944 -7067
rect -910 -7101 -852 -7067
rect -818 -7101 -760 -7067
rect -726 -7101 -668 -7067
rect -634 -7101 -576 -7067
rect -542 -7101 -484 -7067
rect -450 -7101 -392 -7067
rect -358 -7101 -300 -7067
rect -266 -7101 -208 -7067
rect -174 -7101 -116 -7067
rect -82 -7101 -24 -7067
rect 10 -7101 68 -7067
rect 102 -7101 160 -7067
rect 194 -7101 252 -7067
rect 286 -7101 344 -7067
rect 378 -7101 436 -7067
rect 470 -7101 528 -7067
rect 562 -7101 620 -7067
rect 654 -7101 712 -7067
rect 746 -7101 804 -7067
rect 838 -7101 896 -7067
rect 930 -7101 988 -7067
rect 1022 -7101 1080 -7067
rect 1114 -7101 1172 -7067
rect 1206 -7101 1264 -7067
rect 1298 -7101 1356 -7067
rect 1390 -7101 1448 -7067
rect 1482 -7101 1540 -7067
rect 1574 -7101 1632 -7067
rect 1666 -7101 1724 -7067
rect 1758 -7101 1816 -7067
rect 1850 -7101 1908 -7067
rect 1942 -7101 2000 -7067
rect 2034 -7101 2092 -7067
rect 2126 -7101 2184 -7067
rect 2218 -7101 2276 -7067
rect 2310 -7101 2368 -7067
rect 2402 -7101 2460 -7067
rect 2494 -7101 2552 -7067
rect 2586 -7101 2644 -7067
rect 2678 -7101 2736 -7067
rect 2770 -7101 2828 -7067
rect 2862 -7101 2920 -7067
rect 2954 -7101 3012 -7067
rect 3046 -7101 3104 -7067
rect 3138 -7101 3196 -7067
rect 3230 -7101 3288 -7067
rect 3322 -7101 3380 -7067
rect 3414 -7101 3472 -7067
rect 3506 -7101 3564 -7067
rect 3598 -7101 3656 -7067
rect 3690 -7101 3748 -7067
rect 3782 -7101 3840 -7067
rect 3874 -7101 3932 -7067
rect 3966 -7101 4024 -7067
rect 4058 -7101 4116 -7067
rect 4150 -7101 4208 -7067
rect 4242 -7101 4300 -7067
rect 4334 -7101 4392 -7067
rect 4426 -7101 4484 -7067
rect 4518 -7101 4576 -7067
rect 4610 -7101 4668 -7067
rect 4702 -7101 4760 -7067
rect 4794 -7101 4852 -7067
rect 4886 -7101 4944 -7067
rect 4978 -7101 5036 -7067
rect 5070 -7101 5128 -7067
rect 5162 -7101 5220 -7067
rect 5254 -7101 5312 -7067
rect 5346 -7101 5404 -7067
rect 5438 -7101 5496 -7067
rect 5530 -7101 5588 -7067
rect 5622 -7101 5680 -7067
rect 5714 -7101 5772 -7067
rect 5806 -7101 5864 -7067
rect 5898 -7101 5956 -7067
rect 5990 -7101 6048 -7067
rect 6082 -7101 6140 -7067
rect 6174 -7101 6232 -7067
rect 6266 -7101 6324 -7067
rect 6358 -7101 6416 -7067
rect 6450 -7101 6508 -7067
rect 6542 -7101 6600 -7067
rect 6634 -7101 6692 -7067
rect 6726 -7101 6784 -7067
rect 6818 -7101 6876 -7067
rect 6910 -7101 6968 -7067
rect 7002 -7101 7060 -7067
rect 7094 -7101 7152 -7067
rect 7186 -7101 7244 -7067
rect 7278 -7101 7336 -7067
rect 7370 -7101 7428 -7067
rect 7462 -7101 7520 -7067
rect 7554 -7101 7612 -7067
rect 7646 -7101 7704 -7067
rect 7738 -7101 7796 -7067
rect 7830 -7101 7888 -7067
rect 7922 -7101 7980 -7067
rect 8014 -7101 8072 -7067
rect 8106 -7101 8164 -7067
rect 8198 -7101 8256 -7067
rect 8290 -7101 8348 -7067
rect 8382 -7101 8440 -7067
rect 8474 -7101 8532 -7067
rect 8566 -7101 8624 -7067
rect 8658 -7101 8716 -7067
rect 8750 -7101 8808 -7067
rect 8842 -7101 8900 -7067
rect 8934 -7101 8992 -7067
rect 9026 -7101 9084 -7067
rect 9118 -7101 9176 -7067
rect 9210 -7101 9268 -7067
rect 9302 -7101 9360 -7067
rect 9394 -7101 9452 -7067
rect 9486 -7101 9544 -7067
rect 9578 -7101 9636 -7067
rect 9670 -7101 9728 -7067
rect 9762 -7101 9820 -7067
rect 9854 -7101 9912 -7067
rect 9946 -7101 10004 -7067
rect 10038 -7101 10096 -7067
rect 10130 -7101 10188 -7067
rect 10222 -7101 10280 -7067
rect 10314 -7101 10372 -7067
rect 10406 -7101 10464 -7067
rect 10498 -7101 10556 -7067
rect 10590 -7101 10648 -7067
rect 10682 -7101 10740 -7067
rect 10774 -7101 10832 -7067
rect 10866 -7101 10924 -7067
rect 10958 -7101 11016 -7067
rect 11050 -7101 11108 -7067
rect 11142 -7101 11200 -7067
rect 11234 -7101 11292 -7067
rect 11326 -7101 11384 -7067
rect 11418 -7101 11476 -7067
rect 11510 -7101 11568 -7067
rect 11602 -7101 11660 -7067
rect 11694 -7101 11752 -7067
rect 11786 -7101 11844 -7067
rect 11878 -7101 11936 -7067
rect 11970 -7101 12028 -7067
rect 12062 -7101 12120 -7067
rect 12154 -7101 12212 -7067
rect 12246 -7101 12304 -7067
rect 12338 -7101 12396 -7067
rect 12430 -7101 12488 -7067
rect 12522 -7101 12580 -7067
rect 12614 -7101 12672 -7067
rect 12706 -7101 12764 -7067
rect 12798 -7101 12856 -7067
rect 12890 -7101 12948 -7067
rect 12982 -7101 13040 -7067
rect 13074 -7101 13132 -7067
rect 13166 -7101 13224 -7067
rect 13258 -7101 13316 -7067
rect 13350 -7101 13408 -7067
rect 13442 -7101 13500 -7067
rect 13534 -7101 13592 -7067
rect 13626 -7101 13684 -7067
rect 13718 -7101 13776 -7067
rect 13810 -7101 13868 -7067
rect 13902 -7101 13960 -7067
rect 13994 -7101 14052 -7067
rect 14086 -7101 14144 -7067
rect 14178 -7101 14236 -7067
rect 14270 -7101 14328 -7067
rect 14362 -7101 14420 -7067
rect 14454 -7101 14512 -7067
rect 14546 -7101 14604 -7067
rect 14638 -7101 14696 -7067
rect 14730 -7101 14788 -7067
rect 14822 -7101 14880 -7067
rect 14914 -7101 14972 -7067
rect 15006 -7101 15064 -7067
rect 15098 -7101 15156 -7067
rect 15190 -7101 15248 -7067
rect 15282 -7101 15340 -7067
rect 15374 -7101 15432 -7067
rect 15466 -7101 15524 -7067
rect 15558 -7101 15616 -7067
rect 15650 -7101 15708 -7067
rect 15742 -7101 15800 -7067
rect 15834 -7101 15892 -7067
rect 15926 -7101 15984 -7067
rect 16018 -7101 16076 -7067
rect 16110 -7101 16168 -7067
rect 16202 -7101 16260 -7067
rect 16294 -7101 16352 -7067
rect 16386 -7101 16444 -7067
rect 16478 -7101 16536 -7067
rect 16570 -7101 16628 -7067
rect 16662 -7101 16691 -7067
rect -2980 -7162 -2278 -7101
rect -2980 -7196 -2962 -7162
rect -2928 -7196 -2330 -7162
rect -2296 -7196 -2278 -7162
rect -2980 -7255 -2278 -7196
rect -2244 -7195 -2186 -7101
rect -2244 -7229 -2232 -7195
rect -2198 -7229 -2186 -7195
rect -2244 -7246 -2186 -7229
rect -1600 -7162 -898 -7101
rect -1600 -7196 -1582 -7162
rect -1548 -7196 -950 -7162
rect -916 -7196 -898 -7162
rect -2980 -7323 -2902 -7289
rect -2868 -7323 -2799 -7289
rect -2765 -7323 -2696 -7289
rect -2662 -7323 -2642 -7289
rect -2980 -7393 -2642 -7323
rect -2608 -7325 -2278 -7255
rect -2608 -7359 -2588 -7325
rect -2554 -7359 -2489 -7325
rect -2455 -7359 -2390 -7325
rect -2356 -7359 -2278 -7325
rect -1600 -7255 -898 -7196
rect -864 -7162 -162 -7101
rect -864 -7196 -846 -7162
rect -812 -7196 -214 -7162
rect -180 -7196 -162 -7162
rect -864 -7255 -162 -7196
rect -128 -7195 -70 -7101
rect -128 -7229 -116 -7195
rect -82 -7229 -70 -7195
rect -128 -7246 -70 -7229
rect -36 -7162 666 -7101
rect -36 -7196 -18 -7162
rect 16 -7196 614 -7162
rect 648 -7196 666 -7162
rect -36 -7255 666 -7196
rect 700 -7162 1402 -7101
rect 700 -7196 718 -7162
rect 752 -7196 1350 -7162
rect 1384 -7196 1402 -7162
rect 700 -7255 1402 -7196
rect 1436 -7195 1494 -7101
rect 1436 -7229 1448 -7195
rect 1482 -7229 1494 -7195
rect 1436 -7246 1494 -7229
rect 1528 -7162 2230 -7101
rect 1528 -7196 1546 -7162
rect 1580 -7196 2178 -7162
rect 2212 -7196 2230 -7162
rect 1528 -7255 2230 -7196
rect 2264 -7169 2598 -7101
rect 2264 -7203 2282 -7169
rect 2316 -7203 2546 -7169
rect 2580 -7203 2598 -7169
rect 2264 -7255 2598 -7203
rect 2816 -7195 2874 -7101
rect 2816 -7229 2828 -7195
rect 2862 -7229 2874 -7195
rect 2908 -7152 2965 -7101
rect 2908 -7186 2931 -7152
rect 2908 -7202 2965 -7186
rect 2999 -7154 3064 -7135
rect 2999 -7188 3015 -7154
rect 3049 -7188 3064 -7154
rect 2816 -7246 2874 -7229
rect 2999 -7236 3064 -7188
rect -1600 -7325 -1270 -7255
rect -1600 -7359 -1522 -7325
rect -1488 -7359 -1423 -7325
rect -1389 -7359 -1324 -7325
rect -1290 -7359 -1270 -7325
rect -1236 -7323 -1216 -7289
rect -1182 -7323 -1113 -7289
rect -1079 -7323 -1010 -7289
rect -976 -7323 -898 -7289
rect -2980 -7433 -2278 -7393
rect -2980 -7467 -2962 -7433
rect -2928 -7467 -2330 -7433
rect -2296 -7467 -2278 -7433
rect -2980 -7535 -2278 -7467
rect -2980 -7569 -2962 -7535
rect -2928 -7569 -2330 -7535
rect -2296 -7569 -2278 -7535
rect -2980 -7611 -2278 -7569
rect -2244 -7413 -2186 -7378
rect -1236 -7393 -898 -7323
rect -864 -7325 -534 -7255
rect -864 -7359 -786 -7325
rect -752 -7359 -687 -7325
rect -653 -7359 -588 -7325
rect -554 -7359 -534 -7325
rect -500 -7323 -480 -7289
rect -446 -7323 -377 -7289
rect -343 -7323 -274 -7289
rect -240 -7323 -162 -7289
rect -500 -7393 -162 -7323
rect -36 -7325 294 -7255
rect -36 -7359 42 -7325
rect 76 -7359 141 -7325
rect 175 -7359 240 -7325
rect 274 -7359 294 -7325
rect 328 -7323 348 -7289
rect 382 -7323 451 -7289
rect 485 -7323 554 -7289
rect 588 -7323 666 -7289
rect -2244 -7447 -2232 -7413
rect -2198 -7447 -2186 -7413
rect -2244 -7506 -2186 -7447
rect -2244 -7540 -2232 -7506
rect -2198 -7540 -2186 -7506
rect -2244 -7611 -2186 -7540
rect -1600 -7433 -898 -7393
rect -1600 -7467 -1582 -7433
rect -1548 -7467 -950 -7433
rect -916 -7467 -898 -7433
rect -1600 -7535 -898 -7467
rect -1600 -7569 -1582 -7535
rect -1548 -7569 -950 -7535
rect -916 -7569 -898 -7535
rect -1600 -7611 -898 -7569
rect -864 -7433 -162 -7393
rect -864 -7467 -846 -7433
rect -812 -7467 -214 -7433
rect -180 -7467 -162 -7433
rect -864 -7535 -162 -7467
rect -864 -7569 -846 -7535
rect -812 -7569 -214 -7535
rect -180 -7569 -162 -7535
rect -864 -7611 -162 -7569
rect -128 -7413 -70 -7378
rect 328 -7393 666 -7323
rect 700 -7325 1030 -7255
rect 700 -7359 778 -7325
rect 812 -7359 877 -7325
rect 911 -7359 976 -7325
rect 1010 -7359 1030 -7325
rect 1064 -7323 1084 -7289
rect 1118 -7323 1187 -7289
rect 1221 -7323 1290 -7289
rect 1324 -7323 1402 -7289
rect 1064 -7393 1402 -7323
rect 1528 -7325 1858 -7255
rect 1528 -7359 1606 -7325
rect 1640 -7359 1705 -7325
rect 1739 -7359 1804 -7325
rect 1838 -7359 1858 -7325
rect 1892 -7323 1912 -7289
rect 1946 -7323 2015 -7289
rect 2049 -7323 2118 -7289
rect 2152 -7323 2230 -7289
rect -128 -7447 -116 -7413
rect -82 -7447 -70 -7413
rect -128 -7506 -70 -7447
rect -128 -7540 -116 -7506
rect -82 -7540 -70 -7506
rect -128 -7611 -70 -7540
rect -36 -7433 666 -7393
rect -36 -7467 -18 -7433
rect 16 -7467 614 -7433
rect 648 -7467 666 -7433
rect -36 -7535 666 -7467
rect -36 -7569 -18 -7535
rect 16 -7569 614 -7535
rect 648 -7569 666 -7535
rect -36 -7611 666 -7569
rect 700 -7433 1402 -7393
rect 700 -7467 718 -7433
rect 752 -7467 1350 -7433
rect 1384 -7467 1402 -7433
rect 700 -7535 1402 -7467
rect 700 -7569 718 -7535
rect 752 -7569 1350 -7535
rect 1384 -7569 1402 -7535
rect 700 -7611 1402 -7569
rect 1436 -7413 1494 -7378
rect 1892 -7393 2230 -7323
rect 1436 -7447 1448 -7413
rect 1482 -7447 1494 -7413
rect 1436 -7506 1494 -7447
rect 1436 -7540 1448 -7506
rect 1482 -7540 1494 -7506
rect 1436 -7611 1494 -7540
rect 1528 -7433 2230 -7393
rect 1528 -7467 1546 -7433
rect 1580 -7467 2178 -7433
rect 2212 -7467 2230 -7433
rect 1528 -7535 2230 -7467
rect 1528 -7569 1546 -7535
rect 1580 -7569 2178 -7535
rect 2212 -7569 2230 -7535
rect 1528 -7611 2230 -7569
rect 2264 -7323 2284 -7289
rect 2318 -7323 2414 -7289
rect 2264 -7393 2414 -7323
rect 2448 -7325 2598 -7255
rect 2448 -7359 2544 -7325
rect 2578 -7359 2598 -7325
rect 2908 -7270 3064 -7236
rect 2908 -7304 2934 -7270
rect 2968 -7304 3064 -7270
rect 2908 -7342 3064 -7304
rect 2264 -7433 2598 -7393
rect 2264 -7467 2282 -7433
rect 2316 -7467 2546 -7433
rect 2580 -7467 2598 -7433
rect 2264 -7535 2598 -7467
rect 2264 -7569 2282 -7535
rect 2316 -7569 2546 -7535
rect 2580 -7569 2598 -7535
rect 2264 -7611 2598 -7569
rect 2816 -7413 2874 -7378
rect 2816 -7447 2828 -7413
rect 2862 -7447 2874 -7413
rect 2816 -7506 2874 -7447
rect 2816 -7540 2828 -7506
rect 2862 -7540 2874 -7506
rect 2816 -7611 2874 -7540
rect 2908 -7433 2964 -7417
rect 2908 -7467 2930 -7433
rect 2908 -7535 2964 -7467
rect 2908 -7569 2930 -7535
rect 2908 -7611 2964 -7569
rect 2998 -7433 3064 -7342
rect 3102 -7191 3150 -7159
rect 3102 -7225 3111 -7191
rect 3145 -7225 3150 -7191
rect 3102 -7299 3150 -7225
rect 3184 -7195 3242 -7101
rect 3184 -7229 3196 -7195
rect 3230 -7229 3242 -7195
rect 3184 -7246 3242 -7229
rect 3276 -7169 3610 -7101
rect 3276 -7203 3294 -7169
rect 3328 -7203 3558 -7169
rect 3592 -7203 3610 -7169
rect 3276 -7255 3610 -7203
rect 3644 -7195 3702 -7101
rect 3644 -7229 3656 -7195
rect 3690 -7229 3702 -7195
rect 3644 -7246 3702 -7229
rect 3736 -7143 3798 -7101
rect 3736 -7177 3758 -7143
rect 3792 -7177 3798 -7143
rect 3736 -7211 3798 -7177
rect 3736 -7245 3758 -7211
rect 3792 -7245 3798 -7211
rect 3136 -7333 3150 -7299
rect 3102 -7349 3150 -7333
rect 3276 -7323 3296 -7289
rect 3330 -7323 3426 -7289
rect 3184 -7413 3242 -7378
rect 2998 -7467 3014 -7433
rect 3048 -7467 3064 -7433
rect 2998 -7535 3064 -7467
rect 2998 -7569 3014 -7535
rect 3048 -7569 3064 -7535
rect 2998 -7577 3064 -7569
rect 3098 -7433 3150 -7417
rect 3132 -7467 3150 -7433
rect 3098 -7535 3150 -7467
rect 3132 -7569 3150 -7535
rect 3098 -7611 3150 -7569
rect 3184 -7447 3196 -7413
rect 3230 -7447 3242 -7413
rect 3184 -7506 3242 -7447
rect 3184 -7540 3196 -7506
rect 3230 -7540 3242 -7506
rect 3184 -7611 3242 -7540
rect 3276 -7393 3426 -7323
rect 3460 -7325 3610 -7255
rect 3736 -7261 3798 -7245
rect 3839 -7143 3978 -7135
rect 3839 -7177 3926 -7143
rect 3960 -7177 3978 -7143
rect 3839 -7188 3978 -7177
rect 3839 -7222 3852 -7188
rect 3886 -7211 3978 -7188
rect 3886 -7222 3926 -7211
rect 3839 -7245 3926 -7222
rect 3960 -7245 3978 -7211
rect 3839 -7261 3978 -7245
rect 4012 -7195 4070 -7101
rect 4012 -7229 4024 -7195
rect 4058 -7229 4070 -7195
rect 4012 -7246 4070 -7229
rect 4104 -7169 4438 -7101
rect 4104 -7203 4122 -7169
rect 4156 -7203 4386 -7169
rect 4420 -7203 4438 -7169
rect 4104 -7255 4438 -7203
rect 4472 -7195 4530 -7101
rect 4472 -7229 4484 -7195
rect 4518 -7229 4530 -7195
rect 4472 -7246 4530 -7229
rect 4565 -7162 4616 -7135
rect 4565 -7196 4582 -7162
rect 4650 -7143 4716 -7101
rect 4650 -7177 4666 -7143
rect 4700 -7177 4716 -7143
rect 4650 -7181 4716 -7177
rect 4801 -7158 4907 -7135
rect 3460 -7359 3556 -7325
rect 3590 -7359 3610 -7325
rect 3738 -7299 3805 -7295
rect 3738 -7304 3755 -7299
rect 3738 -7338 3747 -7304
rect 3789 -7333 3805 -7299
rect 3781 -7338 3805 -7333
rect 3738 -7349 3805 -7338
rect 3276 -7433 3610 -7393
rect 3276 -7467 3294 -7433
rect 3328 -7467 3558 -7433
rect 3592 -7467 3610 -7433
rect 3276 -7535 3610 -7467
rect 3276 -7569 3294 -7535
rect 3328 -7569 3558 -7535
rect 3592 -7569 3610 -7535
rect 3276 -7611 3610 -7569
rect 3644 -7413 3702 -7378
rect 3839 -7381 3873 -7261
rect 3907 -7333 3923 -7299
rect 3957 -7305 3974 -7299
rect 3907 -7339 3928 -7333
rect 3962 -7339 3974 -7305
rect 3907 -7349 3974 -7339
rect 4104 -7323 4124 -7289
rect 4158 -7323 4254 -7289
rect 3644 -7447 3656 -7413
rect 3690 -7447 3702 -7413
rect 3644 -7506 3702 -7447
rect 3644 -7540 3656 -7506
rect 3690 -7540 3702 -7506
rect 3644 -7611 3702 -7540
rect 3736 -7399 3792 -7383
rect 3736 -7433 3758 -7399
rect 3736 -7467 3792 -7433
rect 3736 -7501 3758 -7467
rect 3736 -7535 3792 -7501
rect 3736 -7569 3758 -7535
rect 3736 -7611 3792 -7569
rect 3826 -7399 3892 -7381
rect 3826 -7433 3842 -7399
rect 3876 -7433 3892 -7399
rect 3826 -7467 3892 -7433
rect 3826 -7501 3842 -7467
rect 3876 -7501 3892 -7467
rect 3826 -7535 3892 -7501
rect 3826 -7569 3842 -7535
rect 3876 -7569 3892 -7535
rect 3826 -7577 3892 -7569
rect 3926 -7399 3978 -7383
rect 3960 -7433 3978 -7399
rect 3926 -7467 3978 -7433
rect 3960 -7501 3978 -7467
rect 3926 -7535 3978 -7501
rect 3960 -7569 3978 -7535
rect 3926 -7611 3978 -7569
rect 4012 -7413 4070 -7378
rect 4012 -7447 4024 -7413
rect 4058 -7447 4070 -7413
rect 4012 -7506 4070 -7447
rect 4012 -7540 4024 -7506
rect 4058 -7540 4070 -7506
rect 4012 -7611 4070 -7540
rect 4104 -7393 4254 -7323
rect 4288 -7325 4438 -7255
rect 4288 -7359 4384 -7325
rect 4418 -7359 4438 -7325
rect 4565 -7249 4616 -7196
rect 4801 -7192 4873 -7158
rect 4801 -7208 4907 -7192
rect 4945 -7204 5000 -7135
rect 4801 -7215 4836 -7208
rect 4650 -7249 4836 -7215
rect 4945 -7238 4955 -7204
rect 4989 -7238 5000 -7204
rect 4565 -7304 4599 -7249
rect 4650 -7283 4684 -7249
rect 4104 -7433 4438 -7393
rect 4104 -7467 4122 -7433
rect 4156 -7467 4386 -7433
rect 4420 -7467 4438 -7433
rect 4104 -7535 4438 -7467
rect 4104 -7569 4122 -7535
rect 4156 -7569 4386 -7535
rect 4420 -7569 4438 -7535
rect 4104 -7611 4438 -7569
rect 4472 -7413 4530 -7378
rect 4472 -7447 4484 -7413
rect 4518 -7447 4530 -7413
rect 4472 -7506 4530 -7447
rect 4472 -7540 4484 -7506
rect 4518 -7540 4530 -7506
rect 4472 -7611 4530 -7540
rect 4565 -7383 4599 -7338
rect 4633 -7299 4684 -7283
rect 4667 -7333 4684 -7299
rect 4633 -7349 4684 -7333
rect 4729 -7299 4768 -7283
rect 4763 -7333 4768 -7299
rect 4729 -7349 4768 -7333
rect 4565 -7399 4632 -7383
rect 4565 -7433 4582 -7399
rect 4616 -7433 4632 -7399
rect 4565 -7467 4632 -7433
rect 4565 -7501 4582 -7467
rect 4616 -7501 4632 -7467
rect 4565 -7535 4632 -7501
rect 4565 -7569 4582 -7535
rect 4616 -7569 4632 -7535
rect 4565 -7577 4632 -7569
rect 4666 -7399 4700 -7383
rect 4666 -7467 4700 -7433
rect 4666 -7535 4700 -7501
rect 4666 -7611 4700 -7569
rect 4734 -7543 4768 -7349
rect 4802 -7475 4836 -7249
rect 4870 -7263 4904 -7247
rect 4870 -7407 4904 -7297
rect 4945 -7263 5000 -7238
rect 4945 -7297 4966 -7263
rect 4945 -7367 5000 -7297
rect 5034 -7306 5072 -7135
rect 5108 -7158 5210 -7101
rect 5142 -7192 5176 -7158
rect 5108 -7208 5210 -7192
rect 5254 -7158 5303 -7142
rect 5254 -7192 5260 -7158
rect 5294 -7192 5303 -7158
rect 5254 -7263 5303 -7192
rect 5392 -7195 5450 -7101
rect 5392 -7229 5404 -7195
rect 5438 -7229 5450 -7195
rect 5392 -7246 5450 -7229
rect 5484 -7169 5818 -7101
rect 5484 -7203 5502 -7169
rect 5536 -7203 5766 -7169
rect 5800 -7203 5818 -7169
rect 5484 -7255 5818 -7203
rect 5852 -7195 5910 -7101
rect 5852 -7229 5864 -7195
rect 5898 -7229 5910 -7195
rect 5852 -7246 5910 -7229
rect 5945 -7181 5996 -7135
rect 5945 -7215 5962 -7181
rect 6030 -7143 6094 -7101
rect 6030 -7177 6046 -7143
rect 6080 -7177 6094 -7143
rect 6229 -7146 6295 -7145
rect 6030 -7193 6094 -7177
rect 6141 -7169 6191 -7153
rect 5112 -7297 5128 -7263
rect 5162 -7297 5358 -7263
rect 5034 -7340 5036 -7306
rect 5070 -7340 5072 -7306
rect 5034 -7376 5072 -7340
rect 5034 -7407 5038 -7376
rect 4870 -7410 5038 -7407
rect 4870 -7441 5072 -7410
rect 5106 -7373 5256 -7372
rect 5106 -7407 5171 -7373
rect 5205 -7376 5256 -7373
rect 5205 -7407 5206 -7376
rect 5106 -7410 5206 -7407
rect 5240 -7410 5256 -7376
rect 4802 -7509 4902 -7475
rect 4936 -7509 4977 -7475
rect 5011 -7509 5027 -7475
rect 5106 -7543 5140 -7410
rect 5290 -7459 5358 -7297
rect 5484 -7323 5504 -7289
rect 5538 -7323 5634 -7289
rect 4734 -7577 5140 -7543
rect 5174 -7475 5208 -7459
rect 5174 -7611 5208 -7509
rect 5255 -7475 5358 -7459
rect 5255 -7509 5260 -7475
rect 5294 -7509 5358 -7475
rect 5255 -7541 5358 -7509
rect 5392 -7413 5450 -7378
rect 5392 -7447 5404 -7413
rect 5438 -7447 5450 -7413
rect 5392 -7506 5450 -7447
rect 5392 -7540 5404 -7506
rect 5438 -7540 5450 -7506
rect 5392 -7611 5450 -7540
rect 5484 -7393 5634 -7323
rect 5668 -7325 5818 -7255
rect 5668 -7359 5764 -7325
rect 5798 -7359 5818 -7325
rect 5945 -7266 5996 -7215
rect 6175 -7203 6191 -7169
rect 6141 -7207 6191 -7203
rect 5484 -7433 5818 -7393
rect 5484 -7467 5502 -7433
rect 5536 -7467 5766 -7433
rect 5800 -7467 5818 -7433
rect 5484 -7535 5818 -7467
rect 5484 -7569 5502 -7535
rect 5536 -7569 5766 -7535
rect 5800 -7569 5818 -7535
rect 5484 -7611 5818 -7569
rect 5852 -7413 5910 -7378
rect 5852 -7447 5864 -7413
rect 5898 -7447 5910 -7413
rect 5852 -7506 5910 -7447
rect 5852 -7540 5864 -7506
rect 5898 -7540 5910 -7506
rect 5852 -7611 5910 -7540
rect 5945 -7380 5992 -7266
rect 6141 -7283 6181 -7207
rect 6229 -7232 6245 -7146
rect 6026 -7299 6181 -7283
rect 6060 -7333 6181 -7299
rect 6026 -7349 6181 -7333
rect 5945 -7393 6012 -7380
rect 5945 -7427 5962 -7393
rect 5996 -7427 6012 -7393
rect 5945 -7464 6012 -7427
rect 5945 -7498 5962 -7464
rect 5996 -7498 6012 -7464
rect 5945 -7535 6012 -7498
rect 5945 -7569 5962 -7535
rect 5996 -7569 6012 -7535
rect 5945 -7577 6012 -7569
rect 6046 -7399 6089 -7383
rect 6080 -7433 6089 -7399
rect 6046 -7467 6089 -7433
rect 6080 -7501 6089 -7467
rect 6046 -7535 6089 -7501
rect 6080 -7569 6089 -7535
rect 6046 -7611 6089 -7569
rect 6127 -7427 6181 -7349
rect 6215 -7248 6245 -7232
rect 6279 -7248 6295 -7146
rect 6329 -7173 6363 -7101
rect 6329 -7223 6363 -7207
rect 6397 -7178 6413 -7144
rect 6447 -7178 6463 -7144
rect 6397 -7212 6463 -7178
rect 6516 -7157 6558 -7101
rect 6921 -7151 6995 -7101
rect 6516 -7191 6519 -7157
rect 6553 -7191 6558 -7157
rect 6516 -7207 6558 -7191
rect 6613 -7191 6717 -7157
rect 6751 -7191 6770 -7157
rect 6804 -7191 6820 -7157
rect 6854 -7191 6885 -7157
rect 6215 -7249 6295 -7248
rect 6397 -7246 6413 -7212
rect 6447 -7246 6463 -7212
rect 6397 -7249 6463 -7246
rect 6215 -7257 6264 -7249
rect 6215 -7373 6253 -7257
rect 6397 -7283 6437 -7249
rect 6613 -7283 6647 -7191
rect 6287 -7299 6437 -7283
rect 6321 -7333 6437 -7299
rect 6287 -7349 6437 -7333
rect 6471 -7299 6647 -7283
rect 6505 -7333 6647 -7299
rect 6471 -7349 6647 -7333
rect 6215 -7383 6262 -7373
rect 6215 -7393 6297 -7383
rect 6215 -7399 6247 -7393
rect 6231 -7427 6247 -7399
rect 6281 -7427 6297 -7393
rect 6399 -7390 6437 -7349
rect 6399 -7393 6579 -7390
rect 6127 -7467 6193 -7427
rect 6127 -7501 6143 -7467
rect 6177 -7501 6193 -7467
rect 6127 -7535 6193 -7501
rect 6127 -7569 6143 -7535
rect 6177 -7569 6193 -7535
rect 6231 -7461 6297 -7427
rect 6231 -7495 6247 -7461
rect 6281 -7495 6297 -7461
rect 6231 -7529 6297 -7495
rect 6231 -7563 6247 -7529
rect 6281 -7563 6297 -7529
rect 6231 -7568 6297 -7563
rect 6331 -7425 6365 -7409
rect 6331 -7505 6365 -7459
rect 6127 -7573 6193 -7569
rect 6331 -7611 6365 -7539
rect 6399 -7427 6417 -7393
rect 6451 -7415 6579 -7393
rect 6451 -7427 6545 -7415
rect 6399 -7449 6545 -7427
rect 6399 -7464 6579 -7449
rect 6399 -7498 6417 -7464
rect 6451 -7465 6579 -7464
rect 6451 -7498 6467 -7465
rect 6399 -7535 6467 -7498
rect 6399 -7569 6417 -7535
rect 6451 -7569 6467 -7535
rect 6399 -7577 6467 -7569
rect 6514 -7527 6577 -7511
rect 6514 -7561 6541 -7527
rect 6575 -7561 6577 -7527
rect 6613 -7517 6647 -7349
rect 6681 -7241 6774 -7225
rect 6681 -7275 6740 -7241
rect 6681 -7291 6774 -7275
rect 6851 -7237 6885 -7191
rect 6921 -7185 6939 -7151
rect 6973 -7185 6995 -7151
rect 7334 -7143 7384 -7101
rect 6921 -7201 6995 -7185
rect 7059 -7191 7138 -7157
rect 7172 -7191 7194 -7157
rect 7233 -7191 7249 -7157
rect 7283 -7191 7300 -7157
rect 6851 -7253 7017 -7237
rect 6851 -7287 6983 -7253
rect 6681 -7373 6745 -7291
rect 6851 -7297 7017 -7287
rect 6681 -7407 6694 -7373
rect 6728 -7407 6745 -7373
rect 6681 -7415 6745 -7407
rect 6715 -7449 6745 -7415
rect 6681 -7483 6745 -7449
rect 6779 -7349 6817 -7333
rect 6779 -7383 6783 -7349
rect 6779 -7441 6817 -7383
rect 6779 -7475 6781 -7441
rect 6815 -7475 6817 -7441
rect 6779 -7477 6817 -7475
rect 6851 -7511 6885 -7297
rect 6977 -7303 7017 -7297
rect 6919 -7347 6953 -7333
rect 7059 -7347 7093 -7191
rect 7266 -7219 7300 -7191
rect 7368 -7177 7384 -7143
rect 7506 -7143 7572 -7101
rect 7334 -7193 7384 -7177
rect 7435 -7169 7472 -7153
rect 7435 -7203 7438 -7169
rect 7506 -7177 7522 -7143
rect 7556 -7177 7572 -7143
rect 7606 -7169 7640 -7153
rect 6919 -7349 7093 -7347
rect 6953 -7381 7093 -7349
rect 7127 -7241 7232 -7231
rect 7127 -7275 7182 -7241
rect 7216 -7275 7232 -7241
rect 7266 -7245 7311 -7219
rect 6953 -7383 7021 -7381
rect 6919 -7399 7021 -7383
rect 6613 -7551 6740 -7517
rect 6774 -7551 6790 -7517
rect 6835 -7527 6885 -7511
rect 6514 -7611 6577 -7561
rect 6869 -7561 6885 -7527
rect 6835 -7577 6885 -7561
rect 6919 -7467 6953 -7451
rect 6919 -7535 6953 -7501
rect 6987 -7522 7021 -7399
rect 7055 -7449 7093 -7415
rect 7127 -7441 7161 -7275
rect 7195 -7337 7243 -7309
rect 7195 -7371 7202 -7337
rect 7236 -7371 7243 -7337
rect 7195 -7373 7243 -7371
rect 7195 -7407 7198 -7373
rect 7232 -7407 7243 -7373
rect 7195 -7428 7243 -7407
rect 7055 -7475 7095 -7449
rect 7129 -7475 7161 -7441
rect 7277 -7466 7311 -7245
rect 7345 -7264 7401 -7227
rect 7345 -7298 7356 -7264
rect 7390 -7298 7401 -7264
rect 7345 -7367 7401 -7298
rect 7379 -7401 7401 -7367
rect 7345 -7417 7401 -7401
rect 7435 -7373 7472 -7203
rect 7606 -7211 7640 -7203
rect 7435 -7407 7436 -7373
rect 7470 -7407 7472 -7373
rect 7055 -7488 7161 -7475
rect 7250 -7492 7311 -7466
rect 7435 -7459 7472 -7407
rect 6987 -7556 7158 -7522
rect 7192 -7556 7208 -7522
rect 7250 -7527 7300 -7492
rect 7435 -7493 7438 -7459
rect 7507 -7245 7640 -7211
rect 7692 -7195 7750 -7101
rect 7692 -7229 7704 -7195
rect 7738 -7229 7750 -7195
rect 7507 -7314 7553 -7245
rect 7692 -7246 7750 -7229
rect 7784 -7162 8486 -7101
rect 7784 -7196 7802 -7162
rect 7836 -7196 8434 -7162
rect 8468 -7196 8486 -7162
rect 7784 -7255 8486 -7196
rect 8520 -7162 9222 -7101
rect 8520 -7196 8538 -7162
rect 8572 -7196 9170 -7162
rect 9204 -7196 9222 -7162
rect 8520 -7255 9222 -7196
rect 9256 -7195 9314 -7101
rect 9256 -7229 9268 -7195
rect 9302 -7229 9314 -7195
rect 9256 -7246 9314 -7229
rect 15880 -7195 15938 -7101
rect 15880 -7229 15892 -7195
rect 15926 -7229 15938 -7195
rect 15880 -7246 15938 -7229
rect 15972 -7162 16674 -7101
rect 15972 -7196 15990 -7162
rect 16024 -7196 16622 -7162
rect 16656 -7196 16674 -7162
rect 15972 -7255 16674 -7196
rect 7541 -7348 7553 -7314
rect 7507 -7441 7553 -7348
rect 7587 -7290 7657 -7279
rect 7587 -7324 7604 -7290
rect 7638 -7299 7657 -7290
rect 7587 -7333 7609 -7324
rect 7643 -7333 7657 -7299
rect 7587 -7364 7657 -7333
rect 7784 -7325 8114 -7255
rect 7784 -7359 7862 -7325
rect 7896 -7359 7961 -7325
rect 7995 -7359 8060 -7325
rect 8094 -7359 8114 -7325
rect 8148 -7323 8168 -7289
rect 8202 -7323 8271 -7289
rect 8305 -7323 8374 -7289
rect 8408 -7323 8486 -7289
rect 7587 -7398 7605 -7364
rect 7639 -7398 7657 -7364
rect 7587 -7409 7657 -7398
rect 7507 -7475 7515 -7441
rect 7549 -7443 7553 -7441
rect 7692 -7413 7750 -7378
rect 8148 -7393 8486 -7323
rect 8520 -7325 8850 -7255
rect 8520 -7359 8598 -7325
rect 8632 -7359 8697 -7325
rect 8731 -7359 8796 -7325
rect 8830 -7359 8850 -7325
rect 8884 -7323 8904 -7289
rect 8938 -7323 9007 -7289
rect 9041 -7323 9110 -7289
rect 9144 -7323 9222 -7289
rect 8884 -7393 9222 -7323
rect 15972 -7325 16302 -7255
rect 15972 -7359 16050 -7325
rect 16084 -7359 16149 -7325
rect 16183 -7359 16248 -7325
rect 16282 -7359 16302 -7325
rect 16336 -7323 16356 -7289
rect 16390 -7323 16459 -7289
rect 16493 -7323 16562 -7289
rect 16596 -7323 16674 -7289
rect 7549 -7459 7640 -7443
rect 7549 -7475 7606 -7459
rect 7507 -7477 7606 -7475
rect 6919 -7611 6953 -7569
rect 7284 -7561 7300 -7527
rect 7250 -7577 7300 -7561
rect 7334 -7535 7387 -7519
rect 7368 -7569 7387 -7535
rect 7334 -7611 7387 -7569
rect 7435 -7527 7472 -7493
rect 7435 -7561 7438 -7527
rect 7435 -7577 7472 -7561
rect 7506 -7545 7522 -7511
rect 7556 -7545 7572 -7511
rect 7506 -7611 7572 -7545
rect 7606 -7527 7640 -7493
rect 7606 -7577 7640 -7561
rect 7692 -7447 7704 -7413
rect 7738 -7447 7750 -7413
rect 7692 -7506 7750 -7447
rect 7692 -7540 7704 -7506
rect 7738 -7540 7750 -7506
rect 7692 -7611 7750 -7540
rect 7784 -7433 8486 -7393
rect 7784 -7467 7802 -7433
rect 7836 -7467 8434 -7433
rect 8468 -7467 8486 -7433
rect 7784 -7535 8486 -7467
rect 7784 -7569 7802 -7535
rect 7836 -7569 8434 -7535
rect 8468 -7569 8486 -7535
rect 7784 -7611 8486 -7569
rect 8520 -7433 9222 -7393
rect 8520 -7467 8538 -7433
rect 8572 -7467 9170 -7433
rect 9204 -7467 9222 -7433
rect 8520 -7535 9222 -7467
rect 8520 -7569 8538 -7535
rect 8572 -7569 9170 -7535
rect 9204 -7569 9222 -7535
rect 8520 -7611 9222 -7569
rect 9256 -7413 9314 -7378
rect 9256 -7447 9268 -7413
rect 9302 -7447 9314 -7413
rect 9256 -7506 9314 -7447
rect 9256 -7540 9268 -7506
rect 9302 -7540 9314 -7506
rect 9256 -7611 9314 -7540
rect 15880 -7413 15938 -7378
rect 16336 -7393 16674 -7323
rect 15880 -7447 15892 -7413
rect 15926 -7447 15938 -7413
rect 15880 -7506 15938 -7447
rect 15880 -7540 15892 -7506
rect 15926 -7540 15938 -7506
rect 15880 -7611 15938 -7540
rect 15972 -7433 16674 -7393
rect 15972 -7467 15990 -7433
rect 16024 -7467 16622 -7433
rect 16656 -7467 16674 -7433
rect 15972 -7535 16674 -7467
rect 15972 -7569 15990 -7535
rect 16024 -7569 16622 -7535
rect 16656 -7569 16674 -7535
rect 15972 -7611 16674 -7569
rect -2997 -7645 -2968 -7611
rect -2934 -7645 -2876 -7611
rect -2842 -7645 -2784 -7611
rect -2750 -7645 -2692 -7611
rect -2658 -7645 -2600 -7611
rect -2566 -7645 -2508 -7611
rect -2474 -7645 -2416 -7611
rect -2382 -7645 -2324 -7611
rect -2290 -7645 -2232 -7611
rect -2198 -7645 -2140 -7611
rect -2106 -7645 -2048 -7611
rect -2014 -7645 -1956 -7611
rect -1922 -7645 -1864 -7611
rect -1830 -7645 -1772 -7611
rect -1738 -7645 -1680 -7611
rect -1646 -7645 -1588 -7611
rect -1554 -7645 -1496 -7611
rect -1462 -7645 -1404 -7611
rect -1370 -7645 -1312 -7611
rect -1278 -7645 -1220 -7611
rect -1186 -7645 -1128 -7611
rect -1094 -7645 -1036 -7611
rect -1002 -7645 -944 -7611
rect -910 -7645 -852 -7611
rect -818 -7645 -760 -7611
rect -726 -7645 -668 -7611
rect -634 -7645 -576 -7611
rect -542 -7645 -484 -7611
rect -450 -7645 -392 -7611
rect -358 -7645 -300 -7611
rect -266 -7645 -208 -7611
rect -174 -7645 -116 -7611
rect -82 -7645 -24 -7611
rect 10 -7645 68 -7611
rect 102 -7645 160 -7611
rect 194 -7645 252 -7611
rect 286 -7645 344 -7611
rect 378 -7645 436 -7611
rect 470 -7645 528 -7611
rect 562 -7645 620 -7611
rect 654 -7645 712 -7611
rect 746 -7645 804 -7611
rect 838 -7645 896 -7611
rect 930 -7645 988 -7611
rect 1022 -7645 1080 -7611
rect 1114 -7645 1172 -7611
rect 1206 -7645 1264 -7611
rect 1298 -7645 1356 -7611
rect 1390 -7645 1448 -7611
rect 1482 -7645 1540 -7611
rect 1574 -7645 1632 -7611
rect 1666 -7645 1724 -7611
rect 1758 -7645 1816 -7611
rect 1850 -7645 1908 -7611
rect 1942 -7645 2000 -7611
rect 2034 -7645 2092 -7611
rect 2126 -7645 2184 -7611
rect 2218 -7645 2276 -7611
rect 2310 -7645 2368 -7611
rect 2402 -7645 2460 -7611
rect 2494 -7645 2552 -7611
rect 2586 -7645 2644 -7611
rect 2678 -7645 2736 -7611
rect 2770 -7645 2828 -7611
rect 2862 -7645 2920 -7611
rect 2954 -7645 3012 -7611
rect 3046 -7645 3104 -7611
rect 3138 -7645 3196 -7611
rect 3230 -7645 3288 -7611
rect 3322 -7645 3380 -7611
rect 3414 -7645 3472 -7611
rect 3506 -7645 3564 -7611
rect 3598 -7645 3656 -7611
rect 3690 -7645 3748 -7611
rect 3782 -7645 3840 -7611
rect 3874 -7645 3932 -7611
rect 3966 -7645 4024 -7611
rect 4058 -7645 4116 -7611
rect 4150 -7645 4208 -7611
rect 4242 -7645 4300 -7611
rect 4334 -7645 4392 -7611
rect 4426 -7645 4484 -7611
rect 4518 -7645 4576 -7611
rect 4610 -7645 4668 -7611
rect 4702 -7645 4760 -7611
rect 4794 -7645 4852 -7611
rect 4886 -7645 4944 -7611
rect 4978 -7645 5036 -7611
rect 5070 -7645 5128 -7611
rect 5162 -7645 5220 -7611
rect 5254 -7645 5312 -7611
rect 5346 -7645 5404 -7611
rect 5438 -7645 5496 -7611
rect 5530 -7645 5588 -7611
rect 5622 -7645 5680 -7611
rect 5714 -7645 5772 -7611
rect 5806 -7645 5864 -7611
rect 5898 -7645 5956 -7611
rect 5990 -7645 6048 -7611
rect 6082 -7645 6140 -7611
rect 6174 -7645 6232 -7611
rect 6266 -7645 6324 -7611
rect 6358 -7645 6416 -7611
rect 6450 -7645 6508 -7611
rect 6542 -7645 6600 -7611
rect 6634 -7645 6692 -7611
rect 6726 -7645 6784 -7611
rect 6818 -7645 6876 -7611
rect 6910 -7645 6968 -7611
rect 7002 -7645 7060 -7611
rect 7094 -7645 7152 -7611
rect 7186 -7645 7244 -7611
rect 7278 -7645 7336 -7611
rect 7370 -7645 7428 -7611
rect 7462 -7645 7520 -7611
rect 7554 -7645 7612 -7611
rect 7646 -7645 7704 -7611
rect 7738 -7645 7796 -7611
rect 7830 -7645 7888 -7611
rect 7922 -7645 7980 -7611
rect 8014 -7645 8072 -7611
rect 8106 -7645 8164 -7611
rect 8198 -7645 8256 -7611
rect 8290 -7645 8348 -7611
rect 8382 -7645 8440 -7611
rect 8474 -7645 8532 -7611
rect 8566 -7645 8624 -7611
rect 8658 -7645 8716 -7611
rect 8750 -7645 8808 -7611
rect 8842 -7645 8900 -7611
rect 8934 -7645 8992 -7611
rect 9026 -7645 9084 -7611
rect 9118 -7645 9176 -7611
rect 9210 -7645 9268 -7611
rect 9302 -7645 9360 -7611
rect 9394 -7645 9452 -7611
rect 9486 -7645 9544 -7611
rect 9578 -7645 9636 -7611
rect 9670 -7645 9728 -7611
rect 9762 -7645 9820 -7611
rect 9854 -7645 9912 -7611
rect 9946 -7645 10004 -7611
rect 10038 -7645 10096 -7611
rect 10130 -7645 10188 -7611
rect 10222 -7645 10280 -7611
rect 10314 -7645 10372 -7611
rect 10406 -7645 10464 -7611
rect 10498 -7645 10556 -7611
rect 10590 -7645 10648 -7611
rect 10682 -7645 10740 -7611
rect 10774 -7645 10832 -7611
rect 10866 -7645 10924 -7611
rect 10958 -7645 11016 -7611
rect 11050 -7645 11108 -7611
rect 11142 -7645 11200 -7611
rect 11234 -7645 11292 -7611
rect 11326 -7645 11384 -7611
rect 11418 -7645 11476 -7611
rect 11510 -7645 11568 -7611
rect 11602 -7645 11660 -7611
rect 11694 -7645 11752 -7611
rect 11786 -7645 11844 -7611
rect 11878 -7645 11936 -7611
rect 11970 -7645 12028 -7611
rect 12062 -7645 12120 -7611
rect 12154 -7645 12212 -7611
rect 12246 -7645 12304 -7611
rect 12338 -7645 12396 -7611
rect 12430 -7645 12488 -7611
rect 12522 -7645 12580 -7611
rect 12614 -7645 12672 -7611
rect 12706 -7645 12764 -7611
rect 12798 -7645 12856 -7611
rect 12890 -7645 12948 -7611
rect 12982 -7645 13040 -7611
rect 13074 -7645 13132 -7611
rect 13166 -7645 13224 -7611
rect 13258 -7645 13316 -7611
rect 13350 -7645 13408 -7611
rect 13442 -7645 13500 -7611
rect 13534 -7645 13592 -7611
rect 13626 -7645 13684 -7611
rect 13718 -7645 13776 -7611
rect 13810 -7645 13868 -7611
rect 13902 -7645 13960 -7611
rect 13994 -7645 14052 -7611
rect 14086 -7645 14144 -7611
rect 14178 -7645 14236 -7611
rect 14270 -7645 14328 -7611
rect 14362 -7645 14420 -7611
rect 14454 -7645 14512 -7611
rect 14546 -7645 14604 -7611
rect 14638 -7645 14696 -7611
rect 14730 -7645 14788 -7611
rect 14822 -7645 14880 -7611
rect 14914 -7645 14972 -7611
rect 15006 -7645 15064 -7611
rect 15098 -7645 15156 -7611
rect 15190 -7645 15248 -7611
rect 15282 -7645 15340 -7611
rect 15374 -7645 15432 -7611
rect 15466 -7645 15524 -7611
rect 15558 -7645 15616 -7611
rect 15650 -7645 15708 -7611
rect 15742 -7645 15800 -7611
rect 15834 -7645 15892 -7611
rect 15926 -7645 15984 -7611
rect 16018 -7645 16076 -7611
rect 16110 -7645 16168 -7611
rect 16202 -7645 16260 -7611
rect 16294 -7645 16352 -7611
rect 16386 -7645 16444 -7611
rect 16478 -7645 16536 -7611
rect 16570 -7645 16628 -7611
rect 16662 -7645 16691 -7611
rect -2980 -7687 -2278 -7645
rect -2980 -7721 -2962 -7687
rect -2928 -7721 -2330 -7687
rect -2296 -7721 -2278 -7687
rect -2980 -7789 -2278 -7721
rect -2980 -7823 -2962 -7789
rect -2928 -7823 -2330 -7789
rect -2296 -7823 -2278 -7789
rect -2980 -7863 -2278 -7823
rect -2980 -7931 -2902 -7897
rect -2868 -7931 -2803 -7897
rect -2769 -7931 -2704 -7897
rect -2670 -7931 -2650 -7897
rect -2980 -8001 -2650 -7931
rect -2616 -7933 -2278 -7863
rect -2244 -7716 -2186 -7645
rect -2244 -7750 -2232 -7716
rect -2198 -7750 -2186 -7716
rect -2244 -7809 -2186 -7750
rect -2244 -7843 -2232 -7809
rect -2198 -7843 -2186 -7809
rect -2244 -7878 -2186 -7843
rect -1416 -7687 -1082 -7645
rect -1416 -7721 -1398 -7687
rect -1364 -7721 -1134 -7687
rect -1100 -7721 -1082 -7687
rect -1416 -7789 -1082 -7721
rect -1416 -7823 -1398 -7789
rect -1364 -7823 -1134 -7789
rect -1100 -7823 -1082 -7789
rect -1416 -7863 -1082 -7823
rect -2616 -7967 -2596 -7933
rect -2562 -7967 -2493 -7933
rect -2459 -7967 -2390 -7933
rect -2356 -7967 -2278 -7933
rect -1416 -7931 -1396 -7897
rect -1362 -7931 -1266 -7897
rect -1416 -8001 -1266 -7931
rect -1232 -7933 -1082 -7863
rect -1048 -7716 -990 -7645
rect -1048 -7750 -1036 -7716
rect -1002 -7750 -990 -7716
rect -1048 -7809 -990 -7750
rect -1048 -7843 -1036 -7809
rect -1002 -7843 -990 -7809
rect -1048 -7878 -990 -7843
rect -956 -7687 -900 -7645
rect -956 -7721 -934 -7687
rect -956 -7755 -900 -7721
rect -956 -7789 -934 -7755
rect -956 -7823 -900 -7789
rect -956 -7857 -934 -7823
rect -956 -7873 -900 -7857
rect -866 -7687 -800 -7679
rect -866 -7721 -850 -7687
rect -816 -7721 -800 -7687
rect -866 -7755 -800 -7721
rect -866 -7789 -850 -7755
rect -816 -7789 -800 -7755
rect -866 -7823 -800 -7789
rect -866 -7857 -850 -7823
rect -816 -7857 -800 -7823
rect -866 -7875 -800 -7857
rect -766 -7687 -714 -7645
rect -732 -7721 -714 -7687
rect -766 -7755 -714 -7721
rect -732 -7789 -714 -7755
rect -766 -7823 -714 -7789
rect -732 -7857 -714 -7823
rect -766 -7873 -714 -7857
rect -680 -7716 -622 -7645
rect -680 -7750 -668 -7716
rect -634 -7750 -622 -7716
rect -680 -7809 -622 -7750
rect -680 -7843 -668 -7809
rect -634 -7843 -622 -7809
rect -1232 -7967 -1136 -7933
rect -1102 -7967 -1082 -7933
rect -954 -7918 -887 -7907
rect -954 -7957 -937 -7918
rect -903 -7957 -887 -7918
rect -954 -7961 -887 -7957
rect -853 -7995 -819 -7875
rect -680 -7878 -622 -7843
rect -588 -7687 -254 -7645
rect -588 -7721 -570 -7687
rect -536 -7721 -306 -7687
rect -272 -7721 -254 -7687
rect -588 -7789 -254 -7721
rect -588 -7823 -570 -7789
rect -536 -7823 -306 -7789
rect -272 -7823 -254 -7789
rect -588 -7863 -254 -7823
rect -785 -7917 -718 -7907
rect -785 -7923 -762 -7917
rect -785 -7957 -769 -7923
rect -728 -7951 -718 -7917
rect -735 -7957 -718 -7951
rect -588 -7931 -568 -7897
rect -534 -7931 -438 -7897
rect -2980 -8060 -2278 -8001
rect -2980 -8094 -2962 -8060
rect -2928 -8094 -2330 -8060
rect -2296 -8094 -2278 -8060
rect -2980 -8155 -2278 -8094
rect -2244 -8027 -2186 -8010
rect -2244 -8061 -2232 -8027
rect -2198 -8061 -2186 -8027
rect -2244 -8155 -2186 -8061
rect -1416 -8053 -1082 -8001
rect -1416 -8087 -1398 -8053
rect -1364 -8087 -1134 -8053
rect -1100 -8087 -1082 -8053
rect -1416 -8155 -1082 -8087
rect -1048 -8027 -990 -8010
rect -1048 -8061 -1036 -8027
rect -1002 -8061 -990 -8027
rect -1048 -8155 -990 -8061
rect -956 -8011 -894 -7995
rect -956 -8045 -934 -8011
rect -900 -8045 -894 -8011
rect -956 -8079 -894 -8045
rect -956 -8113 -934 -8079
rect -900 -8113 -894 -8079
rect -956 -8155 -894 -8113
rect -853 -8011 -714 -7995
rect -588 -8001 -438 -7931
rect -404 -7933 -254 -7863
rect -220 -7716 -162 -7645
rect -220 -7750 -208 -7716
rect -174 -7750 -162 -7716
rect -220 -7809 -162 -7750
rect -220 -7843 -208 -7809
rect -174 -7843 -162 -7809
rect -128 -7694 -59 -7645
rect -128 -7728 -102 -7694
rect -68 -7728 -59 -7694
rect -128 -7762 -59 -7728
rect -128 -7796 -102 -7762
rect -68 -7796 -59 -7762
rect -128 -7812 -59 -7796
rect -24 -7701 27 -7685
rect -24 -7735 -16 -7701
rect 18 -7735 27 -7701
rect -24 -7789 27 -7735
rect -220 -7878 -162 -7843
rect -24 -7823 -16 -7789
rect 18 -7823 27 -7789
rect 61 -7694 113 -7645
rect 61 -7728 70 -7694
rect 104 -7728 113 -7694
rect 61 -7762 113 -7728
rect 61 -7796 70 -7762
rect 104 -7796 113 -7762
rect 61 -7812 113 -7796
rect 148 -7701 199 -7685
rect 148 -7735 156 -7701
rect 190 -7735 199 -7701
rect 148 -7789 199 -7735
rect -24 -7846 27 -7823
rect 148 -7823 156 -7789
rect 190 -7823 199 -7789
rect 233 -7694 285 -7645
rect 233 -7728 242 -7694
rect 276 -7728 285 -7694
rect 233 -7762 285 -7728
rect 233 -7796 242 -7762
rect 276 -7796 285 -7762
rect 233 -7812 285 -7796
rect 319 -7701 371 -7685
rect 319 -7735 328 -7701
rect 362 -7735 371 -7701
rect 319 -7789 371 -7735
rect 148 -7846 199 -7823
rect 319 -7823 328 -7789
rect 362 -7823 371 -7789
rect 405 -7694 482 -7645
rect 405 -7728 414 -7694
rect 448 -7728 482 -7694
rect 405 -7762 482 -7728
rect 405 -7796 414 -7762
rect 448 -7796 482 -7762
rect 405 -7812 482 -7796
rect 516 -7716 574 -7645
rect 516 -7750 528 -7716
rect 562 -7750 574 -7716
rect 516 -7809 574 -7750
rect 319 -7846 371 -7823
rect 516 -7843 528 -7809
rect 562 -7843 574 -7809
rect -404 -7967 -308 -7933
rect -274 -7967 -254 -7933
rect -124 -7880 482 -7846
rect 516 -7878 574 -7843
rect 608 -7687 942 -7645
rect 608 -7721 626 -7687
rect 660 -7721 890 -7687
rect 924 -7721 942 -7687
rect 608 -7789 942 -7721
rect 608 -7823 626 -7789
rect 660 -7823 890 -7789
rect 924 -7823 942 -7789
rect 608 -7863 942 -7823
rect -124 -7993 -90 -7880
rect -56 -7923 387 -7914
rect -56 -7957 -30 -7923
rect 4 -7957 38 -7923
rect 72 -7957 106 -7923
rect 140 -7957 174 -7923
rect 208 -7957 242 -7923
rect 276 -7957 310 -7923
rect 344 -7957 387 -7923
rect -56 -7959 387 -7957
rect 422 -7961 482 -7880
rect 422 -7993 434 -7961
rect -124 -7995 434 -7993
rect 468 -7995 482 -7961
rect -853 -8028 -766 -8011
rect -853 -8062 -848 -8028
rect -814 -8062 -769 -8028
rect -732 -8045 -714 -8011
rect -735 -8062 -714 -8045
rect -853 -8079 -714 -8062
rect -853 -8113 -766 -8079
rect -732 -8113 -714 -8079
rect -853 -8121 -714 -8113
rect -680 -8027 -622 -8010
rect -680 -8061 -668 -8027
rect -634 -8061 -622 -8027
rect -680 -8155 -622 -8061
rect -588 -8053 -254 -8001
rect -588 -8087 -570 -8053
rect -536 -8087 -306 -8053
rect -272 -8087 -254 -8053
rect -588 -8155 -254 -8087
rect -220 -8027 -162 -8010
rect -124 -8027 482 -7995
rect 608 -7931 628 -7897
rect 662 -7931 758 -7897
rect 608 -8001 758 -7931
rect 792 -7933 942 -7863
rect 976 -7716 1034 -7645
rect 976 -7750 988 -7716
rect 1022 -7750 1034 -7716
rect 976 -7809 1034 -7750
rect 976 -7843 988 -7809
rect 1022 -7843 1034 -7809
rect 1068 -7687 1120 -7645
rect 1068 -7721 1086 -7687
rect 1068 -7789 1120 -7721
rect 1068 -7823 1086 -7789
rect 1068 -7839 1120 -7823
rect 1154 -7687 1220 -7679
rect 1154 -7721 1170 -7687
rect 1204 -7721 1220 -7687
rect 1154 -7789 1220 -7721
rect 1154 -7823 1170 -7789
rect 1204 -7823 1220 -7789
rect 976 -7878 1034 -7843
rect 792 -7967 888 -7933
rect 922 -7967 942 -7933
rect 1068 -7923 1116 -7907
rect 1068 -7928 1082 -7923
rect 1068 -7962 1076 -7928
rect 1110 -7962 1116 -7957
rect 1068 -8001 1116 -7962
rect 516 -8027 574 -8010
rect -220 -8061 -208 -8027
rect -174 -8061 -162 -8027
rect -220 -8155 -162 -8061
rect -32 -8077 27 -8061
rect -32 -8111 -16 -8077
rect 18 -8111 27 -8077
rect -32 -8155 27 -8111
rect 61 -8066 113 -8027
rect 61 -8100 70 -8066
rect 104 -8100 113 -8066
rect 61 -8116 113 -8100
rect 147 -8077 199 -8061
rect 147 -8111 156 -8077
rect 190 -8111 199 -8077
rect 147 -8155 199 -8111
rect 233 -8066 284 -8027
rect 516 -8061 528 -8027
rect 562 -8061 574 -8027
rect 233 -8100 242 -8066
rect 276 -8100 284 -8066
rect 233 -8116 284 -8100
rect 318 -8077 378 -8061
rect 318 -8111 328 -8077
rect 362 -8111 378 -8077
rect 318 -8155 378 -8111
rect 516 -8155 574 -8061
rect 608 -8053 942 -8001
rect 608 -8087 626 -8053
rect 660 -8087 890 -8053
rect 924 -8087 942 -8053
rect 608 -8155 942 -8087
rect 976 -8027 1034 -8010
rect 976 -8061 988 -8027
rect 1022 -8061 1034 -8027
rect 976 -8155 1034 -8061
rect 1068 -8035 1076 -8001
rect 1110 -8035 1116 -8001
rect 1068 -8097 1116 -8035
rect 1154 -7914 1220 -7823
rect 1254 -7687 1310 -7645
rect 1288 -7721 1310 -7687
rect 1254 -7789 1310 -7721
rect 1288 -7823 1310 -7789
rect 1254 -7839 1310 -7823
rect 1344 -7716 1402 -7645
rect 1344 -7750 1356 -7716
rect 1390 -7750 1402 -7716
rect 1344 -7809 1402 -7750
rect 1344 -7843 1356 -7809
rect 1390 -7843 1402 -7809
rect 1344 -7878 1402 -7843
rect 1436 -7687 1770 -7645
rect 1436 -7721 1454 -7687
rect 1488 -7721 1718 -7687
rect 1752 -7721 1770 -7687
rect 1436 -7789 1770 -7721
rect 1436 -7823 1454 -7789
rect 1488 -7823 1718 -7789
rect 1752 -7823 1770 -7789
rect 1436 -7863 1770 -7823
rect 1154 -7922 1310 -7914
rect 1154 -7956 1171 -7922
rect 1205 -7956 1263 -7922
rect 1297 -7956 1310 -7922
rect 1154 -8020 1310 -7956
rect 1436 -7931 1456 -7897
rect 1490 -7931 1586 -7897
rect 1436 -8001 1586 -7931
rect 1620 -7933 1770 -7863
rect 1804 -7716 1862 -7645
rect 1804 -7750 1816 -7716
rect 1850 -7750 1862 -7716
rect 1804 -7809 1862 -7750
rect 1804 -7843 1816 -7809
rect 1850 -7843 1862 -7809
rect 1804 -7878 1862 -7843
rect 1896 -7687 2230 -7645
rect 1896 -7721 1914 -7687
rect 1948 -7721 2178 -7687
rect 2212 -7721 2230 -7687
rect 1896 -7789 2230 -7721
rect 1896 -7823 1914 -7789
rect 1948 -7823 2178 -7789
rect 2212 -7823 2230 -7789
rect 1896 -7863 2230 -7823
rect 1620 -7967 1716 -7933
rect 1750 -7967 1770 -7933
rect 1896 -7931 1916 -7897
rect 1950 -7931 2046 -7897
rect 1896 -8001 2046 -7931
rect 2080 -7933 2230 -7863
rect 2264 -7716 2322 -7645
rect 2264 -7750 2276 -7716
rect 2310 -7750 2322 -7716
rect 2264 -7809 2322 -7750
rect 2264 -7843 2276 -7809
rect 2310 -7843 2322 -7809
rect 2264 -7878 2322 -7843
rect 2356 -7694 2425 -7679
rect 2356 -7728 2375 -7694
rect 2409 -7728 2425 -7694
rect 2356 -7762 2425 -7728
rect 2356 -7796 2375 -7762
rect 2409 -7796 2425 -7762
rect 2356 -7846 2425 -7796
rect 2459 -7694 2525 -7645
rect 2459 -7728 2475 -7694
rect 2509 -7728 2525 -7694
rect 2459 -7762 2525 -7728
rect 2459 -7796 2475 -7762
rect 2509 -7796 2525 -7762
rect 2459 -7812 2525 -7796
rect 2615 -7694 2685 -7679
rect 2615 -7728 2633 -7694
rect 2667 -7728 2685 -7694
rect 2615 -7762 2685 -7728
rect 2615 -7796 2633 -7762
rect 2667 -7796 2685 -7762
rect 2356 -7880 2550 -7846
rect 2480 -7909 2550 -7880
rect 2615 -7908 2685 -7796
rect 2737 -7695 2787 -7679
rect 2771 -7729 2787 -7695
rect 2737 -7763 2787 -7729
rect 2771 -7797 2787 -7763
rect 2737 -7839 2787 -7797
rect 2877 -7694 2943 -7645
rect 2877 -7728 2893 -7694
rect 2927 -7728 2943 -7694
rect 2877 -7762 2943 -7728
rect 2877 -7796 2893 -7762
rect 2927 -7796 2943 -7762
rect 2877 -7805 2943 -7796
rect 2977 -7695 3058 -7679
rect 2977 -7729 2991 -7695
rect 3025 -7729 3058 -7695
rect 2977 -7763 3058 -7729
rect 2977 -7797 2991 -7763
rect 3025 -7797 3058 -7763
rect 2977 -7834 3058 -7797
rect 2737 -7873 2855 -7839
rect 2821 -7907 2855 -7873
rect 2080 -7967 2176 -7933
rect 2210 -7967 2230 -7933
rect 2356 -7917 2446 -7914
rect 2356 -7951 2369 -7917
rect 2403 -7923 2446 -7917
rect 2356 -7957 2396 -7951
rect 2430 -7957 2446 -7923
rect 2480 -7923 2566 -7909
rect 2480 -7957 2516 -7923
rect 2550 -7957 2566 -7923
rect 2480 -7967 2566 -7957
rect 2615 -7923 2787 -7908
rect 2615 -7957 2737 -7923
rect 2771 -7957 2787 -7923
rect 2615 -7958 2787 -7957
rect 2821 -7923 2974 -7907
rect 2821 -7957 2937 -7923
rect 2971 -7957 2974 -7923
rect 2480 -7991 2550 -7967
rect 1154 -8068 1219 -8020
rect 1344 -8027 1402 -8010
rect 1154 -8102 1169 -8068
rect 1203 -8102 1219 -8068
rect 1154 -8121 1219 -8102
rect 1253 -8070 1310 -8054
rect 1287 -8104 1310 -8070
rect 1253 -8155 1310 -8104
rect 1344 -8061 1356 -8027
rect 1390 -8061 1402 -8027
rect 1344 -8155 1402 -8061
rect 1436 -8053 1770 -8001
rect 1436 -8087 1454 -8053
rect 1488 -8087 1718 -8053
rect 1752 -8087 1770 -8053
rect 1436 -8155 1770 -8087
rect 1804 -8027 1862 -8010
rect 1804 -8061 1816 -8027
rect 1850 -8061 1862 -8027
rect 1804 -8155 1862 -8061
rect 1896 -8053 2230 -8001
rect 1896 -8087 1914 -8053
rect 1948 -8087 2178 -8053
rect 2212 -8087 2230 -8053
rect 1896 -8155 2230 -8087
rect 2264 -8027 2322 -8010
rect 2264 -8061 2276 -8027
rect 2310 -8061 2322 -8027
rect 2264 -8155 2322 -8061
rect 2356 -8025 2550 -7991
rect 2356 -8068 2422 -8025
rect 2356 -8102 2375 -8068
rect 2409 -8102 2422 -8068
rect 2356 -8121 2422 -8102
rect 2456 -8068 2522 -8059
rect 2456 -8102 2472 -8068
rect 2506 -8102 2522 -8068
rect 2456 -8155 2522 -8102
rect 2615 -8068 2685 -7958
rect 2821 -7973 2974 -7957
rect 3008 -7918 3058 -7834
rect 3092 -7716 3150 -7645
rect 3092 -7750 3104 -7716
rect 3138 -7750 3150 -7716
rect 3092 -7809 3150 -7750
rect 3092 -7843 3104 -7809
rect 3138 -7843 3150 -7809
rect 3092 -7878 3150 -7843
rect 3184 -7687 3518 -7645
rect 3184 -7721 3202 -7687
rect 3236 -7721 3466 -7687
rect 3500 -7721 3518 -7687
rect 3184 -7789 3518 -7721
rect 3184 -7823 3202 -7789
rect 3236 -7823 3466 -7789
rect 3500 -7823 3518 -7789
rect 3184 -7863 3518 -7823
rect 3008 -7952 3015 -7918
rect 3049 -7952 3058 -7918
rect 2821 -7992 2855 -7973
rect 2615 -8102 2632 -8068
rect 2666 -8102 2685 -8068
rect 2615 -8121 2685 -8102
rect 2737 -8026 2855 -7992
rect 2737 -8068 2787 -8026
rect 3008 -8044 3058 -7952
rect 3184 -7931 3204 -7897
rect 3238 -7931 3334 -7897
rect 3184 -8001 3334 -7931
rect 3368 -7933 3518 -7863
rect 3552 -7716 3610 -7645
rect 3552 -7750 3564 -7716
rect 3598 -7750 3610 -7716
rect 3552 -7809 3610 -7750
rect 3552 -7843 3564 -7809
rect 3598 -7843 3610 -7809
rect 3552 -7878 3610 -7843
rect 4380 -7687 5449 -7645
rect 4380 -7721 4398 -7687
rect 4432 -7721 5398 -7687
rect 5432 -7721 5449 -7687
rect 4380 -7789 5449 -7721
rect 4380 -7823 4398 -7789
rect 4432 -7823 5398 -7789
rect 5432 -7823 5449 -7789
rect 4380 -7863 5449 -7823
rect 3368 -7967 3464 -7933
rect 3498 -7967 3518 -7933
rect 4380 -7931 4458 -7897
rect 4492 -7931 4586 -7897
rect 4620 -7931 4714 -7897
rect 4748 -7931 4842 -7897
rect 4876 -7931 4896 -7897
rect 4380 -8001 4896 -7931
rect 4930 -7933 5449 -7863
rect 6312 -7716 6370 -7645
rect 6312 -7750 6324 -7716
rect 6358 -7750 6370 -7716
rect 6312 -7809 6370 -7750
rect 6312 -7843 6324 -7809
rect 6358 -7843 6370 -7809
rect 6312 -7878 6370 -7843
rect 6404 -7687 6738 -7645
rect 6404 -7721 6422 -7687
rect 6456 -7721 6686 -7687
rect 6720 -7721 6738 -7687
rect 6404 -7789 6738 -7721
rect 6404 -7823 6422 -7789
rect 6456 -7823 6686 -7789
rect 6720 -7823 6738 -7789
rect 6404 -7863 6738 -7823
rect 4930 -7967 4950 -7933
rect 4984 -7967 5078 -7933
rect 5112 -7967 5206 -7933
rect 5240 -7967 5334 -7933
rect 5368 -7967 5449 -7933
rect 6404 -7931 6424 -7897
rect 6458 -7931 6554 -7897
rect 6404 -8001 6554 -7931
rect 6588 -7933 6738 -7863
rect 6772 -7716 6830 -7645
rect 6772 -7750 6784 -7716
rect 6818 -7750 6830 -7716
rect 6772 -7809 6830 -7750
rect 6772 -7843 6784 -7809
rect 6818 -7843 6830 -7809
rect 6772 -7878 6830 -7843
rect 6864 -7694 6933 -7679
rect 6864 -7728 6883 -7694
rect 6917 -7728 6933 -7694
rect 6864 -7762 6933 -7728
rect 6864 -7796 6883 -7762
rect 6917 -7796 6933 -7762
rect 6864 -7846 6933 -7796
rect 6967 -7694 7033 -7645
rect 6967 -7728 6983 -7694
rect 7017 -7728 7033 -7694
rect 6967 -7762 7033 -7728
rect 6967 -7796 6983 -7762
rect 7017 -7796 7033 -7762
rect 6967 -7812 7033 -7796
rect 7123 -7694 7193 -7679
rect 7123 -7728 7141 -7694
rect 7175 -7728 7193 -7694
rect 7123 -7762 7193 -7728
rect 7123 -7796 7141 -7762
rect 7175 -7796 7193 -7762
rect 6864 -7880 7058 -7846
rect 6988 -7909 7058 -7880
rect 7123 -7908 7193 -7796
rect 7245 -7695 7295 -7679
rect 7279 -7729 7295 -7695
rect 7245 -7763 7295 -7729
rect 7279 -7797 7295 -7763
rect 7245 -7839 7295 -7797
rect 7385 -7694 7451 -7645
rect 7385 -7728 7401 -7694
rect 7435 -7728 7451 -7694
rect 7385 -7762 7451 -7728
rect 7385 -7796 7401 -7762
rect 7435 -7796 7451 -7762
rect 7385 -7805 7451 -7796
rect 7485 -7695 7566 -7679
rect 7485 -7729 7499 -7695
rect 7533 -7729 7566 -7695
rect 7485 -7763 7566 -7729
rect 7485 -7797 7499 -7763
rect 7533 -7797 7566 -7763
rect 7485 -7834 7566 -7797
rect 7245 -7873 7363 -7839
rect 7329 -7907 7363 -7873
rect 6588 -7967 6684 -7933
rect 6718 -7967 6738 -7933
rect 6864 -7918 6954 -7914
rect 6864 -7952 6876 -7918
rect 6910 -7923 6954 -7918
rect 6864 -7957 6904 -7952
rect 6938 -7957 6954 -7923
rect 6988 -7923 7074 -7909
rect 6988 -7957 7024 -7923
rect 7058 -7957 7074 -7923
rect 6988 -7967 7074 -7957
rect 7123 -7923 7295 -7908
rect 7123 -7957 7245 -7923
rect 7279 -7957 7295 -7923
rect 7123 -7958 7295 -7957
rect 7329 -7923 7482 -7907
rect 7329 -7957 7445 -7923
rect 7479 -7957 7482 -7923
rect 6988 -7991 7058 -7967
rect 2771 -8102 2787 -8068
rect 2737 -8121 2787 -8102
rect 2877 -8068 2943 -8052
rect 2877 -8102 2893 -8068
rect 2927 -8102 2943 -8068
rect 2877 -8155 2943 -8102
rect 2977 -8068 3058 -8044
rect 2977 -8102 2991 -8068
rect 3025 -8102 3058 -8068
rect 2977 -8121 3058 -8102
rect 3092 -8027 3150 -8010
rect 3092 -8061 3104 -8027
rect 3138 -8061 3150 -8027
rect 3092 -8155 3150 -8061
rect 3184 -8053 3518 -8001
rect 3184 -8087 3202 -8053
rect 3236 -8087 3466 -8053
rect 3500 -8087 3518 -8053
rect 3184 -8155 3518 -8087
rect 3552 -8027 3610 -8010
rect 3552 -8061 3564 -8027
rect 3598 -8061 3610 -8027
rect 3552 -8155 3610 -8061
rect 4380 -8060 5449 -8001
rect 4380 -8094 4398 -8060
rect 4432 -8094 5398 -8060
rect 5432 -8094 5449 -8060
rect 4380 -8155 5449 -8094
rect 6312 -8027 6370 -8010
rect 6312 -8061 6324 -8027
rect 6358 -8061 6370 -8027
rect 6312 -8155 6370 -8061
rect 6404 -8053 6738 -8001
rect 6404 -8087 6422 -8053
rect 6456 -8087 6686 -8053
rect 6720 -8087 6738 -8053
rect 6404 -8155 6738 -8087
rect 6772 -8027 6830 -8010
rect 6772 -8061 6784 -8027
rect 6818 -8061 6830 -8027
rect 6772 -8155 6830 -8061
rect 6864 -8025 7058 -7991
rect 6864 -8068 6930 -8025
rect 6864 -8102 6883 -8068
rect 6917 -8102 6930 -8068
rect 6864 -8121 6930 -8102
rect 6964 -8068 7030 -8059
rect 6964 -8102 6980 -8068
rect 7014 -8102 7030 -8068
rect 6964 -8155 7030 -8102
rect 7123 -8068 7193 -7958
rect 7329 -7973 7482 -7957
rect 7516 -7918 7566 -7834
rect 7600 -7716 7658 -7645
rect 7600 -7750 7612 -7716
rect 7646 -7750 7658 -7716
rect 7600 -7809 7658 -7750
rect 7600 -7843 7612 -7809
rect 7646 -7843 7658 -7809
rect 7600 -7878 7658 -7843
rect 7692 -7687 8026 -7645
rect 7692 -7721 7710 -7687
rect 7744 -7721 7974 -7687
rect 8008 -7721 8026 -7687
rect 7692 -7789 8026 -7721
rect 7692 -7823 7710 -7789
rect 7744 -7823 7974 -7789
rect 8008 -7823 8026 -7789
rect 7692 -7863 8026 -7823
rect 7516 -7952 7522 -7918
rect 7556 -7952 7566 -7918
rect 7329 -7992 7363 -7973
rect 7123 -8102 7140 -8068
rect 7174 -8102 7193 -8068
rect 7123 -8121 7193 -8102
rect 7245 -8026 7363 -7992
rect 7245 -8068 7295 -8026
rect 7516 -8044 7566 -7952
rect 7692 -7931 7712 -7897
rect 7746 -7931 7842 -7897
rect 7692 -8001 7842 -7931
rect 7876 -7933 8026 -7863
rect 8060 -7716 8118 -7645
rect 8060 -7750 8072 -7716
rect 8106 -7750 8118 -7716
rect 8060 -7809 8118 -7750
rect 8060 -7843 8072 -7809
rect 8106 -7843 8118 -7809
rect 8060 -7878 8118 -7843
rect 8152 -7694 8221 -7679
rect 8152 -7728 8171 -7694
rect 8205 -7728 8221 -7694
rect 8152 -7762 8221 -7728
rect 8152 -7796 8171 -7762
rect 8205 -7796 8221 -7762
rect 8152 -7846 8221 -7796
rect 8255 -7694 8321 -7645
rect 8255 -7728 8271 -7694
rect 8305 -7728 8321 -7694
rect 8255 -7762 8321 -7728
rect 8255 -7796 8271 -7762
rect 8305 -7796 8321 -7762
rect 8255 -7812 8321 -7796
rect 8411 -7694 8481 -7679
rect 8411 -7728 8429 -7694
rect 8463 -7728 8481 -7694
rect 8411 -7762 8481 -7728
rect 8411 -7796 8429 -7762
rect 8463 -7796 8481 -7762
rect 8152 -7880 8346 -7846
rect 8276 -7909 8346 -7880
rect 8411 -7908 8481 -7796
rect 8533 -7695 8583 -7679
rect 8567 -7729 8583 -7695
rect 8533 -7763 8583 -7729
rect 8567 -7797 8583 -7763
rect 8533 -7839 8583 -7797
rect 8673 -7694 8739 -7645
rect 8673 -7728 8689 -7694
rect 8723 -7728 8739 -7694
rect 8673 -7762 8739 -7728
rect 8673 -7796 8689 -7762
rect 8723 -7796 8739 -7762
rect 8673 -7805 8739 -7796
rect 8773 -7695 8854 -7679
rect 8773 -7729 8787 -7695
rect 8821 -7729 8854 -7695
rect 8773 -7763 8854 -7729
rect 8773 -7797 8787 -7763
rect 8821 -7797 8854 -7763
rect 8773 -7834 8854 -7797
rect 8533 -7873 8651 -7839
rect 8617 -7907 8651 -7873
rect 7876 -7967 7972 -7933
rect 8006 -7967 8026 -7933
rect 8152 -7919 8242 -7914
rect 8152 -7953 8164 -7919
rect 8198 -7923 8242 -7919
rect 8152 -7957 8192 -7953
rect 8226 -7957 8242 -7923
rect 8276 -7923 8362 -7909
rect 8276 -7957 8312 -7923
rect 8346 -7957 8362 -7923
rect 8276 -7967 8362 -7957
rect 8411 -7923 8583 -7908
rect 8411 -7957 8533 -7923
rect 8567 -7957 8583 -7923
rect 8411 -7958 8583 -7957
rect 8617 -7923 8770 -7907
rect 8617 -7957 8733 -7923
rect 8767 -7957 8770 -7923
rect 8276 -7991 8346 -7967
rect 7279 -8102 7295 -8068
rect 7245 -8121 7295 -8102
rect 7385 -8068 7451 -8052
rect 7385 -8102 7401 -8068
rect 7435 -8102 7451 -8068
rect 7385 -8155 7451 -8102
rect 7485 -8068 7566 -8044
rect 7485 -8102 7499 -8068
rect 7533 -8102 7566 -8068
rect 7485 -8121 7566 -8102
rect 7600 -8027 7658 -8010
rect 7600 -8061 7612 -8027
rect 7646 -8061 7658 -8027
rect 7600 -8155 7658 -8061
rect 7692 -8053 8026 -8001
rect 7692 -8087 7710 -8053
rect 7744 -8087 7974 -8053
rect 8008 -8087 8026 -8053
rect 7692 -8155 8026 -8087
rect 8060 -8027 8118 -8010
rect 8060 -8061 8072 -8027
rect 8106 -8061 8118 -8027
rect 8060 -8155 8118 -8061
rect 8152 -8025 8346 -7991
rect 8152 -8068 8218 -8025
rect 8152 -8102 8171 -8068
rect 8205 -8102 8218 -8068
rect 8152 -8121 8218 -8102
rect 8252 -8068 8318 -8059
rect 8252 -8102 8268 -8068
rect 8302 -8102 8318 -8068
rect 8252 -8155 8318 -8102
rect 8411 -8068 8481 -7958
rect 8617 -7973 8770 -7957
rect 8804 -7917 8854 -7834
rect 8888 -7716 8946 -7645
rect 8888 -7750 8900 -7716
rect 8934 -7750 8946 -7716
rect 8888 -7809 8946 -7750
rect 8888 -7843 8900 -7809
rect 8934 -7843 8946 -7809
rect 8888 -7878 8946 -7843
rect 8980 -7687 9314 -7645
rect 8980 -7721 8998 -7687
rect 9032 -7721 9262 -7687
rect 9296 -7721 9314 -7687
rect 8980 -7789 9314 -7721
rect 8980 -7823 8998 -7789
rect 9032 -7823 9262 -7789
rect 9296 -7823 9314 -7789
rect 8980 -7863 9314 -7823
rect 8804 -7951 8811 -7917
rect 8845 -7951 8854 -7917
rect 8617 -7992 8651 -7973
rect 8411 -8102 8428 -8068
rect 8462 -8102 8481 -8068
rect 8411 -8121 8481 -8102
rect 8533 -8026 8651 -7992
rect 8533 -8068 8583 -8026
rect 8804 -8044 8854 -7951
rect 8980 -7931 9000 -7897
rect 9034 -7931 9130 -7897
rect 8980 -8001 9130 -7931
rect 9164 -7933 9314 -7863
rect 9348 -7716 9406 -7645
rect 9348 -7750 9360 -7716
rect 9394 -7750 9406 -7716
rect 9348 -7809 9406 -7750
rect 9348 -7843 9360 -7809
rect 9394 -7843 9406 -7809
rect 9348 -7878 9406 -7843
rect 9440 -7694 9509 -7679
rect 9440 -7728 9459 -7694
rect 9493 -7728 9509 -7694
rect 9440 -7762 9509 -7728
rect 9440 -7796 9459 -7762
rect 9493 -7796 9509 -7762
rect 9440 -7846 9509 -7796
rect 9543 -7694 9609 -7645
rect 9543 -7728 9559 -7694
rect 9593 -7728 9609 -7694
rect 9543 -7762 9609 -7728
rect 9543 -7796 9559 -7762
rect 9593 -7796 9609 -7762
rect 9543 -7812 9609 -7796
rect 9699 -7694 9769 -7679
rect 9699 -7728 9717 -7694
rect 9751 -7728 9769 -7694
rect 9699 -7762 9769 -7728
rect 9699 -7796 9717 -7762
rect 9751 -7796 9769 -7762
rect 9440 -7880 9634 -7846
rect 9564 -7909 9634 -7880
rect 9699 -7908 9769 -7796
rect 9821 -7695 9871 -7679
rect 9855 -7729 9871 -7695
rect 9821 -7763 9871 -7729
rect 9855 -7797 9871 -7763
rect 9821 -7839 9871 -7797
rect 9961 -7694 10027 -7645
rect 9961 -7728 9977 -7694
rect 10011 -7728 10027 -7694
rect 9961 -7762 10027 -7728
rect 9961 -7796 9977 -7762
rect 10011 -7796 10027 -7762
rect 9961 -7805 10027 -7796
rect 10061 -7695 10142 -7679
rect 10061 -7729 10075 -7695
rect 10109 -7729 10142 -7695
rect 10061 -7763 10142 -7729
rect 10061 -7797 10075 -7763
rect 10109 -7797 10142 -7763
rect 10061 -7834 10142 -7797
rect 9821 -7873 9939 -7839
rect 9905 -7907 9939 -7873
rect 9164 -7967 9260 -7933
rect 9294 -7967 9314 -7933
rect 9440 -7917 9530 -7914
rect 9440 -7951 9453 -7917
rect 9487 -7923 9530 -7917
rect 9440 -7957 9480 -7951
rect 9514 -7957 9530 -7923
rect 9564 -7923 9650 -7909
rect 9564 -7957 9600 -7923
rect 9634 -7957 9650 -7923
rect 9564 -7967 9650 -7957
rect 9699 -7923 9871 -7908
rect 9699 -7957 9821 -7923
rect 9855 -7957 9871 -7923
rect 9699 -7958 9871 -7957
rect 9905 -7923 10058 -7907
rect 9905 -7957 10021 -7923
rect 10055 -7957 10058 -7923
rect 9564 -7991 9634 -7967
rect 8567 -8102 8583 -8068
rect 8533 -8121 8583 -8102
rect 8673 -8068 8739 -8052
rect 8673 -8102 8689 -8068
rect 8723 -8102 8739 -8068
rect 8673 -8155 8739 -8102
rect 8773 -8068 8854 -8044
rect 8773 -8102 8787 -8068
rect 8821 -8102 8854 -8068
rect 8773 -8121 8854 -8102
rect 8888 -8027 8946 -8010
rect 8888 -8061 8900 -8027
rect 8934 -8061 8946 -8027
rect 8888 -8155 8946 -8061
rect 8980 -8053 9314 -8001
rect 8980 -8087 8998 -8053
rect 9032 -8087 9262 -8053
rect 9296 -8087 9314 -8053
rect 8980 -8155 9314 -8087
rect 9348 -8027 9406 -8010
rect 9348 -8061 9360 -8027
rect 9394 -8061 9406 -8027
rect 9348 -8155 9406 -8061
rect 9440 -8025 9634 -7991
rect 9440 -8068 9506 -8025
rect 9440 -8102 9459 -8068
rect 9493 -8102 9506 -8068
rect 9440 -8121 9506 -8102
rect 9540 -8068 9606 -8059
rect 9540 -8102 9556 -8068
rect 9590 -8102 9606 -8068
rect 9540 -8155 9606 -8102
rect 9699 -8068 9769 -7958
rect 9905 -7973 10058 -7957
rect 10092 -7916 10142 -7834
rect 10176 -7716 10234 -7645
rect 10176 -7750 10188 -7716
rect 10222 -7750 10234 -7716
rect 10176 -7809 10234 -7750
rect 10176 -7843 10188 -7809
rect 10222 -7843 10234 -7809
rect 10176 -7878 10234 -7843
rect 10268 -7687 10602 -7645
rect 10268 -7721 10286 -7687
rect 10320 -7721 10550 -7687
rect 10584 -7721 10602 -7687
rect 10268 -7789 10602 -7721
rect 10268 -7823 10286 -7789
rect 10320 -7823 10550 -7789
rect 10584 -7823 10602 -7789
rect 10268 -7863 10602 -7823
rect 10092 -7950 10099 -7916
rect 10133 -7950 10142 -7916
rect 9905 -7992 9939 -7973
rect 9699 -8102 9716 -8068
rect 9750 -8102 9769 -8068
rect 9699 -8121 9769 -8102
rect 9821 -8026 9939 -7992
rect 9821 -8068 9871 -8026
rect 10092 -8044 10142 -7950
rect 10268 -7931 10288 -7897
rect 10322 -7931 10418 -7897
rect 10268 -8001 10418 -7931
rect 10452 -7933 10602 -7863
rect 10636 -7716 10694 -7645
rect 10636 -7750 10648 -7716
rect 10682 -7750 10694 -7716
rect 10636 -7809 10694 -7750
rect 10636 -7843 10648 -7809
rect 10682 -7843 10694 -7809
rect 10636 -7878 10694 -7843
rect 10729 -7687 10780 -7645
rect 10729 -7721 10746 -7687
rect 10729 -7755 10780 -7721
rect 10729 -7789 10746 -7755
rect 10729 -7823 10780 -7789
rect 10729 -7857 10746 -7823
rect 10729 -7873 10780 -7857
rect 10814 -7687 10880 -7679
rect 10814 -7721 10830 -7687
rect 10864 -7721 10880 -7687
rect 10814 -7755 10880 -7721
rect 10814 -7789 10830 -7755
rect 10864 -7789 10880 -7755
rect 10814 -7823 10880 -7789
rect 10914 -7687 10948 -7645
rect 10914 -7755 10948 -7721
rect 10914 -7805 10948 -7789
rect 10982 -7687 11048 -7679
rect 10982 -7721 10998 -7687
rect 11032 -7721 11048 -7687
rect 10982 -7755 11048 -7721
rect 10982 -7789 10998 -7755
rect 11032 -7789 11048 -7755
rect 10814 -7857 10830 -7823
rect 10864 -7839 10880 -7823
rect 10982 -7823 11048 -7789
rect 11082 -7687 11116 -7645
rect 11082 -7755 11116 -7721
rect 11082 -7805 11116 -7789
rect 11150 -7687 11216 -7679
rect 11150 -7721 11166 -7687
rect 11200 -7721 11216 -7687
rect 11150 -7755 11216 -7721
rect 11150 -7789 11166 -7755
rect 11200 -7789 11216 -7755
rect 10982 -7839 10998 -7823
rect 10864 -7857 10998 -7839
rect 11032 -7839 11048 -7823
rect 11150 -7823 11216 -7789
rect 11250 -7687 11284 -7645
rect 11250 -7755 11284 -7721
rect 11250 -7805 11284 -7789
rect 11318 -7687 11384 -7679
rect 11318 -7721 11334 -7687
rect 11368 -7721 11384 -7687
rect 11318 -7755 11384 -7721
rect 11318 -7789 11334 -7755
rect 11368 -7789 11384 -7755
rect 11150 -7839 11166 -7823
rect 11032 -7857 11166 -7839
rect 11200 -7839 11216 -7823
rect 11318 -7823 11384 -7789
rect 11418 -7687 11468 -7645
rect 11452 -7721 11468 -7687
rect 11418 -7755 11468 -7721
rect 11452 -7789 11468 -7755
rect 11418 -7805 11468 -7789
rect 11556 -7716 11614 -7645
rect 11556 -7750 11568 -7716
rect 11602 -7750 11614 -7716
rect 11318 -7839 11334 -7823
rect 11200 -7857 11334 -7839
rect 11368 -7857 11384 -7823
rect 10814 -7873 11384 -7857
rect 11556 -7809 11614 -7750
rect 11556 -7843 11568 -7809
rect 11602 -7843 11614 -7809
rect 11093 -7884 11200 -7873
rect 11556 -7878 11614 -7843
rect 11648 -7687 11982 -7645
rect 11648 -7721 11666 -7687
rect 11700 -7721 11930 -7687
rect 11964 -7721 11982 -7687
rect 11648 -7789 11982 -7721
rect 11648 -7823 11666 -7789
rect 11700 -7823 11930 -7789
rect 11964 -7823 11982 -7789
rect 11648 -7863 11982 -7823
rect 10452 -7967 10548 -7933
rect 10582 -7967 10602 -7933
rect 10733 -7917 11057 -7907
rect 10733 -7951 10741 -7917
rect 10775 -7923 10832 -7917
rect 10866 -7918 11057 -7917
rect 10866 -7923 10925 -7918
rect 10959 -7923 11017 -7918
rect 10733 -7957 10749 -7951
rect 10783 -7957 10830 -7923
rect 10866 -7951 10914 -7923
rect 10864 -7957 10914 -7951
rect 10959 -7952 10998 -7923
rect 11051 -7952 11057 -7918
rect 10948 -7957 10998 -7952
rect 11032 -7957 11057 -7952
rect 11093 -7918 11129 -7884
rect 11163 -7918 11200 -7884
rect 11093 -7957 11200 -7918
rect 11234 -7915 11522 -7907
rect 11234 -7957 11250 -7915
rect 11284 -7923 11344 -7915
rect 11284 -7957 11334 -7923
rect 11378 -7949 11522 -7915
rect 11368 -7957 11522 -7949
rect 11648 -7931 11668 -7897
rect 11702 -7931 11798 -7897
rect 9855 -8102 9871 -8068
rect 9821 -8121 9871 -8102
rect 9961 -8068 10027 -8052
rect 9961 -8102 9977 -8068
rect 10011 -8102 10027 -8068
rect 9961 -8155 10027 -8102
rect 10061 -8068 10142 -8044
rect 10061 -8102 10075 -8068
rect 10109 -8102 10142 -8068
rect 10061 -8121 10142 -8102
rect 10176 -8027 10234 -8010
rect 10176 -8061 10188 -8027
rect 10222 -8061 10234 -8027
rect 10176 -8155 10234 -8061
rect 10268 -8053 10602 -8001
rect 10268 -8087 10286 -8053
rect 10320 -8087 10550 -8053
rect 10584 -8087 10602 -8053
rect 10268 -8155 10602 -8087
rect 10636 -8027 10694 -8010
rect 10636 -8061 10648 -8027
rect 10682 -8061 10694 -8027
rect 10636 -8155 10694 -8061
rect 10729 -8011 11116 -7991
rect 10729 -8045 10746 -8011
rect 10780 -8029 10914 -8011
rect 10780 -8045 10796 -8029
rect 10729 -8079 10796 -8045
rect 10898 -8045 10914 -8029
rect 10948 -8029 11082 -8011
rect 10948 -8045 10964 -8029
rect 10729 -8113 10746 -8079
rect 10780 -8113 10796 -8079
rect 10729 -8121 10796 -8113
rect 10830 -8079 10864 -8063
rect 10830 -8155 10864 -8113
rect 10898 -8079 10964 -8045
rect 11066 -8045 11082 -8029
rect 11150 -8011 11200 -7957
rect 11418 -8011 11468 -7995
rect 11648 -8001 11798 -7931
rect 11832 -7933 11982 -7863
rect 13488 -7716 13546 -7645
rect 13488 -7750 13500 -7716
rect 13534 -7750 13546 -7716
rect 13488 -7809 13546 -7750
rect 13488 -7843 13500 -7809
rect 13534 -7843 13546 -7809
rect 13488 -7878 13546 -7843
rect 13580 -7687 14649 -7645
rect 13580 -7721 13598 -7687
rect 13632 -7721 14598 -7687
rect 14632 -7721 14649 -7687
rect 13580 -7789 14649 -7721
rect 13580 -7823 13598 -7789
rect 13632 -7823 14598 -7789
rect 14632 -7823 14649 -7789
rect 13580 -7863 14649 -7823
rect 11832 -7967 11928 -7933
rect 11962 -7967 11982 -7933
rect 13580 -7931 13658 -7897
rect 13692 -7931 13786 -7897
rect 13820 -7931 13914 -7897
rect 13948 -7931 14042 -7897
rect 14076 -7931 14096 -7897
rect 13580 -8001 14096 -7931
rect 14130 -7933 14649 -7863
rect 14684 -7716 14742 -7645
rect 14684 -7750 14696 -7716
rect 14730 -7750 14742 -7716
rect 14684 -7809 14742 -7750
rect 14684 -7843 14696 -7809
rect 14730 -7843 14742 -7809
rect 14684 -7878 14742 -7843
rect 14776 -7687 15845 -7645
rect 14776 -7721 14794 -7687
rect 14828 -7721 15794 -7687
rect 15828 -7721 15845 -7687
rect 14776 -7789 15845 -7721
rect 14776 -7823 14794 -7789
rect 14828 -7823 15794 -7789
rect 15828 -7823 15845 -7789
rect 14776 -7863 15845 -7823
rect 14130 -7967 14150 -7933
rect 14184 -7967 14278 -7933
rect 14312 -7967 14406 -7933
rect 14440 -7967 14534 -7933
rect 14568 -7967 14649 -7933
rect 14776 -7931 14854 -7897
rect 14888 -7931 14982 -7897
rect 15016 -7931 15110 -7897
rect 15144 -7931 15238 -7897
rect 15272 -7931 15292 -7897
rect 14776 -8001 15292 -7931
rect 15326 -7933 15845 -7863
rect 15880 -7716 15938 -7645
rect 15880 -7750 15892 -7716
rect 15926 -7750 15938 -7716
rect 15880 -7809 15938 -7750
rect 15880 -7843 15892 -7809
rect 15926 -7843 15938 -7809
rect 15880 -7878 15938 -7843
rect 15972 -7687 16674 -7645
rect 15972 -7721 15990 -7687
rect 16024 -7721 16622 -7687
rect 16656 -7721 16674 -7687
rect 15972 -7789 16674 -7721
rect 15972 -7823 15990 -7789
rect 16024 -7823 16622 -7789
rect 16656 -7823 16674 -7789
rect 15972 -7863 16674 -7823
rect 15326 -7967 15346 -7933
rect 15380 -7967 15474 -7933
rect 15508 -7967 15602 -7933
rect 15636 -7967 15730 -7933
rect 15764 -7967 15845 -7933
rect 15972 -7931 16050 -7897
rect 16084 -7931 16149 -7897
rect 16183 -7931 16248 -7897
rect 16282 -7931 16302 -7897
rect 15972 -8001 16302 -7931
rect 16336 -7933 16674 -7863
rect 16336 -7967 16356 -7933
rect 16390 -7967 16459 -7933
rect 16493 -7967 16562 -7933
rect 16596 -7967 16674 -7933
rect 11150 -8045 11166 -8011
rect 11200 -8045 11334 -8011
rect 11368 -8045 11384 -8011
rect 11452 -8045 11468 -8011
rect 10898 -8113 10914 -8079
rect 10948 -8113 10964 -8079
rect 10898 -8121 10964 -8113
rect 10998 -8079 11032 -8063
rect 10998 -8155 11032 -8113
rect 11066 -8079 11116 -8045
rect 11418 -8079 11468 -8045
rect 11066 -8113 11082 -8079
rect 11116 -8113 11250 -8079
rect 11284 -8113 11418 -8079
rect 11452 -8113 11468 -8079
rect 11066 -8121 11468 -8113
rect 11556 -8027 11614 -8010
rect 11556 -8061 11568 -8027
rect 11602 -8061 11614 -8027
rect 11556 -8155 11614 -8061
rect 11648 -8053 11982 -8001
rect 11648 -8087 11666 -8053
rect 11700 -8087 11930 -8053
rect 11964 -8087 11982 -8053
rect 11648 -8155 11982 -8087
rect 13488 -8027 13546 -8010
rect 13488 -8061 13500 -8027
rect 13534 -8061 13546 -8027
rect 13488 -8155 13546 -8061
rect 13580 -8060 14649 -8001
rect 13580 -8094 13598 -8060
rect 13632 -8094 14598 -8060
rect 14632 -8094 14649 -8060
rect 13580 -8155 14649 -8094
rect 14684 -8027 14742 -8010
rect 14684 -8061 14696 -8027
rect 14730 -8061 14742 -8027
rect 14684 -8155 14742 -8061
rect 14776 -8060 15845 -8001
rect 14776 -8094 14794 -8060
rect 14828 -8094 15794 -8060
rect 15828 -8094 15845 -8060
rect 14776 -8155 15845 -8094
rect 15880 -8027 15938 -8010
rect 15880 -8061 15892 -8027
rect 15926 -8061 15938 -8027
rect 15880 -8155 15938 -8061
rect 15972 -8060 16674 -8001
rect 15972 -8094 15990 -8060
rect 16024 -8094 16622 -8060
rect 16656 -8094 16674 -8060
rect 15972 -8155 16674 -8094
rect -2997 -8189 -2968 -8155
rect -2934 -8189 -2876 -8155
rect -2842 -8189 -2784 -8155
rect -2750 -8189 -2692 -8155
rect -2658 -8189 -2600 -8155
rect -2566 -8189 -2508 -8155
rect -2474 -8189 -2416 -8155
rect -2382 -8189 -2324 -8155
rect -2290 -8189 -2232 -8155
rect -2198 -8189 -2140 -8155
rect -2106 -8189 -2048 -8155
rect -2014 -8189 -1956 -8155
rect -1922 -8189 -1864 -8155
rect -1830 -8189 -1772 -8155
rect -1738 -8189 -1680 -8155
rect -1646 -8189 -1588 -8155
rect -1554 -8189 -1496 -8155
rect -1462 -8189 -1404 -8155
rect -1370 -8189 -1312 -8155
rect -1278 -8189 -1220 -8155
rect -1186 -8189 -1128 -8155
rect -1094 -8189 -1036 -8155
rect -1002 -8189 -944 -8155
rect -910 -8189 -852 -8155
rect -818 -8189 -760 -8155
rect -726 -8189 -668 -8155
rect -634 -8189 -576 -8155
rect -542 -8189 -484 -8155
rect -450 -8189 -392 -8155
rect -358 -8189 -300 -8155
rect -266 -8189 -208 -8155
rect -174 -8189 -116 -8155
rect -82 -8189 -24 -8155
rect 10 -8189 68 -8155
rect 102 -8189 160 -8155
rect 194 -8189 252 -8155
rect 286 -8189 344 -8155
rect 378 -8189 436 -8155
rect 470 -8189 528 -8155
rect 562 -8189 620 -8155
rect 654 -8189 712 -8155
rect 746 -8189 804 -8155
rect 838 -8189 896 -8155
rect 930 -8189 988 -8155
rect 1022 -8189 1080 -8155
rect 1114 -8189 1172 -8155
rect 1206 -8189 1264 -8155
rect 1298 -8189 1356 -8155
rect 1390 -8189 1448 -8155
rect 1482 -8189 1540 -8155
rect 1574 -8189 1632 -8155
rect 1666 -8189 1724 -8155
rect 1758 -8189 1816 -8155
rect 1850 -8189 1908 -8155
rect 1942 -8189 2000 -8155
rect 2034 -8189 2092 -8155
rect 2126 -8189 2184 -8155
rect 2218 -8189 2276 -8155
rect 2310 -8189 2368 -8155
rect 2402 -8189 2460 -8155
rect 2494 -8189 2552 -8155
rect 2586 -8189 2644 -8155
rect 2678 -8189 2736 -8155
rect 2770 -8189 2828 -8155
rect 2862 -8189 2920 -8155
rect 2954 -8189 3012 -8155
rect 3046 -8189 3104 -8155
rect 3138 -8189 3196 -8155
rect 3230 -8189 3288 -8155
rect 3322 -8189 3380 -8155
rect 3414 -8189 3472 -8155
rect 3506 -8189 3564 -8155
rect 3598 -8189 3656 -8155
rect 3690 -8189 3748 -8155
rect 3782 -8189 3840 -8155
rect 3874 -8189 3932 -8155
rect 3966 -8189 4024 -8155
rect 4058 -8189 4116 -8155
rect 4150 -8189 4208 -8155
rect 4242 -8189 4300 -8155
rect 4334 -8189 4392 -8155
rect 4426 -8189 4484 -8155
rect 4518 -8189 4576 -8155
rect 4610 -8189 4668 -8155
rect 4702 -8189 4760 -8155
rect 4794 -8189 4852 -8155
rect 4886 -8189 4944 -8155
rect 4978 -8189 5036 -8155
rect 5070 -8189 5128 -8155
rect 5162 -8189 5220 -8155
rect 5254 -8189 5312 -8155
rect 5346 -8189 5404 -8155
rect 5438 -8189 5496 -8155
rect 5530 -8189 5588 -8155
rect 5622 -8189 5680 -8155
rect 5714 -8189 5772 -8155
rect 5806 -8189 5864 -8155
rect 5898 -8189 5956 -8155
rect 5990 -8189 6048 -8155
rect 6082 -8189 6140 -8155
rect 6174 -8189 6232 -8155
rect 6266 -8189 6324 -8155
rect 6358 -8189 6416 -8155
rect 6450 -8189 6508 -8155
rect 6542 -8189 6600 -8155
rect 6634 -8189 6692 -8155
rect 6726 -8189 6784 -8155
rect 6818 -8189 6876 -8155
rect 6910 -8189 6968 -8155
rect 7002 -8189 7060 -8155
rect 7094 -8189 7152 -8155
rect 7186 -8189 7244 -8155
rect 7278 -8189 7336 -8155
rect 7370 -8189 7428 -8155
rect 7462 -8189 7520 -8155
rect 7554 -8189 7612 -8155
rect 7646 -8189 7704 -8155
rect 7738 -8189 7796 -8155
rect 7830 -8189 7888 -8155
rect 7922 -8189 7980 -8155
rect 8014 -8189 8072 -8155
rect 8106 -8189 8164 -8155
rect 8198 -8189 8256 -8155
rect 8290 -8189 8348 -8155
rect 8382 -8189 8440 -8155
rect 8474 -8189 8532 -8155
rect 8566 -8189 8624 -8155
rect 8658 -8189 8716 -8155
rect 8750 -8189 8808 -8155
rect 8842 -8189 8900 -8155
rect 8934 -8189 8992 -8155
rect 9026 -8189 9084 -8155
rect 9118 -8189 9176 -8155
rect 9210 -8189 9268 -8155
rect 9302 -8189 9360 -8155
rect 9394 -8189 9452 -8155
rect 9486 -8189 9544 -8155
rect 9578 -8189 9636 -8155
rect 9670 -8189 9728 -8155
rect 9762 -8189 9820 -8155
rect 9854 -8189 9912 -8155
rect 9946 -8189 10004 -8155
rect 10038 -8189 10096 -8155
rect 10130 -8189 10188 -8155
rect 10222 -8189 10280 -8155
rect 10314 -8189 10372 -8155
rect 10406 -8189 10464 -8155
rect 10498 -8189 10556 -8155
rect 10590 -8189 10648 -8155
rect 10682 -8189 10740 -8155
rect 10774 -8189 10832 -8155
rect 10866 -8189 10924 -8155
rect 10958 -8189 11016 -8155
rect 11050 -8189 11108 -8155
rect 11142 -8189 11200 -8155
rect 11234 -8189 11292 -8155
rect 11326 -8189 11384 -8155
rect 11418 -8189 11476 -8155
rect 11510 -8189 11568 -8155
rect 11602 -8189 11660 -8155
rect 11694 -8189 11752 -8155
rect 11786 -8189 11844 -8155
rect 11878 -8189 11936 -8155
rect 11970 -8189 12028 -8155
rect 12062 -8189 12120 -8155
rect 12154 -8189 12212 -8155
rect 12246 -8189 12304 -8155
rect 12338 -8189 12396 -8155
rect 12430 -8189 12488 -8155
rect 12522 -8189 12580 -8155
rect 12614 -8189 12672 -8155
rect 12706 -8189 12764 -8155
rect 12798 -8189 12856 -8155
rect 12890 -8189 12948 -8155
rect 12982 -8189 13040 -8155
rect 13074 -8189 13132 -8155
rect 13166 -8189 13224 -8155
rect 13258 -8189 13316 -8155
rect 13350 -8189 13408 -8155
rect 13442 -8189 13500 -8155
rect 13534 -8189 13592 -8155
rect 13626 -8189 13684 -8155
rect 13718 -8189 13776 -8155
rect 13810 -8189 13868 -8155
rect 13902 -8189 13960 -8155
rect 13994 -8189 14052 -8155
rect 14086 -8189 14144 -8155
rect 14178 -8189 14236 -8155
rect 14270 -8189 14328 -8155
rect 14362 -8189 14420 -8155
rect 14454 -8189 14512 -8155
rect 14546 -8189 14604 -8155
rect 14638 -8189 14696 -8155
rect 14730 -8189 14788 -8155
rect 14822 -8189 14880 -8155
rect 14914 -8189 14972 -8155
rect 15006 -8189 15064 -8155
rect 15098 -8189 15156 -8155
rect 15190 -8189 15248 -8155
rect 15282 -8189 15340 -8155
rect 15374 -8189 15432 -8155
rect 15466 -8189 15524 -8155
rect 15558 -8189 15616 -8155
rect 15650 -8189 15708 -8155
rect 15742 -8189 15800 -8155
rect 15834 -8189 15892 -8155
rect 15926 -8189 15984 -8155
rect 16018 -8189 16076 -8155
rect 16110 -8189 16168 -8155
rect 16202 -8189 16260 -8155
rect 16294 -8189 16352 -8155
rect 16386 -8189 16444 -8155
rect 16478 -8189 16536 -8155
rect 16570 -8189 16628 -8155
rect 16662 -8189 16691 -8155
rect -2980 -8250 -2278 -8189
rect -2980 -8284 -2962 -8250
rect -2928 -8284 -2330 -8250
rect -2296 -8284 -2278 -8250
rect -2980 -8343 -2278 -8284
rect -2244 -8283 -2186 -8189
rect -2244 -8317 -2232 -8283
rect -2198 -8317 -2186 -8283
rect -2244 -8334 -2186 -8317
rect -1600 -8250 -898 -8189
rect -1600 -8284 -1582 -8250
rect -1548 -8284 -950 -8250
rect -916 -8284 -898 -8250
rect -1600 -8343 -898 -8284
rect -864 -8250 -162 -8189
rect -864 -8284 -846 -8250
rect -812 -8284 -214 -8250
rect -180 -8284 -162 -8250
rect -864 -8343 -162 -8284
rect -128 -8283 -70 -8189
rect -128 -8317 -116 -8283
rect -82 -8317 -70 -8283
rect -128 -8334 -70 -8317
rect -36 -8257 298 -8189
rect -36 -8291 -18 -8257
rect 16 -8291 246 -8257
rect 280 -8291 298 -8257
rect -36 -8343 298 -8291
rect 332 -8283 390 -8189
rect 332 -8317 344 -8283
rect 378 -8317 390 -8283
rect 332 -8334 390 -8317
rect 424 -8242 505 -8223
rect 424 -8276 457 -8242
rect 491 -8276 505 -8242
rect 424 -8300 505 -8276
rect 539 -8242 605 -8189
rect 539 -8276 555 -8242
rect 589 -8276 605 -8242
rect 539 -8292 605 -8276
rect 695 -8242 745 -8223
rect 695 -8276 711 -8242
rect -2980 -8411 -2902 -8377
rect -2868 -8411 -2799 -8377
rect -2765 -8411 -2696 -8377
rect -2662 -8411 -2642 -8377
rect -2980 -8481 -2642 -8411
rect -2608 -8413 -2278 -8343
rect -2608 -8447 -2588 -8413
rect -2554 -8447 -2489 -8413
rect -2455 -8447 -2390 -8413
rect -2356 -8447 -2278 -8413
rect -1600 -8411 -1522 -8377
rect -1488 -8411 -1419 -8377
rect -1385 -8411 -1316 -8377
rect -1282 -8411 -1262 -8377
rect -2980 -8521 -2278 -8481
rect -2980 -8555 -2962 -8521
rect -2928 -8555 -2330 -8521
rect -2296 -8555 -2278 -8521
rect -2980 -8623 -2278 -8555
rect -2980 -8657 -2962 -8623
rect -2928 -8657 -2330 -8623
rect -2296 -8657 -2278 -8623
rect -2980 -8699 -2278 -8657
rect -2244 -8501 -2186 -8466
rect -2244 -8535 -2232 -8501
rect -2198 -8535 -2186 -8501
rect -2244 -8594 -2186 -8535
rect -2244 -8628 -2232 -8594
rect -2198 -8628 -2186 -8594
rect -2244 -8699 -2186 -8628
rect -1600 -8481 -1262 -8411
rect -1228 -8413 -898 -8343
rect -1228 -8447 -1208 -8413
rect -1174 -8447 -1109 -8413
rect -1075 -8447 -1010 -8413
rect -976 -8447 -898 -8413
rect -864 -8411 -786 -8377
rect -752 -8411 -683 -8377
rect -649 -8411 -580 -8377
rect -546 -8411 -526 -8377
rect -864 -8481 -526 -8411
rect -492 -8413 -162 -8343
rect -492 -8447 -472 -8413
rect -438 -8447 -373 -8413
rect -339 -8447 -274 -8413
rect -240 -8447 -162 -8413
rect -36 -8411 -16 -8377
rect 18 -8411 114 -8377
rect -1600 -8521 -898 -8481
rect -1600 -8555 -1582 -8521
rect -1548 -8555 -950 -8521
rect -916 -8555 -898 -8521
rect -1600 -8623 -898 -8555
rect -1600 -8657 -1582 -8623
rect -1548 -8657 -950 -8623
rect -916 -8657 -898 -8623
rect -1600 -8699 -898 -8657
rect -864 -8521 -162 -8481
rect -864 -8555 -846 -8521
rect -812 -8555 -214 -8521
rect -180 -8555 -162 -8521
rect -864 -8623 -162 -8555
rect -864 -8657 -846 -8623
rect -812 -8657 -214 -8623
rect -180 -8657 -162 -8623
rect -864 -8699 -162 -8657
rect -128 -8501 -70 -8466
rect -128 -8535 -116 -8501
rect -82 -8535 -70 -8501
rect -128 -8594 -70 -8535
rect -128 -8628 -116 -8594
rect -82 -8628 -70 -8594
rect -128 -8699 -70 -8628
rect -36 -8481 114 -8411
rect 148 -8413 298 -8343
rect 148 -8447 244 -8413
rect 278 -8447 298 -8413
rect 424 -8428 474 -8300
rect 695 -8318 745 -8276
rect 627 -8352 745 -8318
rect 797 -8242 867 -8223
rect 797 -8276 816 -8242
rect 850 -8276 867 -8242
rect 627 -8371 661 -8352
rect 424 -8462 433 -8428
rect 467 -8462 474 -8428
rect 508 -8387 661 -8371
rect 797 -8386 867 -8276
rect 960 -8242 1026 -8189
rect 960 -8276 976 -8242
rect 1010 -8276 1026 -8242
rect 960 -8285 1026 -8276
rect 1060 -8242 1126 -8223
rect 1060 -8276 1073 -8242
rect 1107 -8276 1126 -8242
rect 1060 -8319 1126 -8276
rect 932 -8353 1126 -8319
rect 1160 -8283 1218 -8189
rect 1160 -8317 1172 -8283
rect 1206 -8317 1218 -8283
rect 1160 -8334 1218 -8317
rect 1252 -8257 1586 -8189
rect 1252 -8291 1270 -8257
rect 1304 -8291 1534 -8257
rect 1568 -8291 1586 -8257
rect 1252 -8343 1586 -8291
rect 1620 -8283 1678 -8189
rect 1620 -8317 1632 -8283
rect 1666 -8317 1678 -8283
rect 1620 -8334 1678 -8317
rect 1712 -8250 2414 -8189
rect 1712 -8284 1730 -8250
rect 1764 -8284 2362 -8250
rect 2396 -8284 2414 -8250
rect 1712 -8343 2414 -8284
rect 2448 -8283 2506 -8189
rect 2448 -8317 2460 -8283
rect 2494 -8317 2506 -8283
rect 2448 -8334 2506 -8317
rect 2540 -8257 2874 -8189
rect 2540 -8291 2558 -8257
rect 2592 -8291 2822 -8257
rect 2856 -8291 2874 -8257
rect 2540 -8343 2874 -8291
rect 2908 -8283 2966 -8189
rect 2908 -8317 2920 -8283
rect 2954 -8317 2966 -8283
rect 2908 -8334 2966 -8317
rect 3000 -8242 3081 -8223
rect 3000 -8276 3033 -8242
rect 3067 -8276 3081 -8242
rect 3000 -8300 3081 -8276
rect 3115 -8242 3181 -8189
rect 3115 -8276 3131 -8242
rect 3165 -8276 3181 -8242
rect 3115 -8292 3181 -8276
rect 3271 -8242 3321 -8223
rect 3271 -8276 3287 -8242
rect 932 -8377 1002 -8353
rect 508 -8421 511 -8387
rect 545 -8421 661 -8387
rect 508 -8437 661 -8421
rect 695 -8387 867 -8386
rect 695 -8421 711 -8387
rect 745 -8421 867 -8387
rect 695 -8436 867 -8421
rect 916 -8387 1002 -8377
rect 916 -8421 932 -8387
rect 966 -8421 1002 -8387
rect 916 -8435 1002 -8421
rect 1036 -8425 1052 -8387
rect 1086 -8425 1126 -8387
rect 1036 -8430 1126 -8425
rect 1252 -8411 1272 -8377
rect 1306 -8411 1402 -8377
rect -36 -8521 298 -8481
rect -36 -8555 -18 -8521
rect 16 -8555 246 -8521
rect 280 -8555 298 -8521
rect -36 -8623 298 -8555
rect -36 -8657 -18 -8623
rect 16 -8657 246 -8623
rect 280 -8657 298 -8623
rect -36 -8699 298 -8657
rect 332 -8501 390 -8466
rect 332 -8535 344 -8501
rect 378 -8535 390 -8501
rect 332 -8594 390 -8535
rect 332 -8628 344 -8594
rect 378 -8628 390 -8594
rect 332 -8699 390 -8628
rect 424 -8510 474 -8462
rect 627 -8471 661 -8437
rect 627 -8505 745 -8471
rect 424 -8547 505 -8510
rect 424 -8581 457 -8547
rect 491 -8581 505 -8547
rect 424 -8615 505 -8581
rect 424 -8649 457 -8615
rect 491 -8649 505 -8615
rect 424 -8665 505 -8649
rect 539 -8548 605 -8539
rect 539 -8582 555 -8548
rect 589 -8582 605 -8548
rect 539 -8616 605 -8582
rect 539 -8650 555 -8616
rect 589 -8650 605 -8616
rect 539 -8699 605 -8650
rect 695 -8547 745 -8505
rect 695 -8581 711 -8547
rect 695 -8615 745 -8581
rect 695 -8649 711 -8615
rect 695 -8665 745 -8649
rect 797 -8548 867 -8436
rect 932 -8464 1002 -8435
rect 932 -8498 1126 -8464
rect 797 -8582 815 -8548
rect 849 -8582 867 -8548
rect 797 -8616 867 -8582
rect 797 -8650 815 -8616
rect 849 -8650 867 -8616
rect 797 -8665 867 -8650
rect 957 -8548 1023 -8532
rect 957 -8582 973 -8548
rect 1007 -8582 1023 -8548
rect 957 -8616 1023 -8582
rect 957 -8650 973 -8616
rect 1007 -8650 1023 -8616
rect 957 -8699 1023 -8650
rect 1057 -8548 1126 -8498
rect 1057 -8582 1073 -8548
rect 1107 -8582 1126 -8548
rect 1057 -8616 1126 -8582
rect 1057 -8650 1073 -8616
rect 1107 -8650 1126 -8616
rect 1057 -8665 1126 -8650
rect 1160 -8501 1218 -8466
rect 1160 -8535 1172 -8501
rect 1206 -8535 1218 -8501
rect 1160 -8594 1218 -8535
rect 1160 -8628 1172 -8594
rect 1206 -8628 1218 -8594
rect 1160 -8699 1218 -8628
rect 1252 -8481 1402 -8411
rect 1436 -8413 1586 -8343
rect 1436 -8447 1532 -8413
rect 1566 -8447 1586 -8413
rect 1712 -8411 1790 -8377
rect 1824 -8411 1893 -8377
rect 1927 -8411 1996 -8377
rect 2030 -8411 2050 -8377
rect 1252 -8521 1586 -8481
rect 1252 -8555 1270 -8521
rect 1304 -8555 1534 -8521
rect 1568 -8555 1586 -8521
rect 1252 -8623 1586 -8555
rect 1252 -8657 1270 -8623
rect 1304 -8657 1534 -8623
rect 1568 -8657 1586 -8623
rect 1252 -8699 1586 -8657
rect 1620 -8501 1678 -8466
rect 1620 -8535 1632 -8501
rect 1666 -8535 1678 -8501
rect 1620 -8594 1678 -8535
rect 1620 -8628 1632 -8594
rect 1666 -8628 1678 -8594
rect 1620 -8699 1678 -8628
rect 1712 -8481 2050 -8411
rect 2084 -8413 2414 -8343
rect 2084 -8447 2104 -8413
rect 2138 -8447 2203 -8413
rect 2237 -8447 2302 -8413
rect 2336 -8447 2414 -8413
rect 2540 -8411 2560 -8377
rect 2594 -8411 2690 -8377
rect 1712 -8521 2414 -8481
rect 1712 -8555 1730 -8521
rect 1764 -8555 2362 -8521
rect 2396 -8555 2414 -8521
rect 1712 -8623 2414 -8555
rect 1712 -8657 1730 -8623
rect 1764 -8657 2362 -8623
rect 2396 -8657 2414 -8623
rect 1712 -8699 2414 -8657
rect 2448 -8501 2506 -8466
rect 2448 -8535 2460 -8501
rect 2494 -8535 2506 -8501
rect 2448 -8594 2506 -8535
rect 2448 -8628 2460 -8594
rect 2494 -8628 2506 -8594
rect 2448 -8699 2506 -8628
rect 2540 -8481 2690 -8411
rect 2724 -8413 2874 -8343
rect 2724 -8447 2820 -8413
rect 2854 -8447 2874 -8413
rect 3000 -8391 3050 -8300
rect 3271 -8318 3321 -8276
rect 3203 -8352 3321 -8318
rect 3373 -8242 3443 -8223
rect 3373 -8276 3392 -8242
rect 3426 -8276 3443 -8242
rect 3203 -8371 3237 -8352
rect 3000 -8425 3012 -8391
rect 3046 -8425 3050 -8391
rect 2540 -8521 2874 -8481
rect 2540 -8555 2558 -8521
rect 2592 -8555 2822 -8521
rect 2856 -8555 2874 -8521
rect 2540 -8623 2874 -8555
rect 2540 -8657 2558 -8623
rect 2592 -8657 2822 -8623
rect 2856 -8657 2874 -8623
rect 2540 -8699 2874 -8657
rect 2908 -8501 2966 -8466
rect 2908 -8535 2920 -8501
rect 2954 -8535 2966 -8501
rect 2908 -8594 2966 -8535
rect 2908 -8628 2920 -8594
rect 2954 -8628 2966 -8594
rect 2908 -8699 2966 -8628
rect 3000 -8510 3050 -8425
rect 3084 -8387 3237 -8371
rect 3373 -8386 3443 -8276
rect 3536 -8242 3602 -8189
rect 3536 -8276 3552 -8242
rect 3586 -8276 3602 -8242
rect 3536 -8285 3602 -8276
rect 3636 -8242 3702 -8223
rect 3636 -8276 3649 -8242
rect 3683 -8276 3702 -8242
rect 3636 -8319 3702 -8276
rect 3508 -8353 3702 -8319
rect 3736 -8283 3794 -8189
rect 3736 -8317 3748 -8283
rect 3782 -8317 3794 -8283
rect 3736 -8334 3794 -8317
rect 3828 -8257 4162 -8189
rect 3828 -8291 3846 -8257
rect 3880 -8291 4110 -8257
rect 4144 -8291 4162 -8257
rect 3828 -8343 4162 -8291
rect 4196 -8283 4254 -8189
rect 4196 -8317 4208 -8283
rect 4242 -8317 4254 -8283
rect 4196 -8334 4254 -8317
rect 4288 -8250 4990 -8189
rect 4288 -8284 4306 -8250
rect 4340 -8284 4938 -8250
rect 4972 -8284 4990 -8250
rect 4288 -8343 4990 -8284
rect 5024 -8283 5082 -8189
rect 5024 -8317 5036 -8283
rect 5070 -8317 5082 -8283
rect 5024 -8334 5082 -8317
rect 5116 -8257 5450 -8189
rect 5116 -8291 5134 -8257
rect 5168 -8291 5398 -8257
rect 5432 -8291 5450 -8257
rect 5116 -8343 5450 -8291
rect 5484 -8283 5542 -8189
rect 5484 -8317 5496 -8283
rect 5530 -8317 5542 -8283
rect 5484 -8334 5542 -8317
rect 5576 -8242 5657 -8223
rect 5576 -8276 5609 -8242
rect 5643 -8276 5657 -8242
rect 5576 -8300 5657 -8276
rect 5691 -8242 5757 -8189
rect 5691 -8276 5707 -8242
rect 5741 -8276 5757 -8242
rect 5691 -8292 5757 -8276
rect 5847 -8242 5897 -8223
rect 5847 -8276 5863 -8242
rect 3508 -8377 3578 -8353
rect 3084 -8421 3087 -8387
rect 3121 -8421 3237 -8387
rect 3084 -8437 3237 -8421
rect 3271 -8387 3443 -8386
rect 3271 -8421 3287 -8387
rect 3321 -8421 3443 -8387
rect 3271 -8436 3443 -8421
rect 3492 -8387 3578 -8377
rect 3492 -8421 3508 -8387
rect 3542 -8421 3578 -8387
rect 3492 -8435 3578 -8421
rect 3612 -8391 3628 -8387
rect 3612 -8425 3626 -8391
rect 3662 -8421 3702 -8387
rect 3660 -8425 3702 -8421
rect 3612 -8430 3702 -8425
rect 3828 -8411 3848 -8377
rect 3882 -8411 3978 -8377
rect 3203 -8471 3237 -8437
rect 3203 -8505 3321 -8471
rect 3000 -8547 3081 -8510
rect 3000 -8581 3033 -8547
rect 3067 -8581 3081 -8547
rect 3000 -8615 3081 -8581
rect 3000 -8649 3033 -8615
rect 3067 -8649 3081 -8615
rect 3000 -8665 3081 -8649
rect 3115 -8548 3181 -8539
rect 3115 -8582 3131 -8548
rect 3165 -8582 3181 -8548
rect 3115 -8616 3181 -8582
rect 3115 -8650 3131 -8616
rect 3165 -8650 3181 -8616
rect 3115 -8699 3181 -8650
rect 3271 -8547 3321 -8505
rect 3271 -8581 3287 -8547
rect 3271 -8615 3321 -8581
rect 3271 -8649 3287 -8615
rect 3271 -8665 3321 -8649
rect 3373 -8548 3443 -8436
rect 3508 -8464 3578 -8435
rect 3508 -8498 3702 -8464
rect 3373 -8582 3391 -8548
rect 3425 -8582 3443 -8548
rect 3373 -8616 3443 -8582
rect 3373 -8650 3391 -8616
rect 3425 -8650 3443 -8616
rect 3373 -8665 3443 -8650
rect 3533 -8548 3599 -8532
rect 3533 -8582 3549 -8548
rect 3583 -8582 3599 -8548
rect 3533 -8616 3599 -8582
rect 3533 -8650 3549 -8616
rect 3583 -8650 3599 -8616
rect 3533 -8699 3599 -8650
rect 3633 -8548 3702 -8498
rect 3633 -8582 3649 -8548
rect 3683 -8582 3702 -8548
rect 3633 -8616 3702 -8582
rect 3633 -8650 3649 -8616
rect 3683 -8650 3702 -8616
rect 3633 -8665 3702 -8650
rect 3736 -8501 3794 -8466
rect 3736 -8535 3748 -8501
rect 3782 -8535 3794 -8501
rect 3736 -8594 3794 -8535
rect 3736 -8628 3748 -8594
rect 3782 -8628 3794 -8594
rect 3736 -8699 3794 -8628
rect 3828 -8481 3978 -8411
rect 4012 -8413 4162 -8343
rect 4012 -8447 4108 -8413
rect 4142 -8447 4162 -8413
rect 4288 -8411 4366 -8377
rect 4400 -8411 4469 -8377
rect 4503 -8411 4572 -8377
rect 4606 -8411 4626 -8377
rect 3828 -8521 4162 -8481
rect 3828 -8555 3846 -8521
rect 3880 -8555 4110 -8521
rect 4144 -8555 4162 -8521
rect 3828 -8623 4162 -8555
rect 3828 -8657 3846 -8623
rect 3880 -8657 4110 -8623
rect 4144 -8657 4162 -8623
rect 3828 -8699 4162 -8657
rect 4196 -8501 4254 -8466
rect 4196 -8535 4208 -8501
rect 4242 -8535 4254 -8501
rect 4196 -8594 4254 -8535
rect 4196 -8628 4208 -8594
rect 4242 -8628 4254 -8594
rect 4196 -8699 4254 -8628
rect 4288 -8481 4626 -8411
rect 4660 -8413 4990 -8343
rect 4660 -8447 4680 -8413
rect 4714 -8447 4779 -8413
rect 4813 -8447 4878 -8413
rect 4912 -8447 4990 -8413
rect 5116 -8411 5136 -8377
rect 5170 -8411 5266 -8377
rect 4288 -8521 4990 -8481
rect 4288 -8555 4306 -8521
rect 4340 -8555 4938 -8521
rect 4972 -8555 4990 -8521
rect 4288 -8623 4990 -8555
rect 4288 -8657 4306 -8623
rect 4340 -8657 4938 -8623
rect 4972 -8657 4990 -8623
rect 4288 -8699 4990 -8657
rect 5024 -8501 5082 -8466
rect 5024 -8535 5036 -8501
rect 5070 -8535 5082 -8501
rect 5024 -8594 5082 -8535
rect 5024 -8628 5036 -8594
rect 5070 -8628 5082 -8594
rect 5024 -8699 5082 -8628
rect 5116 -8481 5266 -8411
rect 5300 -8413 5450 -8343
rect 5300 -8447 5396 -8413
rect 5430 -8447 5450 -8413
rect 5576 -8391 5626 -8300
rect 5847 -8318 5897 -8276
rect 5779 -8352 5897 -8318
rect 5949 -8242 6019 -8223
rect 5949 -8276 5968 -8242
rect 6002 -8276 6019 -8242
rect 5779 -8371 5813 -8352
rect 5576 -8425 5586 -8391
rect 5620 -8425 5626 -8391
rect 5116 -8521 5450 -8481
rect 5116 -8555 5134 -8521
rect 5168 -8555 5398 -8521
rect 5432 -8555 5450 -8521
rect 5116 -8623 5450 -8555
rect 5116 -8657 5134 -8623
rect 5168 -8657 5398 -8623
rect 5432 -8657 5450 -8623
rect 5116 -8699 5450 -8657
rect 5484 -8501 5542 -8466
rect 5484 -8535 5496 -8501
rect 5530 -8535 5542 -8501
rect 5484 -8594 5542 -8535
rect 5484 -8628 5496 -8594
rect 5530 -8628 5542 -8594
rect 5484 -8699 5542 -8628
rect 5576 -8510 5626 -8425
rect 5660 -8387 5813 -8371
rect 5949 -8386 6019 -8276
rect 6112 -8242 6178 -8189
rect 6112 -8276 6128 -8242
rect 6162 -8276 6178 -8242
rect 6112 -8285 6178 -8276
rect 6212 -8242 6278 -8223
rect 6212 -8276 6225 -8242
rect 6259 -8276 6278 -8242
rect 6212 -8319 6278 -8276
rect 6084 -8353 6278 -8319
rect 6312 -8283 6370 -8189
rect 6312 -8317 6324 -8283
rect 6358 -8317 6370 -8283
rect 6312 -8334 6370 -8317
rect 6404 -8257 6738 -8189
rect 6404 -8291 6422 -8257
rect 6456 -8291 6686 -8257
rect 6720 -8291 6738 -8257
rect 6404 -8343 6738 -8291
rect 6772 -8283 6830 -8189
rect 6772 -8317 6784 -8283
rect 6818 -8317 6830 -8283
rect 6772 -8334 6830 -8317
rect 6864 -8250 7566 -8189
rect 6864 -8284 6882 -8250
rect 6916 -8284 7514 -8250
rect 7548 -8284 7566 -8250
rect 6864 -8343 7566 -8284
rect 7600 -8283 7658 -8189
rect 7600 -8317 7612 -8283
rect 7646 -8317 7658 -8283
rect 7600 -8334 7658 -8317
rect 7692 -8257 8026 -8189
rect 7692 -8291 7710 -8257
rect 7744 -8291 7974 -8257
rect 8008 -8291 8026 -8257
rect 7692 -8343 8026 -8291
rect 8060 -8283 8118 -8189
rect 8060 -8317 8072 -8283
rect 8106 -8317 8118 -8283
rect 8060 -8334 8118 -8317
rect 8152 -8242 8233 -8223
rect 8152 -8276 8185 -8242
rect 8219 -8276 8233 -8242
rect 8152 -8300 8233 -8276
rect 8267 -8242 8333 -8189
rect 8267 -8276 8283 -8242
rect 8317 -8276 8333 -8242
rect 8267 -8292 8333 -8276
rect 8423 -8242 8473 -8223
rect 8423 -8276 8439 -8242
rect 6084 -8377 6154 -8353
rect 5660 -8421 5663 -8387
rect 5697 -8421 5813 -8387
rect 5660 -8437 5813 -8421
rect 5847 -8387 6019 -8386
rect 5847 -8421 5863 -8387
rect 5897 -8421 6019 -8387
rect 5847 -8436 6019 -8421
rect 6068 -8387 6154 -8377
rect 6068 -8421 6084 -8387
rect 6118 -8421 6154 -8387
rect 6068 -8435 6154 -8421
rect 6188 -8391 6204 -8387
rect 6188 -8425 6200 -8391
rect 6238 -8421 6278 -8387
rect 6234 -8425 6278 -8421
rect 6188 -8430 6278 -8425
rect 6404 -8411 6424 -8377
rect 6458 -8411 6554 -8377
rect 5779 -8471 5813 -8437
rect 5779 -8505 5897 -8471
rect 5576 -8547 5657 -8510
rect 5576 -8581 5609 -8547
rect 5643 -8581 5657 -8547
rect 5576 -8615 5657 -8581
rect 5576 -8649 5609 -8615
rect 5643 -8649 5657 -8615
rect 5576 -8665 5657 -8649
rect 5691 -8548 5757 -8539
rect 5691 -8582 5707 -8548
rect 5741 -8582 5757 -8548
rect 5691 -8616 5757 -8582
rect 5691 -8650 5707 -8616
rect 5741 -8650 5757 -8616
rect 5691 -8699 5757 -8650
rect 5847 -8547 5897 -8505
rect 5847 -8581 5863 -8547
rect 5847 -8615 5897 -8581
rect 5847 -8649 5863 -8615
rect 5847 -8665 5897 -8649
rect 5949 -8548 6019 -8436
rect 6084 -8464 6154 -8435
rect 6084 -8498 6278 -8464
rect 5949 -8582 5967 -8548
rect 6001 -8582 6019 -8548
rect 5949 -8616 6019 -8582
rect 5949 -8650 5967 -8616
rect 6001 -8650 6019 -8616
rect 5949 -8665 6019 -8650
rect 6109 -8548 6175 -8532
rect 6109 -8582 6125 -8548
rect 6159 -8582 6175 -8548
rect 6109 -8616 6175 -8582
rect 6109 -8650 6125 -8616
rect 6159 -8650 6175 -8616
rect 6109 -8699 6175 -8650
rect 6209 -8548 6278 -8498
rect 6209 -8582 6225 -8548
rect 6259 -8582 6278 -8548
rect 6209 -8616 6278 -8582
rect 6209 -8650 6225 -8616
rect 6259 -8650 6278 -8616
rect 6209 -8665 6278 -8650
rect 6312 -8501 6370 -8466
rect 6312 -8535 6324 -8501
rect 6358 -8535 6370 -8501
rect 6312 -8594 6370 -8535
rect 6312 -8628 6324 -8594
rect 6358 -8628 6370 -8594
rect 6312 -8699 6370 -8628
rect 6404 -8481 6554 -8411
rect 6588 -8413 6738 -8343
rect 6588 -8447 6684 -8413
rect 6718 -8447 6738 -8413
rect 6864 -8411 6942 -8377
rect 6976 -8411 7045 -8377
rect 7079 -8411 7148 -8377
rect 7182 -8411 7202 -8377
rect 6404 -8521 6738 -8481
rect 6404 -8555 6422 -8521
rect 6456 -8555 6686 -8521
rect 6720 -8555 6738 -8521
rect 6404 -8623 6738 -8555
rect 6404 -8657 6422 -8623
rect 6456 -8657 6686 -8623
rect 6720 -8657 6738 -8623
rect 6404 -8699 6738 -8657
rect 6772 -8501 6830 -8466
rect 6772 -8535 6784 -8501
rect 6818 -8535 6830 -8501
rect 6772 -8594 6830 -8535
rect 6772 -8628 6784 -8594
rect 6818 -8628 6830 -8594
rect 6772 -8699 6830 -8628
rect 6864 -8481 7202 -8411
rect 7236 -8413 7566 -8343
rect 7236 -8447 7256 -8413
rect 7290 -8447 7355 -8413
rect 7389 -8447 7454 -8413
rect 7488 -8447 7566 -8413
rect 7692 -8411 7712 -8377
rect 7746 -8411 7842 -8377
rect 6864 -8521 7566 -8481
rect 6864 -8555 6882 -8521
rect 6916 -8555 7514 -8521
rect 7548 -8555 7566 -8521
rect 6864 -8623 7566 -8555
rect 6864 -8657 6882 -8623
rect 6916 -8657 7514 -8623
rect 7548 -8657 7566 -8623
rect 6864 -8699 7566 -8657
rect 7600 -8501 7658 -8466
rect 7600 -8535 7612 -8501
rect 7646 -8535 7658 -8501
rect 7600 -8594 7658 -8535
rect 7600 -8628 7612 -8594
rect 7646 -8628 7658 -8594
rect 7600 -8699 7658 -8628
rect 7692 -8481 7842 -8411
rect 7876 -8413 8026 -8343
rect 7876 -8447 7972 -8413
rect 8006 -8447 8026 -8413
rect 8152 -8391 8202 -8300
rect 8423 -8318 8473 -8276
rect 8355 -8352 8473 -8318
rect 8525 -8242 8595 -8223
rect 8525 -8276 8544 -8242
rect 8578 -8276 8595 -8242
rect 8355 -8371 8389 -8352
rect 8152 -8425 8160 -8391
rect 8194 -8425 8202 -8391
rect 7692 -8521 8026 -8481
rect 7692 -8555 7710 -8521
rect 7744 -8555 7974 -8521
rect 8008 -8555 8026 -8521
rect 7692 -8623 8026 -8555
rect 7692 -8657 7710 -8623
rect 7744 -8657 7974 -8623
rect 8008 -8657 8026 -8623
rect 7692 -8699 8026 -8657
rect 8060 -8501 8118 -8466
rect 8060 -8535 8072 -8501
rect 8106 -8535 8118 -8501
rect 8060 -8594 8118 -8535
rect 8060 -8628 8072 -8594
rect 8106 -8628 8118 -8594
rect 8060 -8699 8118 -8628
rect 8152 -8510 8202 -8425
rect 8236 -8387 8389 -8371
rect 8525 -8386 8595 -8276
rect 8688 -8242 8754 -8189
rect 8688 -8276 8704 -8242
rect 8738 -8276 8754 -8242
rect 8688 -8285 8754 -8276
rect 8788 -8242 8854 -8223
rect 8788 -8276 8801 -8242
rect 8835 -8276 8854 -8242
rect 8788 -8319 8854 -8276
rect 8660 -8353 8854 -8319
rect 8888 -8283 8946 -8189
rect 8888 -8317 8900 -8283
rect 8934 -8317 8946 -8283
rect 8888 -8334 8946 -8317
rect 8980 -8257 9314 -8189
rect 8980 -8291 8998 -8257
rect 9032 -8291 9262 -8257
rect 9296 -8291 9314 -8257
rect 8980 -8343 9314 -8291
rect 9348 -8283 9406 -8189
rect 9348 -8317 9360 -8283
rect 9394 -8317 9406 -8283
rect 9348 -8334 9406 -8317
rect 9440 -8250 10142 -8189
rect 9440 -8284 9458 -8250
rect 9492 -8284 10090 -8250
rect 10124 -8284 10142 -8250
rect 9440 -8343 10142 -8284
rect 10176 -8283 10234 -8189
rect 10176 -8317 10188 -8283
rect 10222 -8317 10234 -8283
rect 10176 -8334 10234 -8317
rect 10360 -8257 10694 -8189
rect 10360 -8291 10378 -8257
rect 10412 -8291 10642 -8257
rect 10676 -8291 10694 -8257
rect 10360 -8343 10694 -8291
rect 8660 -8377 8730 -8353
rect 8236 -8421 8239 -8387
rect 8273 -8421 8389 -8387
rect 8236 -8437 8389 -8421
rect 8423 -8387 8595 -8386
rect 8423 -8421 8439 -8387
rect 8473 -8421 8595 -8387
rect 8423 -8436 8595 -8421
rect 8644 -8387 8730 -8377
rect 8644 -8421 8660 -8387
rect 8694 -8421 8730 -8387
rect 8644 -8435 8730 -8421
rect 8764 -8391 8780 -8387
rect 8764 -8425 8774 -8391
rect 8814 -8421 8854 -8387
rect 8808 -8425 8854 -8421
rect 8764 -8430 8854 -8425
rect 8980 -8411 9000 -8377
rect 9034 -8411 9130 -8377
rect 8355 -8471 8389 -8437
rect 8355 -8505 8473 -8471
rect 8152 -8547 8233 -8510
rect 8152 -8581 8185 -8547
rect 8219 -8581 8233 -8547
rect 8152 -8615 8233 -8581
rect 8152 -8649 8185 -8615
rect 8219 -8649 8233 -8615
rect 8152 -8665 8233 -8649
rect 8267 -8548 8333 -8539
rect 8267 -8582 8283 -8548
rect 8317 -8582 8333 -8548
rect 8267 -8616 8333 -8582
rect 8267 -8650 8283 -8616
rect 8317 -8650 8333 -8616
rect 8267 -8699 8333 -8650
rect 8423 -8547 8473 -8505
rect 8423 -8581 8439 -8547
rect 8423 -8615 8473 -8581
rect 8423 -8649 8439 -8615
rect 8423 -8665 8473 -8649
rect 8525 -8548 8595 -8436
rect 8660 -8464 8730 -8435
rect 8660 -8498 8854 -8464
rect 8525 -8582 8543 -8548
rect 8577 -8582 8595 -8548
rect 8525 -8616 8595 -8582
rect 8525 -8650 8543 -8616
rect 8577 -8650 8595 -8616
rect 8525 -8665 8595 -8650
rect 8685 -8548 8751 -8532
rect 8685 -8582 8701 -8548
rect 8735 -8582 8751 -8548
rect 8685 -8616 8751 -8582
rect 8685 -8650 8701 -8616
rect 8735 -8650 8751 -8616
rect 8685 -8699 8751 -8650
rect 8785 -8548 8854 -8498
rect 8785 -8582 8801 -8548
rect 8835 -8582 8854 -8548
rect 8785 -8616 8854 -8582
rect 8785 -8650 8801 -8616
rect 8835 -8650 8854 -8616
rect 8785 -8665 8854 -8650
rect 8888 -8501 8946 -8466
rect 8888 -8535 8900 -8501
rect 8934 -8535 8946 -8501
rect 8888 -8594 8946 -8535
rect 8888 -8628 8900 -8594
rect 8934 -8628 8946 -8594
rect 8888 -8699 8946 -8628
rect 8980 -8481 9130 -8411
rect 9164 -8413 9314 -8343
rect 9164 -8447 9260 -8413
rect 9294 -8447 9314 -8413
rect 9440 -8411 9518 -8377
rect 9552 -8411 9621 -8377
rect 9655 -8411 9724 -8377
rect 9758 -8411 9778 -8377
rect 8980 -8521 9314 -8481
rect 8980 -8555 8998 -8521
rect 9032 -8555 9262 -8521
rect 9296 -8555 9314 -8521
rect 8980 -8623 9314 -8555
rect 8980 -8657 8998 -8623
rect 9032 -8657 9262 -8623
rect 9296 -8657 9314 -8623
rect 8980 -8699 9314 -8657
rect 9348 -8501 9406 -8466
rect 9348 -8535 9360 -8501
rect 9394 -8535 9406 -8501
rect 9348 -8594 9406 -8535
rect 9348 -8628 9360 -8594
rect 9394 -8628 9406 -8594
rect 9348 -8699 9406 -8628
rect 9440 -8481 9778 -8411
rect 9812 -8413 10142 -8343
rect 9812 -8447 9832 -8413
rect 9866 -8447 9931 -8413
rect 9965 -8447 10030 -8413
rect 10064 -8447 10142 -8413
rect 10360 -8411 10380 -8377
rect 10414 -8411 10510 -8377
rect 9440 -8521 10142 -8481
rect 9440 -8555 9458 -8521
rect 9492 -8555 10090 -8521
rect 10124 -8555 10142 -8521
rect 9440 -8623 10142 -8555
rect 9440 -8657 9458 -8623
rect 9492 -8657 10090 -8623
rect 10124 -8657 10142 -8623
rect 9440 -8699 10142 -8657
rect 10176 -8501 10234 -8466
rect 10176 -8535 10188 -8501
rect 10222 -8535 10234 -8501
rect 10176 -8594 10234 -8535
rect 10176 -8628 10188 -8594
rect 10222 -8628 10234 -8594
rect 10176 -8699 10234 -8628
rect 10360 -8481 10510 -8411
rect 10544 -8413 10694 -8343
rect 10544 -8447 10640 -8413
rect 10674 -8447 10694 -8413
rect 10728 -8242 10809 -8223
rect 10728 -8276 10761 -8242
rect 10795 -8276 10809 -8242
rect 10728 -8300 10809 -8276
rect 10843 -8242 10909 -8189
rect 10843 -8276 10859 -8242
rect 10893 -8276 10909 -8242
rect 10843 -8292 10909 -8276
rect 10999 -8242 11049 -8223
rect 10999 -8276 11015 -8242
rect 10728 -8393 10778 -8300
rect 10999 -8318 11049 -8276
rect 10931 -8352 11049 -8318
rect 11101 -8242 11171 -8223
rect 11101 -8276 11120 -8242
rect 11154 -8276 11171 -8242
rect 10931 -8371 10965 -8352
rect 10728 -8427 10737 -8393
rect 10771 -8427 10778 -8393
rect 10360 -8521 10694 -8481
rect 10360 -8555 10378 -8521
rect 10412 -8555 10642 -8521
rect 10676 -8555 10694 -8521
rect 10360 -8623 10694 -8555
rect 10360 -8657 10378 -8623
rect 10412 -8657 10642 -8623
rect 10676 -8657 10694 -8623
rect 10360 -8699 10694 -8657
rect 10728 -8510 10778 -8427
rect 10812 -8387 10965 -8371
rect 11101 -8386 11171 -8276
rect 11264 -8242 11330 -8189
rect 11264 -8276 11280 -8242
rect 11314 -8276 11330 -8242
rect 11264 -8285 11330 -8276
rect 11364 -8242 11430 -8223
rect 11364 -8276 11377 -8242
rect 11411 -8276 11430 -8242
rect 11364 -8319 11430 -8276
rect 11236 -8353 11430 -8319
rect 11464 -8283 11522 -8189
rect 11464 -8317 11476 -8283
rect 11510 -8317 11522 -8283
rect 11464 -8334 11522 -8317
rect 11648 -8257 11982 -8189
rect 11648 -8291 11666 -8257
rect 11700 -8291 11930 -8257
rect 11964 -8291 11982 -8257
rect 11648 -8343 11982 -8291
rect 13580 -8283 13638 -8189
rect 13580 -8317 13592 -8283
rect 13626 -8317 13638 -8283
rect 13672 -8231 13733 -8189
rect 13672 -8265 13690 -8231
rect 13724 -8265 13733 -8231
rect 13672 -8291 13733 -8265
rect 13769 -8244 13819 -8225
rect 13769 -8278 13776 -8244
rect 13810 -8278 13819 -8244
rect 13580 -8334 13638 -8317
rect 11236 -8377 11306 -8353
rect 10812 -8421 10815 -8387
rect 10849 -8421 10965 -8387
rect 10812 -8437 10965 -8421
rect 10999 -8387 11171 -8386
rect 10999 -8421 11015 -8387
rect 11049 -8421 11171 -8387
rect 10999 -8436 11171 -8421
rect 11220 -8387 11306 -8377
rect 11220 -8421 11236 -8387
rect 11270 -8421 11306 -8387
rect 11220 -8435 11306 -8421
rect 11340 -8421 11356 -8387
rect 11390 -8394 11430 -8387
rect 11340 -8428 11369 -8421
rect 11403 -8428 11430 -8394
rect 11340 -8430 11430 -8428
rect 11648 -8411 11668 -8377
rect 11702 -8411 11798 -8377
rect 10931 -8471 10965 -8437
rect 10931 -8505 11049 -8471
rect 10728 -8547 10809 -8510
rect 10728 -8581 10761 -8547
rect 10795 -8581 10809 -8547
rect 10728 -8615 10809 -8581
rect 10728 -8649 10761 -8615
rect 10795 -8649 10809 -8615
rect 10728 -8665 10809 -8649
rect 10843 -8548 10909 -8539
rect 10843 -8582 10859 -8548
rect 10893 -8582 10909 -8548
rect 10843 -8616 10909 -8582
rect 10843 -8650 10859 -8616
rect 10893 -8650 10909 -8616
rect 10843 -8699 10909 -8650
rect 10999 -8547 11049 -8505
rect 10999 -8581 11015 -8547
rect 10999 -8615 11049 -8581
rect 10999 -8649 11015 -8615
rect 10999 -8665 11049 -8649
rect 11101 -8548 11171 -8436
rect 11236 -8464 11306 -8435
rect 11236 -8498 11430 -8464
rect 11101 -8582 11119 -8548
rect 11153 -8582 11171 -8548
rect 11101 -8616 11171 -8582
rect 11101 -8650 11119 -8616
rect 11153 -8650 11171 -8616
rect 11101 -8665 11171 -8650
rect 11261 -8548 11327 -8532
rect 11261 -8582 11277 -8548
rect 11311 -8582 11327 -8548
rect 11261 -8616 11327 -8582
rect 11261 -8650 11277 -8616
rect 11311 -8650 11327 -8616
rect 11261 -8699 11327 -8650
rect 11361 -8548 11430 -8498
rect 11361 -8582 11377 -8548
rect 11411 -8582 11430 -8548
rect 11361 -8616 11430 -8582
rect 11361 -8650 11377 -8616
rect 11411 -8650 11430 -8616
rect 11361 -8665 11430 -8650
rect 11464 -8501 11522 -8466
rect 11464 -8535 11476 -8501
rect 11510 -8535 11522 -8501
rect 11464 -8594 11522 -8535
rect 11464 -8628 11476 -8594
rect 11510 -8628 11522 -8594
rect 11464 -8699 11522 -8628
rect 11648 -8481 11798 -8411
rect 11832 -8413 11982 -8343
rect 11832 -8447 11928 -8413
rect 11962 -8447 11982 -8413
rect 13672 -8362 13735 -8325
rect 13672 -8396 13685 -8362
rect 13719 -8387 13735 -8362
rect 13672 -8421 13692 -8396
rect 13726 -8421 13735 -8387
rect 13672 -8437 13735 -8421
rect 13769 -8387 13819 -8278
rect 13853 -8244 13905 -8189
rect 13853 -8278 13862 -8244
rect 13896 -8278 13905 -8244
rect 13853 -8294 13905 -8278
rect 13941 -8244 13991 -8225
rect 13941 -8278 13948 -8244
rect 13982 -8278 13991 -8244
rect 13941 -8387 13991 -8278
rect 14025 -8244 14077 -8189
rect 14025 -8278 14034 -8244
rect 14068 -8278 14077 -8244
rect 14025 -8301 14077 -8278
rect 14111 -8244 14163 -8228
rect 14111 -8278 14120 -8244
rect 14154 -8278 14163 -8244
rect 14111 -8319 14163 -8278
rect 14197 -8235 14249 -8189
rect 14197 -8269 14206 -8235
rect 14240 -8269 14249 -8235
rect 14197 -8285 14249 -8269
rect 14283 -8244 14335 -8228
rect 14283 -8278 14292 -8244
rect 14326 -8278 14335 -8244
rect 14283 -8319 14335 -8278
rect 14369 -8235 14421 -8189
rect 14369 -8269 14378 -8235
rect 14412 -8269 14421 -8235
rect 14369 -8285 14421 -8269
rect 14455 -8244 14507 -8228
rect 14455 -8278 14464 -8244
rect 14498 -8278 14507 -8244
rect 14455 -8319 14507 -8278
rect 14541 -8235 14590 -8189
rect 14541 -8269 14550 -8235
rect 14584 -8269 14590 -8235
rect 14541 -8285 14590 -8269
rect 14624 -8244 14679 -8228
rect 14624 -8278 14636 -8244
rect 14670 -8278 14679 -8244
rect 14624 -8319 14679 -8278
rect 14713 -8235 14762 -8189
rect 14713 -8269 14722 -8235
rect 14756 -8269 14762 -8235
rect 14713 -8285 14762 -8269
rect 14796 -8244 14848 -8228
rect 14796 -8278 14807 -8244
rect 14841 -8278 14848 -8244
rect 14796 -8319 14848 -8278
rect 14884 -8235 14934 -8189
rect 14884 -8269 14893 -8235
rect 14927 -8269 14934 -8235
rect 14884 -8285 14934 -8269
rect 14968 -8244 15020 -8228
rect 14968 -8278 14979 -8244
rect 15013 -8278 15020 -8244
rect 14968 -8319 15020 -8278
rect 15056 -8235 15106 -8189
rect 15056 -8269 15065 -8235
rect 15099 -8269 15106 -8235
rect 15056 -8285 15106 -8269
rect 15140 -8244 15192 -8228
rect 15140 -8278 15151 -8244
rect 15185 -8278 15192 -8244
rect 15140 -8319 15192 -8278
rect 15228 -8235 15280 -8189
rect 15228 -8269 15237 -8235
rect 15271 -8269 15280 -8235
rect 15228 -8285 15280 -8269
rect 15314 -8244 15366 -8228
rect 15314 -8278 15323 -8244
rect 15357 -8278 15366 -8244
rect 15314 -8319 15366 -8278
rect 15400 -8235 15460 -8189
rect 15400 -8269 15409 -8235
rect 15443 -8269 15460 -8235
rect 15400 -8285 15460 -8269
rect 15512 -8283 15570 -8189
rect 15512 -8317 15524 -8283
rect 15558 -8317 15570 -8283
rect 14111 -8344 15460 -8319
rect 15512 -8334 15570 -8317
rect 15605 -8250 16674 -8189
rect 15605 -8284 15622 -8250
rect 15656 -8284 16622 -8250
rect 16656 -8284 16674 -8250
rect 15605 -8343 16674 -8284
rect 14111 -8353 15248 -8344
rect 15227 -8378 15248 -8353
rect 15282 -8345 15460 -8344
rect 15282 -8378 15340 -8345
rect 15227 -8379 15340 -8378
rect 15374 -8379 15460 -8345
rect 13769 -8421 14119 -8387
rect 14153 -8421 14187 -8387
rect 14221 -8421 14255 -8387
rect 14289 -8421 14323 -8387
rect 14357 -8421 14391 -8387
rect 14425 -8421 14459 -8387
rect 14493 -8421 14527 -8387
rect 14561 -8421 14595 -8387
rect 14629 -8421 14663 -8387
rect 14697 -8421 14731 -8387
rect 14765 -8421 14799 -8387
rect 14833 -8421 14867 -8387
rect 14901 -8421 14935 -8387
rect 14969 -8421 15003 -8387
rect 15037 -8421 15071 -8387
rect 15105 -8421 15139 -8387
rect 15173 -8421 15193 -8387
rect 13769 -8437 15193 -8421
rect 11648 -8521 11982 -8481
rect 11648 -8555 11666 -8521
rect 11700 -8555 11930 -8521
rect 11964 -8555 11982 -8521
rect 11648 -8623 11982 -8555
rect 11648 -8657 11666 -8623
rect 11700 -8657 11930 -8623
rect 11964 -8657 11982 -8623
rect 11648 -8699 11982 -8657
rect 13580 -8501 13638 -8466
rect 13580 -8535 13592 -8501
rect 13626 -8535 13638 -8501
rect 13580 -8594 13638 -8535
rect 13580 -8628 13592 -8594
rect 13626 -8628 13638 -8594
rect 13580 -8699 13638 -8628
rect 13674 -8555 13733 -8537
rect 13674 -8589 13690 -8555
rect 13724 -8589 13733 -8555
rect 13674 -8623 13733 -8589
rect 13674 -8657 13690 -8623
rect 13724 -8657 13733 -8623
rect 13674 -8699 13733 -8657
rect 13769 -8547 13818 -8437
rect 13769 -8581 13776 -8547
rect 13810 -8581 13818 -8547
rect 13769 -8615 13818 -8581
rect 13769 -8649 13776 -8615
rect 13810 -8649 13818 -8615
rect 13769 -8665 13818 -8649
rect 13853 -8555 13905 -8537
rect 13853 -8589 13862 -8555
rect 13896 -8589 13905 -8555
rect 13853 -8623 13905 -8589
rect 13853 -8657 13862 -8623
rect 13896 -8657 13905 -8623
rect 13853 -8699 13905 -8657
rect 13941 -8539 13991 -8437
rect 15227 -8440 15460 -8379
rect 15227 -8471 15248 -8440
rect 14111 -8474 15248 -8471
rect 15282 -8474 15341 -8440
rect 15375 -8474 15460 -8440
rect 15605 -8411 15686 -8377
rect 15720 -8411 15814 -8377
rect 15848 -8411 15942 -8377
rect 15976 -8411 16070 -8377
rect 16104 -8411 16124 -8377
rect 14111 -8493 15460 -8474
rect 14111 -8527 14120 -8493
rect 14154 -8519 14292 -8493
rect 14154 -8527 14163 -8519
rect 13941 -8573 13948 -8539
rect 13982 -8573 13991 -8539
rect 13941 -8607 13991 -8573
rect 13941 -8641 13948 -8607
rect 13982 -8641 13991 -8607
rect 13941 -8664 13991 -8641
rect 14025 -8555 14077 -8539
rect 14025 -8589 14034 -8555
rect 14068 -8589 14077 -8555
rect 14025 -8623 14077 -8589
rect 14025 -8657 14034 -8623
rect 14068 -8657 14077 -8623
rect 14025 -8698 14077 -8657
rect 14111 -8579 14163 -8527
rect 14283 -8527 14292 -8519
rect 14326 -8519 14464 -8493
rect 14326 -8527 14335 -8519
rect 14111 -8613 14120 -8579
rect 14154 -8613 14163 -8579
rect 14111 -8664 14163 -8613
rect 14197 -8599 14249 -8553
rect 14197 -8633 14206 -8599
rect 14240 -8633 14249 -8599
rect 14197 -8698 14249 -8633
rect 14283 -8579 14335 -8527
rect 14455 -8527 14464 -8519
rect 14498 -8519 14636 -8493
rect 14498 -8527 14507 -8519
rect 14283 -8613 14292 -8579
rect 14326 -8613 14335 -8579
rect 14283 -8664 14335 -8613
rect 14369 -8599 14421 -8553
rect 14369 -8633 14378 -8599
rect 14412 -8633 14421 -8599
rect 14369 -8698 14421 -8633
rect 14455 -8579 14507 -8527
rect 14627 -8527 14636 -8519
rect 14670 -8519 14807 -8493
rect 14670 -8527 14679 -8519
rect 14455 -8613 14464 -8579
rect 14498 -8613 14507 -8579
rect 14455 -8664 14507 -8613
rect 14541 -8599 14593 -8553
rect 14541 -8633 14550 -8599
rect 14584 -8633 14593 -8599
rect 14541 -8698 14593 -8633
rect 14627 -8579 14679 -8527
rect 14796 -8527 14807 -8519
rect 14841 -8519 14979 -8493
rect 14841 -8527 14848 -8519
rect 14627 -8613 14636 -8579
rect 14670 -8613 14679 -8579
rect 14627 -8664 14679 -8613
rect 14713 -8599 14762 -8553
rect 14713 -8633 14722 -8599
rect 14756 -8633 14762 -8599
rect 14713 -8698 14762 -8633
rect 14796 -8579 14848 -8527
rect 14968 -8527 14979 -8519
rect 15013 -8519 15151 -8493
rect 15013 -8527 15020 -8519
rect 14796 -8613 14807 -8579
rect 14841 -8613 14848 -8579
rect 14796 -8664 14848 -8613
rect 14885 -8599 14934 -8553
rect 14885 -8633 14893 -8599
rect 14927 -8633 14934 -8599
rect 14885 -8698 14934 -8633
rect 14968 -8579 15020 -8527
rect 15140 -8527 15151 -8519
rect 15185 -8516 15323 -8493
rect 15185 -8527 15192 -8516
rect 14968 -8613 14979 -8579
rect 15013 -8613 15020 -8579
rect 14968 -8664 15020 -8613
rect 15057 -8599 15106 -8553
rect 15057 -8633 15065 -8599
rect 15099 -8633 15106 -8599
rect 15057 -8698 15106 -8633
rect 15140 -8579 15192 -8527
rect 15314 -8527 15323 -8516
rect 15357 -8516 15460 -8493
rect 15512 -8501 15570 -8466
rect 15357 -8527 15372 -8516
rect 15140 -8613 15151 -8579
rect 15185 -8613 15192 -8579
rect 15140 -8664 15192 -8613
rect 15229 -8599 15280 -8553
rect 15229 -8633 15237 -8599
rect 15271 -8633 15280 -8599
rect 15229 -8698 15280 -8633
rect 15314 -8579 15372 -8527
rect 15512 -8535 15524 -8501
rect 15558 -8535 15570 -8501
rect 15314 -8613 15323 -8579
rect 15357 -8613 15372 -8579
rect 15314 -8664 15372 -8613
rect 15406 -8599 15460 -8550
rect 15406 -8633 15409 -8599
rect 15443 -8633 15460 -8599
rect 14025 -8699 15280 -8698
rect 15406 -8699 15460 -8633
rect 15512 -8594 15570 -8535
rect 15512 -8628 15524 -8594
rect 15558 -8628 15570 -8594
rect 15512 -8699 15570 -8628
rect 15605 -8481 16124 -8411
rect 16158 -8413 16674 -8343
rect 16158 -8447 16178 -8413
rect 16212 -8447 16306 -8413
rect 16340 -8447 16434 -8413
rect 16468 -8447 16562 -8413
rect 16596 -8447 16674 -8413
rect 15605 -8521 16674 -8481
rect 15605 -8555 15622 -8521
rect 15656 -8555 16622 -8521
rect 16656 -8555 16674 -8521
rect 15605 -8623 16674 -8555
rect 15605 -8657 15622 -8623
rect 15656 -8657 16622 -8623
rect 16656 -8657 16674 -8623
rect 15605 -8699 16674 -8657
rect -2997 -8733 -2968 -8699
rect -2934 -8733 -2876 -8699
rect -2842 -8733 -2784 -8699
rect -2750 -8733 -2692 -8699
rect -2658 -8733 -2600 -8699
rect -2566 -8733 -2508 -8699
rect -2474 -8733 -2416 -8699
rect -2382 -8733 -2324 -8699
rect -2290 -8733 -2232 -8699
rect -2198 -8733 -2140 -8699
rect -2106 -8733 -2048 -8699
rect -2014 -8733 -1956 -8699
rect -1922 -8733 -1864 -8699
rect -1830 -8733 -1772 -8699
rect -1738 -8733 -1680 -8699
rect -1646 -8733 -1588 -8699
rect -1554 -8733 -1496 -8699
rect -1462 -8733 -1404 -8699
rect -1370 -8733 -1312 -8699
rect -1278 -8733 -1220 -8699
rect -1186 -8733 -1128 -8699
rect -1094 -8733 -1036 -8699
rect -1002 -8733 -944 -8699
rect -910 -8733 -852 -8699
rect -818 -8733 -760 -8699
rect -726 -8733 -668 -8699
rect -634 -8733 -576 -8699
rect -542 -8733 -484 -8699
rect -450 -8733 -392 -8699
rect -358 -8733 -300 -8699
rect -266 -8733 -208 -8699
rect -174 -8733 -116 -8699
rect -82 -8733 -24 -8699
rect 10 -8733 68 -8699
rect 102 -8733 160 -8699
rect 194 -8733 252 -8699
rect 286 -8733 344 -8699
rect 378 -8733 436 -8699
rect 470 -8733 528 -8699
rect 562 -8733 620 -8699
rect 654 -8733 712 -8699
rect 746 -8733 804 -8699
rect 838 -8733 896 -8699
rect 930 -8733 988 -8699
rect 1022 -8733 1080 -8699
rect 1114 -8733 1172 -8699
rect 1206 -8733 1264 -8699
rect 1298 -8733 1356 -8699
rect 1390 -8733 1448 -8699
rect 1482 -8733 1540 -8699
rect 1574 -8733 1632 -8699
rect 1666 -8733 1724 -8699
rect 1758 -8733 1816 -8699
rect 1850 -8733 1908 -8699
rect 1942 -8733 2000 -8699
rect 2034 -8733 2092 -8699
rect 2126 -8733 2184 -8699
rect 2218 -8733 2276 -8699
rect 2310 -8733 2368 -8699
rect 2402 -8733 2460 -8699
rect 2494 -8733 2552 -8699
rect 2586 -8733 2644 -8699
rect 2678 -8733 2736 -8699
rect 2770 -8733 2828 -8699
rect 2862 -8733 2920 -8699
rect 2954 -8733 3012 -8699
rect 3046 -8733 3104 -8699
rect 3138 -8733 3196 -8699
rect 3230 -8733 3288 -8699
rect 3322 -8733 3380 -8699
rect 3414 -8733 3472 -8699
rect 3506 -8733 3564 -8699
rect 3598 -8733 3656 -8699
rect 3690 -8733 3748 -8699
rect 3782 -8733 3840 -8699
rect 3874 -8733 3932 -8699
rect 3966 -8733 4024 -8699
rect 4058 -8733 4116 -8699
rect 4150 -8733 4208 -8699
rect 4242 -8733 4300 -8699
rect 4334 -8733 4392 -8699
rect 4426 -8733 4484 -8699
rect 4518 -8733 4576 -8699
rect 4610 -8733 4668 -8699
rect 4702 -8733 4760 -8699
rect 4794 -8733 4852 -8699
rect 4886 -8733 4944 -8699
rect 4978 -8733 5036 -8699
rect 5070 -8733 5128 -8699
rect 5162 -8733 5220 -8699
rect 5254 -8733 5312 -8699
rect 5346 -8733 5404 -8699
rect 5438 -8733 5496 -8699
rect 5530 -8733 5588 -8699
rect 5622 -8733 5680 -8699
rect 5714 -8733 5772 -8699
rect 5806 -8733 5864 -8699
rect 5898 -8733 5956 -8699
rect 5990 -8733 6048 -8699
rect 6082 -8733 6140 -8699
rect 6174 -8733 6232 -8699
rect 6266 -8733 6324 -8699
rect 6358 -8733 6416 -8699
rect 6450 -8733 6508 -8699
rect 6542 -8733 6600 -8699
rect 6634 -8733 6692 -8699
rect 6726 -8733 6784 -8699
rect 6818 -8733 6876 -8699
rect 6910 -8733 6968 -8699
rect 7002 -8733 7060 -8699
rect 7094 -8733 7152 -8699
rect 7186 -8733 7244 -8699
rect 7278 -8733 7336 -8699
rect 7370 -8733 7428 -8699
rect 7462 -8733 7520 -8699
rect 7554 -8733 7612 -8699
rect 7646 -8733 7704 -8699
rect 7738 -8733 7796 -8699
rect 7830 -8733 7888 -8699
rect 7922 -8733 7980 -8699
rect 8014 -8733 8072 -8699
rect 8106 -8733 8164 -8699
rect 8198 -8733 8256 -8699
rect 8290 -8733 8348 -8699
rect 8382 -8733 8440 -8699
rect 8474 -8733 8532 -8699
rect 8566 -8733 8624 -8699
rect 8658 -8733 8716 -8699
rect 8750 -8733 8808 -8699
rect 8842 -8733 8900 -8699
rect 8934 -8733 8992 -8699
rect 9026 -8733 9084 -8699
rect 9118 -8733 9176 -8699
rect 9210 -8733 9268 -8699
rect 9302 -8733 9360 -8699
rect 9394 -8733 9452 -8699
rect 9486 -8733 9544 -8699
rect 9578 -8733 9636 -8699
rect 9670 -8733 9728 -8699
rect 9762 -8733 9820 -8699
rect 9854 -8733 9912 -8699
rect 9946 -8733 10004 -8699
rect 10038 -8733 10096 -8699
rect 10130 -8733 10188 -8699
rect 10222 -8733 10280 -8699
rect 10314 -8733 10372 -8699
rect 10406 -8733 10464 -8699
rect 10498 -8733 10556 -8699
rect 10590 -8733 10648 -8699
rect 10682 -8733 10740 -8699
rect 10774 -8733 10832 -8699
rect 10866 -8733 10924 -8699
rect 10958 -8733 11016 -8699
rect 11050 -8733 11108 -8699
rect 11142 -8733 11200 -8699
rect 11234 -8733 11292 -8699
rect 11326 -8733 11384 -8699
rect 11418 -8733 11476 -8699
rect 11510 -8733 11568 -8699
rect 11602 -8733 11660 -8699
rect 11694 -8733 11752 -8699
rect 11786 -8733 11844 -8699
rect 11878 -8733 11936 -8699
rect 11970 -8733 12028 -8699
rect 12062 -8733 12120 -8699
rect 12154 -8733 12212 -8699
rect 12246 -8733 12304 -8699
rect 12338 -8733 12396 -8699
rect 12430 -8733 12488 -8699
rect 12522 -8733 12580 -8699
rect 12614 -8733 12672 -8699
rect 12706 -8733 12764 -8699
rect 12798 -8733 12856 -8699
rect 12890 -8733 12948 -8699
rect 12982 -8733 13040 -8699
rect 13074 -8733 13132 -8699
rect 13166 -8733 13224 -8699
rect 13258 -8733 13316 -8699
rect 13350 -8733 13408 -8699
rect 13442 -8733 13500 -8699
rect 13534 -8733 13592 -8699
rect 13626 -8733 13684 -8699
rect 13718 -8733 13776 -8699
rect 13810 -8733 13868 -8699
rect 13902 -8733 13960 -8699
rect 13994 -8733 14052 -8699
rect 14086 -8733 14144 -8699
rect 14178 -8733 14236 -8699
rect 14270 -8733 14328 -8699
rect 14362 -8733 14420 -8699
rect 14454 -8733 14512 -8699
rect 14546 -8733 14604 -8699
rect 14638 -8733 14696 -8699
rect 14730 -8733 14788 -8699
rect 14822 -8733 14880 -8699
rect 14914 -8733 14972 -8699
rect 15006 -8733 15064 -8699
rect 15098 -8733 15156 -8699
rect 15190 -8733 15248 -8699
rect 15282 -8733 15340 -8699
rect 15374 -8733 15432 -8699
rect 15466 -8733 15524 -8699
rect 15558 -8733 15616 -8699
rect 15650 -8733 15708 -8699
rect 15742 -8733 15800 -8699
rect 15834 -8733 15892 -8699
rect 15926 -8733 15984 -8699
rect 16018 -8733 16076 -8699
rect 16110 -8733 16168 -8699
rect 16202 -8733 16260 -8699
rect 16294 -8733 16352 -8699
rect 16386 -8733 16444 -8699
rect 16478 -8733 16536 -8699
rect 16570 -8733 16628 -8699
rect 16662 -8733 16691 -8699
rect -2980 -8775 -2278 -8733
rect -2980 -8809 -2962 -8775
rect -2928 -8809 -2330 -8775
rect -2296 -8809 -2278 -8775
rect -2980 -8877 -2278 -8809
rect -2980 -8911 -2962 -8877
rect -2928 -8911 -2330 -8877
rect -2296 -8911 -2278 -8877
rect -2980 -8951 -2278 -8911
rect -2980 -9019 -2902 -8985
rect -2868 -9019 -2803 -8985
rect -2769 -9019 -2704 -8985
rect -2670 -9019 -2650 -8985
rect -2980 -9089 -2650 -9019
rect -2616 -9021 -2278 -8951
rect -2244 -8804 -2186 -8733
rect -2244 -8838 -2232 -8804
rect -2198 -8838 -2186 -8804
rect -2244 -8897 -2186 -8838
rect -2244 -8931 -2232 -8897
rect -2198 -8931 -2186 -8897
rect -2244 -8966 -2186 -8931
rect -1600 -8775 -898 -8733
rect -1600 -8809 -1582 -8775
rect -1548 -8809 -950 -8775
rect -916 -8809 -898 -8775
rect -1600 -8877 -898 -8809
rect -1600 -8911 -1582 -8877
rect -1548 -8911 -950 -8877
rect -916 -8911 -898 -8877
rect -1600 -8951 -898 -8911
rect -864 -8775 -162 -8733
rect -864 -8809 -846 -8775
rect -812 -8809 -214 -8775
rect -180 -8809 -162 -8775
rect -864 -8877 -162 -8809
rect -864 -8911 -846 -8877
rect -812 -8911 -214 -8877
rect -180 -8911 -162 -8877
rect -864 -8951 -162 -8911
rect -2616 -9055 -2596 -9021
rect -2562 -9055 -2493 -9021
rect -2459 -9055 -2390 -9021
rect -2356 -9055 -2278 -9021
rect -1600 -9019 -1522 -8985
rect -1488 -9019 -1423 -8985
rect -1389 -9019 -1324 -8985
rect -1290 -9019 -1270 -8985
rect -1600 -9089 -1270 -9019
rect -1236 -9021 -898 -8951
rect -1236 -9055 -1216 -9021
rect -1182 -9055 -1113 -9021
rect -1079 -9055 -1010 -9021
rect -976 -9055 -898 -9021
rect -864 -9019 -786 -8985
rect -752 -9019 -687 -8985
rect -653 -9019 -588 -8985
rect -554 -9019 -534 -8985
rect -864 -9089 -534 -9019
rect -500 -9021 -162 -8951
rect -128 -8804 -70 -8733
rect -128 -8838 -116 -8804
rect -82 -8838 -70 -8804
rect -128 -8897 -70 -8838
rect -128 -8931 -116 -8897
rect -82 -8931 -70 -8897
rect -128 -8966 -70 -8931
rect -36 -8775 298 -8733
rect -36 -8809 -18 -8775
rect 16 -8809 246 -8775
rect 280 -8809 298 -8775
rect -36 -8877 298 -8809
rect -36 -8911 -18 -8877
rect 16 -8911 246 -8877
rect 280 -8911 298 -8877
rect -36 -8951 298 -8911
rect 332 -8804 390 -8733
rect 332 -8838 344 -8804
rect 378 -8838 390 -8804
rect 332 -8897 390 -8838
rect 332 -8931 344 -8897
rect 378 -8931 390 -8897
rect -500 -9055 -480 -9021
rect -446 -9055 -377 -9021
rect -343 -9055 -274 -9021
rect -240 -9055 -162 -9021
rect -36 -9021 114 -8951
rect 332 -8966 390 -8931
rect 424 -8782 493 -8767
rect 424 -8816 443 -8782
rect 477 -8816 493 -8782
rect 424 -8850 493 -8816
rect 424 -8884 443 -8850
rect 477 -8884 493 -8850
rect 424 -8934 493 -8884
rect 527 -8782 593 -8733
rect 527 -8816 543 -8782
rect 577 -8816 593 -8782
rect 527 -8850 593 -8816
rect 527 -8884 543 -8850
rect 577 -8884 593 -8850
rect 527 -8900 593 -8884
rect 683 -8782 753 -8767
rect 683 -8816 701 -8782
rect 735 -8816 753 -8782
rect 683 -8850 753 -8816
rect 683 -8884 701 -8850
rect 735 -8884 753 -8850
rect 424 -8968 618 -8934
rect -36 -9055 -16 -9021
rect 18 -9055 114 -9021
rect 148 -9019 244 -8985
rect 278 -9019 298 -8985
rect 548 -8997 618 -8968
rect 683 -8996 753 -8884
rect 805 -8783 855 -8767
rect 839 -8817 855 -8783
rect 805 -8851 855 -8817
rect 839 -8885 855 -8851
rect 805 -8927 855 -8885
rect 945 -8782 1011 -8733
rect 945 -8816 961 -8782
rect 995 -8816 1011 -8782
rect 945 -8850 1011 -8816
rect 945 -8884 961 -8850
rect 995 -8884 1011 -8850
rect 945 -8893 1011 -8884
rect 1045 -8783 1126 -8767
rect 1045 -8817 1059 -8783
rect 1093 -8817 1126 -8783
rect 1045 -8851 1126 -8817
rect 1045 -8885 1059 -8851
rect 1093 -8885 1126 -8851
rect 1045 -8922 1126 -8885
rect 805 -8961 923 -8927
rect 889 -8995 923 -8961
rect 148 -9089 298 -9019
rect 424 -9008 514 -9002
rect 424 -9042 432 -9008
rect 466 -9011 514 -9008
rect 424 -9045 464 -9042
rect 498 -9045 514 -9011
rect 548 -9011 634 -8997
rect 548 -9045 584 -9011
rect 618 -9045 634 -9011
rect 548 -9055 634 -9045
rect 683 -9011 855 -8996
rect 683 -9045 805 -9011
rect 839 -9045 855 -9011
rect 683 -9046 855 -9045
rect 889 -9011 1042 -8995
rect 889 -9045 1005 -9011
rect 1039 -9045 1042 -9011
rect 548 -9079 618 -9055
rect -2980 -9148 -2278 -9089
rect -2980 -9182 -2962 -9148
rect -2928 -9182 -2330 -9148
rect -2296 -9182 -2278 -9148
rect -2980 -9243 -2278 -9182
rect -2244 -9115 -2186 -9098
rect -2244 -9149 -2232 -9115
rect -2198 -9149 -2186 -9115
rect -2244 -9243 -2186 -9149
rect -1600 -9148 -898 -9089
rect -1600 -9182 -1582 -9148
rect -1548 -9182 -950 -9148
rect -916 -9182 -898 -9148
rect -1600 -9243 -898 -9182
rect -864 -9148 -162 -9089
rect -864 -9182 -846 -9148
rect -812 -9182 -214 -9148
rect -180 -9182 -162 -9148
rect -864 -9243 -162 -9182
rect -128 -9115 -70 -9098
rect -128 -9149 -116 -9115
rect -82 -9149 -70 -9115
rect -128 -9243 -70 -9149
rect -36 -9141 298 -9089
rect -36 -9175 -18 -9141
rect 16 -9175 246 -9141
rect 280 -9175 298 -9141
rect -36 -9243 298 -9175
rect 332 -9115 390 -9098
rect 332 -9149 344 -9115
rect 378 -9149 390 -9115
rect 332 -9243 390 -9149
rect 424 -9113 618 -9079
rect 424 -9156 490 -9113
rect 424 -9190 443 -9156
rect 477 -9190 490 -9156
rect 424 -9209 490 -9190
rect 524 -9156 590 -9147
rect 524 -9190 540 -9156
rect 574 -9190 590 -9156
rect 524 -9243 590 -9190
rect 683 -9156 753 -9046
rect 889 -9061 1042 -9045
rect 1076 -9005 1126 -8922
rect 1160 -8804 1218 -8733
rect 1160 -8838 1172 -8804
rect 1206 -8838 1218 -8804
rect 1160 -8897 1218 -8838
rect 1160 -8931 1172 -8897
rect 1206 -8931 1218 -8897
rect 1160 -8966 1218 -8931
rect 1252 -8775 1586 -8733
rect 1252 -8809 1270 -8775
rect 1304 -8809 1534 -8775
rect 1568 -8809 1586 -8775
rect 1252 -8877 1586 -8809
rect 1252 -8911 1270 -8877
rect 1304 -8911 1534 -8877
rect 1568 -8911 1586 -8877
rect 1252 -8951 1586 -8911
rect 1620 -8804 1678 -8733
rect 1620 -8838 1632 -8804
rect 1666 -8838 1678 -8804
rect 1620 -8897 1678 -8838
rect 1620 -8931 1632 -8897
rect 1666 -8931 1678 -8897
rect 1076 -9039 1082 -9005
rect 1116 -9039 1126 -9005
rect 889 -9080 923 -9061
rect 683 -9190 700 -9156
rect 734 -9190 753 -9156
rect 683 -9209 753 -9190
rect 805 -9114 923 -9080
rect 805 -9156 855 -9114
rect 1076 -9132 1126 -9039
rect 1252 -9021 1402 -8951
rect 1620 -8966 1678 -8931
rect 1712 -8775 2414 -8733
rect 1712 -8809 1730 -8775
rect 1764 -8809 2362 -8775
rect 2396 -8809 2414 -8775
rect 1712 -8877 2414 -8809
rect 1712 -8911 1730 -8877
rect 1764 -8911 2362 -8877
rect 2396 -8911 2414 -8877
rect 1712 -8951 2414 -8911
rect 1252 -9055 1272 -9021
rect 1306 -9055 1402 -9021
rect 1436 -9019 1532 -8985
rect 1566 -9019 1586 -8985
rect 1436 -9089 1586 -9019
rect 839 -9190 855 -9156
rect 805 -9209 855 -9190
rect 945 -9156 1011 -9140
rect 945 -9190 961 -9156
rect 995 -9190 1011 -9156
rect 945 -9243 1011 -9190
rect 1045 -9156 1126 -9132
rect 1045 -9190 1059 -9156
rect 1093 -9190 1126 -9156
rect 1045 -9209 1126 -9190
rect 1160 -9115 1218 -9098
rect 1160 -9149 1172 -9115
rect 1206 -9149 1218 -9115
rect 1160 -9243 1218 -9149
rect 1252 -9141 1586 -9089
rect 1712 -9019 1790 -8985
rect 1824 -9019 1889 -8985
rect 1923 -9019 1988 -8985
rect 2022 -9019 2042 -8985
rect 1712 -9089 2042 -9019
rect 2076 -9021 2414 -8951
rect 2448 -8804 2506 -8733
rect 2448 -8838 2460 -8804
rect 2494 -8838 2506 -8804
rect 2448 -8897 2506 -8838
rect 2448 -8931 2460 -8897
rect 2494 -8931 2506 -8897
rect 2448 -8966 2506 -8931
rect 2540 -8775 2874 -8733
rect 2540 -8809 2558 -8775
rect 2592 -8809 2822 -8775
rect 2856 -8809 2874 -8775
rect 2540 -8877 2874 -8809
rect 2540 -8911 2558 -8877
rect 2592 -8911 2822 -8877
rect 2856 -8911 2874 -8877
rect 2540 -8951 2874 -8911
rect 2908 -8804 2966 -8733
rect 2908 -8838 2920 -8804
rect 2954 -8838 2966 -8804
rect 2908 -8897 2966 -8838
rect 2908 -8931 2920 -8897
rect 2954 -8931 2966 -8897
rect 2076 -9055 2096 -9021
rect 2130 -9055 2199 -9021
rect 2233 -9055 2302 -9021
rect 2336 -9055 2414 -9021
rect 2540 -9021 2690 -8951
rect 2908 -8966 2966 -8931
rect 3000 -8782 3069 -8767
rect 3000 -8816 3019 -8782
rect 3053 -8816 3069 -8782
rect 3000 -8850 3069 -8816
rect 3000 -8884 3019 -8850
rect 3053 -8884 3069 -8850
rect 3000 -8934 3069 -8884
rect 3103 -8782 3169 -8733
rect 3103 -8816 3119 -8782
rect 3153 -8816 3169 -8782
rect 3103 -8850 3169 -8816
rect 3103 -8884 3119 -8850
rect 3153 -8884 3169 -8850
rect 3103 -8900 3169 -8884
rect 3259 -8782 3329 -8767
rect 3259 -8816 3277 -8782
rect 3311 -8816 3329 -8782
rect 3259 -8850 3329 -8816
rect 3259 -8884 3277 -8850
rect 3311 -8884 3329 -8850
rect 3000 -8968 3194 -8934
rect 2540 -9055 2560 -9021
rect 2594 -9055 2690 -9021
rect 2724 -9019 2820 -8985
rect 2854 -9019 2874 -8985
rect 3124 -8997 3194 -8968
rect 3259 -8996 3329 -8884
rect 3381 -8783 3431 -8767
rect 3415 -8817 3431 -8783
rect 3381 -8851 3431 -8817
rect 3415 -8885 3431 -8851
rect 3381 -8927 3431 -8885
rect 3521 -8782 3587 -8733
rect 3521 -8816 3537 -8782
rect 3571 -8816 3587 -8782
rect 3521 -8850 3587 -8816
rect 3521 -8884 3537 -8850
rect 3571 -8884 3587 -8850
rect 3521 -8893 3587 -8884
rect 3621 -8783 3702 -8767
rect 3621 -8817 3635 -8783
rect 3669 -8817 3702 -8783
rect 3621 -8851 3702 -8817
rect 3621 -8885 3635 -8851
rect 3669 -8885 3702 -8851
rect 3621 -8922 3702 -8885
rect 3381 -8961 3499 -8927
rect 3465 -8995 3499 -8961
rect 2724 -9089 2874 -9019
rect 3000 -9005 3090 -9002
rect 3000 -9011 3042 -9005
rect 3000 -9045 3040 -9011
rect 3076 -9039 3090 -9005
rect 3074 -9045 3090 -9039
rect 3124 -9011 3210 -8997
rect 3124 -9045 3160 -9011
rect 3194 -9045 3210 -9011
rect 3124 -9055 3210 -9045
rect 3259 -9011 3431 -8996
rect 3259 -9045 3381 -9011
rect 3415 -9045 3431 -9011
rect 3259 -9046 3431 -9045
rect 3465 -9011 3618 -8995
rect 3465 -9045 3581 -9011
rect 3615 -9045 3618 -9011
rect 3124 -9079 3194 -9055
rect 1252 -9175 1270 -9141
rect 1304 -9175 1534 -9141
rect 1568 -9175 1586 -9141
rect 1252 -9243 1586 -9175
rect 1620 -9115 1678 -9098
rect 1620 -9149 1632 -9115
rect 1666 -9149 1678 -9115
rect 1620 -9243 1678 -9149
rect 1712 -9148 2414 -9089
rect 1712 -9182 1730 -9148
rect 1764 -9182 2362 -9148
rect 2396 -9182 2414 -9148
rect 1712 -9243 2414 -9182
rect 2448 -9115 2506 -9098
rect 2448 -9149 2460 -9115
rect 2494 -9149 2506 -9115
rect 2448 -9243 2506 -9149
rect 2540 -9141 2874 -9089
rect 2540 -9175 2558 -9141
rect 2592 -9175 2822 -9141
rect 2856 -9175 2874 -9141
rect 2540 -9243 2874 -9175
rect 2908 -9115 2966 -9098
rect 2908 -9149 2920 -9115
rect 2954 -9149 2966 -9115
rect 2908 -9243 2966 -9149
rect 3000 -9113 3194 -9079
rect 3000 -9156 3066 -9113
rect 3000 -9190 3019 -9156
rect 3053 -9190 3066 -9156
rect 3000 -9209 3066 -9190
rect 3100 -9156 3166 -9147
rect 3100 -9190 3116 -9156
rect 3150 -9190 3166 -9156
rect 3100 -9243 3166 -9190
rect 3259 -9156 3329 -9046
rect 3465 -9061 3618 -9045
rect 3652 -9005 3702 -8922
rect 3736 -8804 3794 -8733
rect 3736 -8838 3748 -8804
rect 3782 -8838 3794 -8804
rect 3736 -8897 3794 -8838
rect 3736 -8931 3748 -8897
rect 3782 -8931 3794 -8897
rect 3736 -8966 3794 -8931
rect 3828 -8775 4162 -8733
rect 3828 -8809 3846 -8775
rect 3880 -8809 4110 -8775
rect 4144 -8809 4162 -8775
rect 3828 -8877 4162 -8809
rect 3828 -8911 3846 -8877
rect 3880 -8911 4110 -8877
rect 4144 -8911 4162 -8877
rect 3828 -8951 4162 -8911
rect 4196 -8804 4254 -8733
rect 4196 -8838 4208 -8804
rect 4242 -8838 4254 -8804
rect 4196 -8897 4254 -8838
rect 4196 -8931 4208 -8897
rect 4242 -8931 4254 -8897
rect 3652 -9039 3656 -9005
rect 3690 -9039 3702 -9005
rect 3465 -9080 3499 -9061
rect 3259 -9190 3276 -9156
rect 3310 -9190 3329 -9156
rect 3259 -9209 3329 -9190
rect 3381 -9114 3499 -9080
rect 3381 -9156 3431 -9114
rect 3652 -9132 3702 -9039
rect 3828 -9021 3978 -8951
rect 4196 -8966 4254 -8931
rect 4288 -8775 4990 -8733
rect 4288 -8809 4306 -8775
rect 4340 -8809 4938 -8775
rect 4972 -8809 4990 -8775
rect 4288 -8877 4990 -8809
rect 4288 -8911 4306 -8877
rect 4340 -8911 4938 -8877
rect 4972 -8911 4990 -8877
rect 4288 -8951 4990 -8911
rect 3828 -9055 3848 -9021
rect 3882 -9055 3978 -9021
rect 4012 -9019 4108 -8985
rect 4142 -9019 4162 -8985
rect 4012 -9089 4162 -9019
rect 3415 -9190 3431 -9156
rect 3381 -9209 3431 -9190
rect 3521 -9156 3587 -9140
rect 3521 -9190 3537 -9156
rect 3571 -9190 3587 -9156
rect 3521 -9243 3587 -9190
rect 3621 -9156 3702 -9132
rect 3621 -9190 3635 -9156
rect 3669 -9190 3702 -9156
rect 3621 -9209 3702 -9190
rect 3736 -9115 3794 -9098
rect 3736 -9149 3748 -9115
rect 3782 -9149 3794 -9115
rect 3736 -9243 3794 -9149
rect 3828 -9141 4162 -9089
rect 4288 -9019 4366 -8985
rect 4400 -9019 4465 -8985
rect 4499 -9019 4564 -8985
rect 4598 -9019 4618 -8985
rect 4288 -9089 4618 -9019
rect 4652 -9021 4990 -8951
rect 5024 -8804 5082 -8733
rect 5024 -8838 5036 -8804
rect 5070 -8838 5082 -8804
rect 5024 -8897 5082 -8838
rect 5024 -8931 5036 -8897
rect 5070 -8931 5082 -8897
rect 5024 -8966 5082 -8931
rect 5116 -8775 5450 -8733
rect 5116 -8809 5134 -8775
rect 5168 -8809 5398 -8775
rect 5432 -8809 5450 -8775
rect 5116 -8877 5450 -8809
rect 5116 -8911 5134 -8877
rect 5168 -8911 5398 -8877
rect 5432 -8911 5450 -8877
rect 5116 -8951 5450 -8911
rect 5484 -8804 5542 -8733
rect 5484 -8838 5496 -8804
rect 5530 -8838 5542 -8804
rect 5484 -8897 5542 -8838
rect 5484 -8931 5496 -8897
rect 5530 -8931 5542 -8897
rect 4652 -9055 4672 -9021
rect 4706 -9055 4775 -9021
rect 4809 -9055 4878 -9021
rect 4912 -9055 4990 -9021
rect 5116 -9021 5266 -8951
rect 5484 -8966 5542 -8931
rect 5576 -8782 5645 -8767
rect 5576 -8816 5595 -8782
rect 5629 -8816 5645 -8782
rect 5576 -8850 5645 -8816
rect 5576 -8884 5595 -8850
rect 5629 -8884 5645 -8850
rect 5576 -8934 5645 -8884
rect 5679 -8782 5745 -8733
rect 5679 -8816 5695 -8782
rect 5729 -8816 5745 -8782
rect 5679 -8850 5745 -8816
rect 5679 -8884 5695 -8850
rect 5729 -8884 5745 -8850
rect 5679 -8900 5745 -8884
rect 5835 -8782 5905 -8767
rect 5835 -8816 5853 -8782
rect 5887 -8816 5905 -8782
rect 5835 -8850 5905 -8816
rect 5835 -8884 5853 -8850
rect 5887 -8884 5905 -8850
rect 5576 -8968 5770 -8934
rect 5116 -9055 5136 -9021
rect 5170 -9055 5266 -9021
rect 5300 -9019 5396 -8985
rect 5430 -9019 5450 -8985
rect 5700 -8997 5770 -8968
rect 5835 -8996 5905 -8884
rect 5957 -8783 6007 -8767
rect 5991 -8817 6007 -8783
rect 5957 -8851 6007 -8817
rect 5991 -8885 6007 -8851
rect 5957 -8927 6007 -8885
rect 6097 -8782 6163 -8733
rect 6097 -8816 6113 -8782
rect 6147 -8816 6163 -8782
rect 6097 -8850 6163 -8816
rect 6097 -8884 6113 -8850
rect 6147 -8884 6163 -8850
rect 6097 -8893 6163 -8884
rect 6197 -8783 6278 -8767
rect 6197 -8817 6211 -8783
rect 6245 -8817 6278 -8783
rect 6197 -8851 6278 -8817
rect 6197 -8885 6211 -8851
rect 6245 -8885 6278 -8851
rect 6197 -8922 6278 -8885
rect 5957 -8961 6075 -8927
rect 6041 -8995 6075 -8961
rect 5300 -9089 5450 -9019
rect 5576 -9005 5666 -9002
rect 5576 -9045 5616 -9005
rect 5650 -9045 5666 -9005
rect 5700 -9011 5786 -8997
rect 5700 -9045 5736 -9011
rect 5770 -9045 5786 -9011
rect 5700 -9055 5786 -9045
rect 5835 -9011 6007 -8996
rect 5835 -9045 5957 -9011
rect 5991 -9045 6007 -9011
rect 5835 -9046 6007 -9045
rect 6041 -9011 6194 -8995
rect 6041 -9045 6157 -9011
rect 6191 -9045 6194 -9011
rect 5700 -9079 5770 -9055
rect 3828 -9175 3846 -9141
rect 3880 -9175 4110 -9141
rect 4144 -9175 4162 -9141
rect 3828 -9243 4162 -9175
rect 4196 -9115 4254 -9098
rect 4196 -9149 4208 -9115
rect 4242 -9149 4254 -9115
rect 4196 -9243 4254 -9149
rect 4288 -9148 4990 -9089
rect 4288 -9182 4306 -9148
rect 4340 -9182 4938 -9148
rect 4972 -9182 4990 -9148
rect 4288 -9243 4990 -9182
rect 5024 -9115 5082 -9098
rect 5024 -9149 5036 -9115
rect 5070 -9149 5082 -9115
rect 5024 -9243 5082 -9149
rect 5116 -9141 5450 -9089
rect 5116 -9175 5134 -9141
rect 5168 -9175 5398 -9141
rect 5432 -9175 5450 -9141
rect 5116 -9243 5450 -9175
rect 5484 -9115 5542 -9098
rect 5484 -9149 5496 -9115
rect 5530 -9149 5542 -9115
rect 5484 -9243 5542 -9149
rect 5576 -9113 5770 -9079
rect 5576 -9156 5642 -9113
rect 5576 -9190 5595 -9156
rect 5629 -9190 5642 -9156
rect 5576 -9209 5642 -9190
rect 5676 -9156 5742 -9147
rect 5676 -9190 5692 -9156
rect 5726 -9190 5742 -9156
rect 5676 -9243 5742 -9190
rect 5835 -9156 5905 -9046
rect 6041 -9061 6194 -9045
rect 6228 -9005 6278 -8922
rect 6312 -8804 6370 -8733
rect 6312 -8838 6324 -8804
rect 6358 -8838 6370 -8804
rect 6312 -8897 6370 -8838
rect 6312 -8931 6324 -8897
rect 6358 -8931 6370 -8897
rect 6312 -8966 6370 -8931
rect 6404 -8775 6738 -8733
rect 6404 -8809 6422 -8775
rect 6456 -8809 6686 -8775
rect 6720 -8809 6738 -8775
rect 6404 -8877 6738 -8809
rect 6404 -8911 6422 -8877
rect 6456 -8911 6686 -8877
rect 6720 -8911 6738 -8877
rect 6404 -8951 6738 -8911
rect 6772 -8804 6830 -8733
rect 6772 -8838 6784 -8804
rect 6818 -8838 6830 -8804
rect 6772 -8897 6830 -8838
rect 6772 -8931 6784 -8897
rect 6818 -8931 6830 -8897
rect 6228 -9039 6230 -9005
rect 6264 -9039 6278 -9005
rect 6041 -9080 6075 -9061
rect 5835 -9190 5852 -9156
rect 5886 -9190 5905 -9156
rect 5835 -9209 5905 -9190
rect 5957 -9114 6075 -9080
rect 5957 -9156 6007 -9114
rect 6228 -9132 6278 -9039
rect 6404 -9021 6554 -8951
rect 6772 -8966 6830 -8931
rect 6864 -8775 7566 -8733
rect 6864 -8809 6882 -8775
rect 6916 -8809 7514 -8775
rect 7548 -8809 7566 -8775
rect 6864 -8877 7566 -8809
rect 6864 -8911 6882 -8877
rect 6916 -8911 7514 -8877
rect 7548 -8911 7566 -8877
rect 6864 -8951 7566 -8911
rect 6404 -9055 6424 -9021
rect 6458 -9055 6554 -9021
rect 6588 -9019 6684 -8985
rect 6718 -9019 6738 -8985
rect 6588 -9089 6738 -9019
rect 5991 -9190 6007 -9156
rect 5957 -9209 6007 -9190
rect 6097 -9156 6163 -9140
rect 6097 -9190 6113 -9156
rect 6147 -9190 6163 -9156
rect 6097 -9243 6163 -9190
rect 6197 -9156 6278 -9132
rect 6197 -9190 6211 -9156
rect 6245 -9190 6278 -9156
rect 6197 -9209 6278 -9190
rect 6312 -9115 6370 -9098
rect 6312 -9149 6324 -9115
rect 6358 -9149 6370 -9115
rect 6312 -9243 6370 -9149
rect 6404 -9141 6738 -9089
rect 6864 -9019 6942 -8985
rect 6976 -9019 7041 -8985
rect 7075 -9019 7140 -8985
rect 7174 -9019 7194 -8985
rect 6864 -9089 7194 -9019
rect 7228 -9021 7566 -8951
rect 7600 -8804 7658 -8733
rect 7600 -8838 7612 -8804
rect 7646 -8838 7658 -8804
rect 7600 -8897 7658 -8838
rect 7600 -8931 7612 -8897
rect 7646 -8931 7658 -8897
rect 7600 -8966 7658 -8931
rect 7692 -8775 8026 -8733
rect 7692 -8809 7710 -8775
rect 7744 -8809 7974 -8775
rect 8008 -8809 8026 -8775
rect 7692 -8877 8026 -8809
rect 7692 -8911 7710 -8877
rect 7744 -8911 7974 -8877
rect 8008 -8911 8026 -8877
rect 7692 -8951 8026 -8911
rect 8060 -8804 8118 -8733
rect 8060 -8838 8072 -8804
rect 8106 -8838 8118 -8804
rect 8060 -8897 8118 -8838
rect 8060 -8931 8072 -8897
rect 8106 -8931 8118 -8897
rect 7228 -9055 7248 -9021
rect 7282 -9055 7351 -9021
rect 7385 -9055 7454 -9021
rect 7488 -9055 7566 -9021
rect 7692 -9021 7842 -8951
rect 8060 -8966 8118 -8931
rect 8152 -8782 8221 -8767
rect 8152 -8816 8171 -8782
rect 8205 -8816 8221 -8782
rect 8152 -8850 8221 -8816
rect 8152 -8884 8171 -8850
rect 8205 -8884 8221 -8850
rect 8152 -8934 8221 -8884
rect 8255 -8782 8321 -8733
rect 8255 -8816 8271 -8782
rect 8305 -8816 8321 -8782
rect 8255 -8850 8321 -8816
rect 8255 -8884 8271 -8850
rect 8305 -8884 8321 -8850
rect 8255 -8900 8321 -8884
rect 8411 -8782 8481 -8767
rect 8411 -8816 8429 -8782
rect 8463 -8816 8481 -8782
rect 8411 -8850 8481 -8816
rect 8411 -8884 8429 -8850
rect 8463 -8884 8481 -8850
rect 8152 -8968 8346 -8934
rect 7692 -9055 7712 -9021
rect 7746 -9055 7842 -9021
rect 7876 -9019 7972 -8985
rect 8006 -9019 8026 -8985
rect 8276 -8997 8346 -8968
rect 8411 -8996 8481 -8884
rect 8533 -8783 8583 -8767
rect 8567 -8817 8583 -8783
rect 8533 -8851 8583 -8817
rect 8567 -8885 8583 -8851
rect 8533 -8927 8583 -8885
rect 8673 -8782 8739 -8733
rect 8673 -8816 8689 -8782
rect 8723 -8816 8739 -8782
rect 8673 -8850 8739 -8816
rect 8673 -8884 8689 -8850
rect 8723 -8884 8739 -8850
rect 8673 -8893 8739 -8884
rect 8773 -8783 8854 -8767
rect 8773 -8817 8787 -8783
rect 8821 -8817 8854 -8783
rect 8773 -8851 8854 -8817
rect 8773 -8885 8787 -8851
rect 8821 -8885 8854 -8851
rect 8773 -8922 8854 -8885
rect 8533 -8961 8651 -8927
rect 8617 -8995 8651 -8961
rect 7876 -9089 8026 -9019
rect 8152 -9005 8242 -9002
rect 8152 -9039 8190 -9005
rect 8224 -9011 8242 -9005
rect 8152 -9045 8192 -9039
rect 8226 -9045 8242 -9011
rect 8276 -9011 8362 -8997
rect 8276 -9045 8312 -9011
rect 8346 -9045 8362 -9011
rect 8276 -9055 8362 -9045
rect 8411 -9011 8583 -8996
rect 8411 -9045 8533 -9011
rect 8567 -9045 8583 -9011
rect 8411 -9046 8583 -9045
rect 8617 -9011 8770 -8995
rect 8617 -9045 8733 -9011
rect 8767 -9045 8770 -9011
rect 8276 -9079 8346 -9055
rect 6404 -9175 6422 -9141
rect 6456 -9175 6686 -9141
rect 6720 -9175 6738 -9141
rect 6404 -9243 6738 -9175
rect 6772 -9115 6830 -9098
rect 6772 -9149 6784 -9115
rect 6818 -9149 6830 -9115
rect 6772 -9243 6830 -9149
rect 6864 -9148 7566 -9089
rect 6864 -9182 6882 -9148
rect 6916 -9182 7514 -9148
rect 7548 -9182 7566 -9148
rect 6864 -9243 7566 -9182
rect 7600 -9115 7658 -9098
rect 7600 -9149 7612 -9115
rect 7646 -9149 7658 -9115
rect 7600 -9243 7658 -9149
rect 7692 -9141 8026 -9089
rect 7692 -9175 7710 -9141
rect 7744 -9175 7974 -9141
rect 8008 -9175 8026 -9141
rect 7692 -9243 8026 -9175
rect 8060 -9115 8118 -9098
rect 8060 -9149 8072 -9115
rect 8106 -9149 8118 -9115
rect 8060 -9243 8118 -9149
rect 8152 -9113 8346 -9079
rect 8152 -9156 8218 -9113
rect 8152 -9190 8171 -9156
rect 8205 -9190 8218 -9156
rect 8152 -9209 8218 -9190
rect 8252 -9156 8318 -9147
rect 8252 -9190 8268 -9156
rect 8302 -9190 8318 -9156
rect 8252 -9243 8318 -9190
rect 8411 -9156 8481 -9046
rect 8617 -9061 8770 -9045
rect 8804 -9005 8854 -8922
rect 8888 -8804 8946 -8733
rect 8888 -8838 8900 -8804
rect 8934 -8838 8946 -8804
rect 8888 -8897 8946 -8838
rect 8888 -8931 8900 -8897
rect 8934 -8931 8946 -8897
rect 8888 -8966 8946 -8931
rect 8980 -8775 9314 -8733
rect 8980 -8809 8998 -8775
rect 9032 -8809 9262 -8775
rect 9296 -8809 9314 -8775
rect 8980 -8877 9314 -8809
rect 8980 -8911 8998 -8877
rect 9032 -8911 9262 -8877
rect 9296 -8911 9314 -8877
rect 8980 -8951 9314 -8911
rect 9348 -8804 9406 -8733
rect 9348 -8838 9360 -8804
rect 9394 -8838 9406 -8804
rect 9348 -8897 9406 -8838
rect 9348 -8931 9360 -8897
rect 9394 -8931 9406 -8897
rect 8838 -9039 8854 -9005
rect 8617 -9080 8651 -9061
rect 8411 -9190 8428 -9156
rect 8462 -9190 8481 -9156
rect 8411 -9209 8481 -9190
rect 8533 -9114 8651 -9080
rect 8533 -9156 8583 -9114
rect 8804 -9132 8854 -9039
rect 8980 -9021 9130 -8951
rect 9348 -8966 9406 -8931
rect 9440 -8775 10142 -8733
rect 9440 -8809 9458 -8775
rect 9492 -8809 10090 -8775
rect 10124 -8809 10142 -8775
rect 9440 -8877 10142 -8809
rect 9440 -8911 9458 -8877
rect 9492 -8911 10090 -8877
rect 10124 -8911 10142 -8877
rect 9440 -8951 10142 -8911
rect 8980 -9055 9000 -9021
rect 9034 -9055 9130 -9021
rect 9164 -9019 9260 -8985
rect 9294 -9019 9314 -8985
rect 9164 -9089 9314 -9019
rect 8567 -9190 8583 -9156
rect 8533 -9209 8583 -9190
rect 8673 -9156 8739 -9140
rect 8673 -9190 8689 -9156
rect 8723 -9190 8739 -9156
rect 8673 -9243 8739 -9190
rect 8773 -9156 8854 -9132
rect 8773 -9190 8787 -9156
rect 8821 -9190 8854 -9156
rect 8773 -9209 8854 -9190
rect 8888 -9115 8946 -9098
rect 8888 -9149 8900 -9115
rect 8934 -9149 8946 -9115
rect 8888 -9243 8946 -9149
rect 8980 -9141 9314 -9089
rect 9440 -9019 9518 -8985
rect 9552 -9019 9617 -8985
rect 9651 -9019 9716 -8985
rect 9750 -9019 9770 -8985
rect 9440 -9089 9770 -9019
rect 9804 -9021 10142 -8951
rect 10176 -8804 10234 -8733
rect 10176 -8838 10188 -8804
rect 10222 -8838 10234 -8804
rect 10176 -8897 10234 -8838
rect 10176 -8931 10188 -8897
rect 10222 -8931 10234 -8897
rect 10176 -8966 10234 -8931
rect 10360 -8775 10694 -8733
rect 10360 -8809 10378 -8775
rect 10412 -8809 10642 -8775
rect 10676 -8809 10694 -8775
rect 10360 -8877 10694 -8809
rect 10360 -8911 10378 -8877
rect 10412 -8911 10642 -8877
rect 10676 -8911 10694 -8877
rect 10360 -8951 10694 -8911
rect 10728 -8782 10797 -8767
rect 10728 -8816 10747 -8782
rect 10781 -8816 10797 -8782
rect 10728 -8850 10797 -8816
rect 10728 -8884 10747 -8850
rect 10781 -8884 10797 -8850
rect 10728 -8934 10797 -8884
rect 10831 -8782 10897 -8733
rect 10831 -8816 10847 -8782
rect 10881 -8816 10897 -8782
rect 10831 -8850 10897 -8816
rect 10831 -8884 10847 -8850
rect 10881 -8884 10897 -8850
rect 10831 -8900 10897 -8884
rect 10987 -8782 11057 -8767
rect 10987 -8816 11005 -8782
rect 11039 -8816 11057 -8782
rect 10987 -8850 11057 -8816
rect 10987 -8884 11005 -8850
rect 11039 -8884 11057 -8850
rect 9804 -9055 9824 -9021
rect 9858 -9055 9927 -9021
rect 9961 -9055 10030 -9021
rect 10064 -9055 10142 -9021
rect 10360 -9021 10510 -8951
rect 10728 -8968 10922 -8934
rect 10360 -9055 10380 -9021
rect 10414 -9055 10510 -9021
rect 10544 -9019 10640 -8985
rect 10674 -9019 10694 -8985
rect 10852 -8997 10922 -8968
rect 10987 -8996 11057 -8884
rect 11109 -8783 11159 -8767
rect 11143 -8817 11159 -8783
rect 11109 -8851 11159 -8817
rect 11143 -8885 11159 -8851
rect 11109 -8927 11159 -8885
rect 11249 -8782 11315 -8733
rect 11249 -8816 11265 -8782
rect 11299 -8816 11315 -8782
rect 11249 -8850 11315 -8816
rect 11249 -8884 11265 -8850
rect 11299 -8884 11315 -8850
rect 11249 -8893 11315 -8884
rect 11349 -8783 11430 -8767
rect 11349 -8817 11363 -8783
rect 11397 -8817 11430 -8783
rect 11349 -8851 11430 -8817
rect 11349 -8885 11363 -8851
rect 11397 -8885 11430 -8851
rect 11349 -8922 11430 -8885
rect 11109 -8961 11227 -8927
rect 11193 -8995 11227 -8961
rect 11380 -8971 11430 -8922
rect 11464 -8804 11522 -8733
rect 11464 -8838 11476 -8804
rect 11510 -8838 11522 -8804
rect 11464 -8897 11522 -8838
rect 11464 -8931 11476 -8897
rect 11510 -8931 11522 -8897
rect 11464 -8966 11522 -8931
rect 11648 -8775 11982 -8733
rect 11648 -8809 11666 -8775
rect 11700 -8809 11930 -8775
rect 11964 -8809 11982 -8775
rect 11648 -8877 11982 -8809
rect 11648 -8911 11666 -8877
rect 11700 -8911 11930 -8877
rect 11964 -8911 11982 -8877
rect 11648 -8951 11982 -8911
rect 12384 -8804 12442 -8733
rect 12384 -8838 12396 -8804
rect 12430 -8838 12442 -8804
rect 12384 -8897 12442 -8838
rect 12384 -8931 12396 -8897
rect 12430 -8931 12442 -8897
rect 12476 -8782 12545 -8733
rect 12476 -8816 12502 -8782
rect 12536 -8816 12545 -8782
rect 12476 -8850 12545 -8816
rect 12476 -8884 12502 -8850
rect 12536 -8884 12545 -8850
rect 12476 -8900 12545 -8884
rect 12580 -8789 12631 -8773
rect 12580 -8823 12588 -8789
rect 12622 -8823 12631 -8789
rect 12580 -8877 12631 -8823
rect 10544 -9089 10694 -9019
rect 10728 -9005 10818 -9002
rect 10728 -9039 10764 -9005
rect 10798 -9011 10818 -9005
rect 10728 -9045 10768 -9039
rect 10802 -9045 10818 -9011
rect 10852 -9011 10938 -8997
rect 10852 -9045 10888 -9011
rect 10922 -9045 10938 -9011
rect 10852 -9055 10938 -9045
rect 10987 -9011 11159 -8996
rect 10987 -9045 11109 -9011
rect 11143 -9045 11159 -9011
rect 10987 -9046 11159 -9045
rect 11193 -9011 11346 -8995
rect 11193 -9045 11309 -9011
rect 11343 -9045 11346 -9011
rect 10852 -9079 10922 -9055
rect 8980 -9175 8998 -9141
rect 9032 -9175 9262 -9141
rect 9296 -9175 9314 -9141
rect 8980 -9243 9314 -9175
rect 9348 -9115 9406 -9098
rect 9348 -9149 9360 -9115
rect 9394 -9149 9406 -9115
rect 9348 -9243 9406 -9149
rect 9440 -9148 10142 -9089
rect 9440 -9182 9458 -9148
rect 9492 -9182 10090 -9148
rect 10124 -9182 10142 -9148
rect 9440 -9243 10142 -9182
rect 10176 -9115 10234 -9098
rect 10176 -9149 10188 -9115
rect 10222 -9149 10234 -9115
rect 10176 -9243 10234 -9149
rect 10360 -9141 10694 -9089
rect 10360 -9175 10378 -9141
rect 10412 -9175 10642 -9141
rect 10676 -9175 10694 -9141
rect 10360 -9243 10694 -9175
rect 10728 -9113 10922 -9079
rect 10728 -9156 10794 -9113
rect 10728 -9190 10747 -9156
rect 10781 -9190 10794 -9156
rect 10728 -9209 10794 -9190
rect 10828 -9156 10894 -9147
rect 10828 -9190 10844 -9156
rect 10878 -9190 10894 -9156
rect 10828 -9243 10894 -9190
rect 10987 -9156 11057 -9046
rect 11193 -9061 11346 -9045
rect 11380 -9005 11387 -8971
rect 11421 -9005 11430 -8971
rect 11193 -9080 11227 -9061
rect 10987 -9190 11004 -9156
rect 11038 -9190 11057 -9156
rect 10987 -9209 11057 -9190
rect 11109 -9114 11227 -9080
rect 11109 -9156 11159 -9114
rect 11380 -9132 11430 -9005
rect 11648 -9021 11798 -8951
rect 12384 -8966 12442 -8931
rect 12580 -8911 12588 -8877
rect 12622 -8911 12631 -8877
rect 12665 -8782 12717 -8733
rect 12665 -8816 12674 -8782
rect 12708 -8816 12717 -8782
rect 12665 -8850 12717 -8816
rect 12665 -8884 12674 -8850
rect 12708 -8884 12717 -8850
rect 12665 -8900 12717 -8884
rect 12752 -8789 12803 -8773
rect 12752 -8823 12760 -8789
rect 12794 -8823 12803 -8789
rect 12752 -8877 12803 -8823
rect 12580 -8934 12631 -8911
rect 12752 -8911 12760 -8877
rect 12794 -8911 12803 -8877
rect 12837 -8782 12889 -8733
rect 12837 -8816 12846 -8782
rect 12880 -8816 12889 -8782
rect 12837 -8850 12889 -8816
rect 12837 -8884 12846 -8850
rect 12880 -8884 12889 -8850
rect 12837 -8900 12889 -8884
rect 12923 -8789 12975 -8773
rect 12923 -8823 12932 -8789
rect 12966 -8823 12975 -8789
rect 12923 -8877 12975 -8823
rect 12752 -8934 12803 -8911
rect 12923 -8911 12932 -8877
rect 12966 -8911 12975 -8877
rect 13009 -8782 13086 -8733
rect 13009 -8816 13018 -8782
rect 13052 -8816 13086 -8782
rect 13009 -8850 13086 -8816
rect 13009 -8884 13018 -8850
rect 13052 -8884 13086 -8850
rect 13009 -8900 13086 -8884
rect 13120 -8804 13178 -8733
rect 13120 -8838 13132 -8804
rect 13166 -8838 13178 -8804
rect 13120 -8897 13178 -8838
rect 12923 -8934 12975 -8911
rect 13120 -8931 13132 -8897
rect 13166 -8931 13178 -8897
rect 12480 -8968 13086 -8934
rect 13120 -8966 13178 -8931
rect 13212 -8775 13546 -8733
rect 13212 -8809 13230 -8775
rect 13264 -8809 13494 -8775
rect 13528 -8809 13546 -8775
rect 13212 -8877 13546 -8809
rect 13212 -8911 13230 -8877
rect 13264 -8911 13494 -8877
rect 13528 -8911 13546 -8877
rect 13212 -8951 13546 -8911
rect 11648 -9055 11668 -9021
rect 11702 -9055 11798 -9021
rect 11832 -9019 11928 -8985
rect 11962 -9019 11982 -8985
rect 11832 -9089 11982 -9019
rect 11143 -9190 11159 -9156
rect 11109 -9209 11159 -9190
rect 11249 -9156 11315 -9140
rect 11249 -9190 11265 -9156
rect 11299 -9190 11315 -9156
rect 11249 -9243 11315 -9190
rect 11349 -9156 11430 -9132
rect 11349 -9190 11363 -9156
rect 11397 -9190 11430 -9156
rect 11349 -9209 11430 -9190
rect 11464 -9115 11522 -9098
rect 11464 -9149 11476 -9115
rect 11510 -9149 11522 -9115
rect 11464 -9243 11522 -9149
rect 11648 -9141 11982 -9089
rect 12480 -9081 12514 -8968
rect 13026 -9001 13086 -8968
rect 12548 -9008 12991 -9002
rect 12548 -9042 12558 -9008
rect 12592 -9011 12642 -9008
rect 12676 -9011 12739 -9008
rect 12773 -9011 12836 -9008
rect 12870 -9011 12942 -9008
rect 12548 -9045 12574 -9042
rect 12608 -9045 12642 -9011
rect 12676 -9045 12710 -9011
rect 12773 -9042 12778 -9011
rect 12744 -9045 12778 -9042
rect 12812 -9042 12836 -9011
rect 12812 -9045 12846 -9042
rect 12880 -9045 12914 -9011
rect 12976 -9042 12991 -9008
rect 12948 -9045 12991 -9042
rect 12548 -9047 12991 -9045
rect 13026 -9035 13038 -9001
rect 13072 -9035 13086 -9001
rect 13026 -9073 13086 -9035
rect 13026 -9081 13038 -9073
rect 11648 -9175 11666 -9141
rect 11700 -9175 11930 -9141
rect 11964 -9175 11982 -9141
rect 11648 -9243 11982 -9175
rect 12384 -9115 12442 -9098
rect 12480 -9107 13038 -9081
rect 13072 -9107 13086 -9073
rect 13212 -9019 13232 -8985
rect 13266 -9019 13362 -8985
rect 13212 -9089 13362 -9019
rect 13396 -9021 13546 -8951
rect 13580 -8804 13638 -8733
rect 13580 -8838 13592 -8804
rect 13626 -8838 13638 -8804
rect 13580 -8897 13638 -8838
rect 13674 -8775 13733 -8733
rect 13674 -8809 13690 -8775
rect 13724 -8809 13733 -8775
rect 13674 -8843 13733 -8809
rect 13674 -8877 13690 -8843
rect 13724 -8877 13733 -8843
rect 13674 -8895 13733 -8877
rect 13769 -8783 13818 -8767
rect 13769 -8817 13776 -8783
rect 13810 -8817 13818 -8783
rect 13769 -8851 13818 -8817
rect 13769 -8885 13776 -8851
rect 13810 -8885 13818 -8851
rect 13580 -8931 13592 -8897
rect 13626 -8931 13638 -8897
rect 13580 -8966 13638 -8931
rect 13769 -8995 13818 -8885
rect 13853 -8775 13905 -8733
rect 14025 -8734 15280 -8733
rect 13853 -8809 13862 -8775
rect 13896 -8809 13905 -8775
rect 13853 -8843 13905 -8809
rect 13853 -8877 13862 -8843
rect 13896 -8877 13905 -8843
rect 13853 -8895 13905 -8877
rect 13941 -8791 13991 -8768
rect 13941 -8825 13948 -8791
rect 13982 -8825 13991 -8791
rect 13941 -8859 13991 -8825
rect 13941 -8893 13948 -8859
rect 13982 -8893 13991 -8859
rect 14025 -8775 14077 -8734
rect 14025 -8809 14034 -8775
rect 14068 -8809 14077 -8775
rect 14025 -8843 14077 -8809
rect 14025 -8877 14034 -8843
rect 14068 -8877 14077 -8843
rect 14025 -8893 14077 -8877
rect 14111 -8819 14163 -8768
rect 14111 -8853 14120 -8819
rect 14154 -8853 14163 -8819
rect 13941 -8995 13991 -8893
rect 14111 -8905 14163 -8853
rect 14197 -8799 14249 -8734
rect 14197 -8833 14206 -8799
rect 14240 -8833 14249 -8799
rect 14197 -8879 14249 -8833
rect 14283 -8819 14335 -8768
rect 14283 -8853 14292 -8819
rect 14326 -8853 14335 -8819
rect 14111 -8939 14120 -8905
rect 14154 -8913 14163 -8905
rect 14283 -8905 14335 -8853
rect 14369 -8799 14421 -8734
rect 14369 -8833 14378 -8799
rect 14412 -8833 14421 -8799
rect 14369 -8879 14421 -8833
rect 14455 -8819 14507 -8768
rect 14455 -8853 14464 -8819
rect 14498 -8853 14507 -8819
rect 14283 -8913 14292 -8905
rect 14154 -8939 14292 -8913
rect 14326 -8913 14335 -8905
rect 14455 -8905 14507 -8853
rect 14541 -8799 14593 -8734
rect 14541 -8833 14550 -8799
rect 14584 -8833 14593 -8799
rect 14541 -8879 14593 -8833
rect 14627 -8819 14679 -8768
rect 14627 -8853 14636 -8819
rect 14670 -8853 14679 -8819
rect 14455 -8913 14464 -8905
rect 14326 -8939 14464 -8913
rect 14498 -8913 14507 -8905
rect 14627 -8905 14679 -8853
rect 14713 -8799 14762 -8734
rect 14713 -8833 14722 -8799
rect 14756 -8833 14762 -8799
rect 14713 -8879 14762 -8833
rect 14796 -8819 14848 -8768
rect 14796 -8853 14807 -8819
rect 14841 -8853 14848 -8819
rect 14627 -8913 14636 -8905
rect 14498 -8939 14636 -8913
rect 14670 -8913 14679 -8905
rect 14796 -8905 14848 -8853
rect 14885 -8799 14934 -8734
rect 14885 -8833 14893 -8799
rect 14927 -8833 14934 -8799
rect 14885 -8879 14934 -8833
rect 14968 -8819 15020 -8768
rect 14968 -8853 14979 -8819
rect 15013 -8853 15020 -8819
rect 14796 -8913 14807 -8905
rect 14670 -8939 14807 -8913
rect 14841 -8913 14848 -8905
rect 14968 -8905 15020 -8853
rect 15057 -8799 15106 -8734
rect 15057 -8833 15065 -8799
rect 15099 -8833 15106 -8799
rect 15057 -8879 15106 -8833
rect 15140 -8819 15192 -8768
rect 15140 -8853 15151 -8819
rect 15185 -8853 15192 -8819
rect 14968 -8913 14979 -8905
rect 14841 -8939 14979 -8913
rect 15013 -8913 15020 -8905
rect 15140 -8905 15192 -8853
rect 15229 -8799 15280 -8734
rect 15229 -8833 15237 -8799
rect 15271 -8833 15280 -8799
rect 15229 -8879 15280 -8833
rect 15314 -8819 15372 -8768
rect 15314 -8853 15323 -8819
rect 15357 -8853 15372 -8819
rect 15140 -8913 15151 -8905
rect 15013 -8939 15151 -8913
rect 15185 -8916 15192 -8905
rect 15314 -8905 15372 -8853
rect 15406 -8799 15460 -8733
rect 15406 -8833 15409 -8799
rect 15443 -8833 15460 -8799
rect 15406 -8882 15460 -8833
rect 15512 -8804 15570 -8733
rect 15512 -8838 15524 -8804
rect 15558 -8838 15570 -8804
rect 15314 -8916 15323 -8905
rect 15185 -8939 15323 -8916
rect 15357 -8916 15372 -8905
rect 15512 -8897 15570 -8838
rect 15357 -8939 15460 -8916
rect 14111 -8954 15460 -8939
rect 14111 -8961 15248 -8954
rect 15227 -8988 15248 -8961
rect 15282 -8955 15460 -8954
rect 15282 -8988 15340 -8955
rect 15227 -8989 15340 -8988
rect 15374 -8989 15460 -8955
rect 15512 -8931 15524 -8897
rect 15558 -8931 15570 -8897
rect 15512 -8966 15570 -8931
rect 15604 -8775 16673 -8733
rect 15604 -8809 15622 -8775
rect 15656 -8809 16622 -8775
rect 16656 -8809 16673 -8775
rect 15604 -8877 16673 -8809
rect 15604 -8911 15622 -8877
rect 15656 -8911 16622 -8877
rect 16656 -8911 16673 -8877
rect 15604 -8951 16673 -8911
rect 13396 -9055 13492 -9021
rect 13526 -9055 13546 -9021
rect 13672 -9011 13735 -8995
rect 13672 -9038 13692 -9011
rect 13672 -9072 13684 -9038
rect 13726 -9045 13735 -9011
rect 13718 -9072 13735 -9045
rect 12480 -9115 13086 -9107
rect 13120 -9115 13178 -9098
rect 12384 -9149 12396 -9115
rect 12430 -9149 12442 -9115
rect 12384 -9243 12442 -9149
rect 12572 -9165 12631 -9149
rect 12572 -9199 12588 -9165
rect 12622 -9199 12631 -9165
rect 12572 -9243 12631 -9199
rect 12665 -9154 12717 -9115
rect 12665 -9188 12674 -9154
rect 12708 -9188 12717 -9154
rect 12665 -9204 12717 -9188
rect 12751 -9165 12803 -9149
rect 12751 -9199 12760 -9165
rect 12794 -9199 12803 -9165
rect 12751 -9243 12803 -9199
rect 12837 -9154 12888 -9115
rect 13120 -9149 13132 -9115
rect 13166 -9149 13178 -9115
rect 12837 -9188 12846 -9154
rect 12880 -9188 12888 -9154
rect 12837 -9204 12888 -9188
rect 12922 -9165 12982 -9149
rect 12922 -9199 12932 -9165
rect 12966 -9199 12982 -9165
rect 12922 -9243 12982 -9199
rect 13120 -9243 13178 -9149
rect 13212 -9141 13546 -9089
rect 13212 -9175 13230 -9141
rect 13264 -9175 13494 -9141
rect 13528 -9175 13546 -9141
rect 13212 -9243 13546 -9175
rect 13580 -9115 13638 -9098
rect 13672 -9107 13735 -9072
rect 13769 -9011 15193 -8995
rect 13769 -9045 14119 -9011
rect 14153 -9045 14187 -9011
rect 14221 -9045 14255 -9011
rect 14289 -9045 14323 -9011
rect 14357 -9045 14391 -9011
rect 14425 -9045 14459 -9011
rect 14493 -9045 14527 -9011
rect 14561 -9045 14595 -9011
rect 14629 -9045 14663 -9011
rect 14697 -9045 14731 -9011
rect 14765 -9045 14799 -9011
rect 14833 -9045 14867 -9011
rect 14901 -9045 14935 -9011
rect 14969 -9045 15003 -9011
rect 15037 -9045 15071 -9011
rect 15105 -9045 15139 -9011
rect 15173 -9045 15193 -9011
rect 13580 -9149 13592 -9115
rect 13626 -9149 13638 -9115
rect 13580 -9243 13638 -9149
rect 13672 -9167 13733 -9141
rect 13672 -9201 13690 -9167
rect 13724 -9201 13733 -9167
rect 13672 -9243 13733 -9201
rect 13769 -9154 13819 -9045
rect 13769 -9188 13776 -9154
rect 13810 -9188 13819 -9154
rect 13769 -9207 13819 -9188
rect 13853 -9154 13905 -9138
rect 13853 -9188 13862 -9154
rect 13896 -9188 13905 -9154
rect 13853 -9243 13905 -9188
rect 13941 -9154 13991 -9045
rect 15227 -9050 15460 -8989
rect 15227 -9079 15248 -9050
rect 14111 -9084 15248 -9079
rect 15282 -9084 15341 -9050
rect 15375 -9084 15460 -9050
rect 14111 -9113 15460 -9084
rect 15604 -9019 15682 -8985
rect 15716 -9019 15810 -8985
rect 15844 -9019 15938 -8985
rect 15972 -9019 16066 -8985
rect 16100 -9019 16120 -8985
rect 15604 -9089 16120 -9019
rect 16154 -9021 16673 -8951
rect 16154 -9055 16174 -9021
rect 16208 -9055 16302 -9021
rect 16336 -9055 16430 -9021
rect 16464 -9055 16558 -9021
rect 16592 -9055 16673 -9021
rect 13941 -9188 13948 -9154
rect 13982 -9188 13991 -9154
rect 13941 -9207 13991 -9188
rect 14025 -9154 14077 -9131
rect 14025 -9188 14034 -9154
rect 14068 -9188 14077 -9154
rect 14025 -9243 14077 -9188
rect 14111 -9154 14163 -9113
rect 14111 -9188 14120 -9154
rect 14154 -9188 14163 -9154
rect 14111 -9204 14163 -9188
rect 14197 -9163 14249 -9147
rect 14197 -9197 14206 -9163
rect 14240 -9197 14249 -9163
rect 14197 -9243 14249 -9197
rect 14283 -9154 14335 -9113
rect 14283 -9188 14292 -9154
rect 14326 -9188 14335 -9154
rect 14283 -9204 14335 -9188
rect 14369 -9163 14421 -9147
rect 14369 -9197 14378 -9163
rect 14412 -9197 14421 -9163
rect 14369 -9243 14421 -9197
rect 14455 -9154 14507 -9113
rect 14455 -9188 14464 -9154
rect 14498 -9188 14507 -9154
rect 14455 -9204 14507 -9188
rect 14541 -9163 14590 -9147
rect 14541 -9197 14550 -9163
rect 14584 -9197 14590 -9163
rect 14541 -9243 14590 -9197
rect 14624 -9154 14679 -9113
rect 14624 -9188 14636 -9154
rect 14670 -9188 14679 -9154
rect 14624 -9204 14679 -9188
rect 14713 -9163 14762 -9147
rect 14713 -9197 14722 -9163
rect 14756 -9197 14762 -9163
rect 14713 -9243 14762 -9197
rect 14796 -9154 14848 -9113
rect 14796 -9188 14807 -9154
rect 14841 -9188 14848 -9154
rect 14796 -9204 14848 -9188
rect 14884 -9163 14934 -9147
rect 14884 -9197 14893 -9163
rect 14927 -9197 14934 -9163
rect 14884 -9243 14934 -9197
rect 14968 -9154 15020 -9113
rect 14968 -9188 14979 -9154
rect 15013 -9188 15020 -9154
rect 14968 -9204 15020 -9188
rect 15056 -9163 15106 -9147
rect 15056 -9197 15065 -9163
rect 15099 -9197 15106 -9163
rect 15056 -9243 15106 -9197
rect 15140 -9154 15192 -9113
rect 15140 -9188 15151 -9154
rect 15185 -9188 15192 -9154
rect 15140 -9204 15192 -9188
rect 15228 -9163 15280 -9147
rect 15228 -9197 15237 -9163
rect 15271 -9197 15280 -9163
rect 15228 -9243 15280 -9197
rect 15314 -9154 15366 -9113
rect 15512 -9115 15570 -9098
rect 15314 -9188 15323 -9154
rect 15357 -9188 15366 -9154
rect 15314 -9204 15366 -9188
rect 15400 -9163 15460 -9147
rect 15400 -9197 15409 -9163
rect 15443 -9197 15460 -9163
rect 15400 -9243 15460 -9197
rect 15512 -9149 15524 -9115
rect 15558 -9149 15570 -9115
rect 15512 -9243 15570 -9149
rect 15604 -9148 16673 -9089
rect 15604 -9182 15622 -9148
rect 15656 -9182 16622 -9148
rect 16656 -9182 16673 -9148
rect 15604 -9243 16673 -9182
rect -2997 -9277 -2968 -9243
rect -2934 -9277 -2876 -9243
rect -2842 -9277 -2784 -9243
rect -2750 -9277 -2692 -9243
rect -2658 -9277 -2600 -9243
rect -2566 -9277 -2508 -9243
rect -2474 -9277 -2416 -9243
rect -2382 -9277 -2324 -9243
rect -2290 -9277 -2232 -9243
rect -2198 -9277 -2140 -9243
rect -2106 -9277 -2048 -9243
rect -2014 -9277 -1956 -9243
rect -1922 -9277 -1864 -9243
rect -1830 -9277 -1772 -9243
rect -1738 -9277 -1680 -9243
rect -1646 -9277 -1588 -9243
rect -1554 -9277 -1496 -9243
rect -1462 -9277 -1404 -9243
rect -1370 -9277 -1312 -9243
rect -1278 -9277 -1220 -9243
rect -1186 -9277 -1128 -9243
rect -1094 -9277 -1036 -9243
rect -1002 -9277 -944 -9243
rect -910 -9277 -852 -9243
rect -818 -9277 -760 -9243
rect -726 -9277 -668 -9243
rect -634 -9277 -576 -9243
rect -542 -9277 -484 -9243
rect -450 -9277 -392 -9243
rect -358 -9277 -300 -9243
rect -266 -9277 -208 -9243
rect -174 -9277 -116 -9243
rect -82 -9277 -24 -9243
rect 10 -9277 68 -9243
rect 102 -9277 160 -9243
rect 194 -9277 252 -9243
rect 286 -9277 344 -9243
rect 378 -9277 436 -9243
rect 470 -9277 528 -9243
rect 562 -9277 620 -9243
rect 654 -9277 712 -9243
rect 746 -9277 804 -9243
rect 838 -9277 896 -9243
rect 930 -9277 988 -9243
rect 1022 -9277 1080 -9243
rect 1114 -9277 1172 -9243
rect 1206 -9277 1264 -9243
rect 1298 -9277 1356 -9243
rect 1390 -9277 1448 -9243
rect 1482 -9277 1540 -9243
rect 1574 -9277 1632 -9243
rect 1666 -9277 1724 -9243
rect 1758 -9277 1816 -9243
rect 1850 -9277 1908 -9243
rect 1942 -9277 2000 -9243
rect 2034 -9277 2092 -9243
rect 2126 -9277 2184 -9243
rect 2218 -9277 2276 -9243
rect 2310 -9277 2368 -9243
rect 2402 -9277 2460 -9243
rect 2494 -9277 2552 -9243
rect 2586 -9277 2644 -9243
rect 2678 -9277 2736 -9243
rect 2770 -9277 2828 -9243
rect 2862 -9277 2920 -9243
rect 2954 -9277 3012 -9243
rect 3046 -9277 3104 -9243
rect 3138 -9277 3196 -9243
rect 3230 -9277 3288 -9243
rect 3322 -9277 3380 -9243
rect 3414 -9277 3472 -9243
rect 3506 -9277 3564 -9243
rect 3598 -9277 3656 -9243
rect 3690 -9277 3748 -9243
rect 3782 -9277 3840 -9243
rect 3874 -9277 3932 -9243
rect 3966 -9277 4024 -9243
rect 4058 -9277 4116 -9243
rect 4150 -9277 4208 -9243
rect 4242 -9277 4300 -9243
rect 4334 -9277 4392 -9243
rect 4426 -9277 4484 -9243
rect 4518 -9277 4576 -9243
rect 4610 -9277 4668 -9243
rect 4702 -9277 4760 -9243
rect 4794 -9277 4852 -9243
rect 4886 -9277 4944 -9243
rect 4978 -9277 5036 -9243
rect 5070 -9277 5128 -9243
rect 5162 -9277 5220 -9243
rect 5254 -9277 5312 -9243
rect 5346 -9277 5404 -9243
rect 5438 -9277 5496 -9243
rect 5530 -9277 5588 -9243
rect 5622 -9277 5680 -9243
rect 5714 -9277 5772 -9243
rect 5806 -9277 5864 -9243
rect 5898 -9277 5956 -9243
rect 5990 -9277 6048 -9243
rect 6082 -9277 6140 -9243
rect 6174 -9277 6232 -9243
rect 6266 -9277 6324 -9243
rect 6358 -9277 6416 -9243
rect 6450 -9277 6508 -9243
rect 6542 -9277 6600 -9243
rect 6634 -9277 6692 -9243
rect 6726 -9277 6784 -9243
rect 6818 -9277 6876 -9243
rect 6910 -9277 6968 -9243
rect 7002 -9277 7060 -9243
rect 7094 -9277 7152 -9243
rect 7186 -9277 7244 -9243
rect 7278 -9277 7336 -9243
rect 7370 -9277 7428 -9243
rect 7462 -9277 7520 -9243
rect 7554 -9277 7612 -9243
rect 7646 -9277 7704 -9243
rect 7738 -9277 7796 -9243
rect 7830 -9277 7888 -9243
rect 7922 -9277 7980 -9243
rect 8014 -9277 8072 -9243
rect 8106 -9277 8164 -9243
rect 8198 -9277 8256 -9243
rect 8290 -9277 8348 -9243
rect 8382 -9277 8440 -9243
rect 8474 -9277 8532 -9243
rect 8566 -9277 8624 -9243
rect 8658 -9277 8716 -9243
rect 8750 -9277 8808 -9243
rect 8842 -9277 8900 -9243
rect 8934 -9277 8992 -9243
rect 9026 -9277 9084 -9243
rect 9118 -9277 9176 -9243
rect 9210 -9277 9268 -9243
rect 9302 -9277 9360 -9243
rect 9394 -9277 9452 -9243
rect 9486 -9277 9544 -9243
rect 9578 -9277 9636 -9243
rect 9670 -9277 9728 -9243
rect 9762 -9277 9820 -9243
rect 9854 -9277 9912 -9243
rect 9946 -9277 10004 -9243
rect 10038 -9277 10096 -9243
rect 10130 -9277 10188 -9243
rect 10222 -9277 10280 -9243
rect 10314 -9277 10372 -9243
rect 10406 -9277 10464 -9243
rect 10498 -9277 10556 -9243
rect 10590 -9277 10648 -9243
rect 10682 -9277 10740 -9243
rect 10774 -9277 10832 -9243
rect 10866 -9277 10924 -9243
rect 10958 -9277 11016 -9243
rect 11050 -9277 11108 -9243
rect 11142 -9277 11200 -9243
rect 11234 -9277 11292 -9243
rect 11326 -9277 11384 -9243
rect 11418 -9277 11476 -9243
rect 11510 -9277 11568 -9243
rect 11602 -9277 11660 -9243
rect 11694 -9277 11752 -9243
rect 11786 -9277 11844 -9243
rect 11878 -9277 11936 -9243
rect 11970 -9277 12028 -9243
rect 12062 -9277 12120 -9243
rect 12154 -9277 12212 -9243
rect 12246 -9277 12304 -9243
rect 12338 -9277 12396 -9243
rect 12430 -9277 12488 -9243
rect 12522 -9277 12580 -9243
rect 12614 -9277 12672 -9243
rect 12706 -9277 12764 -9243
rect 12798 -9277 12856 -9243
rect 12890 -9277 12948 -9243
rect 12982 -9277 13040 -9243
rect 13074 -9277 13132 -9243
rect 13166 -9277 13224 -9243
rect 13258 -9277 13316 -9243
rect 13350 -9277 13408 -9243
rect 13442 -9277 13500 -9243
rect 13534 -9277 13592 -9243
rect 13626 -9277 13684 -9243
rect 13718 -9277 13776 -9243
rect 13810 -9277 13868 -9243
rect 13902 -9277 13960 -9243
rect 13994 -9277 14052 -9243
rect 14086 -9277 14144 -9243
rect 14178 -9277 14236 -9243
rect 14270 -9277 14328 -9243
rect 14362 -9277 14420 -9243
rect 14454 -9277 14512 -9243
rect 14546 -9277 14604 -9243
rect 14638 -9277 14696 -9243
rect 14730 -9277 14788 -9243
rect 14822 -9277 14880 -9243
rect 14914 -9277 14972 -9243
rect 15006 -9277 15064 -9243
rect 15098 -9277 15156 -9243
rect 15190 -9277 15248 -9243
rect 15282 -9277 15340 -9243
rect 15374 -9277 15432 -9243
rect 15466 -9277 15524 -9243
rect 15558 -9277 15616 -9243
rect 15650 -9277 15708 -9243
rect 15742 -9277 15800 -9243
rect 15834 -9277 15892 -9243
rect 15926 -9277 15984 -9243
rect 16018 -9277 16076 -9243
rect 16110 -9277 16168 -9243
rect 16202 -9277 16260 -9243
rect 16294 -9277 16352 -9243
rect 16386 -9277 16444 -9243
rect 16478 -9277 16536 -9243
rect 16570 -9277 16628 -9243
rect 16662 -9277 16691 -9243
rect -2980 -9338 -2278 -9277
rect -2980 -9372 -2962 -9338
rect -2928 -9372 -2330 -9338
rect -2296 -9372 -2278 -9338
rect -2980 -9431 -2278 -9372
rect -2244 -9371 -2186 -9277
rect -2244 -9405 -2232 -9371
rect -2198 -9405 -2186 -9371
rect -2244 -9422 -2186 -9405
rect -1600 -9338 -898 -9277
rect -1600 -9372 -1582 -9338
rect -1548 -9372 -950 -9338
rect -916 -9372 -898 -9338
rect -1600 -9431 -898 -9372
rect -2980 -9499 -2902 -9465
rect -2868 -9499 -2799 -9465
rect -2765 -9499 -2696 -9465
rect -2662 -9499 -2642 -9465
rect -2980 -9569 -2642 -9499
rect -2608 -9501 -2278 -9431
rect -2608 -9535 -2588 -9501
rect -2554 -9535 -2489 -9501
rect -2455 -9535 -2390 -9501
rect -2356 -9535 -2278 -9501
rect -1600 -9499 -1522 -9465
rect -1488 -9499 -1419 -9465
rect -1385 -9499 -1316 -9465
rect -1282 -9499 -1262 -9465
rect -2980 -9609 -2278 -9569
rect -2980 -9643 -2962 -9609
rect -2928 -9643 -2330 -9609
rect -2296 -9643 -2278 -9609
rect -2980 -9711 -2278 -9643
rect -2980 -9745 -2962 -9711
rect -2928 -9745 -2330 -9711
rect -2296 -9745 -2278 -9711
rect -2980 -9787 -2278 -9745
rect -2244 -9589 -2186 -9554
rect -2244 -9623 -2232 -9589
rect -2198 -9623 -2186 -9589
rect -2244 -9682 -2186 -9623
rect -2244 -9716 -2232 -9682
rect -2198 -9716 -2186 -9682
rect -2244 -9787 -2186 -9716
rect -1600 -9569 -1262 -9499
rect -1228 -9501 -898 -9431
rect -1228 -9535 -1208 -9501
rect -1174 -9535 -1109 -9501
rect -1075 -9535 -1010 -9501
rect -976 -9535 -898 -9501
rect -864 -9330 -783 -9311
rect -864 -9364 -831 -9330
rect -797 -9364 -783 -9330
rect -864 -9388 -783 -9364
rect -749 -9330 -683 -9277
rect -749 -9364 -733 -9330
rect -699 -9364 -683 -9330
rect -749 -9380 -683 -9364
rect -593 -9330 -543 -9311
rect -593 -9364 -577 -9330
rect -864 -9516 -814 -9388
rect -593 -9406 -543 -9364
rect -661 -9440 -543 -9406
rect -491 -9330 -421 -9311
rect -491 -9364 -472 -9330
rect -438 -9364 -421 -9330
rect -661 -9459 -627 -9440
rect -864 -9550 -856 -9516
rect -822 -9550 -814 -9516
rect -780 -9475 -627 -9459
rect -491 -9474 -421 -9364
rect -328 -9330 -262 -9277
rect -328 -9364 -312 -9330
rect -278 -9364 -262 -9330
rect -328 -9373 -262 -9364
rect -228 -9330 -162 -9311
rect -228 -9364 -215 -9330
rect -181 -9364 -162 -9330
rect -228 -9407 -162 -9364
rect -356 -9441 -162 -9407
rect -128 -9371 -70 -9277
rect -128 -9405 -116 -9371
rect -82 -9405 -70 -9371
rect -128 -9422 -70 -9405
rect -36 -9345 298 -9277
rect -36 -9379 -18 -9345
rect 16 -9379 246 -9345
rect 280 -9379 298 -9345
rect -36 -9431 298 -9379
rect 332 -9371 390 -9277
rect 332 -9405 344 -9371
rect 378 -9405 390 -9371
rect 332 -9422 390 -9405
rect 424 -9330 505 -9311
rect 424 -9364 457 -9330
rect 491 -9364 505 -9330
rect 424 -9388 505 -9364
rect 539 -9330 605 -9277
rect 539 -9364 555 -9330
rect 589 -9364 605 -9330
rect 539 -9380 605 -9364
rect 695 -9330 745 -9311
rect 695 -9364 711 -9330
rect -356 -9465 -286 -9441
rect -780 -9509 -777 -9475
rect -743 -9509 -627 -9475
rect -780 -9525 -627 -9509
rect -593 -9475 -421 -9474
rect -593 -9509 -577 -9475
rect -543 -9509 -421 -9475
rect -593 -9524 -421 -9509
rect -372 -9475 -286 -9465
rect -372 -9509 -356 -9475
rect -322 -9509 -286 -9475
rect -372 -9523 -286 -9509
rect -252 -9509 -236 -9475
rect -202 -9481 -162 -9475
rect -252 -9515 -210 -9509
rect -176 -9515 -162 -9481
rect -252 -9518 -162 -9515
rect -36 -9499 -16 -9465
rect 18 -9499 114 -9465
rect -1600 -9609 -898 -9569
rect -1600 -9643 -1582 -9609
rect -1548 -9643 -950 -9609
rect -916 -9643 -898 -9609
rect -1600 -9711 -898 -9643
rect -1600 -9745 -1582 -9711
rect -1548 -9745 -950 -9711
rect -916 -9745 -898 -9711
rect -1600 -9787 -898 -9745
rect -864 -9598 -814 -9550
rect -661 -9559 -627 -9525
rect -661 -9593 -543 -9559
rect -864 -9635 -783 -9598
rect -864 -9669 -831 -9635
rect -797 -9669 -783 -9635
rect -864 -9703 -783 -9669
rect -864 -9737 -831 -9703
rect -797 -9737 -783 -9703
rect -864 -9753 -783 -9737
rect -749 -9636 -683 -9627
rect -749 -9670 -733 -9636
rect -699 -9670 -683 -9636
rect -749 -9704 -683 -9670
rect -749 -9738 -733 -9704
rect -699 -9738 -683 -9704
rect -749 -9787 -683 -9738
rect -593 -9635 -543 -9593
rect -593 -9669 -577 -9635
rect -593 -9703 -543 -9669
rect -593 -9737 -577 -9703
rect -593 -9753 -543 -9737
rect -491 -9636 -421 -9524
rect -356 -9552 -286 -9523
rect -356 -9586 -162 -9552
rect -491 -9670 -473 -9636
rect -439 -9670 -421 -9636
rect -491 -9704 -421 -9670
rect -491 -9738 -473 -9704
rect -439 -9738 -421 -9704
rect -491 -9753 -421 -9738
rect -331 -9636 -265 -9620
rect -331 -9670 -315 -9636
rect -281 -9670 -265 -9636
rect -331 -9704 -265 -9670
rect -331 -9738 -315 -9704
rect -281 -9738 -265 -9704
rect -331 -9787 -265 -9738
rect -231 -9636 -162 -9586
rect -231 -9670 -215 -9636
rect -181 -9670 -162 -9636
rect -231 -9704 -162 -9670
rect -231 -9738 -215 -9704
rect -181 -9738 -162 -9704
rect -231 -9753 -162 -9738
rect -128 -9589 -70 -9554
rect -128 -9623 -116 -9589
rect -82 -9623 -70 -9589
rect -128 -9682 -70 -9623
rect -128 -9716 -116 -9682
rect -82 -9716 -70 -9682
rect -128 -9787 -70 -9716
rect -36 -9569 114 -9499
rect 148 -9501 298 -9431
rect 148 -9535 244 -9501
rect 278 -9535 298 -9501
rect 424 -9516 474 -9388
rect 695 -9406 745 -9364
rect 627 -9440 745 -9406
rect 797 -9330 867 -9311
rect 797 -9364 816 -9330
rect 850 -9364 867 -9330
rect 627 -9459 661 -9440
rect 424 -9550 432 -9516
rect 466 -9550 474 -9516
rect 508 -9475 661 -9459
rect 797 -9474 867 -9364
rect 960 -9330 1026 -9277
rect 960 -9364 976 -9330
rect 1010 -9364 1026 -9330
rect 960 -9373 1026 -9364
rect 1060 -9330 1126 -9311
rect 1060 -9364 1073 -9330
rect 1107 -9364 1126 -9330
rect 1060 -9407 1126 -9364
rect 932 -9441 1126 -9407
rect 1160 -9371 1218 -9277
rect 1160 -9405 1172 -9371
rect 1206 -9405 1218 -9371
rect 1160 -9422 1218 -9405
rect 1252 -9345 1586 -9277
rect 1252 -9379 1270 -9345
rect 1304 -9379 1534 -9345
rect 1568 -9379 1586 -9345
rect 1252 -9431 1586 -9379
rect 1620 -9371 1678 -9277
rect 1620 -9405 1632 -9371
rect 1666 -9405 1678 -9371
rect 1620 -9422 1678 -9405
rect 1712 -9338 2414 -9277
rect 1712 -9372 1730 -9338
rect 1764 -9372 2362 -9338
rect 2396 -9372 2414 -9338
rect 1712 -9431 2414 -9372
rect 2448 -9371 2506 -9277
rect 2448 -9405 2460 -9371
rect 2494 -9405 2506 -9371
rect 2448 -9422 2506 -9405
rect 2540 -9345 2874 -9277
rect 2540 -9379 2558 -9345
rect 2592 -9379 2822 -9345
rect 2856 -9379 2874 -9345
rect 2540 -9431 2874 -9379
rect 2908 -9371 2966 -9277
rect 2908 -9405 2920 -9371
rect 2954 -9405 2966 -9371
rect 2908 -9422 2966 -9405
rect 3000 -9330 3081 -9311
rect 3000 -9364 3033 -9330
rect 3067 -9364 3081 -9330
rect 3000 -9388 3081 -9364
rect 3115 -9330 3181 -9277
rect 3115 -9364 3131 -9330
rect 3165 -9364 3181 -9330
rect 3115 -9380 3181 -9364
rect 3271 -9330 3321 -9311
rect 3271 -9364 3287 -9330
rect 932 -9465 1002 -9441
rect 508 -9509 511 -9475
rect 545 -9509 661 -9475
rect 508 -9525 661 -9509
rect 695 -9475 867 -9474
rect 695 -9509 711 -9475
rect 745 -9509 867 -9475
rect 695 -9524 867 -9509
rect 916 -9475 1002 -9465
rect 916 -9509 932 -9475
rect 966 -9509 1002 -9475
rect 916 -9523 1002 -9509
rect 1036 -9509 1052 -9475
rect 1086 -9482 1126 -9475
rect 1036 -9516 1054 -9509
rect 1088 -9516 1126 -9482
rect 1036 -9518 1126 -9516
rect 1252 -9499 1272 -9465
rect 1306 -9499 1402 -9465
rect -36 -9609 298 -9569
rect -36 -9643 -18 -9609
rect 16 -9643 246 -9609
rect 280 -9643 298 -9609
rect -36 -9711 298 -9643
rect -36 -9745 -18 -9711
rect 16 -9745 246 -9711
rect 280 -9745 298 -9711
rect -36 -9787 298 -9745
rect 332 -9589 390 -9554
rect 332 -9623 344 -9589
rect 378 -9623 390 -9589
rect 332 -9682 390 -9623
rect 332 -9716 344 -9682
rect 378 -9716 390 -9682
rect 332 -9787 390 -9716
rect 424 -9598 474 -9550
rect 627 -9559 661 -9525
rect 627 -9593 745 -9559
rect 424 -9635 505 -9598
rect 424 -9669 457 -9635
rect 491 -9669 505 -9635
rect 424 -9703 505 -9669
rect 424 -9737 457 -9703
rect 491 -9737 505 -9703
rect 424 -9753 505 -9737
rect 539 -9636 605 -9627
rect 539 -9670 555 -9636
rect 589 -9670 605 -9636
rect 539 -9704 605 -9670
rect 539 -9738 555 -9704
rect 589 -9738 605 -9704
rect 539 -9787 605 -9738
rect 695 -9635 745 -9593
rect 695 -9669 711 -9635
rect 695 -9703 745 -9669
rect 695 -9737 711 -9703
rect 695 -9753 745 -9737
rect 797 -9636 867 -9524
rect 932 -9552 1002 -9523
rect 932 -9586 1126 -9552
rect 797 -9670 815 -9636
rect 849 -9670 867 -9636
rect 797 -9704 867 -9670
rect 797 -9738 815 -9704
rect 849 -9738 867 -9704
rect 797 -9753 867 -9738
rect 957 -9636 1023 -9620
rect 957 -9670 973 -9636
rect 1007 -9670 1023 -9636
rect 957 -9704 1023 -9670
rect 957 -9738 973 -9704
rect 1007 -9738 1023 -9704
rect 957 -9787 1023 -9738
rect 1057 -9636 1126 -9586
rect 1057 -9670 1073 -9636
rect 1107 -9670 1126 -9636
rect 1057 -9704 1126 -9670
rect 1057 -9738 1073 -9704
rect 1107 -9738 1126 -9704
rect 1057 -9753 1126 -9738
rect 1160 -9589 1218 -9554
rect 1160 -9623 1172 -9589
rect 1206 -9623 1218 -9589
rect 1160 -9682 1218 -9623
rect 1160 -9716 1172 -9682
rect 1206 -9716 1218 -9682
rect 1160 -9787 1218 -9716
rect 1252 -9569 1402 -9499
rect 1436 -9501 1586 -9431
rect 1436 -9535 1532 -9501
rect 1566 -9535 1586 -9501
rect 1712 -9499 1790 -9465
rect 1824 -9499 1893 -9465
rect 1927 -9499 1996 -9465
rect 2030 -9499 2050 -9465
rect 1252 -9609 1586 -9569
rect 1252 -9643 1270 -9609
rect 1304 -9643 1534 -9609
rect 1568 -9643 1586 -9609
rect 1252 -9711 1586 -9643
rect 1252 -9745 1270 -9711
rect 1304 -9745 1534 -9711
rect 1568 -9745 1586 -9711
rect 1252 -9787 1586 -9745
rect 1620 -9589 1678 -9554
rect 1620 -9623 1632 -9589
rect 1666 -9623 1678 -9589
rect 1620 -9682 1678 -9623
rect 1620 -9716 1632 -9682
rect 1666 -9716 1678 -9682
rect 1620 -9787 1678 -9716
rect 1712 -9569 2050 -9499
rect 2084 -9501 2414 -9431
rect 2084 -9535 2104 -9501
rect 2138 -9535 2203 -9501
rect 2237 -9535 2302 -9501
rect 2336 -9535 2414 -9501
rect 2540 -9499 2560 -9465
rect 2594 -9499 2690 -9465
rect 1712 -9609 2414 -9569
rect 1712 -9643 1730 -9609
rect 1764 -9643 2362 -9609
rect 2396 -9643 2414 -9609
rect 1712 -9711 2414 -9643
rect 1712 -9745 1730 -9711
rect 1764 -9745 2362 -9711
rect 2396 -9745 2414 -9711
rect 1712 -9787 2414 -9745
rect 2448 -9589 2506 -9554
rect 2448 -9623 2460 -9589
rect 2494 -9623 2506 -9589
rect 2448 -9682 2506 -9623
rect 2448 -9716 2460 -9682
rect 2494 -9716 2506 -9682
rect 2448 -9787 2506 -9716
rect 2540 -9569 2690 -9499
rect 2724 -9501 2874 -9431
rect 2724 -9535 2820 -9501
rect 2854 -9535 2874 -9501
rect 3000 -9482 3050 -9388
rect 3271 -9406 3321 -9364
rect 3203 -9440 3321 -9406
rect 3373 -9330 3443 -9311
rect 3373 -9364 3392 -9330
rect 3426 -9364 3443 -9330
rect 3203 -9459 3237 -9440
rect 3000 -9516 3014 -9482
rect 3048 -9516 3050 -9482
rect 2540 -9609 2874 -9569
rect 2540 -9643 2558 -9609
rect 2592 -9643 2822 -9609
rect 2856 -9643 2874 -9609
rect 2540 -9711 2874 -9643
rect 2540 -9745 2558 -9711
rect 2592 -9745 2822 -9711
rect 2856 -9745 2874 -9711
rect 2540 -9787 2874 -9745
rect 2908 -9589 2966 -9554
rect 2908 -9623 2920 -9589
rect 2954 -9623 2966 -9589
rect 2908 -9682 2966 -9623
rect 2908 -9716 2920 -9682
rect 2954 -9716 2966 -9682
rect 2908 -9787 2966 -9716
rect 3000 -9598 3050 -9516
rect 3084 -9475 3237 -9459
rect 3373 -9474 3443 -9364
rect 3536 -9330 3602 -9277
rect 3536 -9364 3552 -9330
rect 3586 -9364 3602 -9330
rect 3536 -9373 3602 -9364
rect 3636 -9330 3702 -9311
rect 3636 -9364 3649 -9330
rect 3683 -9364 3702 -9330
rect 3636 -9407 3702 -9364
rect 3508 -9441 3702 -9407
rect 3736 -9371 3794 -9277
rect 3736 -9405 3748 -9371
rect 3782 -9405 3794 -9371
rect 3736 -9422 3794 -9405
rect 3828 -9345 4162 -9277
rect 3828 -9379 3846 -9345
rect 3880 -9379 4110 -9345
rect 4144 -9379 4162 -9345
rect 3828 -9431 4162 -9379
rect 4196 -9371 4254 -9277
rect 4196 -9405 4208 -9371
rect 4242 -9405 4254 -9371
rect 4196 -9422 4254 -9405
rect 4288 -9338 4990 -9277
rect 4288 -9372 4306 -9338
rect 4340 -9372 4938 -9338
rect 4972 -9372 4990 -9338
rect 4288 -9431 4990 -9372
rect 5024 -9371 5082 -9277
rect 5024 -9405 5036 -9371
rect 5070 -9405 5082 -9371
rect 5024 -9422 5082 -9405
rect 5116 -9345 5450 -9277
rect 5116 -9379 5134 -9345
rect 5168 -9379 5398 -9345
rect 5432 -9379 5450 -9345
rect 5116 -9431 5450 -9379
rect 5484 -9371 5542 -9277
rect 5484 -9405 5496 -9371
rect 5530 -9405 5542 -9371
rect 5484 -9422 5542 -9405
rect 5576 -9330 5657 -9311
rect 5576 -9364 5609 -9330
rect 5643 -9364 5657 -9330
rect 5576 -9388 5657 -9364
rect 5691 -9330 5757 -9277
rect 5691 -9364 5707 -9330
rect 5741 -9364 5757 -9330
rect 5691 -9380 5757 -9364
rect 5847 -9330 5897 -9311
rect 5847 -9364 5863 -9330
rect 3508 -9465 3578 -9441
rect 3084 -9509 3087 -9475
rect 3121 -9509 3237 -9475
rect 3084 -9525 3237 -9509
rect 3271 -9475 3443 -9474
rect 3271 -9509 3287 -9475
rect 3321 -9509 3443 -9475
rect 3271 -9524 3443 -9509
rect 3492 -9475 3578 -9465
rect 3492 -9509 3508 -9475
rect 3542 -9509 3578 -9475
rect 3492 -9523 3578 -9509
rect 3612 -9516 3628 -9475
rect 3662 -9516 3702 -9475
rect 3612 -9518 3702 -9516
rect 3828 -9499 3848 -9465
rect 3882 -9499 3978 -9465
rect 3203 -9559 3237 -9525
rect 3203 -9593 3321 -9559
rect 3000 -9635 3081 -9598
rect 3000 -9669 3033 -9635
rect 3067 -9669 3081 -9635
rect 3000 -9703 3081 -9669
rect 3000 -9737 3033 -9703
rect 3067 -9737 3081 -9703
rect 3000 -9753 3081 -9737
rect 3115 -9636 3181 -9627
rect 3115 -9670 3131 -9636
rect 3165 -9670 3181 -9636
rect 3115 -9704 3181 -9670
rect 3115 -9738 3131 -9704
rect 3165 -9738 3181 -9704
rect 3115 -9787 3181 -9738
rect 3271 -9635 3321 -9593
rect 3271 -9669 3287 -9635
rect 3271 -9703 3321 -9669
rect 3271 -9737 3287 -9703
rect 3271 -9753 3321 -9737
rect 3373 -9636 3443 -9524
rect 3508 -9552 3578 -9523
rect 3508 -9586 3702 -9552
rect 3373 -9670 3391 -9636
rect 3425 -9670 3443 -9636
rect 3373 -9704 3443 -9670
rect 3373 -9738 3391 -9704
rect 3425 -9738 3443 -9704
rect 3373 -9753 3443 -9738
rect 3533 -9636 3599 -9620
rect 3533 -9670 3549 -9636
rect 3583 -9670 3599 -9636
rect 3533 -9704 3599 -9670
rect 3533 -9738 3549 -9704
rect 3583 -9738 3599 -9704
rect 3533 -9787 3599 -9738
rect 3633 -9636 3702 -9586
rect 3633 -9670 3649 -9636
rect 3683 -9670 3702 -9636
rect 3633 -9704 3702 -9670
rect 3633 -9738 3649 -9704
rect 3683 -9738 3702 -9704
rect 3633 -9753 3702 -9738
rect 3736 -9589 3794 -9554
rect 3736 -9623 3748 -9589
rect 3782 -9623 3794 -9589
rect 3736 -9682 3794 -9623
rect 3736 -9716 3748 -9682
rect 3782 -9716 3794 -9682
rect 3736 -9787 3794 -9716
rect 3828 -9569 3978 -9499
rect 4012 -9501 4162 -9431
rect 4012 -9535 4108 -9501
rect 4142 -9535 4162 -9501
rect 4288 -9499 4366 -9465
rect 4400 -9499 4469 -9465
rect 4503 -9499 4572 -9465
rect 4606 -9499 4626 -9465
rect 3828 -9609 4162 -9569
rect 3828 -9643 3846 -9609
rect 3880 -9643 4110 -9609
rect 4144 -9643 4162 -9609
rect 3828 -9711 4162 -9643
rect 3828 -9745 3846 -9711
rect 3880 -9745 4110 -9711
rect 4144 -9745 4162 -9711
rect 3828 -9787 4162 -9745
rect 4196 -9589 4254 -9554
rect 4196 -9623 4208 -9589
rect 4242 -9623 4254 -9589
rect 4196 -9682 4254 -9623
rect 4196 -9716 4208 -9682
rect 4242 -9716 4254 -9682
rect 4196 -9787 4254 -9716
rect 4288 -9569 4626 -9499
rect 4660 -9501 4990 -9431
rect 4660 -9535 4680 -9501
rect 4714 -9535 4779 -9501
rect 4813 -9535 4878 -9501
rect 4912 -9535 4990 -9501
rect 5116 -9499 5136 -9465
rect 5170 -9499 5266 -9465
rect 4288 -9609 4990 -9569
rect 4288 -9643 4306 -9609
rect 4340 -9643 4938 -9609
rect 4972 -9643 4990 -9609
rect 4288 -9711 4990 -9643
rect 4288 -9745 4306 -9711
rect 4340 -9745 4938 -9711
rect 4972 -9745 4990 -9711
rect 4288 -9787 4990 -9745
rect 5024 -9589 5082 -9554
rect 5024 -9623 5036 -9589
rect 5070 -9623 5082 -9589
rect 5024 -9682 5082 -9623
rect 5024 -9716 5036 -9682
rect 5070 -9716 5082 -9682
rect 5024 -9787 5082 -9716
rect 5116 -9569 5266 -9499
rect 5300 -9501 5450 -9431
rect 5300 -9535 5396 -9501
rect 5430 -9535 5450 -9501
rect 5576 -9482 5626 -9388
rect 5847 -9406 5897 -9364
rect 5779 -9440 5897 -9406
rect 5949 -9330 6019 -9311
rect 5949 -9364 5968 -9330
rect 6002 -9364 6019 -9330
rect 5779 -9459 5813 -9440
rect 5576 -9516 5588 -9482
rect 5622 -9516 5626 -9482
rect 5116 -9609 5450 -9569
rect 5116 -9643 5134 -9609
rect 5168 -9643 5398 -9609
rect 5432 -9643 5450 -9609
rect 5116 -9711 5450 -9643
rect 5116 -9745 5134 -9711
rect 5168 -9745 5398 -9711
rect 5432 -9745 5450 -9711
rect 5116 -9787 5450 -9745
rect 5484 -9589 5542 -9554
rect 5484 -9623 5496 -9589
rect 5530 -9623 5542 -9589
rect 5484 -9682 5542 -9623
rect 5484 -9716 5496 -9682
rect 5530 -9716 5542 -9682
rect 5484 -9787 5542 -9716
rect 5576 -9598 5626 -9516
rect 5660 -9475 5813 -9459
rect 5949 -9474 6019 -9364
rect 6112 -9330 6178 -9277
rect 6112 -9364 6128 -9330
rect 6162 -9364 6178 -9330
rect 6112 -9373 6178 -9364
rect 6212 -9330 6278 -9311
rect 6212 -9364 6225 -9330
rect 6259 -9364 6278 -9330
rect 6212 -9407 6278 -9364
rect 6084 -9441 6278 -9407
rect 6312 -9371 6370 -9277
rect 6312 -9405 6324 -9371
rect 6358 -9405 6370 -9371
rect 6312 -9422 6370 -9405
rect 6404 -9345 6738 -9277
rect 6404 -9379 6422 -9345
rect 6456 -9379 6686 -9345
rect 6720 -9379 6738 -9345
rect 6404 -9431 6738 -9379
rect 6772 -9371 6830 -9277
rect 6772 -9405 6784 -9371
rect 6818 -9405 6830 -9371
rect 6772 -9422 6830 -9405
rect 6864 -9338 7566 -9277
rect 6864 -9372 6882 -9338
rect 6916 -9372 7514 -9338
rect 7548 -9372 7566 -9338
rect 6864 -9431 7566 -9372
rect 7600 -9371 7658 -9277
rect 7600 -9405 7612 -9371
rect 7646 -9405 7658 -9371
rect 7600 -9422 7658 -9405
rect 7692 -9345 8026 -9277
rect 7692 -9379 7710 -9345
rect 7744 -9379 7974 -9345
rect 8008 -9379 8026 -9345
rect 7692 -9431 8026 -9379
rect 8060 -9371 8118 -9277
rect 8060 -9405 8072 -9371
rect 8106 -9405 8118 -9371
rect 8060 -9422 8118 -9405
rect 8152 -9330 8233 -9311
rect 8152 -9364 8185 -9330
rect 8219 -9364 8233 -9330
rect 8152 -9388 8233 -9364
rect 8267 -9330 8333 -9277
rect 8267 -9364 8283 -9330
rect 8317 -9364 8333 -9330
rect 8267 -9380 8333 -9364
rect 8423 -9330 8473 -9311
rect 8423 -9364 8439 -9330
rect 6084 -9465 6154 -9441
rect 5660 -9509 5663 -9475
rect 5697 -9509 5813 -9475
rect 5660 -9525 5813 -9509
rect 5847 -9475 6019 -9474
rect 5847 -9509 5863 -9475
rect 5897 -9509 6019 -9475
rect 5847 -9524 6019 -9509
rect 6068 -9475 6154 -9465
rect 6068 -9509 6084 -9475
rect 6118 -9509 6154 -9475
rect 6068 -9523 6154 -9509
rect 6188 -9482 6204 -9475
rect 6188 -9516 6202 -9482
rect 6238 -9509 6278 -9475
rect 6236 -9516 6278 -9509
rect 6188 -9518 6278 -9516
rect 6404 -9499 6424 -9465
rect 6458 -9499 6554 -9465
rect 5779 -9559 5813 -9525
rect 5779 -9593 5897 -9559
rect 5576 -9635 5657 -9598
rect 5576 -9669 5609 -9635
rect 5643 -9669 5657 -9635
rect 5576 -9703 5657 -9669
rect 5576 -9737 5609 -9703
rect 5643 -9737 5657 -9703
rect 5576 -9753 5657 -9737
rect 5691 -9636 5757 -9627
rect 5691 -9670 5707 -9636
rect 5741 -9670 5757 -9636
rect 5691 -9704 5757 -9670
rect 5691 -9738 5707 -9704
rect 5741 -9738 5757 -9704
rect 5691 -9787 5757 -9738
rect 5847 -9635 5897 -9593
rect 5847 -9669 5863 -9635
rect 5847 -9703 5897 -9669
rect 5847 -9737 5863 -9703
rect 5847 -9753 5897 -9737
rect 5949 -9636 6019 -9524
rect 6084 -9552 6154 -9523
rect 6084 -9586 6278 -9552
rect 5949 -9670 5967 -9636
rect 6001 -9670 6019 -9636
rect 5949 -9704 6019 -9670
rect 5949 -9738 5967 -9704
rect 6001 -9738 6019 -9704
rect 5949 -9753 6019 -9738
rect 6109 -9636 6175 -9620
rect 6109 -9670 6125 -9636
rect 6159 -9670 6175 -9636
rect 6109 -9704 6175 -9670
rect 6109 -9738 6125 -9704
rect 6159 -9738 6175 -9704
rect 6109 -9787 6175 -9738
rect 6209 -9636 6278 -9586
rect 6209 -9670 6225 -9636
rect 6259 -9670 6278 -9636
rect 6209 -9704 6278 -9670
rect 6209 -9738 6225 -9704
rect 6259 -9738 6278 -9704
rect 6209 -9753 6278 -9738
rect 6312 -9589 6370 -9554
rect 6312 -9623 6324 -9589
rect 6358 -9623 6370 -9589
rect 6312 -9682 6370 -9623
rect 6312 -9716 6324 -9682
rect 6358 -9716 6370 -9682
rect 6312 -9787 6370 -9716
rect 6404 -9569 6554 -9499
rect 6588 -9501 6738 -9431
rect 6588 -9535 6684 -9501
rect 6718 -9535 6738 -9501
rect 6864 -9499 6942 -9465
rect 6976 -9499 7045 -9465
rect 7079 -9499 7148 -9465
rect 7182 -9499 7202 -9465
rect 6404 -9609 6738 -9569
rect 6404 -9643 6422 -9609
rect 6456 -9643 6686 -9609
rect 6720 -9643 6738 -9609
rect 6404 -9711 6738 -9643
rect 6404 -9745 6422 -9711
rect 6456 -9745 6686 -9711
rect 6720 -9745 6738 -9711
rect 6404 -9787 6738 -9745
rect 6772 -9589 6830 -9554
rect 6772 -9623 6784 -9589
rect 6818 -9623 6830 -9589
rect 6772 -9682 6830 -9623
rect 6772 -9716 6784 -9682
rect 6818 -9716 6830 -9682
rect 6772 -9787 6830 -9716
rect 6864 -9569 7202 -9499
rect 7236 -9501 7566 -9431
rect 7236 -9535 7256 -9501
rect 7290 -9535 7355 -9501
rect 7389 -9535 7454 -9501
rect 7488 -9535 7566 -9501
rect 7692 -9499 7712 -9465
rect 7746 -9499 7842 -9465
rect 6864 -9609 7566 -9569
rect 6864 -9643 6882 -9609
rect 6916 -9643 7514 -9609
rect 7548 -9643 7566 -9609
rect 6864 -9711 7566 -9643
rect 6864 -9745 6882 -9711
rect 6916 -9745 7514 -9711
rect 7548 -9745 7566 -9711
rect 6864 -9787 7566 -9745
rect 7600 -9589 7658 -9554
rect 7600 -9623 7612 -9589
rect 7646 -9623 7658 -9589
rect 7600 -9682 7658 -9623
rect 7600 -9716 7612 -9682
rect 7646 -9716 7658 -9682
rect 7600 -9787 7658 -9716
rect 7692 -9569 7842 -9499
rect 7876 -9501 8026 -9431
rect 7876 -9535 7972 -9501
rect 8006 -9535 8026 -9501
rect 8152 -9482 8202 -9388
rect 8423 -9406 8473 -9364
rect 8355 -9440 8473 -9406
rect 8525 -9330 8595 -9311
rect 8525 -9364 8544 -9330
rect 8578 -9364 8595 -9330
rect 8355 -9459 8389 -9440
rect 8152 -9516 8162 -9482
rect 8196 -9516 8202 -9482
rect 7692 -9609 8026 -9569
rect 7692 -9643 7710 -9609
rect 7744 -9643 7974 -9609
rect 8008 -9643 8026 -9609
rect 7692 -9711 8026 -9643
rect 7692 -9745 7710 -9711
rect 7744 -9745 7974 -9711
rect 8008 -9745 8026 -9711
rect 7692 -9787 8026 -9745
rect 8060 -9589 8118 -9554
rect 8060 -9623 8072 -9589
rect 8106 -9623 8118 -9589
rect 8060 -9682 8118 -9623
rect 8060 -9716 8072 -9682
rect 8106 -9716 8118 -9682
rect 8060 -9787 8118 -9716
rect 8152 -9598 8202 -9516
rect 8236 -9475 8389 -9459
rect 8525 -9474 8595 -9364
rect 8688 -9330 8754 -9277
rect 8688 -9364 8704 -9330
rect 8738 -9364 8754 -9330
rect 8688 -9373 8754 -9364
rect 8788 -9330 8854 -9311
rect 8788 -9364 8801 -9330
rect 8835 -9364 8854 -9330
rect 8788 -9407 8854 -9364
rect 8660 -9441 8854 -9407
rect 8888 -9371 8946 -9277
rect 8888 -9405 8900 -9371
rect 8934 -9405 8946 -9371
rect 8888 -9422 8946 -9405
rect 8980 -9345 9314 -9277
rect 8980 -9379 8998 -9345
rect 9032 -9379 9262 -9345
rect 9296 -9379 9314 -9345
rect 8980 -9431 9314 -9379
rect 9348 -9371 9406 -9277
rect 9348 -9405 9360 -9371
rect 9394 -9405 9406 -9371
rect 9348 -9422 9406 -9405
rect 9440 -9338 10142 -9277
rect 9440 -9372 9458 -9338
rect 9492 -9372 10090 -9338
rect 10124 -9372 10142 -9338
rect 9440 -9431 10142 -9372
rect 10176 -9371 10234 -9277
rect 10176 -9405 10188 -9371
rect 10222 -9405 10234 -9371
rect 10176 -9422 10234 -9405
rect 10360 -9345 10694 -9277
rect 10360 -9379 10378 -9345
rect 10412 -9379 10642 -9345
rect 10676 -9379 10694 -9345
rect 10360 -9431 10694 -9379
rect 8660 -9465 8730 -9441
rect 8236 -9509 8239 -9475
rect 8273 -9509 8389 -9475
rect 8236 -9525 8389 -9509
rect 8423 -9475 8595 -9474
rect 8423 -9509 8439 -9475
rect 8473 -9509 8595 -9475
rect 8423 -9524 8595 -9509
rect 8644 -9475 8730 -9465
rect 8644 -9509 8660 -9475
rect 8694 -9509 8730 -9475
rect 8644 -9523 8730 -9509
rect 8764 -9482 8780 -9475
rect 8764 -9516 8776 -9482
rect 8814 -9509 8854 -9475
rect 8810 -9516 8854 -9509
rect 8764 -9518 8854 -9516
rect 8980 -9499 9000 -9465
rect 9034 -9499 9130 -9465
rect 8355 -9559 8389 -9525
rect 8355 -9593 8473 -9559
rect 8152 -9635 8233 -9598
rect 8152 -9669 8185 -9635
rect 8219 -9669 8233 -9635
rect 8152 -9703 8233 -9669
rect 8152 -9737 8185 -9703
rect 8219 -9737 8233 -9703
rect 8152 -9753 8233 -9737
rect 8267 -9636 8333 -9627
rect 8267 -9670 8283 -9636
rect 8317 -9670 8333 -9636
rect 8267 -9704 8333 -9670
rect 8267 -9738 8283 -9704
rect 8317 -9738 8333 -9704
rect 8267 -9787 8333 -9738
rect 8423 -9635 8473 -9593
rect 8423 -9669 8439 -9635
rect 8423 -9703 8473 -9669
rect 8423 -9737 8439 -9703
rect 8423 -9753 8473 -9737
rect 8525 -9636 8595 -9524
rect 8660 -9552 8730 -9523
rect 8660 -9586 8854 -9552
rect 8525 -9670 8543 -9636
rect 8577 -9670 8595 -9636
rect 8525 -9704 8595 -9670
rect 8525 -9738 8543 -9704
rect 8577 -9738 8595 -9704
rect 8525 -9753 8595 -9738
rect 8685 -9636 8751 -9620
rect 8685 -9670 8701 -9636
rect 8735 -9670 8751 -9636
rect 8685 -9704 8751 -9670
rect 8685 -9738 8701 -9704
rect 8735 -9738 8751 -9704
rect 8685 -9787 8751 -9738
rect 8785 -9636 8854 -9586
rect 8785 -9670 8801 -9636
rect 8835 -9670 8854 -9636
rect 8785 -9704 8854 -9670
rect 8785 -9738 8801 -9704
rect 8835 -9738 8854 -9704
rect 8785 -9753 8854 -9738
rect 8888 -9589 8946 -9554
rect 8888 -9623 8900 -9589
rect 8934 -9623 8946 -9589
rect 8888 -9682 8946 -9623
rect 8888 -9716 8900 -9682
rect 8934 -9716 8946 -9682
rect 8888 -9787 8946 -9716
rect 8980 -9569 9130 -9499
rect 9164 -9501 9314 -9431
rect 9164 -9535 9260 -9501
rect 9294 -9535 9314 -9501
rect 9440 -9499 9518 -9465
rect 9552 -9499 9621 -9465
rect 9655 -9499 9724 -9465
rect 9758 -9499 9778 -9465
rect 8980 -9609 9314 -9569
rect 8980 -9643 8998 -9609
rect 9032 -9643 9262 -9609
rect 9296 -9643 9314 -9609
rect 8980 -9711 9314 -9643
rect 8980 -9745 8998 -9711
rect 9032 -9745 9262 -9711
rect 9296 -9745 9314 -9711
rect 8980 -9787 9314 -9745
rect 9348 -9589 9406 -9554
rect 9348 -9623 9360 -9589
rect 9394 -9623 9406 -9589
rect 9348 -9682 9406 -9623
rect 9348 -9716 9360 -9682
rect 9394 -9716 9406 -9682
rect 9348 -9787 9406 -9716
rect 9440 -9569 9778 -9499
rect 9812 -9501 10142 -9431
rect 9812 -9535 9832 -9501
rect 9866 -9535 9931 -9501
rect 9965 -9535 10030 -9501
rect 10064 -9535 10142 -9501
rect 10360 -9499 10380 -9465
rect 10414 -9499 10510 -9465
rect 9440 -9609 10142 -9569
rect 9440 -9643 9458 -9609
rect 9492 -9643 10090 -9609
rect 10124 -9643 10142 -9609
rect 9440 -9711 10142 -9643
rect 9440 -9745 9458 -9711
rect 9492 -9745 10090 -9711
rect 10124 -9745 10142 -9711
rect 9440 -9787 10142 -9745
rect 10176 -9589 10234 -9554
rect 10176 -9623 10188 -9589
rect 10222 -9623 10234 -9589
rect 10176 -9682 10234 -9623
rect 10176 -9716 10188 -9682
rect 10222 -9716 10234 -9682
rect 10176 -9787 10234 -9716
rect 10360 -9569 10510 -9499
rect 10544 -9501 10694 -9431
rect 10544 -9535 10640 -9501
rect 10674 -9535 10694 -9501
rect 10728 -9330 10809 -9311
rect 10728 -9364 10761 -9330
rect 10795 -9364 10809 -9330
rect 10728 -9388 10809 -9364
rect 10843 -9330 10909 -9277
rect 10843 -9364 10859 -9330
rect 10893 -9364 10909 -9330
rect 10843 -9380 10909 -9364
rect 10999 -9330 11049 -9311
rect 10999 -9364 11015 -9330
rect 10728 -9482 10778 -9388
rect 10999 -9406 11049 -9364
rect 10931 -9440 11049 -9406
rect 11101 -9330 11171 -9311
rect 11101 -9364 11120 -9330
rect 11154 -9364 11171 -9330
rect 10931 -9459 10965 -9440
rect 10728 -9516 10736 -9482
rect 10770 -9516 10778 -9482
rect 10360 -9609 10694 -9569
rect 10360 -9643 10378 -9609
rect 10412 -9643 10642 -9609
rect 10676 -9643 10694 -9609
rect 10360 -9711 10694 -9643
rect 10360 -9745 10378 -9711
rect 10412 -9745 10642 -9711
rect 10676 -9745 10694 -9711
rect 10360 -9787 10694 -9745
rect 10728 -9598 10778 -9516
rect 10812 -9475 10965 -9459
rect 11101 -9474 11171 -9364
rect 11264 -9330 11330 -9277
rect 11264 -9364 11280 -9330
rect 11314 -9364 11330 -9330
rect 11264 -9373 11330 -9364
rect 11364 -9330 11430 -9311
rect 11364 -9364 11377 -9330
rect 11411 -9364 11430 -9330
rect 11364 -9407 11430 -9364
rect 11236 -9441 11430 -9407
rect 11464 -9371 11522 -9277
rect 11464 -9405 11476 -9371
rect 11510 -9405 11522 -9371
rect 11464 -9422 11522 -9405
rect 11648 -9345 11982 -9277
rect 11648 -9379 11666 -9345
rect 11700 -9379 11930 -9345
rect 11964 -9379 11982 -9345
rect 11648 -9431 11982 -9379
rect 13580 -9371 13638 -9277
rect 13580 -9405 13592 -9371
rect 13626 -9405 13638 -9371
rect 13672 -9319 13733 -9277
rect 13672 -9353 13690 -9319
rect 13724 -9353 13733 -9319
rect 13672 -9379 13733 -9353
rect 13769 -9332 13819 -9313
rect 13769 -9366 13776 -9332
rect 13810 -9366 13819 -9332
rect 13580 -9422 13638 -9405
rect 11236 -9465 11306 -9441
rect 10812 -9509 10815 -9475
rect 10849 -9509 10965 -9475
rect 10812 -9525 10965 -9509
rect 10999 -9475 11171 -9474
rect 10999 -9509 11015 -9475
rect 11049 -9509 11171 -9475
rect 10999 -9524 11171 -9509
rect 11220 -9475 11306 -9465
rect 11220 -9509 11236 -9475
rect 11270 -9509 11306 -9475
rect 11220 -9523 11306 -9509
rect 11340 -9509 11356 -9475
rect 11390 -9479 11430 -9475
rect 11340 -9513 11386 -9509
rect 11420 -9513 11430 -9479
rect 11340 -9518 11430 -9513
rect 11648 -9499 11668 -9465
rect 11702 -9499 11798 -9465
rect 10931 -9559 10965 -9525
rect 10931 -9593 11049 -9559
rect 10728 -9635 10809 -9598
rect 10728 -9669 10761 -9635
rect 10795 -9669 10809 -9635
rect 10728 -9703 10809 -9669
rect 10728 -9737 10761 -9703
rect 10795 -9737 10809 -9703
rect 10728 -9753 10809 -9737
rect 10843 -9636 10909 -9627
rect 10843 -9670 10859 -9636
rect 10893 -9670 10909 -9636
rect 10843 -9704 10909 -9670
rect 10843 -9738 10859 -9704
rect 10893 -9738 10909 -9704
rect 10843 -9787 10909 -9738
rect 10999 -9635 11049 -9593
rect 10999 -9669 11015 -9635
rect 10999 -9703 11049 -9669
rect 10999 -9737 11015 -9703
rect 10999 -9753 11049 -9737
rect 11101 -9636 11171 -9524
rect 11236 -9552 11306 -9523
rect 11236 -9586 11430 -9552
rect 11101 -9670 11119 -9636
rect 11153 -9670 11171 -9636
rect 11101 -9704 11171 -9670
rect 11101 -9738 11119 -9704
rect 11153 -9738 11171 -9704
rect 11101 -9753 11171 -9738
rect 11261 -9636 11327 -9620
rect 11261 -9670 11277 -9636
rect 11311 -9670 11327 -9636
rect 11261 -9704 11327 -9670
rect 11261 -9738 11277 -9704
rect 11311 -9738 11327 -9704
rect 11261 -9787 11327 -9738
rect 11361 -9636 11430 -9586
rect 11361 -9670 11377 -9636
rect 11411 -9670 11430 -9636
rect 11361 -9704 11430 -9670
rect 11361 -9738 11377 -9704
rect 11411 -9738 11430 -9704
rect 11361 -9753 11430 -9738
rect 11464 -9589 11522 -9554
rect 11464 -9623 11476 -9589
rect 11510 -9623 11522 -9589
rect 11464 -9682 11522 -9623
rect 11464 -9716 11476 -9682
rect 11510 -9716 11522 -9682
rect 11464 -9787 11522 -9716
rect 11648 -9569 11798 -9499
rect 11832 -9501 11982 -9431
rect 11832 -9535 11928 -9501
rect 11962 -9535 11982 -9501
rect 13672 -9448 13735 -9413
rect 13672 -9482 13685 -9448
rect 13719 -9475 13735 -9448
rect 13672 -9509 13692 -9482
rect 13726 -9509 13735 -9475
rect 13672 -9525 13735 -9509
rect 13769 -9475 13819 -9366
rect 13853 -9332 13905 -9277
rect 13853 -9366 13862 -9332
rect 13896 -9366 13905 -9332
rect 13853 -9382 13905 -9366
rect 13941 -9332 13991 -9313
rect 13941 -9366 13948 -9332
rect 13982 -9366 13991 -9332
rect 13941 -9475 13991 -9366
rect 14025 -9332 14077 -9277
rect 14025 -9366 14034 -9332
rect 14068 -9366 14077 -9332
rect 14025 -9389 14077 -9366
rect 14111 -9332 14163 -9316
rect 14111 -9366 14120 -9332
rect 14154 -9366 14163 -9332
rect 14111 -9407 14163 -9366
rect 14197 -9323 14249 -9277
rect 14197 -9357 14206 -9323
rect 14240 -9357 14249 -9323
rect 14197 -9373 14249 -9357
rect 14283 -9332 14335 -9316
rect 14283 -9366 14292 -9332
rect 14326 -9366 14335 -9332
rect 14283 -9407 14335 -9366
rect 14369 -9323 14421 -9277
rect 14369 -9357 14378 -9323
rect 14412 -9357 14421 -9323
rect 14369 -9373 14421 -9357
rect 14455 -9332 14507 -9316
rect 14455 -9366 14464 -9332
rect 14498 -9366 14507 -9332
rect 14455 -9407 14507 -9366
rect 14541 -9323 14590 -9277
rect 14541 -9357 14550 -9323
rect 14584 -9357 14590 -9323
rect 14541 -9373 14590 -9357
rect 14624 -9332 14679 -9316
rect 14624 -9366 14636 -9332
rect 14670 -9366 14679 -9332
rect 14624 -9407 14679 -9366
rect 14713 -9323 14762 -9277
rect 14713 -9357 14722 -9323
rect 14756 -9357 14762 -9323
rect 14713 -9373 14762 -9357
rect 14796 -9332 14848 -9316
rect 14796 -9366 14807 -9332
rect 14841 -9366 14848 -9332
rect 14796 -9407 14848 -9366
rect 14884 -9323 14934 -9277
rect 14884 -9357 14893 -9323
rect 14927 -9357 14934 -9323
rect 14884 -9373 14934 -9357
rect 14968 -9332 15020 -9316
rect 14968 -9366 14979 -9332
rect 15013 -9366 15020 -9332
rect 14968 -9407 15020 -9366
rect 15056 -9323 15106 -9277
rect 15056 -9357 15065 -9323
rect 15099 -9357 15106 -9323
rect 15056 -9373 15106 -9357
rect 15140 -9332 15192 -9316
rect 15140 -9366 15151 -9332
rect 15185 -9366 15192 -9332
rect 15140 -9407 15192 -9366
rect 15228 -9323 15280 -9277
rect 15228 -9357 15237 -9323
rect 15271 -9357 15280 -9323
rect 15228 -9373 15280 -9357
rect 15314 -9332 15366 -9316
rect 15314 -9366 15323 -9332
rect 15357 -9366 15366 -9332
rect 15314 -9407 15366 -9366
rect 15400 -9323 15460 -9277
rect 15400 -9357 15409 -9323
rect 15443 -9357 15460 -9323
rect 15400 -9373 15460 -9357
rect 15512 -9371 15570 -9277
rect 15512 -9405 15524 -9371
rect 15558 -9405 15570 -9371
rect 14111 -9432 15460 -9407
rect 15512 -9422 15570 -9405
rect 15605 -9338 16674 -9277
rect 15605 -9372 15622 -9338
rect 15656 -9372 16622 -9338
rect 16656 -9372 16674 -9338
rect 15605 -9431 16674 -9372
rect 14111 -9441 15248 -9432
rect 15227 -9466 15248 -9441
rect 15282 -9433 15460 -9432
rect 15282 -9466 15340 -9433
rect 15227 -9467 15340 -9466
rect 15374 -9467 15460 -9433
rect 13769 -9509 14119 -9475
rect 14153 -9509 14187 -9475
rect 14221 -9509 14255 -9475
rect 14289 -9509 14323 -9475
rect 14357 -9509 14391 -9475
rect 14425 -9509 14459 -9475
rect 14493 -9509 14527 -9475
rect 14561 -9509 14595 -9475
rect 14629 -9509 14663 -9475
rect 14697 -9509 14731 -9475
rect 14765 -9509 14799 -9475
rect 14833 -9509 14867 -9475
rect 14901 -9509 14935 -9475
rect 14969 -9509 15003 -9475
rect 15037 -9509 15071 -9475
rect 15105 -9509 15139 -9475
rect 15173 -9509 15193 -9475
rect 13769 -9525 15193 -9509
rect 11648 -9609 11982 -9569
rect 11648 -9643 11666 -9609
rect 11700 -9643 11930 -9609
rect 11964 -9643 11982 -9609
rect 11648 -9711 11982 -9643
rect 11648 -9745 11666 -9711
rect 11700 -9745 11930 -9711
rect 11964 -9745 11982 -9711
rect 11648 -9787 11982 -9745
rect 13580 -9589 13638 -9554
rect 13580 -9623 13592 -9589
rect 13626 -9623 13638 -9589
rect 13580 -9682 13638 -9623
rect 13580 -9716 13592 -9682
rect 13626 -9716 13638 -9682
rect 13580 -9787 13638 -9716
rect 13674 -9643 13733 -9625
rect 13674 -9677 13690 -9643
rect 13724 -9677 13733 -9643
rect 13674 -9711 13733 -9677
rect 13674 -9745 13690 -9711
rect 13724 -9745 13733 -9711
rect 13674 -9787 13733 -9745
rect 13769 -9635 13818 -9525
rect 13769 -9669 13776 -9635
rect 13810 -9669 13818 -9635
rect 13769 -9703 13818 -9669
rect 13769 -9737 13776 -9703
rect 13810 -9737 13818 -9703
rect 13769 -9753 13818 -9737
rect 13853 -9643 13905 -9625
rect 13853 -9677 13862 -9643
rect 13896 -9677 13905 -9643
rect 13853 -9711 13905 -9677
rect 13853 -9745 13862 -9711
rect 13896 -9745 13905 -9711
rect 13853 -9787 13905 -9745
rect 13941 -9627 13991 -9525
rect 15227 -9528 15460 -9467
rect 15227 -9559 15248 -9528
rect 14111 -9562 15248 -9559
rect 15282 -9562 15341 -9528
rect 15375 -9562 15460 -9528
rect 15605 -9499 15686 -9465
rect 15720 -9499 15814 -9465
rect 15848 -9499 15942 -9465
rect 15976 -9499 16070 -9465
rect 16104 -9499 16124 -9465
rect 14111 -9581 15460 -9562
rect 14111 -9615 14120 -9581
rect 14154 -9607 14292 -9581
rect 14154 -9615 14163 -9607
rect 13941 -9661 13948 -9627
rect 13982 -9661 13991 -9627
rect 13941 -9695 13991 -9661
rect 13941 -9729 13948 -9695
rect 13982 -9729 13991 -9695
rect 13941 -9752 13991 -9729
rect 14025 -9643 14077 -9627
rect 14025 -9677 14034 -9643
rect 14068 -9677 14077 -9643
rect 14025 -9711 14077 -9677
rect 14025 -9745 14034 -9711
rect 14068 -9745 14077 -9711
rect 14025 -9786 14077 -9745
rect 14111 -9667 14163 -9615
rect 14283 -9615 14292 -9607
rect 14326 -9607 14464 -9581
rect 14326 -9615 14335 -9607
rect 14111 -9701 14120 -9667
rect 14154 -9701 14163 -9667
rect 14111 -9752 14163 -9701
rect 14197 -9687 14249 -9641
rect 14197 -9721 14206 -9687
rect 14240 -9721 14249 -9687
rect 14197 -9786 14249 -9721
rect 14283 -9667 14335 -9615
rect 14455 -9615 14464 -9607
rect 14498 -9607 14636 -9581
rect 14498 -9615 14507 -9607
rect 14283 -9701 14292 -9667
rect 14326 -9701 14335 -9667
rect 14283 -9752 14335 -9701
rect 14369 -9687 14421 -9641
rect 14369 -9721 14378 -9687
rect 14412 -9721 14421 -9687
rect 14369 -9786 14421 -9721
rect 14455 -9667 14507 -9615
rect 14627 -9615 14636 -9607
rect 14670 -9607 14807 -9581
rect 14670 -9615 14679 -9607
rect 14455 -9701 14464 -9667
rect 14498 -9701 14507 -9667
rect 14455 -9752 14507 -9701
rect 14541 -9687 14593 -9641
rect 14541 -9721 14550 -9687
rect 14584 -9721 14593 -9687
rect 14541 -9786 14593 -9721
rect 14627 -9667 14679 -9615
rect 14796 -9615 14807 -9607
rect 14841 -9607 14979 -9581
rect 14841 -9615 14848 -9607
rect 14627 -9701 14636 -9667
rect 14670 -9701 14679 -9667
rect 14627 -9752 14679 -9701
rect 14713 -9687 14762 -9641
rect 14713 -9721 14722 -9687
rect 14756 -9721 14762 -9687
rect 14713 -9786 14762 -9721
rect 14796 -9667 14848 -9615
rect 14968 -9615 14979 -9607
rect 15013 -9607 15151 -9581
rect 15013 -9615 15020 -9607
rect 14796 -9701 14807 -9667
rect 14841 -9701 14848 -9667
rect 14796 -9752 14848 -9701
rect 14885 -9687 14934 -9641
rect 14885 -9721 14893 -9687
rect 14927 -9721 14934 -9687
rect 14885 -9786 14934 -9721
rect 14968 -9667 15020 -9615
rect 15140 -9615 15151 -9607
rect 15185 -9604 15323 -9581
rect 15185 -9615 15192 -9604
rect 14968 -9701 14979 -9667
rect 15013 -9701 15020 -9667
rect 14968 -9752 15020 -9701
rect 15057 -9687 15106 -9641
rect 15057 -9721 15065 -9687
rect 15099 -9721 15106 -9687
rect 15057 -9786 15106 -9721
rect 15140 -9667 15192 -9615
rect 15314 -9615 15323 -9604
rect 15357 -9604 15460 -9581
rect 15512 -9589 15570 -9554
rect 15357 -9615 15372 -9604
rect 15140 -9701 15151 -9667
rect 15185 -9701 15192 -9667
rect 15140 -9752 15192 -9701
rect 15229 -9687 15280 -9641
rect 15229 -9721 15237 -9687
rect 15271 -9721 15280 -9687
rect 15229 -9786 15280 -9721
rect 15314 -9667 15372 -9615
rect 15512 -9623 15524 -9589
rect 15558 -9623 15570 -9589
rect 15314 -9701 15323 -9667
rect 15357 -9701 15372 -9667
rect 15314 -9752 15372 -9701
rect 15406 -9687 15460 -9638
rect 15406 -9721 15409 -9687
rect 15443 -9721 15460 -9687
rect 14025 -9787 15280 -9786
rect 15406 -9787 15460 -9721
rect 15512 -9682 15570 -9623
rect 15512 -9716 15524 -9682
rect 15558 -9716 15570 -9682
rect 15512 -9787 15570 -9716
rect 15605 -9569 16124 -9499
rect 16158 -9501 16674 -9431
rect 16158 -9535 16178 -9501
rect 16212 -9535 16306 -9501
rect 16340 -9535 16434 -9501
rect 16468 -9535 16562 -9501
rect 16596 -9535 16674 -9501
rect 15605 -9609 16674 -9569
rect 15605 -9643 15622 -9609
rect 15656 -9643 16622 -9609
rect 16656 -9643 16674 -9609
rect 15605 -9711 16674 -9643
rect 15605 -9745 15622 -9711
rect 15656 -9745 16622 -9711
rect 16656 -9745 16674 -9711
rect 15605 -9787 16674 -9745
rect -2997 -9821 -2968 -9787
rect -2934 -9821 -2876 -9787
rect -2842 -9821 -2784 -9787
rect -2750 -9821 -2692 -9787
rect -2658 -9821 -2600 -9787
rect -2566 -9821 -2508 -9787
rect -2474 -9821 -2416 -9787
rect -2382 -9821 -2324 -9787
rect -2290 -9821 -2232 -9787
rect -2198 -9821 -2140 -9787
rect -2106 -9821 -2048 -9787
rect -2014 -9821 -1956 -9787
rect -1922 -9821 -1864 -9787
rect -1830 -9821 -1772 -9787
rect -1738 -9821 -1680 -9787
rect -1646 -9821 -1588 -9787
rect -1554 -9821 -1496 -9787
rect -1462 -9821 -1404 -9787
rect -1370 -9821 -1312 -9787
rect -1278 -9821 -1220 -9787
rect -1186 -9821 -1128 -9787
rect -1094 -9821 -1036 -9787
rect -1002 -9821 -944 -9787
rect -910 -9821 -852 -9787
rect -818 -9821 -760 -9787
rect -726 -9821 -668 -9787
rect -634 -9821 -576 -9787
rect -542 -9821 -484 -9787
rect -450 -9821 -392 -9787
rect -358 -9821 -300 -9787
rect -266 -9821 -208 -9787
rect -174 -9821 -116 -9787
rect -82 -9821 -24 -9787
rect 10 -9821 68 -9787
rect 102 -9821 160 -9787
rect 194 -9821 252 -9787
rect 286 -9821 344 -9787
rect 378 -9821 436 -9787
rect 470 -9821 528 -9787
rect 562 -9821 620 -9787
rect 654 -9821 712 -9787
rect 746 -9821 804 -9787
rect 838 -9821 896 -9787
rect 930 -9821 988 -9787
rect 1022 -9821 1080 -9787
rect 1114 -9821 1172 -9787
rect 1206 -9821 1264 -9787
rect 1298 -9821 1356 -9787
rect 1390 -9821 1448 -9787
rect 1482 -9821 1540 -9787
rect 1574 -9821 1632 -9787
rect 1666 -9821 1724 -9787
rect 1758 -9821 1816 -9787
rect 1850 -9821 1908 -9787
rect 1942 -9821 2000 -9787
rect 2034 -9821 2092 -9787
rect 2126 -9821 2184 -9787
rect 2218 -9821 2276 -9787
rect 2310 -9821 2368 -9787
rect 2402 -9821 2460 -9787
rect 2494 -9821 2552 -9787
rect 2586 -9821 2644 -9787
rect 2678 -9821 2736 -9787
rect 2770 -9821 2828 -9787
rect 2862 -9821 2920 -9787
rect 2954 -9821 3012 -9787
rect 3046 -9821 3104 -9787
rect 3138 -9821 3196 -9787
rect 3230 -9821 3288 -9787
rect 3322 -9821 3380 -9787
rect 3414 -9821 3472 -9787
rect 3506 -9821 3564 -9787
rect 3598 -9821 3656 -9787
rect 3690 -9821 3748 -9787
rect 3782 -9821 3840 -9787
rect 3874 -9821 3932 -9787
rect 3966 -9821 4024 -9787
rect 4058 -9821 4116 -9787
rect 4150 -9821 4208 -9787
rect 4242 -9821 4300 -9787
rect 4334 -9821 4392 -9787
rect 4426 -9821 4484 -9787
rect 4518 -9821 4576 -9787
rect 4610 -9821 4668 -9787
rect 4702 -9821 4760 -9787
rect 4794 -9821 4852 -9787
rect 4886 -9821 4944 -9787
rect 4978 -9821 5036 -9787
rect 5070 -9821 5128 -9787
rect 5162 -9821 5220 -9787
rect 5254 -9821 5312 -9787
rect 5346 -9821 5404 -9787
rect 5438 -9821 5496 -9787
rect 5530 -9821 5588 -9787
rect 5622 -9821 5680 -9787
rect 5714 -9821 5772 -9787
rect 5806 -9821 5864 -9787
rect 5898 -9821 5956 -9787
rect 5990 -9821 6048 -9787
rect 6082 -9821 6140 -9787
rect 6174 -9821 6232 -9787
rect 6266 -9821 6324 -9787
rect 6358 -9821 6416 -9787
rect 6450 -9821 6508 -9787
rect 6542 -9821 6600 -9787
rect 6634 -9821 6692 -9787
rect 6726 -9821 6784 -9787
rect 6818 -9821 6876 -9787
rect 6910 -9821 6968 -9787
rect 7002 -9821 7060 -9787
rect 7094 -9821 7152 -9787
rect 7186 -9821 7244 -9787
rect 7278 -9821 7336 -9787
rect 7370 -9821 7428 -9787
rect 7462 -9821 7520 -9787
rect 7554 -9821 7612 -9787
rect 7646 -9821 7704 -9787
rect 7738 -9821 7796 -9787
rect 7830 -9821 7888 -9787
rect 7922 -9821 7980 -9787
rect 8014 -9821 8072 -9787
rect 8106 -9821 8164 -9787
rect 8198 -9821 8256 -9787
rect 8290 -9821 8348 -9787
rect 8382 -9821 8440 -9787
rect 8474 -9821 8532 -9787
rect 8566 -9821 8624 -9787
rect 8658 -9821 8716 -9787
rect 8750 -9821 8808 -9787
rect 8842 -9821 8900 -9787
rect 8934 -9821 8992 -9787
rect 9026 -9821 9084 -9787
rect 9118 -9821 9176 -9787
rect 9210 -9821 9268 -9787
rect 9302 -9821 9360 -9787
rect 9394 -9821 9452 -9787
rect 9486 -9821 9544 -9787
rect 9578 -9821 9636 -9787
rect 9670 -9821 9728 -9787
rect 9762 -9821 9820 -9787
rect 9854 -9821 9912 -9787
rect 9946 -9821 10004 -9787
rect 10038 -9821 10096 -9787
rect 10130 -9821 10188 -9787
rect 10222 -9821 10280 -9787
rect 10314 -9821 10372 -9787
rect 10406 -9821 10464 -9787
rect 10498 -9821 10556 -9787
rect 10590 -9821 10648 -9787
rect 10682 -9821 10740 -9787
rect 10774 -9821 10832 -9787
rect 10866 -9821 10924 -9787
rect 10958 -9821 11016 -9787
rect 11050 -9821 11108 -9787
rect 11142 -9821 11200 -9787
rect 11234 -9821 11292 -9787
rect 11326 -9821 11384 -9787
rect 11418 -9821 11476 -9787
rect 11510 -9821 11568 -9787
rect 11602 -9821 11660 -9787
rect 11694 -9821 11752 -9787
rect 11786 -9821 11844 -9787
rect 11878 -9821 11936 -9787
rect 11970 -9821 12028 -9787
rect 12062 -9821 12120 -9787
rect 12154 -9821 12212 -9787
rect 12246 -9821 12304 -9787
rect 12338 -9821 12396 -9787
rect 12430 -9821 12488 -9787
rect 12522 -9821 12580 -9787
rect 12614 -9821 12672 -9787
rect 12706 -9821 12764 -9787
rect 12798 -9821 12856 -9787
rect 12890 -9821 12948 -9787
rect 12982 -9821 13040 -9787
rect 13074 -9821 13132 -9787
rect 13166 -9821 13224 -9787
rect 13258 -9821 13316 -9787
rect 13350 -9821 13408 -9787
rect 13442 -9821 13500 -9787
rect 13534 -9821 13592 -9787
rect 13626 -9821 13684 -9787
rect 13718 -9821 13776 -9787
rect 13810 -9821 13868 -9787
rect 13902 -9821 13960 -9787
rect 13994 -9821 14052 -9787
rect 14086 -9821 14144 -9787
rect 14178 -9821 14236 -9787
rect 14270 -9821 14328 -9787
rect 14362 -9821 14420 -9787
rect 14454 -9821 14512 -9787
rect 14546 -9821 14604 -9787
rect 14638 -9821 14696 -9787
rect 14730 -9821 14788 -9787
rect 14822 -9821 14880 -9787
rect 14914 -9821 14972 -9787
rect 15006 -9821 15064 -9787
rect 15098 -9821 15156 -9787
rect 15190 -9821 15248 -9787
rect 15282 -9821 15340 -9787
rect 15374 -9821 15432 -9787
rect 15466 -9821 15524 -9787
rect 15558 -9821 15616 -9787
rect 15650 -9821 15708 -9787
rect 15742 -9821 15800 -9787
rect 15834 -9821 15892 -9787
rect 15926 -9821 15984 -9787
rect 16018 -9821 16076 -9787
rect 16110 -9821 16168 -9787
rect 16202 -9821 16260 -9787
rect 16294 -9821 16352 -9787
rect 16386 -9821 16444 -9787
rect 16478 -9821 16536 -9787
rect 16570 -9821 16628 -9787
rect 16662 -9821 16691 -9787
rect -2980 -9863 -2278 -9821
rect -2980 -9897 -2962 -9863
rect -2928 -9897 -2330 -9863
rect -2296 -9897 -2278 -9863
rect -2980 -9965 -2278 -9897
rect -2980 -9999 -2962 -9965
rect -2928 -9999 -2330 -9965
rect -2296 -9999 -2278 -9965
rect -2980 -10039 -2278 -9999
rect -2980 -10107 -2902 -10073
rect -2868 -10107 -2803 -10073
rect -2769 -10107 -2704 -10073
rect -2670 -10107 -2650 -10073
rect -2980 -10177 -2650 -10107
rect -2616 -10109 -2278 -10039
rect -2244 -9892 -2186 -9821
rect -2244 -9926 -2232 -9892
rect -2198 -9926 -2186 -9892
rect -2244 -9985 -2186 -9926
rect -2244 -10019 -2232 -9985
rect -2198 -10019 -2186 -9985
rect -2244 -10054 -2186 -10019
rect -1600 -9863 -898 -9821
rect -1600 -9897 -1582 -9863
rect -1548 -9897 -950 -9863
rect -916 -9897 -898 -9863
rect -1600 -9965 -898 -9897
rect -1600 -9999 -1582 -9965
rect -1548 -9999 -950 -9965
rect -916 -9999 -898 -9965
rect -1600 -10039 -898 -9999
rect -864 -9863 -162 -9821
rect -864 -9897 -846 -9863
rect -812 -9897 -214 -9863
rect -180 -9897 -162 -9863
rect -864 -9965 -162 -9897
rect -864 -9999 -846 -9965
rect -812 -9999 -214 -9965
rect -180 -9999 -162 -9965
rect -864 -10039 -162 -9999
rect -2616 -10143 -2596 -10109
rect -2562 -10143 -2493 -10109
rect -2459 -10143 -2390 -10109
rect -2356 -10143 -2278 -10109
rect -1600 -10107 -1522 -10073
rect -1488 -10107 -1423 -10073
rect -1389 -10107 -1324 -10073
rect -1290 -10107 -1270 -10073
rect -1600 -10177 -1270 -10107
rect -1236 -10109 -898 -10039
rect -1236 -10143 -1216 -10109
rect -1182 -10143 -1113 -10109
rect -1079 -10143 -1010 -10109
rect -976 -10143 -898 -10109
rect -864 -10107 -786 -10073
rect -752 -10107 -687 -10073
rect -653 -10107 -588 -10073
rect -554 -10107 -534 -10073
rect -864 -10177 -534 -10107
rect -500 -10109 -162 -10039
rect -128 -9892 -70 -9821
rect -128 -9926 -116 -9892
rect -82 -9926 -70 -9892
rect -128 -9985 -70 -9926
rect -128 -10019 -116 -9985
rect -82 -10019 -70 -9985
rect -128 -10054 -70 -10019
rect -36 -9863 298 -9821
rect -36 -9897 -18 -9863
rect 16 -9897 246 -9863
rect 280 -9897 298 -9863
rect -36 -9965 298 -9897
rect -36 -9999 -18 -9965
rect 16 -9999 246 -9965
rect 280 -9999 298 -9965
rect -36 -10039 298 -9999
rect 332 -9892 390 -9821
rect 332 -9926 344 -9892
rect 378 -9926 390 -9892
rect 332 -9985 390 -9926
rect 332 -10019 344 -9985
rect 378 -10019 390 -9985
rect -500 -10143 -480 -10109
rect -446 -10143 -377 -10109
rect -343 -10143 -274 -10109
rect -240 -10143 -162 -10109
rect -36 -10109 114 -10039
rect 332 -10054 390 -10019
rect 424 -9870 493 -9855
rect 424 -9904 443 -9870
rect 477 -9904 493 -9870
rect 424 -9938 493 -9904
rect 424 -9972 443 -9938
rect 477 -9972 493 -9938
rect 424 -10022 493 -9972
rect 527 -9870 593 -9821
rect 527 -9904 543 -9870
rect 577 -9904 593 -9870
rect 527 -9938 593 -9904
rect 527 -9972 543 -9938
rect 577 -9972 593 -9938
rect 527 -9988 593 -9972
rect 683 -9870 753 -9855
rect 683 -9904 701 -9870
rect 735 -9904 753 -9870
rect 683 -9938 753 -9904
rect 683 -9972 701 -9938
rect 735 -9972 753 -9938
rect 424 -10056 618 -10022
rect -36 -10143 -16 -10109
rect 18 -10143 114 -10109
rect 148 -10107 244 -10073
rect 278 -10107 298 -10073
rect 548 -10085 618 -10056
rect 683 -10084 753 -9972
rect 805 -9871 855 -9855
rect 839 -9905 855 -9871
rect 805 -9939 855 -9905
rect 839 -9973 855 -9939
rect 805 -10015 855 -9973
rect 945 -9870 1011 -9821
rect 945 -9904 961 -9870
rect 995 -9904 1011 -9870
rect 945 -9938 1011 -9904
rect 945 -9972 961 -9938
rect 995 -9972 1011 -9938
rect 945 -9981 1011 -9972
rect 1045 -9871 1126 -9855
rect 1045 -9905 1059 -9871
rect 1093 -9905 1126 -9871
rect 1045 -9939 1126 -9905
rect 1045 -9973 1059 -9939
rect 1093 -9973 1126 -9939
rect 1045 -10010 1126 -9973
rect 805 -10049 923 -10015
rect 889 -10083 923 -10049
rect 148 -10177 298 -10107
rect 424 -10096 514 -10090
rect 424 -10130 436 -10096
rect 470 -10099 514 -10096
rect 424 -10133 464 -10130
rect 498 -10133 514 -10099
rect 548 -10099 634 -10085
rect 548 -10133 584 -10099
rect 618 -10133 634 -10099
rect 548 -10143 634 -10133
rect 683 -10099 855 -10084
rect 683 -10133 805 -10099
rect 839 -10133 855 -10099
rect 683 -10134 855 -10133
rect 889 -10099 1042 -10083
rect 889 -10133 1005 -10099
rect 1039 -10133 1042 -10099
rect 548 -10167 618 -10143
rect -2980 -10236 -2278 -10177
rect -2980 -10270 -2962 -10236
rect -2928 -10270 -2330 -10236
rect -2296 -10270 -2278 -10236
rect -2980 -10331 -2278 -10270
rect -2244 -10203 -2186 -10186
rect -2244 -10237 -2232 -10203
rect -2198 -10237 -2186 -10203
rect -2244 -10331 -2186 -10237
rect -1600 -10236 -898 -10177
rect -1600 -10270 -1582 -10236
rect -1548 -10270 -950 -10236
rect -916 -10270 -898 -10236
rect -1600 -10331 -898 -10270
rect -864 -10236 -162 -10177
rect -864 -10270 -846 -10236
rect -812 -10270 -214 -10236
rect -180 -10270 -162 -10236
rect -864 -10331 -162 -10270
rect -128 -10203 -70 -10186
rect -128 -10237 -116 -10203
rect -82 -10237 -70 -10203
rect -128 -10331 -70 -10237
rect -36 -10229 298 -10177
rect -36 -10263 -18 -10229
rect 16 -10263 246 -10229
rect 280 -10263 298 -10229
rect -36 -10331 298 -10263
rect 332 -10203 390 -10186
rect 332 -10237 344 -10203
rect 378 -10237 390 -10203
rect 332 -10331 390 -10237
rect 424 -10201 618 -10167
rect 424 -10244 490 -10201
rect 424 -10278 443 -10244
rect 477 -10278 490 -10244
rect 424 -10297 490 -10278
rect 524 -10244 590 -10235
rect 524 -10278 540 -10244
rect 574 -10278 590 -10244
rect 524 -10331 590 -10278
rect 683 -10244 753 -10134
rect 889 -10149 1042 -10133
rect 1076 -10094 1126 -10010
rect 1160 -9892 1218 -9821
rect 1160 -9926 1172 -9892
rect 1206 -9926 1218 -9892
rect 1160 -9985 1218 -9926
rect 1160 -10019 1172 -9985
rect 1206 -10019 1218 -9985
rect 1160 -10054 1218 -10019
rect 1252 -9863 1586 -9821
rect 1252 -9897 1270 -9863
rect 1304 -9897 1534 -9863
rect 1568 -9897 1586 -9863
rect 1252 -9965 1586 -9897
rect 1252 -9999 1270 -9965
rect 1304 -9999 1534 -9965
rect 1568 -9999 1586 -9965
rect 1252 -10039 1586 -9999
rect 1620 -9892 1678 -9821
rect 1620 -9926 1632 -9892
rect 1666 -9926 1678 -9892
rect 1620 -9985 1678 -9926
rect 1620 -10019 1632 -9985
rect 1666 -10019 1678 -9985
rect 1076 -10128 1081 -10094
rect 1115 -10128 1126 -10094
rect 889 -10168 923 -10149
rect 683 -10278 700 -10244
rect 734 -10278 753 -10244
rect 683 -10297 753 -10278
rect 805 -10202 923 -10168
rect 805 -10244 855 -10202
rect 1076 -10220 1126 -10128
rect 1252 -10109 1402 -10039
rect 1620 -10054 1678 -10019
rect 1712 -9863 2414 -9821
rect 1712 -9897 1730 -9863
rect 1764 -9897 2362 -9863
rect 2396 -9897 2414 -9863
rect 1712 -9965 2414 -9897
rect 1712 -9999 1730 -9965
rect 1764 -9999 2362 -9965
rect 2396 -9999 2414 -9965
rect 1712 -10039 2414 -9999
rect 1252 -10143 1272 -10109
rect 1306 -10143 1402 -10109
rect 1436 -10107 1532 -10073
rect 1566 -10107 1586 -10073
rect 1436 -10177 1586 -10107
rect 839 -10278 855 -10244
rect 805 -10297 855 -10278
rect 945 -10244 1011 -10228
rect 945 -10278 961 -10244
rect 995 -10278 1011 -10244
rect 945 -10331 1011 -10278
rect 1045 -10244 1126 -10220
rect 1045 -10278 1059 -10244
rect 1093 -10278 1126 -10244
rect 1045 -10297 1126 -10278
rect 1160 -10203 1218 -10186
rect 1160 -10237 1172 -10203
rect 1206 -10237 1218 -10203
rect 1160 -10331 1218 -10237
rect 1252 -10229 1586 -10177
rect 1712 -10107 1790 -10073
rect 1824 -10107 1889 -10073
rect 1923 -10107 1988 -10073
rect 2022 -10107 2042 -10073
rect 1712 -10177 2042 -10107
rect 2076 -10109 2414 -10039
rect 2448 -9892 2506 -9821
rect 2448 -9926 2460 -9892
rect 2494 -9926 2506 -9892
rect 2448 -9985 2506 -9926
rect 2448 -10019 2460 -9985
rect 2494 -10019 2506 -9985
rect 2448 -10054 2506 -10019
rect 2540 -9863 2874 -9821
rect 2540 -9897 2558 -9863
rect 2592 -9897 2822 -9863
rect 2856 -9897 2874 -9863
rect 2540 -9965 2874 -9897
rect 2540 -9999 2558 -9965
rect 2592 -9999 2822 -9965
rect 2856 -9999 2874 -9965
rect 2540 -10039 2874 -9999
rect 2908 -9892 2966 -9821
rect 2908 -9926 2920 -9892
rect 2954 -9926 2966 -9892
rect 2908 -9985 2966 -9926
rect 2908 -10019 2920 -9985
rect 2954 -10019 2966 -9985
rect 2076 -10143 2096 -10109
rect 2130 -10143 2199 -10109
rect 2233 -10143 2302 -10109
rect 2336 -10143 2414 -10109
rect 2540 -10109 2690 -10039
rect 2908 -10054 2966 -10019
rect 3000 -9870 3069 -9855
rect 3000 -9904 3019 -9870
rect 3053 -9904 3069 -9870
rect 3000 -9938 3069 -9904
rect 3000 -9972 3019 -9938
rect 3053 -9972 3069 -9938
rect 3000 -10022 3069 -9972
rect 3103 -9870 3169 -9821
rect 3103 -9904 3119 -9870
rect 3153 -9904 3169 -9870
rect 3103 -9938 3169 -9904
rect 3103 -9972 3119 -9938
rect 3153 -9972 3169 -9938
rect 3103 -9988 3169 -9972
rect 3259 -9870 3329 -9855
rect 3259 -9904 3277 -9870
rect 3311 -9904 3329 -9870
rect 3259 -9938 3329 -9904
rect 3259 -9972 3277 -9938
rect 3311 -9972 3329 -9938
rect 3000 -10056 3194 -10022
rect 2540 -10143 2560 -10109
rect 2594 -10143 2690 -10109
rect 2724 -10107 2820 -10073
rect 2854 -10107 2874 -10073
rect 3124 -10085 3194 -10056
rect 3259 -10084 3329 -9972
rect 3381 -9871 3431 -9855
rect 3415 -9905 3431 -9871
rect 3381 -9939 3431 -9905
rect 3415 -9973 3431 -9939
rect 3381 -10015 3431 -9973
rect 3521 -9870 3587 -9821
rect 3521 -9904 3537 -9870
rect 3571 -9904 3587 -9870
rect 3521 -9938 3587 -9904
rect 3521 -9972 3537 -9938
rect 3571 -9972 3587 -9938
rect 3521 -9981 3587 -9972
rect 3621 -9871 3702 -9855
rect 3621 -9905 3635 -9871
rect 3669 -9905 3702 -9871
rect 3621 -9939 3702 -9905
rect 3621 -9973 3635 -9939
rect 3669 -9973 3702 -9939
rect 3621 -10010 3702 -9973
rect 3381 -10049 3499 -10015
rect 3465 -10083 3499 -10049
rect 2724 -10177 2874 -10107
rect 3000 -10094 3090 -10090
rect 3000 -10099 3041 -10094
rect 3000 -10133 3040 -10099
rect 3075 -10128 3090 -10094
rect 3074 -10133 3090 -10128
rect 3124 -10099 3210 -10085
rect 3124 -10133 3160 -10099
rect 3194 -10133 3210 -10099
rect 3124 -10143 3210 -10133
rect 3259 -10099 3431 -10084
rect 3259 -10133 3381 -10099
rect 3415 -10133 3431 -10099
rect 3259 -10134 3431 -10133
rect 3465 -10099 3618 -10083
rect 3465 -10133 3581 -10099
rect 3615 -10133 3618 -10099
rect 3124 -10167 3194 -10143
rect 1252 -10263 1270 -10229
rect 1304 -10263 1534 -10229
rect 1568 -10263 1586 -10229
rect 1252 -10331 1586 -10263
rect 1620 -10203 1678 -10186
rect 1620 -10237 1632 -10203
rect 1666 -10237 1678 -10203
rect 1620 -10331 1678 -10237
rect 1712 -10236 2414 -10177
rect 1712 -10270 1730 -10236
rect 1764 -10270 2362 -10236
rect 2396 -10270 2414 -10236
rect 1712 -10331 2414 -10270
rect 2448 -10203 2506 -10186
rect 2448 -10237 2460 -10203
rect 2494 -10237 2506 -10203
rect 2448 -10331 2506 -10237
rect 2540 -10229 2874 -10177
rect 2540 -10263 2558 -10229
rect 2592 -10263 2822 -10229
rect 2856 -10263 2874 -10229
rect 2540 -10331 2874 -10263
rect 2908 -10203 2966 -10186
rect 2908 -10237 2920 -10203
rect 2954 -10237 2966 -10203
rect 2908 -10331 2966 -10237
rect 3000 -10201 3194 -10167
rect 3000 -10244 3066 -10201
rect 3000 -10278 3019 -10244
rect 3053 -10278 3066 -10244
rect 3000 -10297 3066 -10278
rect 3100 -10244 3166 -10235
rect 3100 -10278 3116 -10244
rect 3150 -10278 3166 -10244
rect 3100 -10331 3166 -10278
rect 3259 -10244 3329 -10134
rect 3465 -10149 3618 -10133
rect 3652 -10094 3702 -10010
rect 3736 -9892 3794 -9821
rect 3736 -9926 3748 -9892
rect 3782 -9926 3794 -9892
rect 3736 -9985 3794 -9926
rect 3736 -10019 3748 -9985
rect 3782 -10019 3794 -9985
rect 3736 -10054 3794 -10019
rect 3828 -9863 4162 -9821
rect 3828 -9897 3846 -9863
rect 3880 -9897 4110 -9863
rect 4144 -9897 4162 -9863
rect 3828 -9965 4162 -9897
rect 3828 -9999 3846 -9965
rect 3880 -9999 4110 -9965
rect 4144 -9999 4162 -9965
rect 3828 -10039 4162 -9999
rect 4196 -9892 4254 -9821
rect 4196 -9926 4208 -9892
rect 4242 -9926 4254 -9892
rect 4196 -9985 4254 -9926
rect 4196 -10019 4208 -9985
rect 4242 -10019 4254 -9985
rect 3652 -10128 3655 -10094
rect 3689 -10128 3702 -10094
rect 3465 -10168 3499 -10149
rect 3259 -10278 3276 -10244
rect 3310 -10278 3329 -10244
rect 3259 -10297 3329 -10278
rect 3381 -10202 3499 -10168
rect 3381 -10244 3431 -10202
rect 3652 -10220 3702 -10128
rect 3828 -10109 3978 -10039
rect 4196 -10054 4254 -10019
rect 4288 -9863 4990 -9821
rect 4288 -9897 4306 -9863
rect 4340 -9897 4938 -9863
rect 4972 -9897 4990 -9863
rect 4288 -9965 4990 -9897
rect 4288 -9999 4306 -9965
rect 4340 -9999 4938 -9965
rect 4972 -9999 4990 -9965
rect 4288 -10039 4990 -9999
rect 3828 -10143 3848 -10109
rect 3882 -10143 3978 -10109
rect 4012 -10107 4108 -10073
rect 4142 -10107 4162 -10073
rect 4012 -10177 4162 -10107
rect 3415 -10278 3431 -10244
rect 3381 -10297 3431 -10278
rect 3521 -10244 3587 -10228
rect 3521 -10278 3537 -10244
rect 3571 -10278 3587 -10244
rect 3521 -10331 3587 -10278
rect 3621 -10244 3702 -10220
rect 3621 -10278 3635 -10244
rect 3669 -10278 3702 -10244
rect 3621 -10297 3702 -10278
rect 3736 -10203 3794 -10186
rect 3736 -10237 3748 -10203
rect 3782 -10237 3794 -10203
rect 3736 -10331 3794 -10237
rect 3828 -10229 4162 -10177
rect 4288 -10107 4366 -10073
rect 4400 -10107 4465 -10073
rect 4499 -10107 4564 -10073
rect 4598 -10107 4618 -10073
rect 4288 -10177 4618 -10107
rect 4652 -10109 4990 -10039
rect 5024 -9892 5082 -9821
rect 5024 -9926 5036 -9892
rect 5070 -9926 5082 -9892
rect 5024 -9985 5082 -9926
rect 5024 -10019 5036 -9985
rect 5070 -10019 5082 -9985
rect 5024 -10054 5082 -10019
rect 5116 -9863 5450 -9821
rect 5116 -9897 5134 -9863
rect 5168 -9897 5398 -9863
rect 5432 -9897 5450 -9863
rect 5116 -9965 5450 -9897
rect 5116 -9999 5134 -9965
rect 5168 -9999 5398 -9965
rect 5432 -9999 5450 -9965
rect 5116 -10039 5450 -9999
rect 5484 -9892 5542 -9821
rect 5484 -9926 5496 -9892
rect 5530 -9926 5542 -9892
rect 5484 -9985 5542 -9926
rect 5484 -10019 5496 -9985
rect 5530 -10019 5542 -9985
rect 4652 -10143 4672 -10109
rect 4706 -10143 4775 -10109
rect 4809 -10143 4878 -10109
rect 4912 -10143 4990 -10109
rect 5116 -10109 5266 -10039
rect 5484 -10054 5542 -10019
rect 5576 -9870 5645 -9855
rect 5576 -9904 5595 -9870
rect 5629 -9904 5645 -9870
rect 5576 -9938 5645 -9904
rect 5576 -9972 5595 -9938
rect 5629 -9972 5645 -9938
rect 5576 -10022 5645 -9972
rect 5679 -9870 5745 -9821
rect 5679 -9904 5695 -9870
rect 5729 -9904 5745 -9870
rect 5679 -9938 5745 -9904
rect 5679 -9972 5695 -9938
rect 5729 -9972 5745 -9938
rect 5679 -9988 5745 -9972
rect 5835 -9870 5905 -9855
rect 5835 -9904 5853 -9870
rect 5887 -9904 5905 -9870
rect 5835 -9938 5905 -9904
rect 5835 -9972 5853 -9938
rect 5887 -9972 5905 -9938
rect 5576 -10056 5770 -10022
rect 5116 -10143 5136 -10109
rect 5170 -10143 5266 -10109
rect 5300 -10107 5396 -10073
rect 5430 -10107 5450 -10073
rect 5700 -10085 5770 -10056
rect 5835 -10084 5905 -9972
rect 5957 -9871 6007 -9855
rect 5991 -9905 6007 -9871
rect 5957 -9939 6007 -9905
rect 5991 -9973 6007 -9939
rect 5957 -10015 6007 -9973
rect 6097 -9870 6163 -9821
rect 6097 -9904 6113 -9870
rect 6147 -9904 6163 -9870
rect 6097 -9938 6163 -9904
rect 6097 -9972 6113 -9938
rect 6147 -9972 6163 -9938
rect 6097 -9981 6163 -9972
rect 6197 -9871 6278 -9855
rect 6197 -9905 6211 -9871
rect 6245 -9905 6278 -9871
rect 6197 -9939 6278 -9905
rect 6197 -9973 6211 -9939
rect 6245 -9973 6278 -9939
rect 6197 -10010 6278 -9973
rect 5957 -10049 6075 -10015
rect 6041 -10083 6075 -10049
rect 5300 -10177 5450 -10107
rect 5576 -10094 5666 -10090
rect 5576 -10128 5615 -10094
rect 5649 -10099 5666 -10094
rect 5576 -10133 5616 -10128
rect 5650 -10133 5666 -10099
rect 5700 -10099 5786 -10085
rect 5700 -10133 5736 -10099
rect 5770 -10133 5786 -10099
rect 5700 -10143 5786 -10133
rect 5835 -10099 6007 -10084
rect 5835 -10133 5957 -10099
rect 5991 -10133 6007 -10099
rect 5835 -10134 6007 -10133
rect 6041 -10099 6194 -10083
rect 6041 -10133 6157 -10099
rect 6191 -10133 6194 -10099
rect 5700 -10167 5770 -10143
rect 3828 -10263 3846 -10229
rect 3880 -10263 4110 -10229
rect 4144 -10263 4162 -10229
rect 3828 -10331 4162 -10263
rect 4196 -10203 4254 -10186
rect 4196 -10237 4208 -10203
rect 4242 -10237 4254 -10203
rect 4196 -10331 4254 -10237
rect 4288 -10236 4990 -10177
rect 4288 -10270 4306 -10236
rect 4340 -10270 4938 -10236
rect 4972 -10270 4990 -10236
rect 4288 -10331 4990 -10270
rect 5024 -10203 5082 -10186
rect 5024 -10237 5036 -10203
rect 5070 -10237 5082 -10203
rect 5024 -10331 5082 -10237
rect 5116 -10229 5450 -10177
rect 5116 -10263 5134 -10229
rect 5168 -10263 5398 -10229
rect 5432 -10263 5450 -10229
rect 5116 -10331 5450 -10263
rect 5484 -10203 5542 -10186
rect 5484 -10237 5496 -10203
rect 5530 -10237 5542 -10203
rect 5484 -10331 5542 -10237
rect 5576 -10201 5770 -10167
rect 5576 -10244 5642 -10201
rect 5576 -10278 5595 -10244
rect 5629 -10278 5642 -10244
rect 5576 -10297 5642 -10278
rect 5676 -10244 5742 -10235
rect 5676 -10278 5692 -10244
rect 5726 -10278 5742 -10244
rect 5676 -10331 5742 -10278
rect 5835 -10244 5905 -10134
rect 6041 -10149 6194 -10133
rect 6228 -10094 6278 -10010
rect 6312 -9892 6370 -9821
rect 6312 -9926 6324 -9892
rect 6358 -9926 6370 -9892
rect 6312 -9985 6370 -9926
rect 6312 -10019 6324 -9985
rect 6358 -10019 6370 -9985
rect 6312 -10054 6370 -10019
rect 6404 -9863 6738 -9821
rect 6404 -9897 6422 -9863
rect 6456 -9897 6686 -9863
rect 6720 -9897 6738 -9863
rect 6404 -9965 6738 -9897
rect 6404 -9999 6422 -9965
rect 6456 -9999 6686 -9965
rect 6720 -9999 6738 -9965
rect 6404 -10039 6738 -9999
rect 6772 -9892 6830 -9821
rect 6772 -9926 6784 -9892
rect 6818 -9926 6830 -9892
rect 6772 -9985 6830 -9926
rect 6772 -10019 6784 -9985
rect 6818 -10019 6830 -9985
rect 6228 -10128 6229 -10094
rect 6263 -10128 6278 -10094
rect 6041 -10168 6075 -10149
rect 5835 -10278 5852 -10244
rect 5886 -10278 5905 -10244
rect 5835 -10297 5905 -10278
rect 5957 -10202 6075 -10168
rect 5957 -10244 6007 -10202
rect 6228 -10220 6278 -10128
rect 6404 -10109 6554 -10039
rect 6772 -10054 6830 -10019
rect 6864 -9863 7566 -9821
rect 6864 -9897 6882 -9863
rect 6916 -9897 7514 -9863
rect 7548 -9897 7566 -9863
rect 6864 -9965 7566 -9897
rect 6864 -9999 6882 -9965
rect 6916 -9999 7514 -9965
rect 7548 -9999 7566 -9965
rect 6864 -10039 7566 -9999
rect 6404 -10143 6424 -10109
rect 6458 -10143 6554 -10109
rect 6588 -10107 6684 -10073
rect 6718 -10107 6738 -10073
rect 6588 -10177 6738 -10107
rect 5991 -10278 6007 -10244
rect 5957 -10297 6007 -10278
rect 6097 -10244 6163 -10228
rect 6097 -10278 6113 -10244
rect 6147 -10278 6163 -10244
rect 6097 -10331 6163 -10278
rect 6197 -10244 6278 -10220
rect 6197 -10278 6211 -10244
rect 6245 -10278 6278 -10244
rect 6197 -10297 6278 -10278
rect 6312 -10203 6370 -10186
rect 6312 -10237 6324 -10203
rect 6358 -10237 6370 -10203
rect 6312 -10331 6370 -10237
rect 6404 -10229 6738 -10177
rect 6864 -10107 6942 -10073
rect 6976 -10107 7041 -10073
rect 7075 -10107 7140 -10073
rect 7174 -10107 7194 -10073
rect 6864 -10177 7194 -10107
rect 7228 -10109 7566 -10039
rect 7600 -9892 7658 -9821
rect 7600 -9926 7612 -9892
rect 7646 -9926 7658 -9892
rect 7600 -9985 7658 -9926
rect 7600 -10019 7612 -9985
rect 7646 -10019 7658 -9985
rect 7600 -10054 7658 -10019
rect 7692 -9863 8026 -9821
rect 7692 -9897 7710 -9863
rect 7744 -9897 7974 -9863
rect 8008 -9897 8026 -9863
rect 7692 -9965 8026 -9897
rect 7692 -9999 7710 -9965
rect 7744 -9999 7974 -9965
rect 8008 -9999 8026 -9965
rect 7692 -10039 8026 -9999
rect 8060 -9892 8118 -9821
rect 8060 -9926 8072 -9892
rect 8106 -9926 8118 -9892
rect 8060 -9985 8118 -9926
rect 8060 -10019 8072 -9985
rect 8106 -10019 8118 -9985
rect 7228 -10143 7248 -10109
rect 7282 -10143 7351 -10109
rect 7385 -10143 7454 -10109
rect 7488 -10143 7566 -10109
rect 7692 -10109 7842 -10039
rect 8060 -10054 8118 -10019
rect 8152 -9870 8221 -9855
rect 8152 -9904 8171 -9870
rect 8205 -9904 8221 -9870
rect 8152 -9938 8221 -9904
rect 8152 -9972 8171 -9938
rect 8205 -9972 8221 -9938
rect 8152 -10022 8221 -9972
rect 8255 -9870 8321 -9821
rect 8255 -9904 8271 -9870
rect 8305 -9904 8321 -9870
rect 8255 -9938 8321 -9904
rect 8255 -9972 8271 -9938
rect 8305 -9972 8321 -9938
rect 8255 -9988 8321 -9972
rect 8411 -9870 8481 -9855
rect 8411 -9904 8429 -9870
rect 8463 -9904 8481 -9870
rect 8411 -9938 8481 -9904
rect 8411 -9972 8429 -9938
rect 8463 -9972 8481 -9938
rect 8152 -10056 8346 -10022
rect 7692 -10143 7712 -10109
rect 7746 -10143 7842 -10109
rect 7876 -10107 7972 -10073
rect 8006 -10107 8026 -10073
rect 8276 -10085 8346 -10056
rect 8411 -10084 8481 -9972
rect 8533 -9871 8583 -9855
rect 8567 -9905 8583 -9871
rect 8533 -9939 8583 -9905
rect 8567 -9973 8583 -9939
rect 8533 -10015 8583 -9973
rect 8673 -9870 8739 -9821
rect 8673 -9904 8689 -9870
rect 8723 -9904 8739 -9870
rect 8673 -9938 8739 -9904
rect 8673 -9972 8689 -9938
rect 8723 -9972 8739 -9938
rect 8673 -9981 8739 -9972
rect 8773 -9871 8854 -9855
rect 8773 -9905 8787 -9871
rect 8821 -9905 8854 -9871
rect 8773 -9939 8854 -9905
rect 8773 -9973 8787 -9939
rect 8821 -9973 8854 -9939
rect 8773 -10010 8854 -9973
rect 8533 -10049 8651 -10015
rect 8617 -10083 8651 -10049
rect 7876 -10177 8026 -10107
rect 8152 -10094 8242 -10090
rect 8152 -10128 8189 -10094
rect 8223 -10099 8242 -10094
rect 8152 -10133 8192 -10128
rect 8226 -10133 8242 -10099
rect 8276 -10099 8362 -10085
rect 8276 -10133 8312 -10099
rect 8346 -10133 8362 -10099
rect 8276 -10143 8362 -10133
rect 8411 -10099 8583 -10084
rect 8411 -10133 8533 -10099
rect 8567 -10133 8583 -10099
rect 8411 -10134 8583 -10133
rect 8617 -10099 8770 -10083
rect 8617 -10133 8733 -10099
rect 8767 -10133 8770 -10099
rect 8276 -10167 8346 -10143
rect 6404 -10263 6422 -10229
rect 6456 -10263 6686 -10229
rect 6720 -10263 6738 -10229
rect 6404 -10331 6738 -10263
rect 6772 -10203 6830 -10186
rect 6772 -10237 6784 -10203
rect 6818 -10237 6830 -10203
rect 6772 -10331 6830 -10237
rect 6864 -10236 7566 -10177
rect 6864 -10270 6882 -10236
rect 6916 -10270 7514 -10236
rect 7548 -10270 7566 -10236
rect 6864 -10331 7566 -10270
rect 7600 -10203 7658 -10186
rect 7600 -10237 7612 -10203
rect 7646 -10237 7658 -10203
rect 7600 -10331 7658 -10237
rect 7692 -10229 8026 -10177
rect 7692 -10263 7710 -10229
rect 7744 -10263 7974 -10229
rect 8008 -10263 8026 -10229
rect 7692 -10331 8026 -10263
rect 8060 -10203 8118 -10186
rect 8060 -10237 8072 -10203
rect 8106 -10237 8118 -10203
rect 8060 -10331 8118 -10237
rect 8152 -10201 8346 -10167
rect 8152 -10244 8218 -10201
rect 8152 -10278 8171 -10244
rect 8205 -10278 8218 -10244
rect 8152 -10297 8218 -10278
rect 8252 -10244 8318 -10235
rect 8252 -10278 8268 -10244
rect 8302 -10278 8318 -10244
rect 8252 -10331 8318 -10278
rect 8411 -10244 8481 -10134
rect 8617 -10149 8770 -10133
rect 8804 -10094 8854 -10010
rect 8888 -9892 8946 -9821
rect 8888 -9926 8900 -9892
rect 8934 -9926 8946 -9892
rect 8888 -9985 8946 -9926
rect 8888 -10019 8900 -9985
rect 8934 -10019 8946 -9985
rect 8888 -10054 8946 -10019
rect 8980 -9863 9314 -9821
rect 8980 -9897 8998 -9863
rect 9032 -9897 9262 -9863
rect 9296 -9897 9314 -9863
rect 8980 -9965 9314 -9897
rect 8980 -9999 8998 -9965
rect 9032 -9999 9262 -9965
rect 9296 -9999 9314 -9965
rect 8980 -10039 9314 -9999
rect 9348 -9892 9406 -9821
rect 9348 -9926 9360 -9892
rect 9394 -9926 9406 -9892
rect 9348 -9985 9406 -9926
rect 9348 -10019 9360 -9985
rect 9394 -10019 9406 -9985
rect 8804 -10128 8806 -10094
rect 8840 -10128 8854 -10094
rect 8617 -10168 8651 -10149
rect 8411 -10278 8428 -10244
rect 8462 -10278 8481 -10244
rect 8411 -10297 8481 -10278
rect 8533 -10202 8651 -10168
rect 8533 -10244 8583 -10202
rect 8804 -10220 8854 -10128
rect 8980 -10109 9130 -10039
rect 9348 -10054 9406 -10019
rect 9440 -9863 10142 -9821
rect 9440 -9897 9458 -9863
rect 9492 -9897 10090 -9863
rect 10124 -9897 10142 -9863
rect 9440 -9965 10142 -9897
rect 9440 -9999 9458 -9965
rect 9492 -9999 10090 -9965
rect 10124 -9999 10142 -9965
rect 9440 -10039 10142 -9999
rect 8980 -10143 9000 -10109
rect 9034 -10143 9130 -10109
rect 9164 -10107 9260 -10073
rect 9294 -10107 9314 -10073
rect 9164 -10177 9314 -10107
rect 8567 -10278 8583 -10244
rect 8533 -10297 8583 -10278
rect 8673 -10244 8739 -10228
rect 8673 -10278 8689 -10244
rect 8723 -10278 8739 -10244
rect 8673 -10331 8739 -10278
rect 8773 -10244 8854 -10220
rect 8773 -10278 8787 -10244
rect 8821 -10278 8854 -10244
rect 8773 -10297 8854 -10278
rect 8888 -10203 8946 -10186
rect 8888 -10237 8900 -10203
rect 8934 -10237 8946 -10203
rect 8888 -10331 8946 -10237
rect 8980 -10229 9314 -10177
rect 9440 -10107 9518 -10073
rect 9552 -10107 9617 -10073
rect 9651 -10107 9716 -10073
rect 9750 -10107 9770 -10073
rect 9440 -10177 9770 -10107
rect 9804 -10109 10142 -10039
rect 10176 -9892 10234 -9821
rect 10176 -9926 10188 -9892
rect 10222 -9926 10234 -9892
rect 10176 -9985 10234 -9926
rect 10176 -10019 10188 -9985
rect 10222 -10019 10234 -9985
rect 10176 -10054 10234 -10019
rect 10360 -9863 10694 -9821
rect 10360 -9897 10378 -9863
rect 10412 -9897 10642 -9863
rect 10676 -9897 10694 -9863
rect 10360 -9965 10694 -9897
rect 10360 -9999 10378 -9965
rect 10412 -9999 10642 -9965
rect 10676 -9999 10694 -9965
rect 10360 -10039 10694 -9999
rect 10728 -9870 10797 -9855
rect 10728 -9904 10747 -9870
rect 10781 -9904 10797 -9870
rect 10728 -9938 10797 -9904
rect 10728 -9972 10747 -9938
rect 10781 -9972 10797 -9938
rect 10728 -10022 10797 -9972
rect 10831 -9870 10897 -9821
rect 10831 -9904 10847 -9870
rect 10881 -9904 10897 -9870
rect 10831 -9938 10897 -9904
rect 10831 -9972 10847 -9938
rect 10881 -9972 10897 -9938
rect 10831 -9988 10897 -9972
rect 10987 -9870 11057 -9855
rect 10987 -9904 11005 -9870
rect 11039 -9904 11057 -9870
rect 10987 -9938 11057 -9904
rect 10987 -9972 11005 -9938
rect 11039 -9972 11057 -9938
rect 9804 -10143 9824 -10109
rect 9858 -10143 9927 -10109
rect 9961 -10143 10030 -10109
rect 10064 -10143 10142 -10109
rect 10360 -10109 10510 -10039
rect 10728 -10056 10922 -10022
rect 10360 -10143 10380 -10109
rect 10414 -10143 10510 -10109
rect 10544 -10107 10640 -10073
rect 10674 -10107 10694 -10073
rect 10852 -10085 10922 -10056
rect 10987 -10084 11057 -9972
rect 11109 -9871 11159 -9855
rect 11143 -9905 11159 -9871
rect 11109 -9939 11159 -9905
rect 11143 -9973 11159 -9939
rect 11109 -10015 11159 -9973
rect 11249 -9870 11315 -9821
rect 11249 -9904 11265 -9870
rect 11299 -9904 11315 -9870
rect 11249 -9938 11315 -9904
rect 11249 -9972 11265 -9938
rect 11299 -9972 11315 -9938
rect 11249 -9981 11315 -9972
rect 11349 -9871 11430 -9855
rect 11349 -9905 11363 -9871
rect 11397 -9905 11430 -9871
rect 11349 -9939 11430 -9905
rect 11349 -9973 11363 -9939
rect 11397 -9973 11430 -9939
rect 11349 -10010 11430 -9973
rect 11109 -10049 11227 -10015
rect 11193 -10083 11227 -10049
rect 11380 -10061 11430 -10010
rect 11464 -9892 11522 -9821
rect 11464 -9926 11476 -9892
rect 11510 -9926 11522 -9892
rect 11464 -9985 11522 -9926
rect 11464 -10019 11476 -9985
rect 11510 -10019 11522 -9985
rect 11464 -10054 11522 -10019
rect 11648 -9863 11982 -9821
rect 11648 -9897 11666 -9863
rect 11700 -9897 11930 -9863
rect 11964 -9897 11982 -9863
rect 11648 -9965 11982 -9897
rect 11648 -9999 11666 -9965
rect 11700 -9999 11930 -9965
rect 11964 -9999 11982 -9965
rect 11648 -10039 11982 -9999
rect 12384 -9892 12442 -9821
rect 12384 -9926 12396 -9892
rect 12430 -9926 12442 -9892
rect 12384 -9985 12442 -9926
rect 12384 -10019 12396 -9985
rect 12430 -10019 12442 -9985
rect 12476 -9870 12545 -9821
rect 12476 -9904 12502 -9870
rect 12536 -9904 12545 -9870
rect 12476 -9938 12545 -9904
rect 12476 -9972 12502 -9938
rect 12536 -9972 12545 -9938
rect 12476 -9988 12545 -9972
rect 12580 -9877 12631 -9861
rect 12580 -9911 12588 -9877
rect 12622 -9911 12631 -9877
rect 12580 -9965 12631 -9911
rect 10544 -10177 10694 -10107
rect 10728 -10094 10818 -10090
rect 10728 -10128 10763 -10094
rect 10797 -10099 10818 -10094
rect 10728 -10133 10768 -10128
rect 10802 -10133 10818 -10099
rect 10852 -10099 10938 -10085
rect 10852 -10133 10888 -10099
rect 10922 -10133 10938 -10099
rect 10852 -10143 10938 -10133
rect 10987 -10099 11159 -10084
rect 10987 -10133 11109 -10099
rect 11143 -10133 11159 -10099
rect 10987 -10134 11159 -10133
rect 11193 -10099 11346 -10083
rect 11193 -10133 11309 -10099
rect 11343 -10133 11346 -10099
rect 10852 -10167 10922 -10143
rect 8980 -10263 8998 -10229
rect 9032 -10263 9262 -10229
rect 9296 -10263 9314 -10229
rect 8980 -10331 9314 -10263
rect 9348 -10203 9406 -10186
rect 9348 -10237 9360 -10203
rect 9394 -10237 9406 -10203
rect 9348 -10331 9406 -10237
rect 9440 -10236 10142 -10177
rect 9440 -10270 9458 -10236
rect 9492 -10270 10090 -10236
rect 10124 -10270 10142 -10236
rect 9440 -10331 10142 -10270
rect 10176 -10203 10234 -10186
rect 10176 -10237 10188 -10203
rect 10222 -10237 10234 -10203
rect 10176 -10331 10234 -10237
rect 10360 -10229 10694 -10177
rect 10360 -10263 10378 -10229
rect 10412 -10263 10642 -10229
rect 10676 -10263 10694 -10229
rect 10360 -10331 10694 -10263
rect 10728 -10201 10922 -10167
rect 10728 -10244 10794 -10201
rect 10728 -10278 10747 -10244
rect 10781 -10278 10794 -10244
rect 10728 -10297 10794 -10278
rect 10828 -10244 10894 -10235
rect 10828 -10278 10844 -10244
rect 10878 -10278 10894 -10244
rect 10828 -10331 10894 -10278
rect 10987 -10244 11057 -10134
rect 11193 -10149 11346 -10133
rect 11380 -10095 11386 -10061
rect 11420 -10095 11430 -10061
rect 11193 -10168 11227 -10149
rect 10987 -10278 11004 -10244
rect 11038 -10278 11057 -10244
rect 10987 -10297 11057 -10278
rect 11109 -10202 11227 -10168
rect 11109 -10244 11159 -10202
rect 11380 -10220 11430 -10095
rect 11648 -10109 11798 -10039
rect 12384 -10054 12442 -10019
rect 12580 -9999 12588 -9965
rect 12622 -9999 12631 -9965
rect 12665 -9870 12717 -9821
rect 12665 -9904 12674 -9870
rect 12708 -9904 12717 -9870
rect 12665 -9938 12717 -9904
rect 12665 -9972 12674 -9938
rect 12708 -9972 12717 -9938
rect 12665 -9988 12717 -9972
rect 12752 -9877 12803 -9861
rect 12752 -9911 12760 -9877
rect 12794 -9911 12803 -9877
rect 12752 -9965 12803 -9911
rect 12580 -10022 12631 -9999
rect 12752 -9999 12760 -9965
rect 12794 -9999 12803 -9965
rect 12837 -9870 12889 -9821
rect 12837 -9904 12846 -9870
rect 12880 -9904 12889 -9870
rect 12837 -9938 12889 -9904
rect 12837 -9972 12846 -9938
rect 12880 -9972 12889 -9938
rect 12837 -9988 12889 -9972
rect 12923 -9877 12975 -9861
rect 12923 -9911 12932 -9877
rect 12966 -9911 12975 -9877
rect 12923 -9965 12975 -9911
rect 12752 -10022 12803 -9999
rect 12923 -9999 12932 -9965
rect 12966 -9999 12975 -9965
rect 13009 -9870 13086 -9821
rect 13009 -9904 13018 -9870
rect 13052 -9904 13086 -9870
rect 13009 -9938 13086 -9904
rect 13009 -9972 13018 -9938
rect 13052 -9972 13086 -9938
rect 13009 -9988 13086 -9972
rect 13120 -9892 13178 -9821
rect 13120 -9926 13132 -9892
rect 13166 -9926 13178 -9892
rect 13120 -9985 13178 -9926
rect 12923 -10022 12975 -9999
rect 13120 -10019 13132 -9985
rect 13166 -10019 13178 -9985
rect 12480 -10023 13086 -10022
rect 12514 -10056 13086 -10023
rect 13120 -10054 13178 -10019
rect 13212 -9863 13546 -9821
rect 13212 -9897 13230 -9863
rect 13264 -9897 13494 -9863
rect 13528 -9897 13546 -9863
rect 13212 -9965 13546 -9897
rect 13212 -9999 13230 -9965
rect 13264 -9999 13494 -9965
rect 13528 -9999 13546 -9965
rect 13212 -10039 13546 -9999
rect 11648 -10143 11668 -10109
rect 11702 -10143 11798 -10109
rect 11832 -10107 11928 -10073
rect 11962 -10107 11982 -10073
rect 11832 -10177 11982 -10107
rect 11143 -10278 11159 -10244
rect 11109 -10297 11159 -10278
rect 11249 -10244 11315 -10228
rect 11249 -10278 11265 -10244
rect 11299 -10278 11315 -10244
rect 11249 -10331 11315 -10278
rect 11349 -10244 11430 -10220
rect 11349 -10278 11363 -10244
rect 11397 -10278 11430 -10244
rect 11349 -10297 11430 -10278
rect 11464 -10203 11522 -10186
rect 11464 -10237 11476 -10203
rect 11510 -10237 11522 -10203
rect 11464 -10331 11522 -10237
rect 11648 -10229 11982 -10177
rect 12480 -10097 12514 -10057
rect 13026 -10082 13086 -10056
rect 12480 -10169 12514 -10131
rect 12548 -10093 12991 -10090
rect 12548 -10095 12858 -10093
rect 12548 -10129 12568 -10095
rect 12602 -10099 12659 -10095
rect 12693 -10099 12765 -10095
rect 12799 -10099 12858 -10095
rect 12892 -10099 12942 -10093
rect 12548 -10133 12574 -10129
rect 12608 -10133 12642 -10099
rect 12693 -10129 12710 -10099
rect 12676 -10133 12710 -10129
rect 12744 -10129 12765 -10099
rect 12744 -10133 12778 -10129
rect 12812 -10133 12846 -10099
rect 12892 -10127 12914 -10099
rect 12976 -10127 12991 -10093
rect 12880 -10133 12914 -10127
rect 12948 -10133 12991 -10127
rect 12548 -10135 12991 -10133
rect 13026 -10116 13039 -10082
rect 13073 -10116 13086 -10082
rect 13026 -10159 13086 -10116
rect 13026 -10169 13042 -10159
rect 11648 -10263 11666 -10229
rect 11700 -10263 11930 -10229
rect 11964 -10263 11982 -10229
rect 11648 -10331 11982 -10263
rect 12384 -10203 12442 -10186
rect 12514 -10193 13042 -10169
rect 13076 -10193 13086 -10159
rect 13212 -10107 13232 -10073
rect 13266 -10107 13362 -10073
rect 13212 -10177 13362 -10107
rect 13396 -10109 13546 -10039
rect 13580 -9892 13638 -9821
rect 13580 -9926 13592 -9892
rect 13626 -9926 13638 -9892
rect 13580 -9985 13638 -9926
rect 13674 -9863 13733 -9821
rect 13674 -9897 13690 -9863
rect 13724 -9897 13733 -9863
rect 13674 -9931 13733 -9897
rect 13674 -9965 13690 -9931
rect 13724 -9965 13733 -9931
rect 13674 -9983 13733 -9965
rect 13769 -9871 13818 -9855
rect 13769 -9905 13776 -9871
rect 13810 -9905 13818 -9871
rect 13769 -9939 13818 -9905
rect 13769 -9973 13776 -9939
rect 13810 -9973 13818 -9939
rect 13580 -10019 13592 -9985
rect 13626 -10019 13638 -9985
rect 13580 -10054 13638 -10019
rect 13769 -10083 13818 -9973
rect 13853 -9863 13905 -9821
rect 14025 -9822 15280 -9821
rect 13853 -9897 13862 -9863
rect 13896 -9897 13905 -9863
rect 13853 -9931 13905 -9897
rect 13853 -9965 13862 -9931
rect 13896 -9965 13905 -9931
rect 13853 -9983 13905 -9965
rect 13941 -9879 13991 -9856
rect 13941 -9913 13948 -9879
rect 13982 -9913 13991 -9879
rect 13941 -9947 13991 -9913
rect 13941 -9981 13948 -9947
rect 13982 -9981 13991 -9947
rect 14025 -9863 14077 -9822
rect 14025 -9897 14034 -9863
rect 14068 -9897 14077 -9863
rect 14025 -9931 14077 -9897
rect 14025 -9965 14034 -9931
rect 14068 -9965 14077 -9931
rect 14025 -9981 14077 -9965
rect 14111 -9907 14163 -9856
rect 14111 -9941 14120 -9907
rect 14154 -9941 14163 -9907
rect 13941 -10083 13991 -9981
rect 14111 -9993 14163 -9941
rect 14197 -9887 14249 -9822
rect 14197 -9921 14206 -9887
rect 14240 -9921 14249 -9887
rect 14197 -9967 14249 -9921
rect 14283 -9907 14335 -9856
rect 14283 -9941 14292 -9907
rect 14326 -9941 14335 -9907
rect 14111 -10027 14120 -9993
rect 14154 -10001 14163 -9993
rect 14283 -9993 14335 -9941
rect 14369 -9887 14421 -9822
rect 14369 -9921 14378 -9887
rect 14412 -9921 14421 -9887
rect 14369 -9967 14421 -9921
rect 14455 -9907 14507 -9856
rect 14455 -9941 14464 -9907
rect 14498 -9941 14507 -9907
rect 14283 -10001 14292 -9993
rect 14154 -10027 14292 -10001
rect 14326 -10001 14335 -9993
rect 14455 -9993 14507 -9941
rect 14541 -9887 14593 -9822
rect 14541 -9921 14550 -9887
rect 14584 -9921 14593 -9887
rect 14541 -9967 14593 -9921
rect 14627 -9907 14679 -9856
rect 14627 -9941 14636 -9907
rect 14670 -9941 14679 -9907
rect 14455 -10001 14464 -9993
rect 14326 -10027 14464 -10001
rect 14498 -10001 14507 -9993
rect 14627 -9993 14679 -9941
rect 14713 -9887 14762 -9822
rect 14713 -9921 14722 -9887
rect 14756 -9921 14762 -9887
rect 14713 -9967 14762 -9921
rect 14796 -9907 14848 -9856
rect 14796 -9941 14807 -9907
rect 14841 -9941 14848 -9907
rect 14627 -10001 14636 -9993
rect 14498 -10027 14636 -10001
rect 14670 -10001 14679 -9993
rect 14796 -9993 14848 -9941
rect 14885 -9887 14934 -9822
rect 14885 -9921 14893 -9887
rect 14927 -9921 14934 -9887
rect 14885 -9967 14934 -9921
rect 14968 -9907 15020 -9856
rect 14968 -9941 14979 -9907
rect 15013 -9941 15020 -9907
rect 14796 -10001 14807 -9993
rect 14670 -10027 14807 -10001
rect 14841 -10001 14848 -9993
rect 14968 -9993 15020 -9941
rect 15057 -9887 15106 -9822
rect 15057 -9921 15065 -9887
rect 15099 -9921 15106 -9887
rect 15057 -9967 15106 -9921
rect 15140 -9907 15192 -9856
rect 15140 -9941 15151 -9907
rect 15185 -9941 15192 -9907
rect 14968 -10001 14979 -9993
rect 14841 -10027 14979 -10001
rect 15013 -10001 15020 -9993
rect 15140 -9993 15192 -9941
rect 15229 -9887 15280 -9822
rect 15229 -9921 15237 -9887
rect 15271 -9921 15280 -9887
rect 15229 -9967 15280 -9921
rect 15314 -9907 15372 -9856
rect 15314 -9941 15323 -9907
rect 15357 -9941 15372 -9907
rect 15140 -10001 15151 -9993
rect 15013 -10027 15151 -10001
rect 15185 -10004 15192 -9993
rect 15314 -9993 15372 -9941
rect 15406 -9887 15460 -9821
rect 15406 -9921 15409 -9887
rect 15443 -9921 15460 -9887
rect 15406 -9970 15460 -9921
rect 15512 -9892 15570 -9821
rect 15512 -9926 15524 -9892
rect 15558 -9926 15570 -9892
rect 15314 -10004 15323 -9993
rect 15185 -10027 15323 -10004
rect 15357 -10004 15372 -9993
rect 15512 -9985 15570 -9926
rect 15357 -10027 15460 -10004
rect 14111 -10042 15460 -10027
rect 14111 -10049 15248 -10042
rect 15227 -10076 15248 -10049
rect 15282 -10076 15340 -10042
rect 15374 -10076 15460 -10042
rect 15512 -10019 15524 -9985
rect 15558 -10019 15570 -9985
rect 15512 -10054 15570 -10019
rect 15604 -9863 16673 -9821
rect 15604 -9897 15622 -9863
rect 15656 -9897 16622 -9863
rect 16656 -9897 16673 -9863
rect 15604 -9965 16673 -9897
rect 15604 -9999 15622 -9965
rect 15656 -9999 16622 -9965
rect 16656 -9999 16673 -9965
rect 15604 -10039 16673 -9999
rect 13396 -10143 13492 -10109
rect 13526 -10143 13546 -10109
rect 13672 -10099 13735 -10083
rect 13672 -10126 13692 -10099
rect 13672 -10160 13685 -10126
rect 13726 -10133 13735 -10099
rect 13719 -10160 13735 -10133
rect 12514 -10203 13086 -10193
rect 13120 -10203 13178 -10186
rect 12384 -10237 12396 -10203
rect 12430 -10237 12442 -10203
rect 12384 -10331 12442 -10237
rect 12572 -10253 12631 -10237
rect 12572 -10287 12588 -10253
rect 12622 -10287 12631 -10253
rect 12572 -10331 12631 -10287
rect 12665 -10242 12717 -10203
rect 12665 -10276 12674 -10242
rect 12708 -10276 12717 -10242
rect 12665 -10292 12717 -10276
rect 12751 -10253 12803 -10237
rect 12751 -10287 12760 -10253
rect 12794 -10287 12803 -10253
rect 12751 -10331 12803 -10287
rect 12837 -10242 12888 -10203
rect 13120 -10237 13132 -10203
rect 13166 -10237 13178 -10203
rect 12837 -10276 12846 -10242
rect 12880 -10276 12888 -10242
rect 12837 -10292 12888 -10276
rect 12922 -10253 12982 -10237
rect 12922 -10287 12932 -10253
rect 12966 -10287 12982 -10253
rect 12922 -10331 12982 -10287
rect 13120 -10331 13178 -10237
rect 13212 -10229 13546 -10177
rect 13212 -10263 13230 -10229
rect 13264 -10263 13494 -10229
rect 13528 -10263 13546 -10229
rect 13212 -10331 13546 -10263
rect 13580 -10203 13638 -10186
rect 13672 -10195 13735 -10160
rect 13769 -10099 15193 -10083
rect 13769 -10133 14119 -10099
rect 14153 -10133 14187 -10099
rect 14221 -10133 14255 -10099
rect 14289 -10133 14323 -10099
rect 14357 -10133 14391 -10099
rect 14425 -10133 14459 -10099
rect 14493 -10133 14527 -10099
rect 14561 -10133 14595 -10099
rect 14629 -10133 14663 -10099
rect 14697 -10133 14731 -10099
rect 14765 -10133 14799 -10099
rect 14833 -10133 14867 -10099
rect 14901 -10133 14935 -10099
rect 14969 -10133 15003 -10099
rect 15037 -10133 15071 -10099
rect 15105 -10133 15139 -10099
rect 15173 -10133 15193 -10099
rect 13580 -10237 13592 -10203
rect 13626 -10237 13638 -10203
rect 13580 -10331 13638 -10237
rect 13672 -10255 13733 -10229
rect 13672 -10289 13690 -10255
rect 13724 -10289 13733 -10255
rect 13672 -10331 13733 -10289
rect 13769 -10242 13819 -10133
rect 13769 -10276 13776 -10242
rect 13810 -10276 13819 -10242
rect 13769 -10295 13819 -10276
rect 13853 -10242 13905 -10226
rect 13853 -10276 13862 -10242
rect 13896 -10276 13905 -10242
rect 13853 -10331 13905 -10276
rect 13941 -10242 13991 -10133
rect 15227 -10138 15460 -10076
rect 15227 -10167 15248 -10138
rect 14111 -10172 15248 -10167
rect 15282 -10172 15341 -10138
rect 15375 -10172 15460 -10138
rect 14111 -10201 15460 -10172
rect 15604 -10107 15682 -10073
rect 15716 -10107 15810 -10073
rect 15844 -10107 15938 -10073
rect 15972 -10107 16066 -10073
rect 16100 -10107 16120 -10073
rect 15604 -10177 16120 -10107
rect 16154 -10109 16673 -10039
rect 16154 -10143 16174 -10109
rect 16208 -10143 16302 -10109
rect 16336 -10143 16430 -10109
rect 16464 -10143 16558 -10109
rect 16592 -10143 16673 -10109
rect 13941 -10276 13948 -10242
rect 13982 -10276 13991 -10242
rect 13941 -10295 13991 -10276
rect 14025 -10242 14077 -10219
rect 14025 -10276 14034 -10242
rect 14068 -10276 14077 -10242
rect 14025 -10331 14077 -10276
rect 14111 -10242 14163 -10201
rect 14111 -10276 14120 -10242
rect 14154 -10276 14163 -10242
rect 14111 -10292 14163 -10276
rect 14197 -10251 14249 -10235
rect 14197 -10285 14206 -10251
rect 14240 -10285 14249 -10251
rect 14197 -10331 14249 -10285
rect 14283 -10242 14335 -10201
rect 14283 -10276 14292 -10242
rect 14326 -10276 14335 -10242
rect 14283 -10292 14335 -10276
rect 14369 -10251 14421 -10235
rect 14369 -10285 14378 -10251
rect 14412 -10285 14421 -10251
rect 14369 -10331 14421 -10285
rect 14455 -10242 14507 -10201
rect 14455 -10276 14464 -10242
rect 14498 -10276 14507 -10242
rect 14455 -10292 14507 -10276
rect 14541 -10251 14590 -10235
rect 14541 -10285 14550 -10251
rect 14584 -10285 14590 -10251
rect 14541 -10331 14590 -10285
rect 14624 -10242 14679 -10201
rect 14624 -10276 14636 -10242
rect 14670 -10276 14679 -10242
rect 14624 -10292 14679 -10276
rect 14713 -10251 14762 -10235
rect 14713 -10285 14722 -10251
rect 14756 -10285 14762 -10251
rect 14713 -10331 14762 -10285
rect 14796 -10242 14848 -10201
rect 14796 -10276 14807 -10242
rect 14841 -10276 14848 -10242
rect 14796 -10292 14848 -10276
rect 14884 -10251 14934 -10235
rect 14884 -10285 14893 -10251
rect 14927 -10285 14934 -10251
rect 14884 -10331 14934 -10285
rect 14968 -10242 15020 -10201
rect 14968 -10276 14979 -10242
rect 15013 -10276 15020 -10242
rect 14968 -10292 15020 -10276
rect 15056 -10251 15106 -10235
rect 15056 -10285 15065 -10251
rect 15099 -10285 15106 -10251
rect 15056 -10331 15106 -10285
rect 15140 -10242 15192 -10201
rect 15140 -10276 15151 -10242
rect 15185 -10276 15192 -10242
rect 15140 -10292 15192 -10276
rect 15228 -10251 15280 -10235
rect 15228 -10285 15237 -10251
rect 15271 -10285 15280 -10251
rect 15228 -10331 15280 -10285
rect 15314 -10242 15366 -10201
rect 15512 -10203 15570 -10186
rect 15314 -10276 15323 -10242
rect 15357 -10276 15366 -10242
rect 15314 -10292 15366 -10276
rect 15400 -10251 15460 -10235
rect 15400 -10285 15409 -10251
rect 15443 -10285 15460 -10251
rect 15400 -10331 15460 -10285
rect 15512 -10237 15524 -10203
rect 15558 -10237 15570 -10203
rect 15512 -10331 15570 -10237
rect 15604 -10236 16673 -10177
rect 15604 -10270 15622 -10236
rect 15656 -10270 16622 -10236
rect 16656 -10270 16673 -10236
rect 15604 -10331 16673 -10270
rect -2997 -10365 -2968 -10331
rect -2934 -10365 -2876 -10331
rect -2842 -10365 -2784 -10331
rect -2750 -10365 -2692 -10331
rect -2658 -10365 -2600 -10331
rect -2566 -10365 -2508 -10331
rect -2474 -10365 -2416 -10331
rect -2382 -10365 -2324 -10331
rect -2290 -10365 -2232 -10331
rect -2198 -10365 -2140 -10331
rect -2106 -10365 -2048 -10331
rect -2014 -10365 -1956 -10331
rect -1922 -10365 -1864 -10331
rect -1830 -10365 -1772 -10331
rect -1738 -10365 -1680 -10331
rect -1646 -10365 -1588 -10331
rect -1554 -10365 -1496 -10331
rect -1462 -10365 -1404 -10331
rect -1370 -10365 -1312 -10331
rect -1278 -10365 -1220 -10331
rect -1186 -10365 -1128 -10331
rect -1094 -10365 -1036 -10331
rect -1002 -10365 -944 -10331
rect -910 -10365 -852 -10331
rect -818 -10365 -760 -10331
rect -726 -10365 -668 -10331
rect -634 -10365 -576 -10331
rect -542 -10365 -484 -10331
rect -450 -10365 -392 -10331
rect -358 -10365 -300 -10331
rect -266 -10365 -208 -10331
rect -174 -10365 -116 -10331
rect -82 -10365 -24 -10331
rect 10 -10365 68 -10331
rect 102 -10365 160 -10331
rect 194 -10365 252 -10331
rect 286 -10365 344 -10331
rect 378 -10365 436 -10331
rect 470 -10365 528 -10331
rect 562 -10365 620 -10331
rect 654 -10365 712 -10331
rect 746 -10365 804 -10331
rect 838 -10365 896 -10331
rect 930 -10365 988 -10331
rect 1022 -10365 1080 -10331
rect 1114 -10365 1172 -10331
rect 1206 -10365 1264 -10331
rect 1298 -10365 1356 -10331
rect 1390 -10365 1448 -10331
rect 1482 -10365 1540 -10331
rect 1574 -10365 1632 -10331
rect 1666 -10365 1724 -10331
rect 1758 -10365 1816 -10331
rect 1850 -10365 1908 -10331
rect 1942 -10365 2000 -10331
rect 2034 -10365 2092 -10331
rect 2126 -10365 2184 -10331
rect 2218 -10365 2276 -10331
rect 2310 -10365 2368 -10331
rect 2402 -10365 2460 -10331
rect 2494 -10365 2552 -10331
rect 2586 -10365 2644 -10331
rect 2678 -10365 2736 -10331
rect 2770 -10365 2828 -10331
rect 2862 -10365 2920 -10331
rect 2954 -10365 3012 -10331
rect 3046 -10365 3104 -10331
rect 3138 -10365 3196 -10331
rect 3230 -10365 3288 -10331
rect 3322 -10365 3380 -10331
rect 3414 -10365 3472 -10331
rect 3506 -10365 3564 -10331
rect 3598 -10365 3656 -10331
rect 3690 -10365 3748 -10331
rect 3782 -10365 3840 -10331
rect 3874 -10365 3932 -10331
rect 3966 -10365 4024 -10331
rect 4058 -10365 4116 -10331
rect 4150 -10365 4208 -10331
rect 4242 -10365 4300 -10331
rect 4334 -10365 4392 -10331
rect 4426 -10365 4484 -10331
rect 4518 -10365 4576 -10331
rect 4610 -10365 4668 -10331
rect 4702 -10365 4760 -10331
rect 4794 -10365 4852 -10331
rect 4886 -10365 4944 -10331
rect 4978 -10365 5036 -10331
rect 5070 -10365 5128 -10331
rect 5162 -10365 5220 -10331
rect 5254 -10365 5312 -10331
rect 5346 -10365 5404 -10331
rect 5438 -10365 5496 -10331
rect 5530 -10365 5588 -10331
rect 5622 -10365 5680 -10331
rect 5714 -10365 5772 -10331
rect 5806 -10365 5864 -10331
rect 5898 -10365 5956 -10331
rect 5990 -10365 6048 -10331
rect 6082 -10365 6140 -10331
rect 6174 -10365 6232 -10331
rect 6266 -10365 6324 -10331
rect 6358 -10365 6416 -10331
rect 6450 -10365 6508 -10331
rect 6542 -10365 6600 -10331
rect 6634 -10365 6692 -10331
rect 6726 -10365 6784 -10331
rect 6818 -10365 6876 -10331
rect 6910 -10365 6968 -10331
rect 7002 -10365 7060 -10331
rect 7094 -10365 7152 -10331
rect 7186 -10365 7244 -10331
rect 7278 -10365 7336 -10331
rect 7370 -10365 7428 -10331
rect 7462 -10365 7520 -10331
rect 7554 -10365 7612 -10331
rect 7646 -10365 7704 -10331
rect 7738 -10365 7796 -10331
rect 7830 -10365 7888 -10331
rect 7922 -10365 7980 -10331
rect 8014 -10365 8072 -10331
rect 8106 -10365 8164 -10331
rect 8198 -10365 8256 -10331
rect 8290 -10365 8348 -10331
rect 8382 -10365 8440 -10331
rect 8474 -10365 8532 -10331
rect 8566 -10365 8624 -10331
rect 8658 -10365 8716 -10331
rect 8750 -10365 8808 -10331
rect 8842 -10365 8900 -10331
rect 8934 -10365 8992 -10331
rect 9026 -10365 9084 -10331
rect 9118 -10365 9176 -10331
rect 9210 -10365 9268 -10331
rect 9302 -10365 9360 -10331
rect 9394 -10365 9452 -10331
rect 9486 -10365 9544 -10331
rect 9578 -10365 9636 -10331
rect 9670 -10365 9728 -10331
rect 9762 -10365 9820 -10331
rect 9854 -10365 9912 -10331
rect 9946 -10365 10004 -10331
rect 10038 -10365 10096 -10331
rect 10130 -10365 10188 -10331
rect 10222 -10365 10280 -10331
rect 10314 -10365 10372 -10331
rect 10406 -10365 10464 -10331
rect 10498 -10365 10556 -10331
rect 10590 -10365 10648 -10331
rect 10682 -10365 10740 -10331
rect 10774 -10365 10832 -10331
rect 10866 -10365 10924 -10331
rect 10958 -10365 11016 -10331
rect 11050 -10365 11108 -10331
rect 11142 -10365 11200 -10331
rect 11234 -10365 11292 -10331
rect 11326 -10365 11384 -10331
rect 11418 -10365 11476 -10331
rect 11510 -10365 11568 -10331
rect 11602 -10365 11660 -10331
rect 11694 -10365 11752 -10331
rect 11786 -10365 11844 -10331
rect 11878 -10365 11936 -10331
rect 11970 -10365 12028 -10331
rect 12062 -10365 12120 -10331
rect 12154 -10365 12212 -10331
rect 12246 -10365 12304 -10331
rect 12338 -10365 12396 -10331
rect 12430 -10365 12488 -10331
rect 12522 -10365 12580 -10331
rect 12614 -10365 12672 -10331
rect 12706 -10365 12764 -10331
rect 12798 -10365 12856 -10331
rect 12890 -10365 12948 -10331
rect 12982 -10365 13040 -10331
rect 13074 -10365 13132 -10331
rect 13166 -10365 13224 -10331
rect 13258 -10365 13316 -10331
rect 13350 -10365 13408 -10331
rect 13442 -10365 13500 -10331
rect 13534 -10365 13592 -10331
rect 13626 -10365 13684 -10331
rect 13718 -10365 13776 -10331
rect 13810 -10365 13868 -10331
rect 13902 -10365 13960 -10331
rect 13994 -10365 14052 -10331
rect 14086 -10365 14144 -10331
rect 14178 -10365 14236 -10331
rect 14270 -10365 14328 -10331
rect 14362 -10365 14420 -10331
rect 14454 -10365 14512 -10331
rect 14546 -10365 14604 -10331
rect 14638 -10365 14696 -10331
rect 14730 -10365 14788 -10331
rect 14822 -10365 14880 -10331
rect 14914 -10365 14972 -10331
rect 15006 -10365 15064 -10331
rect 15098 -10365 15156 -10331
rect 15190 -10365 15248 -10331
rect 15282 -10365 15340 -10331
rect 15374 -10365 15432 -10331
rect 15466 -10365 15524 -10331
rect 15558 -10365 15616 -10331
rect 15650 -10365 15708 -10331
rect 15742 -10365 15800 -10331
rect 15834 -10365 15892 -10331
rect 15926 -10365 15984 -10331
rect 16018 -10365 16076 -10331
rect 16110 -10365 16168 -10331
rect 16202 -10365 16260 -10331
rect 16294 -10365 16352 -10331
rect 16386 -10365 16444 -10331
rect 16478 -10365 16536 -10331
rect 16570 -10365 16628 -10331
rect 16662 -10365 16691 -10331
rect -2980 -10426 -2278 -10365
rect -2980 -10460 -2962 -10426
rect -2928 -10460 -2330 -10426
rect -2296 -10460 -2278 -10426
rect -2980 -10519 -2278 -10460
rect -2244 -10459 -2186 -10365
rect -1882 -10418 -1817 -10399
rect -2244 -10493 -2232 -10459
rect -2198 -10493 -2186 -10459
rect -2244 -10510 -2186 -10493
rect -1968 -10499 -1920 -10423
rect -2980 -10587 -2902 -10553
rect -2868 -10587 -2799 -10553
rect -2765 -10587 -2696 -10553
rect -2662 -10587 -2642 -10553
rect -2980 -10657 -2642 -10587
rect -2608 -10589 -2278 -10519
rect -2608 -10623 -2588 -10589
rect -2554 -10623 -2489 -10589
rect -2455 -10623 -2390 -10589
rect -2356 -10623 -2278 -10589
rect -1968 -10533 -1961 -10499
rect -1927 -10533 -1920 -10499
rect -1968 -10563 -1920 -10533
rect -1968 -10597 -1954 -10563
rect -1968 -10613 -1920 -10597
rect -1882 -10452 -1867 -10418
rect -1833 -10452 -1817 -10418
rect -1882 -10500 -1817 -10452
rect -1783 -10416 -1726 -10365
rect -1749 -10450 -1726 -10416
rect -1783 -10466 -1726 -10450
rect -1692 -10459 -1634 -10365
rect -1692 -10493 -1680 -10459
rect -1646 -10493 -1634 -10459
rect -1882 -10534 -1726 -10500
rect -1692 -10510 -1634 -10493
rect -1600 -10426 -898 -10365
rect -1600 -10460 -1582 -10426
rect -1548 -10460 -950 -10426
rect -916 -10460 -898 -10426
rect -1600 -10519 -898 -10460
rect -864 -10426 -162 -10365
rect -864 -10460 -846 -10426
rect -812 -10460 -214 -10426
rect -180 -10460 -162 -10426
rect -864 -10519 -162 -10460
rect -128 -10459 -70 -10365
rect -128 -10493 -116 -10459
rect -82 -10493 -70 -10459
rect -128 -10510 -70 -10493
rect -36 -10433 298 -10365
rect -36 -10467 -18 -10433
rect 16 -10467 246 -10433
rect 280 -10467 298 -10433
rect -36 -10519 298 -10467
rect 332 -10459 390 -10365
rect 332 -10493 344 -10459
rect 378 -10493 390 -10459
rect 332 -10510 390 -10493
rect 424 -10418 505 -10399
rect 424 -10452 457 -10418
rect 491 -10452 505 -10418
rect 424 -10476 505 -10452
rect 539 -10418 605 -10365
rect 539 -10452 555 -10418
rect 589 -10452 605 -10418
rect 539 -10468 605 -10452
rect 695 -10418 745 -10399
rect 695 -10452 711 -10418
rect -1882 -10568 -1813 -10534
rect -1779 -10568 -1726 -10534
rect -1882 -10606 -1726 -10568
rect -1600 -10587 -1522 -10553
rect -1488 -10587 -1419 -10553
rect -1385 -10587 -1316 -10553
rect -1282 -10587 -1262 -10553
rect -2980 -10697 -2278 -10657
rect -2980 -10731 -2962 -10697
rect -2928 -10731 -2330 -10697
rect -2296 -10731 -2278 -10697
rect -2980 -10799 -2278 -10731
rect -2980 -10833 -2962 -10799
rect -2928 -10833 -2330 -10799
rect -2296 -10833 -2278 -10799
rect -2980 -10875 -2278 -10833
rect -2244 -10677 -2186 -10642
rect -2244 -10711 -2232 -10677
rect -2198 -10711 -2186 -10677
rect -2244 -10770 -2186 -10711
rect -2244 -10804 -2232 -10770
rect -2198 -10804 -2186 -10770
rect -2244 -10875 -2186 -10804
rect -1968 -10697 -1916 -10681
rect -1968 -10731 -1950 -10697
rect -1968 -10799 -1916 -10731
rect -1968 -10833 -1950 -10799
rect -1968 -10875 -1916 -10833
rect -1882 -10697 -1816 -10606
rect -1692 -10677 -1634 -10642
rect -1882 -10731 -1866 -10697
rect -1832 -10731 -1816 -10697
rect -1882 -10799 -1816 -10731
rect -1882 -10833 -1866 -10799
rect -1832 -10833 -1816 -10799
rect -1882 -10841 -1816 -10833
rect -1782 -10697 -1726 -10681
rect -1748 -10731 -1726 -10697
rect -1782 -10799 -1726 -10731
rect -1748 -10833 -1726 -10799
rect -1782 -10875 -1726 -10833
rect -1692 -10711 -1680 -10677
rect -1646 -10711 -1634 -10677
rect -1692 -10770 -1634 -10711
rect -1692 -10804 -1680 -10770
rect -1646 -10804 -1634 -10770
rect -1692 -10875 -1634 -10804
rect -1600 -10657 -1262 -10587
rect -1228 -10589 -898 -10519
rect -1228 -10623 -1208 -10589
rect -1174 -10623 -1109 -10589
rect -1075 -10623 -1010 -10589
rect -976 -10623 -898 -10589
rect -864 -10587 -786 -10553
rect -752 -10587 -683 -10553
rect -649 -10587 -580 -10553
rect -546 -10587 -526 -10553
rect -864 -10657 -526 -10587
rect -492 -10589 -162 -10519
rect -492 -10623 -472 -10589
rect -438 -10623 -373 -10589
rect -339 -10623 -274 -10589
rect -240 -10623 -162 -10589
rect -36 -10587 -16 -10553
rect 18 -10587 114 -10553
rect -1600 -10697 -898 -10657
rect -1600 -10731 -1582 -10697
rect -1548 -10731 -950 -10697
rect -916 -10731 -898 -10697
rect -1600 -10799 -898 -10731
rect -1600 -10833 -1582 -10799
rect -1548 -10833 -950 -10799
rect -916 -10833 -898 -10799
rect -1600 -10875 -898 -10833
rect -864 -10697 -162 -10657
rect -864 -10731 -846 -10697
rect -812 -10731 -214 -10697
rect -180 -10731 -162 -10697
rect -864 -10799 -162 -10731
rect -864 -10833 -846 -10799
rect -812 -10833 -214 -10799
rect -180 -10833 -162 -10799
rect -864 -10875 -162 -10833
rect -128 -10677 -70 -10642
rect -128 -10711 -116 -10677
rect -82 -10711 -70 -10677
rect -128 -10770 -70 -10711
rect -128 -10804 -116 -10770
rect -82 -10804 -70 -10770
rect -128 -10875 -70 -10804
rect -36 -10657 114 -10587
rect 148 -10589 298 -10519
rect 148 -10623 244 -10589
rect 278 -10623 298 -10589
rect 424 -10603 474 -10476
rect 695 -10494 745 -10452
rect 627 -10528 745 -10494
rect 797 -10418 867 -10399
rect 797 -10452 816 -10418
rect 850 -10452 867 -10418
rect 627 -10547 661 -10528
rect 424 -10637 429 -10603
rect 463 -10637 474 -10603
rect 508 -10563 661 -10547
rect 797 -10562 867 -10452
rect 960 -10418 1026 -10365
rect 960 -10452 976 -10418
rect 1010 -10452 1026 -10418
rect 960 -10461 1026 -10452
rect 1060 -10418 1126 -10399
rect 1060 -10452 1073 -10418
rect 1107 -10452 1126 -10418
rect 1060 -10495 1126 -10452
rect 932 -10529 1126 -10495
rect 1160 -10459 1218 -10365
rect 1160 -10493 1172 -10459
rect 1206 -10493 1218 -10459
rect 1160 -10510 1218 -10493
rect 1252 -10433 1586 -10365
rect 1252 -10467 1270 -10433
rect 1304 -10467 1534 -10433
rect 1568 -10467 1586 -10433
rect 1252 -10519 1586 -10467
rect 1620 -10459 1678 -10365
rect 1620 -10493 1632 -10459
rect 1666 -10493 1678 -10459
rect 1620 -10510 1678 -10493
rect 1712 -10426 2414 -10365
rect 1712 -10460 1730 -10426
rect 1764 -10460 2362 -10426
rect 2396 -10460 2414 -10426
rect 1712 -10519 2414 -10460
rect 2448 -10459 2506 -10365
rect 2448 -10493 2460 -10459
rect 2494 -10493 2506 -10459
rect 2448 -10510 2506 -10493
rect 2540 -10433 2874 -10365
rect 2540 -10467 2558 -10433
rect 2592 -10467 2822 -10433
rect 2856 -10467 2874 -10433
rect 2540 -10519 2874 -10467
rect 2908 -10459 2966 -10365
rect 2908 -10493 2920 -10459
rect 2954 -10493 2966 -10459
rect 2908 -10510 2966 -10493
rect 3000 -10418 3081 -10399
rect 3000 -10452 3033 -10418
rect 3067 -10452 3081 -10418
rect 3000 -10476 3081 -10452
rect 3115 -10418 3181 -10365
rect 3115 -10452 3131 -10418
rect 3165 -10452 3181 -10418
rect 3115 -10468 3181 -10452
rect 3271 -10418 3321 -10399
rect 3271 -10452 3287 -10418
rect 932 -10553 1002 -10529
rect 508 -10597 511 -10563
rect 545 -10597 661 -10563
rect 508 -10613 661 -10597
rect 695 -10563 867 -10562
rect 695 -10597 711 -10563
rect 745 -10597 867 -10563
rect 695 -10612 867 -10597
rect 916 -10563 1002 -10553
rect 916 -10597 932 -10563
rect 966 -10597 1002 -10563
rect 916 -10611 1002 -10597
rect 1036 -10597 1052 -10563
rect 1086 -10568 1126 -10563
rect 1036 -10602 1072 -10597
rect 1106 -10602 1126 -10568
rect 1036 -10606 1126 -10602
rect 1252 -10587 1272 -10553
rect 1306 -10587 1402 -10553
rect -36 -10697 298 -10657
rect -36 -10731 -18 -10697
rect 16 -10731 246 -10697
rect 280 -10731 298 -10697
rect -36 -10799 298 -10731
rect -36 -10833 -18 -10799
rect 16 -10833 246 -10799
rect 280 -10833 298 -10799
rect -36 -10875 298 -10833
rect 332 -10677 390 -10642
rect 332 -10711 344 -10677
rect 378 -10711 390 -10677
rect 332 -10770 390 -10711
rect 332 -10804 344 -10770
rect 378 -10804 390 -10770
rect 332 -10875 390 -10804
rect 424 -10686 474 -10637
rect 627 -10647 661 -10613
rect 627 -10681 745 -10647
rect 424 -10723 505 -10686
rect 424 -10757 457 -10723
rect 491 -10757 505 -10723
rect 424 -10791 505 -10757
rect 424 -10825 457 -10791
rect 491 -10825 505 -10791
rect 424 -10841 505 -10825
rect 539 -10724 605 -10715
rect 539 -10758 555 -10724
rect 589 -10758 605 -10724
rect 539 -10792 605 -10758
rect 539 -10826 555 -10792
rect 589 -10826 605 -10792
rect 539 -10875 605 -10826
rect 695 -10723 745 -10681
rect 695 -10757 711 -10723
rect 695 -10791 745 -10757
rect 695 -10825 711 -10791
rect 695 -10841 745 -10825
rect 797 -10724 867 -10612
rect 932 -10640 1002 -10611
rect 932 -10674 1126 -10640
rect 797 -10758 815 -10724
rect 849 -10758 867 -10724
rect 797 -10792 867 -10758
rect 797 -10826 815 -10792
rect 849 -10826 867 -10792
rect 797 -10841 867 -10826
rect 957 -10724 1023 -10708
rect 957 -10758 973 -10724
rect 1007 -10758 1023 -10724
rect 957 -10792 1023 -10758
rect 957 -10826 973 -10792
rect 1007 -10826 1023 -10792
rect 957 -10875 1023 -10826
rect 1057 -10724 1126 -10674
rect 1057 -10758 1073 -10724
rect 1107 -10758 1126 -10724
rect 1057 -10792 1126 -10758
rect 1057 -10826 1073 -10792
rect 1107 -10826 1126 -10792
rect 1057 -10841 1126 -10826
rect 1160 -10677 1218 -10642
rect 1160 -10711 1172 -10677
rect 1206 -10711 1218 -10677
rect 1160 -10770 1218 -10711
rect 1160 -10804 1172 -10770
rect 1206 -10804 1218 -10770
rect 1160 -10875 1218 -10804
rect 1252 -10657 1402 -10587
rect 1436 -10589 1586 -10519
rect 1436 -10623 1532 -10589
rect 1566 -10623 1586 -10589
rect 1712 -10587 1790 -10553
rect 1824 -10587 1893 -10553
rect 1927 -10587 1996 -10553
rect 2030 -10587 2050 -10553
rect 1252 -10697 1586 -10657
rect 1252 -10731 1270 -10697
rect 1304 -10731 1534 -10697
rect 1568 -10731 1586 -10697
rect 1252 -10799 1586 -10731
rect 1252 -10833 1270 -10799
rect 1304 -10833 1534 -10799
rect 1568 -10833 1586 -10799
rect 1252 -10875 1586 -10833
rect 1620 -10677 1678 -10642
rect 1620 -10711 1632 -10677
rect 1666 -10711 1678 -10677
rect 1620 -10770 1678 -10711
rect 1620 -10804 1632 -10770
rect 1666 -10804 1678 -10770
rect 1620 -10875 1678 -10804
rect 1712 -10657 2050 -10587
rect 2084 -10589 2414 -10519
rect 2084 -10623 2104 -10589
rect 2138 -10623 2203 -10589
rect 2237 -10623 2302 -10589
rect 2336 -10623 2414 -10589
rect 2540 -10587 2560 -10553
rect 2594 -10587 2690 -10553
rect 1712 -10697 2414 -10657
rect 1712 -10731 1730 -10697
rect 1764 -10731 2362 -10697
rect 2396 -10731 2414 -10697
rect 1712 -10799 2414 -10731
rect 1712 -10833 1730 -10799
rect 1764 -10833 2362 -10799
rect 2396 -10833 2414 -10799
rect 1712 -10875 2414 -10833
rect 2448 -10677 2506 -10642
rect 2448 -10711 2460 -10677
rect 2494 -10711 2506 -10677
rect 2448 -10770 2506 -10711
rect 2448 -10804 2460 -10770
rect 2494 -10804 2506 -10770
rect 2448 -10875 2506 -10804
rect 2540 -10657 2690 -10587
rect 2724 -10589 2874 -10519
rect 2724 -10623 2820 -10589
rect 2854 -10623 2874 -10589
rect 3000 -10569 3050 -10476
rect 3271 -10494 3321 -10452
rect 3203 -10528 3321 -10494
rect 3373 -10418 3443 -10399
rect 3373 -10452 3392 -10418
rect 3426 -10452 3443 -10418
rect 3203 -10547 3237 -10528
rect 3000 -10603 3016 -10569
rect 2540 -10697 2874 -10657
rect 2540 -10731 2558 -10697
rect 2592 -10731 2822 -10697
rect 2856 -10731 2874 -10697
rect 2540 -10799 2874 -10731
rect 2540 -10833 2558 -10799
rect 2592 -10833 2822 -10799
rect 2856 -10833 2874 -10799
rect 2540 -10875 2874 -10833
rect 2908 -10677 2966 -10642
rect 2908 -10711 2920 -10677
rect 2954 -10711 2966 -10677
rect 2908 -10770 2966 -10711
rect 2908 -10804 2920 -10770
rect 2954 -10804 2966 -10770
rect 2908 -10875 2966 -10804
rect 3000 -10686 3050 -10603
rect 3084 -10563 3237 -10547
rect 3373 -10562 3443 -10452
rect 3536 -10418 3602 -10365
rect 3536 -10452 3552 -10418
rect 3586 -10452 3602 -10418
rect 3536 -10461 3602 -10452
rect 3636 -10418 3702 -10399
rect 3636 -10452 3649 -10418
rect 3683 -10452 3702 -10418
rect 3636 -10495 3702 -10452
rect 3508 -10529 3702 -10495
rect 3736 -10459 3794 -10365
rect 3736 -10493 3748 -10459
rect 3782 -10493 3794 -10459
rect 3736 -10510 3794 -10493
rect 3828 -10433 4162 -10365
rect 3828 -10467 3846 -10433
rect 3880 -10467 4110 -10433
rect 4144 -10467 4162 -10433
rect 3828 -10519 4162 -10467
rect 4196 -10459 4254 -10365
rect 4196 -10493 4208 -10459
rect 4242 -10493 4254 -10459
rect 4196 -10510 4254 -10493
rect 4288 -10426 4990 -10365
rect 4288 -10460 4306 -10426
rect 4340 -10460 4938 -10426
rect 4972 -10460 4990 -10426
rect 4288 -10519 4990 -10460
rect 5024 -10459 5082 -10365
rect 5024 -10493 5036 -10459
rect 5070 -10493 5082 -10459
rect 5024 -10510 5082 -10493
rect 5116 -10433 5450 -10365
rect 5116 -10467 5134 -10433
rect 5168 -10467 5398 -10433
rect 5432 -10467 5450 -10433
rect 5116 -10519 5450 -10467
rect 5484 -10459 5542 -10365
rect 5484 -10493 5496 -10459
rect 5530 -10493 5542 -10459
rect 5484 -10510 5542 -10493
rect 5576 -10418 5657 -10399
rect 5576 -10452 5609 -10418
rect 5643 -10452 5657 -10418
rect 5576 -10476 5657 -10452
rect 5691 -10418 5757 -10365
rect 5691 -10452 5707 -10418
rect 5741 -10452 5757 -10418
rect 5691 -10468 5757 -10452
rect 5847 -10418 5897 -10399
rect 5847 -10452 5863 -10418
rect 3508 -10553 3578 -10529
rect 3084 -10597 3087 -10563
rect 3121 -10597 3237 -10563
rect 3084 -10613 3237 -10597
rect 3271 -10563 3443 -10562
rect 3271 -10597 3287 -10563
rect 3321 -10597 3443 -10563
rect 3271 -10612 3443 -10597
rect 3492 -10563 3578 -10553
rect 3492 -10597 3508 -10563
rect 3542 -10597 3578 -10563
rect 3492 -10611 3578 -10597
rect 3612 -10597 3628 -10563
rect 3662 -10569 3702 -10563
rect 3612 -10603 3630 -10597
rect 3664 -10603 3702 -10569
rect 3612 -10606 3702 -10603
rect 3828 -10587 3848 -10553
rect 3882 -10587 3978 -10553
rect 3203 -10647 3237 -10613
rect 3203 -10681 3321 -10647
rect 3000 -10723 3081 -10686
rect 3000 -10757 3033 -10723
rect 3067 -10757 3081 -10723
rect 3000 -10791 3081 -10757
rect 3000 -10825 3033 -10791
rect 3067 -10825 3081 -10791
rect 3000 -10841 3081 -10825
rect 3115 -10724 3181 -10715
rect 3115 -10758 3131 -10724
rect 3165 -10758 3181 -10724
rect 3115 -10792 3181 -10758
rect 3115 -10826 3131 -10792
rect 3165 -10826 3181 -10792
rect 3115 -10875 3181 -10826
rect 3271 -10723 3321 -10681
rect 3271 -10757 3287 -10723
rect 3271 -10791 3321 -10757
rect 3271 -10825 3287 -10791
rect 3271 -10841 3321 -10825
rect 3373 -10724 3443 -10612
rect 3508 -10640 3578 -10611
rect 3508 -10674 3702 -10640
rect 3373 -10758 3391 -10724
rect 3425 -10758 3443 -10724
rect 3373 -10792 3443 -10758
rect 3373 -10826 3391 -10792
rect 3425 -10826 3443 -10792
rect 3373 -10841 3443 -10826
rect 3533 -10724 3599 -10708
rect 3533 -10758 3549 -10724
rect 3583 -10758 3599 -10724
rect 3533 -10792 3599 -10758
rect 3533 -10826 3549 -10792
rect 3583 -10826 3599 -10792
rect 3533 -10875 3599 -10826
rect 3633 -10724 3702 -10674
rect 3633 -10758 3649 -10724
rect 3683 -10758 3702 -10724
rect 3633 -10792 3702 -10758
rect 3633 -10826 3649 -10792
rect 3683 -10826 3702 -10792
rect 3633 -10841 3702 -10826
rect 3736 -10677 3794 -10642
rect 3736 -10711 3748 -10677
rect 3782 -10711 3794 -10677
rect 3736 -10770 3794 -10711
rect 3736 -10804 3748 -10770
rect 3782 -10804 3794 -10770
rect 3736 -10875 3794 -10804
rect 3828 -10657 3978 -10587
rect 4012 -10589 4162 -10519
rect 4012 -10623 4108 -10589
rect 4142 -10623 4162 -10589
rect 4288 -10587 4366 -10553
rect 4400 -10587 4469 -10553
rect 4503 -10587 4572 -10553
rect 4606 -10587 4626 -10553
rect 3828 -10697 4162 -10657
rect 3828 -10731 3846 -10697
rect 3880 -10731 4110 -10697
rect 4144 -10731 4162 -10697
rect 3828 -10799 4162 -10731
rect 3828 -10833 3846 -10799
rect 3880 -10833 4110 -10799
rect 4144 -10833 4162 -10799
rect 3828 -10875 4162 -10833
rect 4196 -10677 4254 -10642
rect 4196 -10711 4208 -10677
rect 4242 -10711 4254 -10677
rect 4196 -10770 4254 -10711
rect 4196 -10804 4208 -10770
rect 4242 -10804 4254 -10770
rect 4196 -10875 4254 -10804
rect 4288 -10657 4626 -10587
rect 4660 -10589 4990 -10519
rect 4660 -10623 4680 -10589
rect 4714 -10623 4779 -10589
rect 4813 -10623 4878 -10589
rect 4912 -10623 4990 -10589
rect 5116 -10587 5136 -10553
rect 5170 -10587 5266 -10553
rect 4288 -10697 4990 -10657
rect 4288 -10731 4306 -10697
rect 4340 -10731 4938 -10697
rect 4972 -10731 4990 -10697
rect 4288 -10799 4990 -10731
rect 4288 -10833 4306 -10799
rect 4340 -10833 4938 -10799
rect 4972 -10833 4990 -10799
rect 4288 -10875 4990 -10833
rect 5024 -10677 5082 -10642
rect 5024 -10711 5036 -10677
rect 5070 -10711 5082 -10677
rect 5024 -10770 5082 -10711
rect 5024 -10804 5036 -10770
rect 5070 -10804 5082 -10770
rect 5024 -10875 5082 -10804
rect 5116 -10657 5266 -10587
rect 5300 -10589 5450 -10519
rect 5300 -10623 5396 -10589
rect 5430 -10623 5450 -10589
rect 5576 -10569 5626 -10476
rect 5847 -10494 5897 -10452
rect 5779 -10528 5897 -10494
rect 5949 -10418 6019 -10399
rect 5949 -10452 5968 -10418
rect 6002 -10452 6019 -10418
rect 5779 -10547 5813 -10528
rect 5576 -10603 5590 -10569
rect 5624 -10603 5626 -10569
rect 5116 -10697 5450 -10657
rect 5116 -10731 5134 -10697
rect 5168 -10731 5398 -10697
rect 5432 -10731 5450 -10697
rect 5116 -10799 5450 -10731
rect 5116 -10833 5134 -10799
rect 5168 -10833 5398 -10799
rect 5432 -10833 5450 -10799
rect 5116 -10875 5450 -10833
rect 5484 -10677 5542 -10642
rect 5484 -10711 5496 -10677
rect 5530 -10711 5542 -10677
rect 5484 -10770 5542 -10711
rect 5484 -10804 5496 -10770
rect 5530 -10804 5542 -10770
rect 5484 -10875 5542 -10804
rect 5576 -10686 5626 -10603
rect 5660 -10563 5813 -10547
rect 5949 -10562 6019 -10452
rect 6112 -10418 6178 -10365
rect 6112 -10452 6128 -10418
rect 6162 -10452 6178 -10418
rect 6112 -10461 6178 -10452
rect 6212 -10418 6278 -10399
rect 6212 -10452 6225 -10418
rect 6259 -10452 6278 -10418
rect 6212 -10495 6278 -10452
rect 6084 -10529 6278 -10495
rect 6312 -10459 6370 -10365
rect 6312 -10493 6324 -10459
rect 6358 -10493 6370 -10459
rect 6312 -10510 6370 -10493
rect 6404 -10433 6738 -10365
rect 6404 -10467 6422 -10433
rect 6456 -10467 6686 -10433
rect 6720 -10467 6738 -10433
rect 6404 -10519 6738 -10467
rect 6772 -10459 6830 -10365
rect 6772 -10493 6784 -10459
rect 6818 -10493 6830 -10459
rect 6772 -10510 6830 -10493
rect 6864 -10426 7566 -10365
rect 6864 -10460 6882 -10426
rect 6916 -10460 7514 -10426
rect 7548 -10460 7566 -10426
rect 6864 -10519 7566 -10460
rect 7600 -10459 7658 -10365
rect 7600 -10493 7612 -10459
rect 7646 -10493 7658 -10459
rect 7600 -10510 7658 -10493
rect 7692 -10433 8026 -10365
rect 7692 -10467 7710 -10433
rect 7744 -10467 7974 -10433
rect 8008 -10467 8026 -10433
rect 7692 -10519 8026 -10467
rect 8060 -10459 8118 -10365
rect 8060 -10493 8072 -10459
rect 8106 -10493 8118 -10459
rect 8060 -10510 8118 -10493
rect 8152 -10418 8233 -10399
rect 8152 -10452 8185 -10418
rect 8219 -10452 8233 -10418
rect 8152 -10476 8233 -10452
rect 8267 -10418 8333 -10365
rect 8267 -10452 8283 -10418
rect 8317 -10452 8333 -10418
rect 8267 -10468 8333 -10452
rect 8423 -10418 8473 -10399
rect 8423 -10452 8439 -10418
rect 6084 -10553 6154 -10529
rect 5660 -10597 5663 -10563
rect 5697 -10597 5813 -10563
rect 5660 -10613 5813 -10597
rect 5847 -10563 6019 -10562
rect 5847 -10597 5863 -10563
rect 5897 -10597 6019 -10563
rect 5847 -10612 6019 -10597
rect 6068 -10563 6154 -10553
rect 6068 -10597 6084 -10563
rect 6118 -10597 6154 -10563
rect 6068 -10611 6154 -10597
rect 6188 -10603 6204 -10563
rect 6238 -10603 6278 -10563
rect 6188 -10606 6278 -10603
rect 6404 -10587 6424 -10553
rect 6458 -10587 6554 -10553
rect 5779 -10647 5813 -10613
rect 5779 -10681 5897 -10647
rect 5576 -10723 5657 -10686
rect 5576 -10757 5609 -10723
rect 5643 -10757 5657 -10723
rect 5576 -10791 5657 -10757
rect 5576 -10825 5609 -10791
rect 5643 -10825 5657 -10791
rect 5576 -10841 5657 -10825
rect 5691 -10724 5757 -10715
rect 5691 -10758 5707 -10724
rect 5741 -10758 5757 -10724
rect 5691 -10792 5757 -10758
rect 5691 -10826 5707 -10792
rect 5741 -10826 5757 -10792
rect 5691 -10875 5757 -10826
rect 5847 -10723 5897 -10681
rect 5847 -10757 5863 -10723
rect 5847 -10791 5897 -10757
rect 5847 -10825 5863 -10791
rect 5847 -10841 5897 -10825
rect 5949 -10724 6019 -10612
rect 6084 -10640 6154 -10611
rect 6084 -10674 6278 -10640
rect 5949 -10758 5967 -10724
rect 6001 -10758 6019 -10724
rect 5949 -10792 6019 -10758
rect 5949 -10826 5967 -10792
rect 6001 -10826 6019 -10792
rect 5949 -10841 6019 -10826
rect 6109 -10724 6175 -10708
rect 6109 -10758 6125 -10724
rect 6159 -10758 6175 -10724
rect 6109 -10792 6175 -10758
rect 6109 -10826 6125 -10792
rect 6159 -10826 6175 -10792
rect 6109 -10875 6175 -10826
rect 6209 -10724 6278 -10674
rect 6209 -10758 6225 -10724
rect 6259 -10758 6278 -10724
rect 6209 -10792 6278 -10758
rect 6209 -10826 6225 -10792
rect 6259 -10826 6278 -10792
rect 6209 -10841 6278 -10826
rect 6312 -10677 6370 -10642
rect 6312 -10711 6324 -10677
rect 6358 -10711 6370 -10677
rect 6312 -10770 6370 -10711
rect 6312 -10804 6324 -10770
rect 6358 -10804 6370 -10770
rect 6312 -10875 6370 -10804
rect 6404 -10657 6554 -10587
rect 6588 -10589 6738 -10519
rect 6588 -10623 6684 -10589
rect 6718 -10623 6738 -10589
rect 6864 -10587 6942 -10553
rect 6976 -10587 7045 -10553
rect 7079 -10587 7148 -10553
rect 7182 -10587 7202 -10553
rect 6404 -10697 6738 -10657
rect 6404 -10731 6422 -10697
rect 6456 -10731 6686 -10697
rect 6720 -10731 6738 -10697
rect 6404 -10799 6738 -10731
rect 6404 -10833 6422 -10799
rect 6456 -10833 6686 -10799
rect 6720 -10833 6738 -10799
rect 6404 -10875 6738 -10833
rect 6772 -10677 6830 -10642
rect 6772 -10711 6784 -10677
rect 6818 -10711 6830 -10677
rect 6772 -10770 6830 -10711
rect 6772 -10804 6784 -10770
rect 6818 -10804 6830 -10770
rect 6772 -10875 6830 -10804
rect 6864 -10657 7202 -10587
rect 7236 -10589 7566 -10519
rect 7236 -10623 7256 -10589
rect 7290 -10623 7355 -10589
rect 7389 -10623 7454 -10589
rect 7488 -10623 7566 -10589
rect 7692 -10587 7712 -10553
rect 7746 -10587 7842 -10553
rect 6864 -10697 7566 -10657
rect 6864 -10731 6882 -10697
rect 6916 -10731 7514 -10697
rect 7548 -10731 7566 -10697
rect 6864 -10799 7566 -10731
rect 6864 -10833 6882 -10799
rect 6916 -10833 7514 -10799
rect 7548 -10833 7566 -10799
rect 6864 -10875 7566 -10833
rect 7600 -10677 7658 -10642
rect 7600 -10711 7612 -10677
rect 7646 -10711 7658 -10677
rect 7600 -10770 7658 -10711
rect 7600 -10804 7612 -10770
rect 7646 -10804 7658 -10770
rect 7600 -10875 7658 -10804
rect 7692 -10657 7842 -10587
rect 7876 -10589 8026 -10519
rect 7876 -10623 7972 -10589
rect 8006 -10623 8026 -10589
rect 8152 -10569 8202 -10476
rect 8423 -10494 8473 -10452
rect 8355 -10528 8473 -10494
rect 8525 -10418 8595 -10399
rect 8525 -10452 8544 -10418
rect 8578 -10452 8595 -10418
rect 8355 -10547 8389 -10528
rect 8152 -10603 8164 -10569
rect 8198 -10603 8202 -10569
rect 7692 -10697 8026 -10657
rect 7692 -10731 7710 -10697
rect 7744 -10731 7974 -10697
rect 8008 -10731 8026 -10697
rect 7692 -10799 8026 -10731
rect 7692 -10833 7710 -10799
rect 7744 -10833 7974 -10799
rect 8008 -10833 8026 -10799
rect 7692 -10875 8026 -10833
rect 8060 -10677 8118 -10642
rect 8060 -10711 8072 -10677
rect 8106 -10711 8118 -10677
rect 8060 -10770 8118 -10711
rect 8060 -10804 8072 -10770
rect 8106 -10804 8118 -10770
rect 8060 -10875 8118 -10804
rect 8152 -10686 8202 -10603
rect 8236 -10563 8389 -10547
rect 8525 -10562 8595 -10452
rect 8688 -10418 8754 -10365
rect 8688 -10452 8704 -10418
rect 8738 -10452 8754 -10418
rect 8688 -10461 8754 -10452
rect 8788 -10418 8854 -10399
rect 8788 -10452 8801 -10418
rect 8835 -10452 8854 -10418
rect 8788 -10495 8854 -10452
rect 8660 -10529 8854 -10495
rect 8888 -10459 8946 -10365
rect 8888 -10493 8900 -10459
rect 8934 -10493 8946 -10459
rect 8888 -10510 8946 -10493
rect 8980 -10433 9314 -10365
rect 8980 -10467 8998 -10433
rect 9032 -10467 9262 -10433
rect 9296 -10467 9314 -10433
rect 8980 -10519 9314 -10467
rect 9348 -10459 9406 -10365
rect 9348 -10493 9360 -10459
rect 9394 -10493 9406 -10459
rect 9348 -10510 9406 -10493
rect 9440 -10426 10142 -10365
rect 9440 -10460 9458 -10426
rect 9492 -10460 10090 -10426
rect 10124 -10460 10142 -10426
rect 9440 -10519 10142 -10460
rect 10176 -10459 10234 -10365
rect 10176 -10493 10188 -10459
rect 10222 -10493 10234 -10459
rect 10176 -10510 10234 -10493
rect 10360 -10433 10694 -10365
rect 10360 -10467 10378 -10433
rect 10412 -10467 10642 -10433
rect 10676 -10467 10694 -10433
rect 10360 -10519 10694 -10467
rect 8660 -10553 8730 -10529
rect 8236 -10597 8239 -10563
rect 8273 -10597 8389 -10563
rect 8236 -10613 8389 -10597
rect 8423 -10563 8595 -10562
rect 8423 -10597 8439 -10563
rect 8473 -10597 8595 -10563
rect 8423 -10612 8595 -10597
rect 8644 -10563 8730 -10553
rect 8644 -10597 8660 -10563
rect 8694 -10597 8730 -10563
rect 8644 -10611 8730 -10597
rect 8764 -10569 8780 -10563
rect 8764 -10603 8778 -10569
rect 8814 -10597 8854 -10563
rect 8812 -10603 8854 -10597
rect 8764 -10606 8854 -10603
rect 8980 -10587 9000 -10553
rect 9034 -10587 9130 -10553
rect 8355 -10647 8389 -10613
rect 8355 -10681 8473 -10647
rect 8152 -10723 8233 -10686
rect 8152 -10757 8185 -10723
rect 8219 -10757 8233 -10723
rect 8152 -10791 8233 -10757
rect 8152 -10825 8185 -10791
rect 8219 -10825 8233 -10791
rect 8152 -10841 8233 -10825
rect 8267 -10724 8333 -10715
rect 8267 -10758 8283 -10724
rect 8317 -10758 8333 -10724
rect 8267 -10792 8333 -10758
rect 8267 -10826 8283 -10792
rect 8317 -10826 8333 -10792
rect 8267 -10875 8333 -10826
rect 8423 -10723 8473 -10681
rect 8423 -10757 8439 -10723
rect 8423 -10791 8473 -10757
rect 8423 -10825 8439 -10791
rect 8423 -10841 8473 -10825
rect 8525 -10724 8595 -10612
rect 8660 -10640 8730 -10611
rect 8660 -10674 8854 -10640
rect 8525 -10758 8543 -10724
rect 8577 -10758 8595 -10724
rect 8525 -10792 8595 -10758
rect 8525 -10826 8543 -10792
rect 8577 -10826 8595 -10792
rect 8525 -10841 8595 -10826
rect 8685 -10724 8751 -10708
rect 8685 -10758 8701 -10724
rect 8735 -10758 8751 -10724
rect 8685 -10792 8751 -10758
rect 8685 -10826 8701 -10792
rect 8735 -10826 8751 -10792
rect 8685 -10875 8751 -10826
rect 8785 -10724 8854 -10674
rect 8785 -10758 8801 -10724
rect 8835 -10758 8854 -10724
rect 8785 -10792 8854 -10758
rect 8785 -10826 8801 -10792
rect 8835 -10826 8854 -10792
rect 8785 -10841 8854 -10826
rect 8888 -10677 8946 -10642
rect 8888 -10711 8900 -10677
rect 8934 -10711 8946 -10677
rect 8888 -10770 8946 -10711
rect 8888 -10804 8900 -10770
rect 8934 -10804 8946 -10770
rect 8888 -10875 8946 -10804
rect 8980 -10657 9130 -10587
rect 9164 -10589 9314 -10519
rect 9164 -10623 9260 -10589
rect 9294 -10623 9314 -10589
rect 9440 -10587 9518 -10553
rect 9552 -10587 9621 -10553
rect 9655 -10587 9724 -10553
rect 9758 -10587 9778 -10553
rect 8980 -10697 9314 -10657
rect 8980 -10731 8998 -10697
rect 9032 -10731 9262 -10697
rect 9296 -10731 9314 -10697
rect 8980 -10799 9314 -10731
rect 8980 -10833 8998 -10799
rect 9032 -10833 9262 -10799
rect 9296 -10833 9314 -10799
rect 8980 -10875 9314 -10833
rect 9348 -10677 9406 -10642
rect 9348 -10711 9360 -10677
rect 9394 -10711 9406 -10677
rect 9348 -10770 9406 -10711
rect 9348 -10804 9360 -10770
rect 9394 -10804 9406 -10770
rect 9348 -10875 9406 -10804
rect 9440 -10657 9778 -10587
rect 9812 -10589 10142 -10519
rect 9812 -10623 9832 -10589
rect 9866 -10623 9931 -10589
rect 9965 -10623 10030 -10589
rect 10064 -10623 10142 -10589
rect 10360 -10587 10380 -10553
rect 10414 -10587 10510 -10553
rect 9440 -10697 10142 -10657
rect 9440 -10731 9458 -10697
rect 9492 -10731 10090 -10697
rect 10124 -10731 10142 -10697
rect 9440 -10799 10142 -10731
rect 9440 -10833 9458 -10799
rect 9492 -10833 10090 -10799
rect 10124 -10833 10142 -10799
rect 9440 -10875 10142 -10833
rect 10176 -10677 10234 -10642
rect 10176 -10711 10188 -10677
rect 10222 -10711 10234 -10677
rect 10176 -10770 10234 -10711
rect 10176 -10804 10188 -10770
rect 10222 -10804 10234 -10770
rect 10176 -10875 10234 -10804
rect 10360 -10657 10510 -10587
rect 10544 -10589 10694 -10519
rect 10544 -10623 10640 -10589
rect 10674 -10623 10694 -10589
rect 10728 -10418 10809 -10399
rect 10728 -10452 10761 -10418
rect 10795 -10452 10809 -10418
rect 10728 -10476 10809 -10452
rect 10843 -10418 10909 -10365
rect 10843 -10452 10859 -10418
rect 10893 -10452 10909 -10418
rect 10843 -10468 10909 -10452
rect 10999 -10418 11049 -10399
rect 10999 -10452 11015 -10418
rect 10728 -10570 10778 -10476
rect 10999 -10494 11049 -10452
rect 10931 -10528 11049 -10494
rect 11101 -10418 11171 -10399
rect 11101 -10452 11120 -10418
rect 11154 -10452 11171 -10418
rect 10931 -10547 10965 -10528
rect 10728 -10604 10738 -10570
rect 10772 -10604 10778 -10570
rect 10360 -10697 10694 -10657
rect 10360 -10731 10378 -10697
rect 10412 -10731 10642 -10697
rect 10676 -10731 10694 -10697
rect 10360 -10799 10694 -10731
rect 10360 -10833 10378 -10799
rect 10412 -10833 10642 -10799
rect 10676 -10833 10694 -10799
rect 10360 -10875 10694 -10833
rect 10728 -10686 10778 -10604
rect 10812 -10563 10965 -10547
rect 11101 -10562 11171 -10452
rect 11264 -10418 11330 -10365
rect 11264 -10452 11280 -10418
rect 11314 -10452 11330 -10418
rect 11264 -10461 11330 -10452
rect 11364 -10418 11430 -10399
rect 11364 -10452 11377 -10418
rect 11411 -10452 11430 -10418
rect 11364 -10495 11430 -10452
rect 11236 -10529 11430 -10495
rect 11464 -10459 11522 -10365
rect 11464 -10493 11476 -10459
rect 11510 -10493 11522 -10459
rect 11464 -10510 11522 -10493
rect 11648 -10433 11982 -10365
rect 11648 -10467 11666 -10433
rect 11700 -10467 11930 -10433
rect 11964 -10467 11982 -10433
rect 11648 -10519 11982 -10467
rect 13488 -10459 13546 -10365
rect 13488 -10493 13500 -10459
rect 13534 -10493 13546 -10459
rect 13488 -10510 13546 -10493
rect 13581 -10426 14650 -10365
rect 13581 -10460 13598 -10426
rect 13632 -10460 14598 -10426
rect 14632 -10460 14650 -10426
rect 13581 -10519 14650 -10460
rect 14684 -10459 14742 -10365
rect 14684 -10493 14696 -10459
rect 14730 -10493 14742 -10459
rect 14684 -10510 14742 -10493
rect 14777 -10426 15846 -10365
rect 14777 -10460 14794 -10426
rect 14828 -10460 15794 -10426
rect 15828 -10460 15846 -10426
rect 14777 -10519 15846 -10460
rect 15880 -10459 15938 -10365
rect 15880 -10493 15892 -10459
rect 15926 -10493 15938 -10459
rect 15880 -10510 15938 -10493
rect 15972 -10426 16674 -10365
rect 15972 -10460 15990 -10426
rect 16024 -10460 16622 -10426
rect 16656 -10460 16674 -10426
rect 15972 -10519 16674 -10460
rect 11236 -10553 11306 -10529
rect 10812 -10597 10815 -10563
rect 10849 -10597 10965 -10563
rect 10812 -10613 10965 -10597
rect 10999 -10563 11171 -10562
rect 10999 -10597 11015 -10563
rect 11049 -10597 11171 -10563
rect 10999 -10612 11171 -10597
rect 11220 -10563 11306 -10553
rect 11220 -10597 11236 -10563
rect 11270 -10597 11306 -10563
rect 11220 -10611 11306 -10597
rect 11340 -10597 11356 -10563
rect 11390 -10568 11430 -10563
rect 11340 -10602 11384 -10597
rect 11418 -10602 11430 -10568
rect 11340 -10606 11430 -10602
rect 11648 -10587 11668 -10553
rect 11702 -10587 11798 -10553
rect 10931 -10647 10965 -10613
rect 10931 -10681 11049 -10647
rect 10728 -10723 10809 -10686
rect 10728 -10757 10761 -10723
rect 10795 -10757 10809 -10723
rect 10728 -10791 10809 -10757
rect 10728 -10825 10761 -10791
rect 10795 -10825 10809 -10791
rect 10728 -10841 10809 -10825
rect 10843 -10724 10909 -10715
rect 10843 -10758 10859 -10724
rect 10893 -10758 10909 -10724
rect 10843 -10792 10909 -10758
rect 10843 -10826 10859 -10792
rect 10893 -10826 10909 -10792
rect 10843 -10875 10909 -10826
rect 10999 -10723 11049 -10681
rect 10999 -10757 11015 -10723
rect 10999 -10791 11049 -10757
rect 10999 -10825 11015 -10791
rect 10999 -10841 11049 -10825
rect 11101 -10724 11171 -10612
rect 11236 -10640 11306 -10611
rect 11236 -10674 11430 -10640
rect 11101 -10758 11119 -10724
rect 11153 -10758 11171 -10724
rect 11101 -10792 11171 -10758
rect 11101 -10826 11119 -10792
rect 11153 -10826 11171 -10792
rect 11101 -10841 11171 -10826
rect 11261 -10724 11327 -10708
rect 11261 -10758 11277 -10724
rect 11311 -10758 11327 -10724
rect 11261 -10792 11327 -10758
rect 11261 -10826 11277 -10792
rect 11311 -10826 11327 -10792
rect 11261 -10875 11327 -10826
rect 11361 -10724 11430 -10674
rect 11361 -10758 11377 -10724
rect 11411 -10758 11430 -10724
rect 11361 -10792 11430 -10758
rect 11361 -10826 11377 -10792
rect 11411 -10826 11430 -10792
rect 11361 -10841 11430 -10826
rect 11464 -10677 11522 -10642
rect 11464 -10711 11476 -10677
rect 11510 -10711 11522 -10677
rect 11464 -10770 11522 -10711
rect 11464 -10804 11476 -10770
rect 11510 -10804 11522 -10770
rect 11464 -10875 11522 -10804
rect 11648 -10657 11798 -10587
rect 11832 -10589 11982 -10519
rect 11832 -10623 11928 -10589
rect 11962 -10623 11982 -10589
rect 13581 -10587 13662 -10553
rect 13696 -10587 13790 -10553
rect 13824 -10587 13918 -10553
rect 13952 -10587 14046 -10553
rect 14080 -10587 14100 -10553
rect 11648 -10697 11982 -10657
rect 11648 -10731 11666 -10697
rect 11700 -10731 11930 -10697
rect 11964 -10731 11982 -10697
rect 11648 -10799 11982 -10731
rect 11648 -10833 11666 -10799
rect 11700 -10833 11930 -10799
rect 11964 -10833 11982 -10799
rect 11648 -10875 11982 -10833
rect 13488 -10677 13546 -10642
rect 13488 -10711 13500 -10677
rect 13534 -10711 13546 -10677
rect 13488 -10770 13546 -10711
rect 13488 -10804 13500 -10770
rect 13534 -10804 13546 -10770
rect 13488 -10875 13546 -10804
rect 13581 -10657 14100 -10587
rect 14134 -10589 14650 -10519
rect 14134 -10623 14154 -10589
rect 14188 -10623 14282 -10589
rect 14316 -10623 14410 -10589
rect 14444 -10623 14538 -10589
rect 14572 -10623 14650 -10589
rect 14777 -10587 14858 -10553
rect 14892 -10587 14986 -10553
rect 15020 -10587 15114 -10553
rect 15148 -10587 15242 -10553
rect 15276 -10587 15296 -10553
rect 13581 -10697 14650 -10657
rect 13581 -10731 13598 -10697
rect 13632 -10731 14598 -10697
rect 14632 -10731 14650 -10697
rect 13581 -10799 14650 -10731
rect 13581 -10833 13598 -10799
rect 13632 -10833 14598 -10799
rect 14632 -10833 14650 -10799
rect 13581 -10875 14650 -10833
rect 14684 -10677 14742 -10642
rect 14684 -10711 14696 -10677
rect 14730 -10711 14742 -10677
rect 14684 -10770 14742 -10711
rect 14684 -10804 14696 -10770
rect 14730 -10804 14742 -10770
rect 14684 -10875 14742 -10804
rect 14777 -10657 15296 -10587
rect 15330 -10589 15846 -10519
rect 15330 -10623 15350 -10589
rect 15384 -10623 15478 -10589
rect 15512 -10623 15606 -10589
rect 15640 -10623 15734 -10589
rect 15768 -10623 15846 -10589
rect 15972 -10587 16050 -10553
rect 16084 -10587 16153 -10553
rect 16187 -10587 16256 -10553
rect 16290 -10587 16310 -10553
rect 14777 -10697 15846 -10657
rect 14777 -10731 14794 -10697
rect 14828 -10731 15794 -10697
rect 15828 -10731 15846 -10697
rect 14777 -10799 15846 -10731
rect 14777 -10833 14794 -10799
rect 14828 -10833 15794 -10799
rect 15828 -10833 15846 -10799
rect 14777 -10875 15846 -10833
rect 15880 -10677 15938 -10642
rect 15880 -10711 15892 -10677
rect 15926 -10711 15938 -10677
rect 15880 -10770 15938 -10711
rect 15880 -10804 15892 -10770
rect 15926 -10804 15938 -10770
rect 15880 -10875 15938 -10804
rect 15972 -10657 16310 -10587
rect 16344 -10589 16674 -10519
rect 16344 -10623 16364 -10589
rect 16398 -10623 16463 -10589
rect 16497 -10623 16562 -10589
rect 16596 -10623 16674 -10589
rect 15972 -10697 16674 -10657
rect 15972 -10731 15990 -10697
rect 16024 -10731 16622 -10697
rect 16656 -10731 16674 -10697
rect 15972 -10799 16674 -10731
rect 15972 -10833 15990 -10799
rect 16024 -10833 16622 -10799
rect 16656 -10833 16674 -10799
rect 15972 -10875 16674 -10833
rect -2997 -10909 -2968 -10875
rect -2934 -10909 -2876 -10875
rect -2842 -10909 -2784 -10875
rect -2750 -10909 -2692 -10875
rect -2658 -10909 -2600 -10875
rect -2566 -10909 -2508 -10875
rect -2474 -10909 -2416 -10875
rect -2382 -10909 -2324 -10875
rect -2290 -10909 -2232 -10875
rect -2198 -10909 -2140 -10875
rect -2106 -10909 -2048 -10875
rect -2014 -10909 -1956 -10875
rect -1922 -10909 -1864 -10875
rect -1830 -10909 -1772 -10875
rect -1738 -10909 -1680 -10875
rect -1646 -10909 -1588 -10875
rect -1554 -10909 -1496 -10875
rect -1462 -10909 -1404 -10875
rect -1370 -10909 -1312 -10875
rect -1278 -10909 -1220 -10875
rect -1186 -10909 -1128 -10875
rect -1094 -10909 -1036 -10875
rect -1002 -10909 -944 -10875
rect -910 -10909 -852 -10875
rect -818 -10909 -760 -10875
rect -726 -10909 -668 -10875
rect -634 -10909 -576 -10875
rect -542 -10909 -484 -10875
rect -450 -10909 -392 -10875
rect -358 -10909 -300 -10875
rect -266 -10909 -208 -10875
rect -174 -10909 -116 -10875
rect -82 -10909 -24 -10875
rect 10 -10909 68 -10875
rect 102 -10909 160 -10875
rect 194 -10909 252 -10875
rect 286 -10909 344 -10875
rect 378 -10909 436 -10875
rect 470 -10909 528 -10875
rect 562 -10909 620 -10875
rect 654 -10909 712 -10875
rect 746 -10909 804 -10875
rect 838 -10909 896 -10875
rect 930 -10909 988 -10875
rect 1022 -10909 1080 -10875
rect 1114 -10909 1172 -10875
rect 1206 -10909 1264 -10875
rect 1298 -10909 1356 -10875
rect 1390 -10909 1448 -10875
rect 1482 -10909 1540 -10875
rect 1574 -10909 1632 -10875
rect 1666 -10909 1724 -10875
rect 1758 -10909 1816 -10875
rect 1850 -10909 1908 -10875
rect 1942 -10909 2000 -10875
rect 2034 -10909 2092 -10875
rect 2126 -10909 2184 -10875
rect 2218 -10909 2276 -10875
rect 2310 -10909 2368 -10875
rect 2402 -10909 2460 -10875
rect 2494 -10909 2552 -10875
rect 2586 -10909 2644 -10875
rect 2678 -10909 2736 -10875
rect 2770 -10909 2828 -10875
rect 2862 -10909 2920 -10875
rect 2954 -10909 3012 -10875
rect 3046 -10909 3104 -10875
rect 3138 -10909 3196 -10875
rect 3230 -10909 3288 -10875
rect 3322 -10909 3380 -10875
rect 3414 -10909 3472 -10875
rect 3506 -10909 3564 -10875
rect 3598 -10909 3656 -10875
rect 3690 -10909 3748 -10875
rect 3782 -10909 3840 -10875
rect 3874 -10909 3932 -10875
rect 3966 -10909 4024 -10875
rect 4058 -10909 4116 -10875
rect 4150 -10909 4208 -10875
rect 4242 -10909 4300 -10875
rect 4334 -10909 4392 -10875
rect 4426 -10909 4484 -10875
rect 4518 -10909 4576 -10875
rect 4610 -10909 4668 -10875
rect 4702 -10909 4760 -10875
rect 4794 -10909 4852 -10875
rect 4886 -10909 4944 -10875
rect 4978 -10909 5036 -10875
rect 5070 -10909 5128 -10875
rect 5162 -10909 5220 -10875
rect 5254 -10909 5312 -10875
rect 5346 -10909 5404 -10875
rect 5438 -10909 5496 -10875
rect 5530 -10909 5588 -10875
rect 5622 -10909 5680 -10875
rect 5714 -10909 5772 -10875
rect 5806 -10909 5864 -10875
rect 5898 -10909 5956 -10875
rect 5990 -10909 6048 -10875
rect 6082 -10909 6140 -10875
rect 6174 -10909 6232 -10875
rect 6266 -10909 6324 -10875
rect 6358 -10909 6416 -10875
rect 6450 -10909 6508 -10875
rect 6542 -10909 6600 -10875
rect 6634 -10909 6692 -10875
rect 6726 -10909 6784 -10875
rect 6818 -10909 6876 -10875
rect 6910 -10909 6968 -10875
rect 7002 -10909 7060 -10875
rect 7094 -10909 7152 -10875
rect 7186 -10909 7244 -10875
rect 7278 -10909 7336 -10875
rect 7370 -10909 7428 -10875
rect 7462 -10909 7520 -10875
rect 7554 -10909 7612 -10875
rect 7646 -10909 7704 -10875
rect 7738 -10909 7796 -10875
rect 7830 -10909 7888 -10875
rect 7922 -10909 7980 -10875
rect 8014 -10909 8072 -10875
rect 8106 -10909 8164 -10875
rect 8198 -10909 8256 -10875
rect 8290 -10909 8348 -10875
rect 8382 -10909 8440 -10875
rect 8474 -10909 8532 -10875
rect 8566 -10909 8624 -10875
rect 8658 -10909 8716 -10875
rect 8750 -10909 8808 -10875
rect 8842 -10909 8900 -10875
rect 8934 -10909 8992 -10875
rect 9026 -10909 9084 -10875
rect 9118 -10909 9176 -10875
rect 9210 -10909 9268 -10875
rect 9302 -10909 9360 -10875
rect 9394 -10909 9452 -10875
rect 9486 -10909 9544 -10875
rect 9578 -10909 9636 -10875
rect 9670 -10909 9728 -10875
rect 9762 -10909 9820 -10875
rect 9854 -10909 9912 -10875
rect 9946 -10909 10004 -10875
rect 10038 -10909 10096 -10875
rect 10130 -10909 10188 -10875
rect 10222 -10909 10280 -10875
rect 10314 -10909 10372 -10875
rect 10406 -10909 10464 -10875
rect 10498 -10909 10556 -10875
rect 10590 -10909 10648 -10875
rect 10682 -10909 10740 -10875
rect 10774 -10909 10832 -10875
rect 10866 -10909 10924 -10875
rect 10958 -10909 11016 -10875
rect 11050 -10909 11108 -10875
rect 11142 -10909 11200 -10875
rect 11234 -10909 11292 -10875
rect 11326 -10909 11384 -10875
rect 11418 -10909 11476 -10875
rect 11510 -10909 11568 -10875
rect 11602 -10909 11660 -10875
rect 11694 -10909 11752 -10875
rect 11786 -10909 11844 -10875
rect 11878 -10909 11936 -10875
rect 11970 -10909 12028 -10875
rect 12062 -10909 12120 -10875
rect 12154 -10909 12212 -10875
rect 12246 -10909 12304 -10875
rect 12338 -10909 12396 -10875
rect 12430 -10909 12488 -10875
rect 12522 -10909 12580 -10875
rect 12614 -10909 12672 -10875
rect 12706 -10909 12764 -10875
rect 12798 -10909 12856 -10875
rect 12890 -10909 12948 -10875
rect 12982 -10909 13040 -10875
rect 13074 -10909 13132 -10875
rect 13166 -10909 13224 -10875
rect 13258 -10909 13316 -10875
rect 13350 -10909 13408 -10875
rect 13442 -10909 13500 -10875
rect 13534 -10909 13592 -10875
rect 13626 -10909 13684 -10875
rect 13718 -10909 13776 -10875
rect 13810 -10909 13868 -10875
rect 13902 -10909 13960 -10875
rect 13994 -10909 14052 -10875
rect 14086 -10909 14144 -10875
rect 14178 -10909 14236 -10875
rect 14270 -10909 14328 -10875
rect 14362 -10909 14420 -10875
rect 14454 -10909 14512 -10875
rect 14546 -10909 14604 -10875
rect 14638 -10909 14696 -10875
rect 14730 -10909 14788 -10875
rect 14822 -10909 14880 -10875
rect 14914 -10909 14972 -10875
rect 15006 -10909 15064 -10875
rect 15098 -10909 15156 -10875
rect 15190 -10909 15248 -10875
rect 15282 -10909 15340 -10875
rect 15374 -10909 15432 -10875
rect 15466 -10909 15524 -10875
rect 15558 -10909 15616 -10875
rect 15650 -10909 15708 -10875
rect 15742 -10909 15800 -10875
rect 15834 -10909 15892 -10875
rect 15926 -10909 15984 -10875
rect 16018 -10909 16076 -10875
rect 16110 -10909 16168 -10875
rect 16202 -10909 16260 -10875
rect 16294 -10909 16352 -10875
rect 16386 -10909 16444 -10875
rect 16478 -10909 16536 -10875
rect 16570 -10909 16628 -10875
rect 16662 -10909 16691 -10875
rect -2980 -10951 -2278 -10909
rect -2980 -10985 -2962 -10951
rect -2928 -10985 -2330 -10951
rect -2296 -10985 -2278 -10951
rect -2980 -11053 -2278 -10985
rect -2980 -11087 -2962 -11053
rect -2928 -11087 -2330 -11053
rect -2296 -11087 -2278 -11053
rect -2980 -11127 -2278 -11087
rect -2980 -11195 -2902 -11161
rect -2868 -11195 -2803 -11161
rect -2769 -11195 -2704 -11161
rect -2670 -11195 -2650 -11161
rect -2980 -11265 -2650 -11195
rect -2616 -11197 -2278 -11127
rect -2244 -10980 -2186 -10909
rect -2244 -11014 -2232 -10980
rect -2198 -11014 -2186 -10980
rect -2244 -11073 -2186 -11014
rect -2244 -11107 -2232 -11073
rect -2198 -11107 -2186 -11073
rect -2244 -11142 -2186 -11107
rect -1600 -10951 -898 -10909
rect -1600 -10985 -1582 -10951
rect -1548 -10985 -950 -10951
rect -916 -10985 -898 -10951
rect -1600 -11053 -898 -10985
rect -1600 -11087 -1582 -11053
rect -1548 -11087 -950 -11053
rect -916 -11087 -898 -11053
rect -1600 -11127 -898 -11087
rect -864 -10951 -162 -10909
rect -864 -10985 -846 -10951
rect -812 -10985 -214 -10951
rect -180 -10985 -162 -10951
rect -864 -11053 -162 -10985
rect -864 -11087 -846 -11053
rect -812 -11087 -214 -11053
rect -180 -11087 -162 -11053
rect -864 -11127 -162 -11087
rect -128 -10980 -70 -10909
rect -128 -11014 -116 -10980
rect -82 -11014 -70 -10980
rect -128 -11073 -70 -11014
rect -128 -11107 -116 -11073
rect -82 -11107 -70 -11073
rect -2616 -11231 -2596 -11197
rect -2562 -11231 -2493 -11197
rect -2459 -11231 -2390 -11197
rect -2356 -11231 -2278 -11197
rect -1600 -11197 -1262 -11127
rect -1600 -11231 -1522 -11197
rect -1488 -11231 -1419 -11197
rect -1385 -11231 -1316 -11197
rect -1282 -11231 -1262 -11197
rect -1228 -11195 -1208 -11161
rect -1174 -11195 -1109 -11161
rect -1075 -11195 -1010 -11161
rect -976 -11195 -898 -11161
rect -1228 -11265 -898 -11195
rect -864 -11197 -526 -11127
rect -128 -11142 -70 -11107
rect -36 -10951 298 -10909
rect -36 -10985 -18 -10951
rect 16 -10985 246 -10951
rect 280 -10985 298 -10951
rect -36 -11053 298 -10985
rect -36 -11087 -18 -11053
rect 16 -11087 246 -11053
rect 280 -11087 298 -11053
rect -36 -11127 298 -11087
rect 332 -10980 390 -10909
rect 332 -11014 344 -10980
rect 378 -11014 390 -10980
rect 332 -11073 390 -11014
rect 332 -11107 344 -11073
rect 378 -11107 390 -11073
rect -864 -11231 -786 -11197
rect -752 -11231 -683 -11197
rect -649 -11231 -580 -11197
rect -546 -11231 -526 -11197
rect -492 -11195 -472 -11161
rect -438 -11195 -373 -11161
rect -339 -11195 -274 -11161
rect -240 -11195 -162 -11161
rect -492 -11265 -162 -11195
rect -36 -11197 114 -11127
rect 332 -11142 390 -11107
rect 424 -10959 505 -10943
rect 424 -10993 457 -10959
rect 491 -10993 505 -10959
rect 424 -11027 505 -10993
rect 424 -11061 457 -11027
rect 491 -11061 505 -11027
rect 424 -11098 505 -11061
rect 539 -10958 605 -10909
rect 539 -10992 555 -10958
rect 589 -10992 605 -10958
rect 539 -11026 605 -10992
rect 539 -11060 555 -11026
rect 589 -11060 605 -11026
rect 539 -11069 605 -11060
rect 695 -10959 745 -10943
rect 695 -10993 711 -10959
rect 695 -11027 745 -10993
rect 695 -11061 711 -11027
rect 424 -11147 474 -11098
rect 695 -11103 745 -11061
rect -36 -11231 -16 -11197
rect 18 -11231 114 -11197
rect 148 -11195 244 -11161
rect 278 -11195 298 -11161
rect 148 -11265 298 -11195
rect -2980 -11324 -2278 -11265
rect -2980 -11358 -2962 -11324
rect -2928 -11358 -2330 -11324
rect -2296 -11358 -2278 -11324
rect -2980 -11419 -2278 -11358
rect -2244 -11291 -2186 -11274
rect -2244 -11325 -2232 -11291
rect -2198 -11325 -2186 -11291
rect -2244 -11419 -2186 -11325
rect -1600 -11324 -898 -11265
rect -1600 -11358 -1582 -11324
rect -1548 -11358 -950 -11324
rect -916 -11358 -898 -11324
rect -1600 -11419 -898 -11358
rect -864 -11324 -162 -11265
rect -864 -11358 -846 -11324
rect -812 -11358 -214 -11324
rect -180 -11358 -162 -11324
rect -864 -11419 -162 -11358
rect -128 -11291 -70 -11274
rect -128 -11325 -116 -11291
rect -82 -11325 -70 -11291
rect -128 -11419 -70 -11325
rect -36 -11317 298 -11265
rect 424 -11181 432 -11147
rect 466 -11181 474 -11147
rect 627 -11137 745 -11103
rect 797 -10958 867 -10943
rect 797 -10992 815 -10958
rect 849 -10992 867 -10958
rect 797 -11026 867 -10992
rect 797 -11060 815 -11026
rect 849 -11060 867 -11026
rect 627 -11171 661 -11137
rect -36 -11351 -18 -11317
rect 16 -11351 246 -11317
rect 280 -11351 298 -11317
rect -36 -11419 298 -11351
rect 332 -11291 390 -11274
rect 332 -11325 344 -11291
rect 378 -11325 390 -11291
rect 332 -11419 390 -11325
rect 424 -11308 474 -11181
rect 508 -11187 661 -11171
rect 797 -11172 867 -11060
rect 957 -10958 1023 -10909
rect 957 -10992 973 -10958
rect 1007 -10992 1023 -10958
rect 957 -11026 1023 -10992
rect 957 -11060 973 -11026
rect 1007 -11060 1023 -11026
rect 957 -11076 1023 -11060
rect 1057 -10958 1126 -10943
rect 1057 -10992 1073 -10958
rect 1107 -10992 1126 -10958
rect 1057 -11026 1126 -10992
rect 1057 -11060 1073 -11026
rect 1107 -11060 1126 -11026
rect 1057 -11110 1126 -11060
rect 508 -11221 511 -11187
rect 545 -11221 661 -11187
rect 508 -11237 661 -11221
rect 695 -11187 867 -11172
rect 932 -11144 1126 -11110
rect 1160 -10980 1218 -10909
rect 1160 -11014 1172 -10980
rect 1206 -11014 1218 -10980
rect 1160 -11073 1218 -11014
rect 1160 -11107 1172 -11073
rect 1206 -11107 1218 -11073
rect 1160 -11142 1218 -11107
rect 1252 -10951 1586 -10909
rect 1252 -10985 1270 -10951
rect 1304 -10985 1534 -10951
rect 1568 -10985 1586 -10951
rect 1252 -11053 1586 -10985
rect 1252 -11087 1270 -11053
rect 1304 -11087 1534 -11053
rect 1568 -11087 1586 -11053
rect 1252 -11127 1586 -11087
rect 1620 -10980 1678 -10909
rect 1620 -11014 1632 -10980
rect 1666 -11014 1678 -10980
rect 1620 -11073 1678 -11014
rect 1620 -11107 1632 -11073
rect 1666 -11107 1678 -11073
rect 932 -11173 1002 -11144
rect 695 -11221 711 -11187
rect 745 -11221 867 -11187
rect 695 -11222 867 -11221
rect 627 -11256 661 -11237
rect 627 -11290 745 -11256
rect 424 -11332 505 -11308
rect 424 -11366 457 -11332
rect 491 -11366 505 -11332
rect 424 -11385 505 -11366
rect 539 -11332 605 -11316
rect 539 -11366 555 -11332
rect 589 -11366 605 -11332
rect 539 -11419 605 -11366
rect 695 -11332 745 -11290
rect 695 -11366 711 -11332
rect 695 -11385 745 -11366
rect 797 -11332 867 -11222
rect 916 -11187 1002 -11173
rect 916 -11221 932 -11187
rect 966 -11221 1002 -11187
rect 1036 -11184 1126 -11178
rect 1036 -11187 1070 -11184
rect 1036 -11221 1052 -11187
rect 1104 -11218 1126 -11184
rect 1086 -11221 1126 -11218
rect 1252 -11197 1402 -11127
rect 1620 -11142 1678 -11107
rect 1712 -10951 2414 -10909
rect 1712 -10985 1730 -10951
rect 1764 -10985 2362 -10951
rect 2396 -10985 2414 -10951
rect 1712 -11053 2414 -10985
rect 1712 -11087 1730 -11053
rect 1764 -11087 2362 -11053
rect 2396 -11087 2414 -11053
rect 1712 -11127 2414 -11087
rect 916 -11231 1002 -11221
rect 1252 -11231 1272 -11197
rect 1306 -11231 1402 -11197
rect 1436 -11195 1532 -11161
rect 1566 -11195 1586 -11161
rect 932 -11255 1002 -11231
rect 932 -11289 1126 -11255
rect 1436 -11265 1586 -11195
rect 797 -11366 816 -11332
rect 850 -11366 867 -11332
rect 797 -11385 867 -11366
rect 960 -11332 1026 -11323
rect 960 -11366 976 -11332
rect 1010 -11366 1026 -11332
rect 960 -11419 1026 -11366
rect 1060 -11332 1126 -11289
rect 1060 -11366 1073 -11332
rect 1107 -11366 1126 -11332
rect 1060 -11385 1126 -11366
rect 1160 -11291 1218 -11274
rect 1160 -11325 1172 -11291
rect 1206 -11325 1218 -11291
rect 1160 -11419 1218 -11325
rect 1252 -11317 1586 -11265
rect 1712 -11195 1790 -11161
rect 1824 -11195 1889 -11161
rect 1923 -11195 1988 -11161
rect 2022 -11195 2042 -11161
rect 1712 -11265 2042 -11195
rect 2076 -11197 2414 -11127
rect 2448 -10980 2506 -10909
rect 2448 -11014 2460 -10980
rect 2494 -11014 2506 -10980
rect 2448 -11073 2506 -11014
rect 2448 -11107 2460 -11073
rect 2494 -11107 2506 -11073
rect 2448 -11142 2506 -11107
rect 2540 -10951 2874 -10909
rect 2540 -10985 2558 -10951
rect 2592 -10985 2822 -10951
rect 2856 -10985 2874 -10951
rect 2540 -11053 2874 -10985
rect 2540 -11087 2558 -11053
rect 2592 -11087 2822 -11053
rect 2856 -11087 2874 -11053
rect 2540 -11127 2874 -11087
rect 2908 -10980 2966 -10909
rect 2908 -11014 2920 -10980
rect 2954 -11014 2966 -10980
rect 2908 -11073 2966 -11014
rect 2908 -11107 2920 -11073
rect 2954 -11107 2966 -11073
rect 2076 -11231 2096 -11197
rect 2130 -11231 2199 -11197
rect 2233 -11231 2302 -11197
rect 2336 -11231 2414 -11197
rect 2540 -11197 2690 -11127
rect 2908 -11142 2966 -11107
rect 3000 -10959 3081 -10943
rect 3000 -10993 3033 -10959
rect 3067 -10993 3081 -10959
rect 3000 -11027 3081 -10993
rect 3000 -11061 3033 -11027
rect 3067 -11061 3081 -11027
rect 3000 -11098 3081 -11061
rect 3115 -10958 3181 -10909
rect 3115 -10992 3131 -10958
rect 3165 -10992 3181 -10958
rect 3115 -11026 3181 -10992
rect 3115 -11060 3131 -11026
rect 3165 -11060 3181 -11026
rect 3115 -11069 3181 -11060
rect 3271 -10959 3321 -10943
rect 3271 -10993 3287 -10959
rect 3271 -11027 3321 -10993
rect 3271 -11061 3287 -11027
rect 2540 -11231 2560 -11197
rect 2594 -11231 2690 -11197
rect 2724 -11195 2820 -11161
rect 2854 -11195 2874 -11161
rect 2724 -11265 2874 -11195
rect 1252 -11351 1270 -11317
rect 1304 -11351 1534 -11317
rect 1568 -11351 1586 -11317
rect 1252 -11419 1586 -11351
rect 1620 -11291 1678 -11274
rect 1620 -11325 1632 -11291
rect 1666 -11325 1678 -11291
rect 1620 -11419 1678 -11325
rect 1712 -11324 2414 -11265
rect 1712 -11358 1730 -11324
rect 1764 -11358 2362 -11324
rect 2396 -11358 2414 -11324
rect 1712 -11419 2414 -11358
rect 2448 -11291 2506 -11274
rect 2448 -11325 2460 -11291
rect 2494 -11325 2506 -11291
rect 2448 -11419 2506 -11325
rect 2540 -11317 2874 -11265
rect 3000 -11181 3050 -11098
rect 3271 -11103 3321 -11061
rect 3203 -11137 3321 -11103
rect 3373 -10958 3443 -10943
rect 3373 -10992 3391 -10958
rect 3425 -10992 3443 -10958
rect 3373 -11026 3443 -10992
rect 3373 -11060 3391 -11026
rect 3425 -11060 3443 -11026
rect 3203 -11171 3237 -11137
rect 3000 -11215 3016 -11181
rect 2540 -11351 2558 -11317
rect 2592 -11351 2822 -11317
rect 2856 -11351 2874 -11317
rect 2540 -11419 2874 -11351
rect 2908 -11291 2966 -11274
rect 2908 -11325 2920 -11291
rect 2954 -11325 2966 -11291
rect 2908 -11419 2966 -11325
rect 3000 -11308 3050 -11215
rect 3084 -11187 3237 -11171
rect 3373 -11172 3443 -11060
rect 3533 -10958 3599 -10909
rect 3533 -10992 3549 -10958
rect 3583 -10992 3599 -10958
rect 3533 -11026 3599 -10992
rect 3533 -11060 3549 -11026
rect 3583 -11060 3599 -11026
rect 3533 -11076 3599 -11060
rect 3633 -10958 3702 -10943
rect 3633 -10992 3649 -10958
rect 3683 -10992 3702 -10958
rect 3633 -11026 3702 -10992
rect 3633 -11060 3649 -11026
rect 3683 -11060 3702 -11026
rect 3633 -11110 3702 -11060
rect 3084 -11221 3087 -11187
rect 3121 -11221 3237 -11187
rect 3084 -11237 3237 -11221
rect 3271 -11187 3443 -11172
rect 3508 -11144 3702 -11110
rect 3736 -10980 3794 -10909
rect 3736 -11014 3748 -10980
rect 3782 -11014 3794 -10980
rect 3736 -11073 3794 -11014
rect 3736 -11107 3748 -11073
rect 3782 -11107 3794 -11073
rect 3736 -11142 3794 -11107
rect 3828 -10951 4162 -10909
rect 3828 -10985 3846 -10951
rect 3880 -10985 4110 -10951
rect 4144 -10985 4162 -10951
rect 3828 -11053 4162 -10985
rect 3828 -11087 3846 -11053
rect 3880 -11087 4110 -11053
rect 4144 -11087 4162 -11053
rect 3828 -11127 4162 -11087
rect 4196 -10980 4254 -10909
rect 4196 -11014 4208 -10980
rect 4242 -11014 4254 -10980
rect 4196 -11073 4254 -11014
rect 4196 -11107 4208 -11073
rect 4242 -11107 4254 -11073
rect 3508 -11173 3578 -11144
rect 3271 -11221 3287 -11187
rect 3321 -11221 3443 -11187
rect 3271 -11222 3443 -11221
rect 3203 -11256 3237 -11237
rect 3203 -11290 3321 -11256
rect 3000 -11332 3081 -11308
rect 3000 -11366 3033 -11332
rect 3067 -11366 3081 -11332
rect 3000 -11385 3081 -11366
rect 3115 -11332 3181 -11316
rect 3115 -11366 3131 -11332
rect 3165 -11366 3181 -11332
rect 3115 -11419 3181 -11366
rect 3271 -11332 3321 -11290
rect 3271 -11366 3287 -11332
rect 3271 -11385 3321 -11366
rect 3373 -11332 3443 -11222
rect 3492 -11187 3578 -11173
rect 3492 -11221 3508 -11187
rect 3542 -11221 3578 -11187
rect 3612 -11181 3702 -11178
rect 3612 -11187 3630 -11181
rect 3612 -11221 3628 -11187
rect 3664 -11215 3702 -11181
rect 3662 -11221 3702 -11215
rect 3828 -11197 3978 -11127
rect 4196 -11142 4254 -11107
rect 4288 -10951 4990 -10909
rect 4288 -10985 4306 -10951
rect 4340 -10985 4938 -10951
rect 4972 -10985 4990 -10951
rect 4288 -11053 4990 -10985
rect 4288 -11087 4306 -11053
rect 4340 -11087 4938 -11053
rect 4972 -11087 4990 -11053
rect 4288 -11127 4990 -11087
rect 3492 -11231 3578 -11221
rect 3828 -11231 3848 -11197
rect 3882 -11231 3978 -11197
rect 4012 -11195 4108 -11161
rect 4142 -11195 4162 -11161
rect 3508 -11255 3578 -11231
rect 3508 -11289 3702 -11255
rect 4012 -11265 4162 -11195
rect 3373 -11366 3392 -11332
rect 3426 -11366 3443 -11332
rect 3373 -11385 3443 -11366
rect 3536 -11332 3602 -11323
rect 3536 -11366 3552 -11332
rect 3586 -11366 3602 -11332
rect 3536 -11419 3602 -11366
rect 3636 -11332 3702 -11289
rect 3636 -11366 3649 -11332
rect 3683 -11366 3702 -11332
rect 3636 -11385 3702 -11366
rect 3736 -11291 3794 -11274
rect 3736 -11325 3748 -11291
rect 3782 -11325 3794 -11291
rect 3736 -11419 3794 -11325
rect 3828 -11317 4162 -11265
rect 4288 -11195 4366 -11161
rect 4400 -11195 4465 -11161
rect 4499 -11195 4564 -11161
rect 4598 -11195 4618 -11161
rect 4288 -11265 4618 -11195
rect 4652 -11197 4990 -11127
rect 5024 -10980 5082 -10909
rect 5024 -11014 5036 -10980
rect 5070 -11014 5082 -10980
rect 5024 -11073 5082 -11014
rect 5024 -11107 5036 -11073
rect 5070 -11107 5082 -11073
rect 5024 -11142 5082 -11107
rect 5116 -10951 5450 -10909
rect 5116 -10985 5134 -10951
rect 5168 -10985 5398 -10951
rect 5432 -10985 5450 -10951
rect 5116 -11053 5450 -10985
rect 5116 -11087 5134 -11053
rect 5168 -11087 5398 -11053
rect 5432 -11087 5450 -11053
rect 5116 -11127 5450 -11087
rect 5484 -10980 5542 -10909
rect 5484 -11014 5496 -10980
rect 5530 -11014 5542 -10980
rect 5484 -11073 5542 -11014
rect 5484 -11107 5496 -11073
rect 5530 -11107 5542 -11073
rect 4652 -11231 4672 -11197
rect 4706 -11231 4775 -11197
rect 4809 -11231 4878 -11197
rect 4912 -11231 4990 -11197
rect 5116 -11197 5266 -11127
rect 5484 -11142 5542 -11107
rect 5576 -10959 5657 -10943
rect 5576 -10993 5609 -10959
rect 5643 -10993 5657 -10959
rect 5576 -11027 5657 -10993
rect 5576 -11061 5609 -11027
rect 5643 -11061 5657 -11027
rect 5576 -11098 5657 -11061
rect 5691 -10958 5757 -10909
rect 5691 -10992 5707 -10958
rect 5741 -10992 5757 -10958
rect 5691 -11026 5757 -10992
rect 5691 -11060 5707 -11026
rect 5741 -11060 5757 -11026
rect 5691 -11069 5757 -11060
rect 5847 -10959 5897 -10943
rect 5847 -10993 5863 -10959
rect 5847 -11027 5897 -10993
rect 5847 -11061 5863 -11027
rect 5116 -11231 5136 -11197
rect 5170 -11231 5266 -11197
rect 5300 -11195 5396 -11161
rect 5430 -11195 5450 -11161
rect 5300 -11265 5450 -11195
rect 3828 -11351 3846 -11317
rect 3880 -11351 4110 -11317
rect 4144 -11351 4162 -11317
rect 3828 -11419 4162 -11351
rect 4196 -11291 4254 -11274
rect 4196 -11325 4208 -11291
rect 4242 -11325 4254 -11291
rect 4196 -11419 4254 -11325
rect 4288 -11324 4990 -11265
rect 4288 -11358 4306 -11324
rect 4340 -11358 4938 -11324
rect 4972 -11358 4990 -11324
rect 4288 -11419 4990 -11358
rect 5024 -11291 5082 -11274
rect 5024 -11325 5036 -11291
rect 5070 -11325 5082 -11291
rect 5024 -11419 5082 -11325
rect 5116 -11317 5450 -11265
rect 5576 -11181 5626 -11098
rect 5847 -11103 5897 -11061
rect 5779 -11137 5897 -11103
rect 5949 -10958 6019 -10943
rect 5949 -10992 5967 -10958
rect 6001 -10992 6019 -10958
rect 5949 -11026 6019 -10992
rect 5949 -11060 5967 -11026
rect 6001 -11060 6019 -11026
rect 5779 -11171 5813 -11137
rect 5576 -11215 5590 -11181
rect 5624 -11215 5626 -11181
rect 5116 -11351 5134 -11317
rect 5168 -11351 5398 -11317
rect 5432 -11351 5450 -11317
rect 5116 -11419 5450 -11351
rect 5484 -11291 5542 -11274
rect 5484 -11325 5496 -11291
rect 5530 -11325 5542 -11291
rect 5484 -11419 5542 -11325
rect 5576 -11308 5626 -11215
rect 5660 -11187 5813 -11171
rect 5949 -11172 6019 -11060
rect 6109 -10958 6175 -10909
rect 6109 -10992 6125 -10958
rect 6159 -10992 6175 -10958
rect 6109 -11026 6175 -10992
rect 6109 -11060 6125 -11026
rect 6159 -11060 6175 -11026
rect 6109 -11076 6175 -11060
rect 6209 -10958 6278 -10943
rect 6209 -10992 6225 -10958
rect 6259 -10992 6278 -10958
rect 6209 -11026 6278 -10992
rect 6209 -11060 6225 -11026
rect 6259 -11060 6278 -11026
rect 6209 -11110 6278 -11060
rect 5660 -11221 5663 -11187
rect 5697 -11221 5813 -11187
rect 5660 -11237 5813 -11221
rect 5847 -11187 6019 -11172
rect 6084 -11144 6278 -11110
rect 6312 -10980 6370 -10909
rect 6312 -11014 6324 -10980
rect 6358 -11014 6370 -10980
rect 6312 -11073 6370 -11014
rect 6312 -11107 6324 -11073
rect 6358 -11107 6370 -11073
rect 6312 -11142 6370 -11107
rect 6404 -10951 6738 -10909
rect 6404 -10985 6422 -10951
rect 6456 -10985 6686 -10951
rect 6720 -10985 6738 -10951
rect 6404 -11053 6738 -10985
rect 6404 -11087 6422 -11053
rect 6456 -11087 6686 -11053
rect 6720 -11087 6738 -11053
rect 6404 -11127 6738 -11087
rect 6772 -10980 6830 -10909
rect 6772 -11014 6784 -10980
rect 6818 -11014 6830 -10980
rect 6772 -11073 6830 -11014
rect 6772 -11107 6784 -11073
rect 6818 -11107 6830 -11073
rect 6084 -11173 6154 -11144
rect 5847 -11221 5863 -11187
rect 5897 -11221 6019 -11187
rect 5847 -11222 6019 -11221
rect 5779 -11256 5813 -11237
rect 5779 -11290 5897 -11256
rect 5576 -11332 5657 -11308
rect 5576 -11366 5609 -11332
rect 5643 -11366 5657 -11332
rect 5576 -11385 5657 -11366
rect 5691 -11332 5757 -11316
rect 5691 -11366 5707 -11332
rect 5741 -11366 5757 -11332
rect 5691 -11419 5757 -11366
rect 5847 -11332 5897 -11290
rect 5847 -11366 5863 -11332
rect 5847 -11385 5897 -11366
rect 5949 -11332 6019 -11222
rect 6068 -11187 6154 -11173
rect 6068 -11221 6084 -11187
rect 6118 -11221 6154 -11187
rect 6188 -11181 6278 -11178
rect 6188 -11221 6204 -11181
rect 6238 -11221 6278 -11181
rect 6404 -11197 6554 -11127
rect 6772 -11142 6830 -11107
rect 6864 -10951 7566 -10909
rect 6864 -10985 6882 -10951
rect 6916 -10985 7514 -10951
rect 7548 -10985 7566 -10951
rect 6864 -11053 7566 -10985
rect 6864 -11087 6882 -11053
rect 6916 -11087 7514 -11053
rect 7548 -11087 7566 -11053
rect 6864 -11127 7566 -11087
rect 6068 -11231 6154 -11221
rect 6404 -11231 6424 -11197
rect 6458 -11231 6554 -11197
rect 6588 -11195 6684 -11161
rect 6718 -11195 6738 -11161
rect 6084 -11255 6154 -11231
rect 6084 -11289 6278 -11255
rect 6588 -11265 6738 -11195
rect 5949 -11366 5968 -11332
rect 6002 -11366 6019 -11332
rect 5949 -11385 6019 -11366
rect 6112 -11332 6178 -11323
rect 6112 -11366 6128 -11332
rect 6162 -11366 6178 -11332
rect 6112 -11419 6178 -11366
rect 6212 -11332 6278 -11289
rect 6212 -11366 6225 -11332
rect 6259 -11366 6278 -11332
rect 6212 -11385 6278 -11366
rect 6312 -11291 6370 -11274
rect 6312 -11325 6324 -11291
rect 6358 -11325 6370 -11291
rect 6312 -11419 6370 -11325
rect 6404 -11317 6738 -11265
rect 6864 -11195 6942 -11161
rect 6976 -11195 7041 -11161
rect 7075 -11195 7140 -11161
rect 7174 -11195 7194 -11161
rect 6864 -11265 7194 -11195
rect 7228 -11197 7566 -11127
rect 7600 -10980 7658 -10909
rect 7600 -11014 7612 -10980
rect 7646 -11014 7658 -10980
rect 7600 -11073 7658 -11014
rect 7600 -11107 7612 -11073
rect 7646 -11107 7658 -11073
rect 7600 -11142 7658 -11107
rect 7692 -10951 8026 -10909
rect 7692 -10985 7710 -10951
rect 7744 -10985 7974 -10951
rect 8008 -10985 8026 -10951
rect 7692 -11053 8026 -10985
rect 7692 -11087 7710 -11053
rect 7744 -11087 7974 -11053
rect 8008 -11087 8026 -11053
rect 7692 -11127 8026 -11087
rect 8060 -10980 8118 -10909
rect 8060 -11014 8072 -10980
rect 8106 -11014 8118 -10980
rect 8060 -11073 8118 -11014
rect 8060 -11107 8072 -11073
rect 8106 -11107 8118 -11073
rect 7228 -11231 7248 -11197
rect 7282 -11231 7351 -11197
rect 7385 -11231 7454 -11197
rect 7488 -11231 7566 -11197
rect 7692 -11197 7842 -11127
rect 8060 -11142 8118 -11107
rect 8152 -10959 8233 -10943
rect 8152 -10993 8185 -10959
rect 8219 -10993 8233 -10959
rect 8152 -11027 8233 -10993
rect 8152 -11061 8185 -11027
rect 8219 -11061 8233 -11027
rect 8152 -11098 8233 -11061
rect 8267 -10958 8333 -10909
rect 8267 -10992 8283 -10958
rect 8317 -10992 8333 -10958
rect 8267 -11026 8333 -10992
rect 8267 -11060 8283 -11026
rect 8317 -11060 8333 -11026
rect 8267 -11069 8333 -11060
rect 8423 -10959 8473 -10943
rect 8423 -10993 8439 -10959
rect 8423 -11027 8473 -10993
rect 8423 -11061 8439 -11027
rect 7692 -11231 7712 -11197
rect 7746 -11231 7842 -11197
rect 7876 -11195 7972 -11161
rect 8006 -11195 8026 -11161
rect 7876 -11265 8026 -11195
rect 6404 -11351 6422 -11317
rect 6456 -11351 6686 -11317
rect 6720 -11351 6738 -11317
rect 6404 -11419 6738 -11351
rect 6772 -11291 6830 -11274
rect 6772 -11325 6784 -11291
rect 6818 -11325 6830 -11291
rect 6772 -11419 6830 -11325
rect 6864 -11324 7566 -11265
rect 6864 -11358 6882 -11324
rect 6916 -11358 7514 -11324
rect 7548 -11358 7566 -11324
rect 6864 -11419 7566 -11358
rect 7600 -11291 7658 -11274
rect 7600 -11325 7612 -11291
rect 7646 -11325 7658 -11291
rect 7600 -11419 7658 -11325
rect 7692 -11317 8026 -11265
rect 8152 -11181 8202 -11098
rect 8423 -11103 8473 -11061
rect 8355 -11137 8473 -11103
rect 8525 -10958 8595 -10943
rect 8525 -10992 8543 -10958
rect 8577 -10992 8595 -10958
rect 8525 -11026 8595 -10992
rect 8525 -11060 8543 -11026
rect 8577 -11060 8595 -11026
rect 8355 -11171 8389 -11137
rect 8152 -11215 8164 -11181
rect 8198 -11215 8202 -11181
rect 7692 -11351 7710 -11317
rect 7744 -11351 7974 -11317
rect 8008 -11351 8026 -11317
rect 7692 -11419 8026 -11351
rect 8060 -11291 8118 -11274
rect 8060 -11325 8072 -11291
rect 8106 -11325 8118 -11291
rect 8060 -11419 8118 -11325
rect 8152 -11308 8202 -11215
rect 8236 -11187 8389 -11171
rect 8525 -11172 8595 -11060
rect 8685 -10958 8751 -10909
rect 8685 -10992 8701 -10958
rect 8735 -10992 8751 -10958
rect 8685 -11026 8751 -10992
rect 8685 -11060 8701 -11026
rect 8735 -11060 8751 -11026
rect 8685 -11076 8751 -11060
rect 8785 -10958 8854 -10943
rect 8785 -10992 8801 -10958
rect 8835 -10992 8854 -10958
rect 8785 -11026 8854 -10992
rect 8785 -11060 8801 -11026
rect 8835 -11060 8854 -11026
rect 8785 -11110 8854 -11060
rect 8236 -11221 8239 -11187
rect 8273 -11221 8389 -11187
rect 8236 -11237 8389 -11221
rect 8423 -11187 8595 -11172
rect 8660 -11144 8854 -11110
rect 8888 -10980 8946 -10909
rect 8888 -11014 8900 -10980
rect 8934 -11014 8946 -10980
rect 8888 -11073 8946 -11014
rect 8888 -11107 8900 -11073
rect 8934 -11107 8946 -11073
rect 8888 -11142 8946 -11107
rect 8980 -10951 9314 -10909
rect 8980 -10985 8998 -10951
rect 9032 -10985 9262 -10951
rect 9296 -10985 9314 -10951
rect 8980 -11053 9314 -10985
rect 8980 -11087 8998 -11053
rect 9032 -11087 9262 -11053
rect 9296 -11087 9314 -11053
rect 8980 -11127 9314 -11087
rect 9348 -10980 9406 -10909
rect 9348 -11014 9360 -10980
rect 9394 -11014 9406 -10980
rect 9348 -11073 9406 -11014
rect 9348 -11107 9360 -11073
rect 9394 -11107 9406 -11073
rect 8660 -11173 8730 -11144
rect 8423 -11221 8439 -11187
rect 8473 -11221 8595 -11187
rect 8423 -11222 8595 -11221
rect 8355 -11256 8389 -11237
rect 8355 -11290 8473 -11256
rect 8152 -11332 8233 -11308
rect 8152 -11366 8185 -11332
rect 8219 -11366 8233 -11332
rect 8152 -11385 8233 -11366
rect 8267 -11332 8333 -11316
rect 8267 -11366 8283 -11332
rect 8317 -11366 8333 -11332
rect 8267 -11419 8333 -11366
rect 8423 -11332 8473 -11290
rect 8423 -11366 8439 -11332
rect 8423 -11385 8473 -11366
rect 8525 -11332 8595 -11222
rect 8644 -11187 8730 -11173
rect 8644 -11221 8660 -11187
rect 8694 -11221 8730 -11187
rect 8764 -11181 8854 -11178
rect 8764 -11215 8778 -11181
rect 8812 -11187 8854 -11181
rect 8764 -11221 8780 -11215
rect 8814 -11221 8854 -11187
rect 8980 -11197 9130 -11127
rect 9348 -11142 9406 -11107
rect 9440 -10951 10142 -10909
rect 9440 -10985 9458 -10951
rect 9492 -10985 10090 -10951
rect 10124 -10985 10142 -10951
rect 9440 -11053 10142 -10985
rect 9440 -11087 9458 -11053
rect 9492 -11087 10090 -11053
rect 10124 -11087 10142 -11053
rect 9440 -11127 10142 -11087
rect 8644 -11231 8730 -11221
rect 8980 -11231 9000 -11197
rect 9034 -11231 9130 -11197
rect 9164 -11195 9260 -11161
rect 9294 -11195 9314 -11161
rect 8660 -11255 8730 -11231
rect 8660 -11289 8854 -11255
rect 9164 -11265 9314 -11195
rect 8525 -11366 8544 -11332
rect 8578 -11366 8595 -11332
rect 8525 -11385 8595 -11366
rect 8688 -11332 8754 -11323
rect 8688 -11366 8704 -11332
rect 8738 -11366 8754 -11332
rect 8688 -11419 8754 -11366
rect 8788 -11332 8854 -11289
rect 8788 -11366 8801 -11332
rect 8835 -11366 8854 -11332
rect 8788 -11385 8854 -11366
rect 8888 -11291 8946 -11274
rect 8888 -11325 8900 -11291
rect 8934 -11325 8946 -11291
rect 8888 -11419 8946 -11325
rect 8980 -11317 9314 -11265
rect 9440 -11195 9518 -11161
rect 9552 -11195 9617 -11161
rect 9651 -11195 9716 -11161
rect 9750 -11195 9770 -11161
rect 9440 -11265 9770 -11195
rect 9804 -11197 10142 -11127
rect 10176 -10980 10234 -10909
rect 10176 -11014 10188 -10980
rect 10222 -11014 10234 -10980
rect 10176 -11073 10234 -11014
rect 10176 -11107 10188 -11073
rect 10222 -11107 10234 -11073
rect 10176 -11142 10234 -11107
rect 10360 -10951 10694 -10909
rect 10360 -10985 10378 -10951
rect 10412 -10985 10642 -10951
rect 10676 -10985 10694 -10951
rect 10360 -11053 10694 -10985
rect 10360 -11087 10378 -11053
rect 10412 -11087 10642 -11053
rect 10676 -11087 10694 -11053
rect 10360 -11127 10694 -11087
rect 10728 -10959 10809 -10943
rect 10728 -10993 10761 -10959
rect 10795 -10993 10809 -10959
rect 10728 -11027 10809 -10993
rect 10728 -11061 10761 -11027
rect 10795 -11061 10809 -11027
rect 10728 -11098 10809 -11061
rect 10843 -10958 10909 -10909
rect 10843 -10992 10859 -10958
rect 10893 -10992 10909 -10958
rect 10843 -11026 10909 -10992
rect 10843 -11060 10859 -11026
rect 10893 -11060 10909 -11026
rect 10843 -11069 10909 -11060
rect 10999 -10959 11049 -10943
rect 10999 -10993 11015 -10959
rect 10999 -11027 11049 -10993
rect 10999 -11061 11015 -11027
rect 9804 -11231 9824 -11197
rect 9858 -11231 9927 -11197
rect 9961 -11231 10030 -11197
rect 10064 -11231 10142 -11197
rect 10360 -11197 10510 -11127
rect 10360 -11231 10380 -11197
rect 10414 -11231 10510 -11197
rect 10544 -11195 10640 -11161
rect 10674 -11195 10694 -11161
rect 10544 -11265 10694 -11195
rect 8980 -11351 8998 -11317
rect 9032 -11351 9262 -11317
rect 9296 -11351 9314 -11317
rect 8980 -11419 9314 -11351
rect 9348 -11291 9406 -11274
rect 9348 -11325 9360 -11291
rect 9394 -11325 9406 -11291
rect 9348 -11419 9406 -11325
rect 9440 -11324 10142 -11265
rect 9440 -11358 9458 -11324
rect 9492 -11358 10090 -11324
rect 10124 -11358 10142 -11324
rect 9440 -11419 10142 -11358
rect 10176 -11291 10234 -11274
rect 10176 -11325 10188 -11291
rect 10222 -11325 10234 -11291
rect 10176 -11419 10234 -11325
rect 10360 -11317 10694 -11265
rect 10360 -11351 10378 -11317
rect 10412 -11351 10642 -11317
rect 10676 -11351 10694 -11317
rect 10360 -11419 10694 -11351
rect 10728 -11184 10778 -11098
rect 10999 -11103 11049 -11061
rect 10931 -11137 11049 -11103
rect 11101 -10958 11171 -10943
rect 11101 -10992 11119 -10958
rect 11153 -10992 11171 -10958
rect 11101 -11026 11171 -10992
rect 11101 -11060 11119 -11026
rect 11153 -11060 11171 -11026
rect 10931 -11171 10965 -11137
rect 10728 -11218 10735 -11184
rect 10769 -11218 10778 -11184
rect 10728 -11308 10778 -11218
rect 10812 -11187 10965 -11171
rect 11101 -11172 11171 -11060
rect 11261 -10958 11327 -10909
rect 11261 -10992 11277 -10958
rect 11311 -10992 11327 -10958
rect 11261 -11026 11327 -10992
rect 11261 -11060 11277 -11026
rect 11311 -11060 11327 -11026
rect 11261 -11076 11327 -11060
rect 11361 -10958 11430 -10943
rect 11361 -10992 11377 -10958
rect 11411 -10992 11430 -10958
rect 11361 -11026 11430 -10992
rect 11361 -11060 11377 -11026
rect 11411 -11060 11430 -11026
rect 11361 -11110 11430 -11060
rect 10812 -11221 10815 -11187
rect 10849 -11221 10965 -11187
rect 10812 -11237 10965 -11221
rect 10999 -11187 11171 -11172
rect 11236 -11144 11430 -11110
rect 11464 -10980 11522 -10909
rect 11464 -11014 11476 -10980
rect 11510 -11014 11522 -10980
rect 11464 -11073 11522 -11014
rect 11464 -11107 11476 -11073
rect 11510 -11107 11522 -11073
rect 11464 -11142 11522 -11107
rect 11648 -10951 11982 -10909
rect 11648 -10985 11666 -10951
rect 11700 -10985 11930 -10951
rect 11964 -10985 11982 -10951
rect 11648 -11053 11982 -10985
rect 11648 -11087 11666 -11053
rect 11700 -11087 11930 -11053
rect 11964 -11087 11982 -11053
rect 11648 -11127 11982 -11087
rect 13488 -10980 13546 -10909
rect 13488 -11014 13500 -10980
rect 13534 -11014 13546 -10980
rect 13488 -11073 13546 -11014
rect 13488 -11107 13500 -11073
rect 13534 -11107 13546 -11073
rect 11236 -11173 11306 -11144
rect 10999 -11221 11015 -11187
rect 11049 -11221 11171 -11187
rect 10999 -11222 11171 -11221
rect 10931 -11256 10965 -11237
rect 10931 -11290 11049 -11256
rect 10728 -11332 10809 -11308
rect 10728 -11366 10761 -11332
rect 10795 -11366 10809 -11332
rect 10728 -11385 10809 -11366
rect 10843 -11332 10909 -11316
rect 10843 -11366 10859 -11332
rect 10893 -11366 10909 -11332
rect 10843 -11419 10909 -11366
rect 10999 -11332 11049 -11290
rect 10999 -11366 11015 -11332
rect 10999 -11385 11049 -11366
rect 11101 -11332 11171 -11222
rect 11220 -11187 11306 -11173
rect 11220 -11221 11236 -11187
rect 11270 -11221 11306 -11187
rect 11340 -11183 11430 -11178
rect 11340 -11187 11383 -11183
rect 11340 -11221 11356 -11187
rect 11417 -11217 11430 -11183
rect 11390 -11221 11430 -11217
rect 11648 -11197 11798 -11127
rect 13488 -11142 13546 -11107
rect 13581 -10951 14650 -10909
rect 13581 -10985 13598 -10951
rect 13632 -10985 14598 -10951
rect 14632 -10985 14650 -10951
rect 13581 -11053 14650 -10985
rect 13581 -11087 13598 -11053
rect 13632 -11087 14598 -11053
rect 14632 -11087 14650 -11053
rect 13581 -11127 14650 -11087
rect 14684 -10980 14742 -10909
rect 14684 -11014 14696 -10980
rect 14730 -11014 14742 -10980
rect 14684 -11073 14742 -11014
rect 14684 -11107 14696 -11073
rect 14730 -11107 14742 -11073
rect 11220 -11231 11306 -11221
rect 11648 -11231 11668 -11197
rect 11702 -11231 11798 -11197
rect 11832 -11195 11928 -11161
rect 11962 -11195 11982 -11161
rect 11236 -11255 11306 -11231
rect 11236 -11289 11430 -11255
rect 11832 -11265 11982 -11195
rect 13581 -11197 14100 -11127
rect 14684 -11142 14742 -11107
rect 14777 -10951 15846 -10909
rect 14777 -10985 14794 -10951
rect 14828 -10985 15794 -10951
rect 15828 -10985 15846 -10951
rect 14777 -11053 15846 -10985
rect 14777 -11087 14794 -11053
rect 14828 -11087 15794 -11053
rect 15828 -11087 15846 -11053
rect 14777 -11127 15846 -11087
rect 15880 -10980 15938 -10909
rect 15880 -11014 15892 -10980
rect 15926 -11014 15938 -10980
rect 15880 -11073 15938 -11014
rect 15880 -11107 15892 -11073
rect 15926 -11107 15938 -11073
rect 13581 -11231 13662 -11197
rect 13696 -11231 13790 -11197
rect 13824 -11231 13918 -11197
rect 13952 -11231 14046 -11197
rect 14080 -11231 14100 -11197
rect 14134 -11195 14154 -11161
rect 14188 -11195 14282 -11161
rect 14316 -11195 14410 -11161
rect 14444 -11195 14538 -11161
rect 14572 -11195 14650 -11161
rect 14134 -11265 14650 -11195
rect 14777 -11197 15296 -11127
rect 15880 -11142 15938 -11107
rect 15972 -10951 16674 -10909
rect 15972 -10985 15990 -10951
rect 16024 -10985 16622 -10951
rect 16656 -10985 16674 -10951
rect 15972 -11053 16674 -10985
rect 15972 -11087 15990 -11053
rect 16024 -11087 16622 -11053
rect 16656 -11087 16674 -11053
rect 15972 -11127 16674 -11087
rect 14777 -11231 14858 -11197
rect 14892 -11231 14986 -11197
rect 15020 -11231 15114 -11197
rect 15148 -11231 15242 -11197
rect 15276 -11231 15296 -11197
rect 15330 -11195 15350 -11161
rect 15384 -11195 15478 -11161
rect 15512 -11195 15606 -11161
rect 15640 -11195 15734 -11161
rect 15768 -11195 15846 -11161
rect 15330 -11265 15846 -11195
rect 15972 -11197 16310 -11127
rect 15972 -11231 16050 -11197
rect 16084 -11231 16153 -11197
rect 16187 -11231 16256 -11197
rect 16290 -11231 16310 -11197
rect 16344 -11195 16364 -11161
rect 16398 -11195 16463 -11161
rect 16497 -11195 16562 -11161
rect 16596 -11195 16674 -11161
rect 16344 -11265 16674 -11195
rect 11101 -11366 11120 -11332
rect 11154 -11366 11171 -11332
rect 11101 -11385 11171 -11366
rect 11264 -11332 11330 -11323
rect 11264 -11366 11280 -11332
rect 11314 -11366 11330 -11332
rect 11264 -11419 11330 -11366
rect 11364 -11332 11430 -11289
rect 11364 -11366 11377 -11332
rect 11411 -11366 11430 -11332
rect 11364 -11385 11430 -11366
rect 11464 -11291 11522 -11274
rect 11464 -11325 11476 -11291
rect 11510 -11325 11522 -11291
rect 11464 -11419 11522 -11325
rect 11648 -11317 11982 -11265
rect 11648 -11351 11666 -11317
rect 11700 -11351 11930 -11317
rect 11964 -11351 11982 -11317
rect 11648 -11419 11982 -11351
rect 13488 -11291 13546 -11274
rect 13488 -11325 13500 -11291
rect 13534 -11325 13546 -11291
rect 13488 -11419 13546 -11325
rect 13581 -11324 14650 -11265
rect 13581 -11358 13598 -11324
rect 13632 -11358 14598 -11324
rect 14632 -11358 14650 -11324
rect 13581 -11419 14650 -11358
rect 14684 -11291 14742 -11274
rect 14684 -11325 14696 -11291
rect 14730 -11325 14742 -11291
rect 14684 -11419 14742 -11325
rect 14777 -11324 15846 -11265
rect 14777 -11358 14794 -11324
rect 14828 -11358 15794 -11324
rect 15828 -11358 15846 -11324
rect 14777 -11419 15846 -11358
rect 15880 -11291 15938 -11274
rect 15880 -11325 15892 -11291
rect 15926 -11325 15938 -11291
rect 15880 -11419 15938 -11325
rect 15972 -11324 16674 -11265
rect 15972 -11358 15990 -11324
rect 16024 -11358 16622 -11324
rect 16656 -11358 16674 -11324
rect 15972 -11419 16674 -11358
rect -2997 -11453 -2968 -11419
rect -2934 -11453 -2876 -11419
rect -2842 -11453 -2784 -11419
rect -2750 -11453 -2692 -11419
rect -2658 -11453 -2600 -11419
rect -2566 -11453 -2508 -11419
rect -2474 -11453 -2416 -11419
rect -2382 -11453 -2324 -11419
rect -2290 -11453 -2232 -11419
rect -2198 -11453 -2140 -11419
rect -2106 -11453 -2048 -11419
rect -2014 -11453 -1956 -11419
rect -1922 -11453 -1864 -11419
rect -1830 -11453 -1772 -11419
rect -1738 -11453 -1680 -11419
rect -1646 -11453 -1588 -11419
rect -1554 -11453 -1496 -11419
rect -1462 -11453 -1404 -11419
rect -1370 -11453 -1312 -11419
rect -1278 -11453 -1220 -11419
rect -1186 -11453 -1128 -11419
rect -1094 -11453 -1036 -11419
rect -1002 -11453 -944 -11419
rect -910 -11453 -852 -11419
rect -818 -11453 -760 -11419
rect -726 -11453 -668 -11419
rect -634 -11453 -576 -11419
rect -542 -11453 -484 -11419
rect -450 -11453 -392 -11419
rect -358 -11453 -300 -11419
rect -266 -11453 -208 -11419
rect -174 -11453 -116 -11419
rect -82 -11453 -24 -11419
rect 10 -11453 68 -11419
rect 102 -11453 160 -11419
rect 194 -11453 252 -11419
rect 286 -11453 344 -11419
rect 378 -11453 436 -11419
rect 470 -11453 528 -11419
rect 562 -11453 620 -11419
rect 654 -11453 712 -11419
rect 746 -11453 804 -11419
rect 838 -11453 896 -11419
rect 930 -11453 988 -11419
rect 1022 -11453 1080 -11419
rect 1114 -11453 1172 -11419
rect 1206 -11453 1264 -11419
rect 1298 -11453 1356 -11419
rect 1390 -11453 1448 -11419
rect 1482 -11453 1540 -11419
rect 1574 -11453 1632 -11419
rect 1666 -11453 1724 -11419
rect 1758 -11453 1816 -11419
rect 1850 -11453 1908 -11419
rect 1942 -11453 2000 -11419
rect 2034 -11453 2092 -11419
rect 2126 -11453 2184 -11419
rect 2218 -11453 2276 -11419
rect 2310 -11453 2368 -11419
rect 2402 -11453 2460 -11419
rect 2494 -11453 2552 -11419
rect 2586 -11453 2644 -11419
rect 2678 -11453 2736 -11419
rect 2770 -11453 2828 -11419
rect 2862 -11453 2920 -11419
rect 2954 -11453 3012 -11419
rect 3046 -11453 3104 -11419
rect 3138 -11453 3196 -11419
rect 3230 -11453 3288 -11419
rect 3322 -11453 3380 -11419
rect 3414 -11453 3472 -11419
rect 3506 -11453 3564 -11419
rect 3598 -11453 3656 -11419
rect 3690 -11453 3748 -11419
rect 3782 -11453 3840 -11419
rect 3874 -11453 3932 -11419
rect 3966 -11453 4024 -11419
rect 4058 -11453 4116 -11419
rect 4150 -11453 4208 -11419
rect 4242 -11453 4300 -11419
rect 4334 -11453 4392 -11419
rect 4426 -11453 4484 -11419
rect 4518 -11453 4576 -11419
rect 4610 -11453 4668 -11419
rect 4702 -11453 4760 -11419
rect 4794 -11453 4852 -11419
rect 4886 -11453 4944 -11419
rect 4978 -11453 5036 -11419
rect 5070 -11453 5128 -11419
rect 5162 -11453 5220 -11419
rect 5254 -11453 5312 -11419
rect 5346 -11453 5404 -11419
rect 5438 -11453 5496 -11419
rect 5530 -11453 5588 -11419
rect 5622 -11453 5680 -11419
rect 5714 -11453 5772 -11419
rect 5806 -11453 5864 -11419
rect 5898 -11453 5956 -11419
rect 5990 -11453 6048 -11419
rect 6082 -11453 6140 -11419
rect 6174 -11453 6232 -11419
rect 6266 -11453 6324 -11419
rect 6358 -11453 6416 -11419
rect 6450 -11453 6508 -11419
rect 6542 -11453 6600 -11419
rect 6634 -11453 6692 -11419
rect 6726 -11453 6784 -11419
rect 6818 -11453 6876 -11419
rect 6910 -11453 6968 -11419
rect 7002 -11453 7060 -11419
rect 7094 -11453 7152 -11419
rect 7186 -11453 7244 -11419
rect 7278 -11453 7336 -11419
rect 7370 -11453 7428 -11419
rect 7462 -11453 7520 -11419
rect 7554 -11453 7612 -11419
rect 7646 -11453 7704 -11419
rect 7738 -11453 7796 -11419
rect 7830 -11453 7888 -11419
rect 7922 -11453 7980 -11419
rect 8014 -11453 8072 -11419
rect 8106 -11453 8164 -11419
rect 8198 -11453 8256 -11419
rect 8290 -11453 8348 -11419
rect 8382 -11453 8440 -11419
rect 8474 -11453 8532 -11419
rect 8566 -11453 8624 -11419
rect 8658 -11453 8716 -11419
rect 8750 -11453 8808 -11419
rect 8842 -11453 8900 -11419
rect 8934 -11453 8992 -11419
rect 9026 -11453 9084 -11419
rect 9118 -11453 9176 -11419
rect 9210 -11453 9268 -11419
rect 9302 -11453 9360 -11419
rect 9394 -11453 9452 -11419
rect 9486 -11453 9544 -11419
rect 9578 -11453 9636 -11419
rect 9670 -11453 9728 -11419
rect 9762 -11453 9820 -11419
rect 9854 -11453 9912 -11419
rect 9946 -11453 10004 -11419
rect 10038 -11453 10096 -11419
rect 10130 -11453 10188 -11419
rect 10222 -11453 10280 -11419
rect 10314 -11453 10372 -11419
rect 10406 -11453 10464 -11419
rect 10498 -11453 10556 -11419
rect 10590 -11453 10648 -11419
rect 10682 -11453 10740 -11419
rect 10774 -11453 10832 -11419
rect 10866 -11453 10924 -11419
rect 10958 -11453 11016 -11419
rect 11050 -11453 11108 -11419
rect 11142 -11453 11200 -11419
rect 11234 -11453 11292 -11419
rect 11326 -11453 11384 -11419
rect 11418 -11453 11476 -11419
rect 11510 -11453 11568 -11419
rect 11602 -11453 11660 -11419
rect 11694 -11453 11752 -11419
rect 11786 -11453 11844 -11419
rect 11878 -11453 11936 -11419
rect 11970 -11453 12028 -11419
rect 12062 -11453 12120 -11419
rect 12154 -11453 12212 -11419
rect 12246 -11453 12304 -11419
rect 12338 -11453 12396 -11419
rect 12430 -11453 12488 -11419
rect 12522 -11453 12580 -11419
rect 12614 -11453 12672 -11419
rect 12706 -11453 12764 -11419
rect 12798 -11453 12856 -11419
rect 12890 -11453 12948 -11419
rect 12982 -11453 13040 -11419
rect 13074 -11453 13132 -11419
rect 13166 -11453 13224 -11419
rect 13258 -11453 13316 -11419
rect 13350 -11453 13408 -11419
rect 13442 -11453 13500 -11419
rect 13534 -11453 13592 -11419
rect 13626 -11453 13684 -11419
rect 13718 -11453 13776 -11419
rect 13810 -11453 13868 -11419
rect 13902 -11453 13960 -11419
rect 13994 -11453 14052 -11419
rect 14086 -11453 14144 -11419
rect 14178 -11453 14236 -11419
rect 14270 -11453 14328 -11419
rect 14362 -11453 14420 -11419
rect 14454 -11453 14512 -11419
rect 14546 -11453 14604 -11419
rect 14638 -11453 14696 -11419
rect 14730 -11453 14788 -11419
rect 14822 -11453 14880 -11419
rect 14914 -11453 14972 -11419
rect 15006 -11453 15064 -11419
rect 15098 -11453 15156 -11419
rect 15190 -11453 15248 -11419
rect 15282 -11453 15340 -11419
rect 15374 -11453 15432 -11419
rect 15466 -11453 15524 -11419
rect 15558 -11453 15616 -11419
rect 15650 -11453 15708 -11419
rect 15742 -11453 15800 -11419
rect 15834 -11453 15892 -11419
rect 15926 -11453 15984 -11419
rect 16018 -11453 16076 -11419
rect 16110 -11453 16168 -11419
rect 16202 -11453 16260 -11419
rect 16294 -11453 16352 -11419
rect 16386 -11453 16444 -11419
rect 16478 -11453 16536 -11419
rect 16570 -11453 16628 -11419
rect 16662 -11453 16691 -11419
rect -2980 -11514 -2278 -11453
rect -2980 -11548 -2962 -11514
rect -2928 -11548 -2330 -11514
rect -2296 -11548 -2278 -11514
rect -2980 -11607 -2278 -11548
rect -2244 -11547 -2186 -11453
rect -2244 -11581 -2232 -11547
rect -2198 -11581 -2186 -11547
rect -2244 -11598 -2186 -11581
rect -1600 -11514 -898 -11453
rect -1600 -11548 -1582 -11514
rect -1548 -11548 -950 -11514
rect -916 -11548 -898 -11514
rect -2980 -11675 -2902 -11641
rect -2868 -11675 -2799 -11641
rect -2765 -11675 -2696 -11641
rect -2662 -11675 -2642 -11641
rect -2980 -11745 -2642 -11675
rect -2608 -11677 -2278 -11607
rect -2608 -11711 -2588 -11677
rect -2554 -11711 -2489 -11677
rect -2455 -11711 -2390 -11677
rect -2356 -11711 -2278 -11677
rect -1600 -11607 -898 -11548
rect -864 -11514 -162 -11453
rect -864 -11548 -846 -11514
rect -812 -11548 -214 -11514
rect -180 -11548 -162 -11514
rect -864 -11607 -162 -11548
rect -128 -11547 -70 -11453
rect -128 -11581 -116 -11547
rect -82 -11581 -70 -11547
rect -128 -11598 -70 -11581
rect -36 -11521 298 -11453
rect -36 -11555 -18 -11521
rect 16 -11555 246 -11521
rect 280 -11555 298 -11521
rect -36 -11607 298 -11555
rect 332 -11547 390 -11453
rect 332 -11581 344 -11547
rect 378 -11581 390 -11547
rect 332 -11598 390 -11581
rect 424 -11506 490 -11487
rect 424 -11540 443 -11506
rect 477 -11540 490 -11506
rect 424 -11583 490 -11540
rect 524 -11506 590 -11453
rect 524 -11540 540 -11506
rect 574 -11540 590 -11506
rect 524 -11549 590 -11540
rect 683 -11506 753 -11487
rect 683 -11540 700 -11506
rect 734 -11540 753 -11506
rect -1600 -11677 -1270 -11607
rect -1600 -11711 -1522 -11677
rect -1488 -11711 -1423 -11677
rect -1389 -11711 -1324 -11677
rect -1290 -11711 -1270 -11677
rect -1236 -11675 -1216 -11641
rect -1182 -11675 -1113 -11641
rect -1079 -11675 -1010 -11641
rect -976 -11675 -898 -11641
rect -2980 -11785 -2278 -11745
rect -2980 -11819 -2962 -11785
rect -2928 -11819 -2330 -11785
rect -2296 -11819 -2278 -11785
rect -2980 -11887 -2278 -11819
rect -2980 -11921 -2962 -11887
rect -2928 -11921 -2330 -11887
rect -2296 -11921 -2278 -11887
rect -2980 -11963 -2278 -11921
rect -2244 -11765 -2186 -11730
rect -1236 -11745 -898 -11675
rect -864 -11677 -534 -11607
rect -864 -11711 -786 -11677
rect -752 -11711 -687 -11677
rect -653 -11711 -588 -11677
rect -554 -11711 -534 -11677
rect -500 -11675 -480 -11641
rect -446 -11675 -377 -11641
rect -343 -11675 -274 -11641
rect -240 -11675 -162 -11641
rect -500 -11745 -162 -11675
rect -36 -11675 -16 -11641
rect 18 -11675 114 -11641
rect -2244 -11799 -2232 -11765
rect -2198 -11799 -2186 -11765
rect -2244 -11858 -2186 -11799
rect -2244 -11892 -2232 -11858
rect -2198 -11892 -2186 -11858
rect -2244 -11963 -2186 -11892
rect -1600 -11785 -898 -11745
rect -1600 -11819 -1582 -11785
rect -1548 -11819 -950 -11785
rect -916 -11819 -898 -11785
rect -1600 -11887 -898 -11819
rect -1600 -11921 -1582 -11887
rect -1548 -11921 -950 -11887
rect -916 -11921 -898 -11887
rect -1600 -11963 -898 -11921
rect -864 -11785 -162 -11745
rect -864 -11819 -846 -11785
rect -812 -11819 -214 -11785
rect -180 -11819 -162 -11785
rect -864 -11887 -162 -11819
rect -864 -11921 -846 -11887
rect -812 -11921 -214 -11887
rect -180 -11921 -162 -11887
rect -864 -11963 -162 -11921
rect -128 -11765 -70 -11730
rect -128 -11799 -116 -11765
rect -82 -11799 -70 -11765
rect -128 -11858 -70 -11799
rect -128 -11892 -116 -11858
rect -82 -11892 -70 -11858
rect -128 -11963 -70 -11892
rect -36 -11745 114 -11675
rect 148 -11677 298 -11607
rect 424 -11617 618 -11583
rect 548 -11641 618 -11617
rect 548 -11651 634 -11641
rect 148 -11711 244 -11677
rect 278 -11711 298 -11677
rect 424 -11656 464 -11651
rect 424 -11690 436 -11656
rect 498 -11685 514 -11651
rect 470 -11690 514 -11685
rect 424 -11694 514 -11690
rect 548 -11685 584 -11651
rect 618 -11685 634 -11651
rect 548 -11699 634 -11685
rect 683 -11650 753 -11540
rect 805 -11506 855 -11487
rect 839 -11540 855 -11506
rect 805 -11582 855 -11540
rect 945 -11506 1011 -11453
rect 945 -11540 961 -11506
rect 995 -11540 1011 -11506
rect 945 -11556 1011 -11540
rect 1045 -11506 1126 -11487
rect 1045 -11540 1059 -11506
rect 1093 -11540 1126 -11506
rect 1045 -11564 1126 -11540
rect 805 -11616 923 -11582
rect 889 -11635 923 -11616
rect 683 -11651 855 -11650
rect 683 -11685 805 -11651
rect 839 -11685 855 -11651
rect 548 -11728 618 -11699
rect -36 -11785 298 -11745
rect -36 -11819 -18 -11785
rect 16 -11819 246 -11785
rect 280 -11819 298 -11785
rect -36 -11887 298 -11819
rect -36 -11921 -18 -11887
rect 16 -11921 246 -11887
rect 280 -11921 298 -11887
rect -36 -11963 298 -11921
rect 332 -11765 390 -11730
rect 332 -11799 344 -11765
rect 378 -11799 390 -11765
rect 332 -11858 390 -11799
rect 332 -11892 344 -11858
rect 378 -11892 390 -11858
rect 332 -11963 390 -11892
rect 424 -11762 618 -11728
rect 683 -11700 855 -11685
rect 889 -11651 1042 -11635
rect 889 -11685 1005 -11651
rect 1039 -11685 1042 -11651
rect 424 -11812 493 -11762
rect 424 -11846 443 -11812
rect 477 -11846 493 -11812
rect 424 -11880 493 -11846
rect 424 -11914 443 -11880
rect 477 -11914 493 -11880
rect 424 -11929 493 -11914
rect 527 -11812 593 -11796
rect 527 -11846 543 -11812
rect 577 -11846 593 -11812
rect 527 -11880 593 -11846
rect 527 -11914 543 -11880
rect 577 -11914 593 -11880
rect 527 -11963 593 -11914
rect 683 -11812 753 -11700
rect 889 -11701 1042 -11685
rect 1076 -11656 1126 -11564
rect 1160 -11547 1218 -11453
rect 1160 -11581 1172 -11547
rect 1206 -11581 1218 -11547
rect 1160 -11598 1218 -11581
rect 1252 -11521 1586 -11453
rect 1252 -11555 1270 -11521
rect 1304 -11555 1534 -11521
rect 1568 -11555 1586 -11521
rect 1252 -11607 1586 -11555
rect 1620 -11547 1678 -11453
rect 1620 -11581 1632 -11547
rect 1666 -11581 1678 -11547
rect 1620 -11598 1678 -11581
rect 1712 -11514 2414 -11453
rect 1712 -11548 1730 -11514
rect 1764 -11548 2362 -11514
rect 2396 -11548 2414 -11514
rect 1712 -11607 2414 -11548
rect 2448 -11547 2506 -11453
rect 2448 -11581 2460 -11547
rect 2494 -11581 2506 -11547
rect 2448 -11598 2506 -11581
rect 2540 -11521 2874 -11453
rect 2540 -11555 2558 -11521
rect 2592 -11555 2822 -11521
rect 2856 -11555 2874 -11521
rect 2540 -11607 2874 -11555
rect 2908 -11547 2966 -11453
rect 2908 -11581 2920 -11547
rect 2954 -11581 2966 -11547
rect 2908 -11598 2966 -11581
rect 3000 -11506 3066 -11487
rect 3000 -11540 3019 -11506
rect 3053 -11540 3066 -11506
rect 3000 -11583 3066 -11540
rect 3100 -11506 3166 -11453
rect 3100 -11540 3116 -11506
rect 3150 -11540 3166 -11506
rect 3100 -11549 3166 -11540
rect 3259 -11506 3329 -11487
rect 3259 -11540 3276 -11506
rect 3310 -11540 3329 -11506
rect 1076 -11690 1081 -11656
rect 1115 -11690 1126 -11656
rect 889 -11735 923 -11701
rect 683 -11846 701 -11812
rect 735 -11846 753 -11812
rect 683 -11880 753 -11846
rect 683 -11914 701 -11880
rect 735 -11914 753 -11880
rect 683 -11929 753 -11914
rect 805 -11769 923 -11735
rect 805 -11811 855 -11769
rect 1076 -11774 1126 -11690
rect 1252 -11675 1272 -11641
rect 1306 -11675 1402 -11641
rect 839 -11845 855 -11811
rect 805 -11879 855 -11845
rect 839 -11913 855 -11879
rect 805 -11929 855 -11913
rect 945 -11812 1011 -11803
rect 945 -11846 961 -11812
rect 995 -11846 1011 -11812
rect 945 -11880 1011 -11846
rect 945 -11914 961 -11880
rect 995 -11914 1011 -11880
rect 945 -11963 1011 -11914
rect 1045 -11811 1126 -11774
rect 1045 -11845 1059 -11811
rect 1093 -11845 1126 -11811
rect 1045 -11879 1126 -11845
rect 1045 -11913 1059 -11879
rect 1093 -11913 1126 -11879
rect 1045 -11929 1126 -11913
rect 1160 -11765 1218 -11730
rect 1160 -11799 1172 -11765
rect 1206 -11799 1218 -11765
rect 1160 -11858 1218 -11799
rect 1160 -11892 1172 -11858
rect 1206 -11892 1218 -11858
rect 1160 -11963 1218 -11892
rect 1252 -11745 1402 -11675
rect 1436 -11677 1586 -11607
rect 1436 -11711 1532 -11677
rect 1566 -11711 1586 -11677
rect 1712 -11675 1790 -11641
rect 1824 -11675 1893 -11641
rect 1927 -11675 1996 -11641
rect 2030 -11675 2050 -11641
rect 1252 -11785 1586 -11745
rect 1252 -11819 1270 -11785
rect 1304 -11819 1534 -11785
rect 1568 -11819 1586 -11785
rect 1252 -11887 1586 -11819
rect 1252 -11921 1270 -11887
rect 1304 -11921 1534 -11887
rect 1568 -11921 1586 -11887
rect 1252 -11963 1586 -11921
rect 1620 -11765 1678 -11730
rect 1620 -11799 1632 -11765
rect 1666 -11799 1678 -11765
rect 1620 -11858 1678 -11799
rect 1620 -11892 1632 -11858
rect 1666 -11892 1678 -11858
rect 1620 -11963 1678 -11892
rect 1712 -11745 2050 -11675
rect 2084 -11677 2414 -11607
rect 2084 -11711 2104 -11677
rect 2138 -11711 2203 -11677
rect 2237 -11711 2302 -11677
rect 2336 -11711 2414 -11677
rect 2540 -11675 2560 -11641
rect 2594 -11675 2690 -11641
rect 1712 -11785 2414 -11745
rect 1712 -11819 1730 -11785
rect 1764 -11819 2362 -11785
rect 2396 -11819 2414 -11785
rect 1712 -11887 2414 -11819
rect 1712 -11921 1730 -11887
rect 1764 -11921 2362 -11887
rect 2396 -11921 2414 -11887
rect 1712 -11963 2414 -11921
rect 2448 -11765 2506 -11730
rect 2448 -11799 2460 -11765
rect 2494 -11799 2506 -11765
rect 2448 -11858 2506 -11799
rect 2448 -11892 2460 -11858
rect 2494 -11892 2506 -11858
rect 2448 -11963 2506 -11892
rect 2540 -11745 2690 -11675
rect 2724 -11677 2874 -11607
rect 3000 -11617 3194 -11583
rect 3124 -11641 3194 -11617
rect 3124 -11651 3210 -11641
rect 2724 -11711 2820 -11677
rect 2854 -11711 2874 -11677
rect 3000 -11685 3040 -11651
rect 3074 -11656 3090 -11651
rect 3000 -11690 3041 -11685
rect 3075 -11690 3090 -11656
rect 3000 -11694 3090 -11690
rect 3124 -11685 3160 -11651
rect 3194 -11685 3210 -11651
rect 3124 -11699 3210 -11685
rect 3259 -11650 3329 -11540
rect 3381 -11506 3431 -11487
rect 3415 -11540 3431 -11506
rect 3381 -11582 3431 -11540
rect 3521 -11506 3587 -11453
rect 3521 -11540 3537 -11506
rect 3571 -11540 3587 -11506
rect 3521 -11556 3587 -11540
rect 3621 -11506 3702 -11487
rect 3621 -11540 3635 -11506
rect 3669 -11540 3702 -11506
rect 3621 -11564 3702 -11540
rect 3381 -11616 3499 -11582
rect 3465 -11635 3499 -11616
rect 3259 -11651 3431 -11650
rect 3259 -11685 3381 -11651
rect 3415 -11685 3431 -11651
rect 3124 -11728 3194 -11699
rect 2540 -11785 2874 -11745
rect 2540 -11819 2558 -11785
rect 2592 -11819 2822 -11785
rect 2856 -11819 2874 -11785
rect 2540 -11887 2874 -11819
rect 2540 -11921 2558 -11887
rect 2592 -11921 2822 -11887
rect 2856 -11921 2874 -11887
rect 2540 -11963 2874 -11921
rect 2908 -11765 2966 -11730
rect 2908 -11799 2920 -11765
rect 2954 -11799 2966 -11765
rect 2908 -11858 2966 -11799
rect 2908 -11892 2920 -11858
rect 2954 -11892 2966 -11858
rect 2908 -11963 2966 -11892
rect 3000 -11762 3194 -11728
rect 3259 -11700 3431 -11685
rect 3465 -11651 3618 -11635
rect 3465 -11685 3581 -11651
rect 3615 -11685 3618 -11651
rect 3000 -11812 3069 -11762
rect 3000 -11846 3019 -11812
rect 3053 -11846 3069 -11812
rect 3000 -11880 3069 -11846
rect 3000 -11914 3019 -11880
rect 3053 -11914 3069 -11880
rect 3000 -11929 3069 -11914
rect 3103 -11812 3169 -11796
rect 3103 -11846 3119 -11812
rect 3153 -11846 3169 -11812
rect 3103 -11880 3169 -11846
rect 3103 -11914 3119 -11880
rect 3153 -11914 3169 -11880
rect 3103 -11963 3169 -11914
rect 3259 -11812 3329 -11700
rect 3465 -11701 3618 -11685
rect 3652 -11656 3702 -11564
rect 3736 -11547 3794 -11453
rect 3736 -11581 3748 -11547
rect 3782 -11581 3794 -11547
rect 3736 -11598 3794 -11581
rect 3828 -11521 4162 -11453
rect 3828 -11555 3846 -11521
rect 3880 -11555 4110 -11521
rect 4144 -11555 4162 -11521
rect 3828 -11607 4162 -11555
rect 4196 -11547 4254 -11453
rect 4196 -11581 4208 -11547
rect 4242 -11581 4254 -11547
rect 4196 -11598 4254 -11581
rect 4288 -11514 4990 -11453
rect 4288 -11548 4306 -11514
rect 4340 -11548 4938 -11514
rect 4972 -11548 4990 -11514
rect 4288 -11607 4990 -11548
rect 5024 -11547 5082 -11453
rect 5024 -11581 5036 -11547
rect 5070 -11581 5082 -11547
rect 5024 -11598 5082 -11581
rect 5116 -11521 5450 -11453
rect 5116 -11555 5134 -11521
rect 5168 -11555 5398 -11521
rect 5432 -11555 5450 -11521
rect 5116 -11607 5450 -11555
rect 5484 -11547 5542 -11453
rect 5484 -11581 5496 -11547
rect 5530 -11581 5542 -11547
rect 5484 -11598 5542 -11581
rect 5576 -11506 5642 -11487
rect 5576 -11540 5595 -11506
rect 5629 -11540 5642 -11506
rect 5576 -11583 5642 -11540
rect 5676 -11506 5742 -11453
rect 5676 -11540 5692 -11506
rect 5726 -11540 5742 -11506
rect 5676 -11549 5742 -11540
rect 5835 -11506 5905 -11487
rect 5835 -11540 5852 -11506
rect 5886 -11540 5905 -11506
rect 3652 -11690 3655 -11656
rect 3689 -11690 3702 -11656
rect 3465 -11735 3499 -11701
rect 3259 -11846 3277 -11812
rect 3311 -11846 3329 -11812
rect 3259 -11880 3329 -11846
rect 3259 -11914 3277 -11880
rect 3311 -11914 3329 -11880
rect 3259 -11929 3329 -11914
rect 3381 -11769 3499 -11735
rect 3381 -11811 3431 -11769
rect 3652 -11774 3702 -11690
rect 3828 -11675 3848 -11641
rect 3882 -11675 3978 -11641
rect 3415 -11845 3431 -11811
rect 3381 -11879 3431 -11845
rect 3415 -11913 3431 -11879
rect 3381 -11929 3431 -11913
rect 3521 -11812 3587 -11803
rect 3521 -11846 3537 -11812
rect 3571 -11846 3587 -11812
rect 3521 -11880 3587 -11846
rect 3521 -11914 3537 -11880
rect 3571 -11914 3587 -11880
rect 3521 -11963 3587 -11914
rect 3621 -11811 3702 -11774
rect 3621 -11845 3635 -11811
rect 3669 -11845 3702 -11811
rect 3621 -11879 3702 -11845
rect 3621 -11913 3635 -11879
rect 3669 -11913 3702 -11879
rect 3621 -11929 3702 -11913
rect 3736 -11765 3794 -11730
rect 3736 -11799 3748 -11765
rect 3782 -11799 3794 -11765
rect 3736 -11858 3794 -11799
rect 3736 -11892 3748 -11858
rect 3782 -11892 3794 -11858
rect 3736 -11963 3794 -11892
rect 3828 -11745 3978 -11675
rect 4012 -11677 4162 -11607
rect 4012 -11711 4108 -11677
rect 4142 -11711 4162 -11677
rect 4288 -11675 4366 -11641
rect 4400 -11675 4469 -11641
rect 4503 -11675 4572 -11641
rect 4606 -11675 4626 -11641
rect 3828 -11785 4162 -11745
rect 3828 -11819 3846 -11785
rect 3880 -11819 4110 -11785
rect 4144 -11819 4162 -11785
rect 3828 -11887 4162 -11819
rect 3828 -11921 3846 -11887
rect 3880 -11921 4110 -11887
rect 4144 -11921 4162 -11887
rect 3828 -11963 4162 -11921
rect 4196 -11765 4254 -11730
rect 4196 -11799 4208 -11765
rect 4242 -11799 4254 -11765
rect 4196 -11858 4254 -11799
rect 4196 -11892 4208 -11858
rect 4242 -11892 4254 -11858
rect 4196 -11963 4254 -11892
rect 4288 -11745 4626 -11675
rect 4660 -11677 4990 -11607
rect 4660 -11711 4680 -11677
rect 4714 -11711 4779 -11677
rect 4813 -11711 4878 -11677
rect 4912 -11711 4990 -11677
rect 5116 -11675 5136 -11641
rect 5170 -11675 5266 -11641
rect 4288 -11785 4990 -11745
rect 4288 -11819 4306 -11785
rect 4340 -11819 4938 -11785
rect 4972 -11819 4990 -11785
rect 4288 -11887 4990 -11819
rect 4288 -11921 4306 -11887
rect 4340 -11921 4938 -11887
rect 4972 -11921 4990 -11887
rect 4288 -11963 4990 -11921
rect 5024 -11765 5082 -11730
rect 5024 -11799 5036 -11765
rect 5070 -11799 5082 -11765
rect 5024 -11858 5082 -11799
rect 5024 -11892 5036 -11858
rect 5070 -11892 5082 -11858
rect 5024 -11963 5082 -11892
rect 5116 -11745 5266 -11675
rect 5300 -11677 5450 -11607
rect 5576 -11617 5770 -11583
rect 5700 -11641 5770 -11617
rect 5700 -11651 5786 -11641
rect 5300 -11711 5396 -11677
rect 5430 -11711 5450 -11677
rect 5576 -11656 5616 -11651
rect 5576 -11690 5615 -11656
rect 5650 -11685 5666 -11651
rect 5649 -11690 5666 -11685
rect 5576 -11694 5666 -11690
rect 5700 -11685 5736 -11651
rect 5770 -11685 5786 -11651
rect 5700 -11699 5786 -11685
rect 5835 -11650 5905 -11540
rect 5957 -11506 6007 -11487
rect 5991 -11540 6007 -11506
rect 5957 -11582 6007 -11540
rect 6097 -11506 6163 -11453
rect 6097 -11540 6113 -11506
rect 6147 -11540 6163 -11506
rect 6097 -11556 6163 -11540
rect 6197 -11506 6278 -11487
rect 6197 -11540 6211 -11506
rect 6245 -11540 6278 -11506
rect 6197 -11564 6278 -11540
rect 5957 -11616 6075 -11582
rect 6041 -11635 6075 -11616
rect 5835 -11651 6007 -11650
rect 5835 -11685 5957 -11651
rect 5991 -11685 6007 -11651
rect 5700 -11728 5770 -11699
rect 5116 -11785 5450 -11745
rect 5116 -11819 5134 -11785
rect 5168 -11819 5398 -11785
rect 5432 -11819 5450 -11785
rect 5116 -11887 5450 -11819
rect 5116 -11921 5134 -11887
rect 5168 -11921 5398 -11887
rect 5432 -11921 5450 -11887
rect 5116 -11963 5450 -11921
rect 5484 -11765 5542 -11730
rect 5484 -11799 5496 -11765
rect 5530 -11799 5542 -11765
rect 5484 -11858 5542 -11799
rect 5484 -11892 5496 -11858
rect 5530 -11892 5542 -11858
rect 5484 -11963 5542 -11892
rect 5576 -11762 5770 -11728
rect 5835 -11700 6007 -11685
rect 6041 -11651 6194 -11635
rect 6041 -11685 6157 -11651
rect 6191 -11685 6194 -11651
rect 5576 -11812 5645 -11762
rect 5576 -11846 5595 -11812
rect 5629 -11846 5645 -11812
rect 5576 -11880 5645 -11846
rect 5576 -11914 5595 -11880
rect 5629 -11914 5645 -11880
rect 5576 -11929 5645 -11914
rect 5679 -11812 5745 -11796
rect 5679 -11846 5695 -11812
rect 5729 -11846 5745 -11812
rect 5679 -11880 5745 -11846
rect 5679 -11914 5695 -11880
rect 5729 -11914 5745 -11880
rect 5679 -11963 5745 -11914
rect 5835 -11812 5905 -11700
rect 6041 -11701 6194 -11685
rect 6228 -11656 6278 -11564
rect 6312 -11547 6370 -11453
rect 6312 -11581 6324 -11547
rect 6358 -11581 6370 -11547
rect 6312 -11598 6370 -11581
rect 6404 -11521 6738 -11453
rect 6404 -11555 6422 -11521
rect 6456 -11555 6686 -11521
rect 6720 -11555 6738 -11521
rect 6404 -11607 6738 -11555
rect 6772 -11547 6830 -11453
rect 6772 -11581 6784 -11547
rect 6818 -11581 6830 -11547
rect 6772 -11598 6830 -11581
rect 6864 -11514 7566 -11453
rect 6864 -11548 6882 -11514
rect 6916 -11548 7514 -11514
rect 7548 -11548 7566 -11514
rect 6864 -11607 7566 -11548
rect 7600 -11547 7658 -11453
rect 7600 -11581 7612 -11547
rect 7646 -11581 7658 -11547
rect 7600 -11598 7658 -11581
rect 7692 -11521 8026 -11453
rect 7692 -11555 7710 -11521
rect 7744 -11555 7974 -11521
rect 8008 -11555 8026 -11521
rect 7692 -11607 8026 -11555
rect 8060 -11547 8118 -11453
rect 8060 -11581 8072 -11547
rect 8106 -11581 8118 -11547
rect 8060 -11598 8118 -11581
rect 8152 -11506 8218 -11487
rect 8152 -11540 8171 -11506
rect 8205 -11540 8218 -11506
rect 8152 -11583 8218 -11540
rect 8252 -11506 8318 -11453
rect 8252 -11540 8268 -11506
rect 8302 -11540 8318 -11506
rect 8252 -11549 8318 -11540
rect 8411 -11506 8481 -11487
rect 8411 -11540 8428 -11506
rect 8462 -11540 8481 -11506
rect 6228 -11690 6229 -11656
rect 6263 -11690 6278 -11656
rect 6041 -11735 6075 -11701
rect 5835 -11846 5853 -11812
rect 5887 -11846 5905 -11812
rect 5835 -11880 5905 -11846
rect 5835 -11914 5853 -11880
rect 5887 -11914 5905 -11880
rect 5835 -11929 5905 -11914
rect 5957 -11769 6075 -11735
rect 5957 -11811 6007 -11769
rect 6228 -11774 6278 -11690
rect 6404 -11675 6424 -11641
rect 6458 -11675 6554 -11641
rect 5991 -11845 6007 -11811
rect 5957 -11879 6007 -11845
rect 5991 -11913 6007 -11879
rect 5957 -11929 6007 -11913
rect 6097 -11812 6163 -11803
rect 6097 -11846 6113 -11812
rect 6147 -11846 6163 -11812
rect 6097 -11880 6163 -11846
rect 6097 -11914 6113 -11880
rect 6147 -11914 6163 -11880
rect 6097 -11963 6163 -11914
rect 6197 -11811 6278 -11774
rect 6197 -11845 6211 -11811
rect 6245 -11845 6278 -11811
rect 6197 -11879 6278 -11845
rect 6197 -11913 6211 -11879
rect 6245 -11913 6278 -11879
rect 6197 -11929 6278 -11913
rect 6312 -11765 6370 -11730
rect 6312 -11799 6324 -11765
rect 6358 -11799 6370 -11765
rect 6312 -11858 6370 -11799
rect 6312 -11892 6324 -11858
rect 6358 -11892 6370 -11858
rect 6312 -11963 6370 -11892
rect 6404 -11745 6554 -11675
rect 6588 -11677 6738 -11607
rect 6588 -11711 6684 -11677
rect 6718 -11711 6738 -11677
rect 6864 -11675 6942 -11641
rect 6976 -11675 7045 -11641
rect 7079 -11675 7148 -11641
rect 7182 -11675 7202 -11641
rect 6404 -11785 6738 -11745
rect 6404 -11819 6422 -11785
rect 6456 -11819 6686 -11785
rect 6720 -11819 6738 -11785
rect 6404 -11887 6738 -11819
rect 6404 -11921 6422 -11887
rect 6456 -11921 6686 -11887
rect 6720 -11921 6738 -11887
rect 6404 -11963 6738 -11921
rect 6772 -11765 6830 -11730
rect 6772 -11799 6784 -11765
rect 6818 -11799 6830 -11765
rect 6772 -11858 6830 -11799
rect 6772 -11892 6784 -11858
rect 6818 -11892 6830 -11858
rect 6772 -11963 6830 -11892
rect 6864 -11745 7202 -11675
rect 7236 -11677 7566 -11607
rect 7236 -11711 7256 -11677
rect 7290 -11711 7355 -11677
rect 7389 -11711 7454 -11677
rect 7488 -11711 7566 -11677
rect 7692 -11675 7712 -11641
rect 7746 -11675 7842 -11641
rect 6864 -11785 7566 -11745
rect 6864 -11819 6882 -11785
rect 6916 -11819 7514 -11785
rect 7548 -11819 7566 -11785
rect 6864 -11887 7566 -11819
rect 6864 -11921 6882 -11887
rect 6916 -11921 7514 -11887
rect 7548 -11921 7566 -11887
rect 6864 -11963 7566 -11921
rect 7600 -11765 7658 -11730
rect 7600 -11799 7612 -11765
rect 7646 -11799 7658 -11765
rect 7600 -11858 7658 -11799
rect 7600 -11892 7612 -11858
rect 7646 -11892 7658 -11858
rect 7600 -11963 7658 -11892
rect 7692 -11745 7842 -11675
rect 7876 -11677 8026 -11607
rect 8152 -11617 8346 -11583
rect 8276 -11641 8346 -11617
rect 8276 -11651 8362 -11641
rect 7876 -11711 7972 -11677
rect 8006 -11711 8026 -11677
rect 8152 -11656 8192 -11651
rect 8152 -11690 8189 -11656
rect 8226 -11685 8242 -11651
rect 8223 -11690 8242 -11685
rect 8152 -11694 8242 -11690
rect 8276 -11685 8312 -11651
rect 8346 -11685 8362 -11651
rect 8276 -11699 8362 -11685
rect 8411 -11650 8481 -11540
rect 8533 -11506 8583 -11487
rect 8567 -11540 8583 -11506
rect 8533 -11582 8583 -11540
rect 8673 -11506 8739 -11453
rect 8673 -11540 8689 -11506
rect 8723 -11540 8739 -11506
rect 8673 -11556 8739 -11540
rect 8773 -11506 8854 -11487
rect 8773 -11540 8787 -11506
rect 8821 -11540 8854 -11506
rect 8773 -11564 8854 -11540
rect 8533 -11616 8651 -11582
rect 8617 -11635 8651 -11616
rect 8411 -11651 8583 -11650
rect 8411 -11685 8533 -11651
rect 8567 -11685 8583 -11651
rect 8276 -11728 8346 -11699
rect 7692 -11785 8026 -11745
rect 7692 -11819 7710 -11785
rect 7744 -11819 7974 -11785
rect 8008 -11819 8026 -11785
rect 7692 -11887 8026 -11819
rect 7692 -11921 7710 -11887
rect 7744 -11921 7974 -11887
rect 8008 -11921 8026 -11887
rect 7692 -11963 8026 -11921
rect 8060 -11765 8118 -11730
rect 8060 -11799 8072 -11765
rect 8106 -11799 8118 -11765
rect 8060 -11858 8118 -11799
rect 8060 -11892 8072 -11858
rect 8106 -11892 8118 -11858
rect 8060 -11963 8118 -11892
rect 8152 -11762 8346 -11728
rect 8411 -11700 8583 -11685
rect 8617 -11651 8770 -11635
rect 8617 -11685 8733 -11651
rect 8767 -11685 8770 -11651
rect 8152 -11812 8221 -11762
rect 8152 -11846 8171 -11812
rect 8205 -11846 8221 -11812
rect 8152 -11880 8221 -11846
rect 8152 -11914 8171 -11880
rect 8205 -11914 8221 -11880
rect 8152 -11929 8221 -11914
rect 8255 -11812 8321 -11796
rect 8255 -11846 8271 -11812
rect 8305 -11846 8321 -11812
rect 8255 -11880 8321 -11846
rect 8255 -11914 8271 -11880
rect 8305 -11914 8321 -11880
rect 8255 -11963 8321 -11914
rect 8411 -11812 8481 -11700
rect 8617 -11701 8770 -11685
rect 8804 -11656 8854 -11564
rect 8888 -11547 8946 -11453
rect 8888 -11581 8900 -11547
rect 8934 -11581 8946 -11547
rect 8888 -11598 8946 -11581
rect 8980 -11521 9314 -11453
rect 8980 -11555 8998 -11521
rect 9032 -11555 9262 -11521
rect 9296 -11555 9314 -11521
rect 8980 -11607 9314 -11555
rect 9348 -11547 9406 -11453
rect 9348 -11581 9360 -11547
rect 9394 -11581 9406 -11547
rect 9348 -11598 9406 -11581
rect 9440 -11514 10142 -11453
rect 9440 -11548 9458 -11514
rect 9492 -11548 10090 -11514
rect 10124 -11548 10142 -11514
rect 9440 -11607 10142 -11548
rect 10176 -11547 10234 -11453
rect 10176 -11581 10188 -11547
rect 10222 -11581 10234 -11547
rect 10176 -11598 10234 -11581
rect 10360 -11521 10694 -11453
rect 10360 -11555 10378 -11521
rect 10412 -11555 10642 -11521
rect 10676 -11555 10694 -11521
rect 10360 -11607 10694 -11555
rect 8804 -11690 8806 -11656
rect 8840 -11690 8854 -11656
rect 8617 -11735 8651 -11701
rect 8411 -11846 8429 -11812
rect 8463 -11846 8481 -11812
rect 8411 -11880 8481 -11846
rect 8411 -11914 8429 -11880
rect 8463 -11914 8481 -11880
rect 8411 -11929 8481 -11914
rect 8533 -11769 8651 -11735
rect 8533 -11811 8583 -11769
rect 8804 -11774 8854 -11690
rect 8980 -11675 9000 -11641
rect 9034 -11675 9130 -11641
rect 8567 -11845 8583 -11811
rect 8533 -11879 8583 -11845
rect 8567 -11913 8583 -11879
rect 8533 -11929 8583 -11913
rect 8673 -11812 8739 -11803
rect 8673 -11846 8689 -11812
rect 8723 -11846 8739 -11812
rect 8673 -11880 8739 -11846
rect 8673 -11914 8689 -11880
rect 8723 -11914 8739 -11880
rect 8673 -11963 8739 -11914
rect 8773 -11811 8854 -11774
rect 8773 -11845 8787 -11811
rect 8821 -11845 8854 -11811
rect 8773 -11879 8854 -11845
rect 8773 -11913 8787 -11879
rect 8821 -11913 8854 -11879
rect 8773 -11929 8854 -11913
rect 8888 -11765 8946 -11730
rect 8888 -11799 8900 -11765
rect 8934 -11799 8946 -11765
rect 8888 -11858 8946 -11799
rect 8888 -11892 8900 -11858
rect 8934 -11892 8946 -11858
rect 8888 -11963 8946 -11892
rect 8980 -11745 9130 -11675
rect 9164 -11677 9314 -11607
rect 9164 -11711 9260 -11677
rect 9294 -11711 9314 -11677
rect 9440 -11675 9518 -11641
rect 9552 -11675 9621 -11641
rect 9655 -11675 9724 -11641
rect 9758 -11675 9778 -11641
rect 8980 -11785 9314 -11745
rect 8980 -11819 8998 -11785
rect 9032 -11819 9262 -11785
rect 9296 -11819 9314 -11785
rect 8980 -11887 9314 -11819
rect 8980 -11921 8998 -11887
rect 9032 -11921 9262 -11887
rect 9296 -11921 9314 -11887
rect 8980 -11963 9314 -11921
rect 9348 -11765 9406 -11730
rect 9348 -11799 9360 -11765
rect 9394 -11799 9406 -11765
rect 9348 -11858 9406 -11799
rect 9348 -11892 9360 -11858
rect 9394 -11892 9406 -11858
rect 9348 -11963 9406 -11892
rect 9440 -11745 9778 -11675
rect 9812 -11677 10142 -11607
rect 9812 -11711 9832 -11677
rect 9866 -11711 9931 -11677
rect 9965 -11711 10030 -11677
rect 10064 -11711 10142 -11677
rect 10360 -11675 10380 -11641
rect 10414 -11675 10510 -11641
rect 9440 -11785 10142 -11745
rect 9440 -11819 9458 -11785
rect 9492 -11819 10090 -11785
rect 10124 -11819 10142 -11785
rect 9440 -11887 10142 -11819
rect 9440 -11921 9458 -11887
rect 9492 -11921 10090 -11887
rect 10124 -11921 10142 -11887
rect 9440 -11963 10142 -11921
rect 10176 -11765 10234 -11730
rect 10176 -11799 10188 -11765
rect 10222 -11799 10234 -11765
rect 10176 -11858 10234 -11799
rect 10176 -11892 10188 -11858
rect 10222 -11892 10234 -11858
rect 10176 -11963 10234 -11892
rect 10360 -11745 10510 -11675
rect 10544 -11677 10694 -11607
rect 10728 -11506 10794 -11487
rect 10728 -11540 10747 -11506
rect 10781 -11540 10794 -11506
rect 10728 -11583 10794 -11540
rect 10828 -11506 10894 -11453
rect 10828 -11540 10844 -11506
rect 10878 -11540 10894 -11506
rect 10828 -11549 10894 -11540
rect 10987 -11506 11057 -11487
rect 10987 -11540 11004 -11506
rect 11038 -11540 11057 -11506
rect 10728 -11617 10922 -11583
rect 10852 -11641 10922 -11617
rect 10852 -11651 10938 -11641
rect 10544 -11711 10640 -11677
rect 10674 -11711 10694 -11677
rect 10728 -11656 10768 -11651
rect 10728 -11690 10763 -11656
rect 10802 -11685 10818 -11651
rect 10797 -11690 10818 -11685
rect 10728 -11694 10818 -11690
rect 10852 -11685 10888 -11651
rect 10922 -11685 10938 -11651
rect 10852 -11699 10938 -11685
rect 10987 -11650 11057 -11540
rect 11109 -11506 11159 -11487
rect 11143 -11540 11159 -11506
rect 11109 -11582 11159 -11540
rect 11249 -11506 11315 -11453
rect 11249 -11540 11265 -11506
rect 11299 -11540 11315 -11506
rect 11249 -11556 11315 -11540
rect 11349 -11506 11430 -11487
rect 11349 -11540 11363 -11506
rect 11397 -11540 11430 -11506
rect 11349 -11564 11430 -11540
rect 11109 -11616 11227 -11582
rect 11193 -11635 11227 -11616
rect 10987 -11651 11159 -11650
rect 10987 -11685 11109 -11651
rect 11143 -11685 11159 -11651
rect 10852 -11728 10922 -11699
rect 10360 -11785 10694 -11745
rect 10360 -11819 10378 -11785
rect 10412 -11819 10642 -11785
rect 10676 -11819 10694 -11785
rect 10360 -11887 10694 -11819
rect 10360 -11921 10378 -11887
rect 10412 -11921 10642 -11887
rect 10676 -11921 10694 -11887
rect 10360 -11963 10694 -11921
rect 10728 -11762 10922 -11728
rect 10987 -11700 11159 -11685
rect 11193 -11651 11346 -11635
rect 11193 -11685 11309 -11651
rect 11343 -11685 11346 -11651
rect 10728 -11812 10797 -11762
rect 10728 -11846 10747 -11812
rect 10781 -11846 10797 -11812
rect 10728 -11880 10797 -11846
rect 10728 -11914 10747 -11880
rect 10781 -11914 10797 -11880
rect 10728 -11929 10797 -11914
rect 10831 -11812 10897 -11796
rect 10831 -11846 10847 -11812
rect 10881 -11846 10897 -11812
rect 10831 -11880 10897 -11846
rect 10831 -11914 10847 -11880
rect 10881 -11914 10897 -11880
rect 10831 -11963 10897 -11914
rect 10987 -11812 11057 -11700
rect 11193 -11701 11346 -11685
rect 11380 -11693 11430 -11564
rect 11464 -11547 11522 -11453
rect 11464 -11581 11476 -11547
rect 11510 -11581 11522 -11547
rect 11464 -11598 11522 -11581
rect 11648 -11521 11982 -11453
rect 11648 -11555 11666 -11521
rect 11700 -11555 11930 -11521
rect 11964 -11555 11982 -11521
rect 11648 -11607 11982 -11555
rect 12384 -11547 12442 -11453
rect 12572 -11497 12631 -11453
rect 12572 -11531 12588 -11497
rect 12622 -11531 12631 -11497
rect 12572 -11547 12631 -11531
rect 12665 -11508 12717 -11492
rect 12665 -11542 12674 -11508
rect 12708 -11542 12717 -11508
rect 12384 -11581 12396 -11547
rect 12430 -11581 12442 -11547
rect 12665 -11581 12717 -11542
rect 12751 -11497 12803 -11453
rect 12751 -11531 12760 -11497
rect 12794 -11531 12803 -11497
rect 12751 -11547 12803 -11531
rect 12837 -11508 12888 -11492
rect 12837 -11542 12846 -11508
rect 12880 -11542 12888 -11508
rect 12837 -11581 12888 -11542
rect 12922 -11497 12982 -11453
rect 12922 -11531 12932 -11497
rect 12966 -11531 12982 -11497
rect 12922 -11547 12982 -11531
rect 13120 -11547 13178 -11453
rect 13120 -11581 13132 -11547
rect 13166 -11581 13178 -11547
rect 12384 -11598 12442 -11581
rect 11193 -11735 11227 -11701
rect 10987 -11846 11005 -11812
rect 11039 -11846 11057 -11812
rect 10987 -11880 11057 -11846
rect 10987 -11914 11005 -11880
rect 11039 -11914 11057 -11880
rect 10987 -11929 11057 -11914
rect 11109 -11769 11227 -11735
rect 11380 -11727 11386 -11693
rect 11420 -11727 11430 -11693
rect 11109 -11811 11159 -11769
rect 11380 -11774 11430 -11727
rect 11648 -11675 11668 -11641
rect 11702 -11675 11798 -11641
rect 11143 -11845 11159 -11811
rect 11109 -11879 11159 -11845
rect 11143 -11913 11159 -11879
rect 11109 -11929 11159 -11913
rect 11249 -11812 11315 -11803
rect 11249 -11846 11265 -11812
rect 11299 -11846 11315 -11812
rect 11249 -11880 11315 -11846
rect 11249 -11914 11265 -11880
rect 11299 -11914 11315 -11880
rect 11249 -11963 11315 -11914
rect 11349 -11811 11430 -11774
rect 11349 -11845 11363 -11811
rect 11397 -11845 11430 -11811
rect 11349 -11879 11430 -11845
rect 11349 -11913 11363 -11879
rect 11397 -11913 11430 -11879
rect 11349 -11929 11430 -11913
rect 11464 -11765 11522 -11730
rect 11464 -11799 11476 -11765
rect 11510 -11799 11522 -11765
rect 11464 -11858 11522 -11799
rect 11464 -11892 11476 -11858
rect 11510 -11892 11522 -11858
rect 11464 -11963 11522 -11892
rect 11648 -11745 11798 -11675
rect 11832 -11677 11982 -11607
rect 11832 -11711 11928 -11677
rect 11962 -11711 11982 -11677
rect 12514 -11591 13086 -11581
rect 12514 -11615 13042 -11591
rect 12480 -11653 12514 -11615
rect 13026 -11625 13042 -11615
rect 13076 -11625 13086 -11591
rect 13120 -11598 13178 -11581
rect 13212 -11521 13546 -11453
rect 13212 -11555 13230 -11521
rect 13264 -11555 13494 -11521
rect 13528 -11555 13546 -11521
rect 12480 -11727 12514 -11687
rect 12548 -11651 12991 -11649
rect 12548 -11655 12574 -11651
rect 12548 -11689 12568 -11655
rect 12608 -11685 12642 -11651
rect 12676 -11655 12710 -11651
rect 12693 -11685 12710 -11655
rect 12744 -11655 12778 -11651
rect 12744 -11685 12765 -11655
rect 12812 -11685 12846 -11651
rect 12880 -11657 12914 -11651
rect 12948 -11657 12991 -11651
rect 12892 -11685 12914 -11657
rect 12602 -11689 12659 -11685
rect 12693 -11689 12765 -11685
rect 12799 -11689 12858 -11685
rect 12548 -11691 12858 -11689
rect 12892 -11691 12942 -11685
rect 12976 -11691 12991 -11657
rect 12548 -11694 12991 -11691
rect 13026 -11668 13086 -11625
rect 11648 -11785 11982 -11745
rect 11648 -11819 11666 -11785
rect 11700 -11819 11930 -11785
rect 11964 -11819 11982 -11785
rect 11648 -11887 11982 -11819
rect 11648 -11921 11666 -11887
rect 11700 -11921 11930 -11887
rect 11964 -11921 11982 -11887
rect 11648 -11963 11982 -11921
rect 12384 -11765 12442 -11730
rect 13026 -11702 13039 -11668
rect 13073 -11702 13086 -11668
rect 13026 -11728 13086 -11702
rect 13212 -11607 13546 -11555
rect 13580 -11547 13638 -11453
rect 13580 -11581 13592 -11547
rect 13626 -11581 13638 -11547
rect 13672 -11495 13733 -11453
rect 13672 -11529 13690 -11495
rect 13724 -11529 13733 -11495
rect 13672 -11555 13733 -11529
rect 13769 -11508 13819 -11489
rect 13769 -11542 13776 -11508
rect 13810 -11542 13819 -11508
rect 13580 -11598 13638 -11581
rect 13212 -11677 13362 -11607
rect 13672 -11624 13735 -11589
rect 13212 -11711 13232 -11677
rect 13266 -11711 13362 -11677
rect 13396 -11675 13492 -11641
rect 13526 -11675 13546 -11641
rect 12514 -11761 13086 -11728
rect 12480 -11762 13086 -11761
rect 12384 -11799 12396 -11765
rect 12430 -11799 12442 -11765
rect 12580 -11785 12631 -11762
rect 12384 -11858 12442 -11799
rect 12384 -11892 12396 -11858
rect 12430 -11892 12442 -11858
rect 12384 -11963 12442 -11892
rect 12476 -11812 12545 -11796
rect 12476 -11846 12502 -11812
rect 12536 -11846 12545 -11812
rect 12476 -11880 12545 -11846
rect 12476 -11914 12502 -11880
rect 12536 -11914 12545 -11880
rect 12476 -11963 12545 -11914
rect 12580 -11819 12588 -11785
rect 12622 -11819 12631 -11785
rect 12752 -11785 12803 -11762
rect 12580 -11873 12631 -11819
rect 12580 -11907 12588 -11873
rect 12622 -11907 12631 -11873
rect 12580 -11923 12631 -11907
rect 12665 -11812 12717 -11796
rect 12665 -11846 12674 -11812
rect 12708 -11846 12717 -11812
rect 12665 -11880 12717 -11846
rect 12665 -11914 12674 -11880
rect 12708 -11914 12717 -11880
rect 12665 -11963 12717 -11914
rect 12752 -11819 12760 -11785
rect 12794 -11819 12803 -11785
rect 12923 -11785 12975 -11762
rect 12752 -11873 12803 -11819
rect 12752 -11907 12760 -11873
rect 12794 -11907 12803 -11873
rect 12752 -11923 12803 -11907
rect 12837 -11812 12889 -11796
rect 12837 -11846 12846 -11812
rect 12880 -11846 12889 -11812
rect 12837 -11880 12889 -11846
rect 12837 -11914 12846 -11880
rect 12880 -11914 12889 -11880
rect 12837 -11963 12889 -11914
rect 12923 -11819 12932 -11785
rect 12966 -11819 12975 -11785
rect 13120 -11765 13178 -11730
rect 13396 -11745 13546 -11675
rect 13672 -11658 13685 -11624
rect 13719 -11651 13735 -11624
rect 13672 -11685 13692 -11658
rect 13726 -11685 13735 -11651
rect 13672 -11701 13735 -11685
rect 13769 -11651 13819 -11542
rect 13853 -11508 13905 -11453
rect 13853 -11542 13862 -11508
rect 13896 -11542 13905 -11508
rect 13853 -11558 13905 -11542
rect 13941 -11508 13991 -11489
rect 13941 -11542 13948 -11508
rect 13982 -11542 13991 -11508
rect 13941 -11651 13991 -11542
rect 14025 -11508 14077 -11453
rect 14025 -11542 14034 -11508
rect 14068 -11542 14077 -11508
rect 14025 -11565 14077 -11542
rect 14111 -11508 14163 -11492
rect 14111 -11542 14120 -11508
rect 14154 -11542 14163 -11508
rect 14111 -11583 14163 -11542
rect 14197 -11499 14249 -11453
rect 14197 -11533 14206 -11499
rect 14240 -11533 14249 -11499
rect 14197 -11549 14249 -11533
rect 14283 -11508 14335 -11492
rect 14283 -11542 14292 -11508
rect 14326 -11542 14335 -11508
rect 14283 -11583 14335 -11542
rect 14369 -11499 14421 -11453
rect 14369 -11533 14378 -11499
rect 14412 -11533 14421 -11499
rect 14369 -11549 14421 -11533
rect 14455 -11508 14507 -11492
rect 14455 -11542 14464 -11508
rect 14498 -11542 14507 -11508
rect 14455 -11583 14507 -11542
rect 14541 -11499 14590 -11453
rect 14541 -11533 14550 -11499
rect 14584 -11533 14590 -11499
rect 14541 -11549 14590 -11533
rect 14624 -11508 14679 -11492
rect 14624 -11542 14636 -11508
rect 14670 -11542 14679 -11508
rect 14624 -11583 14679 -11542
rect 14713 -11499 14762 -11453
rect 14713 -11533 14722 -11499
rect 14756 -11533 14762 -11499
rect 14713 -11549 14762 -11533
rect 14796 -11508 14848 -11492
rect 14796 -11542 14807 -11508
rect 14841 -11542 14848 -11508
rect 14796 -11583 14848 -11542
rect 14884 -11499 14934 -11453
rect 14884 -11533 14893 -11499
rect 14927 -11533 14934 -11499
rect 14884 -11549 14934 -11533
rect 14968 -11508 15020 -11492
rect 14968 -11542 14979 -11508
rect 15013 -11542 15020 -11508
rect 14968 -11583 15020 -11542
rect 15056 -11499 15106 -11453
rect 15056 -11533 15065 -11499
rect 15099 -11533 15106 -11499
rect 15056 -11549 15106 -11533
rect 15140 -11508 15192 -11492
rect 15140 -11542 15151 -11508
rect 15185 -11542 15192 -11508
rect 15140 -11583 15192 -11542
rect 15228 -11499 15280 -11453
rect 15228 -11533 15237 -11499
rect 15271 -11533 15280 -11499
rect 15228 -11549 15280 -11533
rect 15314 -11508 15366 -11492
rect 15314 -11542 15323 -11508
rect 15357 -11542 15366 -11508
rect 15314 -11583 15366 -11542
rect 15400 -11499 15460 -11453
rect 15400 -11533 15409 -11499
rect 15443 -11533 15460 -11499
rect 15400 -11549 15460 -11533
rect 15512 -11547 15570 -11453
rect 15512 -11581 15524 -11547
rect 15558 -11581 15570 -11547
rect 14111 -11612 15460 -11583
rect 15512 -11598 15570 -11581
rect 15604 -11514 16673 -11453
rect 15604 -11548 15622 -11514
rect 15656 -11548 16622 -11514
rect 16656 -11548 16673 -11514
rect 14111 -11617 15248 -11612
rect 15227 -11646 15248 -11617
rect 15282 -11646 15341 -11612
rect 15375 -11646 15460 -11612
rect 13769 -11685 14119 -11651
rect 14153 -11685 14187 -11651
rect 14221 -11685 14255 -11651
rect 14289 -11685 14323 -11651
rect 14357 -11685 14391 -11651
rect 14425 -11685 14459 -11651
rect 14493 -11685 14527 -11651
rect 14561 -11685 14595 -11651
rect 14629 -11685 14663 -11651
rect 14697 -11685 14731 -11651
rect 14765 -11685 14799 -11651
rect 14833 -11685 14867 -11651
rect 14901 -11685 14935 -11651
rect 14969 -11685 15003 -11651
rect 15037 -11685 15071 -11651
rect 15105 -11685 15139 -11651
rect 15173 -11685 15193 -11651
rect 13769 -11701 15193 -11685
rect 12923 -11873 12975 -11819
rect 12923 -11907 12932 -11873
rect 12966 -11907 12975 -11873
rect 12923 -11923 12975 -11907
rect 13009 -11812 13086 -11796
rect 13009 -11846 13018 -11812
rect 13052 -11846 13086 -11812
rect 13009 -11880 13086 -11846
rect 13009 -11914 13018 -11880
rect 13052 -11914 13086 -11880
rect 13009 -11963 13086 -11914
rect 13120 -11799 13132 -11765
rect 13166 -11799 13178 -11765
rect 13120 -11858 13178 -11799
rect 13120 -11892 13132 -11858
rect 13166 -11892 13178 -11858
rect 13120 -11963 13178 -11892
rect 13212 -11785 13546 -11745
rect 13212 -11819 13230 -11785
rect 13264 -11819 13494 -11785
rect 13528 -11819 13546 -11785
rect 13212 -11887 13546 -11819
rect 13212 -11921 13230 -11887
rect 13264 -11921 13494 -11887
rect 13528 -11921 13546 -11887
rect 13212 -11963 13546 -11921
rect 13580 -11765 13638 -11730
rect 13580 -11799 13592 -11765
rect 13626 -11799 13638 -11765
rect 13580 -11858 13638 -11799
rect 13580 -11892 13592 -11858
rect 13626 -11892 13638 -11858
rect 13580 -11963 13638 -11892
rect 13674 -11819 13733 -11801
rect 13674 -11853 13690 -11819
rect 13724 -11853 13733 -11819
rect 13674 -11887 13733 -11853
rect 13674 -11921 13690 -11887
rect 13724 -11921 13733 -11887
rect 13674 -11963 13733 -11921
rect 13769 -11811 13818 -11701
rect 13769 -11845 13776 -11811
rect 13810 -11845 13818 -11811
rect 13769 -11879 13818 -11845
rect 13769 -11913 13776 -11879
rect 13810 -11913 13818 -11879
rect 13769 -11929 13818 -11913
rect 13853 -11819 13905 -11801
rect 13853 -11853 13862 -11819
rect 13896 -11853 13905 -11819
rect 13853 -11887 13905 -11853
rect 13853 -11921 13862 -11887
rect 13896 -11921 13905 -11887
rect 13853 -11963 13905 -11921
rect 13941 -11803 13991 -11701
rect 15227 -11708 15460 -11646
rect 15227 -11735 15248 -11708
rect 14111 -11742 15248 -11735
rect 15282 -11742 15340 -11708
rect 15374 -11742 15460 -11708
rect 15604 -11607 16673 -11548
rect 15604 -11677 16120 -11607
rect 15604 -11711 15682 -11677
rect 15716 -11711 15810 -11677
rect 15844 -11711 15938 -11677
rect 15972 -11711 16066 -11677
rect 16100 -11711 16120 -11677
rect 16154 -11675 16174 -11641
rect 16208 -11675 16302 -11641
rect 16336 -11675 16430 -11641
rect 16464 -11675 16558 -11641
rect 16592 -11675 16673 -11641
rect 14111 -11757 15460 -11742
rect 14111 -11791 14120 -11757
rect 14154 -11783 14292 -11757
rect 14154 -11791 14163 -11783
rect 13941 -11837 13948 -11803
rect 13982 -11837 13991 -11803
rect 13941 -11871 13991 -11837
rect 13941 -11905 13948 -11871
rect 13982 -11905 13991 -11871
rect 13941 -11928 13991 -11905
rect 14025 -11819 14077 -11803
rect 14025 -11853 14034 -11819
rect 14068 -11853 14077 -11819
rect 14025 -11887 14077 -11853
rect 14025 -11921 14034 -11887
rect 14068 -11921 14077 -11887
rect 14025 -11962 14077 -11921
rect 14111 -11843 14163 -11791
rect 14283 -11791 14292 -11783
rect 14326 -11783 14464 -11757
rect 14326 -11791 14335 -11783
rect 14111 -11877 14120 -11843
rect 14154 -11877 14163 -11843
rect 14111 -11928 14163 -11877
rect 14197 -11863 14249 -11817
rect 14197 -11897 14206 -11863
rect 14240 -11897 14249 -11863
rect 14197 -11962 14249 -11897
rect 14283 -11843 14335 -11791
rect 14455 -11791 14464 -11783
rect 14498 -11783 14636 -11757
rect 14498 -11791 14507 -11783
rect 14283 -11877 14292 -11843
rect 14326 -11877 14335 -11843
rect 14283 -11928 14335 -11877
rect 14369 -11863 14421 -11817
rect 14369 -11897 14378 -11863
rect 14412 -11897 14421 -11863
rect 14369 -11962 14421 -11897
rect 14455 -11843 14507 -11791
rect 14627 -11791 14636 -11783
rect 14670 -11783 14807 -11757
rect 14670 -11791 14679 -11783
rect 14455 -11877 14464 -11843
rect 14498 -11877 14507 -11843
rect 14455 -11928 14507 -11877
rect 14541 -11863 14593 -11817
rect 14541 -11897 14550 -11863
rect 14584 -11897 14593 -11863
rect 14541 -11962 14593 -11897
rect 14627 -11843 14679 -11791
rect 14796 -11791 14807 -11783
rect 14841 -11783 14979 -11757
rect 14841 -11791 14848 -11783
rect 14627 -11877 14636 -11843
rect 14670 -11877 14679 -11843
rect 14627 -11928 14679 -11877
rect 14713 -11863 14762 -11817
rect 14713 -11897 14722 -11863
rect 14756 -11897 14762 -11863
rect 14713 -11962 14762 -11897
rect 14796 -11843 14848 -11791
rect 14968 -11791 14979 -11783
rect 15013 -11783 15151 -11757
rect 15013 -11791 15020 -11783
rect 14796 -11877 14807 -11843
rect 14841 -11877 14848 -11843
rect 14796 -11928 14848 -11877
rect 14885 -11863 14934 -11817
rect 14885 -11897 14893 -11863
rect 14927 -11897 14934 -11863
rect 14885 -11962 14934 -11897
rect 14968 -11843 15020 -11791
rect 15140 -11791 15151 -11783
rect 15185 -11780 15323 -11757
rect 15185 -11791 15192 -11780
rect 14968 -11877 14979 -11843
rect 15013 -11877 15020 -11843
rect 14968 -11928 15020 -11877
rect 15057 -11863 15106 -11817
rect 15057 -11897 15065 -11863
rect 15099 -11897 15106 -11863
rect 15057 -11962 15106 -11897
rect 15140 -11843 15192 -11791
rect 15314 -11791 15323 -11780
rect 15357 -11780 15460 -11757
rect 15512 -11765 15570 -11730
rect 16154 -11745 16673 -11675
rect 15357 -11791 15372 -11780
rect 15140 -11877 15151 -11843
rect 15185 -11877 15192 -11843
rect 15140 -11928 15192 -11877
rect 15229 -11863 15280 -11817
rect 15229 -11897 15237 -11863
rect 15271 -11897 15280 -11863
rect 15229 -11962 15280 -11897
rect 15314 -11843 15372 -11791
rect 15512 -11799 15524 -11765
rect 15558 -11799 15570 -11765
rect 15314 -11877 15323 -11843
rect 15357 -11877 15372 -11843
rect 15314 -11928 15372 -11877
rect 15406 -11863 15460 -11814
rect 15406 -11897 15409 -11863
rect 15443 -11897 15460 -11863
rect 14025 -11963 15280 -11962
rect 15406 -11963 15460 -11897
rect 15512 -11858 15570 -11799
rect 15512 -11892 15524 -11858
rect 15558 -11892 15570 -11858
rect 15512 -11963 15570 -11892
rect 15604 -11785 16673 -11745
rect 15604 -11819 15622 -11785
rect 15656 -11819 16622 -11785
rect 16656 -11819 16673 -11785
rect 15604 -11887 16673 -11819
rect 15604 -11921 15622 -11887
rect 15656 -11921 16622 -11887
rect 16656 -11921 16673 -11887
rect 15604 -11963 16673 -11921
rect -2997 -11997 -2968 -11963
rect -2934 -11997 -2876 -11963
rect -2842 -11997 -2784 -11963
rect -2750 -11997 -2692 -11963
rect -2658 -11997 -2600 -11963
rect -2566 -11997 -2508 -11963
rect -2474 -11997 -2416 -11963
rect -2382 -11997 -2324 -11963
rect -2290 -11997 -2232 -11963
rect -2198 -11997 -2140 -11963
rect -2106 -11997 -2048 -11963
rect -2014 -11997 -1956 -11963
rect -1922 -11997 -1864 -11963
rect -1830 -11997 -1772 -11963
rect -1738 -11997 -1680 -11963
rect -1646 -11997 -1588 -11963
rect -1554 -11997 -1496 -11963
rect -1462 -11997 -1404 -11963
rect -1370 -11997 -1312 -11963
rect -1278 -11997 -1220 -11963
rect -1186 -11997 -1128 -11963
rect -1094 -11997 -1036 -11963
rect -1002 -11997 -944 -11963
rect -910 -11997 -852 -11963
rect -818 -11997 -760 -11963
rect -726 -11997 -668 -11963
rect -634 -11997 -576 -11963
rect -542 -11997 -484 -11963
rect -450 -11997 -392 -11963
rect -358 -11997 -300 -11963
rect -266 -11997 -208 -11963
rect -174 -11997 -116 -11963
rect -82 -11997 -24 -11963
rect 10 -11997 68 -11963
rect 102 -11997 160 -11963
rect 194 -11997 252 -11963
rect 286 -11997 344 -11963
rect 378 -11997 436 -11963
rect 470 -11997 528 -11963
rect 562 -11997 620 -11963
rect 654 -11997 712 -11963
rect 746 -11997 804 -11963
rect 838 -11997 896 -11963
rect 930 -11997 988 -11963
rect 1022 -11997 1080 -11963
rect 1114 -11997 1172 -11963
rect 1206 -11997 1264 -11963
rect 1298 -11997 1356 -11963
rect 1390 -11997 1448 -11963
rect 1482 -11997 1540 -11963
rect 1574 -11997 1632 -11963
rect 1666 -11997 1724 -11963
rect 1758 -11997 1816 -11963
rect 1850 -11997 1908 -11963
rect 1942 -11997 2000 -11963
rect 2034 -11997 2092 -11963
rect 2126 -11997 2184 -11963
rect 2218 -11997 2276 -11963
rect 2310 -11997 2368 -11963
rect 2402 -11997 2460 -11963
rect 2494 -11997 2552 -11963
rect 2586 -11997 2644 -11963
rect 2678 -11997 2736 -11963
rect 2770 -11997 2828 -11963
rect 2862 -11997 2920 -11963
rect 2954 -11997 3012 -11963
rect 3046 -11997 3104 -11963
rect 3138 -11997 3196 -11963
rect 3230 -11997 3288 -11963
rect 3322 -11997 3380 -11963
rect 3414 -11997 3472 -11963
rect 3506 -11997 3564 -11963
rect 3598 -11997 3656 -11963
rect 3690 -11997 3748 -11963
rect 3782 -11997 3840 -11963
rect 3874 -11997 3932 -11963
rect 3966 -11997 4024 -11963
rect 4058 -11997 4116 -11963
rect 4150 -11997 4208 -11963
rect 4242 -11997 4300 -11963
rect 4334 -11997 4392 -11963
rect 4426 -11997 4484 -11963
rect 4518 -11997 4576 -11963
rect 4610 -11997 4668 -11963
rect 4702 -11997 4760 -11963
rect 4794 -11997 4852 -11963
rect 4886 -11997 4944 -11963
rect 4978 -11997 5036 -11963
rect 5070 -11997 5128 -11963
rect 5162 -11997 5220 -11963
rect 5254 -11997 5312 -11963
rect 5346 -11997 5404 -11963
rect 5438 -11997 5496 -11963
rect 5530 -11997 5588 -11963
rect 5622 -11997 5680 -11963
rect 5714 -11997 5772 -11963
rect 5806 -11997 5864 -11963
rect 5898 -11997 5956 -11963
rect 5990 -11997 6048 -11963
rect 6082 -11997 6140 -11963
rect 6174 -11997 6232 -11963
rect 6266 -11997 6324 -11963
rect 6358 -11997 6416 -11963
rect 6450 -11997 6508 -11963
rect 6542 -11997 6600 -11963
rect 6634 -11997 6692 -11963
rect 6726 -11997 6784 -11963
rect 6818 -11997 6876 -11963
rect 6910 -11997 6968 -11963
rect 7002 -11997 7060 -11963
rect 7094 -11997 7152 -11963
rect 7186 -11997 7244 -11963
rect 7278 -11997 7336 -11963
rect 7370 -11997 7428 -11963
rect 7462 -11997 7520 -11963
rect 7554 -11997 7612 -11963
rect 7646 -11997 7704 -11963
rect 7738 -11997 7796 -11963
rect 7830 -11997 7888 -11963
rect 7922 -11997 7980 -11963
rect 8014 -11997 8072 -11963
rect 8106 -11997 8164 -11963
rect 8198 -11997 8256 -11963
rect 8290 -11997 8348 -11963
rect 8382 -11997 8440 -11963
rect 8474 -11997 8532 -11963
rect 8566 -11997 8624 -11963
rect 8658 -11997 8716 -11963
rect 8750 -11997 8808 -11963
rect 8842 -11997 8900 -11963
rect 8934 -11997 8992 -11963
rect 9026 -11997 9084 -11963
rect 9118 -11997 9176 -11963
rect 9210 -11997 9268 -11963
rect 9302 -11997 9360 -11963
rect 9394 -11997 9452 -11963
rect 9486 -11997 9544 -11963
rect 9578 -11997 9636 -11963
rect 9670 -11997 9728 -11963
rect 9762 -11997 9820 -11963
rect 9854 -11997 9912 -11963
rect 9946 -11997 10004 -11963
rect 10038 -11997 10096 -11963
rect 10130 -11997 10188 -11963
rect 10222 -11997 10280 -11963
rect 10314 -11997 10372 -11963
rect 10406 -11997 10464 -11963
rect 10498 -11997 10556 -11963
rect 10590 -11997 10648 -11963
rect 10682 -11997 10740 -11963
rect 10774 -11997 10832 -11963
rect 10866 -11997 10924 -11963
rect 10958 -11997 11016 -11963
rect 11050 -11997 11108 -11963
rect 11142 -11997 11200 -11963
rect 11234 -11997 11292 -11963
rect 11326 -11997 11384 -11963
rect 11418 -11997 11476 -11963
rect 11510 -11997 11568 -11963
rect 11602 -11997 11660 -11963
rect 11694 -11997 11752 -11963
rect 11786 -11997 11844 -11963
rect 11878 -11997 11936 -11963
rect 11970 -11997 12028 -11963
rect 12062 -11997 12120 -11963
rect 12154 -11997 12212 -11963
rect 12246 -11997 12304 -11963
rect 12338 -11997 12396 -11963
rect 12430 -11997 12488 -11963
rect 12522 -11997 12580 -11963
rect 12614 -11997 12672 -11963
rect 12706 -11997 12764 -11963
rect 12798 -11997 12856 -11963
rect 12890 -11997 12948 -11963
rect 12982 -11997 13040 -11963
rect 13074 -11997 13132 -11963
rect 13166 -11997 13224 -11963
rect 13258 -11997 13316 -11963
rect 13350 -11997 13408 -11963
rect 13442 -11997 13500 -11963
rect 13534 -11997 13592 -11963
rect 13626 -11997 13684 -11963
rect 13718 -11997 13776 -11963
rect 13810 -11997 13868 -11963
rect 13902 -11997 13960 -11963
rect 13994 -11997 14052 -11963
rect 14086 -11997 14144 -11963
rect 14178 -11997 14236 -11963
rect 14270 -11997 14328 -11963
rect 14362 -11997 14420 -11963
rect 14454 -11997 14512 -11963
rect 14546 -11997 14604 -11963
rect 14638 -11997 14696 -11963
rect 14730 -11997 14788 -11963
rect 14822 -11997 14880 -11963
rect 14914 -11997 14972 -11963
rect 15006 -11997 15064 -11963
rect 15098 -11997 15156 -11963
rect 15190 -11997 15248 -11963
rect 15282 -11997 15340 -11963
rect 15374 -11997 15432 -11963
rect 15466 -11997 15524 -11963
rect 15558 -11997 15616 -11963
rect 15650 -11997 15708 -11963
rect 15742 -11997 15800 -11963
rect 15834 -11997 15892 -11963
rect 15926 -11997 15984 -11963
rect 16018 -11997 16076 -11963
rect 16110 -11997 16168 -11963
rect 16202 -11997 16260 -11963
rect 16294 -11997 16352 -11963
rect 16386 -11997 16444 -11963
rect 16478 -11997 16536 -11963
rect 16570 -11997 16628 -11963
rect 16662 -11997 16691 -11963
rect -2980 -12039 -2278 -11997
rect -2980 -12073 -2962 -12039
rect -2928 -12073 -2330 -12039
rect -2296 -12073 -2278 -12039
rect -2980 -12141 -2278 -12073
rect -2980 -12175 -2962 -12141
rect -2928 -12175 -2330 -12141
rect -2296 -12175 -2278 -12141
rect -2980 -12215 -2278 -12175
rect -2980 -12283 -2902 -12249
rect -2868 -12283 -2803 -12249
rect -2769 -12283 -2704 -12249
rect -2670 -12283 -2650 -12249
rect -2980 -12353 -2650 -12283
rect -2616 -12285 -2278 -12215
rect -2244 -12068 -2186 -11997
rect -2244 -12102 -2232 -12068
rect -2198 -12102 -2186 -12068
rect -2244 -12161 -2186 -12102
rect -2244 -12195 -2232 -12161
rect -2198 -12195 -2186 -12161
rect -2244 -12230 -2186 -12195
rect -1600 -12039 -898 -11997
rect -1600 -12073 -1582 -12039
rect -1548 -12073 -950 -12039
rect -916 -12073 -898 -12039
rect -1600 -12141 -898 -12073
rect -1600 -12175 -1582 -12141
rect -1548 -12175 -950 -12141
rect -916 -12175 -898 -12141
rect -1600 -12215 -898 -12175
rect -864 -12047 -783 -12031
rect -864 -12081 -831 -12047
rect -797 -12081 -783 -12047
rect -864 -12115 -783 -12081
rect -864 -12149 -831 -12115
rect -797 -12149 -783 -12115
rect -864 -12186 -783 -12149
rect -749 -12046 -683 -11997
rect -749 -12080 -733 -12046
rect -699 -12080 -683 -12046
rect -749 -12114 -683 -12080
rect -749 -12148 -733 -12114
rect -699 -12148 -683 -12114
rect -749 -12157 -683 -12148
rect -593 -12047 -543 -12031
rect -593 -12081 -577 -12047
rect -593 -12115 -543 -12081
rect -593 -12149 -577 -12115
rect -2616 -12319 -2596 -12285
rect -2562 -12319 -2493 -12285
rect -2459 -12319 -2390 -12285
rect -2356 -12319 -2278 -12285
rect -1600 -12285 -1262 -12215
rect -864 -12235 -814 -12186
rect -593 -12191 -543 -12149
rect -1600 -12319 -1522 -12285
rect -1488 -12319 -1419 -12285
rect -1385 -12319 -1316 -12285
rect -1282 -12319 -1262 -12285
rect -1228 -12283 -1208 -12249
rect -1174 -12283 -1109 -12249
rect -1075 -12283 -1010 -12249
rect -976 -12283 -898 -12249
rect -1228 -12353 -898 -12283
rect -2980 -12412 -2278 -12353
rect -2980 -12446 -2962 -12412
rect -2928 -12446 -2330 -12412
rect -2296 -12446 -2278 -12412
rect -2980 -12507 -2278 -12446
rect -2244 -12379 -2186 -12362
rect -2244 -12413 -2232 -12379
rect -2198 -12413 -2186 -12379
rect -2244 -12507 -2186 -12413
rect -1600 -12412 -898 -12353
rect -1600 -12446 -1582 -12412
rect -1548 -12446 -950 -12412
rect -916 -12446 -898 -12412
rect -1600 -12507 -898 -12446
rect -864 -12269 -855 -12235
rect -821 -12269 -814 -12235
rect -661 -12225 -543 -12191
rect -491 -12046 -421 -12031
rect -491 -12080 -473 -12046
rect -439 -12080 -421 -12046
rect -491 -12114 -421 -12080
rect -491 -12148 -473 -12114
rect -439 -12148 -421 -12114
rect -661 -12259 -627 -12225
rect -864 -12396 -814 -12269
rect -780 -12275 -627 -12259
rect -491 -12260 -421 -12148
rect -331 -12046 -265 -11997
rect -331 -12080 -315 -12046
rect -281 -12080 -265 -12046
rect -331 -12114 -265 -12080
rect -331 -12148 -315 -12114
rect -281 -12148 -265 -12114
rect -331 -12164 -265 -12148
rect -231 -12046 -162 -12031
rect -231 -12080 -215 -12046
rect -181 -12080 -162 -12046
rect -231 -12114 -162 -12080
rect -231 -12148 -215 -12114
rect -181 -12148 -162 -12114
rect -231 -12198 -162 -12148
rect -780 -12309 -777 -12275
rect -743 -12309 -627 -12275
rect -780 -12325 -627 -12309
rect -593 -12275 -421 -12260
rect -356 -12232 -162 -12198
rect -128 -12068 -70 -11997
rect -128 -12102 -116 -12068
rect -82 -12102 -70 -12068
rect -128 -12161 -70 -12102
rect -128 -12195 -116 -12161
rect -82 -12195 -70 -12161
rect -128 -12230 -70 -12195
rect -36 -12039 298 -11997
rect -36 -12073 -18 -12039
rect 16 -12073 246 -12039
rect 280 -12073 298 -12039
rect -36 -12141 298 -12073
rect -36 -12175 -18 -12141
rect 16 -12175 246 -12141
rect 280 -12175 298 -12141
rect -36 -12215 298 -12175
rect 332 -12068 390 -11997
rect 332 -12102 344 -12068
rect 378 -12102 390 -12068
rect 332 -12161 390 -12102
rect 332 -12195 344 -12161
rect 378 -12195 390 -12161
rect -356 -12261 -286 -12232
rect -593 -12309 -577 -12275
rect -543 -12309 -421 -12275
rect -593 -12310 -421 -12309
rect -661 -12344 -627 -12325
rect -661 -12378 -543 -12344
rect -864 -12420 -783 -12396
rect -864 -12454 -831 -12420
rect -797 -12454 -783 -12420
rect -864 -12473 -783 -12454
rect -749 -12420 -683 -12404
rect -749 -12454 -733 -12420
rect -699 -12454 -683 -12420
rect -749 -12507 -683 -12454
rect -593 -12420 -543 -12378
rect -593 -12454 -577 -12420
rect -593 -12473 -543 -12454
rect -491 -12420 -421 -12310
rect -372 -12275 -286 -12261
rect -372 -12309 -356 -12275
rect -322 -12309 -286 -12275
rect -252 -12272 -162 -12266
rect -252 -12275 -210 -12272
rect -252 -12309 -236 -12275
rect -176 -12306 -162 -12272
rect -202 -12309 -162 -12306
rect -36 -12285 114 -12215
rect 332 -12230 390 -12195
rect 424 -12047 505 -12031
rect 424 -12081 457 -12047
rect 491 -12081 505 -12047
rect 424 -12115 505 -12081
rect 424 -12149 457 -12115
rect 491 -12149 505 -12115
rect 424 -12186 505 -12149
rect 539 -12046 605 -11997
rect 539 -12080 555 -12046
rect 589 -12080 605 -12046
rect 539 -12114 605 -12080
rect 539 -12148 555 -12114
rect 589 -12148 605 -12114
rect 539 -12157 605 -12148
rect 695 -12047 745 -12031
rect 695 -12081 711 -12047
rect 695 -12115 745 -12081
rect 695 -12149 711 -12115
rect 424 -12235 474 -12186
rect 695 -12191 745 -12149
rect -372 -12319 -286 -12309
rect -36 -12319 -16 -12285
rect 18 -12319 114 -12285
rect 148 -12283 244 -12249
rect 278 -12283 298 -12249
rect -356 -12343 -286 -12319
rect -356 -12377 -162 -12343
rect 148 -12353 298 -12283
rect -491 -12454 -472 -12420
rect -438 -12454 -421 -12420
rect -491 -12473 -421 -12454
rect -328 -12420 -262 -12411
rect -328 -12454 -312 -12420
rect -278 -12454 -262 -12420
rect -328 -12507 -262 -12454
rect -228 -12420 -162 -12377
rect -228 -12454 -215 -12420
rect -181 -12454 -162 -12420
rect -228 -12473 -162 -12454
rect -128 -12379 -70 -12362
rect -128 -12413 -116 -12379
rect -82 -12413 -70 -12379
rect -128 -12507 -70 -12413
rect -36 -12405 298 -12353
rect 424 -12269 433 -12235
rect 467 -12269 474 -12235
rect 627 -12225 745 -12191
rect 797 -12046 867 -12031
rect 797 -12080 815 -12046
rect 849 -12080 867 -12046
rect 797 -12114 867 -12080
rect 797 -12148 815 -12114
rect 849 -12148 867 -12114
rect 627 -12259 661 -12225
rect -36 -12439 -18 -12405
rect 16 -12439 246 -12405
rect 280 -12439 298 -12405
rect -36 -12507 298 -12439
rect 332 -12379 390 -12362
rect 332 -12413 344 -12379
rect 378 -12413 390 -12379
rect 332 -12507 390 -12413
rect 424 -12396 474 -12269
rect 508 -12275 661 -12259
rect 797 -12260 867 -12148
rect 957 -12046 1023 -11997
rect 957 -12080 973 -12046
rect 1007 -12080 1023 -12046
rect 957 -12114 1023 -12080
rect 957 -12148 973 -12114
rect 1007 -12148 1023 -12114
rect 957 -12164 1023 -12148
rect 1057 -12046 1126 -12031
rect 1057 -12080 1073 -12046
rect 1107 -12080 1126 -12046
rect 1057 -12114 1126 -12080
rect 1057 -12148 1073 -12114
rect 1107 -12148 1126 -12114
rect 1057 -12198 1126 -12148
rect 508 -12309 511 -12275
rect 545 -12309 661 -12275
rect 508 -12325 661 -12309
rect 695 -12275 867 -12260
rect 932 -12232 1126 -12198
rect 1160 -12068 1218 -11997
rect 1160 -12102 1172 -12068
rect 1206 -12102 1218 -12068
rect 1160 -12161 1218 -12102
rect 1160 -12195 1172 -12161
rect 1206 -12195 1218 -12161
rect 1160 -12230 1218 -12195
rect 1252 -12039 1586 -11997
rect 1252 -12073 1270 -12039
rect 1304 -12073 1534 -12039
rect 1568 -12073 1586 -12039
rect 1252 -12141 1586 -12073
rect 1252 -12175 1270 -12141
rect 1304 -12175 1534 -12141
rect 1568 -12175 1586 -12141
rect 1252 -12215 1586 -12175
rect 1620 -12068 1678 -11997
rect 1620 -12102 1632 -12068
rect 1666 -12102 1678 -12068
rect 1620 -12161 1678 -12102
rect 1620 -12195 1632 -12161
rect 1666 -12195 1678 -12161
rect 932 -12261 1002 -12232
rect 695 -12309 711 -12275
rect 745 -12309 867 -12275
rect 695 -12310 867 -12309
rect 627 -12344 661 -12325
rect 627 -12378 745 -12344
rect 424 -12420 505 -12396
rect 424 -12454 457 -12420
rect 491 -12454 505 -12420
rect 424 -12473 505 -12454
rect 539 -12420 605 -12404
rect 539 -12454 555 -12420
rect 589 -12454 605 -12420
rect 539 -12507 605 -12454
rect 695 -12420 745 -12378
rect 695 -12454 711 -12420
rect 695 -12473 745 -12454
rect 797 -12420 867 -12310
rect 916 -12275 1002 -12261
rect 916 -12309 932 -12275
rect 966 -12309 1002 -12275
rect 1036 -12268 1126 -12266
rect 1036 -12275 1054 -12268
rect 1036 -12309 1052 -12275
rect 1088 -12302 1126 -12268
rect 1086 -12309 1126 -12302
rect 1252 -12285 1402 -12215
rect 1620 -12230 1678 -12195
rect 1712 -12039 2414 -11997
rect 1712 -12073 1730 -12039
rect 1764 -12073 2362 -12039
rect 2396 -12073 2414 -12039
rect 1712 -12141 2414 -12073
rect 1712 -12175 1730 -12141
rect 1764 -12175 2362 -12141
rect 2396 -12175 2414 -12141
rect 1712 -12215 2414 -12175
rect 916 -12319 1002 -12309
rect 1252 -12319 1272 -12285
rect 1306 -12319 1402 -12285
rect 1436 -12283 1532 -12249
rect 1566 -12283 1586 -12249
rect 932 -12343 1002 -12319
rect 932 -12377 1126 -12343
rect 1436 -12353 1586 -12283
rect 797 -12454 816 -12420
rect 850 -12454 867 -12420
rect 797 -12473 867 -12454
rect 960 -12420 1026 -12411
rect 960 -12454 976 -12420
rect 1010 -12454 1026 -12420
rect 960 -12507 1026 -12454
rect 1060 -12420 1126 -12377
rect 1060 -12454 1073 -12420
rect 1107 -12454 1126 -12420
rect 1060 -12473 1126 -12454
rect 1160 -12379 1218 -12362
rect 1160 -12413 1172 -12379
rect 1206 -12413 1218 -12379
rect 1160 -12507 1218 -12413
rect 1252 -12405 1586 -12353
rect 1712 -12283 1790 -12249
rect 1824 -12283 1889 -12249
rect 1923 -12283 1988 -12249
rect 2022 -12283 2042 -12249
rect 1712 -12353 2042 -12283
rect 2076 -12285 2414 -12215
rect 2448 -12068 2506 -11997
rect 2448 -12102 2460 -12068
rect 2494 -12102 2506 -12068
rect 2448 -12161 2506 -12102
rect 2448 -12195 2460 -12161
rect 2494 -12195 2506 -12161
rect 2448 -12230 2506 -12195
rect 2540 -12039 2874 -11997
rect 2540 -12073 2558 -12039
rect 2592 -12073 2822 -12039
rect 2856 -12073 2874 -12039
rect 2540 -12141 2874 -12073
rect 2540 -12175 2558 -12141
rect 2592 -12175 2822 -12141
rect 2856 -12175 2874 -12141
rect 2540 -12215 2874 -12175
rect 2908 -12068 2966 -11997
rect 2908 -12102 2920 -12068
rect 2954 -12102 2966 -12068
rect 2908 -12161 2966 -12102
rect 2908 -12195 2920 -12161
rect 2954 -12195 2966 -12161
rect 2076 -12319 2096 -12285
rect 2130 -12319 2199 -12285
rect 2233 -12319 2302 -12285
rect 2336 -12319 2414 -12285
rect 2540 -12285 2690 -12215
rect 2908 -12230 2966 -12195
rect 3000 -12047 3081 -12031
rect 3000 -12081 3033 -12047
rect 3067 -12081 3081 -12047
rect 3000 -12115 3081 -12081
rect 3000 -12149 3033 -12115
rect 3067 -12149 3081 -12115
rect 3000 -12186 3081 -12149
rect 3115 -12046 3181 -11997
rect 3115 -12080 3131 -12046
rect 3165 -12080 3181 -12046
rect 3115 -12114 3181 -12080
rect 3115 -12148 3131 -12114
rect 3165 -12148 3181 -12114
rect 3115 -12157 3181 -12148
rect 3271 -12047 3321 -12031
rect 3271 -12081 3287 -12047
rect 3271 -12115 3321 -12081
rect 3271 -12149 3287 -12115
rect 2540 -12319 2560 -12285
rect 2594 -12319 2690 -12285
rect 2724 -12283 2820 -12249
rect 2854 -12283 2874 -12249
rect 2724 -12353 2874 -12283
rect 1252 -12439 1270 -12405
rect 1304 -12439 1534 -12405
rect 1568 -12439 1586 -12405
rect 1252 -12507 1586 -12439
rect 1620 -12379 1678 -12362
rect 1620 -12413 1632 -12379
rect 1666 -12413 1678 -12379
rect 1620 -12507 1678 -12413
rect 1712 -12412 2414 -12353
rect 1712 -12446 1730 -12412
rect 1764 -12446 2362 -12412
rect 2396 -12446 2414 -12412
rect 1712 -12507 2414 -12446
rect 2448 -12379 2506 -12362
rect 2448 -12413 2460 -12379
rect 2494 -12413 2506 -12379
rect 2448 -12507 2506 -12413
rect 2540 -12405 2874 -12353
rect 3000 -12268 3050 -12186
rect 3271 -12191 3321 -12149
rect 3203 -12225 3321 -12191
rect 3373 -12046 3443 -12031
rect 3373 -12080 3391 -12046
rect 3425 -12080 3443 -12046
rect 3373 -12114 3443 -12080
rect 3373 -12148 3391 -12114
rect 3425 -12148 3443 -12114
rect 3203 -12259 3237 -12225
rect 3000 -12302 3014 -12268
rect 3048 -12302 3050 -12268
rect 2540 -12439 2558 -12405
rect 2592 -12439 2822 -12405
rect 2856 -12439 2874 -12405
rect 2540 -12507 2874 -12439
rect 2908 -12379 2966 -12362
rect 2908 -12413 2920 -12379
rect 2954 -12413 2966 -12379
rect 2908 -12507 2966 -12413
rect 3000 -12396 3050 -12302
rect 3084 -12275 3237 -12259
rect 3373 -12260 3443 -12148
rect 3533 -12046 3599 -11997
rect 3533 -12080 3549 -12046
rect 3583 -12080 3599 -12046
rect 3533 -12114 3599 -12080
rect 3533 -12148 3549 -12114
rect 3583 -12148 3599 -12114
rect 3533 -12164 3599 -12148
rect 3633 -12046 3702 -12031
rect 3633 -12080 3649 -12046
rect 3683 -12080 3702 -12046
rect 3633 -12114 3702 -12080
rect 3633 -12148 3649 -12114
rect 3683 -12148 3702 -12114
rect 3633 -12198 3702 -12148
rect 3084 -12309 3087 -12275
rect 3121 -12309 3237 -12275
rect 3084 -12325 3237 -12309
rect 3271 -12275 3443 -12260
rect 3508 -12232 3702 -12198
rect 3736 -12068 3794 -11997
rect 3736 -12102 3748 -12068
rect 3782 -12102 3794 -12068
rect 3736 -12161 3794 -12102
rect 3736 -12195 3748 -12161
rect 3782 -12195 3794 -12161
rect 3736 -12230 3794 -12195
rect 3828 -12039 4162 -11997
rect 3828 -12073 3846 -12039
rect 3880 -12073 4110 -12039
rect 4144 -12073 4162 -12039
rect 3828 -12141 4162 -12073
rect 3828 -12175 3846 -12141
rect 3880 -12175 4110 -12141
rect 4144 -12175 4162 -12141
rect 3828 -12215 4162 -12175
rect 4196 -12068 4254 -11997
rect 4196 -12102 4208 -12068
rect 4242 -12102 4254 -12068
rect 4196 -12161 4254 -12102
rect 4196 -12195 4208 -12161
rect 4242 -12195 4254 -12161
rect 3508 -12261 3578 -12232
rect 3271 -12309 3287 -12275
rect 3321 -12309 3443 -12275
rect 3271 -12310 3443 -12309
rect 3203 -12344 3237 -12325
rect 3203 -12378 3321 -12344
rect 3000 -12420 3081 -12396
rect 3000 -12454 3033 -12420
rect 3067 -12454 3081 -12420
rect 3000 -12473 3081 -12454
rect 3115 -12420 3181 -12404
rect 3115 -12454 3131 -12420
rect 3165 -12454 3181 -12420
rect 3115 -12507 3181 -12454
rect 3271 -12420 3321 -12378
rect 3271 -12454 3287 -12420
rect 3271 -12473 3321 -12454
rect 3373 -12420 3443 -12310
rect 3492 -12275 3578 -12261
rect 3492 -12309 3508 -12275
rect 3542 -12309 3578 -12275
rect 3612 -12268 3702 -12266
rect 3612 -12309 3628 -12268
rect 3662 -12309 3702 -12268
rect 3828 -12285 3978 -12215
rect 4196 -12230 4254 -12195
rect 4288 -12039 4990 -11997
rect 4288 -12073 4306 -12039
rect 4340 -12073 4938 -12039
rect 4972 -12073 4990 -12039
rect 4288 -12141 4990 -12073
rect 4288 -12175 4306 -12141
rect 4340 -12175 4938 -12141
rect 4972 -12175 4990 -12141
rect 4288 -12215 4990 -12175
rect 3492 -12319 3578 -12309
rect 3828 -12319 3848 -12285
rect 3882 -12319 3978 -12285
rect 4012 -12283 4108 -12249
rect 4142 -12283 4162 -12249
rect 3508 -12343 3578 -12319
rect 3508 -12377 3702 -12343
rect 4012 -12353 4162 -12283
rect 3373 -12454 3392 -12420
rect 3426 -12454 3443 -12420
rect 3373 -12473 3443 -12454
rect 3536 -12420 3602 -12411
rect 3536 -12454 3552 -12420
rect 3586 -12454 3602 -12420
rect 3536 -12507 3602 -12454
rect 3636 -12420 3702 -12377
rect 3636 -12454 3649 -12420
rect 3683 -12454 3702 -12420
rect 3636 -12473 3702 -12454
rect 3736 -12379 3794 -12362
rect 3736 -12413 3748 -12379
rect 3782 -12413 3794 -12379
rect 3736 -12507 3794 -12413
rect 3828 -12405 4162 -12353
rect 4288 -12283 4366 -12249
rect 4400 -12283 4465 -12249
rect 4499 -12283 4564 -12249
rect 4598 -12283 4618 -12249
rect 4288 -12353 4618 -12283
rect 4652 -12285 4990 -12215
rect 5024 -12068 5082 -11997
rect 5024 -12102 5036 -12068
rect 5070 -12102 5082 -12068
rect 5024 -12161 5082 -12102
rect 5024 -12195 5036 -12161
rect 5070 -12195 5082 -12161
rect 5024 -12230 5082 -12195
rect 5116 -12039 5450 -11997
rect 5116 -12073 5134 -12039
rect 5168 -12073 5398 -12039
rect 5432 -12073 5450 -12039
rect 5116 -12141 5450 -12073
rect 5116 -12175 5134 -12141
rect 5168 -12175 5398 -12141
rect 5432 -12175 5450 -12141
rect 5116 -12215 5450 -12175
rect 5484 -12068 5542 -11997
rect 5484 -12102 5496 -12068
rect 5530 -12102 5542 -12068
rect 5484 -12161 5542 -12102
rect 5484 -12195 5496 -12161
rect 5530 -12195 5542 -12161
rect 4652 -12319 4672 -12285
rect 4706 -12319 4775 -12285
rect 4809 -12319 4878 -12285
rect 4912 -12319 4990 -12285
rect 5116 -12285 5266 -12215
rect 5484 -12230 5542 -12195
rect 5576 -12047 5657 -12031
rect 5576 -12081 5609 -12047
rect 5643 -12081 5657 -12047
rect 5576 -12115 5657 -12081
rect 5576 -12149 5609 -12115
rect 5643 -12149 5657 -12115
rect 5576 -12186 5657 -12149
rect 5691 -12046 5757 -11997
rect 5691 -12080 5707 -12046
rect 5741 -12080 5757 -12046
rect 5691 -12114 5757 -12080
rect 5691 -12148 5707 -12114
rect 5741 -12148 5757 -12114
rect 5691 -12157 5757 -12148
rect 5847 -12047 5897 -12031
rect 5847 -12081 5863 -12047
rect 5847 -12115 5897 -12081
rect 5847 -12149 5863 -12115
rect 5116 -12319 5136 -12285
rect 5170 -12319 5266 -12285
rect 5300 -12283 5396 -12249
rect 5430 -12283 5450 -12249
rect 5300 -12353 5450 -12283
rect 3828 -12439 3846 -12405
rect 3880 -12439 4110 -12405
rect 4144 -12439 4162 -12405
rect 3828 -12507 4162 -12439
rect 4196 -12379 4254 -12362
rect 4196 -12413 4208 -12379
rect 4242 -12413 4254 -12379
rect 4196 -12507 4254 -12413
rect 4288 -12412 4990 -12353
rect 4288 -12446 4306 -12412
rect 4340 -12446 4938 -12412
rect 4972 -12446 4990 -12412
rect 4288 -12507 4990 -12446
rect 5024 -12379 5082 -12362
rect 5024 -12413 5036 -12379
rect 5070 -12413 5082 -12379
rect 5024 -12507 5082 -12413
rect 5116 -12405 5450 -12353
rect 5576 -12268 5626 -12186
rect 5847 -12191 5897 -12149
rect 5779 -12225 5897 -12191
rect 5949 -12046 6019 -12031
rect 5949 -12080 5967 -12046
rect 6001 -12080 6019 -12046
rect 5949 -12114 6019 -12080
rect 5949 -12148 5967 -12114
rect 6001 -12148 6019 -12114
rect 5779 -12259 5813 -12225
rect 5576 -12302 5588 -12268
rect 5622 -12302 5626 -12268
rect 5116 -12439 5134 -12405
rect 5168 -12439 5398 -12405
rect 5432 -12439 5450 -12405
rect 5116 -12507 5450 -12439
rect 5484 -12379 5542 -12362
rect 5484 -12413 5496 -12379
rect 5530 -12413 5542 -12379
rect 5484 -12507 5542 -12413
rect 5576 -12396 5626 -12302
rect 5660 -12275 5813 -12259
rect 5949 -12260 6019 -12148
rect 6109 -12046 6175 -11997
rect 6109 -12080 6125 -12046
rect 6159 -12080 6175 -12046
rect 6109 -12114 6175 -12080
rect 6109 -12148 6125 -12114
rect 6159 -12148 6175 -12114
rect 6109 -12164 6175 -12148
rect 6209 -12046 6278 -12031
rect 6209 -12080 6225 -12046
rect 6259 -12080 6278 -12046
rect 6209 -12114 6278 -12080
rect 6209 -12148 6225 -12114
rect 6259 -12148 6278 -12114
rect 6209 -12198 6278 -12148
rect 5660 -12309 5663 -12275
rect 5697 -12309 5813 -12275
rect 5660 -12325 5813 -12309
rect 5847 -12275 6019 -12260
rect 6084 -12232 6278 -12198
rect 6312 -12068 6370 -11997
rect 6312 -12102 6324 -12068
rect 6358 -12102 6370 -12068
rect 6312 -12161 6370 -12102
rect 6312 -12195 6324 -12161
rect 6358 -12195 6370 -12161
rect 6312 -12230 6370 -12195
rect 6404 -12039 6738 -11997
rect 6404 -12073 6422 -12039
rect 6456 -12073 6686 -12039
rect 6720 -12073 6738 -12039
rect 6404 -12141 6738 -12073
rect 6404 -12175 6422 -12141
rect 6456 -12175 6686 -12141
rect 6720 -12175 6738 -12141
rect 6404 -12215 6738 -12175
rect 6772 -12068 6830 -11997
rect 6772 -12102 6784 -12068
rect 6818 -12102 6830 -12068
rect 6772 -12161 6830 -12102
rect 6772 -12195 6784 -12161
rect 6818 -12195 6830 -12161
rect 6084 -12261 6154 -12232
rect 5847 -12309 5863 -12275
rect 5897 -12309 6019 -12275
rect 5847 -12310 6019 -12309
rect 5779 -12344 5813 -12325
rect 5779 -12378 5897 -12344
rect 5576 -12420 5657 -12396
rect 5576 -12454 5609 -12420
rect 5643 -12454 5657 -12420
rect 5576 -12473 5657 -12454
rect 5691 -12420 5757 -12404
rect 5691 -12454 5707 -12420
rect 5741 -12454 5757 -12420
rect 5691 -12507 5757 -12454
rect 5847 -12420 5897 -12378
rect 5847 -12454 5863 -12420
rect 5847 -12473 5897 -12454
rect 5949 -12420 6019 -12310
rect 6068 -12275 6154 -12261
rect 6068 -12309 6084 -12275
rect 6118 -12309 6154 -12275
rect 6188 -12268 6278 -12266
rect 6188 -12302 6202 -12268
rect 6236 -12275 6278 -12268
rect 6188 -12309 6204 -12302
rect 6238 -12309 6278 -12275
rect 6404 -12285 6554 -12215
rect 6772 -12230 6830 -12195
rect 6864 -12039 7566 -11997
rect 6864 -12073 6882 -12039
rect 6916 -12073 7514 -12039
rect 7548 -12073 7566 -12039
rect 6864 -12141 7566 -12073
rect 6864 -12175 6882 -12141
rect 6916 -12175 7514 -12141
rect 7548 -12175 7566 -12141
rect 6864 -12215 7566 -12175
rect 6068 -12319 6154 -12309
rect 6404 -12319 6424 -12285
rect 6458 -12319 6554 -12285
rect 6588 -12283 6684 -12249
rect 6718 -12283 6738 -12249
rect 6084 -12343 6154 -12319
rect 6084 -12377 6278 -12343
rect 6588 -12353 6738 -12283
rect 5949 -12454 5968 -12420
rect 6002 -12454 6019 -12420
rect 5949 -12473 6019 -12454
rect 6112 -12420 6178 -12411
rect 6112 -12454 6128 -12420
rect 6162 -12454 6178 -12420
rect 6112 -12507 6178 -12454
rect 6212 -12420 6278 -12377
rect 6212 -12454 6225 -12420
rect 6259 -12454 6278 -12420
rect 6212 -12473 6278 -12454
rect 6312 -12379 6370 -12362
rect 6312 -12413 6324 -12379
rect 6358 -12413 6370 -12379
rect 6312 -12507 6370 -12413
rect 6404 -12405 6738 -12353
rect 6864 -12283 6942 -12249
rect 6976 -12283 7041 -12249
rect 7075 -12283 7140 -12249
rect 7174 -12283 7194 -12249
rect 6864 -12353 7194 -12283
rect 7228 -12285 7566 -12215
rect 7600 -12068 7658 -11997
rect 7600 -12102 7612 -12068
rect 7646 -12102 7658 -12068
rect 7600 -12161 7658 -12102
rect 7600 -12195 7612 -12161
rect 7646 -12195 7658 -12161
rect 7600 -12230 7658 -12195
rect 7692 -12039 8026 -11997
rect 7692 -12073 7710 -12039
rect 7744 -12073 7974 -12039
rect 8008 -12073 8026 -12039
rect 7692 -12141 8026 -12073
rect 7692 -12175 7710 -12141
rect 7744 -12175 7974 -12141
rect 8008 -12175 8026 -12141
rect 7692 -12215 8026 -12175
rect 8060 -12068 8118 -11997
rect 8060 -12102 8072 -12068
rect 8106 -12102 8118 -12068
rect 8060 -12161 8118 -12102
rect 8060 -12195 8072 -12161
rect 8106 -12195 8118 -12161
rect 7228 -12319 7248 -12285
rect 7282 -12319 7351 -12285
rect 7385 -12319 7454 -12285
rect 7488 -12319 7566 -12285
rect 7692 -12285 7842 -12215
rect 8060 -12230 8118 -12195
rect 8152 -12047 8233 -12031
rect 8152 -12081 8185 -12047
rect 8219 -12081 8233 -12047
rect 8152 -12115 8233 -12081
rect 8152 -12149 8185 -12115
rect 8219 -12149 8233 -12115
rect 8152 -12186 8233 -12149
rect 8267 -12046 8333 -11997
rect 8267 -12080 8283 -12046
rect 8317 -12080 8333 -12046
rect 8267 -12114 8333 -12080
rect 8267 -12148 8283 -12114
rect 8317 -12148 8333 -12114
rect 8267 -12157 8333 -12148
rect 8423 -12047 8473 -12031
rect 8423 -12081 8439 -12047
rect 8423 -12115 8473 -12081
rect 8423 -12149 8439 -12115
rect 7692 -12319 7712 -12285
rect 7746 -12319 7842 -12285
rect 7876 -12283 7972 -12249
rect 8006 -12283 8026 -12249
rect 7876 -12353 8026 -12283
rect 6404 -12439 6422 -12405
rect 6456 -12439 6686 -12405
rect 6720 -12439 6738 -12405
rect 6404 -12507 6738 -12439
rect 6772 -12379 6830 -12362
rect 6772 -12413 6784 -12379
rect 6818 -12413 6830 -12379
rect 6772 -12507 6830 -12413
rect 6864 -12412 7566 -12353
rect 6864 -12446 6882 -12412
rect 6916 -12446 7514 -12412
rect 7548 -12446 7566 -12412
rect 6864 -12507 7566 -12446
rect 7600 -12379 7658 -12362
rect 7600 -12413 7612 -12379
rect 7646 -12413 7658 -12379
rect 7600 -12507 7658 -12413
rect 7692 -12405 8026 -12353
rect 8152 -12268 8202 -12186
rect 8423 -12191 8473 -12149
rect 8355 -12225 8473 -12191
rect 8525 -12046 8595 -12031
rect 8525 -12080 8543 -12046
rect 8577 -12080 8595 -12046
rect 8525 -12114 8595 -12080
rect 8525 -12148 8543 -12114
rect 8577 -12148 8595 -12114
rect 8355 -12259 8389 -12225
rect 8152 -12302 8162 -12268
rect 8196 -12302 8202 -12268
rect 7692 -12439 7710 -12405
rect 7744 -12439 7974 -12405
rect 8008 -12439 8026 -12405
rect 7692 -12507 8026 -12439
rect 8060 -12379 8118 -12362
rect 8060 -12413 8072 -12379
rect 8106 -12413 8118 -12379
rect 8060 -12507 8118 -12413
rect 8152 -12396 8202 -12302
rect 8236 -12275 8389 -12259
rect 8525 -12260 8595 -12148
rect 8685 -12046 8751 -11997
rect 8685 -12080 8701 -12046
rect 8735 -12080 8751 -12046
rect 8685 -12114 8751 -12080
rect 8685 -12148 8701 -12114
rect 8735 -12148 8751 -12114
rect 8685 -12164 8751 -12148
rect 8785 -12046 8854 -12031
rect 8785 -12080 8801 -12046
rect 8835 -12080 8854 -12046
rect 8785 -12114 8854 -12080
rect 8785 -12148 8801 -12114
rect 8835 -12148 8854 -12114
rect 8785 -12198 8854 -12148
rect 8236 -12309 8239 -12275
rect 8273 -12309 8389 -12275
rect 8236 -12325 8389 -12309
rect 8423 -12275 8595 -12260
rect 8660 -12232 8854 -12198
rect 8888 -12068 8946 -11997
rect 8888 -12102 8900 -12068
rect 8934 -12102 8946 -12068
rect 8888 -12161 8946 -12102
rect 8888 -12195 8900 -12161
rect 8934 -12195 8946 -12161
rect 8888 -12230 8946 -12195
rect 8980 -12039 9314 -11997
rect 8980 -12073 8998 -12039
rect 9032 -12073 9262 -12039
rect 9296 -12073 9314 -12039
rect 8980 -12141 9314 -12073
rect 8980 -12175 8998 -12141
rect 9032 -12175 9262 -12141
rect 9296 -12175 9314 -12141
rect 8980 -12215 9314 -12175
rect 9348 -12068 9406 -11997
rect 9348 -12102 9360 -12068
rect 9394 -12102 9406 -12068
rect 9348 -12161 9406 -12102
rect 9348 -12195 9360 -12161
rect 9394 -12195 9406 -12161
rect 8660 -12261 8730 -12232
rect 8423 -12309 8439 -12275
rect 8473 -12309 8595 -12275
rect 8423 -12310 8595 -12309
rect 8355 -12344 8389 -12325
rect 8355 -12378 8473 -12344
rect 8152 -12420 8233 -12396
rect 8152 -12454 8185 -12420
rect 8219 -12454 8233 -12420
rect 8152 -12473 8233 -12454
rect 8267 -12420 8333 -12404
rect 8267 -12454 8283 -12420
rect 8317 -12454 8333 -12420
rect 8267 -12507 8333 -12454
rect 8423 -12420 8473 -12378
rect 8423 -12454 8439 -12420
rect 8423 -12473 8473 -12454
rect 8525 -12420 8595 -12310
rect 8644 -12275 8730 -12261
rect 8644 -12309 8660 -12275
rect 8694 -12309 8730 -12275
rect 8764 -12268 8854 -12266
rect 8764 -12302 8776 -12268
rect 8810 -12275 8854 -12268
rect 8764 -12309 8780 -12302
rect 8814 -12309 8854 -12275
rect 8980 -12285 9130 -12215
rect 9348 -12230 9406 -12195
rect 9440 -12039 10142 -11997
rect 9440 -12073 9458 -12039
rect 9492 -12073 10090 -12039
rect 10124 -12073 10142 -12039
rect 9440 -12141 10142 -12073
rect 9440 -12175 9458 -12141
rect 9492 -12175 10090 -12141
rect 10124 -12175 10142 -12141
rect 9440 -12215 10142 -12175
rect 8644 -12319 8730 -12309
rect 8980 -12319 9000 -12285
rect 9034 -12319 9130 -12285
rect 9164 -12283 9260 -12249
rect 9294 -12283 9314 -12249
rect 8660 -12343 8730 -12319
rect 8660 -12377 8854 -12343
rect 9164 -12353 9314 -12283
rect 8525 -12454 8544 -12420
rect 8578 -12454 8595 -12420
rect 8525 -12473 8595 -12454
rect 8688 -12420 8754 -12411
rect 8688 -12454 8704 -12420
rect 8738 -12454 8754 -12420
rect 8688 -12507 8754 -12454
rect 8788 -12420 8854 -12377
rect 8788 -12454 8801 -12420
rect 8835 -12454 8854 -12420
rect 8788 -12473 8854 -12454
rect 8888 -12379 8946 -12362
rect 8888 -12413 8900 -12379
rect 8934 -12413 8946 -12379
rect 8888 -12507 8946 -12413
rect 8980 -12405 9314 -12353
rect 9440 -12283 9518 -12249
rect 9552 -12283 9617 -12249
rect 9651 -12283 9716 -12249
rect 9750 -12283 9770 -12249
rect 9440 -12353 9770 -12283
rect 9804 -12285 10142 -12215
rect 10176 -12068 10234 -11997
rect 10176 -12102 10188 -12068
rect 10222 -12102 10234 -12068
rect 10176 -12161 10234 -12102
rect 10176 -12195 10188 -12161
rect 10222 -12195 10234 -12161
rect 10176 -12230 10234 -12195
rect 10360 -12039 10694 -11997
rect 10360 -12073 10378 -12039
rect 10412 -12073 10642 -12039
rect 10676 -12073 10694 -12039
rect 10360 -12141 10694 -12073
rect 10360 -12175 10378 -12141
rect 10412 -12175 10642 -12141
rect 10676 -12175 10694 -12141
rect 10360 -12215 10694 -12175
rect 10728 -12047 10809 -12031
rect 10728 -12081 10761 -12047
rect 10795 -12081 10809 -12047
rect 10728 -12115 10809 -12081
rect 10728 -12149 10761 -12115
rect 10795 -12149 10809 -12115
rect 10728 -12186 10809 -12149
rect 10843 -12046 10909 -11997
rect 10843 -12080 10859 -12046
rect 10893 -12080 10909 -12046
rect 10843 -12114 10909 -12080
rect 10843 -12148 10859 -12114
rect 10893 -12148 10909 -12114
rect 10843 -12157 10909 -12148
rect 10999 -12047 11049 -12031
rect 10999 -12081 11015 -12047
rect 10999 -12115 11049 -12081
rect 10999 -12149 11015 -12115
rect 9804 -12319 9824 -12285
rect 9858 -12319 9927 -12285
rect 9961 -12319 10030 -12285
rect 10064 -12319 10142 -12285
rect 10360 -12285 10510 -12215
rect 10360 -12319 10380 -12285
rect 10414 -12319 10510 -12285
rect 10544 -12283 10640 -12249
rect 10674 -12283 10694 -12249
rect 10544 -12353 10694 -12283
rect 8980 -12439 8998 -12405
rect 9032 -12439 9262 -12405
rect 9296 -12439 9314 -12405
rect 8980 -12507 9314 -12439
rect 9348 -12379 9406 -12362
rect 9348 -12413 9360 -12379
rect 9394 -12413 9406 -12379
rect 9348 -12507 9406 -12413
rect 9440 -12412 10142 -12353
rect 9440 -12446 9458 -12412
rect 9492 -12446 10090 -12412
rect 10124 -12446 10142 -12412
rect 9440 -12507 10142 -12446
rect 10176 -12379 10234 -12362
rect 10176 -12413 10188 -12379
rect 10222 -12413 10234 -12379
rect 10176 -12507 10234 -12413
rect 10360 -12405 10694 -12353
rect 10360 -12439 10378 -12405
rect 10412 -12439 10642 -12405
rect 10676 -12439 10694 -12405
rect 10360 -12507 10694 -12439
rect 10728 -12268 10778 -12186
rect 10999 -12191 11049 -12149
rect 10931 -12225 11049 -12191
rect 11101 -12046 11171 -12031
rect 11101 -12080 11119 -12046
rect 11153 -12080 11171 -12046
rect 11101 -12114 11171 -12080
rect 11101 -12148 11119 -12114
rect 11153 -12148 11171 -12114
rect 10931 -12259 10965 -12225
rect 10728 -12302 10736 -12268
rect 10770 -12302 10778 -12268
rect 10728 -12396 10778 -12302
rect 10812 -12275 10965 -12259
rect 11101 -12260 11171 -12148
rect 11261 -12046 11327 -11997
rect 11261 -12080 11277 -12046
rect 11311 -12080 11327 -12046
rect 11261 -12114 11327 -12080
rect 11261 -12148 11277 -12114
rect 11311 -12148 11327 -12114
rect 11261 -12164 11327 -12148
rect 11361 -12046 11430 -12031
rect 11361 -12080 11377 -12046
rect 11411 -12080 11430 -12046
rect 11361 -12114 11430 -12080
rect 11361 -12148 11377 -12114
rect 11411 -12148 11430 -12114
rect 11361 -12198 11430 -12148
rect 10812 -12309 10815 -12275
rect 10849 -12309 10965 -12275
rect 10812 -12325 10965 -12309
rect 10999 -12275 11171 -12260
rect 11236 -12232 11430 -12198
rect 11464 -12068 11522 -11997
rect 11464 -12102 11476 -12068
rect 11510 -12102 11522 -12068
rect 11464 -12161 11522 -12102
rect 11464 -12195 11476 -12161
rect 11510 -12195 11522 -12161
rect 11464 -12230 11522 -12195
rect 11648 -12039 11982 -11997
rect 11648 -12073 11666 -12039
rect 11700 -12073 11930 -12039
rect 11964 -12073 11982 -12039
rect 11648 -12141 11982 -12073
rect 11648 -12175 11666 -12141
rect 11700 -12175 11930 -12141
rect 11964 -12175 11982 -12141
rect 11648 -12215 11982 -12175
rect 13580 -12068 13638 -11997
rect 13580 -12102 13592 -12068
rect 13626 -12102 13638 -12068
rect 13580 -12161 13638 -12102
rect 13674 -12039 13733 -11997
rect 13674 -12073 13690 -12039
rect 13724 -12073 13733 -12039
rect 13674 -12107 13733 -12073
rect 13674 -12141 13690 -12107
rect 13724 -12141 13733 -12107
rect 13674 -12159 13733 -12141
rect 13769 -12047 13818 -12031
rect 13769 -12081 13776 -12047
rect 13810 -12081 13818 -12047
rect 13769 -12115 13818 -12081
rect 13769 -12149 13776 -12115
rect 13810 -12149 13818 -12115
rect 13580 -12195 13592 -12161
rect 13626 -12195 13638 -12161
rect 11236 -12261 11306 -12232
rect 10999 -12309 11015 -12275
rect 11049 -12309 11171 -12275
rect 10999 -12310 11171 -12309
rect 10931 -12344 10965 -12325
rect 10931 -12378 11049 -12344
rect 10728 -12420 10809 -12396
rect 10728 -12454 10761 -12420
rect 10795 -12454 10809 -12420
rect 10728 -12473 10809 -12454
rect 10843 -12420 10909 -12404
rect 10843 -12454 10859 -12420
rect 10893 -12454 10909 -12420
rect 10843 -12507 10909 -12454
rect 10999 -12420 11049 -12378
rect 10999 -12454 11015 -12420
rect 10999 -12473 11049 -12454
rect 11101 -12420 11171 -12310
rect 11220 -12275 11306 -12261
rect 11220 -12309 11236 -12275
rect 11270 -12309 11306 -12275
rect 11340 -12273 11430 -12266
rect 11340 -12275 11384 -12273
rect 11340 -12309 11356 -12275
rect 11418 -12307 11430 -12273
rect 11390 -12309 11430 -12307
rect 11648 -12285 11798 -12215
rect 13580 -12230 13638 -12195
rect 11220 -12319 11306 -12309
rect 11648 -12319 11668 -12285
rect 11702 -12319 11798 -12285
rect 11832 -12283 11928 -12249
rect 11962 -12283 11982 -12249
rect 13769 -12259 13818 -12149
rect 13853 -12039 13905 -11997
rect 14025 -11998 15280 -11997
rect 13853 -12073 13862 -12039
rect 13896 -12073 13905 -12039
rect 13853 -12107 13905 -12073
rect 13853 -12141 13862 -12107
rect 13896 -12141 13905 -12107
rect 13853 -12159 13905 -12141
rect 13941 -12055 13991 -12032
rect 13941 -12089 13948 -12055
rect 13982 -12089 13991 -12055
rect 13941 -12123 13991 -12089
rect 13941 -12157 13948 -12123
rect 13982 -12157 13991 -12123
rect 14025 -12039 14077 -11998
rect 14025 -12073 14034 -12039
rect 14068 -12073 14077 -12039
rect 14025 -12107 14077 -12073
rect 14025 -12141 14034 -12107
rect 14068 -12141 14077 -12107
rect 14025 -12157 14077 -12141
rect 14111 -12083 14163 -12032
rect 14111 -12117 14120 -12083
rect 14154 -12117 14163 -12083
rect 13941 -12259 13991 -12157
rect 14111 -12169 14163 -12117
rect 14197 -12063 14249 -11998
rect 14197 -12097 14206 -12063
rect 14240 -12097 14249 -12063
rect 14197 -12143 14249 -12097
rect 14283 -12083 14335 -12032
rect 14283 -12117 14292 -12083
rect 14326 -12117 14335 -12083
rect 14111 -12203 14120 -12169
rect 14154 -12177 14163 -12169
rect 14283 -12169 14335 -12117
rect 14369 -12063 14421 -11998
rect 14369 -12097 14378 -12063
rect 14412 -12097 14421 -12063
rect 14369 -12143 14421 -12097
rect 14455 -12083 14507 -12032
rect 14455 -12117 14464 -12083
rect 14498 -12117 14507 -12083
rect 14283 -12177 14292 -12169
rect 14154 -12203 14292 -12177
rect 14326 -12177 14335 -12169
rect 14455 -12169 14507 -12117
rect 14541 -12063 14593 -11998
rect 14541 -12097 14550 -12063
rect 14584 -12097 14593 -12063
rect 14541 -12143 14593 -12097
rect 14627 -12083 14679 -12032
rect 14627 -12117 14636 -12083
rect 14670 -12117 14679 -12083
rect 14455 -12177 14464 -12169
rect 14326 -12203 14464 -12177
rect 14498 -12177 14507 -12169
rect 14627 -12169 14679 -12117
rect 14713 -12063 14762 -11998
rect 14713 -12097 14722 -12063
rect 14756 -12097 14762 -12063
rect 14713 -12143 14762 -12097
rect 14796 -12083 14848 -12032
rect 14796 -12117 14807 -12083
rect 14841 -12117 14848 -12083
rect 14627 -12177 14636 -12169
rect 14498 -12203 14636 -12177
rect 14670 -12177 14679 -12169
rect 14796 -12169 14848 -12117
rect 14885 -12063 14934 -11998
rect 14885 -12097 14893 -12063
rect 14927 -12097 14934 -12063
rect 14885 -12143 14934 -12097
rect 14968 -12083 15020 -12032
rect 14968 -12117 14979 -12083
rect 15013 -12117 15020 -12083
rect 14796 -12177 14807 -12169
rect 14670 -12203 14807 -12177
rect 14841 -12177 14848 -12169
rect 14968 -12169 15020 -12117
rect 15057 -12063 15106 -11998
rect 15057 -12097 15065 -12063
rect 15099 -12097 15106 -12063
rect 15057 -12143 15106 -12097
rect 15140 -12083 15192 -12032
rect 15140 -12117 15151 -12083
rect 15185 -12117 15192 -12083
rect 14968 -12177 14979 -12169
rect 14841 -12203 14979 -12177
rect 15013 -12177 15020 -12169
rect 15140 -12169 15192 -12117
rect 15229 -12063 15280 -11998
rect 15229 -12097 15237 -12063
rect 15271 -12097 15280 -12063
rect 15229 -12143 15280 -12097
rect 15314 -12083 15372 -12032
rect 15314 -12117 15323 -12083
rect 15357 -12117 15372 -12083
rect 15140 -12177 15151 -12169
rect 15013 -12203 15151 -12177
rect 15185 -12180 15192 -12169
rect 15314 -12169 15372 -12117
rect 15406 -12063 15460 -11997
rect 15406 -12097 15409 -12063
rect 15443 -12097 15460 -12063
rect 15406 -12146 15460 -12097
rect 15512 -12068 15570 -11997
rect 15512 -12102 15524 -12068
rect 15558 -12102 15570 -12068
rect 15314 -12180 15323 -12169
rect 15185 -12203 15323 -12180
rect 15357 -12180 15372 -12169
rect 15512 -12161 15570 -12102
rect 15357 -12203 15460 -12180
rect 14111 -12222 15460 -12203
rect 14111 -12225 15248 -12222
rect 15227 -12256 15248 -12225
rect 15282 -12256 15341 -12222
rect 15375 -12256 15460 -12222
rect 15512 -12195 15524 -12161
rect 15558 -12195 15570 -12161
rect 15512 -12230 15570 -12195
rect 15605 -12039 16674 -11997
rect 15605 -12073 15622 -12039
rect 15656 -12073 16622 -12039
rect 16656 -12073 16674 -12039
rect 15605 -12141 16674 -12073
rect 15605 -12175 15622 -12141
rect 15656 -12175 16622 -12141
rect 16656 -12175 16674 -12141
rect 15605 -12215 16674 -12175
rect 11236 -12343 11306 -12319
rect 11236 -12377 11430 -12343
rect 11832 -12353 11982 -12283
rect 11101 -12454 11120 -12420
rect 11154 -12454 11171 -12420
rect 11101 -12473 11171 -12454
rect 11264 -12420 11330 -12411
rect 11264 -12454 11280 -12420
rect 11314 -12454 11330 -12420
rect 11264 -12507 11330 -12454
rect 11364 -12420 11430 -12377
rect 11364 -12454 11377 -12420
rect 11411 -12454 11430 -12420
rect 11364 -12473 11430 -12454
rect 11464 -12379 11522 -12362
rect 11464 -12413 11476 -12379
rect 11510 -12413 11522 -12379
rect 11464 -12507 11522 -12413
rect 11648 -12405 11982 -12353
rect 13672 -12275 13735 -12259
rect 13672 -12302 13692 -12275
rect 13672 -12336 13685 -12302
rect 13726 -12309 13735 -12275
rect 13719 -12336 13735 -12309
rect 11648 -12439 11666 -12405
rect 11700 -12439 11930 -12405
rect 11964 -12439 11982 -12405
rect 11648 -12507 11982 -12439
rect 13580 -12379 13638 -12362
rect 13672 -12371 13735 -12336
rect 13769 -12275 15193 -12259
rect 13769 -12309 14119 -12275
rect 14153 -12309 14187 -12275
rect 14221 -12309 14255 -12275
rect 14289 -12309 14323 -12275
rect 14357 -12309 14391 -12275
rect 14425 -12309 14459 -12275
rect 14493 -12309 14527 -12275
rect 14561 -12309 14595 -12275
rect 14629 -12309 14663 -12275
rect 14697 -12309 14731 -12275
rect 14765 -12309 14799 -12275
rect 14833 -12309 14867 -12275
rect 14901 -12309 14935 -12275
rect 14969 -12309 15003 -12275
rect 15037 -12309 15071 -12275
rect 15105 -12309 15139 -12275
rect 15173 -12309 15193 -12275
rect 13580 -12413 13592 -12379
rect 13626 -12413 13638 -12379
rect 13580 -12507 13638 -12413
rect 13672 -12431 13733 -12405
rect 13672 -12465 13690 -12431
rect 13724 -12465 13733 -12431
rect 13672 -12507 13733 -12465
rect 13769 -12418 13819 -12309
rect 13769 -12452 13776 -12418
rect 13810 -12452 13819 -12418
rect 13769 -12471 13819 -12452
rect 13853 -12418 13905 -12402
rect 13853 -12452 13862 -12418
rect 13896 -12452 13905 -12418
rect 13853 -12507 13905 -12452
rect 13941 -12418 13991 -12309
rect 15227 -12317 15460 -12256
rect 15227 -12318 15340 -12317
rect 15227 -12343 15248 -12318
rect 14111 -12352 15248 -12343
rect 15282 -12351 15340 -12318
rect 15374 -12351 15460 -12317
rect 15605 -12285 16124 -12215
rect 15605 -12319 15686 -12285
rect 15720 -12319 15814 -12285
rect 15848 -12319 15942 -12285
rect 15976 -12319 16070 -12285
rect 16104 -12319 16124 -12285
rect 16158 -12283 16178 -12249
rect 16212 -12283 16306 -12249
rect 16340 -12283 16434 -12249
rect 16468 -12283 16562 -12249
rect 16596 -12283 16674 -12249
rect 15282 -12352 15460 -12351
rect 14111 -12377 15460 -12352
rect 16158 -12353 16674 -12283
rect 13941 -12452 13948 -12418
rect 13982 -12452 13991 -12418
rect 13941 -12471 13991 -12452
rect 14025 -12418 14077 -12395
rect 14025 -12452 14034 -12418
rect 14068 -12452 14077 -12418
rect 14025 -12507 14077 -12452
rect 14111 -12418 14163 -12377
rect 14111 -12452 14120 -12418
rect 14154 -12452 14163 -12418
rect 14111 -12468 14163 -12452
rect 14197 -12427 14249 -12411
rect 14197 -12461 14206 -12427
rect 14240 -12461 14249 -12427
rect 14197 -12507 14249 -12461
rect 14283 -12418 14335 -12377
rect 14283 -12452 14292 -12418
rect 14326 -12452 14335 -12418
rect 14283 -12468 14335 -12452
rect 14369 -12427 14421 -12411
rect 14369 -12461 14378 -12427
rect 14412 -12461 14421 -12427
rect 14369 -12507 14421 -12461
rect 14455 -12418 14507 -12377
rect 14455 -12452 14464 -12418
rect 14498 -12452 14507 -12418
rect 14455 -12468 14507 -12452
rect 14541 -12427 14590 -12411
rect 14541 -12461 14550 -12427
rect 14584 -12461 14590 -12427
rect 14541 -12507 14590 -12461
rect 14624 -12418 14679 -12377
rect 14624 -12452 14636 -12418
rect 14670 -12452 14679 -12418
rect 14624 -12468 14679 -12452
rect 14713 -12427 14762 -12411
rect 14713 -12461 14722 -12427
rect 14756 -12461 14762 -12427
rect 14713 -12507 14762 -12461
rect 14796 -12418 14848 -12377
rect 14796 -12452 14807 -12418
rect 14841 -12452 14848 -12418
rect 14796 -12468 14848 -12452
rect 14884 -12427 14934 -12411
rect 14884 -12461 14893 -12427
rect 14927 -12461 14934 -12427
rect 14884 -12507 14934 -12461
rect 14968 -12418 15020 -12377
rect 14968 -12452 14979 -12418
rect 15013 -12452 15020 -12418
rect 14968 -12468 15020 -12452
rect 15056 -12427 15106 -12411
rect 15056 -12461 15065 -12427
rect 15099 -12461 15106 -12427
rect 15056 -12507 15106 -12461
rect 15140 -12418 15192 -12377
rect 15140 -12452 15151 -12418
rect 15185 -12452 15192 -12418
rect 15140 -12468 15192 -12452
rect 15228 -12427 15280 -12411
rect 15228 -12461 15237 -12427
rect 15271 -12461 15280 -12427
rect 15228 -12507 15280 -12461
rect 15314 -12418 15366 -12377
rect 15512 -12379 15570 -12362
rect 15314 -12452 15323 -12418
rect 15357 -12452 15366 -12418
rect 15314 -12468 15366 -12452
rect 15400 -12427 15460 -12411
rect 15400 -12461 15409 -12427
rect 15443 -12461 15460 -12427
rect 15400 -12507 15460 -12461
rect 15512 -12413 15524 -12379
rect 15558 -12413 15570 -12379
rect 15512 -12507 15570 -12413
rect 15605 -12412 16674 -12353
rect 15605 -12446 15622 -12412
rect 15656 -12446 16622 -12412
rect 16656 -12446 16674 -12412
rect 15605 -12507 16674 -12446
rect -2997 -12541 -2968 -12507
rect -2934 -12541 -2876 -12507
rect -2842 -12541 -2784 -12507
rect -2750 -12541 -2692 -12507
rect -2658 -12541 -2600 -12507
rect -2566 -12541 -2508 -12507
rect -2474 -12541 -2416 -12507
rect -2382 -12541 -2324 -12507
rect -2290 -12541 -2232 -12507
rect -2198 -12541 -2140 -12507
rect -2106 -12541 -2048 -12507
rect -2014 -12541 -1956 -12507
rect -1922 -12541 -1864 -12507
rect -1830 -12541 -1772 -12507
rect -1738 -12541 -1680 -12507
rect -1646 -12541 -1588 -12507
rect -1554 -12541 -1496 -12507
rect -1462 -12541 -1404 -12507
rect -1370 -12541 -1312 -12507
rect -1278 -12541 -1220 -12507
rect -1186 -12541 -1128 -12507
rect -1094 -12541 -1036 -12507
rect -1002 -12541 -944 -12507
rect -910 -12541 -852 -12507
rect -818 -12541 -760 -12507
rect -726 -12541 -668 -12507
rect -634 -12541 -576 -12507
rect -542 -12541 -484 -12507
rect -450 -12541 -392 -12507
rect -358 -12541 -300 -12507
rect -266 -12541 -208 -12507
rect -174 -12541 -116 -12507
rect -82 -12541 -24 -12507
rect 10 -12541 68 -12507
rect 102 -12541 160 -12507
rect 194 -12541 252 -12507
rect 286 -12541 344 -12507
rect 378 -12541 436 -12507
rect 470 -12541 528 -12507
rect 562 -12541 620 -12507
rect 654 -12541 712 -12507
rect 746 -12541 804 -12507
rect 838 -12541 896 -12507
rect 930 -12541 988 -12507
rect 1022 -12541 1080 -12507
rect 1114 -12541 1172 -12507
rect 1206 -12541 1264 -12507
rect 1298 -12541 1356 -12507
rect 1390 -12541 1448 -12507
rect 1482 -12541 1540 -12507
rect 1574 -12541 1632 -12507
rect 1666 -12541 1724 -12507
rect 1758 -12541 1816 -12507
rect 1850 -12541 1908 -12507
rect 1942 -12541 2000 -12507
rect 2034 -12541 2092 -12507
rect 2126 -12541 2184 -12507
rect 2218 -12541 2276 -12507
rect 2310 -12541 2368 -12507
rect 2402 -12541 2460 -12507
rect 2494 -12541 2552 -12507
rect 2586 -12541 2644 -12507
rect 2678 -12541 2736 -12507
rect 2770 -12541 2828 -12507
rect 2862 -12541 2920 -12507
rect 2954 -12541 3012 -12507
rect 3046 -12541 3104 -12507
rect 3138 -12541 3196 -12507
rect 3230 -12541 3288 -12507
rect 3322 -12541 3380 -12507
rect 3414 -12541 3472 -12507
rect 3506 -12541 3564 -12507
rect 3598 -12541 3656 -12507
rect 3690 -12541 3748 -12507
rect 3782 -12541 3840 -12507
rect 3874 -12541 3932 -12507
rect 3966 -12541 4024 -12507
rect 4058 -12541 4116 -12507
rect 4150 -12541 4208 -12507
rect 4242 -12541 4300 -12507
rect 4334 -12541 4392 -12507
rect 4426 -12541 4484 -12507
rect 4518 -12541 4576 -12507
rect 4610 -12541 4668 -12507
rect 4702 -12541 4760 -12507
rect 4794 -12541 4852 -12507
rect 4886 -12541 4944 -12507
rect 4978 -12541 5036 -12507
rect 5070 -12541 5128 -12507
rect 5162 -12541 5220 -12507
rect 5254 -12541 5312 -12507
rect 5346 -12541 5404 -12507
rect 5438 -12541 5496 -12507
rect 5530 -12541 5588 -12507
rect 5622 -12541 5680 -12507
rect 5714 -12541 5772 -12507
rect 5806 -12541 5864 -12507
rect 5898 -12541 5956 -12507
rect 5990 -12541 6048 -12507
rect 6082 -12541 6140 -12507
rect 6174 -12541 6232 -12507
rect 6266 -12541 6324 -12507
rect 6358 -12541 6416 -12507
rect 6450 -12541 6508 -12507
rect 6542 -12541 6600 -12507
rect 6634 -12541 6692 -12507
rect 6726 -12541 6784 -12507
rect 6818 -12541 6876 -12507
rect 6910 -12541 6968 -12507
rect 7002 -12541 7060 -12507
rect 7094 -12541 7152 -12507
rect 7186 -12541 7244 -12507
rect 7278 -12541 7336 -12507
rect 7370 -12541 7428 -12507
rect 7462 -12541 7520 -12507
rect 7554 -12541 7612 -12507
rect 7646 -12541 7704 -12507
rect 7738 -12541 7796 -12507
rect 7830 -12541 7888 -12507
rect 7922 -12541 7980 -12507
rect 8014 -12541 8072 -12507
rect 8106 -12541 8164 -12507
rect 8198 -12541 8256 -12507
rect 8290 -12541 8348 -12507
rect 8382 -12541 8440 -12507
rect 8474 -12541 8532 -12507
rect 8566 -12541 8624 -12507
rect 8658 -12541 8716 -12507
rect 8750 -12541 8808 -12507
rect 8842 -12541 8900 -12507
rect 8934 -12541 8992 -12507
rect 9026 -12541 9084 -12507
rect 9118 -12541 9176 -12507
rect 9210 -12541 9268 -12507
rect 9302 -12541 9360 -12507
rect 9394 -12541 9452 -12507
rect 9486 -12541 9544 -12507
rect 9578 -12541 9636 -12507
rect 9670 -12541 9728 -12507
rect 9762 -12541 9820 -12507
rect 9854 -12541 9912 -12507
rect 9946 -12541 10004 -12507
rect 10038 -12541 10096 -12507
rect 10130 -12541 10188 -12507
rect 10222 -12541 10280 -12507
rect 10314 -12541 10372 -12507
rect 10406 -12541 10464 -12507
rect 10498 -12541 10556 -12507
rect 10590 -12541 10648 -12507
rect 10682 -12541 10740 -12507
rect 10774 -12541 10832 -12507
rect 10866 -12541 10924 -12507
rect 10958 -12541 11016 -12507
rect 11050 -12541 11108 -12507
rect 11142 -12541 11200 -12507
rect 11234 -12541 11292 -12507
rect 11326 -12541 11384 -12507
rect 11418 -12541 11476 -12507
rect 11510 -12541 11568 -12507
rect 11602 -12541 11660 -12507
rect 11694 -12541 11752 -12507
rect 11786 -12541 11844 -12507
rect 11878 -12541 11936 -12507
rect 11970 -12541 12028 -12507
rect 12062 -12541 12120 -12507
rect 12154 -12541 12212 -12507
rect 12246 -12541 12304 -12507
rect 12338 -12541 12396 -12507
rect 12430 -12541 12488 -12507
rect 12522 -12541 12580 -12507
rect 12614 -12541 12672 -12507
rect 12706 -12541 12764 -12507
rect 12798 -12541 12856 -12507
rect 12890 -12541 12948 -12507
rect 12982 -12541 13040 -12507
rect 13074 -12541 13132 -12507
rect 13166 -12541 13224 -12507
rect 13258 -12541 13316 -12507
rect 13350 -12541 13408 -12507
rect 13442 -12541 13500 -12507
rect 13534 -12541 13592 -12507
rect 13626 -12541 13684 -12507
rect 13718 -12541 13776 -12507
rect 13810 -12541 13868 -12507
rect 13902 -12541 13960 -12507
rect 13994 -12541 14052 -12507
rect 14086 -12541 14144 -12507
rect 14178 -12541 14236 -12507
rect 14270 -12541 14328 -12507
rect 14362 -12541 14420 -12507
rect 14454 -12541 14512 -12507
rect 14546 -12541 14604 -12507
rect 14638 -12541 14696 -12507
rect 14730 -12541 14788 -12507
rect 14822 -12541 14880 -12507
rect 14914 -12541 14972 -12507
rect 15006 -12541 15064 -12507
rect 15098 -12541 15156 -12507
rect 15190 -12541 15248 -12507
rect 15282 -12541 15340 -12507
rect 15374 -12541 15432 -12507
rect 15466 -12541 15524 -12507
rect 15558 -12541 15616 -12507
rect 15650 -12541 15708 -12507
rect 15742 -12541 15800 -12507
rect 15834 -12541 15892 -12507
rect 15926 -12541 15984 -12507
rect 16018 -12541 16076 -12507
rect 16110 -12541 16168 -12507
rect 16202 -12541 16260 -12507
rect 16294 -12541 16352 -12507
rect 16386 -12541 16444 -12507
rect 16478 -12541 16536 -12507
rect 16570 -12541 16628 -12507
rect 16662 -12541 16691 -12507
rect -2980 -12602 -2278 -12541
rect -2980 -12636 -2962 -12602
rect -2928 -12636 -2330 -12602
rect -2296 -12636 -2278 -12602
rect -2980 -12695 -2278 -12636
rect -2244 -12635 -2186 -12541
rect -2244 -12669 -2232 -12635
rect -2198 -12669 -2186 -12635
rect -2244 -12686 -2186 -12669
rect -1600 -12602 -898 -12541
rect -1600 -12636 -1582 -12602
rect -1548 -12636 -950 -12602
rect -916 -12636 -898 -12602
rect -2980 -12763 -2902 -12729
rect -2868 -12763 -2799 -12729
rect -2765 -12763 -2696 -12729
rect -2662 -12763 -2642 -12729
rect -2980 -12833 -2642 -12763
rect -2608 -12765 -2278 -12695
rect -2608 -12799 -2588 -12765
rect -2554 -12799 -2489 -12765
rect -2455 -12799 -2390 -12765
rect -2356 -12799 -2278 -12765
rect -1600 -12695 -898 -12636
rect -864 -12602 -162 -12541
rect -864 -12636 -846 -12602
rect -812 -12636 -214 -12602
rect -180 -12636 -162 -12602
rect -864 -12695 -162 -12636
rect -128 -12635 -70 -12541
rect -128 -12669 -116 -12635
rect -82 -12669 -70 -12635
rect -128 -12686 -70 -12669
rect -36 -12609 298 -12541
rect -36 -12643 -18 -12609
rect 16 -12643 246 -12609
rect 280 -12643 298 -12609
rect -36 -12695 298 -12643
rect 332 -12635 390 -12541
rect 332 -12669 344 -12635
rect 378 -12669 390 -12635
rect 332 -12686 390 -12669
rect 424 -12594 490 -12575
rect 424 -12628 443 -12594
rect 477 -12628 490 -12594
rect 424 -12671 490 -12628
rect 524 -12594 590 -12541
rect 524 -12628 540 -12594
rect 574 -12628 590 -12594
rect 524 -12637 590 -12628
rect 683 -12594 753 -12575
rect 683 -12628 700 -12594
rect 734 -12628 753 -12594
rect -1600 -12765 -1270 -12695
rect -1600 -12799 -1522 -12765
rect -1488 -12799 -1423 -12765
rect -1389 -12799 -1324 -12765
rect -1290 -12799 -1270 -12765
rect -1236 -12763 -1216 -12729
rect -1182 -12763 -1113 -12729
rect -1079 -12763 -1010 -12729
rect -976 -12763 -898 -12729
rect -2980 -12873 -2278 -12833
rect -2980 -12907 -2962 -12873
rect -2928 -12907 -2330 -12873
rect -2296 -12907 -2278 -12873
rect -2980 -12975 -2278 -12907
rect -2980 -13009 -2962 -12975
rect -2928 -13009 -2330 -12975
rect -2296 -13009 -2278 -12975
rect -2980 -13051 -2278 -13009
rect -2244 -12853 -2186 -12818
rect -1236 -12833 -898 -12763
rect -864 -12765 -534 -12695
rect -864 -12799 -786 -12765
rect -752 -12799 -687 -12765
rect -653 -12799 -588 -12765
rect -554 -12799 -534 -12765
rect -500 -12763 -480 -12729
rect -446 -12763 -377 -12729
rect -343 -12763 -274 -12729
rect -240 -12763 -162 -12729
rect -500 -12833 -162 -12763
rect -36 -12763 -16 -12729
rect 18 -12763 114 -12729
rect -2244 -12887 -2232 -12853
rect -2198 -12887 -2186 -12853
rect -2244 -12946 -2186 -12887
rect -2244 -12980 -2232 -12946
rect -2198 -12980 -2186 -12946
rect -2244 -13051 -2186 -12980
rect -1600 -12873 -898 -12833
rect -1600 -12907 -1582 -12873
rect -1548 -12907 -950 -12873
rect -916 -12907 -898 -12873
rect -1600 -12975 -898 -12907
rect -1600 -13009 -1582 -12975
rect -1548 -13009 -950 -12975
rect -916 -13009 -898 -12975
rect -1600 -13051 -898 -13009
rect -864 -12873 -162 -12833
rect -864 -12907 -846 -12873
rect -812 -12907 -214 -12873
rect -180 -12907 -162 -12873
rect -864 -12975 -162 -12907
rect -864 -13009 -846 -12975
rect -812 -13009 -214 -12975
rect -180 -13009 -162 -12975
rect -864 -13051 -162 -13009
rect -128 -12853 -70 -12818
rect -128 -12887 -116 -12853
rect -82 -12887 -70 -12853
rect -128 -12946 -70 -12887
rect -128 -12980 -116 -12946
rect -82 -12980 -70 -12946
rect -128 -13051 -70 -12980
rect -36 -12833 114 -12763
rect 148 -12765 298 -12695
rect 424 -12705 618 -12671
rect 548 -12729 618 -12705
rect 548 -12739 634 -12729
rect 148 -12799 244 -12765
rect 278 -12799 298 -12765
rect 424 -12744 464 -12739
rect 424 -12778 436 -12744
rect 498 -12773 514 -12739
rect 470 -12778 514 -12773
rect 424 -12782 514 -12778
rect 548 -12773 584 -12739
rect 618 -12773 634 -12739
rect 548 -12787 634 -12773
rect 683 -12738 753 -12628
rect 805 -12594 855 -12575
rect 839 -12628 855 -12594
rect 805 -12670 855 -12628
rect 945 -12594 1011 -12541
rect 945 -12628 961 -12594
rect 995 -12628 1011 -12594
rect 945 -12644 1011 -12628
rect 1045 -12594 1126 -12575
rect 1045 -12628 1059 -12594
rect 1093 -12628 1126 -12594
rect 1045 -12652 1126 -12628
rect 805 -12704 923 -12670
rect 889 -12723 923 -12704
rect 683 -12739 855 -12738
rect 683 -12773 805 -12739
rect 839 -12773 855 -12739
rect 548 -12816 618 -12787
rect -36 -12873 298 -12833
rect -36 -12907 -18 -12873
rect 16 -12907 246 -12873
rect 280 -12907 298 -12873
rect -36 -12975 298 -12907
rect -36 -13009 -18 -12975
rect 16 -13009 246 -12975
rect 280 -13009 298 -12975
rect -36 -13051 298 -13009
rect 332 -12853 390 -12818
rect 332 -12887 344 -12853
rect 378 -12887 390 -12853
rect 332 -12946 390 -12887
rect 332 -12980 344 -12946
rect 378 -12980 390 -12946
rect 332 -13051 390 -12980
rect 424 -12850 618 -12816
rect 683 -12788 855 -12773
rect 889 -12739 1042 -12723
rect 889 -12773 1005 -12739
rect 1039 -12773 1042 -12739
rect 424 -12900 493 -12850
rect 424 -12934 443 -12900
rect 477 -12934 493 -12900
rect 424 -12968 493 -12934
rect 424 -13002 443 -12968
rect 477 -13002 493 -12968
rect 424 -13017 493 -13002
rect 527 -12900 593 -12884
rect 527 -12934 543 -12900
rect 577 -12934 593 -12900
rect 527 -12968 593 -12934
rect 527 -13002 543 -12968
rect 577 -13002 593 -12968
rect 527 -13051 593 -13002
rect 683 -12900 753 -12788
rect 889 -12789 1042 -12773
rect 1076 -12745 1126 -12652
rect 1160 -12635 1218 -12541
rect 1160 -12669 1172 -12635
rect 1206 -12669 1218 -12635
rect 1160 -12686 1218 -12669
rect 1252 -12609 1586 -12541
rect 1252 -12643 1270 -12609
rect 1304 -12643 1534 -12609
rect 1568 -12643 1586 -12609
rect 1252 -12695 1586 -12643
rect 1620 -12635 1678 -12541
rect 1620 -12669 1632 -12635
rect 1666 -12669 1678 -12635
rect 1620 -12686 1678 -12669
rect 1712 -12602 2414 -12541
rect 1712 -12636 1730 -12602
rect 1764 -12636 2362 -12602
rect 2396 -12636 2414 -12602
rect 1712 -12695 2414 -12636
rect 2448 -12635 2506 -12541
rect 2448 -12669 2460 -12635
rect 2494 -12669 2506 -12635
rect 2448 -12686 2506 -12669
rect 2540 -12609 2874 -12541
rect 2540 -12643 2558 -12609
rect 2592 -12643 2822 -12609
rect 2856 -12643 2874 -12609
rect 2540 -12695 2874 -12643
rect 2908 -12635 2966 -12541
rect 2908 -12669 2920 -12635
rect 2954 -12669 2966 -12635
rect 2908 -12686 2966 -12669
rect 3000 -12594 3066 -12575
rect 3000 -12628 3019 -12594
rect 3053 -12628 3066 -12594
rect 3000 -12671 3066 -12628
rect 3100 -12594 3166 -12541
rect 3100 -12628 3116 -12594
rect 3150 -12628 3166 -12594
rect 3100 -12637 3166 -12628
rect 3259 -12594 3329 -12575
rect 3259 -12628 3276 -12594
rect 3310 -12628 3329 -12594
rect 1076 -12779 1082 -12745
rect 1116 -12779 1126 -12745
rect 889 -12823 923 -12789
rect 683 -12934 701 -12900
rect 735 -12934 753 -12900
rect 683 -12968 753 -12934
rect 683 -13002 701 -12968
rect 735 -13002 753 -12968
rect 683 -13017 753 -13002
rect 805 -12857 923 -12823
rect 805 -12899 855 -12857
rect 1076 -12862 1126 -12779
rect 1252 -12763 1272 -12729
rect 1306 -12763 1402 -12729
rect 839 -12933 855 -12899
rect 805 -12967 855 -12933
rect 839 -13001 855 -12967
rect 805 -13017 855 -13001
rect 945 -12900 1011 -12891
rect 945 -12934 961 -12900
rect 995 -12934 1011 -12900
rect 945 -12968 1011 -12934
rect 945 -13002 961 -12968
rect 995 -13002 1011 -12968
rect 945 -13051 1011 -13002
rect 1045 -12899 1126 -12862
rect 1045 -12933 1059 -12899
rect 1093 -12933 1126 -12899
rect 1045 -12967 1126 -12933
rect 1045 -13001 1059 -12967
rect 1093 -13001 1126 -12967
rect 1045 -13017 1126 -13001
rect 1160 -12853 1218 -12818
rect 1160 -12887 1172 -12853
rect 1206 -12887 1218 -12853
rect 1160 -12946 1218 -12887
rect 1160 -12980 1172 -12946
rect 1206 -12980 1218 -12946
rect 1160 -13051 1218 -12980
rect 1252 -12833 1402 -12763
rect 1436 -12765 1586 -12695
rect 1436 -12799 1532 -12765
rect 1566 -12799 1586 -12765
rect 1712 -12763 1790 -12729
rect 1824 -12763 1893 -12729
rect 1927 -12763 1996 -12729
rect 2030 -12763 2050 -12729
rect 1252 -12873 1586 -12833
rect 1252 -12907 1270 -12873
rect 1304 -12907 1534 -12873
rect 1568 -12907 1586 -12873
rect 1252 -12975 1586 -12907
rect 1252 -13009 1270 -12975
rect 1304 -13009 1534 -12975
rect 1568 -13009 1586 -12975
rect 1252 -13051 1586 -13009
rect 1620 -12853 1678 -12818
rect 1620 -12887 1632 -12853
rect 1666 -12887 1678 -12853
rect 1620 -12946 1678 -12887
rect 1620 -12980 1632 -12946
rect 1666 -12980 1678 -12946
rect 1620 -13051 1678 -12980
rect 1712 -12833 2050 -12763
rect 2084 -12765 2414 -12695
rect 2084 -12799 2104 -12765
rect 2138 -12799 2203 -12765
rect 2237 -12799 2302 -12765
rect 2336 -12799 2414 -12765
rect 2540 -12763 2560 -12729
rect 2594 -12763 2690 -12729
rect 1712 -12873 2414 -12833
rect 1712 -12907 1730 -12873
rect 1764 -12907 2362 -12873
rect 2396 -12907 2414 -12873
rect 1712 -12975 2414 -12907
rect 1712 -13009 1730 -12975
rect 1764 -13009 2362 -12975
rect 2396 -13009 2414 -12975
rect 1712 -13051 2414 -13009
rect 2448 -12853 2506 -12818
rect 2448 -12887 2460 -12853
rect 2494 -12887 2506 -12853
rect 2448 -12946 2506 -12887
rect 2448 -12980 2460 -12946
rect 2494 -12980 2506 -12946
rect 2448 -13051 2506 -12980
rect 2540 -12833 2690 -12763
rect 2724 -12765 2874 -12695
rect 3000 -12705 3194 -12671
rect 3124 -12729 3194 -12705
rect 3124 -12739 3210 -12729
rect 2724 -12799 2820 -12765
rect 2854 -12799 2874 -12765
rect 3000 -12773 3040 -12739
rect 3074 -12745 3090 -12739
rect 3000 -12779 3042 -12773
rect 3076 -12779 3090 -12745
rect 3000 -12782 3090 -12779
rect 3124 -12773 3160 -12739
rect 3194 -12773 3210 -12739
rect 3124 -12787 3210 -12773
rect 3259 -12738 3329 -12628
rect 3381 -12594 3431 -12575
rect 3415 -12628 3431 -12594
rect 3381 -12670 3431 -12628
rect 3521 -12594 3587 -12541
rect 3521 -12628 3537 -12594
rect 3571 -12628 3587 -12594
rect 3521 -12644 3587 -12628
rect 3621 -12594 3702 -12575
rect 3621 -12628 3635 -12594
rect 3669 -12628 3702 -12594
rect 3621 -12652 3702 -12628
rect 3381 -12704 3499 -12670
rect 3465 -12723 3499 -12704
rect 3259 -12739 3431 -12738
rect 3259 -12773 3381 -12739
rect 3415 -12773 3431 -12739
rect 3124 -12816 3194 -12787
rect 2540 -12873 2874 -12833
rect 2540 -12907 2558 -12873
rect 2592 -12907 2822 -12873
rect 2856 -12907 2874 -12873
rect 2540 -12975 2874 -12907
rect 2540 -13009 2558 -12975
rect 2592 -13009 2822 -12975
rect 2856 -13009 2874 -12975
rect 2540 -13051 2874 -13009
rect 2908 -12853 2966 -12818
rect 2908 -12887 2920 -12853
rect 2954 -12887 2966 -12853
rect 2908 -12946 2966 -12887
rect 2908 -12980 2920 -12946
rect 2954 -12980 2966 -12946
rect 2908 -13051 2966 -12980
rect 3000 -12850 3194 -12816
rect 3259 -12788 3431 -12773
rect 3465 -12739 3618 -12723
rect 3465 -12773 3581 -12739
rect 3615 -12773 3618 -12739
rect 3000 -12900 3069 -12850
rect 3000 -12934 3019 -12900
rect 3053 -12934 3069 -12900
rect 3000 -12968 3069 -12934
rect 3000 -13002 3019 -12968
rect 3053 -13002 3069 -12968
rect 3000 -13017 3069 -13002
rect 3103 -12900 3169 -12884
rect 3103 -12934 3119 -12900
rect 3153 -12934 3169 -12900
rect 3103 -12968 3169 -12934
rect 3103 -13002 3119 -12968
rect 3153 -13002 3169 -12968
rect 3103 -13051 3169 -13002
rect 3259 -12900 3329 -12788
rect 3465 -12789 3618 -12773
rect 3652 -12745 3702 -12652
rect 3736 -12635 3794 -12541
rect 3736 -12669 3748 -12635
rect 3782 -12669 3794 -12635
rect 3736 -12686 3794 -12669
rect 3828 -12609 4162 -12541
rect 3828 -12643 3846 -12609
rect 3880 -12643 4110 -12609
rect 4144 -12643 4162 -12609
rect 3828 -12695 4162 -12643
rect 4196 -12635 4254 -12541
rect 4196 -12669 4208 -12635
rect 4242 -12669 4254 -12635
rect 4196 -12686 4254 -12669
rect 4288 -12602 4990 -12541
rect 4288 -12636 4306 -12602
rect 4340 -12636 4938 -12602
rect 4972 -12636 4990 -12602
rect 4288 -12695 4990 -12636
rect 5024 -12635 5082 -12541
rect 5024 -12669 5036 -12635
rect 5070 -12669 5082 -12635
rect 5024 -12686 5082 -12669
rect 5116 -12609 5450 -12541
rect 5116 -12643 5134 -12609
rect 5168 -12643 5398 -12609
rect 5432 -12643 5450 -12609
rect 5116 -12695 5450 -12643
rect 5484 -12635 5542 -12541
rect 5484 -12669 5496 -12635
rect 5530 -12669 5542 -12635
rect 5484 -12686 5542 -12669
rect 5576 -12594 5642 -12575
rect 5576 -12628 5595 -12594
rect 5629 -12628 5642 -12594
rect 5576 -12671 5642 -12628
rect 5676 -12594 5742 -12541
rect 5676 -12628 5692 -12594
rect 5726 -12628 5742 -12594
rect 5676 -12637 5742 -12628
rect 5835 -12594 5905 -12575
rect 5835 -12628 5852 -12594
rect 5886 -12628 5905 -12594
rect 3652 -12779 3656 -12745
rect 3690 -12779 3702 -12745
rect 3465 -12823 3499 -12789
rect 3259 -12934 3277 -12900
rect 3311 -12934 3329 -12900
rect 3259 -12968 3329 -12934
rect 3259 -13002 3277 -12968
rect 3311 -13002 3329 -12968
rect 3259 -13017 3329 -13002
rect 3381 -12857 3499 -12823
rect 3381 -12899 3431 -12857
rect 3652 -12862 3702 -12779
rect 3828 -12763 3848 -12729
rect 3882 -12763 3978 -12729
rect 3415 -12933 3431 -12899
rect 3381 -12967 3431 -12933
rect 3415 -13001 3431 -12967
rect 3381 -13017 3431 -13001
rect 3521 -12900 3587 -12891
rect 3521 -12934 3537 -12900
rect 3571 -12934 3587 -12900
rect 3521 -12968 3587 -12934
rect 3521 -13002 3537 -12968
rect 3571 -13002 3587 -12968
rect 3521 -13051 3587 -13002
rect 3621 -12899 3702 -12862
rect 3621 -12933 3635 -12899
rect 3669 -12933 3702 -12899
rect 3621 -12967 3702 -12933
rect 3621 -13001 3635 -12967
rect 3669 -13001 3702 -12967
rect 3621 -13017 3702 -13001
rect 3736 -12853 3794 -12818
rect 3736 -12887 3748 -12853
rect 3782 -12887 3794 -12853
rect 3736 -12946 3794 -12887
rect 3736 -12980 3748 -12946
rect 3782 -12980 3794 -12946
rect 3736 -13051 3794 -12980
rect 3828 -12833 3978 -12763
rect 4012 -12765 4162 -12695
rect 4012 -12799 4108 -12765
rect 4142 -12799 4162 -12765
rect 4288 -12763 4366 -12729
rect 4400 -12763 4469 -12729
rect 4503 -12763 4572 -12729
rect 4606 -12763 4626 -12729
rect 3828 -12873 4162 -12833
rect 3828 -12907 3846 -12873
rect 3880 -12907 4110 -12873
rect 4144 -12907 4162 -12873
rect 3828 -12975 4162 -12907
rect 3828 -13009 3846 -12975
rect 3880 -13009 4110 -12975
rect 4144 -13009 4162 -12975
rect 3828 -13051 4162 -13009
rect 4196 -12853 4254 -12818
rect 4196 -12887 4208 -12853
rect 4242 -12887 4254 -12853
rect 4196 -12946 4254 -12887
rect 4196 -12980 4208 -12946
rect 4242 -12980 4254 -12946
rect 4196 -13051 4254 -12980
rect 4288 -12833 4626 -12763
rect 4660 -12765 4990 -12695
rect 4660 -12799 4680 -12765
rect 4714 -12799 4779 -12765
rect 4813 -12799 4878 -12765
rect 4912 -12799 4990 -12765
rect 5116 -12763 5136 -12729
rect 5170 -12763 5266 -12729
rect 4288 -12873 4990 -12833
rect 4288 -12907 4306 -12873
rect 4340 -12907 4938 -12873
rect 4972 -12907 4990 -12873
rect 4288 -12975 4990 -12907
rect 4288 -13009 4306 -12975
rect 4340 -13009 4938 -12975
rect 4972 -13009 4990 -12975
rect 4288 -13051 4990 -13009
rect 5024 -12853 5082 -12818
rect 5024 -12887 5036 -12853
rect 5070 -12887 5082 -12853
rect 5024 -12946 5082 -12887
rect 5024 -12980 5036 -12946
rect 5070 -12980 5082 -12946
rect 5024 -13051 5082 -12980
rect 5116 -12833 5266 -12763
rect 5300 -12765 5450 -12695
rect 5576 -12705 5770 -12671
rect 5700 -12729 5770 -12705
rect 5700 -12739 5786 -12729
rect 5300 -12799 5396 -12765
rect 5430 -12799 5450 -12765
rect 5576 -12779 5616 -12739
rect 5650 -12779 5666 -12739
rect 5576 -12782 5666 -12779
rect 5700 -12773 5736 -12739
rect 5770 -12773 5786 -12739
rect 5700 -12787 5786 -12773
rect 5835 -12738 5905 -12628
rect 5957 -12594 6007 -12575
rect 5991 -12628 6007 -12594
rect 5957 -12670 6007 -12628
rect 6097 -12594 6163 -12541
rect 6097 -12628 6113 -12594
rect 6147 -12628 6163 -12594
rect 6097 -12644 6163 -12628
rect 6197 -12594 6278 -12575
rect 6197 -12628 6211 -12594
rect 6245 -12628 6278 -12594
rect 6197 -12652 6278 -12628
rect 5957 -12704 6075 -12670
rect 6041 -12723 6075 -12704
rect 5835 -12739 6007 -12738
rect 5835 -12773 5957 -12739
rect 5991 -12773 6007 -12739
rect 5700 -12816 5770 -12787
rect 5116 -12873 5450 -12833
rect 5116 -12907 5134 -12873
rect 5168 -12907 5398 -12873
rect 5432 -12907 5450 -12873
rect 5116 -12975 5450 -12907
rect 5116 -13009 5134 -12975
rect 5168 -13009 5398 -12975
rect 5432 -13009 5450 -12975
rect 5116 -13051 5450 -13009
rect 5484 -12853 5542 -12818
rect 5484 -12887 5496 -12853
rect 5530 -12887 5542 -12853
rect 5484 -12946 5542 -12887
rect 5484 -12980 5496 -12946
rect 5530 -12980 5542 -12946
rect 5484 -13051 5542 -12980
rect 5576 -12850 5770 -12816
rect 5835 -12788 6007 -12773
rect 6041 -12739 6194 -12723
rect 6041 -12773 6157 -12739
rect 6191 -12773 6194 -12739
rect 5576 -12900 5645 -12850
rect 5576 -12934 5595 -12900
rect 5629 -12934 5645 -12900
rect 5576 -12968 5645 -12934
rect 5576 -13002 5595 -12968
rect 5629 -13002 5645 -12968
rect 5576 -13017 5645 -13002
rect 5679 -12900 5745 -12884
rect 5679 -12934 5695 -12900
rect 5729 -12934 5745 -12900
rect 5679 -12968 5745 -12934
rect 5679 -13002 5695 -12968
rect 5729 -13002 5745 -12968
rect 5679 -13051 5745 -13002
rect 5835 -12900 5905 -12788
rect 6041 -12789 6194 -12773
rect 6228 -12745 6278 -12652
rect 6312 -12635 6370 -12541
rect 6312 -12669 6324 -12635
rect 6358 -12669 6370 -12635
rect 6312 -12686 6370 -12669
rect 6404 -12609 6738 -12541
rect 6404 -12643 6422 -12609
rect 6456 -12643 6686 -12609
rect 6720 -12643 6738 -12609
rect 6404 -12695 6738 -12643
rect 6772 -12635 6830 -12541
rect 6772 -12669 6784 -12635
rect 6818 -12669 6830 -12635
rect 6772 -12686 6830 -12669
rect 6864 -12602 7566 -12541
rect 6864 -12636 6882 -12602
rect 6916 -12636 7514 -12602
rect 7548 -12636 7566 -12602
rect 6864 -12695 7566 -12636
rect 7600 -12635 7658 -12541
rect 7600 -12669 7612 -12635
rect 7646 -12669 7658 -12635
rect 7600 -12686 7658 -12669
rect 7692 -12609 8026 -12541
rect 7692 -12643 7710 -12609
rect 7744 -12643 7974 -12609
rect 8008 -12643 8026 -12609
rect 7692 -12695 8026 -12643
rect 8060 -12635 8118 -12541
rect 8060 -12669 8072 -12635
rect 8106 -12669 8118 -12635
rect 8060 -12686 8118 -12669
rect 8152 -12594 8218 -12575
rect 8152 -12628 8171 -12594
rect 8205 -12628 8218 -12594
rect 8152 -12671 8218 -12628
rect 8252 -12594 8318 -12541
rect 8252 -12628 8268 -12594
rect 8302 -12628 8318 -12594
rect 8252 -12637 8318 -12628
rect 8411 -12594 8481 -12575
rect 8411 -12628 8428 -12594
rect 8462 -12628 8481 -12594
rect 6228 -12779 6230 -12745
rect 6264 -12779 6278 -12745
rect 6041 -12823 6075 -12789
rect 5835 -12934 5853 -12900
rect 5887 -12934 5905 -12900
rect 5835 -12968 5905 -12934
rect 5835 -13002 5853 -12968
rect 5887 -13002 5905 -12968
rect 5835 -13017 5905 -13002
rect 5957 -12857 6075 -12823
rect 5957 -12899 6007 -12857
rect 6228 -12862 6278 -12779
rect 6404 -12763 6424 -12729
rect 6458 -12763 6554 -12729
rect 5991 -12933 6007 -12899
rect 5957 -12967 6007 -12933
rect 5991 -13001 6007 -12967
rect 5957 -13017 6007 -13001
rect 6097 -12900 6163 -12891
rect 6097 -12934 6113 -12900
rect 6147 -12934 6163 -12900
rect 6097 -12968 6163 -12934
rect 6097 -13002 6113 -12968
rect 6147 -13002 6163 -12968
rect 6097 -13051 6163 -13002
rect 6197 -12899 6278 -12862
rect 6197 -12933 6211 -12899
rect 6245 -12933 6278 -12899
rect 6197 -12967 6278 -12933
rect 6197 -13001 6211 -12967
rect 6245 -13001 6278 -12967
rect 6197 -13017 6278 -13001
rect 6312 -12853 6370 -12818
rect 6312 -12887 6324 -12853
rect 6358 -12887 6370 -12853
rect 6312 -12946 6370 -12887
rect 6312 -12980 6324 -12946
rect 6358 -12980 6370 -12946
rect 6312 -13051 6370 -12980
rect 6404 -12833 6554 -12763
rect 6588 -12765 6738 -12695
rect 6588 -12799 6684 -12765
rect 6718 -12799 6738 -12765
rect 6864 -12763 6942 -12729
rect 6976 -12763 7045 -12729
rect 7079 -12763 7148 -12729
rect 7182 -12763 7202 -12729
rect 6404 -12873 6738 -12833
rect 6404 -12907 6422 -12873
rect 6456 -12907 6686 -12873
rect 6720 -12907 6738 -12873
rect 6404 -12975 6738 -12907
rect 6404 -13009 6422 -12975
rect 6456 -13009 6686 -12975
rect 6720 -13009 6738 -12975
rect 6404 -13051 6738 -13009
rect 6772 -12853 6830 -12818
rect 6772 -12887 6784 -12853
rect 6818 -12887 6830 -12853
rect 6772 -12946 6830 -12887
rect 6772 -12980 6784 -12946
rect 6818 -12980 6830 -12946
rect 6772 -13051 6830 -12980
rect 6864 -12833 7202 -12763
rect 7236 -12765 7566 -12695
rect 7236 -12799 7256 -12765
rect 7290 -12799 7355 -12765
rect 7389 -12799 7454 -12765
rect 7488 -12799 7566 -12765
rect 7692 -12763 7712 -12729
rect 7746 -12763 7842 -12729
rect 6864 -12873 7566 -12833
rect 6864 -12907 6882 -12873
rect 6916 -12907 7514 -12873
rect 7548 -12907 7566 -12873
rect 6864 -12975 7566 -12907
rect 6864 -13009 6882 -12975
rect 6916 -13009 7514 -12975
rect 7548 -13009 7566 -12975
rect 6864 -13051 7566 -13009
rect 7600 -12853 7658 -12818
rect 7600 -12887 7612 -12853
rect 7646 -12887 7658 -12853
rect 7600 -12946 7658 -12887
rect 7600 -12980 7612 -12946
rect 7646 -12980 7658 -12946
rect 7600 -13051 7658 -12980
rect 7692 -12833 7842 -12763
rect 7876 -12765 8026 -12695
rect 8152 -12705 8346 -12671
rect 8276 -12729 8346 -12705
rect 8276 -12739 8362 -12729
rect 7876 -12799 7972 -12765
rect 8006 -12799 8026 -12765
rect 8152 -12745 8192 -12739
rect 8152 -12779 8190 -12745
rect 8226 -12773 8242 -12739
rect 8224 -12779 8242 -12773
rect 8152 -12782 8242 -12779
rect 8276 -12773 8312 -12739
rect 8346 -12773 8362 -12739
rect 8276 -12787 8362 -12773
rect 8411 -12738 8481 -12628
rect 8533 -12594 8583 -12575
rect 8567 -12628 8583 -12594
rect 8533 -12670 8583 -12628
rect 8673 -12594 8739 -12541
rect 8673 -12628 8689 -12594
rect 8723 -12628 8739 -12594
rect 8673 -12644 8739 -12628
rect 8773 -12594 8854 -12575
rect 8773 -12628 8787 -12594
rect 8821 -12628 8854 -12594
rect 8773 -12652 8854 -12628
rect 8533 -12704 8651 -12670
rect 8617 -12723 8651 -12704
rect 8411 -12739 8583 -12738
rect 8411 -12773 8533 -12739
rect 8567 -12773 8583 -12739
rect 8276 -12816 8346 -12787
rect 7692 -12873 8026 -12833
rect 7692 -12907 7710 -12873
rect 7744 -12907 7974 -12873
rect 8008 -12907 8026 -12873
rect 7692 -12975 8026 -12907
rect 7692 -13009 7710 -12975
rect 7744 -13009 7974 -12975
rect 8008 -13009 8026 -12975
rect 7692 -13051 8026 -13009
rect 8060 -12853 8118 -12818
rect 8060 -12887 8072 -12853
rect 8106 -12887 8118 -12853
rect 8060 -12946 8118 -12887
rect 8060 -12980 8072 -12946
rect 8106 -12980 8118 -12946
rect 8060 -13051 8118 -12980
rect 8152 -12850 8346 -12816
rect 8411 -12788 8583 -12773
rect 8617 -12739 8770 -12723
rect 8617 -12773 8733 -12739
rect 8767 -12773 8770 -12739
rect 8152 -12900 8221 -12850
rect 8152 -12934 8171 -12900
rect 8205 -12934 8221 -12900
rect 8152 -12968 8221 -12934
rect 8152 -13002 8171 -12968
rect 8205 -13002 8221 -12968
rect 8152 -13017 8221 -13002
rect 8255 -12900 8321 -12884
rect 8255 -12934 8271 -12900
rect 8305 -12934 8321 -12900
rect 8255 -12968 8321 -12934
rect 8255 -13002 8271 -12968
rect 8305 -13002 8321 -12968
rect 8255 -13051 8321 -13002
rect 8411 -12900 8481 -12788
rect 8617 -12789 8770 -12773
rect 8804 -12745 8854 -12652
rect 8888 -12635 8946 -12541
rect 8888 -12669 8900 -12635
rect 8934 -12669 8946 -12635
rect 8888 -12686 8946 -12669
rect 8980 -12609 9314 -12541
rect 8980 -12643 8998 -12609
rect 9032 -12643 9262 -12609
rect 9296 -12643 9314 -12609
rect 8980 -12695 9314 -12643
rect 9348 -12635 9406 -12541
rect 9348 -12669 9360 -12635
rect 9394 -12669 9406 -12635
rect 9348 -12686 9406 -12669
rect 9440 -12602 10142 -12541
rect 9440 -12636 9458 -12602
rect 9492 -12636 10090 -12602
rect 10124 -12636 10142 -12602
rect 9440 -12695 10142 -12636
rect 10176 -12635 10234 -12541
rect 10176 -12669 10188 -12635
rect 10222 -12669 10234 -12635
rect 10176 -12686 10234 -12669
rect 10360 -12609 10694 -12541
rect 10360 -12643 10378 -12609
rect 10412 -12643 10642 -12609
rect 10676 -12643 10694 -12609
rect 10360 -12695 10694 -12643
rect 8838 -12779 8854 -12745
rect 8617 -12823 8651 -12789
rect 8411 -12934 8429 -12900
rect 8463 -12934 8481 -12900
rect 8411 -12968 8481 -12934
rect 8411 -13002 8429 -12968
rect 8463 -13002 8481 -12968
rect 8411 -13017 8481 -13002
rect 8533 -12857 8651 -12823
rect 8533 -12899 8583 -12857
rect 8804 -12862 8854 -12779
rect 8980 -12763 9000 -12729
rect 9034 -12763 9130 -12729
rect 8567 -12933 8583 -12899
rect 8533 -12967 8583 -12933
rect 8567 -13001 8583 -12967
rect 8533 -13017 8583 -13001
rect 8673 -12900 8739 -12891
rect 8673 -12934 8689 -12900
rect 8723 -12934 8739 -12900
rect 8673 -12968 8739 -12934
rect 8673 -13002 8689 -12968
rect 8723 -13002 8739 -12968
rect 8673 -13051 8739 -13002
rect 8773 -12899 8854 -12862
rect 8773 -12933 8787 -12899
rect 8821 -12933 8854 -12899
rect 8773 -12967 8854 -12933
rect 8773 -13001 8787 -12967
rect 8821 -13001 8854 -12967
rect 8773 -13017 8854 -13001
rect 8888 -12853 8946 -12818
rect 8888 -12887 8900 -12853
rect 8934 -12887 8946 -12853
rect 8888 -12946 8946 -12887
rect 8888 -12980 8900 -12946
rect 8934 -12980 8946 -12946
rect 8888 -13051 8946 -12980
rect 8980 -12833 9130 -12763
rect 9164 -12765 9314 -12695
rect 9164 -12799 9260 -12765
rect 9294 -12799 9314 -12765
rect 9440 -12763 9518 -12729
rect 9552 -12763 9621 -12729
rect 9655 -12763 9724 -12729
rect 9758 -12763 9778 -12729
rect 8980 -12873 9314 -12833
rect 8980 -12907 8998 -12873
rect 9032 -12907 9262 -12873
rect 9296 -12907 9314 -12873
rect 8980 -12975 9314 -12907
rect 8980 -13009 8998 -12975
rect 9032 -13009 9262 -12975
rect 9296 -13009 9314 -12975
rect 8980 -13051 9314 -13009
rect 9348 -12853 9406 -12818
rect 9348 -12887 9360 -12853
rect 9394 -12887 9406 -12853
rect 9348 -12946 9406 -12887
rect 9348 -12980 9360 -12946
rect 9394 -12980 9406 -12946
rect 9348 -13051 9406 -12980
rect 9440 -12833 9778 -12763
rect 9812 -12765 10142 -12695
rect 9812 -12799 9832 -12765
rect 9866 -12799 9931 -12765
rect 9965 -12799 10030 -12765
rect 10064 -12799 10142 -12765
rect 10360 -12763 10380 -12729
rect 10414 -12763 10510 -12729
rect 9440 -12873 10142 -12833
rect 9440 -12907 9458 -12873
rect 9492 -12907 10090 -12873
rect 10124 -12907 10142 -12873
rect 9440 -12975 10142 -12907
rect 9440 -13009 9458 -12975
rect 9492 -13009 10090 -12975
rect 10124 -13009 10142 -12975
rect 9440 -13051 10142 -13009
rect 10176 -12853 10234 -12818
rect 10176 -12887 10188 -12853
rect 10222 -12887 10234 -12853
rect 10176 -12946 10234 -12887
rect 10176 -12980 10188 -12946
rect 10222 -12980 10234 -12946
rect 10176 -13051 10234 -12980
rect 10360 -12833 10510 -12763
rect 10544 -12765 10694 -12695
rect 10728 -12594 10794 -12575
rect 10728 -12628 10747 -12594
rect 10781 -12628 10794 -12594
rect 10728 -12671 10794 -12628
rect 10828 -12594 10894 -12541
rect 10828 -12628 10844 -12594
rect 10878 -12628 10894 -12594
rect 10828 -12637 10894 -12628
rect 10987 -12594 11057 -12575
rect 10987 -12628 11004 -12594
rect 11038 -12628 11057 -12594
rect 10728 -12705 10922 -12671
rect 10852 -12729 10922 -12705
rect 10852 -12739 10938 -12729
rect 10544 -12799 10640 -12765
rect 10674 -12799 10694 -12765
rect 10728 -12745 10768 -12739
rect 10728 -12779 10764 -12745
rect 10802 -12773 10818 -12739
rect 10798 -12779 10818 -12773
rect 10728 -12782 10818 -12779
rect 10852 -12773 10888 -12739
rect 10922 -12773 10938 -12739
rect 10852 -12787 10938 -12773
rect 10987 -12738 11057 -12628
rect 11109 -12594 11159 -12575
rect 11143 -12628 11159 -12594
rect 11109 -12670 11159 -12628
rect 11249 -12594 11315 -12541
rect 11249 -12628 11265 -12594
rect 11299 -12628 11315 -12594
rect 11249 -12644 11315 -12628
rect 11349 -12594 11430 -12575
rect 11349 -12628 11363 -12594
rect 11397 -12628 11430 -12594
rect 11349 -12652 11430 -12628
rect 11109 -12704 11227 -12670
rect 11193 -12723 11227 -12704
rect 10987 -12739 11159 -12738
rect 10987 -12773 11109 -12739
rect 11143 -12773 11159 -12739
rect 10852 -12816 10922 -12787
rect 10360 -12873 10694 -12833
rect 10360 -12907 10378 -12873
rect 10412 -12907 10642 -12873
rect 10676 -12907 10694 -12873
rect 10360 -12975 10694 -12907
rect 10360 -13009 10378 -12975
rect 10412 -13009 10642 -12975
rect 10676 -13009 10694 -12975
rect 10360 -13051 10694 -13009
rect 10728 -12850 10922 -12816
rect 10987 -12788 11159 -12773
rect 11193 -12739 11346 -12723
rect 11193 -12773 11309 -12739
rect 11343 -12773 11346 -12739
rect 10728 -12900 10797 -12850
rect 10728 -12934 10747 -12900
rect 10781 -12934 10797 -12900
rect 10728 -12968 10797 -12934
rect 10728 -13002 10747 -12968
rect 10781 -13002 10797 -12968
rect 10728 -13017 10797 -13002
rect 10831 -12900 10897 -12884
rect 10831 -12934 10847 -12900
rect 10881 -12934 10897 -12900
rect 10831 -12968 10897 -12934
rect 10831 -13002 10847 -12968
rect 10881 -13002 10897 -12968
rect 10831 -13051 10897 -13002
rect 10987 -12900 11057 -12788
rect 11193 -12789 11346 -12773
rect 11380 -12778 11430 -12652
rect 11464 -12635 11522 -12541
rect 11464 -12669 11476 -12635
rect 11510 -12669 11522 -12635
rect 11464 -12686 11522 -12669
rect 11648 -12609 11982 -12541
rect 11648 -12643 11666 -12609
rect 11700 -12643 11930 -12609
rect 11964 -12643 11982 -12609
rect 11648 -12695 11982 -12643
rect 12384 -12635 12442 -12541
rect 12572 -12585 12631 -12541
rect 12572 -12619 12588 -12585
rect 12622 -12619 12631 -12585
rect 12572 -12635 12631 -12619
rect 12665 -12596 12717 -12580
rect 12665 -12630 12674 -12596
rect 12708 -12630 12717 -12596
rect 12384 -12669 12396 -12635
rect 12430 -12669 12442 -12635
rect 12665 -12669 12717 -12630
rect 12751 -12585 12803 -12541
rect 12751 -12619 12760 -12585
rect 12794 -12619 12803 -12585
rect 12751 -12635 12803 -12619
rect 12837 -12596 12888 -12580
rect 12837 -12630 12846 -12596
rect 12880 -12630 12888 -12596
rect 12837 -12669 12888 -12630
rect 12922 -12585 12982 -12541
rect 12922 -12619 12932 -12585
rect 12966 -12619 12982 -12585
rect 12922 -12635 12982 -12619
rect 13120 -12635 13178 -12541
rect 13120 -12669 13132 -12635
rect 13166 -12669 13178 -12635
rect 12384 -12686 12442 -12669
rect 12480 -12677 13086 -12669
rect 11193 -12823 11227 -12789
rect 10987 -12934 11005 -12900
rect 11039 -12934 11057 -12900
rect 10987 -12968 11057 -12934
rect 10987 -13002 11005 -12968
rect 11039 -13002 11057 -12968
rect 10987 -13017 11057 -13002
rect 11109 -12857 11227 -12823
rect 11380 -12812 11389 -12778
rect 11423 -12812 11430 -12778
rect 11109 -12899 11159 -12857
rect 11380 -12862 11430 -12812
rect 11648 -12763 11668 -12729
rect 11702 -12763 11798 -12729
rect 11143 -12933 11159 -12899
rect 11109 -12967 11159 -12933
rect 11143 -13001 11159 -12967
rect 11109 -13017 11159 -13001
rect 11249 -12900 11315 -12891
rect 11249 -12934 11265 -12900
rect 11299 -12934 11315 -12900
rect 11249 -12968 11315 -12934
rect 11249 -13002 11265 -12968
rect 11299 -13002 11315 -12968
rect 11249 -13051 11315 -13002
rect 11349 -12899 11430 -12862
rect 11349 -12933 11363 -12899
rect 11397 -12933 11430 -12899
rect 11349 -12967 11430 -12933
rect 11349 -13001 11363 -12967
rect 11397 -13001 11430 -12967
rect 11349 -13017 11430 -13001
rect 11464 -12853 11522 -12818
rect 11464 -12887 11476 -12853
rect 11510 -12887 11522 -12853
rect 11464 -12946 11522 -12887
rect 11464 -12980 11476 -12946
rect 11510 -12980 11522 -12946
rect 11464 -13051 11522 -12980
rect 11648 -12833 11798 -12763
rect 11832 -12765 11982 -12695
rect 11832 -12799 11928 -12765
rect 11962 -12799 11982 -12765
rect 12480 -12703 13038 -12677
rect 12480 -12816 12514 -12703
rect 13026 -12711 13038 -12703
rect 13072 -12711 13086 -12677
rect 13120 -12686 13178 -12669
rect 13212 -12609 13546 -12541
rect 13212 -12643 13230 -12609
rect 13264 -12643 13494 -12609
rect 13528 -12643 13546 -12609
rect 12548 -12739 12991 -12737
rect 12548 -12742 12574 -12739
rect 12548 -12776 12558 -12742
rect 12608 -12773 12642 -12739
rect 12676 -12773 12710 -12739
rect 12744 -12742 12778 -12739
rect 12773 -12773 12778 -12742
rect 12812 -12742 12846 -12739
rect 12812 -12773 12836 -12742
rect 12880 -12773 12914 -12739
rect 12948 -12742 12991 -12739
rect 12592 -12776 12642 -12773
rect 12676 -12776 12739 -12773
rect 12773 -12776 12836 -12773
rect 12870 -12776 12942 -12773
rect 12976 -12776 12991 -12742
rect 12548 -12782 12991 -12776
rect 13026 -12749 13086 -12711
rect 13026 -12783 13038 -12749
rect 13072 -12783 13086 -12749
rect 13026 -12816 13086 -12783
rect 13212 -12695 13546 -12643
rect 13580 -12635 13638 -12541
rect 13580 -12669 13592 -12635
rect 13626 -12669 13638 -12635
rect 13672 -12583 13733 -12541
rect 13672 -12617 13690 -12583
rect 13724 -12617 13733 -12583
rect 13672 -12643 13733 -12617
rect 13769 -12596 13819 -12577
rect 13769 -12630 13776 -12596
rect 13810 -12630 13819 -12596
rect 13580 -12686 13638 -12669
rect 13212 -12765 13362 -12695
rect 13672 -12712 13735 -12677
rect 13212 -12799 13232 -12765
rect 13266 -12799 13362 -12765
rect 13396 -12763 13492 -12729
rect 13526 -12763 13546 -12729
rect 11648 -12873 11982 -12833
rect 11648 -12907 11666 -12873
rect 11700 -12907 11930 -12873
rect 11964 -12907 11982 -12873
rect 11648 -12975 11982 -12907
rect 11648 -13009 11666 -12975
rect 11700 -13009 11930 -12975
rect 11964 -13009 11982 -12975
rect 11648 -13051 11982 -13009
rect 12384 -12853 12442 -12818
rect 12480 -12850 13086 -12816
rect 12384 -12887 12396 -12853
rect 12430 -12887 12442 -12853
rect 12580 -12873 12631 -12850
rect 12384 -12946 12442 -12887
rect 12384 -12980 12396 -12946
rect 12430 -12980 12442 -12946
rect 12384 -13051 12442 -12980
rect 12476 -12900 12545 -12884
rect 12476 -12934 12502 -12900
rect 12536 -12934 12545 -12900
rect 12476 -12968 12545 -12934
rect 12476 -13002 12502 -12968
rect 12536 -13002 12545 -12968
rect 12476 -13051 12545 -13002
rect 12580 -12907 12588 -12873
rect 12622 -12907 12631 -12873
rect 12752 -12873 12803 -12850
rect 12580 -12961 12631 -12907
rect 12580 -12995 12588 -12961
rect 12622 -12995 12631 -12961
rect 12580 -13011 12631 -12995
rect 12665 -12900 12717 -12884
rect 12665 -12934 12674 -12900
rect 12708 -12934 12717 -12900
rect 12665 -12968 12717 -12934
rect 12665 -13002 12674 -12968
rect 12708 -13002 12717 -12968
rect 12665 -13051 12717 -13002
rect 12752 -12907 12760 -12873
rect 12794 -12907 12803 -12873
rect 12923 -12873 12975 -12850
rect 12752 -12961 12803 -12907
rect 12752 -12995 12760 -12961
rect 12794 -12995 12803 -12961
rect 12752 -13011 12803 -12995
rect 12837 -12900 12889 -12884
rect 12837 -12934 12846 -12900
rect 12880 -12934 12889 -12900
rect 12837 -12968 12889 -12934
rect 12837 -13002 12846 -12968
rect 12880 -13002 12889 -12968
rect 12837 -13051 12889 -13002
rect 12923 -12907 12932 -12873
rect 12966 -12907 12975 -12873
rect 13120 -12853 13178 -12818
rect 13396 -12833 13546 -12763
rect 13672 -12746 13684 -12712
rect 13718 -12739 13735 -12712
rect 13672 -12773 13692 -12746
rect 13726 -12773 13735 -12739
rect 13672 -12789 13735 -12773
rect 13769 -12739 13819 -12630
rect 13853 -12596 13905 -12541
rect 13853 -12630 13862 -12596
rect 13896 -12630 13905 -12596
rect 13853 -12646 13905 -12630
rect 13941 -12596 13991 -12577
rect 13941 -12630 13948 -12596
rect 13982 -12630 13991 -12596
rect 13941 -12739 13991 -12630
rect 14025 -12596 14077 -12541
rect 14025 -12630 14034 -12596
rect 14068 -12630 14077 -12596
rect 14025 -12653 14077 -12630
rect 14111 -12596 14163 -12580
rect 14111 -12630 14120 -12596
rect 14154 -12630 14163 -12596
rect 14111 -12671 14163 -12630
rect 14197 -12587 14249 -12541
rect 14197 -12621 14206 -12587
rect 14240 -12621 14249 -12587
rect 14197 -12637 14249 -12621
rect 14283 -12596 14335 -12580
rect 14283 -12630 14292 -12596
rect 14326 -12630 14335 -12596
rect 14283 -12671 14335 -12630
rect 14369 -12587 14421 -12541
rect 14369 -12621 14378 -12587
rect 14412 -12621 14421 -12587
rect 14369 -12637 14421 -12621
rect 14455 -12596 14507 -12580
rect 14455 -12630 14464 -12596
rect 14498 -12630 14507 -12596
rect 14455 -12671 14507 -12630
rect 14541 -12587 14590 -12541
rect 14541 -12621 14550 -12587
rect 14584 -12621 14590 -12587
rect 14541 -12637 14590 -12621
rect 14624 -12596 14679 -12580
rect 14624 -12630 14636 -12596
rect 14670 -12630 14679 -12596
rect 14624 -12671 14679 -12630
rect 14713 -12587 14762 -12541
rect 14713 -12621 14722 -12587
rect 14756 -12621 14762 -12587
rect 14713 -12637 14762 -12621
rect 14796 -12596 14848 -12580
rect 14796 -12630 14807 -12596
rect 14841 -12630 14848 -12596
rect 14796 -12671 14848 -12630
rect 14884 -12587 14934 -12541
rect 14884 -12621 14893 -12587
rect 14927 -12621 14934 -12587
rect 14884 -12637 14934 -12621
rect 14968 -12596 15020 -12580
rect 14968 -12630 14979 -12596
rect 15013 -12630 15020 -12596
rect 14968 -12671 15020 -12630
rect 15056 -12587 15106 -12541
rect 15056 -12621 15065 -12587
rect 15099 -12621 15106 -12587
rect 15056 -12637 15106 -12621
rect 15140 -12596 15192 -12580
rect 15140 -12630 15151 -12596
rect 15185 -12630 15192 -12596
rect 15140 -12671 15192 -12630
rect 15228 -12587 15280 -12541
rect 15228 -12621 15237 -12587
rect 15271 -12621 15280 -12587
rect 15228 -12637 15280 -12621
rect 15314 -12596 15366 -12580
rect 15314 -12630 15323 -12596
rect 15357 -12630 15366 -12596
rect 15314 -12671 15366 -12630
rect 15400 -12587 15460 -12541
rect 15400 -12621 15409 -12587
rect 15443 -12621 15460 -12587
rect 15400 -12637 15460 -12621
rect 15512 -12635 15570 -12541
rect 15512 -12669 15524 -12635
rect 15558 -12669 15570 -12635
rect 14111 -12700 15460 -12671
rect 15512 -12686 15570 -12669
rect 15604 -12602 16673 -12541
rect 15604 -12636 15622 -12602
rect 15656 -12636 16622 -12602
rect 16656 -12636 16673 -12602
rect 14111 -12705 15248 -12700
rect 15227 -12734 15248 -12705
rect 15282 -12734 15341 -12700
rect 15375 -12734 15460 -12700
rect 13769 -12773 14119 -12739
rect 14153 -12773 14187 -12739
rect 14221 -12773 14255 -12739
rect 14289 -12773 14323 -12739
rect 14357 -12773 14391 -12739
rect 14425 -12773 14459 -12739
rect 14493 -12773 14527 -12739
rect 14561 -12773 14595 -12739
rect 14629 -12773 14663 -12739
rect 14697 -12773 14731 -12739
rect 14765 -12773 14799 -12739
rect 14833 -12773 14867 -12739
rect 14901 -12773 14935 -12739
rect 14969 -12773 15003 -12739
rect 15037 -12773 15071 -12739
rect 15105 -12773 15139 -12739
rect 15173 -12773 15193 -12739
rect 13769 -12789 15193 -12773
rect 12923 -12961 12975 -12907
rect 12923 -12995 12932 -12961
rect 12966 -12995 12975 -12961
rect 12923 -13011 12975 -12995
rect 13009 -12900 13086 -12884
rect 13009 -12934 13018 -12900
rect 13052 -12934 13086 -12900
rect 13009 -12968 13086 -12934
rect 13009 -13002 13018 -12968
rect 13052 -13002 13086 -12968
rect 13009 -13051 13086 -13002
rect 13120 -12887 13132 -12853
rect 13166 -12887 13178 -12853
rect 13120 -12946 13178 -12887
rect 13120 -12980 13132 -12946
rect 13166 -12980 13178 -12946
rect 13120 -13051 13178 -12980
rect 13212 -12873 13546 -12833
rect 13212 -12907 13230 -12873
rect 13264 -12907 13494 -12873
rect 13528 -12907 13546 -12873
rect 13212 -12975 13546 -12907
rect 13212 -13009 13230 -12975
rect 13264 -13009 13494 -12975
rect 13528 -13009 13546 -12975
rect 13212 -13051 13546 -13009
rect 13580 -12853 13638 -12818
rect 13580 -12887 13592 -12853
rect 13626 -12887 13638 -12853
rect 13580 -12946 13638 -12887
rect 13580 -12980 13592 -12946
rect 13626 -12980 13638 -12946
rect 13580 -13051 13638 -12980
rect 13674 -12907 13733 -12889
rect 13674 -12941 13690 -12907
rect 13724 -12941 13733 -12907
rect 13674 -12975 13733 -12941
rect 13674 -13009 13690 -12975
rect 13724 -13009 13733 -12975
rect 13674 -13051 13733 -13009
rect 13769 -12899 13818 -12789
rect 13769 -12933 13776 -12899
rect 13810 -12933 13818 -12899
rect 13769 -12967 13818 -12933
rect 13769 -13001 13776 -12967
rect 13810 -13001 13818 -12967
rect 13769 -13017 13818 -13001
rect 13853 -12907 13905 -12889
rect 13853 -12941 13862 -12907
rect 13896 -12941 13905 -12907
rect 13853 -12975 13905 -12941
rect 13853 -13009 13862 -12975
rect 13896 -13009 13905 -12975
rect 13853 -13051 13905 -13009
rect 13941 -12891 13991 -12789
rect 15227 -12795 15460 -12734
rect 15227 -12796 15340 -12795
rect 15227 -12823 15248 -12796
rect 14111 -12830 15248 -12823
rect 15282 -12829 15340 -12796
rect 15374 -12829 15460 -12795
rect 15604 -12695 16673 -12636
rect 15604 -12765 16120 -12695
rect 15604 -12799 15682 -12765
rect 15716 -12799 15810 -12765
rect 15844 -12799 15938 -12765
rect 15972 -12799 16066 -12765
rect 16100 -12799 16120 -12765
rect 16154 -12763 16174 -12729
rect 16208 -12763 16302 -12729
rect 16336 -12763 16430 -12729
rect 16464 -12763 16558 -12729
rect 16592 -12763 16673 -12729
rect 15282 -12830 15460 -12829
rect 14111 -12845 15460 -12830
rect 14111 -12879 14120 -12845
rect 14154 -12871 14292 -12845
rect 14154 -12879 14163 -12871
rect 13941 -12925 13948 -12891
rect 13982 -12925 13991 -12891
rect 13941 -12959 13991 -12925
rect 13941 -12993 13948 -12959
rect 13982 -12993 13991 -12959
rect 13941 -13016 13991 -12993
rect 14025 -12907 14077 -12891
rect 14025 -12941 14034 -12907
rect 14068 -12941 14077 -12907
rect 14025 -12975 14077 -12941
rect 14025 -13009 14034 -12975
rect 14068 -13009 14077 -12975
rect 14025 -13050 14077 -13009
rect 14111 -12931 14163 -12879
rect 14283 -12879 14292 -12871
rect 14326 -12871 14464 -12845
rect 14326 -12879 14335 -12871
rect 14111 -12965 14120 -12931
rect 14154 -12965 14163 -12931
rect 14111 -13016 14163 -12965
rect 14197 -12951 14249 -12905
rect 14197 -12985 14206 -12951
rect 14240 -12985 14249 -12951
rect 14197 -13050 14249 -12985
rect 14283 -12931 14335 -12879
rect 14455 -12879 14464 -12871
rect 14498 -12871 14636 -12845
rect 14498 -12879 14507 -12871
rect 14283 -12965 14292 -12931
rect 14326 -12965 14335 -12931
rect 14283 -13016 14335 -12965
rect 14369 -12951 14421 -12905
rect 14369 -12985 14378 -12951
rect 14412 -12985 14421 -12951
rect 14369 -13050 14421 -12985
rect 14455 -12931 14507 -12879
rect 14627 -12879 14636 -12871
rect 14670 -12871 14807 -12845
rect 14670 -12879 14679 -12871
rect 14455 -12965 14464 -12931
rect 14498 -12965 14507 -12931
rect 14455 -13016 14507 -12965
rect 14541 -12951 14593 -12905
rect 14541 -12985 14550 -12951
rect 14584 -12985 14593 -12951
rect 14541 -13050 14593 -12985
rect 14627 -12931 14679 -12879
rect 14796 -12879 14807 -12871
rect 14841 -12871 14979 -12845
rect 14841 -12879 14848 -12871
rect 14627 -12965 14636 -12931
rect 14670 -12965 14679 -12931
rect 14627 -13016 14679 -12965
rect 14713 -12951 14762 -12905
rect 14713 -12985 14722 -12951
rect 14756 -12985 14762 -12951
rect 14713 -13050 14762 -12985
rect 14796 -12931 14848 -12879
rect 14968 -12879 14979 -12871
rect 15013 -12871 15151 -12845
rect 15013 -12879 15020 -12871
rect 14796 -12965 14807 -12931
rect 14841 -12965 14848 -12931
rect 14796 -13016 14848 -12965
rect 14885 -12951 14934 -12905
rect 14885 -12985 14893 -12951
rect 14927 -12985 14934 -12951
rect 14885 -13050 14934 -12985
rect 14968 -12931 15020 -12879
rect 15140 -12879 15151 -12871
rect 15185 -12868 15323 -12845
rect 15185 -12879 15192 -12868
rect 14968 -12965 14979 -12931
rect 15013 -12965 15020 -12931
rect 14968 -13016 15020 -12965
rect 15057 -12951 15106 -12905
rect 15057 -12985 15065 -12951
rect 15099 -12985 15106 -12951
rect 15057 -13050 15106 -12985
rect 15140 -12931 15192 -12879
rect 15314 -12879 15323 -12868
rect 15357 -12868 15460 -12845
rect 15512 -12853 15570 -12818
rect 16154 -12833 16673 -12763
rect 15357 -12879 15372 -12868
rect 15140 -12965 15151 -12931
rect 15185 -12965 15192 -12931
rect 15140 -13016 15192 -12965
rect 15229 -12951 15280 -12905
rect 15229 -12985 15237 -12951
rect 15271 -12985 15280 -12951
rect 15229 -13050 15280 -12985
rect 15314 -12931 15372 -12879
rect 15512 -12887 15524 -12853
rect 15558 -12887 15570 -12853
rect 15314 -12965 15323 -12931
rect 15357 -12965 15372 -12931
rect 15314 -13016 15372 -12965
rect 15406 -12951 15460 -12902
rect 15406 -12985 15409 -12951
rect 15443 -12985 15460 -12951
rect 14025 -13051 15280 -13050
rect 15406 -13051 15460 -12985
rect 15512 -12946 15570 -12887
rect 15512 -12980 15524 -12946
rect 15558 -12980 15570 -12946
rect 15512 -13051 15570 -12980
rect 15604 -12873 16673 -12833
rect 15604 -12907 15622 -12873
rect 15656 -12907 16622 -12873
rect 16656 -12907 16673 -12873
rect 15604 -12975 16673 -12907
rect 15604 -13009 15622 -12975
rect 15656 -13009 16622 -12975
rect 16656 -13009 16673 -12975
rect 15604 -13051 16673 -13009
rect -2997 -13085 -2968 -13051
rect -2934 -13085 -2876 -13051
rect -2842 -13085 -2784 -13051
rect -2750 -13085 -2692 -13051
rect -2658 -13085 -2600 -13051
rect -2566 -13085 -2508 -13051
rect -2474 -13085 -2416 -13051
rect -2382 -13085 -2324 -13051
rect -2290 -13085 -2232 -13051
rect -2198 -13085 -2140 -13051
rect -2106 -13085 -2048 -13051
rect -2014 -13085 -1956 -13051
rect -1922 -13085 -1864 -13051
rect -1830 -13085 -1772 -13051
rect -1738 -13085 -1680 -13051
rect -1646 -13085 -1588 -13051
rect -1554 -13085 -1496 -13051
rect -1462 -13085 -1404 -13051
rect -1370 -13085 -1312 -13051
rect -1278 -13085 -1220 -13051
rect -1186 -13085 -1128 -13051
rect -1094 -13085 -1036 -13051
rect -1002 -13085 -944 -13051
rect -910 -13085 -852 -13051
rect -818 -13085 -760 -13051
rect -726 -13085 -668 -13051
rect -634 -13085 -576 -13051
rect -542 -13085 -484 -13051
rect -450 -13085 -392 -13051
rect -358 -13085 -300 -13051
rect -266 -13085 -208 -13051
rect -174 -13085 -116 -13051
rect -82 -13085 -24 -13051
rect 10 -13085 68 -13051
rect 102 -13085 160 -13051
rect 194 -13085 252 -13051
rect 286 -13085 344 -13051
rect 378 -13085 436 -13051
rect 470 -13085 528 -13051
rect 562 -13085 620 -13051
rect 654 -13085 712 -13051
rect 746 -13085 804 -13051
rect 838 -13085 896 -13051
rect 930 -13085 988 -13051
rect 1022 -13085 1080 -13051
rect 1114 -13085 1172 -13051
rect 1206 -13085 1264 -13051
rect 1298 -13085 1356 -13051
rect 1390 -13085 1448 -13051
rect 1482 -13085 1540 -13051
rect 1574 -13085 1632 -13051
rect 1666 -13085 1724 -13051
rect 1758 -13085 1816 -13051
rect 1850 -13085 1908 -13051
rect 1942 -13085 2000 -13051
rect 2034 -13085 2092 -13051
rect 2126 -13085 2184 -13051
rect 2218 -13085 2276 -13051
rect 2310 -13085 2368 -13051
rect 2402 -13085 2460 -13051
rect 2494 -13085 2552 -13051
rect 2586 -13085 2644 -13051
rect 2678 -13085 2736 -13051
rect 2770 -13085 2828 -13051
rect 2862 -13085 2920 -13051
rect 2954 -13085 3012 -13051
rect 3046 -13085 3104 -13051
rect 3138 -13085 3196 -13051
rect 3230 -13085 3288 -13051
rect 3322 -13085 3380 -13051
rect 3414 -13085 3472 -13051
rect 3506 -13085 3564 -13051
rect 3598 -13085 3656 -13051
rect 3690 -13085 3748 -13051
rect 3782 -13085 3840 -13051
rect 3874 -13085 3932 -13051
rect 3966 -13085 4024 -13051
rect 4058 -13085 4116 -13051
rect 4150 -13085 4208 -13051
rect 4242 -13085 4300 -13051
rect 4334 -13085 4392 -13051
rect 4426 -13085 4484 -13051
rect 4518 -13085 4576 -13051
rect 4610 -13085 4668 -13051
rect 4702 -13085 4760 -13051
rect 4794 -13085 4852 -13051
rect 4886 -13085 4944 -13051
rect 4978 -13085 5036 -13051
rect 5070 -13085 5128 -13051
rect 5162 -13085 5220 -13051
rect 5254 -13085 5312 -13051
rect 5346 -13085 5404 -13051
rect 5438 -13085 5496 -13051
rect 5530 -13085 5588 -13051
rect 5622 -13085 5680 -13051
rect 5714 -13085 5772 -13051
rect 5806 -13085 5864 -13051
rect 5898 -13085 5956 -13051
rect 5990 -13085 6048 -13051
rect 6082 -13085 6140 -13051
rect 6174 -13085 6232 -13051
rect 6266 -13085 6324 -13051
rect 6358 -13085 6416 -13051
rect 6450 -13085 6508 -13051
rect 6542 -13085 6600 -13051
rect 6634 -13085 6692 -13051
rect 6726 -13085 6784 -13051
rect 6818 -13085 6876 -13051
rect 6910 -13085 6968 -13051
rect 7002 -13085 7060 -13051
rect 7094 -13085 7152 -13051
rect 7186 -13085 7244 -13051
rect 7278 -13085 7336 -13051
rect 7370 -13085 7428 -13051
rect 7462 -13085 7520 -13051
rect 7554 -13085 7612 -13051
rect 7646 -13085 7704 -13051
rect 7738 -13085 7796 -13051
rect 7830 -13085 7888 -13051
rect 7922 -13085 7980 -13051
rect 8014 -13085 8072 -13051
rect 8106 -13085 8164 -13051
rect 8198 -13085 8256 -13051
rect 8290 -13085 8348 -13051
rect 8382 -13085 8440 -13051
rect 8474 -13085 8532 -13051
rect 8566 -13085 8624 -13051
rect 8658 -13085 8716 -13051
rect 8750 -13085 8808 -13051
rect 8842 -13085 8900 -13051
rect 8934 -13085 8992 -13051
rect 9026 -13085 9084 -13051
rect 9118 -13085 9176 -13051
rect 9210 -13085 9268 -13051
rect 9302 -13085 9360 -13051
rect 9394 -13085 9452 -13051
rect 9486 -13085 9544 -13051
rect 9578 -13085 9636 -13051
rect 9670 -13085 9728 -13051
rect 9762 -13085 9820 -13051
rect 9854 -13085 9912 -13051
rect 9946 -13085 10004 -13051
rect 10038 -13085 10096 -13051
rect 10130 -13085 10188 -13051
rect 10222 -13085 10280 -13051
rect 10314 -13085 10372 -13051
rect 10406 -13085 10464 -13051
rect 10498 -13085 10556 -13051
rect 10590 -13085 10648 -13051
rect 10682 -13085 10740 -13051
rect 10774 -13085 10832 -13051
rect 10866 -13085 10924 -13051
rect 10958 -13085 11016 -13051
rect 11050 -13085 11108 -13051
rect 11142 -13085 11200 -13051
rect 11234 -13085 11292 -13051
rect 11326 -13085 11384 -13051
rect 11418 -13085 11476 -13051
rect 11510 -13085 11568 -13051
rect 11602 -13085 11660 -13051
rect 11694 -13085 11752 -13051
rect 11786 -13085 11844 -13051
rect 11878 -13085 11936 -13051
rect 11970 -13085 12028 -13051
rect 12062 -13085 12120 -13051
rect 12154 -13085 12212 -13051
rect 12246 -13085 12304 -13051
rect 12338 -13085 12396 -13051
rect 12430 -13085 12488 -13051
rect 12522 -13085 12580 -13051
rect 12614 -13085 12672 -13051
rect 12706 -13085 12764 -13051
rect 12798 -13085 12856 -13051
rect 12890 -13085 12948 -13051
rect 12982 -13085 13040 -13051
rect 13074 -13085 13132 -13051
rect 13166 -13085 13224 -13051
rect 13258 -13085 13316 -13051
rect 13350 -13085 13408 -13051
rect 13442 -13085 13500 -13051
rect 13534 -13085 13592 -13051
rect 13626 -13085 13684 -13051
rect 13718 -13085 13776 -13051
rect 13810 -13085 13868 -13051
rect 13902 -13085 13960 -13051
rect 13994 -13085 14052 -13051
rect 14086 -13085 14144 -13051
rect 14178 -13085 14236 -13051
rect 14270 -13085 14328 -13051
rect 14362 -13085 14420 -13051
rect 14454 -13085 14512 -13051
rect 14546 -13085 14604 -13051
rect 14638 -13085 14696 -13051
rect 14730 -13085 14788 -13051
rect 14822 -13085 14880 -13051
rect 14914 -13085 14972 -13051
rect 15006 -13085 15064 -13051
rect 15098 -13085 15156 -13051
rect 15190 -13085 15248 -13051
rect 15282 -13085 15340 -13051
rect 15374 -13085 15432 -13051
rect 15466 -13085 15524 -13051
rect 15558 -13085 15616 -13051
rect 15650 -13085 15708 -13051
rect 15742 -13085 15800 -13051
rect 15834 -13085 15892 -13051
rect 15926 -13085 15984 -13051
rect 16018 -13085 16076 -13051
rect 16110 -13085 16168 -13051
rect 16202 -13085 16260 -13051
rect 16294 -13085 16352 -13051
rect 16386 -13085 16444 -13051
rect 16478 -13085 16536 -13051
rect 16570 -13085 16628 -13051
rect 16662 -13085 16691 -13051
rect -2980 -13127 -2278 -13085
rect -2980 -13161 -2962 -13127
rect -2928 -13161 -2330 -13127
rect -2296 -13161 -2278 -13127
rect -2980 -13229 -2278 -13161
rect -2980 -13263 -2962 -13229
rect -2928 -13263 -2330 -13229
rect -2296 -13263 -2278 -13229
rect -2980 -13303 -2278 -13263
rect -2980 -13371 -2902 -13337
rect -2868 -13371 -2803 -13337
rect -2769 -13371 -2704 -13337
rect -2670 -13371 -2650 -13337
rect -2980 -13441 -2650 -13371
rect -2616 -13373 -2278 -13303
rect -2244 -13156 -2186 -13085
rect -2244 -13190 -2232 -13156
rect -2198 -13190 -2186 -13156
rect -2244 -13249 -2186 -13190
rect -2244 -13283 -2232 -13249
rect -2198 -13283 -2186 -13249
rect -2244 -13318 -2186 -13283
rect -1600 -13127 -898 -13085
rect -1600 -13161 -1582 -13127
rect -1548 -13161 -950 -13127
rect -916 -13161 -898 -13127
rect -1600 -13229 -898 -13161
rect -1600 -13263 -1582 -13229
rect -1548 -13263 -950 -13229
rect -916 -13263 -898 -13229
rect -1600 -13303 -898 -13263
rect -864 -13127 -162 -13085
rect -864 -13161 -846 -13127
rect -812 -13161 -214 -13127
rect -180 -13161 -162 -13127
rect -864 -13229 -162 -13161
rect -864 -13263 -846 -13229
rect -812 -13263 -214 -13229
rect -180 -13263 -162 -13229
rect -864 -13303 -162 -13263
rect -128 -13156 -70 -13085
rect -128 -13190 -116 -13156
rect -82 -13190 -70 -13156
rect -128 -13249 -70 -13190
rect -128 -13283 -116 -13249
rect -82 -13283 -70 -13249
rect -2616 -13407 -2596 -13373
rect -2562 -13407 -2493 -13373
rect -2459 -13407 -2390 -13373
rect -2356 -13407 -2278 -13373
rect -1600 -13373 -1262 -13303
rect -1600 -13407 -1522 -13373
rect -1488 -13407 -1419 -13373
rect -1385 -13407 -1316 -13373
rect -1282 -13407 -1262 -13373
rect -1228 -13371 -1208 -13337
rect -1174 -13371 -1109 -13337
rect -1075 -13371 -1010 -13337
rect -976 -13371 -898 -13337
rect -1228 -13441 -898 -13371
rect -864 -13373 -526 -13303
rect -128 -13318 -70 -13283
rect -36 -13127 298 -13085
rect -36 -13161 -18 -13127
rect 16 -13161 246 -13127
rect 280 -13161 298 -13127
rect -36 -13229 298 -13161
rect -36 -13263 -18 -13229
rect 16 -13263 246 -13229
rect 280 -13263 298 -13229
rect -36 -13303 298 -13263
rect 332 -13156 390 -13085
rect 332 -13190 344 -13156
rect 378 -13190 390 -13156
rect 332 -13249 390 -13190
rect 332 -13283 344 -13249
rect 378 -13283 390 -13249
rect -864 -13407 -786 -13373
rect -752 -13407 -683 -13373
rect -649 -13407 -580 -13373
rect -546 -13407 -526 -13373
rect -492 -13371 -472 -13337
rect -438 -13371 -373 -13337
rect -339 -13371 -274 -13337
rect -240 -13371 -162 -13337
rect -492 -13441 -162 -13371
rect -36 -13373 114 -13303
rect 332 -13318 390 -13283
rect 424 -13135 505 -13119
rect 424 -13169 457 -13135
rect 491 -13169 505 -13135
rect 424 -13203 505 -13169
rect 424 -13237 457 -13203
rect 491 -13237 505 -13203
rect 424 -13274 505 -13237
rect 539 -13134 605 -13085
rect 539 -13168 555 -13134
rect 589 -13168 605 -13134
rect 539 -13202 605 -13168
rect 539 -13236 555 -13202
rect 589 -13236 605 -13202
rect 539 -13245 605 -13236
rect 695 -13135 745 -13119
rect 695 -13169 711 -13135
rect 695 -13203 745 -13169
rect 695 -13237 711 -13203
rect 424 -13324 474 -13274
rect 695 -13279 745 -13237
rect -36 -13407 -16 -13373
rect 18 -13407 114 -13373
rect 148 -13371 244 -13337
rect 278 -13371 298 -13337
rect 148 -13441 298 -13371
rect -2980 -13500 -2278 -13441
rect -2980 -13534 -2962 -13500
rect -2928 -13534 -2330 -13500
rect -2296 -13534 -2278 -13500
rect -2980 -13595 -2278 -13534
rect -2244 -13467 -2186 -13450
rect -2244 -13501 -2232 -13467
rect -2198 -13501 -2186 -13467
rect -2244 -13595 -2186 -13501
rect -1600 -13500 -898 -13441
rect -1600 -13534 -1582 -13500
rect -1548 -13534 -950 -13500
rect -916 -13534 -898 -13500
rect -1600 -13595 -898 -13534
rect -864 -13500 -162 -13441
rect -864 -13534 -846 -13500
rect -812 -13534 -214 -13500
rect -180 -13534 -162 -13500
rect -864 -13595 -162 -13534
rect -128 -13467 -70 -13450
rect -128 -13501 -116 -13467
rect -82 -13501 -70 -13467
rect -128 -13595 -70 -13501
rect -36 -13493 298 -13441
rect 424 -13358 432 -13324
rect 466 -13358 474 -13324
rect 627 -13313 745 -13279
rect 797 -13134 867 -13119
rect 797 -13168 815 -13134
rect 849 -13168 867 -13134
rect 797 -13202 867 -13168
rect 797 -13236 815 -13202
rect 849 -13236 867 -13202
rect 627 -13347 661 -13313
rect -36 -13527 -18 -13493
rect 16 -13527 246 -13493
rect 280 -13527 298 -13493
rect -36 -13595 298 -13527
rect 332 -13467 390 -13450
rect 332 -13501 344 -13467
rect 378 -13501 390 -13467
rect 332 -13595 390 -13501
rect 424 -13484 474 -13358
rect 508 -13363 661 -13347
rect 797 -13348 867 -13236
rect 957 -13134 1023 -13085
rect 957 -13168 973 -13134
rect 1007 -13168 1023 -13134
rect 957 -13202 1023 -13168
rect 957 -13236 973 -13202
rect 1007 -13236 1023 -13202
rect 957 -13252 1023 -13236
rect 1057 -13134 1126 -13119
rect 1057 -13168 1073 -13134
rect 1107 -13168 1126 -13134
rect 1057 -13202 1126 -13168
rect 1057 -13236 1073 -13202
rect 1107 -13236 1126 -13202
rect 1057 -13286 1126 -13236
rect 508 -13397 511 -13363
rect 545 -13397 661 -13363
rect 508 -13413 661 -13397
rect 695 -13363 867 -13348
rect 932 -13320 1126 -13286
rect 1160 -13156 1218 -13085
rect 1160 -13190 1172 -13156
rect 1206 -13190 1218 -13156
rect 1160 -13249 1218 -13190
rect 1160 -13283 1172 -13249
rect 1206 -13283 1218 -13249
rect 1160 -13318 1218 -13283
rect 1252 -13127 1586 -13085
rect 1252 -13161 1270 -13127
rect 1304 -13161 1534 -13127
rect 1568 -13161 1586 -13127
rect 1252 -13229 1586 -13161
rect 1252 -13263 1270 -13229
rect 1304 -13263 1534 -13229
rect 1568 -13263 1586 -13229
rect 1252 -13303 1586 -13263
rect 1620 -13156 1678 -13085
rect 1620 -13190 1632 -13156
rect 1666 -13190 1678 -13156
rect 1620 -13249 1678 -13190
rect 1620 -13283 1632 -13249
rect 1666 -13283 1678 -13249
rect 932 -13349 1002 -13320
rect 695 -13397 711 -13363
rect 745 -13397 867 -13363
rect 695 -13398 867 -13397
rect 627 -13432 661 -13413
rect 627 -13466 745 -13432
rect 424 -13508 505 -13484
rect 424 -13542 457 -13508
rect 491 -13542 505 -13508
rect 424 -13561 505 -13542
rect 539 -13508 605 -13492
rect 539 -13542 555 -13508
rect 589 -13542 605 -13508
rect 539 -13595 605 -13542
rect 695 -13508 745 -13466
rect 695 -13542 711 -13508
rect 695 -13561 745 -13542
rect 797 -13508 867 -13398
rect 916 -13363 1002 -13349
rect 916 -13397 932 -13363
rect 966 -13397 1002 -13363
rect 1036 -13359 1126 -13354
rect 1036 -13397 1052 -13359
rect 1086 -13397 1126 -13359
rect 1252 -13373 1402 -13303
rect 1620 -13318 1678 -13283
rect 1712 -13127 2414 -13085
rect 1712 -13161 1730 -13127
rect 1764 -13161 2362 -13127
rect 2396 -13161 2414 -13127
rect 1712 -13229 2414 -13161
rect 1712 -13263 1730 -13229
rect 1764 -13263 2362 -13229
rect 2396 -13263 2414 -13229
rect 1712 -13303 2414 -13263
rect 916 -13407 1002 -13397
rect 1252 -13407 1272 -13373
rect 1306 -13407 1402 -13373
rect 1436 -13371 1532 -13337
rect 1566 -13371 1586 -13337
rect 932 -13431 1002 -13407
rect 932 -13465 1126 -13431
rect 1436 -13441 1586 -13371
rect 797 -13542 816 -13508
rect 850 -13542 867 -13508
rect 797 -13561 867 -13542
rect 960 -13508 1026 -13499
rect 960 -13542 976 -13508
rect 1010 -13542 1026 -13508
rect 960 -13595 1026 -13542
rect 1060 -13508 1126 -13465
rect 1060 -13542 1073 -13508
rect 1107 -13542 1126 -13508
rect 1060 -13561 1126 -13542
rect 1160 -13467 1218 -13450
rect 1160 -13501 1172 -13467
rect 1206 -13501 1218 -13467
rect 1160 -13595 1218 -13501
rect 1252 -13493 1586 -13441
rect 1712 -13371 1790 -13337
rect 1824 -13371 1889 -13337
rect 1923 -13371 1988 -13337
rect 2022 -13371 2042 -13337
rect 1712 -13441 2042 -13371
rect 2076 -13373 2414 -13303
rect 2448 -13156 2506 -13085
rect 2448 -13190 2460 -13156
rect 2494 -13190 2506 -13156
rect 2448 -13249 2506 -13190
rect 2448 -13283 2460 -13249
rect 2494 -13283 2506 -13249
rect 2448 -13318 2506 -13283
rect 2540 -13127 2874 -13085
rect 2540 -13161 2558 -13127
rect 2592 -13161 2822 -13127
rect 2856 -13161 2874 -13127
rect 2540 -13229 2874 -13161
rect 2540 -13263 2558 -13229
rect 2592 -13263 2822 -13229
rect 2856 -13263 2874 -13229
rect 2540 -13303 2874 -13263
rect 2908 -13156 2966 -13085
rect 2908 -13190 2920 -13156
rect 2954 -13190 2966 -13156
rect 2908 -13249 2966 -13190
rect 2908 -13283 2920 -13249
rect 2954 -13283 2966 -13249
rect 2076 -13407 2096 -13373
rect 2130 -13407 2199 -13373
rect 2233 -13407 2302 -13373
rect 2336 -13407 2414 -13373
rect 2540 -13373 2690 -13303
rect 2908 -13318 2966 -13283
rect 3000 -13135 3081 -13119
rect 3000 -13169 3033 -13135
rect 3067 -13169 3081 -13135
rect 3000 -13203 3081 -13169
rect 3000 -13237 3033 -13203
rect 3067 -13237 3081 -13203
rect 3000 -13274 3081 -13237
rect 3115 -13134 3181 -13085
rect 3115 -13168 3131 -13134
rect 3165 -13168 3181 -13134
rect 3115 -13202 3181 -13168
rect 3115 -13236 3131 -13202
rect 3165 -13236 3181 -13202
rect 3115 -13245 3181 -13236
rect 3271 -13135 3321 -13119
rect 3271 -13169 3287 -13135
rect 3271 -13203 3321 -13169
rect 3271 -13237 3287 -13203
rect 2540 -13407 2560 -13373
rect 2594 -13407 2690 -13373
rect 2724 -13371 2820 -13337
rect 2854 -13371 2874 -13337
rect 2724 -13441 2874 -13371
rect 1252 -13527 1270 -13493
rect 1304 -13527 1534 -13493
rect 1568 -13527 1586 -13493
rect 1252 -13595 1586 -13527
rect 1620 -13467 1678 -13450
rect 1620 -13501 1632 -13467
rect 1666 -13501 1678 -13467
rect 1620 -13595 1678 -13501
rect 1712 -13500 2414 -13441
rect 1712 -13534 1730 -13500
rect 1764 -13534 2362 -13500
rect 2396 -13534 2414 -13500
rect 1712 -13595 2414 -13534
rect 2448 -13467 2506 -13450
rect 2448 -13501 2460 -13467
rect 2494 -13501 2506 -13467
rect 2448 -13595 2506 -13501
rect 2540 -13493 2874 -13441
rect 3000 -13359 3050 -13274
rect 3271 -13279 3321 -13237
rect 3203 -13313 3321 -13279
rect 3373 -13134 3443 -13119
rect 3373 -13168 3391 -13134
rect 3425 -13168 3443 -13134
rect 3373 -13202 3443 -13168
rect 3373 -13236 3391 -13202
rect 3425 -13236 3443 -13202
rect 3203 -13347 3237 -13313
rect 3000 -13393 3012 -13359
rect 3046 -13393 3050 -13359
rect 2540 -13527 2558 -13493
rect 2592 -13527 2822 -13493
rect 2856 -13527 2874 -13493
rect 2540 -13595 2874 -13527
rect 2908 -13467 2966 -13450
rect 2908 -13501 2920 -13467
rect 2954 -13501 2966 -13467
rect 2908 -13595 2966 -13501
rect 3000 -13484 3050 -13393
rect 3084 -13363 3237 -13347
rect 3373 -13348 3443 -13236
rect 3533 -13134 3599 -13085
rect 3533 -13168 3549 -13134
rect 3583 -13168 3599 -13134
rect 3533 -13202 3599 -13168
rect 3533 -13236 3549 -13202
rect 3583 -13236 3599 -13202
rect 3533 -13252 3599 -13236
rect 3633 -13134 3702 -13119
rect 3633 -13168 3649 -13134
rect 3683 -13168 3702 -13134
rect 3633 -13202 3702 -13168
rect 3633 -13236 3649 -13202
rect 3683 -13236 3702 -13202
rect 3633 -13286 3702 -13236
rect 3084 -13397 3087 -13363
rect 3121 -13397 3237 -13363
rect 3084 -13413 3237 -13397
rect 3271 -13363 3443 -13348
rect 3508 -13320 3702 -13286
rect 3736 -13156 3794 -13085
rect 3736 -13190 3748 -13156
rect 3782 -13190 3794 -13156
rect 3736 -13249 3794 -13190
rect 3736 -13283 3748 -13249
rect 3782 -13283 3794 -13249
rect 3736 -13318 3794 -13283
rect 3828 -13127 4162 -13085
rect 3828 -13161 3846 -13127
rect 3880 -13161 4110 -13127
rect 4144 -13161 4162 -13127
rect 3828 -13229 4162 -13161
rect 3828 -13263 3846 -13229
rect 3880 -13263 4110 -13229
rect 4144 -13263 4162 -13229
rect 3828 -13303 4162 -13263
rect 4196 -13156 4254 -13085
rect 4196 -13190 4208 -13156
rect 4242 -13190 4254 -13156
rect 4196 -13249 4254 -13190
rect 4196 -13283 4208 -13249
rect 4242 -13283 4254 -13249
rect 3508 -13349 3578 -13320
rect 3271 -13397 3287 -13363
rect 3321 -13397 3443 -13363
rect 3271 -13398 3443 -13397
rect 3203 -13432 3237 -13413
rect 3203 -13466 3321 -13432
rect 3000 -13508 3081 -13484
rect 3000 -13542 3033 -13508
rect 3067 -13542 3081 -13508
rect 3000 -13561 3081 -13542
rect 3115 -13508 3181 -13492
rect 3115 -13542 3131 -13508
rect 3165 -13542 3181 -13508
rect 3115 -13595 3181 -13542
rect 3271 -13508 3321 -13466
rect 3271 -13542 3287 -13508
rect 3271 -13561 3321 -13542
rect 3373 -13508 3443 -13398
rect 3492 -13363 3578 -13349
rect 3492 -13397 3508 -13363
rect 3542 -13397 3578 -13363
rect 3612 -13359 3702 -13354
rect 3612 -13393 3626 -13359
rect 3660 -13363 3702 -13359
rect 3612 -13397 3628 -13393
rect 3662 -13397 3702 -13363
rect 3828 -13373 3978 -13303
rect 4196 -13318 4254 -13283
rect 4288 -13127 4990 -13085
rect 4288 -13161 4306 -13127
rect 4340 -13161 4938 -13127
rect 4972 -13161 4990 -13127
rect 4288 -13229 4990 -13161
rect 4288 -13263 4306 -13229
rect 4340 -13263 4938 -13229
rect 4972 -13263 4990 -13229
rect 4288 -13303 4990 -13263
rect 3492 -13407 3578 -13397
rect 3828 -13407 3848 -13373
rect 3882 -13407 3978 -13373
rect 4012 -13371 4108 -13337
rect 4142 -13371 4162 -13337
rect 3508 -13431 3578 -13407
rect 3508 -13465 3702 -13431
rect 4012 -13441 4162 -13371
rect 3373 -13542 3392 -13508
rect 3426 -13542 3443 -13508
rect 3373 -13561 3443 -13542
rect 3536 -13508 3602 -13499
rect 3536 -13542 3552 -13508
rect 3586 -13542 3602 -13508
rect 3536 -13595 3602 -13542
rect 3636 -13508 3702 -13465
rect 3636 -13542 3649 -13508
rect 3683 -13542 3702 -13508
rect 3636 -13561 3702 -13542
rect 3736 -13467 3794 -13450
rect 3736 -13501 3748 -13467
rect 3782 -13501 3794 -13467
rect 3736 -13595 3794 -13501
rect 3828 -13493 4162 -13441
rect 4288 -13371 4366 -13337
rect 4400 -13371 4465 -13337
rect 4499 -13371 4564 -13337
rect 4598 -13371 4618 -13337
rect 4288 -13441 4618 -13371
rect 4652 -13373 4990 -13303
rect 5024 -13156 5082 -13085
rect 5024 -13190 5036 -13156
rect 5070 -13190 5082 -13156
rect 5024 -13249 5082 -13190
rect 5024 -13283 5036 -13249
rect 5070 -13283 5082 -13249
rect 5024 -13318 5082 -13283
rect 5116 -13127 5450 -13085
rect 5116 -13161 5134 -13127
rect 5168 -13161 5398 -13127
rect 5432 -13161 5450 -13127
rect 5116 -13229 5450 -13161
rect 5116 -13263 5134 -13229
rect 5168 -13263 5398 -13229
rect 5432 -13263 5450 -13229
rect 5116 -13303 5450 -13263
rect 5484 -13156 5542 -13085
rect 5484 -13190 5496 -13156
rect 5530 -13190 5542 -13156
rect 5484 -13249 5542 -13190
rect 5484 -13283 5496 -13249
rect 5530 -13283 5542 -13249
rect 4652 -13407 4672 -13373
rect 4706 -13407 4775 -13373
rect 4809 -13407 4878 -13373
rect 4912 -13407 4990 -13373
rect 5116 -13373 5266 -13303
rect 5484 -13318 5542 -13283
rect 5576 -13135 5657 -13119
rect 5576 -13169 5609 -13135
rect 5643 -13169 5657 -13135
rect 5576 -13203 5657 -13169
rect 5576 -13237 5609 -13203
rect 5643 -13237 5657 -13203
rect 5576 -13274 5657 -13237
rect 5691 -13134 5757 -13085
rect 5691 -13168 5707 -13134
rect 5741 -13168 5757 -13134
rect 5691 -13202 5757 -13168
rect 5691 -13236 5707 -13202
rect 5741 -13236 5757 -13202
rect 5691 -13245 5757 -13236
rect 5847 -13135 5897 -13119
rect 5847 -13169 5863 -13135
rect 5847 -13203 5897 -13169
rect 5847 -13237 5863 -13203
rect 5116 -13407 5136 -13373
rect 5170 -13407 5266 -13373
rect 5300 -13371 5396 -13337
rect 5430 -13371 5450 -13337
rect 5300 -13441 5450 -13371
rect 3828 -13527 3846 -13493
rect 3880 -13527 4110 -13493
rect 4144 -13527 4162 -13493
rect 3828 -13595 4162 -13527
rect 4196 -13467 4254 -13450
rect 4196 -13501 4208 -13467
rect 4242 -13501 4254 -13467
rect 4196 -13595 4254 -13501
rect 4288 -13500 4990 -13441
rect 4288 -13534 4306 -13500
rect 4340 -13534 4938 -13500
rect 4972 -13534 4990 -13500
rect 4288 -13595 4990 -13534
rect 5024 -13467 5082 -13450
rect 5024 -13501 5036 -13467
rect 5070 -13501 5082 -13467
rect 5024 -13595 5082 -13501
rect 5116 -13493 5450 -13441
rect 5576 -13359 5626 -13274
rect 5847 -13279 5897 -13237
rect 5779 -13313 5897 -13279
rect 5949 -13134 6019 -13119
rect 5949 -13168 5967 -13134
rect 6001 -13168 6019 -13134
rect 5949 -13202 6019 -13168
rect 5949 -13236 5967 -13202
rect 6001 -13236 6019 -13202
rect 5779 -13347 5813 -13313
rect 5576 -13393 5586 -13359
rect 5620 -13393 5626 -13359
rect 5116 -13527 5134 -13493
rect 5168 -13527 5398 -13493
rect 5432 -13527 5450 -13493
rect 5116 -13595 5450 -13527
rect 5484 -13467 5542 -13450
rect 5484 -13501 5496 -13467
rect 5530 -13501 5542 -13467
rect 5484 -13595 5542 -13501
rect 5576 -13484 5626 -13393
rect 5660 -13363 5813 -13347
rect 5949 -13348 6019 -13236
rect 6109 -13134 6175 -13085
rect 6109 -13168 6125 -13134
rect 6159 -13168 6175 -13134
rect 6109 -13202 6175 -13168
rect 6109 -13236 6125 -13202
rect 6159 -13236 6175 -13202
rect 6109 -13252 6175 -13236
rect 6209 -13134 6278 -13119
rect 6209 -13168 6225 -13134
rect 6259 -13168 6278 -13134
rect 6209 -13202 6278 -13168
rect 6209 -13236 6225 -13202
rect 6259 -13236 6278 -13202
rect 6209 -13286 6278 -13236
rect 5660 -13397 5663 -13363
rect 5697 -13397 5813 -13363
rect 5660 -13413 5813 -13397
rect 5847 -13363 6019 -13348
rect 6084 -13320 6278 -13286
rect 6312 -13156 6370 -13085
rect 6312 -13190 6324 -13156
rect 6358 -13190 6370 -13156
rect 6312 -13249 6370 -13190
rect 6312 -13283 6324 -13249
rect 6358 -13283 6370 -13249
rect 6312 -13318 6370 -13283
rect 6404 -13127 6738 -13085
rect 6404 -13161 6422 -13127
rect 6456 -13161 6686 -13127
rect 6720 -13161 6738 -13127
rect 6404 -13229 6738 -13161
rect 6404 -13263 6422 -13229
rect 6456 -13263 6686 -13229
rect 6720 -13263 6738 -13229
rect 6404 -13303 6738 -13263
rect 6772 -13156 6830 -13085
rect 6772 -13190 6784 -13156
rect 6818 -13190 6830 -13156
rect 6772 -13249 6830 -13190
rect 6772 -13283 6784 -13249
rect 6818 -13283 6830 -13249
rect 6084 -13349 6154 -13320
rect 5847 -13397 5863 -13363
rect 5897 -13397 6019 -13363
rect 5847 -13398 6019 -13397
rect 5779 -13432 5813 -13413
rect 5779 -13466 5897 -13432
rect 5576 -13508 5657 -13484
rect 5576 -13542 5609 -13508
rect 5643 -13542 5657 -13508
rect 5576 -13561 5657 -13542
rect 5691 -13508 5757 -13492
rect 5691 -13542 5707 -13508
rect 5741 -13542 5757 -13508
rect 5691 -13595 5757 -13542
rect 5847 -13508 5897 -13466
rect 5847 -13542 5863 -13508
rect 5847 -13561 5897 -13542
rect 5949 -13508 6019 -13398
rect 6068 -13363 6154 -13349
rect 6068 -13397 6084 -13363
rect 6118 -13397 6154 -13363
rect 6188 -13359 6278 -13354
rect 6188 -13393 6200 -13359
rect 6234 -13363 6278 -13359
rect 6188 -13397 6204 -13393
rect 6238 -13397 6278 -13363
rect 6404 -13373 6554 -13303
rect 6772 -13318 6830 -13283
rect 6864 -13127 7566 -13085
rect 6864 -13161 6882 -13127
rect 6916 -13161 7514 -13127
rect 7548 -13161 7566 -13127
rect 6864 -13229 7566 -13161
rect 6864 -13263 6882 -13229
rect 6916 -13263 7514 -13229
rect 7548 -13263 7566 -13229
rect 6864 -13303 7566 -13263
rect 6068 -13407 6154 -13397
rect 6404 -13407 6424 -13373
rect 6458 -13407 6554 -13373
rect 6588 -13371 6684 -13337
rect 6718 -13371 6738 -13337
rect 6084 -13431 6154 -13407
rect 6084 -13465 6278 -13431
rect 6588 -13441 6738 -13371
rect 5949 -13542 5968 -13508
rect 6002 -13542 6019 -13508
rect 5949 -13561 6019 -13542
rect 6112 -13508 6178 -13499
rect 6112 -13542 6128 -13508
rect 6162 -13542 6178 -13508
rect 6112 -13595 6178 -13542
rect 6212 -13508 6278 -13465
rect 6212 -13542 6225 -13508
rect 6259 -13542 6278 -13508
rect 6212 -13561 6278 -13542
rect 6312 -13467 6370 -13450
rect 6312 -13501 6324 -13467
rect 6358 -13501 6370 -13467
rect 6312 -13595 6370 -13501
rect 6404 -13493 6738 -13441
rect 6864 -13371 6942 -13337
rect 6976 -13371 7041 -13337
rect 7075 -13371 7140 -13337
rect 7174 -13371 7194 -13337
rect 6864 -13441 7194 -13371
rect 7228 -13373 7566 -13303
rect 7600 -13156 7658 -13085
rect 7600 -13190 7612 -13156
rect 7646 -13190 7658 -13156
rect 7600 -13249 7658 -13190
rect 7600 -13283 7612 -13249
rect 7646 -13283 7658 -13249
rect 7600 -13318 7658 -13283
rect 7692 -13127 8026 -13085
rect 7692 -13161 7710 -13127
rect 7744 -13161 7974 -13127
rect 8008 -13161 8026 -13127
rect 7692 -13229 8026 -13161
rect 7692 -13263 7710 -13229
rect 7744 -13263 7974 -13229
rect 8008 -13263 8026 -13229
rect 7692 -13303 8026 -13263
rect 8060 -13156 8118 -13085
rect 8060 -13190 8072 -13156
rect 8106 -13190 8118 -13156
rect 8060 -13249 8118 -13190
rect 8060 -13283 8072 -13249
rect 8106 -13283 8118 -13249
rect 7228 -13407 7248 -13373
rect 7282 -13407 7351 -13373
rect 7385 -13407 7454 -13373
rect 7488 -13407 7566 -13373
rect 7692 -13373 7842 -13303
rect 8060 -13318 8118 -13283
rect 8152 -13135 8233 -13119
rect 8152 -13169 8185 -13135
rect 8219 -13169 8233 -13135
rect 8152 -13203 8233 -13169
rect 8152 -13237 8185 -13203
rect 8219 -13237 8233 -13203
rect 8152 -13274 8233 -13237
rect 8267 -13134 8333 -13085
rect 8267 -13168 8283 -13134
rect 8317 -13168 8333 -13134
rect 8267 -13202 8333 -13168
rect 8267 -13236 8283 -13202
rect 8317 -13236 8333 -13202
rect 8267 -13245 8333 -13236
rect 8423 -13135 8473 -13119
rect 8423 -13169 8439 -13135
rect 8423 -13203 8473 -13169
rect 8423 -13237 8439 -13203
rect 7692 -13407 7712 -13373
rect 7746 -13407 7842 -13373
rect 7876 -13371 7972 -13337
rect 8006 -13371 8026 -13337
rect 7876 -13441 8026 -13371
rect 6404 -13527 6422 -13493
rect 6456 -13527 6686 -13493
rect 6720 -13527 6738 -13493
rect 6404 -13595 6738 -13527
rect 6772 -13467 6830 -13450
rect 6772 -13501 6784 -13467
rect 6818 -13501 6830 -13467
rect 6772 -13595 6830 -13501
rect 6864 -13500 7566 -13441
rect 6864 -13534 6882 -13500
rect 6916 -13534 7514 -13500
rect 7548 -13534 7566 -13500
rect 6864 -13595 7566 -13534
rect 7600 -13467 7658 -13450
rect 7600 -13501 7612 -13467
rect 7646 -13501 7658 -13467
rect 7600 -13595 7658 -13501
rect 7692 -13493 8026 -13441
rect 8152 -13359 8202 -13274
rect 8423 -13279 8473 -13237
rect 8355 -13313 8473 -13279
rect 8525 -13134 8595 -13119
rect 8525 -13168 8543 -13134
rect 8577 -13168 8595 -13134
rect 8525 -13202 8595 -13168
rect 8525 -13236 8543 -13202
rect 8577 -13236 8595 -13202
rect 8355 -13347 8389 -13313
rect 8152 -13393 8160 -13359
rect 8194 -13393 8202 -13359
rect 7692 -13527 7710 -13493
rect 7744 -13527 7974 -13493
rect 8008 -13527 8026 -13493
rect 7692 -13595 8026 -13527
rect 8060 -13467 8118 -13450
rect 8060 -13501 8072 -13467
rect 8106 -13501 8118 -13467
rect 8060 -13595 8118 -13501
rect 8152 -13484 8202 -13393
rect 8236 -13363 8389 -13347
rect 8525 -13348 8595 -13236
rect 8685 -13134 8751 -13085
rect 8685 -13168 8701 -13134
rect 8735 -13168 8751 -13134
rect 8685 -13202 8751 -13168
rect 8685 -13236 8701 -13202
rect 8735 -13236 8751 -13202
rect 8685 -13252 8751 -13236
rect 8785 -13134 8854 -13119
rect 8785 -13168 8801 -13134
rect 8835 -13168 8854 -13134
rect 8785 -13202 8854 -13168
rect 8785 -13236 8801 -13202
rect 8835 -13236 8854 -13202
rect 8785 -13286 8854 -13236
rect 8236 -13397 8239 -13363
rect 8273 -13397 8389 -13363
rect 8236 -13413 8389 -13397
rect 8423 -13363 8595 -13348
rect 8660 -13320 8854 -13286
rect 8888 -13156 8946 -13085
rect 8888 -13190 8900 -13156
rect 8934 -13190 8946 -13156
rect 8888 -13249 8946 -13190
rect 8888 -13283 8900 -13249
rect 8934 -13283 8946 -13249
rect 8888 -13318 8946 -13283
rect 8980 -13127 9314 -13085
rect 8980 -13161 8998 -13127
rect 9032 -13161 9262 -13127
rect 9296 -13161 9314 -13127
rect 8980 -13229 9314 -13161
rect 8980 -13263 8998 -13229
rect 9032 -13263 9262 -13229
rect 9296 -13263 9314 -13229
rect 8980 -13303 9314 -13263
rect 9348 -13156 9406 -13085
rect 9348 -13190 9360 -13156
rect 9394 -13190 9406 -13156
rect 9348 -13249 9406 -13190
rect 9348 -13283 9360 -13249
rect 9394 -13283 9406 -13249
rect 8660 -13349 8730 -13320
rect 8423 -13397 8439 -13363
rect 8473 -13397 8595 -13363
rect 8423 -13398 8595 -13397
rect 8355 -13432 8389 -13413
rect 8355 -13466 8473 -13432
rect 8152 -13508 8233 -13484
rect 8152 -13542 8185 -13508
rect 8219 -13542 8233 -13508
rect 8152 -13561 8233 -13542
rect 8267 -13508 8333 -13492
rect 8267 -13542 8283 -13508
rect 8317 -13542 8333 -13508
rect 8267 -13595 8333 -13542
rect 8423 -13508 8473 -13466
rect 8423 -13542 8439 -13508
rect 8423 -13561 8473 -13542
rect 8525 -13508 8595 -13398
rect 8644 -13363 8730 -13349
rect 8644 -13397 8660 -13363
rect 8694 -13397 8730 -13363
rect 8764 -13359 8854 -13354
rect 8764 -13393 8774 -13359
rect 8808 -13363 8854 -13359
rect 8764 -13397 8780 -13393
rect 8814 -13397 8854 -13363
rect 8980 -13373 9130 -13303
rect 9348 -13318 9406 -13283
rect 9440 -13127 10142 -13085
rect 9440 -13161 9458 -13127
rect 9492 -13161 10090 -13127
rect 10124 -13161 10142 -13127
rect 9440 -13229 10142 -13161
rect 9440 -13263 9458 -13229
rect 9492 -13263 10090 -13229
rect 10124 -13263 10142 -13229
rect 9440 -13303 10142 -13263
rect 8644 -13407 8730 -13397
rect 8980 -13407 9000 -13373
rect 9034 -13407 9130 -13373
rect 9164 -13371 9260 -13337
rect 9294 -13371 9314 -13337
rect 8660 -13431 8730 -13407
rect 8660 -13465 8854 -13431
rect 9164 -13441 9314 -13371
rect 8525 -13542 8544 -13508
rect 8578 -13542 8595 -13508
rect 8525 -13561 8595 -13542
rect 8688 -13508 8754 -13499
rect 8688 -13542 8704 -13508
rect 8738 -13542 8754 -13508
rect 8688 -13595 8754 -13542
rect 8788 -13508 8854 -13465
rect 8788 -13542 8801 -13508
rect 8835 -13542 8854 -13508
rect 8788 -13561 8854 -13542
rect 8888 -13467 8946 -13450
rect 8888 -13501 8900 -13467
rect 8934 -13501 8946 -13467
rect 8888 -13595 8946 -13501
rect 8980 -13493 9314 -13441
rect 9440 -13371 9518 -13337
rect 9552 -13371 9617 -13337
rect 9651 -13371 9716 -13337
rect 9750 -13371 9770 -13337
rect 9440 -13441 9770 -13371
rect 9804 -13373 10142 -13303
rect 10176 -13156 10234 -13085
rect 10176 -13190 10188 -13156
rect 10222 -13190 10234 -13156
rect 10176 -13249 10234 -13190
rect 10176 -13283 10188 -13249
rect 10222 -13283 10234 -13249
rect 10176 -13318 10234 -13283
rect 10360 -13127 10694 -13085
rect 10360 -13161 10378 -13127
rect 10412 -13161 10642 -13127
rect 10676 -13161 10694 -13127
rect 10360 -13229 10694 -13161
rect 10360 -13263 10378 -13229
rect 10412 -13263 10642 -13229
rect 10676 -13263 10694 -13229
rect 10360 -13303 10694 -13263
rect 10728 -13135 10809 -13119
rect 10728 -13169 10761 -13135
rect 10795 -13169 10809 -13135
rect 10728 -13203 10809 -13169
rect 10728 -13237 10761 -13203
rect 10795 -13237 10809 -13203
rect 10728 -13274 10809 -13237
rect 10843 -13134 10909 -13085
rect 10843 -13168 10859 -13134
rect 10893 -13168 10909 -13134
rect 10843 -13202 10909 -13168
rect 10843 -13236 10859 -13202
rect 10893 -13236 10909 -13202
rect 10843 -13245 10909 -13236
rect 10999 -13135 11049 -13119
rect 10999 -13169 11015 -13135
rect 10999 -13203 11049 -13169
rect 10999 -13237 11015 -13203
rect 9804 -13407 9824 -13373
rect 9858 -13407 9927 -13373
rect 9961 -13407 10030 -13373
rect 10064 -13407 10142 -13373
rect 10360 -13373 10510 -13303
rect 10360 -13407 10380 -13373
rect 10414 -13407 10510 -13373
rect 10544 -13371 10640 -13337
rect 10674 -13371 10694 -13337
rect 10544 -13441 10694 -13371
rect 8980 -13527 8998 -13493
rect 9032 -13527 9262 -13493
rect 9296 -13527 9314 -13493
rect 8980 -13595 9314 -13527
rect 9348 -13467 9406 -13450
rect 9348 -13501 9360 -13467
rect 9394 -13501 9406 -13467
rect 9348 -13595 9406 -13501
rect 9440 -13500 10142 -13441
rect 9440 -13534 9458 -13500
rect 9492 -13534 10090 -13500
rect 10124 -13534 10142 -13500
rect 9440 -13595 10142 -13534
rect 10176 -13467 10234 -13450
rect 10176 -13501 10188 -13467
rect 10222 -13501 10234 -13467
rect 10176 -13595 10234 -13501
rect 10360 -13493 10694 -13441
rect 10360 -13527 10378 -13493
rect 10412 -13527 10642 -13493
rect 10676 -13527 10694 -13493
rect 10360 -13595 10694 -13527
rect 10728 -13357 10778 -13274
rect 10999 -13279 11049 -13237
rect 10931 -13313 11049 -13279
rect 11101 -13134 11171 -13119
rect 11101 -13168 11119 -13134
rect 11153 -13168 11171 -13134
rect 11101 -13202 11171 -13168
rect 11101 -13236 11119 -13202
rect 11153 -13236 11171 -13202
rect 10931 -13347 10965 -13313
rect 10728 -13391 10737 -13357
rect 10771 -13391 10778 -13357
rect 10728 -13484 10778 -13391
rect 10812 -13363 10965 -13347
rect 11101 -13348 11171 -13236
rect 11261 -13134 11327 -13085
rect 11261 -13168 11277 -13134
rect 11311 -13168 11327 -13134
rect 11261 -13202 11327 -13168
rect 11261 -13236 11277 -13202
rect 11311 -13236 11327 -13202
rect 11261 -13252 11327 -13236
rect 11361 -13134 11430 -13119
rect 11361 -13168 11377 -13134
rect 11411 -13168 11430 -13134
rect 11361 -13202 11430 -13168
rect 11361 -13236 11377 -13202
rect 11411 -13236 11430 -13202
rect 11361 -13286 11430 -13236
rect 10812 -13397 10815 -13363
rect 10849 -13397 10965 -13363
rect 10812 -13413 10965 -13397
rect 10999 -13363 11171 -13348
rect 11236 -13320 11430 -13286
rect 11464 -13156 11522 -13085
rect 11464 -13190 11476 -13156
rect 11510 -13190 11522 -13156
rect 11464 -13249 11522 -13190
rect 11464 -13283 11476 -13249
rect 11510 -13283 11522 -13249
rect 11464 -13318 11522 -13283
rect 11648 -13127 11982 -13085
rect 11648 -13161 11666 -13127
rect 11700 -13161 11930 -13127
rect 11964 -13161 11982 -13127
rect 11648 -13229 11982 -13161
rect 11648 -13263 11666 -13229
rect 11700 -13263 11930 -13229
rect 11964 -13263 11982 -13229
rect 11648 -13303 11982 -13263
rect 13580 -13156 13638 -13085
rect 13580 -13190 13592 -13156
rect 13626 -13190 13638 -13156
rect 13580 -13249 13638 -13190
rect 13674 -13127 13733 -13085
rect 13674 -13161 13690 -13127
rect 13724 -13161 13733 -13127
rect 13674 -13195 13733 -13161
rect 13674 -13229 13690 -13195
rect 13724 -13229 13733 -13195
rect 13674 -13247 13733 -13229
rect 13769 -13135 13818 -13119
rect 13769 -13169 13776 -13135
rect 13810 -13169 13818 -13135
rect 13769 -13203 13818 -13169
rect 13769 -13237 13776 -13203
rect 13810 -13237 13818 -13203
rect 13580 -13283 13592 -13249
rect 13626 -13283 13638 -13249
rect 11236 -13349 11306 -13320
rect 10999 -13397 11015 -13363
rect 11049 -13397 11171 -13363
rect 10999 -13398 11171 -13397
rect 10931 -13432 10965 -13413
rect 10931 -13466 11049 -13432
rect 10728 -13508 10809 -13484
rect 10728 -13542 10761 -13508
rect 10795 -13542 10809 -13508
rect 10728 -13561 10809 -13542
rect 10843 -13508 10909 -13492
rect 10843 -13542 10859 -13508
rect 10893 -13542 10909 -13508
rect 10843 -13595 10909 -13542
rect 10999 -13508 11049 -13466
rect 10999 -13542 11015 -13508
rect 10999 -13561 11049 -13542
rect 11101 -13508 11171 -13398
rect 11220 -13363 11306 -13349
rect 11220 -13397 11236 -13363
rect 11270 -13397 11306 -13363
rect 11340 -13356 11430 -13354
rect 11340 -13363 11369 -13356
rect 11340 -13397 11356 -13363
rect 11403 -13390 11430 -13356
rect 11390 -13397 11430 -13390
rect 11648 -13373 11798 -13303
rect 13580 -13318 13638 -13283
rect 11220 -13407 11306 -13397
rect 11648 -13407 11668 -13373
rect 11702 -13407 11798 -13373
rect 11832 -13371 11928 -13337
rect 11962 -13371 11982 -13337
rect 13769 -13347 13818 -13237
rect 13853 -13127 13905 -13085
rect 14025 -13086 15280 -13085
rect 13853 -13161 13862 -13127
rect 13896 -13161 13905 -13127
rect 13853 -13195 13905 -13161
rect 13853 -13229 13862 -13195
rect 13896 -13229 13905 -13195
rect 13853 -13247 13905 -13229
rect 13941 -13143 13991 -13120
rect 13941 -13177 13948 -13143
rect 13982 -13177 13991 -13143
rect 13941 -13211 13991 -13177
rect 13941 -13245 13948 -13211
rect 13982 -13245 13991 -13211
rect 14025 -13127 14077 -13086
rect 14025 -13161 14034 -13127
rect 14068 -13161 14077 -13127
rect 14025 -13195 14077 -13161
rect 14025 -13229 14034 -13195
rect 14068 -13229 14077 -13195
rect 14025 -13245 14077 -13229
rect 14111 -13171 14163 -13120
rect 14111 -13205 14120 -13171
rect 14154 -13205 14163 -13171
rect 13941 -13347 13991 -13245
rect 14111 -13257 14163 -13205
rect 14197 -13151 14249 -13086
rect 14197 -13185 14206 -13151
rect 14240 -13185 14249 -13151
rect 14197 -13231 14249 -13185
rect 14283 -13171 14335 -13120
rect 14283 -13205 14292 -13171
rect 14326 -13205 14335 -13171
rect 14111 -13291 14120 -13257
rect 14154 -13265 14163 -13257
rect 14283 -13257 14335 -13205
rect 14369 -13151 14421 -13086
rect 14369 -13185 14378 -13151
rect 14412 -13185 14421 -13151
rect 14369 -13231 14421 -13185
rect 14455 -13171 14507 -13120
rect 14455 -13205 14464 -13171
rect 14498 -13205 14507 -13171
rect 14283 -13265 14292 -13257
rect 14154 -13291 14292 -13265
rect 14326 -13265 14335 -13257
rect 14455 -13257 14507 -13205
rect 14541 -13151 14593 -13086
rect 14541 -13185 14550 -13151
rect 14584 -13185 14593 -13151
rect 14541 -13231 14593 -13185
rect 14627 -13171 14679 -13120
rect 14627 -13205 14636 -13171
rect 14670 -13205 14679 -13171
rect 14455 -13265 14464 -13257
rect 14326 -13291 14464 -13265
rect 14498 -13265 14507 -13257
rect 14627 -13257 14679 -13205
rect 14713 -13151 14762 -13086
rect 14713 -13185 14722 -13151
rect 14756 -13185 14762 -13151
rect 14713 -13231 14762 -13185
rect 14796 -13171 14848 -13120
rect 14796 -13205 14807 -13171
rect 14841 -13205 14848 -13171
rect 14627 -13265 14636 -13257
rect 14498 -13291 14636 -13265
rect 14670 -13265 14679 -13257
rect 14796 -13257 14848 -13205
rect 14885 -13151 14934 -13086
rect 14885 -13185 14893 -13151
rect 14927 -13185 14934 -13151
rect 14885 -13231 14934 -13185
rect 14968 -13171 15020 -13120
rect 14968 -13205 14979 -13171
rect 15013 -13205 15020 -13171
rect 14796 -13265 14807 -13257
rect 14670 -13291 14807 -13265
rect 14841 -13265 14848 -13257
rect 14968 -13257 15020 -13205
rect 15057 -13151 15106 -13086
rect 15057 -13185 15065 -13151
rect 15099 -13185 15106 -13151
rect 15057 -13231 15106 -13185
rect 15140 -13171 15192 -13120
rect 15140 -13205 15151 -13171
rect 15185 -13205 15192 -13171
rect 14968 -13265 14979 -13257
rect 14841 -13291 14979 -13265
rect 15013 -13265 15020 -13257
rect 15140 -13257 15192 -13205
rect 15229 -13151 15280 -13086
rect 15229 -13185 15237 -13151
rect 15271 -13185 15280 -13151
rect 15229 -13231 15280 -13185
rect 15314 -13171 15372 -13120
rect 15314 -13205 15323 -13171
rect 15357 -13205 15372 -13171
rect 15140 -13265 15151 -13257
rect 15013 -13291 15151 -13265
rect 15185 -13268 15192 -13257
rect 15314 -13257 15372 -13205
rect 15406 -13151 15460 -13085
rect 15406 -13185 15409 -13151
rect 15443 -13185 15460 -13151
rect 15406 -13234 15460 -13185
rect 15512 -13156 15570 -13085
rect 15512 -13190 15524 -13156
rect 15558 -13190 15570 -13156
rect 15314 -13268 15323 -13257
rect 15185 -13291 15323 -13268
rect 15357 -13268 15372 -13257
rect 15512 -13249 15570 -13190
rect 15357 -13291 15460 -13268
rect 14111 -13310 15460 -13291
rect 14111 -13313 15248 -13310
rect 15227 -13344 15248 -13313
rect 15282 -13344 15341 -13310
rect 15375 -13344 15460 -13310
rect 15512 -13283 15524 -13249
rect 15558 -13283 15570 -13249
rect 15512 -13318 15570 -13283
rect 15605 -13127 16674 -13085
rect 15605 -13161 15622 -13127
rect 15656 -13161 16622 -13127
rect 16656 -13161 16674 -13127
rect 15605 -13229 16674 -13161
rect 15605 -13263 15622 -13229
rect 15656 -13263 16622 -13229
rect 16656 -13263 16674 -13229
rect 15605 -13303 16674 -13263
rect 11236 -13431 11306 -13407
rect 11236 -13465 11430 -13431
rect 11832 -13441 11982 -13371
rect 11101 -13542 11120 -13508
rect 11154 -13542 11171 -13508
rect 11101 -13561 11171 -13542
rect 11264 -13508 11330 -13499
rect 11264 -13542 11280 -13508
rect 11314 -13542 11330 -13508
rect 11264 -13595 11330 -13542
rect 11364 -13508 11430 -13465
rect 11364 -13542 11377 -13508
rect 11411 -13542 11430 -13508
rect 11364 -13561 11430 -13542
rect 11464 -13467 11522 -13450
rect 11464 -13501 11476 -13467
rect 11510 -13501 11522 -13467
rect 11464 -13595 11522 -13501
rect 11648 -13493 11982 -13441
rect 13672 -13363 13735 -13347
rect 13672 -13388 13692 -13363
rect 13672 -13422 13685 -13388
rect 13726 -13397 13735 -13363
rect 13719 -13422 13735 -13397
rect 11648 -13527 11666 -13493
rect 11700 -13527 11930 -13493
rect 11964 -13527 11982 -13493
rect 11648 -13595 11982 -13527
rect 13580 -13467 13638 -13450
rect 13672 -13459 13735 -13422
rect 13769 -13363 15193 -13347
rect 13769 -13397 14119 -13363
rect 14153 -13397 14187 -13363
rect 14221 -13397 14255 -13363
rect 14289 -13397 14323 -13363
rect 14357 -13397 14391 -13363
rect 14425 -13397 14459 -13363
rect 14493 -13397 14527 -13363
rect 14561 -13397 14595 -13363
rect 14629 -13397 14663 -13363
rect 14697 -13397 14731 -13363
rect 14765 -13397 14799 -13363
rect 14833 -13397 14867 -13363
rect 14901 -13397 14935 -13363
rect 14969 -13397 15003 -13363
rect 15037 -13397 15071 -13363
rect 15105 -13397 15139 -13363
rect 15173 -13397 15193 -13363
rect 13580 -13501 13592 -13467
rect 13626 -13501 13638 -13467
rect 13580 -13595 13638 -13501
rect 13672 -13519 13733 -13493
rect 13672 -13553 13690 -13519
rect 13724 -13553 13733 -13519
rect 13672 -13595 13733 -13553
rect 13769 -13506 13819 -13397
rect 13769 -13540 13776 -13506
rect 13810 -13540 13819 -13506
rect 13769 -13559 13819 -13540
rect 13853 -13506 13905 -13490
rect 13853 -13540 13862 -13506
rect 13896 -13540 13905 -13506
rect 13853 -13595 13905 -13540
rect 13941 -13506 13991 -13397
rect 15227 -13405 15460 -13344
rect 15227 -13406 15340 -13405
rect 15227 -13431 15248 -13406
rect 14111 -13440 15248 -13431
rect 15282 -13439 15340 -13406
rect 15374 -13439 15460 -13405
rect 15605 -13373 16124 -13303
rect 15605 -13407 15686 -13373
rect 15720 -13407 15814 -13373
rect 15848 -13407 15942 -13373
rect 15976 -13407 16070 -13373
rect 16104 -13407 16124 -13373
rect 16158 -13371 16178 -13337
rect 16212 -13371 16306 -13337
rect 16340 -13371 16434 -13337
rect 16468 -13371 16562 -13337
rect 16596 -13371 16674 -13337
rect 15282 -13440 15460 -13439
rect 14111 -13465 15460 -13440
rect 16158 -13441 16674 -13371
rect 13941 -13540 13948 -13506
rect 13982 -13540 13991 -13506
rect 13941 -13559 13991 -13540
rect 14025 -13506 14077 -13483
rect 14025 -13540 14034 -13506
rect 14068 -13540 14077 -13506
rect 14025 -13595 14077 -13540
rect 14111 -13506 14163 -13465
rect 14111 -13540 14120 -13506
rect 14154 -13540 14163 -13506
rect 14111 -13556 14163 -13540
rect 14197 -13515 14249 -13499
rect 14197 -13549 14206 -13515
rect 14240 -13549 14249 -13515
rect 14197 -13595 14249 -13549
rect 14283 -13506 14335 -13465
rect 14283 -13540 14292 -13506
rect 14326 -13540 14335 -13506
rect 14283 -13556 14335 -13540
rect 14369 -13515 14421 -13499
rect 14369 -13549 14378 -13515
rect 14412 -13549 14421 -13515
rect 14369 -13595 14421 -13549
rect 14455 -13506 14507 -13465
rect 14455 -13540 14464 -13506
rect 14498 -13540 14507 -13506
rect 14455 -13556 14507 -13540
rect 14541 -13515 14590 -13499
rect 14541 -13549 14550 -13515
rect 14584 -13549 14590 -13515
rect 14541 -13595 14590 -13549
rect 14624 -13506 14679 -13465
rect 14624 -13540 14636 -13506
rect 14670 -13540 14679 -13506
rect 14624 -13556 14679 -13540
rect 14713 -13515 14762 -13499
rect 14713 -13549 14722 -13515
rect 14756 -13549 14762 -13515
rect 14713 -13595 14762 -13549
rect 14796 -13506 14848 -13465
rect 14796 -13540 14807 -13506
rect 14841 -13540 14848 -13506
rect 14796 -13556 14848 -13540
rect 14884 -13515 14934 -13499
rect 14884 -13549 14893 -13515
rect 14927 -13549 14934 -13515
rect 14884 -13595 14934 -13549
rect 14968 -13506 15020 -13465
rect 14968 -13540 14979 -13506
rect 15013 -13540 15020 -13506
rect 14968 -13556 15020 -13540
rect 15056 -13515 15106 -13499
rect 15056 -13549 15065 -13515
rect 15099 -13549 15106 -13515
rect 15056 -13595 15106 -13549
rect 15140 -13506 15192 -13465
rect 15140 -13540 15151 -13506
rect 15185 -13540 15192 -13506
rect 15140 -13556 15192 -13540
rect 15228 -13515 15280 -13499
rect 15228 -13549 15237 -13515
rect 15271 -13549 15280 -13515
rect 15228 -13595 15280 -13549
rect 15314 -13506 15366 -13465
rect 15512 -13467 15570 -13450
rect 15314 -13540 15323 -13506
rect 15357 -13540 15366 -13506
rect 15314 -13556 15366 -13540
rect 15400 -13515 15460 -13499
rect 15400 -13549 15409 -13515
rect 15443 -13549 15460 -13515
rect 15400 -13595 15460 -13549
rect 15512 -13501 15524 -13467
rect 15558 -13501 15570 -13467
rect 15512 -13595 15570 -13501
rect 15605 -13500 16674 -13441
rect 15605 -13534 15622 -13500
rect 15656 -13534 16622 -13500
rect 16656 -13534 16674 -13500
rect 15605 -13595 16674 -13534
rect -2997 -13629 -2968 -13595
rect -2934 -13629 -2876 -13595
rect -2842 -13629 -2784 -13595
rect -2750 -13629 -2692 -13595
rect -2658 -13629 -2600 -13595
rect -2566 -13629 -2508 -13595
rect -2474 -13629 -2416 -13595
rect -2382 -13629 -2324 -13595
rect -2290 -13629 -2232 -13595
rect -2198 -13629 -2140 -13595
rect -2106 -13629 -2048 -13595
rect -2014 -13629 -1956 -13595
rect -1922 -13629 -1864 -13595
rect -1830 -13629 -1772 -13595
rect -1738 -13629 -1680 -13595
rect -1646 -13629 -1588 -13595
rect -1554 -13629 -1496 -13595
rect -1462 -13629 -1404 -13595
rect -1370 -13629 -1312 -13595
rect -1278 -13629 -1220 -13595
rect -1186 -13629 -1128 -13595
rect -1094 -13629 -1036 -13595
rect -1002 -13629 -944 -13595
rect -910 -13629 -852 -13595
rect -818 -13629 -760 -13595
rect -726 -13629 -668 -13595
rect -634 -13629 -576 -13595
rect -542 -13629 -484 -13595
rect -450 -13629 -392 -13595
rect -358 -13629 -300 -13595
rect -266 -13629 -208 -13595
rect -174 -13629 -116 -13595
rect -82 -13629 -24 -13595
rect 10 -13629 68 -13595
rect 102 -13629 160 -13595
rect 194 -13629 252 -13595
rect 286 -13629 344 -13595
rect 378 -13629 436 -13595
rect 470 -13629 528 -13595
rect 562 -13629 620 -13595
rect 654 -13629 712 -13595
rect 746 -13629 804 -13595
rect 838 -13629 896 -13595
rect 930 -13629 988 -13595
rect 1022 -13629 1080 -13595
rect 1114 -13629 1172 -13595
rect 1206 -13629 1264 -13595
rect 1298 -13629 1356 -13595
rect 1390 -13629 1448 -13595
rect 1482 -13629 1540 -13595
rect 1574 -13629 1632 -13595
rect 1666 -13629 1724 -13595
rect 1758 -13629 1816 -13595
rect 1850 -13629 1908 -13595
rect 1942 -13629 2000 -13595
rect 2034 -13629 2092 -13595
rect 2126 -13629 2184 -13595
rect 2218 -13629 2276 -13595
rect 2310 -13629 2368 -13595
rect 2402 -13629 2460 -13595
rect 2494 -13629 2552 -13595
rect 2586 -13629 2644 -13595
rect 2678 -13629 2736 -13595
rect 2770 -13629 2828 -13595
rect 2862 -13629 2920 -13595
rect 2954 -13629 3012 -13595
rect 3046 -13629 3104 -13595
rect 3138 -13629 3196 -13595
rect 3230 -13629 3288 -13595
rect 3322 -13629 3380 -13595
rect 3414 -13629 3472 -13595
rect 3506 -13629 3564 -13595
rect 3598 -13629 3656 -13595
rect 3690 -13629 3748 -13595
rect 3782 -13629 3840 -13595
rect 3874 -13629 3932 -13595
rect 3966 -13629 4024 -13595
rect 4058 -13629 4116 -13595
rect 4150 -13629 4208 -13595
rect 4242 -13629 4300 -13595
rect 4334 -13629 4392 -13595
rect 4426 -13629 4484 -13595
rect 4518 -13629 4576 -13595
rect 4610 -13629 4668 -13595
rect 4702 -13629 4760 -13595
rect 4794 -13629 4852 -13595
rect 4886 -13629 4944 -13595
rect 4978 -13629 5036 -13595
rect 5070 -13629 5128 -13595
rect 5162 -13629 5220 -13595
rect 5254 -13629 5312 -13595
rect 5346 -13629 5404 -13595
rect 5438 -13629 5496 -13595
rect 5530 -13629 5588 -13595
rect 5622 -13629 5680 -13595
rect 5714 -13629 5772 -13595
rect 5806 -13629 5864 -13595
rect 5898 -13629 5956 -13595
rect 5990 -13629 6048 -13595
rect 6082 -13629 6140 -13595
rect 6174 -13629 6232 -13595
rect 6266 -13629 6324 -13595
rect 6358 -13629 6416 -13595
rect 6450 -13629 6508 -13595
rect 6542 -13629 6600 -13595
rect 6634 -13629 6692 -13595
rect 6726 -13629 6784 -13595
rect 6818 -13629 6876 -13595
rect 6910 -13629 6968 -13595
rect 7002 -13629 7060 -13595
rect 7094 -13629 7152 -13595
rect 7186 -13629 7244 -13595
rect 7278 -13629 7336 -13595
rect 7370 -13629 7428 -13595
rect 7462 -13629 7520 -13595
rect 7554 -13629 7612 -13595
rect 7646 -13629 7704 -13595
rect 7738 -13629 7796 -13595
rect 7830 -13629 7888 -13595
rect 7922 -13629 7980 -13595
rect 8014 -13629 8072 -13595
rect 8106 -13629 8164 -13595
rect 8198 -13629 8256 -13595
rect 8290 -13629 8348 -13595
rect 8382 -13629 8440 -13595
rect 8474 -13629 8532 -13595
rect 8566 -13629 8624 -13595
rect 8658 -13629 8716 -13595
rect 8750 -13629 8808 -13595
rect 8842 -13629 8900 -13595
rect 8934 -13629 8992 -13595
rect 9026 -13629 9084 -13595
rect 9118 -13629 9176 -13595
rect 9210 -13629 9268 -13595
rect 9302 -13629 9360 -13595
rect 9394 -13629 9452 -13595
rect 9486 -13629 9544 -13595
rect 9578 -13629 9636 -13595
rect 9670 -13629 9728 -13595
rect 9762 -13629 9820 -13595
rect 9854 -13629 9912 -13595
rect 9946 -13629 10004 -13595
rect 10038 -13629 10096 -13595
rect 10130 -13629 10188 -13595
rect 10222 -13629 10280 -13595
rect 10314 -13629 10372 -13595
rect 10406 -13629 10464 -13595
rect 10498 -13629 10556 -13595
rect 10590 -13629 10648 -13595
rect 10682 -13629 10740 -13595
rect 10774 -13629 10832 -13595
rect 10866 -13629 10924 -13595
rect 10958 -13629 11016 -13595
rect 11050 -13629 11108 -13595
rect 11142 -13629 11200 -13595
rect 11234 -13629 11292 -13595
rect 11326 -13629 11384 -13595
rect 11418 -13629 11476 -13595
rect 11510 -13629 11568 -13595
rect 11602 -13629 11660 -13595
rect 11694 -13629 11752 -13595
rect 11786 -13629 11844 -13595
rect 11878 -13629 11936 -13595
rect 11970 -13629 12028 -13595
rect 12062 -13629 12120 -13595
rect 12154 -13629 12212 -13595
rect 12246 -13629 12304 -13595
rect 12338 -13629 12396 -13595
rect 12430 -13629 12488 -13595
rect 12522 -13629 12580 -13595
rect 12614 -13629 12672 -13595
rect 12706 -13629 12764 -13595
rect 12798 -13629 12856 -13595
rect 12890 -13629 12948 -13595
rect 12982 -13629 13040 -13595
rect 13074 -13629 13132 -13595
rect 13166 -13629 13224 -13595
rect 13258 -13629 13316 -13595
rect 13350 -13629 13408 -13595
rect 13442 -13629 13500 -13595
rect 13534 -13629 13592 -13595
rect 13626 -13629 13684 -13595
rect 13718 -13629 13776 -13595
rect 13810 -13629 13868 -13595
rect 13902 -13629 13960 -13595
rect 13994 -13629 14052 -13595
rect 14086 -13629 14144 -13595
rect 14178 -13629 14236 -13595
rect 14270 -13629 14328 -13595
rect 14362 -13629 14420 -13595
rect 14454 -13629 14512 -13595
rect 14546 -13629 14604 -13595
rect 14638 -13629 14696 -13595
rect 14730 -13629 14788 -13595
rect 14822 -13629 14880 -13595
rect 14914 -13629 14972 -13595
rect 15006 -13629 15064 -13595
rect 15098 -13629 15156 -13595
rect 15190 -13629 15248 -13595
rect 15282 -13629 15340 -13595
rect 15374 -13629 15432 -13595
rect 15466 -13629 15524 -13595
rect 15558 -13629 15616 -13595
rect 15650 -13629 15708 -13595
rect 15742 -13629 15800 -13595
rect 15834 -13629 15892 -13595
rect 15926 -13629 15984 -13595
rect 16018 -13629 16076 -13595
rect 16110 -13629 16168 -13595
rect 16202 -13629 16260 -13595
rect 16294 -13629 16352 -13595
rect 16386 -13629 16444 -13595
rect 16478 -13629 16536 -13595
rect 16570 -13629 16628 -13595
rect 16662 -13629 16691 -13595
rect -2980 -13690 -2278 -13629
rect -2980 -13724 -2962 -13690
rect -2928 -13724 -2330 -13690
rect -2296 -13724 -2278 -13690
rect -2980 -13783 -2278 -13724
rect -2244 -13723 -2186 -13629
rect -2244 -13757 -2232 -13723
rect -2198 -13757 -2186 -13723
rect -2244 -13774 -2186 -13757
rect -1416 -13697 -1082 -13629
rect -1416 -13731 -1398 -13697
rect -1364 -13731 -1134 -13697
rect -1100 -13731 -1082 -13697
rect -2980 -13851 -2902 -13817
rect -2868 -13851 -2799 -13817
rect -2765 -13851 -2696 -13817
rect -2662 -13851 -2642 -13817
rect -2980 -13921 -2642 -13851
rect -2608 -13853 -2278 -13783
rect -2608 -13887 -2588 -13853
rect -2554 -13887 -2489 -13853
rect -2455 -13887 -2390 -13853
rect -2356 -13887 -2278 -13853
rect -1416 -13783 -1082 -13731
rect -1048 -13723 -990 -13629
rect -1048 -13757 -1036 -13723
rect -1002 -13757 -990 -13723
rect -1048 -13774 -990 -13757
rect -956 -13671 -894 -13629
rect -956 -13705 -934 -13671
rect -900 -13705 -894 -13671
rect -956 -13739 -894 -13705
rect -956 -13773 -934 -13739
rect -900 -13773 -894 -13739
rect -1416 -13853 -1266 -13783
rect -956 -13789 -894 -13773
rect -853 -13671 -714 -13663
rect -853 -13705 -766 -13671
rect -732 -13705 -714 -13671
rect -853 -13722 -714 -13705
rect -853 -13756 -848 -13722
rect -814 -13756 -769 -13722
rect -735 -13739 -714 -13722
rect -853 -13773 -766 -13756
rect -732 -13773 -714 -13739
rect -853 -13789 -714 -13773
rect -680 -13723 -622 -13629
rect -680 -13757 -668 -13723
rect -634 -13757 -622 -13723
rect -680 -13774 -622 -13757
rect -588 -13697 -254 -13629
rect -588 -13731 -570 -13697
rect -536 -13731 -306 -13697
rect -272 -13731 -254 -13697
rect -588 -13783 -254 -13731
rect -220 -13723 -162 -13629
rect -32 -13673 27 -13629
rect -32 -13707 -16 -13673
rect 18 -13707 27 -13673
rect -32 -13723 27 -13707
rect 61 -13684 113 -13668
rect 61 -13718 70 -13684
rect 104 -13718 113 -13684
rect -220 -13757 -208 -13723
rect -174 -13757 -162 -13723
rect 61 -13757 113 -13718
rect 147 -13673 199 -13629
rect 147 -13707 156 -13673
rect 190 -13707 199 -13673
rect 147 -13723 199 -13707
rect 233 -13684 284 -13668
rect 233 -13718 242 -13684
rect 276 -13718 284 -13684
rect 233 -13757 284 -13718
rect 318 -13673 378 -13629
rect 318 -13707 328 -13673
rect 362 -13707 378 -13673
rect 318 -13723 378 -13707
rect 516 -13723 574 -13629
rect 516 -13757 528 -13723
rect 562 -13757 574 -13723
rect -220 -13774 -162 -13757
rect -1416 -13887 -1396 -13853
rect -1362 -13887 -1266 -13853
rect -1232 -13851 -1136 -13817
rect -1102 -13851 -1082 -13817
rect -2980 -13961 -2278 -13921
rect -2980 -13995 -2962 -13961
rect -2928 -13995 -2330 -13961
rect -2296 -13995 -2278 -13961
rect -2980 -14063 -2278 -13995
rect -2980 -14097 -2962 -14063
rect -2928 -14097 -2330 -14063
rect -2296 -14097 -2278 -14063
rect -2980 -14139 -2278 -14097
rect -2244 -13941 -2186 -13906
rect -1232 -13921 -1082 -13851
rect -954 -13827 -887 -13823
rect -954 -13861 -937 -13827
rect -903 -13834 -887 -13827
rect -954 -13868 -932 -13861
rect -898 -13868 -887 -13834
rect -954 -13877 -887 -13868
rect -2244 -13975 -2232 -13941
rect -2198 -13975 -2186 -13941
rect -2244 -14034 -2186 -13975
rect -2244 -14068 -2232 -14034
rect -2198 -14068 -2186 -14034
rect -2244 -14139 -2186 -14068
rect -1416 -13961 -1082 -13921
rect -1416 -13995 -1398 -13961
rect -1364 -13995 -1134 -13961
rect -1100 -13995 -1082 -13961
rect -1416 -14063 -1082 -13995
rect -1416 -14097 -1398 -14063
rect -1364 -14097 -1134 -14063
rect -1100 -14097 -1082 -14063
rect -1416 -14139 -1082 -14097
rect -1048 -13941 -990 -13906
rect -853 -13909 -819 -13789
rect -785 -13861 -769 -13827
rect -735 -13835 -718 -13827
rect -785 -13869 -764 -13861
rect -730 -13869 -718 -13835
rect -785 -13877 -718 -13869
rect -588 -13853 -438 -13783
rect -124 -13789 482 -13757
rect 516 -13774 574 -13757
rect 608 -13697 942 -13629
rect 608 -13731 626 -13697
rect 660 -13731 890 -13697
rect 924 -13731 942 -13697
rect -124 -13791 434 -13789
rect -588 -13887 -568 -13853
rect -534 -13887 -438 -13853
rect -404 -13851 -308 -13817
rect -274 -13851 -254 -13817
rect -1048 -13975 -1036 -13941
rect -1002 -13975 -990 -13941
rect -1048 -14034 -990 -13975
rect -1048 -14068 -1036 -14034
rect -1002 -14068 -990 -14034
rect -1048 -14139 -990 -14068
rect -956 -13927 -900 -13911
rect -956 -13961 -934 -13927
rect -956 -13995 -900 -13961
rect -956 -14029 -934 -13995
rect -956 -14063 -900 -14029
rect -956 -14097 -934 -14063
rect -956 -14139 -900 -14097
rect -866 -13927 -800 -13909
rect -866 -13961 -850 -13927
rect -816 -13961 -800 -13927
rect -866 -13995 -800 -13961
rect -866 -14029 -850 -13995
rect -816 -14029 -800 -13995
rect -866 -14063 -800 -14029
rect -866 -14097 -850 -14063
rect -816 -14097 -800 -14063
rect -866 -14105 -800 -14097
rect -766 -13927 -714 -13911
rect -732 -13961 -714 -13927
rect -766 -13995 -714 -13961
rect -732 -14029 -714 -13995
rect -766 -14063 -714 -14029
rect -732 -14097 -714 -14063
rect -766 -14139 -714 -14097
rect -680 -13941 -622 -13906
rect -404 -13921 -254 -13851
rect -124 -13904 -90 -13791
rect 422 -13823 434 -13791
rect 468 -13823 482 -13789
rect -56 -13827 387 -13825
rect -56 -13861 -30 -13827
rect 4 -13861 38 -13827
rect 72 -13861 106 -13827
rect 140 -13861 174 -13827
rect 208 -13861 242 -13827
rect 276 -13861 310 -13827
rect 344 -13861 387 -13827
rect -56 -13870 387 -13861
rect 422 -13904 482 -13823
rect 608 -13783 942 -13731
rect 976 -13723 1034 -13629
rect 1154 -13682 1219 -13663
rect 976 -13757 988 -13723
rect 1022 -13757 1034 -13723
rect 976 -13774 1034 -13757
rect 1068 -13749 1116 -13687
rect 1068 -13783 1076 -13749
rect 1110 -13783 1116 -13749
rect 608 -13853 758 -13783
rect 608 -13887 628 -13853
rect 662 -13887 758 -13853
rect 792 -13851 888 -13817
rect 922 -13851 942 -13817
rect -680 -13975 -668 -13941
rect -634 -13975 -622 -13941
rect -680 -14034 -622 -13975
rect -680 -14068 -668 -14034
rect -634 -14068 -622 -14034
rect -680 -14139 -622 -14068
rect -588 -13961 -254 -13921
rect -588 -13995 -570 -13961
rect -536 -13995 -306 -13961
rect -272 -13995 -254 -13961
rect -588 -14063 -254 -13995
rect -588 -14097 -570 -14063
rect -536 -14097 -306 -14063
rect -272 -14097 -254 -14063
rect -588 -14139 -254 -14097
rect -220 -13941 -162 -13906
rect -124 -13938 482 -13904
rect -220 -13975 -208 -13941
rect -174 -13975 -162 -13941
rect -24 -13961 27 -13938
rect -220 -14034 -162 -13975
rect -220 -14068 -208 -14034
rect -174 -14068 -162 -14034
rect -220 -14139 -162 -14068
rect -128 -13988 -59 -13972
rect -128 -14022 -102 -13988
rect -68 -14022 -59 -13988
rect -128 -14056 -59 -14022
rect -128 -14090 -102 -14056
rect -68 -14090 -59 -14056
rect -128 -14139 -59 -14090
rect -24 -13995 -16 -13961
rect 18 -13995 27 -13961
rect 148 -13961 199 -13938
rect -24 -14049 27 -13995
rect -24 -14083 -16 -14049
rect 18 -14083 27 -14049
rect -24 -14099 27 -14083
rect 61 -13988 113 -13972
rect 61 -14022 70 -13988
rect 104 -14022 113 -13988
rect 61 -14056 113 -14022
rect 61 -14090 70 -14056
rect 104 -14090 113 -14056
rect 61 -14139 113 -14090
rect 148 -13995 156 -13961
rect 190 -13995 199 -13961
rect 319 -13961 371 -13938
rect 148 -14049 199 -13995
rect 148 -14083 156 -14049
rect 190 -14083 199 -14049
rect 148 -14099 199 -14083
rect 233 -13988 285 -13972
rect 233 -14022 242 -13988
rect 276 -14022 285 -13988
rect 233 -14056 285 -14022
rect 233 -14090 242 -14056
rect 276 -14090 285 -14056
rect 233 -14139 285 -14090
rect 319 -13995 328 -13961
rect 362 -13995 371 -13961
rect 516 -13941 574 -13906
rect 792 -13921 942 -13851
rect 1068 -13822 1116 -13783
rect 1068 -13856 1076 -13822
rect 1110 -13827 1116 -13822
rect 1068 -13861 1082 -13856
rect 1068 -13877 1116 -13861
rect 1154 -13716 1169 -13682
rect 1203 -13716 1219 -13682
rect 1154 -13764 1219 -13716
rect 1253 -13680 1310 -13629
rect 1287 -13714 1310 -13680
rect 1253 -13730 1310 -13714
rect 1344 -13723 1402 -13629
rect 1344 -13757 1356 -13723
rect 1390 -13757 1402 -13723
rect 1154 -13828 1310 -13764
rect 1344 -13774 1402 -13757
rect 1436 -13697 1770 -13629
rect 1436 -13731 1454 -13697
rect 1488 -13731 1718 -13697
rect 1752 -13731 1770 -13697
rect 1154 -13862 1171 -13828
rect 1205 -13862 1263 -13828
rect 1297 -13862 1310 -13828
rect 1154 -13870 1310 -13862
rect 1436 -13783 1770 -13731
rect 1804 -13723 1862 -13629
rect 1804 -13757 1816 -13723
rect 1850 -13757 1862 -13723
rect 1804 -13774 1862 -13757
rect 1896 -13697 2230 -13629
rect 1896 -13731 1914 -13697
rect 1948 -13731 2178 -13697
rect 2212 -13731 2230 -13697
rect 1896 -13783 2230 -13731
rect 2264 -13723 2322 -13629
rect 2264 -13757 2276 -13723
rect 2310 -13757 2322 -13723
rect 2264 -13774 2322 -13757
rect 2356 -13682 2422 -13663
rect 2356 -13716 2375 -13682
rect 2409 -13716 2422 -13682
rect 2356 -13759 2422 -13716
rect 2456 -13682 2522 -13629
rect 2456 -13716 2472 -13682
rect 2506 -13716 2522 -13682
rect 2456 -13725 2522 -13716
rect 2615 -13682 2685 -13663
rect 2615 -13716 2632 -13682
rect 2666 -13716 2685 -13682
rect 1436 -13853 1586 -13783
rect 319 -14049 371 -13995
rect 319 -14083 328 -14049
rect 362 -14083 371 -14049
rect 319 -14099 371 -14083
rect 405 -13988 482 -13972
rect 405 -14022 414 -13988
rect 448 -14022 482 -13988
rect 405 -14056 482 -14022
rect 405 -14090 414 -14056
rect 448 -14090 482 -14056
rect 405 -14139 482 -14090
rect 516 -13975 528 -13941
rect 562 -13975 574 -13941
rect 516 -14034 574 -13975
rect 516 -14068 528 -14034
rect 562 -14068 574 -14034
rect 516 -14139 574 -14068
rect 608 -13961 942 -13921
rect 608 -13995 626 -13961
rect 660 -13995 890 -13961
rect 924 -13995 942 -13961
rect 608 -14063 942 -13995
rect 608 -14097 626 -14063
rect 660 -14097 890 -14063
rect 924 -14097 942 -14063
rect 608 -14139 942 -14097
rect 976 -13941 1034 -13906
rect 976 -13975 988 -13941
rect 1022 -13975 1034 -13941
rect 976 -14034 1034 -13975
rect 976 -14068 988 -14034
rect 1022 -14068 1034 -14034
rect 976 -14139 1034 -14068
rect 1068 -13961 1120 -13945
rect 1068 -13995 1086 -13961
rect 1068 -14063 1120 -13995
rect 1068 -14097 1086 -14063
rect 1068 -14139 1120 -14097
rect 1154 -13961 1220 -13870
rect 1436 -13887 1456 -13853
rect 1490 -13887 1586 -13853
rect 1620 -13851 1716 -13817
rect 1750 -13851 1770 -13817
rect 1344 -13941 1402 -13906
rect 1620 -13921 1770 -13851
rect 1896 -13853 2046 -13783
rect 2356 -13793 2550 -13759
rect 2480 -13817 2550 -13793
rect 1896 -13887 1916 -13853
rect 1950 -13887 2046 -13853
rect 2080 -13851 2176 -13817
rect 2210 -13851 2230 -13817
rect 2480 -13827 2566 -13817
rect 1154 -13995 1170 -13961
rect 1204 -13995 1220 -13961
rect 1154 -14063 1220 -13995
rect 1154 -14097 1170 -14063
rect 1204 -14097 1220 -14063
rect 1154 -14105 1220 -14097
rect 1254 -13961 1310 -13945
rect 1288 -13995 1310 -13961
rect 1254 -14063 1310 -13995
rect 1288 -14097 1310 -14063
rect 1254 -14139 1310 -14097
rect 1344 -13975 1356 -13941
rect 1390 -13975 1402 -13941
rect 1344 -14034 1402 -13975
rect 1344 -14068 1356 -14034
rect 1390 -14068 1402 -14034
rect 1344 -14139 1402 -14068
rect 1436 -13961 1770 -13921
rect 1436 -13995 1454 -13961
rect 1488 -13995 1718 -13961
rect 1752 -13995 1770 -13961
rect 1436 -14063 1770 -13995
rect 1436 -14097 1454 -14063
rect 1488 -14097 1718 -14063
rect 1752 -14097 1770 -14063
rect 1436 -14139 1770 -14097
rect 1804 -13941 1862 -13906
rect 2080 -13921 2230 -13851
rect 2356 -13833 2396 -13827
rect 2356 -13867 2369 -13833
rect 2430 -13861 2446 -13827
rect 2403 -13867 2446 -13861
rect 2356 -13870 2446 -13867
rect 2480 -13861 2516 -13827
rect 2550 -13861 2566 -13827
rect 2480 -13875 2566 -13861
rect 2615 -13826 2685 -13716
rect 2737 -13682 2787 -13663
rect 2771 -13716 2787 -13682
rect 2737 -13758 2787 -13716
rect 2877 -13682 2943 -13629
rect 2877 -13716 2893 -13682
rect 2927 -13716 2943 -13682
rect 2877 -13732 2943 -13716
rect 2977 -13682 3058 -13663
rect 2977 -13716 2991 -13682
rect 3025 -13716 3058 -13682
rect 2977 -13740 3058 -13716
rect 2737 -13792 2855 -13758
rect 2821 -13811 2855 -13792
rect 2615 -13827 2787 -13826
rect 2615 -13861 2737 -13827
rect 2771 -13861 2787 -13827
rect 2480 -13904 2550 -13875
rect 1804 -13975 1816 -13941
rect 1850 -13975 1862 -13941
rect 1804 -14034 1862 -13975
rect 1804 -14068 1816 -14034
rect 1850 -14068 1862 -14034
rect 1804 -14139 1862 -14068
rect 1896 -13961 2230 -13921
rect 1896 -13995 1914 -13961
rect 1948 -13995 2178 -13961
rect 2212 -13995 2230 -13961
rect 1896 -14063 2230 -13995
rect 1896 -14097 1914 -14063
rect 1948 -14097 2178 -14063
rect 2212 -14097 2230 -14063
rect 1896 -14139 2230 -14097
rect 2264 -13941 2322 -13906
rect 2264 -13975 2276 -13941
rect 2310 -13975 2322 -13941
rect 2264 -14034 2322 -13975
rect 2264 -14068 2276 -14034
rect 2310 -14068 2322 -14034
rect 2264 -14139 2322 -14068
rect 2356 -13938 2550 -13904
rect 2615 -13876 2787 -13861
rect 2821 -13827 2974 -13811
rect 2821 -13861 2937 -13827
rect 2971 -13861 2974 -13827
rect 2356 -13988 2425 -13938
rect 2356 -14022 2375 -13988
rect 2409 -14022 2425 -13988
rect 2356 -14056 2425 -14022
rect 2356 -14090 2375 -14056
rect 2409 -14090 2425 -14056
rect 2356 -14105 2425 -14090
rect 2459 -13988 2525 -13972
rect 2459 -14022 2475 -13988
rect 2509 -14022 2525 -13988
rect 2459 -14056 2525 -14022
rect 2459 -14090 2475 -14056
rect 2509 -14090 2525 -14056
rect 2459 -14139 2525 -14090
rect 2615 -13988 2685 -13876
rect 2821 -13877 2974 -13861
rect 3008 -13832 3058 -13740
rect 3092 -13723 3150 -13629
rect 3092 -13757 3104 -13723
rect 3138 -13757 3150 -13723
rect 3092 -13774 3150 -13757
rect 3184 -13697 3518 -13629
rect 3184 -13731 3202 -13697
rect 3236 -13731 3466 -13697
rect 3500 -13731 3518 -13697
rect 3008 -13866 3015 -13832
rect 3049 -13866 3058 -13832
rect 2821 -13911 2855 -13877
rect 2615 -14022 2633 -13988
rect 2667 -14022 2685 -13988
rect 2615 -14056 2685 -14022
rect 2615 -14090 2633 -14056
rect 2667 -14090 2685 -14056
rect 2615 -14105 2685 -14090
rect 2737 -13945 2855 -13911
rect 2737 -13987 2787 -13945
rect 3008 -13950 3058 -13866
rect 3184 -13783 3518 -13731
rect 3552 -13723 3610 -13629
rect 3552 -13757 3564 -13723
rect 3598 -13757 3610 -13723
rect 3552 -13774 3610 -13757
rect 4380 -13690 5449 -13629
rect 4380 -13724 4398 -13690
rect 4432 -13724 5398 -13690
rect 5432 -13724 5449 -13690
rect 4380 -13783 5449 -13724
rect 6312 -13723 6370 -13629
rect 6312 -13757 6324 -13723
rect 6358 -13757 6370 -13723
rect 6312 -13774 6370 -13757
rect 6404 -13697 6738 -13629
rect 6404 -13731 6422 -13697
rect 6456 -13731 6686 -13697
rect 6720 -13731 6738 -13697
rect 6404 -13783 6738 -13731
rect 6772 -13723 6830 -13629
rect 6772 -13757 6784 -13723
rect 6818 -13757 6830 -13723
rect 6772 -13774 6830 -13757
rect 6864 -13682 6930 -13663
rect 6864 -13716 6883 -13682
rect 6917 -13716 6930 -13682
rect 6864 -13759 6930 -13716
rect 6964 -13682 7030 -13629
rect 6964 -13716 6980 -13682
rect 7014 -13716 7030 -13682
rect 6964 -13725 7030 -13716
rect 7123 -13682 7193 -13663
rect 7123 -13716 7140 -13682
rect 7174 -13716 7193 -13682
rect 3184 -13853 3334 -13783
rect 3184 -13887 3204 -13853
rect 3238 -13887 3334 -13853
rect 3368 -13851 3464 -13817
rect 3498 -13851 3518 -13817
rect 2771 -14021 2787 -13987
rect 2737 -14055 2787 -14021
rect 2771 -14089 2787 -14055
rect 2737 -14105 2787 -14089
rect 2877 -13988 2943 -13979
rect 2877 -14022 2893 -13988
rect 2927 -14022 2943 -13988
rect 2877 -14056 2943 -14022
rect 2877 -14090 2893 -14056
rect 2927 -14090 2943 -14056
rect 2877 -14139 2943 -14090
rect 2977 -13987 3058 -13950
rect 2977 -14021 2991 -13987
rect 3025 -14021 3058 -13987
rect 2977 -14055 3058 -14021
rect 2977 -14089 2991 -14055
rect 3025 -14089 3058 -14055
rect 2977 -14105 3058 -14089
rect 3092 -13941 3150 -13906
rect 3368 -13921 3518 -13851
rect 4380 -13853 4896 -13783
rect 4380 -13887 4458 -13853
rect 4492 -13887 4586 -13853
rect 4620 -13887 4714 -13853
rect 4748 -13887 4842 -13853
rect 4876 -13887 4896 -13853
rect 4930 -13851 4950 -13817
rect 4984 -13851 5078 -13817
rect 5112 -13851 5206 -13817
rect 5240 -13851 5334 -13817
rect 5368 -13851 5449 -13817
rect 3092 -13975 3104 -13941
rect 3138 -13975 3150 -13941
rect 3092 -14034 3150 -13975
rect 3092 -14068 3104 -14034
rect 3138 -14068 3150 -14034
rect 3092 -14139 3150 -14068
rect 3184 -13961 3518 -13921
rect 3184 -13995 3202 -13961
rect 3236 -13995 3466 -13961
rect 3500 -13995 3518 -13961
rect 3184 -14063 3518 -13995
rect 3184 -14097 3202 -14063
rect 3236 -14097 3466 -14063
rect 3500 -14097 3518 -14063
rect 3184 -14139 3518 -14097
rect 3552 -13941 3610 -13906
rect 4930 -13921 5449 -13851
rect 6404 -13853 6554 -13783
rect 6864 -13793 7058 -13759
rect 6988 -13817 7058 -13793
rect 6404 -13887 6424 -13853
rect 6458 -13887 6554 -13853
rect 6588 -13851 6684 -13817
rect 6718 -13851 6738 -13817
rect 6988 -13827 7074 -13817
rect 3552 -13975 3564 -13941
rect 3598 -13975 3610 -13941
rect 3552 -14034 3610 -13975
rect 3552 -14068 3564 -14034
rect 3598 -14068 3610 -14034
rect 3552 -14139 3610 -14068
rect 4380 -13961 5449 -13921
rect 4380 -13995 4398 -13961
rect 4432 -13995 5398 -13961
rect 5432 -13995 5449 -13961
rect 4380 -14063 5449 -13995
rect 4380 -14097 4398 -14063
rect 4432 -14097 5398 -14063
rect 5432 -14097 5449 -14063
rect 4380 -14139 5449 -14097
rect 6312 -13941 6370 -13906
rect 6588 -13921 6738 -13851
rect 6864 -13832 6904 -13827
rect 6864 -13866 6876 -13832
rect 6938 -13861 6954 -13827
rect 6910 -13866 6954 -13861
rect 6864 -13870 6954 -13866
rect 6988 -13861 7024 -13827
rect 7058 -13861 7074 -13827
rect 6988 -13875 7074 -13861
rect 7123 -13826 7193 -13716
rect 7245 -13682 7295 -13663
rect 7279 -13716 7295 -13682
rect 7245 -13758 7295 -13716
rect 7385 -13682 7451 -13629
rect 7385 -13716 7401 -13682
rect 7435 -13716 7451 -13682
rect 7385 -13732 7451 -13716
rect 7485 -13682 7566 -13663
rect 7485 -13716 7499 -13682
rect 7533 -13716 7566 -13682
rect 7485 -13740 7566 -13716
rect 7245 -13792 7363 -13758
rect 7329 -13811 7363 -13792
rect 7123 -13827 7295 -13826
rect 7123 -13861 7245 -13827
rect 7279 -13861 7295 -13827
rect 6988 -13904 7058 -13875
rect 6312 -13975 6324 -13941
rect 6358 -13975 6370 -13941
rect 6312 -14034 6370 -13975
rect 6312 -14068 6324 -14034
rect 6358 -14068 6370 -14034
rect 6312 -14139 6370 -14068
rect 6404 -13961 6738 -13921
rect 6404 -13995 6422 -13961
rect 6456 -13995 6686 -13961
rect 6720 -13995 6738 -13961
rect 6404 -14063 6738 -13995
rect 6404 -14097 6422 -14063
rect 6456 -14097 6686 -14063
rect 6720 -14097 6738 -14063
rect 6404 -14139 6738 -14097
rect 6772 -13941 6830 -13906
rect 6772 -13975 6784 -13941
rect 6818 -13975 6830 -13941
rect 6772 -14034 6830 -13975
rect 6772 -14068 6784 -14034
rect 6818 -14068 6830 -14034
rect 6772 -14139 6830 -14068
rect 6864 -13938 7058 -13904
rect 7123 -13876 7295 -13861
rect 7329 -13827 7482 -13811
rect 7329 -13861 7445 -13827
rect 7479 -13861 7482 -13827
rect 6864 -13988 6933 -13938
rect 6864 -14022 6883 -13988
rect 6917 -14022 6933 -13988
rect 6864 -14056 6933 -14022
rect 6864 -14090 6883 -14056
rect 6917 -14090 6933 -14056
rect 6864 -14105 6933 -14090
rect 6967 -13988 7033 -13972
rect 6967 -14022 6983 -13988
rect 7017 -14022 7033 -13988
rect 6967 -14056 7033 -14022
rect 6967 -14090 6983 -14056
rect 7017 -14090 7033 -14056
rect 6967 -14139 7033 -14090
rect 7123 -13988 7193 -13876
rect 7329 -13877 7482 -13861
rect 7516 -13832 7566 -13740
rect 7600 -13723 7658 -13629
rect 7600 -13757 7612 -13723
rect 7646 -13757 7658 -13723
rect 7600 -13774 7658 -13757
rect 7692 -13697 8026 -13629
rect 7692 -13731 7710 -13697
rect 7744 -13731 7974 -13697
rect 8008 -13731 8026 -13697
rect 7516 -13866 7522 -13832
rect 7556 -13866 7566 -13832
rect 7329 -13911 7363 -13877
rect 7123 -14022 7141 -13988
rect 7175 -14022 7193 -13988
rect 7123 -14056 7193 -14022
rect 7123 -14090 7141 -14056
rect 7175 -14090 7193 -14056
rect 7123 -14105 7193 -14090
rect 7245 -13945 7363 -13911
rect 7245 -13987 7295 -13945
rect 7516 -13950 7566 -13866
rect 7692 -13783 8026 -13731
rect 8060 -13723 8118 -13629
rect 8060 -13757 8072 -13723
rect 8106 -13757 8118 -13723
rect 8060 -13774 8118 -13757
rect 8152 -13682 8218 -13663
rect 8152 -13716 8171 -13682
rect 8205 -13716 8218 -13682
rect 8152 -13759 8218 -13716
rect 8252 -13682 8318 -13629
rect 8252 -13716 8268 -13682
rect 8302 -13716 8318 -13682
rect 8252 -13725 8318 -13716
rect 8411 -13682 8481 -13663
rect 8411 -13716 8428 -13682
rect 8462 -13716 8481 -13682
rect 7692 -13853 7842 -13783
rect 8152 -13793 8346 -13759
rect 8276 -13817 8346 -13793
rect 7692 -13887 7712 -13853
rect 7746 -13887 7842 -13853
rect 7876 -13851 7972 -13817
rect 8006 -13851 8026 -13817
rect 8276 -13827 8362 -13817
rect 7279 -14021 7295 -13987
rect 7245 -14055 7295 -14021
rect 7279 -14089 7295 -14055
rect 7245 -14105 7295 -14089
rect 7385 -13988 7451 -13979
rect 7385 -14022 7401 -13988
rect 7435 -14022 7451 -13988
rect 7385 -14056 7451 -14022
rect 7385 -14090 7401 -14056
rect 7435 -14090 7451 -14056
rect 7385 -14139 7451 -14090
rect 7485 -13987 7566 -13950
rect 7485 -14021 7499 -13987
rect 7533 -14021 7566 -13987
rect 7485 -14055 7566 -14021
rect 7485 -14089 7499 -14055
rect 7533 -14089 7566 -14055
rect 7485 -14105 7566 -14089
rect 7600 -13941 7658 -13906
rect 7876 -13921 8026 -13851
rect 8152 -13831 8192 -13827
rect 8152 -13865 8164 -13831
rect 8226 -13861 8242 -13827
rect 8198 -13865 8242 -13861
rect 8152 -13870 8242 -13865
rect 8276 -13861 8312 -13827
rect 8346 -13861 8362 -13827
rect 8276 -13875 8362 -13861
rect 8411 -13826 8481 -13716
rect 8533 -13682 8583 -13663
rect 8567 -13716 8583 -13682
rect 8533 -13758 8583 -13716
rect 8673 -13682 8739 -13629
rect 8673 -13716 8689 -13682
rect 8723 -13716 8739 -13682
rect 8673 -13732 8739 -13716
rect 8773 -13682 8854 -13663
rect 8773 -13716 8787 -13682
rect 8821 -13716 8854 -13682
rect 8773 -13740 8854 -13716
rect 8533 -13792 8651 -13758
rect 8617 -13811 8651 -13792
rect 8411 -13827 8583 -13826
rect 8411 -13861 8533 -13827
rect 8567 -13861 8583 -13827
rect 8276 -13904 8346 -13875
rect 7600 -13975 7612 -13941
rect 7646 -13975 7658 -13941
rect 7600 -14034 7658 -13975
rect 7600 -14068 7612 -14034
rect 7646 -14068 7658 -14034
rect 7600 -14139 7658 -14068
rect 7692 -13961 8026 -13921
rect 7692 -13995 7710 -13961
rect 7744 -13995 7974 -13961
rect 8008 -13995 8026 -13961
rect 7692 -14063 8026 -13995
rect 7692 -14097 7710 -14063
rect 7744 -14097 7974 -14063
rect 8008 -14097 8026 -14063
rect 7692 -14139 8026 -14097
rect 8060 -13941 8118 -13906
rect 8060 -13975 8072 -13941
rect 8106 -13975 8118 -13941
rect 8060 -14034 8118 -13975
rect 8060 -14068 8072 -14034
rect 8106 -14068 8118 -14034
rect 8060 -14139 8118 -14068
rect 8152 -13938 8346 -13904
rect 8411 -13876 8583 -13861
rect 8617 -13827 8770 -13811
rect 8617 -13861 8733 -13827
rect 8767 -13861 8770 -13827
rect 8152 -13988 8221 -13938
rect 8152 -14022 8171 -13988
rect 8205 -14022 8221 -13988
rect 8152 -14056 8221 -14022
rect 8152 -14090 8171 -14056
rect 8205 -14090 8221 -14056
rect 8152 -14105 8221 -14090
rect 8255 -13988 8321 -13972
rect 8255 -14022 8271 -13988
rect 8305 -14022 8321 -13988
rect 8255 -14056 8321 -14022
rect 8255 -14090 8271 -14056
rect 8305 -14090 8321 -14056
rect 8255 -14139 8321 -14090
rect 8411 -13988 8481 -13876
rect 8617 -13877 8770 -13861
rect 8804 -13833 8854 -13740
rect 8888 -13723 8946 -13629
rect 8888 -13757 8900 -13723
rect 8934 -13757 8946 -13723
rect 8888 -13774 8946 -13757
rect 8980 -13697 9314 -13629
rect 8980 -13731 8998 -13697
rect 9032 -13731 9262 -13697
rect 9296 -13731 9314 -13697
rect 8804 -13867 8811 -13833
rect 8845 -13867 8854 -13833
rect 8617 -13911 8651 -13877
rect 8411 -14022 8429 -13988
rect 8463 -14022 8481 -13988
rect 8411 -14056 8481 -14022
rect 8411 -14090 8429 -14056
rect 8463 -14090 8481 -14056
rect 8411 -14105 8481 -14090
rect 8533 -13945 8651 -13911
rect 8533 -13987 8583 -13945
rect 8804 -13950 8854 -13867
rect 8980 -13783 9314 -13731
rect 9348 -13723 9406 -13629
rect 9348 -13757 9360 -13723
rect 9394 -13757 9406 -13723
rect 9348 -13774 9406 -13757
rect 9440 -13682 9506 -13663
rect 9440 -13716 9459 -13682
rect 9493 -13716 9506 -13682
rect 9440 -13759 9506 -13716
rect 9540 -13682 9606 -13629
rect 9540 -13716 9556 -13682
rect 9590 -13716 9606 -13682
rect 9540 -13725 9606 -13716
rect 9699 -13682 9769 -13663
rect 9699 -13716 9716 -13682
rect 9750 -13716 9769 -13682
rect 8980 -13853 9130 -13783
rect 9440 -13793 9634 -13759
rect 9564 -13817 9634 -13793
rect 8980 -13887 9000 -13853
rect 9034 -13887 9130 -13853
rect 9164 -13851 9260 -13817
rect 9294 -13851 9314 -13817
rect 9564 -13827 9650 -13817
rect 8567 -14021 8583 -13987
rect 8533 -14055 8583 -14021
rect 8567 -14089 8583 -14055
rect 8533 -14105 8583 -14089
rect 8673 -13988 8739 -13979
rect 8673 -14022 8689 -13988
rect 8723 -14022 8739 -13988
rect 8673 -14056 8739 -14022
rect 8673 -14090 8689 -14056
rect 8723 -14090 8739 -14056
rect 8673 -14139 8739 -14090
rect 8773 -13987 8854 -13950
rect 8773 -14021 8787 -13987
rect 8821 -14021 8854 -13987
rect 8773 -14055 8854 -14021
rect 8773 -14089 8787 -14055
rect 8821 -14089 8854 -14055
rect 8773 -14105 8854 -14089
rect 8888 -13941 8946 -13906
rect 9164 -13921 9314 -13851
rect 9440 -13833 9480 -13827
rect 9440 -13867 9453 -13833
rect 9514 -13861 9530 -13827
rect 9487 -13867 9530 -13861
rect 9440 -13870 9530 -13867
rect 9564 -13861 9600 -13827
rect 9634 -13861 9650 -13827
rect 9564 -13875 9650 -13861
rect 9699 -13826 9769 -13716
rect 9821 -13682 9871 -13663
rect 9855 -13716 9871 -13682
rect 9821 -13758 9871 -13716
rect 9961 -13682 10027 -13629
rect 9961 -13716 9977 -13682
rect 10011 -13716 10027 -13682
rect 9961 -13732 10027 -13716
rect 10061 -13682 10142 -13663
rect 10061 -13716 10075 -13682
rect 10109 -13716 10142 -13682
rect 10061 -13740 10142 -13716
rect 9821 -13792 9939 -13758
rect 9905 -13811 9939 -13792
rect 9699 -13827 9871 -13826
rect 9699 -13861 9821 -13827
rect 9855 -13861 9871 -13827
rect 9564 -13904 9634 -13875
rect 8888 -13975 8900 -13941
rect 8934 -13975 8946 -13941
rect 8888 -14034 8946 -13975
rect 8888 -14068 8900 -14034
rect 8934 -14068 8946 -14034
rect 8888 -14139 8946 -14068
rect 8980 -13961 9314 -13921
rect 8980 -13995 8998 -13961
rect 9032 -13995 9262 -13961
rect 9296 -13995 9314 -13961
rect 8980 -14063 9314 -13995
rect 8980 -14097 8998 -14063
rect 9032 -14097 9262 -14063
rect 9296 -14097 9314 -14063
rect 8980 -14139 9314 -14097
rect 9348 -13941 9406 -13906
rect 9348 -13975 9360 -13941
rect 9394 -13975 9406 -13941
rect 9348 -14034 9406 -13975
rect 9348 -14068 9360 -14034
rect 9394 -14068 9406 -14034
rect 9348 -14139 9406 -14068
rect 9440 -13938 9634 -13904
rect 9699 -13876 9871 -13861
rect 9905 -13827 10058 -13811
rect 9905 -13861 10021 -13827
rect 10055 -13861 10058 -13827
rect 9440 -13988 9509 -13938
rect 9440 -14022 9459 -13988
rect 9493 -14022 9509 -13988
rect 9440 -14056 9509 -14022
rect 9440 -14090 9459 -14056
rect 9493 -14090 9509 -14056
rect 9440 -14105 9509 -14090
rect 9543 -13988 9609 -13972
rect 9543 -14022 9559 -13988
rect 9593 -14022 9609 -13988
rect 9543 -14056 9609 -14022
rect 9543 -14090 9559 -14056
rect 9593 -14090 9609 -14056
rect 9543 -14139 9609 -14090
rect 9699 -13988 9769 -13876
rect 9905 -13877 10058 -13861
rect 10092 -13834 10142 -13740
rect 10176 -13723 10234 -13629
rect 10176 -13757 10188 -13723
rect 10222 -13757 10234 -13723
rect 10176 -13774 10234 -13757
rect 10268 -13697 10602 -13629
rect 10268 -13731 10286 -13697
rect 10320 -13731 10550 -13697
rect 10584 -13731 10602 -13697
rect 10092 -13868 10099 -13834
rect 10133 -13868 10142 -13834
rect 9905 -13911 9939 -13877
rect 9699 -14022 9717 -13988
rect 9751 -14022 9769 -13988
rect 9699 -14056 9769 -14022
rect 9699 -14090 9717 -14056
rect 9751 -14090 9769 -14056
rect 9699 -14105 9769 -14090
rect 9821 -13945 9939 -13911
rect 9821 -13987 9871 -13945
rect 10092 -13950 10142 -13868
rect 10268 -13783 10602 -13731
rect 10636 -13723 10694 -13629
rect 10636 -13757 10648 -13723
rect 10682 -13757 10694 -13723
rect 10636 -13774 10694 -13757
rect 10729 -13671 10796 -13663
rect 10729 -13705 10746 -13671
rect 10780 -13705 10796 -13671
rect 10729 -13739 10796 -13705
rect 10830 -13671 10864 -13629
rect 10830 -13721 10864 -13705
rect 10898 -13671 10964 -13663
rect 10898 -13705 10914 -13671
rect 10948 -13705 10964 -13671
rect 10729 -13773 10746 -13739
rect 10780 -13755 10796 -13739
rect 10898 -13739 10964 -13705
rect 10998 -13671 11032 -13629
rect 10998 -13721 11032 -13705
rect 11066 -13671 11468 -13663
rect 11066 -13705 11082 -13671
rect 11116 -13705 11250 -13671
rect 11284 -13705 11418 -13671
rect 11452 -13705 11468 -13671
rect 10898 -13755 10914 -13739
rect 10780 -13773 10914 -13755
rect 10948 -13755 10964 -13739
rect 11066 -13739 11116 -13705
rect 11418 -13739 11468 -13705
rect 11066 -13755 11082 -13739
rect 10948 -13773 11082 -13755
rect 10268 -13853 10418 -13783
rect 10729 -13793 11116 -13773
rect 11150 -13773 11166 -13739
rect 11200 -13773 11334 -13739
rect 11368 -13773 11384 -13739
rect 11452 -13773 11468 -13739
rect 10268 -13887 10288 -13853
rect 10322 -13887 10418 -13853
rect 10452 -13851 10548 -13817
rect 10582 -13851 10602 -13817
rect 11150 -13827 11200 -13773
rect 11418 -13789 11468 -13773
rect 11556 -13723 11614 -13629
rect 11556 -13757 11568 -13723
rect 11602 -13757 11614 -13723
rect 11556 -13774 11614 -13757
rect 11648 -13697 11982 -13629
rect 11648 -13731 11666 -13697
rect 11700 -13731 11930 -13697
rect 11964 -13731 11982 -13697
rect 11648 -13783 11982 -13731
rect 13488 -13723 13546 -13629
rect 13488 -13757 13500 -13723
rect 13534 -13757 13546 -13723
rect 13488 -13774 13546 -13757
rect 13580 -13690 14649 -13629
rect 13580 -13724 13598 -13690
rect 13632 -13724 14598 -13690
rect 14632 -13724 14649 -13690
rect 13580 -13783 14649 -13724
rect 14684 -13723 14742 -13629
rect 14684 -13757 14696 -13723
rect 14730 -13757 14742 -13723
rect 14684 -13774 14742 -13757
rect 14776 -13690 15845 -13629
rect 14776 -13724 14794 -13690
rect 14828 -13724 15794 -13690
rect 15828 -13724 15845 -13690
rect 14776 -13783 15845 -13724
rect 15880 -13723 15938 -13629
rect 15880 -13757 15892 -13723
rect 15926 -13757 15938 -13723
rect 15880 -13774 15938 -13757
rect 15972 -13690 16674 -13629
rect 15972 -13724 15990 -13690
rect 16024 -13724 16622 -13690
rect 16656 -13724 16674 -13690
rect 15972 -13783 16674 -13724
rect 9855 -14021 9871 -13987
rect 9821 -14055 9871 -14021
rect 9855 -14089 9871 -14055
rect 9821 -14105 9871 -14089
rect 9961 -13988 10027 -13979
rect 9961 -14022 9977 -13988
rect 10011 -14022 10027 -13988
rect 9961 -14056 10027 -14022
rect 9961 -14090 9977 -14056
rect 10011 -14090 10027 -14056
rect 9961 -14139 10027 -14090
rect 10061 -13987 10142 -13950
rect 10061 -14021 10075 -13987
rect 10109 -14021 10142 -13987
rect 10061 -14055 10142 -14021
rect 10061 -14089 10075 -14055
rect 10109 -14089 10142 -14055
rect 10061 -14105 10142 -14089
rect 10176 -13941 10234 -13906
rect 10452 -13921 10602 -13851
rect 10733 -13833 10749 -13827
rect 10733 -13867 10741 -13833
rect 10783 -13861 10830 -13827
rect 10864 -13833 10914 -13827
rect 10948 -13832 10998 -13827
rect 11032 -13832 11057 -13827
rect 10866 -13861 10914 -13833
rect 10959 -13861 10998 -13832
rect 10775 -13867 10832 -13861
rect 10866 -13866 10925 -13861
rect 10959 -13866 11017 -13861
rect 11051 -13866 11057 -13832
rect 10866 -13867 11057 -13866
rect 10733 -13877 11057 -13867
rect 11093 -13866 11200 -13827
rect 11093 -13900 11129 -13866
rect 11163 -13900 11200 -13866
rect 11234 -13869 11250 -13827
rect 11284 -13861 11334 -13827
rect 11368 -13835 11522 -13827
rect 11284 -13869 11344 -13861
rect 11378 -13869 11522 -13835
rect 11234 -13877 11522 -13869
rect 11648 -13853 11798 -13783
rect 11648 -13887 11668 -13853
rect 11702 -13887 11798 -13853
rect 11832 -13851 11928 -13817
rect 11962 -13851 11982 -13817
rect 10176 -13975 10188 -13941
rect 10222 -13975 10234 -13941
rect 10176 -14034 10234 -13975
rect 10176 -14068 10188 -14034
rect 10222 -14068 10234 -14034
rect 10176 -14139 10234 -14068
rect 10268 -13961 10602 -13921
rect 10268 -13995 10286 -13961
rect 10320 -13995 10550 -13961
rect 10584 -13995 10602 -13961
rect 10268 -14063 10602 -13995
rect 10268 -14097 10286 -14063
rect 10320 -14097 10550 -14063
rect 10584 -14097 10602 -14063
rect 10268 -14139 10602 -14097
rect 10636 -13941 10694 -13906
rect 11093 -13911 11200 -13900
rect 10636 -13975 10648 -13941
rect 10682 -13975 10694 -13941
rect 10636 -14034 10694 -13975
rect 10636 -14068 10648 -14034
rect 10682 -14068 10694 -14034
rect 10636 -14139 10694 -14068
rect 10729 -13927 10780 -13911
rect 10729 -13961 10746 -13927
rect 10729 -13995 10780 -13961
rect 10729 -14029 10746 -13995
rect 10729 -14063 10780 -14029
rect 10729 -14097 10746 -14063
rect 10729 -14139 10780 -14097
rect 10814 -13927 11384 -13911
rect 10814 -13961 10830 -13927
rect 10864 -13945 10998 -13927
rect 10864 -13961 10880 -13945
rect 10814 -13995 10880 -13961
rect 10982 -13961 10998 -13945
rect 11032 -13945 11166 -13927
rect 11032 -13961 11048 -13945
rect 10814 -14029 10830 -13995
rect 10864 -14029 10880 -13995
rect 10814 -14063 10880 -14029
rect 10814 -14097 10830 -14063
rect 10864 -14097 10880 -14063
rect 10814 -14105 10880 -14097
rect 10914 -13995 10948 -13979
rect 10914 -14063 10948 -14029
rect 10914 -14139 10948 -14097
rect 10982 -13995 11048 -13961
rect 11150 -13961 11166 -13945
rect 11200 -13945 11334 -13927
rect 11200 -13961 11216 -13945
rect 10982 -14029 10998 -13995
rect 11032 -14029 11048 -13995
rect 10982 -14063 11048 -14029
rect 10982 -14097 10998 -14063
rect 11032 -14097 11048 -14063
rect 10982 -14105 11048 -14097
rect 11082 -13995 11116 -13979
rect 11082 -14063 11116 -14029
rect 11082 -14139 11116 -14097
rect 11150 -13995 11216 -13961
rect 11318 -13961 11334 -13945
rect 11368 -13961 11384 -13927
rect 11150 -14029 11166 -13995
rect 11200 -14029 11216 -13995
rect 11150 -14063 11216 -14029
rect 11150 -14097 11166 -14063
rect 11200 -14097 11216 -14063
rect 11150 -14105 11216 -14097
rect 11250 -13995 11284 -13979
rect 11250 -14063 11284 -14029
rect 11250 -14139 11284 -14097
rect 11318 -13995 11384 -13961
rect 11556 -13941 11614 -13906
rect 11832 -13921 11982 -13851
rect 13580 -13853 14096 -13783
rect 13580 -13887 13658 -13853
rect 13692 -13887 13786 -13853
rect 13820 -13887 13914 -13853
rect 13948 -13887 14042 -13853
rect 14076 -13887 14096 -13853
rect 14130 -13851 14150 -13817
rect 14184 -13851 14278 -13817
rect 14312 -13851 14406 -13817
rect 14440 -13851 14534 -13817
rect 14568 -13851 14649 -13817
rect 11556 -13975 11568 -13941
rect 11602 -13975 11614 -13941
rect 11318 -14029 11334 -13995
rect 11368 -14029 11384 -13995
rect 11318 -14063 11384 -14029
rect 11318 -14097 11334 -14063
rect 11368 -14097 11384 -14063
rect 11318 -14105 11384 -14097
rect 11418 -13995 11468 -13979
rect 11452 -14029 11468 -13995
rect 11418 -14063 11468 -14029
rect 11452 -14097 11468 -14063
rect 11418 -14139 11468 -14097
rect 11556 -14034 11614 -13975
rect 11556 -14068 11568 -14034
rect 11602 -14068 11614 -14034
rect 11556 -14139 11614 -14068
rect 11648 -13961 11982 -13921
rect 11648 -13995 11666 -13961
rect 11700 -13995 11930 -13961
rect 11964 -13995 11982 -13961
rect 11648 -14063 11982 -13995
rect 11648 -14097 11666 -14063
rect 11700 -14097 11930 -14063
rect 11964 -14097 11982 -14063
rect 11648 -14139 11982 -14097
rect 13488 -13941 13546 -13906
rect 14130 -13921 14649 -13851
rect 14776 -13853 15292 -13783
rect 14776 -13887 14854 -13853
rect 14888 -13887 14982 -13853
rect 15016 -13887 15110 -13853
rect 15144 -13887 15238 -13853
rect 15272 -13887 15292 -13853
rect 15326 -13851 15346 -13817
rect 15380 -13851 15474 -13817
rect 15508 -13851 15602 -13817
rect 15636 -13851 15730 -13817
rect 15764 -13851 15845 -13817
rect 13488 -13975 13500 -13941
rect 13534 -13975 13546 -13941
rect 13488 -14034 13546 -13975
rect 13488 -14068 13500 -14034
rect 13534 -14068 13546 -14034
rect 13488 -14139 13546 -14068
rect 13580 -13961 14649 -13921
rect 13580 -13995 13598 -13961
rect 13632 -13995 14598 -13961
rect 14632 -13995 14649 -13961
rect 13580 -14063 14649 -13995
rect 13580 -14097 13598 -14063
rect 13632 -14097 14598 -14063
rect 14632 -14097 14649 -14063
rect 13580 -14139 14649 -14097
rect 14684 -13941 14742 -13906
rect 15326 -13921 15845 -13851
rect 15972 -13853 16302 -13783
rect 15972 -13887 16050 -13853
rect 16084 -13887 16149 -13853
rect 16183 -13887 16248 -13853
rect 16282 -13887 16302 -13853
rect 16336 -13851 16356 -13817
rect 16390 -13851 16459 -13817
rect 16493 -13851 16562 -13817
rect 16596 -13851 16674 -13817
rect 14684 -13975 14696 -13941
rect 14730 -13975 14742 -13941
rect 14684 -14034 14742 -13975
rect 14684 -14068 14696 -14034
rect 14730 -14068 14742 -14034
rect 14684 -14139 14742 -14068
rect 14776 -13961 15845 -13921
rect 14776 -13995 14794 -13961
rect 14828 -13995 15794 -13961
rect 15828 -13995 15845 -13961
rect 14776 -14063 15845 -13995
rect 14776 -14097 14794 -14063
rect 14828 -14097 15794 -14063
rect 15828 -14097 15845 -14063
rect 14776 -14139 15845 -14097
rect 15880 -13941 15938 -13906
rect 16336 -13921 16674 -13851
rect 15880 -13975 15892 -13941
rect 15926 -13975 15938 -13941
rect 15880 -14034 15938 -13975
rect 15880 -14068 15892 -14034
rect 15926 -14068 15938 -14034
rect 15880 -14139 15938 -14068
rect 15972 -13961 16674 -13921
rect 15972 -13995 15990 -13961
rect 16024 -13995 16622 -13961
rect 16656 -13995 16674 -13961
rect 15972 -14063 16674 -13995
rect 15972 -14097 15990 -14063
rect 16024 -14097 16622 -14063
rect 16656 -14097 16674 -14063
rect 15972 -14139 16674 -14097
rect -2997 -14173 -2968 -14139
rect -2934 -14173 -2876 -14139
rect -2842 -14173 -2784 -14139
rect -2750 -14173 -2692 -14139
rect -2658 -14173 -2600 -14139
rect -2566 -14173 -2508 -14139
rect -2474 -14173 -2416 -14139
rect -2382 -14173 -2324 -14139
rect -2290 -14173 -2232 -14139
rect -2198 -14173 -2140 -14139
rect -2106 -14173 -2048 -14139
rect -2014 -14173 -1956 -14139
rect -1922 -14173 -1864 -14139
rect -1830 -14173 -1772 -14139
rect -1738 -14173 -1680 -14139
rect -1646 -14173 -1588 -14139
rect -1554 -14173 -1496 -14139
rect -1462 -14173 -1404 -14139
rect -1370 -14173 -1312 -14139
rect -1278 -14173 -1220 -14139
rect -1186 -14173 -1128 -14139
rect -1094 -14173 -1036 -14139
rect -1002 -14173 -944 -14139
rect -910 -14173 -852 -14139
rect -818 -14173 -760 -14139
rect -726 -14173 -668 -14139
rect -634 -14173 -576 -14139
rect -542 -14173 -484 -14139
rect -450 -14173 -392 -14139
rect -358 -14173 -300 -14139
rect -266 -14173 -208 -14139
rect -174 -14173 -116 -14139
rect -82 -14173 -24 -14139
rect 10 -14173 68 -14139
rect 102 -14173 160 -14139
rect 194 -14173 252 -14139
rect 286 -14173 344 -14139
rect 378 -14173 436 -14139
rect 470 -14173 528 -14139
rect 562 -14173 620 -14139
rect 654 -14173 712 -14139
rect 746 -14173 804 -14139
rect 838 -14173 896 -14139
rect 930 -14173 988 -14139
rect 1022 -14173 1080 -14139
rect 1114 -14173 1172 -14139
rect 1206 -14173 1264 -14139
rect 1298 -14173 1356 -14139
rect 1390 -14173 1448 -14139
rect 1482 -14173 1540 -14139
rect 1574 -14173 1632 -14139
rect 1666 -14173 1724 -14139
rect 1758 -14173 1816 -14139
rect 1850 -14173 1908 -14139
rect 1942 -14173 2000 -14139
rect 2034 -14173 2092 -14139
rect 2126 -14173 2184 -14139
rect 2218 -14173 2276 -14139
rect 2310 -14173 2368 -14139
rect 2402 -14173 2460 -14139
rect 2494 -14173 2552 -14139
rect 2586 -14173 2644 -14139
rect 2678 -14173 2736 -14139
rect 2770 -14173 2828 -14139
rect 2862 -14173 2920 -14139
rect 2954 -14173 3012 -14139
rect 3046 -14173 3104 -14139
rect 3138 -14173 3196 -14139
rect 3230 -14173 3288 -14139
rect 3322 -14173 3380 -14139
rect 3414 -14173 3472 -14139
rect 3506 -14173 3564 -14139
rect 3598 -14173 3656 -14139
rect 3690 -14173 3748 -14139
rect 3782 -14173 3840 -14139
rect 3874 -14173 3932 -14139
rect 3966 -14173 4024 -14139
rect 4058 -14173 4116 -14139
rect 4150 -14173 4208 -14139
rect 4242 -14173 4300 -14139
rect 4334 -14173 4392 -14139
rect 4426 -14173 4484 -14139
rect 4518 -14173 4576 -14139
rect 4610 -14173 4668 -14139
rect 4702 -14173 4760 -14139
rect 4794 -14173 4852 -14139
rect 4886 -14173 4944 -14139
rect 4978 -14173 5036 -14139
rect 5070 -14173 5128 -14139
rect 5162 -14173 5220 -14139
rect 5254 -14173 5312 -14139
rect 5346 -14173 5404 -14139
rect 5438 -14173 5496 -14139
rect 5530 -14173 5588 -14139
rect 5622 -14173 5680 -14139
rect 5714 -14173 5772 -14139
rect 5806 -14173 5864 -14139
rect 5898 -14173 5956 -14139
rect 5990 -14173 6048 -14139
rect 6082 -14173 6140 -14139
rect 6174 -14173 6232 -14139
rect 6266 -14173 6324 -14139
rect 6358 -14173 6416 -14139
rect 6450 -14173 6508 -14139
rect 6542 -14173 6600 -14139
rect 6634 -14173 6692 -14139
rect 6726 -14173 6784 -14139
rect 6818 -14173 6876 -14139
rect 6910 -14173 6968 -14139
rect 7002 -14173 7060 -14139
rect 7094 -14173 7152 -14139
rect 7186 -14173 7244 -14139
rect 7278 -14173 7336 -14139
rect 7370 -14173 7428 -14139
rect 7462 -14173 7520 -14139
rect 7554 -14173 7612 -14139
rect 7646 -14173 7704 -14139
rect 7738 -14173 7796 -14139
rect 7830 -14173 7888 -14139
rect 7922 -14173 7980 -14139
rect 8014 -14173 8072 -14139
rect 8106 -14173 8164 -14139
rect 8198 -14173 8256 -14139
rect 8290 -14173 8348 -14139
rect 8382 -14173 8440 -14139
rect 8474 -14173 8532 -14139
rect 8566 -14173 8624 -14139
rect 8658 -14173 8716 -14139
rect 8750 -14173 8808 -14139
rect 8842 -14173 8900 -14139
rect 8934 -14173 8992 -14139
rect 9026 -14173 9084 -14139
rect 9118 -14173 9176 -14139
rect 9210 -14173 9268 -14139
rect 9302 -14173 9360 -14139
rect 9394 -14173 9452 -14139
rect 9486 -14173 9544 -14139
rect 9578 -14173 9636 -14139
rect 9670 -14173 9728 -14139
rect 9762 -14173 9820 -14139
rect 9854 -14173 9912 -14139
rect 9946 -14173 10004 -14139
rect 10038 -14173 10096 -14139
rect 10130 -14173 10188 -14139
rect 10222 -14173 10280 -14139
rect 10314 -14173 10372 -14139
rect 10406 -14173 10464 -14139
rect 10498 -14173 10556 -14139
rect 10590 -14173 10648 -14139
rect 10682 -14173 10740 -14139
rect 10774 -14173 10832 -14139
rect 10866 -14173 10924 -14139
rect 10958 -14173 11016 -14139
rect 11050 -14173 11108 -14139
rect 11142 -14173 11200 -14139
rect 11234 -14173 11292 -14139
rect 11326 -14173 11384 -14139
rect 11418 -14173 11476 -14139
rect 11510 -14173 11568 -14139
rect 11602 -14173 11660 -14139
rect 11694 -14173 11752 -14139
rect 11786 -14173 11844 -14139
rect 11878 -14173 11936 -14139
rect 11970 -14173 12028 -14139
rect 12062 -14173 12120 -14139
rect 12154 -14173 12212 -14139
rect 12246 -14173 12304 -14139
rect 12338 -14173 12396 -14139
rect 12430 -14173 12488 -14139
rect 12522 -14173 12580 -14139
rect 12614 -14173 12672 -14139
rect 12706 -14173 12764 -14139
rect 12798 -14173 12856 -14139
rect 12890 -14173 12948 -14139
rect 12982 -14173 13040 -14139
rect 13074 -14173 13132 -14139
rect 13166 -14173 13224 -14139
rect 13258 -14173 13316 -14139
rect 13350 -14173 13408 -14139
rect 13442 -14173 13500 -14139
rect 13534 -14173 13592 -14139
rect 13626 -14173 13684 -14139
rect 13718 -14173 13776 -14139
rect 13810 -14173 13868 -14139
rect 13902 -14173 13960 -14139
rect 13994 -14173 14052 -14139
rect 14086 -14173 14144 -14139
rect 14178 -14173 14236 -14139
rect 14270 -14173 14328 -14139
rect 14362 -14173 14420 -14139
rect 14454 -14173 14512 -14139
rect 14546 -14173 14604 -14139
rect 14638 -14173 14696 -14139
rect 14730 -14173 14788 -14139
rect 14822 -14173 14880 -14139
rect 14914 -14173 14972 -14139
rect 15006 -14173 15064 -14139
rect 15098 -14173 15156 -14139
rect 15190 -14173 15248 -14139
rect 15282 -14173 15340 -14139
rect 15374 -14173 15432 -14139
rect 15466 -14173 15524 -14139
rect 15558 -14173 15616 -14139
rect 15650 -14173 15708 -14139
rect 15742 -14173 15800 -14139
rect 15834 -14173 15892 -14139
rect 15926 -14173 15984 -14139
rect 16018 -14173 16076 -14139
rect 16110 -14173 16168 -14139
rect 16202 -14173 16260 -14139
rect 16294 -14173 16352 -14139
rect 16386 -14173 16444 -14139
rect 16478 -14173 16536 -14139
rect 16570 -14173 16628 -14139
rect 16662 -14173 16691 -14139
<< viali >>
rect -2968 -29 -2934 5
rect -2876 -29 -2842 5
rect -2784 -29 -2750 5
rect -2692 -29 -2658 5
rect -2600 -29 -2566 5
rect -2508 -29 -2474 5
rect -2416 -29 -2382 5
rect -2324 -29 -2290 5
rect -2232 -29 -2198 5
rect -2140 -29 -2106 5
rect -2048 -29 -2014 5
rect -1956 -29 -1922 5
rect -1864 -29 -1830 5
rect -1772 -29 -1738 5
rect -1680 -29 -1646 5
rect -1588 -29 -1554 5
rect -1496 -29 -1462 5
rect -1404 -29 -1370 5
rect -1312 -29 -1278 5
rect -1220 -29 -1186 5
rect -1128 -29 -1094 5
rect -1036 -29 -1002 5
rect -944 -29 -910 5
rect -852 -29 -818 5
rect -760 -29 -726 5
rect -668 -29 -634 5
rect -576 -29 -542 5
rect -484 -29 -450 5
rect -392 -29 -358 5
rect -300 -29 -266 5
rect -208 -29 -174 5
rect -116 -29 -82 5
rect -24 -29 10 5
rect 68 -29 102 5
rect 160 -29 194 5
rect 252 -29 286 5
rect 344 -29 378 5
rect 436 -29 470 5
rect 528 -29 562 5
rect 620 -29 654 5
rect 712 -29 746 5
rect 804 -29 838 5
rect 896 -29 930 5
rect 988 -29 1022 5
rect 1080 -29 1114 5
rect 1172 -29 1206 5
rect 1264 -29 1298 5
rect 1356 -29 1390 5
rect 1448 -29 1482 5
rect 1540 -29 1574 5
rect 1632 -29 1666 5
rect 1724 -29 1758 5
rect 1816 -29 1850 5
rect 1908 -29 1942 5
rect 2000 -29 2034 5
rect 2092 -29 2126 5
rect 2184 -29 2218 5
rect 2276 -29 2310 5
rect 2368 -29 2402 5
rect 2460 -29 2494 5
rect 2552 -29 2586 5
rect 2644 -29 2678 5
rect 2736 -29 2770 5
rect 2828 -29 2862 5
rect 2920 -29 2954 5
rect 3012 -29 3046 5
rect 3104 -29 3138 5
rect 3196 -29 3230 5
rect 3288 -29 3322 5
rect 3380 -29 3414 5
rect 3472 -29 3506 5
rect 3564 -29 3598 5
rect 3656 -29 3690 5
rect 3748 -29 3782 5
rect 3840 -29 3874 5
rect 3932 -29 3966 5
rect 4024 -29 4058 5
rect 4116 -29 4150 5
rect 4208 -29 4242 5
rect 4300 -29 4334 5
rect 4392 -29 4426 5
rect 4484 -29 4518 5
rect 4576 -29 4610 5
rect 4668 -29 4702 5
rect 4760 -29 4794 5
rect 4852 -29 4886 5
rect 4944 -29 4978 5
rect 5036 -29 5070 5
rect 5128 -29 5162 5
rect 5220 -29 5254 5
rect 5312 -29 5346 5
rect 5404 -29 5438 5
rect 5496 -29 5530 5
rect 5588 -29 5622 5
rect 5680 -29 5714 5
rect 5772 -29 5806 5
rect 5864 -29 5898 5
rect 5956 -29 5990 5
rect 6048 -29 6082 5
rect 6140 -29 6174 5
rect 6232 -29 6266 5
rect 6324 -29 6358 5
rect 6416 -29 6450 5
rect 6508 -29 6542 5
rect 6600 -29 6634 5
rect 6692 -29 6726 5
rect 6784 -29 6818 5
rect 6876 -29 6910 5
rect 6968 -29 7002 5
rect 7060 -29 7094 5
rect 7152 -29 7186 5
rect 7244 -29 7278 5
rect 7336 -29 7370 5
rect 7428 -29 7462 5
rect 7520 -29 7554 5
rect 7612 -29 7646 5
rect 7704 -29 7738 5
rect 7796 -29 7830 5
rect 7888 -29 7922 5
rect 7980 -29 8014 5
rect 8072 -29 8106 5
rect 8164 -29 8198 5
rect 8256 -29 8290 5
rect 8348 -29 8382 5
rect 8440 -29 8474 5
rect 8532 -29 8566 5
rect 8624 -29 8658 5
rect 8716 -29 8750 5
rect 8808 -29 8842 5
rect 8900 -29 8934 5
rect 8992 -29 9026 5
rect 9084 -29 9118 5
rect 9176 -29 9210 5
rect 9268 -29 9302 5
rect 9360 -29 9394 5
rect 9452 -29 9486 5
rect 9544 -29 9578 5
rect 9636 -29 9670 5
rect 9728 -29 9762 5
rect 9820 -29 9854 5
rect 9912 -29 9946 5
rect 10004 -29 10038 5
rect 10096 -29 10130 5
rect 10188 -29 10222 5
rect 10280 -29 10314 5
rect 10372 -29 10406 5
rect 10464 -29 10498 5
rect 10556 -29 10590 5
rect 10648 -29 10682 5
rect 10740 -29 10774 5
rect 10832 -29 10866 5
rect 10924 -29 10958 5
rect 11016 -29 11050 5
rect 11108 -29 11142 5
rect 11200 -29 11234 5
rect 11292 -29 11326 5
rect 11384 -29 11418 5
rect 11476 -29 11510 5
rect 11568 -29 11602 5
rect 11660 -29 11694 5
rect 11752 -29 11786 5
rect 11844 -29 11878 5
rect 11936 -29 11970 5
rect 12028 -29 12062 5
rect 12120 -29 12154 5
rect 12212 -29 12246 5
rect 12304 -29 12338 5
rect 12396 -29 12430 5
rect 12488 -29 12522 5
rect 12580 -29 12614 5
rect 12672 -29 12706 5
rect 12764 -29 12798 5
rect 12856 -29 12890 5
rect 12948 -29 12982 5
rect 13040 -29 13074 5
rect 13132 -29 13166 5
rect 13224 -29 13258 5
rect 13316 -29 13350 5
rect 13408 -29 13442 5
rect 13500 -29 13534 5
rect 13592 -29 13626 5
rect 13684 -29 13718 5
rect 13776 -29 13810 5
rect 13868 -29 13902 5
rect 13960 -29 13994 5
rect 14052 -29 14086 5
rect 14144 -29 14178 5
rect 14236 -29 14270 5
rect 14328 -29 14362 5
rect 14420 -29 14454 5
rect 14512 -29 14546 5
rect 14604 -29 14638 5
rect 14696 -29 14730 5
rect 14788 -29 14822 5
rect 14880 -29 14914 5
rect 14972 -29 15006 5
rect 15064 -29 15098 5
rect 15156 -29 15190 5
rect 15248 -29 15282 5
rect 15340 -29 15374 5
rect 15432 -29 15466 5
rect 15524 -29 15558 5
rect 15616 -29 15650 5
rect 15708 -29 15742 5
rect 15800 -29 15834 5
rect 15892 -29 15926 5
rect 15984 -29 16018 5
rect 16076 -29 16110 5
rect 16168 -29 16202 5
rect 16260 -29 16294 5
rect 16352 -29 16386 5
rect 16444 -29 16478 5
rect 16536 -29 16570 5
rect 16628 -29 16662 5
rect -943 -307 -909 -301
rect -943 -335 -937 -307
rect -937 -335 -909 -307
rect -762 -307 -728 -301
rect -762 -335 -735 -307
rect -735 -335 -728 -307
rect -30 -341 4 -307
rect 106 -341 140 -307
rect 242 -341 276 -307
rect 434 -379 468 -345
rect -848 -446 -814 -412
rect -769 -429 -766 -412
rect -766 -429 -735 -412
rect -769 -446 -735 -429
rect 1076 -341 1082 -312
rect 1082 -341 1110 -312
rect 1076 -346 1110 -341
rect 1076 -419 1110 -385
rect 1171 -340 1205 -306
rect 1263 -340 1297 -306
rect 2369 -307 2403 -301
rect 2369 -335 2396 -307
rect 2396 -335 2403 -307
rect 3015 -336 3049 -302
rect 6876 -307 6910 -302
rect 6876 -336 6904 -307
rect 6904 -336 6910 -307
rect 7522 -336 7556 -302
rect 8164 -307 8198 -303
rect 8164 -337 8192 -307
rect 8192 -337 8198 -307
rect 8811 -335 8845 -301
rect 9453 -307 9487 -301
rect 9453 -335 9480 -307
rect 9480 -335 9487 -307
rect 10099 -334 10133 -300
rect 10741 -307 10775 -301
rect 10832 -307 10866 -301
rect 10925 -307 10959 -302
rect 11017 -307 11051 -302
rect 10741 -335 10749 -307
rect 10749 -335 10775 -307
rect 10832 -335 10864 -307
rect 10864 -335 10866 -307
rect 10925 -336 10948 -307
rect 10948 -336 10959 -307
rect 11017 -336 11032 -307
rect 11032 -336 11051 -307
rect 11129 -302 11163 -268
rect 11250 -307 11284 -299
rect 11344 -307 11378 -299
rect 11250 -333 11284 -307
rect 11344 -333 11368 -307
rect 11368 -333 11378 -307
rect -2968 -573 -2934 -539
rect -2876 -573 -2842 -539
rect -2784 -573 -2750 -539
rect -2692 -573 -2658 -539
rect -2600 -573 -2566 -539
rect -2508 -573 -2474 -539
rect -2416 -573 -2382 -539
rect -2324 -573 -2290 -539
rect -2232 -573 -2198 -539
rect -2140 -573 -2106 -539
rect -2048 -573 -2014 -539
rect -1956 -573 -1922 -539
rect -1864 -573 -1830 -539
rect -1772 -573 -1738 -539
rect -1680 -573 -1646 -539
rect -1588 -573 -1554 -539
rect -1496 -573 -1462 -539
rect -1404 -573 -1370 -539
rect -1312 -573 -1278 -539
rect -1220 -573 -1186 -539
rect -1128 -573 -1094 -539
rect -1036 -573 -1002 -539
rect -944 -573 -910 -539
rect -852 -573 -818 -539
rect -760 -573 -726 -539
rect -668 -573 -634 -539
rect -576 -573 -542 -539
rect -484 -573 -450 -539
rect -392 -573 -358 -539
rect -300 -573 -266 -539
rect -208 -573 -174 -539
rect -116 -573 -82 -539
rect -24 -573 10 -539
rect 68 -573 102 -539
rect 160 -573 194 -539
rect 252 -573 286 -539
rect 344 -573 378 -539
rect 436 -573 470 -539
rect 528 -573 562 -539
rect 620 -573 654 -539
rect 712 -573 746 -539
rect 804 -573 838 -539
rect 896 -573 930 -539
rect 988 -573 1022 -539
rect 1080 -573 1114 -539
rect 1172 -573 1206 -539
rect 1264 -573 1298 -539
rect 1356 -573 1390 -539
rect 1448 -573 1482 -539
rect 1540 -573 1574 -539
rect 1632 -573 1666 -539
rect 1724 -573 1758 -539
rect 1816 -573 1850 -539
rect 1908 -573 1942 -539
rect 2000 -573 2034 -539
rect 2092 -573 2126 -539
rect 2184 -573 2218 -539
rect 2276 -573 2310 -539
rect 2368 -573 2402 -539
rect 2460 -573 2494 -539
rect 2552 -573 2586 -539
rect 2644 -573 2678 -539
rect 2736 -573 2770 -539
rect 2828 -573 2862 -539
rect 2920 -573 2954 -539
rect 3012 -573 3046 -539
rect 3104 -573 3138 -539
rect 3196 -573 3230 -539
rect 3288 -573 3322 -539
rect 3380 -573 3414 -539
rect 3472 -573 3506 -539
rect 3564 -573 3598 -539
rect 3656 -573 3690 -539
rect 3748 -573 3782 -539
rect 3840 -573 3874 -539
rect 3932 -573 3966 -539
rect 4024 -573 4058 -539
rect 4116 -573 4150 -539
rect 4208 -573 4242 -539
rect 4300 -573 4334 -539
rect 4392 -573 4426 -539
rect 4484 -573 4518 -539
rect 4576 -573 4610 -539
rect 4668 -573 4702 -539
rect 4760 -573 4794 -539
rect 4852 -573 4886 -539
rect 4944 -573 4978 -539
rect 5036 -573 5070 -539
rect 5128 -573 5162 -539
rect 5220 -573 5254 -539
rect 5312 -573 5346 -539
rect 5404 -573 5438 -539
rect 5496 -573 5530 -539
rect 5588 -573 5622 -539
rect 5680 -573 5714 -539
rect 5772 -573 5806 -539
rect 5864 -573 5898 -539
rect 5956 -573 5990 -539
rect 6048 -573 6082 -539
rect 6140 -573 6174 -539
rect 6232 -573 6266 -539
rect 6324 -573 6358 -539
rect 6416 -573 6450 -539
rect 6508 -573 6542 -539
rect 6600 -573 6634 -539
rect 6692 -573 6726 -539
rect 6784 -573 6818 -539
rect 6876 -573 6910 -539
rect 6968 -573 7002 -539
rect 7060 -573 7094 -539
rect 7152 -573 7186 -539
rect 7244 -573 7278 -539
rect 7336 -573 7370 -539
rect 7428 -573 7462 -539
rect 7520 -573 7554 -539
rect 7612 -573 7646 -539
rect 7704 -573 7738 -539
rect 7796 -573 7830 -539
rect 7888 -573 7922 -539
rect 7980 -573 8014 -539
rect 8072 -573 8106 -539
rect 8164 -573 8198 -539
rect 8256 -573 8290 -539
rect 8348 -573 8382 -539
rect 8440 -573 8474 -539
rect 8532 -573 8566 -539
rect 8624 -573 8658 -539
rect 8716 -573 8750 -539
rect 8808 -573 8842 -539
rect 8900 -573 8934 -539
rect 8992 -573 9026 -539
rect 9084 -573 9118 -539
rect 9176 -573 9210 -539
rect 9268 -573 9302 -539
rect 9360 -573 9394 -539
rect 9452 -573 9486 -539
rect 9544 -573 9578 -539
rect 9636 -573 9670 -539
rect 9728 -573 9762 -539
rect 9820 -573 9854 -539
rect 9912 -573 9946 -539
rect 10004 -573 10038 -539
rect 10096 -573 10130 -539
rect 10188 -573 10222 -539
rect 10280 -573 10314 -539
rect 10372 -573 10406 -539
rect 10464 -573 10498 -539
rect 10556 -573 10590 -539
rect 10648 -573 10682 -539
rect 10740 -573 10774 -539
rect 10832 -573 10866 -539
rect 10924 -573 10958 -539
rect 11016 -573 11050 -539
rect 11108 -573 11142 -539
rect 11200 -573 11234 -539
rect 11292 -573 11326 -539
rect 11384 -573 11418 -539
rect 11476 -573 11510 -539
rect 11568 -573 11602 -539
rect 11660 -573 11694 -539
rect 11752 -573 11786 -539
rect 11844 -573 11878 -539
rect 11936 -573 11970 -539
rect 12028 -573 12062 -539
rect 12120 -573 12154 -539
rect 12212 -573 12246 -539
rect 12304 -573 12338 -539
rect 12396 -573 12430 -539
rect 12488 -573 12522 -539
rect 12580 -573 12614 -539
rect 12672 -573 12706 -539
rect 12764 -573 12798 -539
rect 12856 -573 12890 -539
rect 12948 -573 12982 -539
rect 13040 -573 13074 -539
rect 13132 -573 13166 -539
rect 13224 -573 13258 -539
rect 13316 -573 13350 -539
rect 13408 -573 13442 -539
rect 13500 -573 13534 -539
rect 13592 -573 13626 -539
rect 13684 -573 13718 -539
rect 13776 -573 13810 -539
rect 13868 -573 13902 -539
rect 13960 -573 13994 -539
rect 14052 -573 14086 -539
rect 14144 -573 14178 -539
rect 14236 -573 14270 -539
rect 14328 -573 14362 -539
rect 14420 -573 14454 -539
rect 14512 -573 14546 -539
rect 14604 -573 14638 -539
rect 14696 -573 14730 -539
rect 14788 -573 14822 -539
rect 14880 -573 14914 -539
rect 14972 -573 15006 -539
rect 15064 -573 15098 -539
rect 15156 -573 15190 -539
rect 15248 -573 15282 -539
rect 15340 -573 15374 -539
rect 15432 -573 15466 -539
rect 15524 -573 15558 -539
rect 15616 -573 15650 -539
rect 15708 -573 15742 -539
rect 15800 -573 15834 -539
rect 15892 -573 15926 -539
rect 15984 -573 16018 -539
rect 16076 -573 16110 -539
rect 16168 -573 16202 -539
rect 16260 -573 16294 -539
rect 16352 -573 16386 -539
rect 16444 -573 16478 -539
rect 16536 -573 16570 -539
rect 16628 -573 16662 -539
rect 433 -846 467 -812
rect 1052 -805 1086 -775
rect 1052 -809 1086 -805
rect 3012 -809 3046 -775
rect 3626 -805 3628 -775
rect 3628 -805 3660 -775
rect 3626 -809 3660 -805
rect 5586 -809 5620 -775
rect 6200 -805 6204 -775
rect 6204 -805 6234 -775
rect 6200 -809 6234 -805
rect 8160 -809 8194 -775
rect 8774 -805 8780 -775
rect 8780 -805 8808 -775
rect 8774 -809 8808 -805
rect 10737 -811 10771 -777
rect 11369 -805 11390 -778
rect 11390 -805 11403 -778
rect 11369 -812 11403 -805
rect 13685 -771 13719 -746
rect 13685 -780 13692 -771
rect 13692 -780 13719 -771
rect 15248 -762 15282 -728
rect 15340 -763 15374 -729
rect 15248 -858 15282 -824
rect 15341 -858 15375 -824
rect -2968 -1117 -2934 -1083
rect -2876 -1117 -2842 -1083
rect -2784 -1117 -2750 -1083
rect -2692 -1117 -2658 -1083
rect -2600 -1117 -2566 -1083
rect -2508 -1117 -2474 -1083
rect -2416 -1117 -2382 -1083
rect -2324 -1117 -2290 -1083
rect -2232 -1117 -2198 -1083
rect -2140 -1117 -2106 -1083
rect -2048 -1117 -2014 -1083
rect -1956 -1117 -1922 -1083
rect -1864 -1117 -1830 -1083
rect -1772 -1117 -1738 -1083
rect -1680 -1117 -1646 -1083
rect -1588 -1117 -1554 -1083
rect -1496 -1117 -1462 -1083
rect -1404 -1117 -1370 -1083
rect -1312 -1117 -1278 -1083
rect -1220 -1117 -1186 -1083
rect -1128 -1117 -1094 -1083
rect -1036 -1117 -1002 -1083
rect -944 -1117 -910 -1083
rect -852 -1117 -818 -1083
rect -760 -1117 -726 -1083
rect -668 -1117 -634 -1083
rect -576 -1117 -542 -1083
rect -484 -1117 -450 -1083
rect -392 -1117 -358 -1083
rect -300 -1117 -266 -1083
rect -208 -1117 -174 -1083
rect -116 -1117 -82 -1083
rect -24 -1117 10 -1083
rect 68 -1117 102 -1083
rect 160 -1117 194 -1083
rect 252 -1117 286 -1083
rect 344 -1117 378 -1083
rect 436 -1117 470 -1083
rect 528 -1117 562 -1083
rect 620 -1117 654 -1083
rect 712 -1117 746 -1083
rect 804 -1117 838 -1083
rect 896 -1117 930 -1083
rect 988 -1117 1022 -1083
rect 1080 -1117 1114 -1083
rect 1172 -1117 1206 -1083
rect 1264 -1117 1298 -1083
rect 1356 -1117 1390 -1083
rect 1448 -1117 1482 -1083
rect 1540 -1117 1574 -1083
rect 1632 -1117 1666 -1083
rect 1724 -1117 1758 -1083
rect 1816 -1117 1850 -1083
rect 1908 -1117 1942 -1083
rect 2000 -1117 2034 -1083
rect 2092 -1117 2126 -1083
rect 2184 -1117 2218 -1083
rect 2276 -1117 2310 -1083
rect 2368 -1117 2402 -1083
rect 2460 -1117 2494 -1083
rect 2552 -1117 2586 -1083
rect 2644 -1117 2678 -1083
rect 2736 -1117 2770 -1083
rect 2828 -1117 2862 -1083
rect 2920 -1117 2954 -1083
rect 3012 -1117 3046 -1083
rect 3104 -1117 3138 -1083
rect 3196 -1117 3230 -1083
rect 3288 -1117 3322 -1083
rect 3380 -1117 3414 -1083
rect 3472 -1117 3506 -1083
rect 3564 -1117 3598 -1083
rect 3656 -1117 3690 -1083
rect 3748 -1117 3782 -1083
rect 3840 -1117 3874 -1083
rect 3932 -1117 3966 -1083
rect 4024 -1117 4058 -1083
rect 4116 -1117 4150 -1083
rect 4208 -1117 4242 -1083
rect 4300 -1117 4334 -1083
rect 4392 -1117 4426 -1083
rect 4484 -1117 4518 -1083
rect 4576 -1117 4610 -1083
rect 4668 -1117 4702 -1083
rect 4760 -1117 4794 -1083
rect 4852 -1117 4886 -1083
rect 4944 -1117 4978 -1083
rect 5036 -1117 5070 -1083
rect 5128 -1117 5162 -1083
rect 5220 -1117 5254 -1083
rect 5312 -1117 5346 -1083
rect 5404 -1117 5438 -1083
rect 5496 -1117 5530 -1083
rect 5588 -1117 5622 -1083
rect 5680 -1117 5714 -1083
rect 5772 -1117 5806 -1083
rect 5864 -1117 5898 -1083
rect 5956 -1117 5990 -1083
rect 6048 -1117 6082 -1083
rect 6140 -1117 6174 -1083
rect 6232 -1117 6266 -1083
rect 6324 -1117 6358 -1083
rect 6416 -1117 6450 -1083
rect 6508 -1117 6542 -1083
rect 6600 -1117 6634 -1083
rect 6692 -1117 6726 -1083
rect 6784 -1117 6818 -1083
rect 6876 -1117 6910 -1083
rect 6968 -1117 7002 -1083
rect 7060 -1117 7094 -1083
rect 7152 -1117 7186 -1083
rect 7244 -1117 7278 -1083
rect 7336 -1117 7370 -1083
rect 7428 -1117 7462 -1083
rect 7520 -1117 7554 -1083
rect 7612 -1117 7646 -1083
rect 7704 -1117 7738 -1083
rect 7796 -1117 7830 -1083
rect 7888 -1117 7922 -1083
rect 7980 -1117 8014 -1083
rect 8072 -1117 8106 -1083
rect 8164 -1117 8198 -1083
rect 8256 -1117 8290 -1083
rect 8348 -1117 8382 -1083
rect 8440 -1117 8474 -1083
rect 8532 -1117 8566 -1083
rect 8624 -1117 8658 -1083
rect 8716 -1117 8750 -1083
rect 8808 -1117 8842 -1083
rect 8900 -1117 8934 -1083
rect 8992 -1117 9026 -1083
rect 9084 -1117 9118 -1083
rect 9176 -1117 9210 -1083
rect 9268 -1117 9302 -1083
rect 9360 -1117 9394 -1083
rect 9452 -1117 9486 -1083
rect 9544 -1117 9578 -1083
rect 9636 -1117 9670 -1083
rect 9728 -1117 9762 -1083
rect 9820 -1117 9854 -1083
rect 9912 -1117 9946 -1083
rect 10004 -1117 10038 -1083
rect 10096 -1117 10130 -1083
rect 10188 -1117 10222 -1083
rect 10280 -1117 10314 -1083
rect 10372 -1117 10406 -1083
rect 10464 -1117 10498 -1083
rect 10556 -1117 10590 -1083
rect 10648 -1117 10682 -1083
rect 10740 -1117 10774 -1083
rect 10832 -1117 10866 -1083
rect 10924 -1117 10958 -1083
rect 11016 -1117 11050 -1083
rect 11108 -1117 11142 -1083
rect 11200 -1117 11234 -1083
rect 11292 -1117 11326 -1083
rect 11384 -1117 11418 -1083
rect 11476 -1117 11510 -1083
rect 11568 -1117 11602 -1083
rect 11660 -1117 11694 -1083
rect 11752 -1117 11786 -1083
rect 11844 -1117 11878 -1083
rect 11936 -1117 11970 -1083
rect 12028 -1117 12062 -1083
rect 12120 -1117 12154 -1083
rect 12212 -1117 12246 -1083
rect 12304 -1117 12338 -1083
rect 12396 -1117 12430 -1083
rect 12488 -1117 12522 -1083
rect 12580 -1117 12614 -1083
rect 12672 -1117 12706 -1083
rect 12764 -1117 12798 -1083
rect 12856 -1117 12890 -1083
rect 12948 -1117 12982 -1083
rect 13040 -1117 13074 -1083
rect 13132 -1117 13166 -1083
rect 13224 -1117 13258 -1083
rect 13316 -1117 13350 -1083
rect 13408 -1117 13442 -1083
rect 13500 -1117 13534 -1083
rect 13592 -1117 13626 -1083
rect 13684 -1117 13718 -1083
rect 13776 -1117 13810 -1083
rect 13868 -1117 13902 -1083
rect 13960 -1117 13994 -1083
rect 14052 -1117 14086 -1083
rect 14144 -1117 14178 -1083
rect 14236 -1117 14270 -1083
rect 14328 -1117 14362 -1083
rect 14420 -1117 14454 -1083
rect 14512 -1117 14546 -1083
rect 14604 -1117 14638 -1083
rect 14696 -1117 14730 -1083
rect 14788 -1117 14822 -1083
rect 14880 -1117 14914 -1083
rect 14972 -1117 15006 -1083
rect 15064 -1117 15098 -1083
rect 15156 -1117 15190 -1083
rect 15248 -1117 15282 -1083
rect 15340 -1117 15374 -1083
rect 15432 -1117 15466 -1083
rect 15524 -1117 15558 -1083
rect 15616 -1117 15650 -1083
rect 15708 -1117 15742 -1083
rect 15800 -1117 15834 -1083
rect 15892 -1117 15926 -1083
rect 15984 -1117 16018 -1083
rect 16076 -1117 16110 -1083
rect 16168 -1117 16202 -1083
rect 16260 -1117 16294 -1083
rect 16352 -1117 16386 -1083
rect 16444 -1117 16478 -1083
rect 16536 -1117 16570 -1083
rect 16628 -1117 16662 -1083
rect 432 -1395 466 -1392
rect 432 -1426 464 -1395
rect 464 -1426 466 -1395
rect 1082 -1423 1116 -1389
rect 3042 -1395 3076 -1389
rect 3042 -1423 3074 -1395
rect 3074 -1423 3076 -1395
rect 3656 -1423 3690 -1389
rect 5616 -1395 5650 -1389
rect 5616 -1423 5650 -1395
rect 6230 -1423 6264 -1389
rect 8190 -1395 8224 -1389
rect 8190 -1423 8192 -1395
rect 8192 -1423 8224 -1395
rect 8804 -1423 8838 -1389
rect 10764 -1395 10798 -1389
rect 10764 -1423 10768 -1395
rect 10768 -1423 10798 -1395
rect 11387 -1389 11421 -1355
rect 12558 -1395 12592 -1392
rect 12642 -1395 12676 -1392
rect 12739 -1395 12773 -1392
rect 12836 -1395 12870 -1392
rect 12942 -1395 12976 -1392
rect 12558 -1426 12574 -1395
rect 12574 -1426 12592 -1395
rect 12642 -1426 12676 -1395
rect 12739 -1426 12744 -1395
rect 12744 -1426 12773 -1395
rect 12836 -1426 12846 -1395
rect 12846 -1426 12870 -1395
rect 12942 -1426 12948 -1395
rect 12948 -1426 12976 -1395
rect 13038 -1419 13072 -1385
rect 13038 -1491 13072 -1457
rect 15248 -1372 15282 -1338
rect 15340 -1373 15374 -1339
rect 13684 -1429 13692 -1422
rect 13692 -1429 13718 -1422
rect 13684 -1456 13718 -1429
rect 15248 -1468 15282 -1434
rect 15341 -1468 15375 -1434
rect -2968 -1661 -2934 -1627
rect -2876 -1661 -2842 -1627
rect -2784 -1661 -2750 -1627
rect -2692 -1661 -2658 -1627
rect -2600 -1661 -2566 -1627
rect -2508 -1661 -2474 -1627
rect -2416 -1661 -2382 -1627
rect -2324 -1661 -2290 -1627
rect -2232 -1661 -2198 -1627
rect -2140 -1661 -2106 -1627
rect -2048 -1661 -2014 -1627
rect -1956 -1661 -1922 -1627
rect -1864 -1661 -1830 -1627
rect -1772 -1661 -1738 -1627
rect -1680 -1661 -1646 -1627
rect -1588 -1661 -1554 -1627
rect -1496 -1661 -1462 -1627
rect -1404 -1661 -1370 -1627
rect -1312 -1661 -1278 -1627
rect -1220 -1661 -1186 -1627
rect -1128 -1661 -1094 -1627
rect -1036 -1661 -1002 -1627
rect -944 -1661 -910 -1627
rect -852 -1661 -818 -1627
rect -760 -1661 -726 -1627
rect -668 -1661 -634 -1627
rect -576 -1661 -542 -1627
rect -484 -1661 -450 -1627
rect -392 -1661 -358 -1627
rect -300 -1661 -266 -1627
rect -208 -1661 -174 -1627
rect -116 -1661 -82 -1627
rect -24 -1661 10 -1627
rect 68 -1661 102 -1627
rect 160 -1661 194 -1627
rect 252 -1661 286 -1627
rect 344 -1661 378 -1627
rect 436 -1661 470 -1627
rect 528 -1661 562 -1627
rect 620 -1661 654 -1627
rect 712 -1661 746 -1627
rect 804 -1661 838 -1627
rect 896 -1661 930 -1627
rect 988 -1661 1022 -1627
rect 1080 -1661 1114 -1627
rect 1172 -1661 1206 -1627
rect 1264 -1661 1298 -1627
rect 1356 -1661 1390 -1627
rect 1448 -1661 1482 -1627
rect 1540 -1661 1574 -1627
rect 1632 -1661 1666 -1627
rect 1724 -1661 1758 -1627
rect 1816 -1661 1850 -1627
rect 1908 -1661 1942 -1627
rect 2000 -1661 2034 -1627
rect 2092 -1661 2126 -1627
rect 2184 -1661 2218 -1627
rect 2276 -1661 2310 -1627
rect 2368 -1661 2402 -1627
rect 2460 -1661 2494 -1627
rect 2552 -1661 2586 -1627
rect 2644 -1661 2678 -1627
rect 2736 -1661 2770 -1627
rect 2828 -1661 2862 -1627
rect 2920 -1661 2954 -1627
rect 3012 -1661 3046 -1627
rect 3104 -1661 3138 -1627
rect 3196 -1661 3230 -1627
rect 3288 -1661 3322 -1627
rect 3380 -1661 3414 -1627
rect 3472 -1661 3506 -1627
rect 3564 -1661 3598 -1627
rect 3656 -1661 3690 -1627
rect 3748 -1661 3782 -1627
rect 3840 -1661 3874 -1627
rect 3932 -1661 3966 -1627
rect 4024 -1661 4058 -1627
rect 4116 -1661 4150 -1627
rect 4208 -1661 4242 -1627
rect 4300 -1661 4334 -1627
rect 4392 -1661 4426 -1627
rect 4484 -1661 4518 -1627
rect 4576 -1661 4610 -1627
rect 4668 -1661 4702 -1627
rect 4760 -1661 4794 -1627
rect 4852 -1661 4886 -1627
rect 4944 -1661 4978 -1627
rect 5036 -1661 5070 -1627
rect 5128 -1661 5162 -1627
rect 5220 -1661 5254 -1627
rect 5312 -1661 5346 -1627
rect 5404 -1661 5438 -1627
rect 5496 -1661 5530 -1627
rect 5588 -1661 5622 -1627
rect 5680 -1661 5714 -1627
rect 5772 -1661 5806 -1627
rect 5864 -1661 5898 -1627
rect 5956 -1661 5990 -1627
rect 6048 -1661 6082 -1627
rect 6140 -1661 6174 -1627
rect 6232 -1661 6266 -1627
rect 6324 -1661 6358 -1627
rect 6416 -1661 6450 -1627
rect 6508 -1661 6542 -1627
rect 6600 -1661 6634 -1627
rect 6692 -1661 6726 -1627
rect 6784 -1661 6818 -1627
rect 6876 -1661 6910 -1627
rect 6968 -1661 7002 -1627
rect 7060 -1661 7094 -1627
rect 7152 -1661 7186 -1627
rect 7244 -1661 7278 -1627
rect 7336 -1661 7370 -1627
rect 7428 -1661 7462 -1627
rect 7520 -1661 7554 -1627
rect 7612 -1661 7646 -1627
rect 7704 -1661 7738 -1627
rect 7796 -1661 7830 -1627
rect 7888 -1661 7922 -1627
rect 7980 -1661 8014 -1627
rect 8072 -1661 8106 -1627
rect 8164 -1661 8198 -1627
rect 8256 -1661 8290 -1627
rect 8348 -1661 8382 -1627
rect 8440 -1661 8474 -1627
rect 8532 -1661 8566 -1627
rect 8624 -1661 8658 -1627
rect 8716 -1661 8750 -1627
rect 8808 -1661 8842 -1627
rect 8900 -1661 8934 -1627
rect 8992 -1661 9026 -1627
rect 9084 -1661 9118 -1627
rect 9176 -1661 9210 -1627
rect 9268 -1661 9302 -1627
rect 9360 -1661 9394 -1627
rect 9452 -1661 9486 -1627
rect 9544 -1661 9578 -1627
rect 9636 -1661 9670 -1627
rect 9728 -1661 9762 -1627
rect 9820 -1661 9854 -1627
rect 9912 -1661 9946 -1627
rect 10004 -1661 10038 -1627
rect 10096 -1661 10130 -1627
rect 10188 -1661 10222 -1627
rect 10280 -1661 10314 -1627
rect 10372 -1661 10406 -1627
rect 10464 -1661 10498 -1627
rect 10556 -1661 10590 -1627
rect 10648 -1661 10682 -1627
rect 10740 -1661 10774 -1627
rect 10832 -1661 10866 -1627
rect 10924 -1661 10958 -1627
rect 11016 -1661 11050 -1627
rect 11108 -1661 11142 -1627
rect 11200 -1661 11234 -1627
rect 11292 -1661 11326 -1627
rect 11384 -1661 11418 -1627
rect 11476 -1661 11510 -1627
rect 11568 -1661 11602 -1627
rect 11660 -1661 11694 -1627
rect 11752 -1661 11786 -1627
rect 11844 -1661 11878 -1627
rect 11936 -1661 11970 -1627
rect 12028 -1661 12062 -1627
rect 12120 -1661 12154 -1627
rect 12212 -1661 12246 -1627
rect 12304 -1661 12338 -1627
rect 12396 -1661 12430 -1627
rect 12488 -1661 12522 -1627
rect 12580 -1661 12614 -1627
rect 12672 -1661 12706 -1627
rect 12764 -1661 12798 -1627
rect 12856 -1661 12890 -1627
rect 12948 -1661 12982 -1627
rect 13040 -1661 13074 -1627
rect 13132 -1661 13166 -1627
rect 13224 -1661 13258 -1627
rect 13316 -1661 13350 -1627
rect 13408 -1661 13442 -1627
rect 13500 -1661 13534 -1627
rect 13592 -1661 13626 -1627
rect 13684 -1661 13718 -1627
rect 13776 -1661 13810 -1627
rect 13868 -1661 13902 -1627
rect 13960 -1661 13994 -1627
rect 14052 -1661 14086 -1627
rect 14144 -1661 14178 -1627
rect 14236 -1661 14270 -1627
rect 14328 -1661 14362 -1627
rect 14420 -1661 14454 -1627
rect 14512 -1661 14546 -1627
rect 14604 -1661 14638 -1627
rect 14696 -1661 14730 -1627
rect 14788 -1661 14822 -1627
rect 14880 -1661 14914 -1627
rect 14972 -1661 15006 -1627
rect 15064 -1661 15098 -1627
rect 15156 -1661 15190 -1627
rect 15248 -1661 15282 -1627
rect 15340 -1661 15374 -1627
rect 15432 -1661 15466 -1627
rect 15524 -1661 15558 -1627
rect 15616 -1661 15650 -1627
rect 15708 -1661 15742 -1627
rect 15800 -1661 15834 -1627
rect 15892 -1661 15926 -1627
rect 15984 -1661 16018 -1627
rect 16076 -1661 16110 -1627
rect 16168 -1661 16202 -1627
rect 16260 -1661 16294 -1627
rect 16352 -1661 16386 -1627
rect 16444 -1661 16478 -1627
rect 16536 -1661 16570 -1627
rect 16628 -1661 16662 -1627
rect -856 -1934 -822 -1900
rect -210 -1893 -202 -1865
rect -202 -1893 -176 -1865
rect -210 -1899 -176 -1893
rect 432 -1934 466 -1900
rect 1054 -1893 1086 -1866
rect 1086 -1893 1088 -1866
rect 1054 -1900 1088 -1893
rect 3014 -1900 3048 -1866
rect 3628 -1893 3662 -1866
rect 3628 -1900 3662 -1893
rect 5588 -1900 5622 -1866
rect 6202 -1893 6204 -1866
rect 6204 -1893 6236 -1866
rect 6202 -1900 6236 -1893
rect 8162 -1900 8196 -1866
rect 8776 -1893 8780 -1866
rect 8780 -1893 8810 -1866
rect 8776 -1900 8810 -1893
rect 10736 -1900 10770 -1866
rect 11386 -1893 11390 -1863
rect 11390 -1893 11420 -1863
rect 11386 -1897 11420 -1893
rect 13685 -1859 13719 -1832
rect 13685 -1866 13692 -1859
rect 13692 -1866 13719 -1859
rect 15248 -1850 15282 -1816
rect 15340 -1851 15374 -1817
rect 15248 -1946 15282 -1912
rect 15341 -1946 15375 -1912
rect -2968 -2205 -2934 -2171
rect -2876 -2205 -2842 -2171
rect -2784 -2205 -2750 -2171
rect -2692 -2205 -2658 -2171
rect -2600 -2205 -2566 -2171
rect -2508 -2205 -2474 -2171
rect -2416 -2205 -2382 -2171
rect -2324 -2205 -2290 -2171
rect -2232 -2205 -2198 -2171
rect -2140 -2205 -2106 -2171
rect -2048 -2205 -2014 -2171
rect -1956 -2205 -1922 -2171
rect -1864 -2205 -1830 -2171
rect -1772 -2205 -1738 -2171
rect -1680 -2205 -1646 -2171
rect -1588 -2205 -1554 -2171
rect -1496 -2205 -1462 -2171
rect -1404 -2205 -1370 -2171
rect -1312 -2205 -1278 -2171
rect -1220 -2205 -1186 -2171
rect -1128 -2205 -1094 -2171
rect -1036 -2205 -1002 -2171
rect -944 -2205 -910 -2171
rect -852 -2205 -818 -2171
rect -760 -2205 -726 -2171
rect -668 -2205 -634 -2171
rect -576 -2205 -542 -2171
rect -484 -2205 -450 -2171
rect -392 -2205 -358 -2171
rect -300 -2205 -266 -2171
rect -208 -2205 -174 -2171
rect -116 -2205 -82 -2171
rect -24 -2205 10 -2171
rect 68 -2205 102 -2171
rect 160 -2205 194 -2171
rect 252 -2205 286 -2171
rect 344 -2205 378 -2171
rect 436 -2205 470 -2171
rect 528 -2205 562 -2171
rect 620 -2205 654 -2171
rect 712 -2205 746 -2171
rect 804 -2205 838 -2171
rect 896 -2205 930 -2171
rect 988 -2205 1022 -2171
rect 1080 -2205 1114 -2171
rect 1172 -2205 1206 -2171
rect 1264 -2205 1298 -2171
rect 1356 -2205 1390 -2171
rect 1448 -2205 1482 -2171
rect 1540 -2205 1574 -2171
rect 1632 -2205 1666 -2171
rect 1724 -2205 1758 -2171
rect 1816 -2205 1850 -2171
rect 1908 -2205 1942 -2171
rect 2000 -2205 2034 -2171
rect 2092 -2205 2126 -2171
rect 2184 -2205 2218 -2171
rect 2276 -2205 2310 -2171
rect 2368 -2205 2402 -2171
rect 2460 -2205 2494 -2171
rect 2552 -2205 2586 -2171
rect 2644 -2205 2678 -2171
rect 2736 -2205 2770 -2171
rect 2828 -2205 2862 -2171
rect 2920 -2205 2954 -2171
rect 3012 -2205 3046 -2171
rect 3104 -2205 3138 -2171
rect 3196 -2205 3230 -2171
rect 3288 -2205 3322 -2171
rect 3380 -2205 3414 -2171
rect 3472 -2205 3506 -2171
rect 3564 -2205 3598 -2171
rect 3656 -2205 3690 -2171
rect 3748 -2205 3782 -2171
rect 3840 -2205 3874 -2171
rect 3932 -2205 3966 -2171
rect 4024 -2205 4058 -2171
rect 4116 -2205 4150 -2171
rect 4208 -2205 4242 -2171
rect 4300 -2205 4334 -2171
rect 4392 -2205 4426 -2171
rect 4484 -2205 4518 -2171
rect 4576 -2205 4610 -2171
rect 4668 -2205 4702 -2171
rect 4760 -2205 4794 -2171
rect 4852 -2205 4886 -2171
rect 4944 -2205 4978 -2171
rect 5036 -2205 5070 -2171
rect 5128 -2205 5162 -2171
rect 5220 -2205 5254 -2171
rect 5312 -2205 5346 -2171
rect 5404 -2205 5438 -2171
rect 5496 -2205 5530 -2171
rect 5588 -2205 5622 -2171
rect 5680 -2205 5714 -2171
rect 5772 -2205 5806 -2171
rect 5864 -2205 5898 -2171
rect 5956 -2205 5990 -2171
rect 6048 -2205 6082 -2171
rect 6140 -2205 6174 -2171
rect 6232 -2205 6266 -2171
rect 6324 -2205 6358 -2171
rect 6416 -2205 6450 -2171
rect 6508 -2205 6542 -2171
rect 6600 -2205 6634 -2171
rect 6692 -2205 6726 -2171
rect 6784 -2205 6818 -2171
rect 6876 -2205 6910 -2171
rect 6968 -2205 7002 -2171
rect 7060 -2205 7094 -2171
rect 7152 -2205 7186 -2171
rect 7244 -2205 7278 -2171
rect 7336 -2205 7370 -2171
rect 7428 -2205 7462 -2171
rect 7520 -2205 7554 -2171
rect 7612 -2205 7646 -2171
rect 7704 -2205 7738 -2171
rect 7796 -2205 7830 -2171
rect 7888 -2205 7922 -2171
rect 7980 -2205 8014 -2171
rect 8072 -2205 8106 -2171
rect 8164 -2205 8198 -2171
rect 8256 -2205 8290 -2171
rect 8348 -2205 8382 -2171
rect 8440 -2205 8474 -2171
rect 8532 -2205 8566 -2171
rect 8624 -2205 8658 -2171
rect 8716 -2205 8750 -2171
rect 8808 -2205 8842 -2171
rect 8900 -2205 8934 -2171
rect 8992 -2205 9026 -2171
rect 9084 -2205 9118 -2171
rect 9176 -2205 9210 -2171
rect 9268 -2205 9302 -2171
rect 9360 -2205 9394 -2171
rect 9452 -2205 9486 -2171
rect 9544 -2205 9578 -2171
rect 9636 -2205 9670 -2171
rect 9728 -2205 9762 -2171
rect 9820 -2205 9854 -2171
rect 9912 -2205 9946 -2171
rect 10004 -2205 10038 -2171
rect 10096 -2205 10130 -2171
rect 10188 -2205 10222 -2171
rect 10280 -2205 10314 -2171
rect 10372 -2205 10406 -2171
rect 10464 -2205 10498 -2171
rect 10556 -2205 10590 -2171
rect 10648 -2205 10682 -2171
rect 10740 -2205 10774 -2171
rect 10832 -2205 10866 -2171
rect 10924 -2205 10958 -2171
rect 11016 -2205 11050 -2171
rect 11108 -2205 11142 -2171
rect 11200 -2205 11234 -2171
rect 11292 -2205 11326 -2171
rect 11384 -2205 11418 -2171
rect 11476 -2205 11510 -2171
rect 11568 -2205 11602 -2171
rect 11660 -2205 11694 -2171
rect 11752 -2205 11786 -2171
rect 11844 -2205 11878 -2171
rect 11936 -2205 11970 -2171
rect 12028 -2205 12062 -2171
rect 12120 -2205 12154 -2171
rect 12212 -2205 12246 -2171
rect 12304 -2205 12338 -2171
rect 12396 -2205 12430 -2171
rect 12488 -2205 12522 -2171
rect 12580 -2205 12614 -2171
rect 12672 -2205 12706 -2171
rect 12764 -2205 12798 -2171
rect 12856 -2205 12890 -2171
rect 12948 -2205 12982 -2171
rect 13040 -2205 13074 -2171
rect 13132 -2205 13166 -2171
rect 13224 -2205 13258 -2171
rect 13316 -2205 13350 -2171
rect 13408 -2205 13442 -2171
rect 13500 -2205 13534 -2171
rect 13592 -2205 13626 -2171
rect 13684 -2205 13718 -2171
rect 13776 -2205 13810 -2171
rect 13868 -2205 13902 -2171
rect 13960 -2205 13994 -2171
rect 14052 -2205 14086 -2171
rect 14144 -2205 14178 -2171
rect 14236 -2205 14270 -2171
rect 14328 -2205 14362 -2171
rect 14420 -2205 14454 -2171
rect 14512 -2205 14546 -2171
rect 14604 -2205 14638 -2171
rect 14696 -2205 14730 -2171
rect 14788 -2205 14822 -2171
rect 14880 -2205 14914 -2171
rect 14972 -2205 15006 -2171
rect 15064 -2205 15098 -2171
rect 15156 -2205 15190 -2171
rect 15248 -2205 15282 -2171
rect 15340 -2205 15374 -2171
rect 15432 -2205 15466 -2171
rect 15524 -2205 15558 -2171
rect 15616 -2205 15650 -2171
rect 15708 -2205 15742 -2171
rect 15800 -2205 15834 -2171
rect 15892 -2205 15926 -2171
rect 15984 -2205 16018 -2171
rect 16076 -2205 16110 -2171
rect 16168 -2205 16202 -2171
rect 16260 -2205 16294 -2171
rect 16352 -2205 16386 -2171
rect 16444 -2205 16478 -2171
rect 16536 -2205 16570 -2171
rect 16628 -2205 16662 -2171
rect 436 -2483 470 -2480
rect 436 -2514 464 -2483
rect 464 -2514 470 -2483
rect 1081 -2512 1115 -2478
rect 3041 -2483 3075 -2478
rect 3041 -2512 3074 -2483
rect 3074 -2512 3075 -2483
rect 3655 -2512 3689 -2478
rect 5615 -2483 5649 -2478
rect 5615 -2512 5616 -2483
rect 5616 -2512 5649 -2483
rect 6229 -2512 6263 -2478
rect 8189 -2483 8223 -2478
rect 8189 -2512 8192 -2483
rect 8192 -2512 8223 -2483
rect 8806 -2512 8840 -2478
rect 10763 -2483 10797 -2478
rect 10763 -2512 10768 -2483
rect 10768 -2512 10797 -2483
rect 11386 -2479 11420 -2445
rect 12480 -2441 12514 -2407
rect 12480 -2515 12514 -2481
rect 12568 -2483 12602 -2479
rect 12659 -2483 12693 -2479
rect 12765 -2483 12799 -2479
rect 12858 -2483 12892 -2477
rect 12942 -2483 12976 -2477
rect 12568 -2513 12574 -2483
rect 12574 -2513 12602 -2483
rect 12659 -2513 12676 -2483
rect 12676 -2513 12693 -2483
rect 12765 -2513 12778 -2483
rect 12778 -2513 12799 -2483
rect 12858 -2511 12880 -2483
rect 12880 -2511 12892 -2483
rect 12942 -2511 12948 -2483
rect 12948 -2511 12976 -2483
rect 13039 -2500 13073 -2466
rect 12480 -2587 12514 -2553
rect 13042 -2577 13076 -2543
rect 15248 -2460 15282 -2426
rect 15340 -2460 15374 -2426
rect 13685 -2517 13692 -2510
rect 13692 -2517 13719 -2510
rect 13685 -2544 13719 -2517
rect 15248 -2556 15282 -2522
rect 15341 -2556 15375 -2522
rect -2968 -2749 -2934 -2715
rect -2876 -2749 -2842 -2715
rect -2784 -2749 -2750 -2715
rect -2692 -2749 -2658 -2715
rect -2600 -2749 -2566 -2715
rect -2508 -2749 -2474 -2715
rect -2416 -2749 -2382 -2715
rect -2324 -2749 -2290 -2715
rect -2232 -2749 -2198 -2715
rect -2140 -2749 -2106 -2715
rect -2048 -2749 -2014 -2715
rect -1956 -2749 -1922 -2715
rect -1864 -2749 -1830 -2715
rect -1772 -2749 -1738 -2715
rect -1680 -2749 -1646 -2715
rect -1588 -2749 -1554 -2715
rect -1496 -2749 -1462 -2715
rect -1404 -2749 -1370 -2715
rect -1312 -2749 -1278 -2715
rect -1220 -2749 -1186 -2715
rect -1128 -2749 -1094 -2715
rect -1036 -2749 -1002 -2715
rect -944 -2749 -910 -2715
rect -852 -2749 -818 -2715
rect -760 -2749 -726 -2715
rect -668 -2749 -634 -2715
rect -576 -2749 -542 -2715
rect -484 -2749 -450 -2715
rect -392 -2749 -358 -2715
rect -300 -2749 -266 -2715
rect -208 -2749 -174 -2715
rect -116 -2749 -82 -2715
rect -24 -2749 10 -2715
rect 68 -2749 102 -2715
rect 160 -2749 194 -2715
rect 252 -2749 286 -2715
rect 344 -2749 378 -2715
rect 436 -2749 470 -2715
rect 528 -2749 562 -2715
rect 620 -2749 654 -2715
rect 712 -2749 746 -2715
rect 804 -2749 838 -2715
rect 896 -2749 930 -2715
rect 988 -2749 1022 -2715
rect 1080 -2749 1114 -2715
rect 1172 -2749 1206 -2715
rect 1264 -2749 1298 -2715
rect 1356 -2749 1390 -2715
rect 1448 -2749 1482 -2715
rect 1540 -2749 1574 -2715
rect 1632 -2749 1666 -2715
rect 1724 -2749 1758 -2715
rect 1816 -2749 1850 -2715
rect 1908 -2749 1942 -2715
rect 2000 -2749 2034 -2715
rect 2092 -2749 2126 -2715
rect 2184 -2749 2218 -2715
rect 2276 -2749 2310 -2715
rect 2368 -2749 2402 -2715
rect 2460 -2749 2494 -2715
rect 2552 -2749 2586 -2715
rect 2644 -2749 2678 -2715
rect 2736 -2749 2770 -2715
rect 2828 -2749 2862 -2715
rect 2920 -2749 2954 -2715
rect 3012 -2749 3046 -2715
rect 3104 -2749 3138 -2715
rect 3196 -2749 3230 -2715
rect 3288 -2749 3322 -2715
rect 3380 -2749 3414 -2715
rect 3472 -2749 3506 -2715
rect 3564 -2749 3598 -2715
rect 3656 -2749 3690 -2715
rect 3748 -2749 3782 -2715
rect 3840 -2749 3874 -2715
rect 3932 -2749 3966 -2715
rect 4024 -2749 4058 -2715
rect 4116 -2749 4150 -2715
rect 4208 -2749 4242 -2715
rect 4300 -2749 4334 -2715
rect 4392 -2749 4426 -2715
rect 4484 -2749 4518 -2715
rect 4576 -2749 4610 -2715
rect 4668 -2749 4702 -2715
rect 4760 -2749 4794 -2715
rect 4852 -2749 4886 -2715
rect 4944 -2749 4978 -2715
rect 5036 -2749 5070 -2715
rect 5128 -2749 5162 -2715
rect 5220 -2749 5254 -2715
rect 5312 -2749 5346 -2715
rect 5404 -2749 5438 -2715
rect 5496 -2749 5530 -2715
rect 5588 -2749 5622 -2715
rect 5680 -2749 5714 -2715
rect 5772 -2749 5806 -2715
rect 5864 -2749 5898 -2715
rect 5956 -2749 5990 -2715
rect 6048 -2749 6082 -2715
rect 6140 -2749 6174 -2715
rect 6232 -2749 6266 -2715
rect 6324 -2749 6358 -2715
rect 6416 -2749 6450 -2715
rect 6508 -2749 6542 -2715
rect 6600 -2749 6634 -2715
rect 6692 -2749 6726 -2715
rect 6784 -2749 6818 -2715
rect 6876 -2749 6910 -2715
rect 6968 -2749 7002 -2715
rect 7060 -2749 7094 -2715
rect 7152 -2749 7186 -2715
rect 7244 -2749 7278 -2715
rect 7336 -2749 7370 -2715
rect 7428 -2749 7462 -2715
rect 7520 -2749 7554 -2715
rect 7612 -2749 7646 -2715
rect 7704 -2749 7738 -2715
rect 7796 -2749 7830 -2715
rect 7888 -2749 7922 -2715
rect 7980 -2749 8014 -2715
rect 8072 -2749 8106 -2715
rect 8164 -2749 8198 -2715
rect 8256 -2749 8290 -2715
rect 8348 -2749 8382 -2715
rect 8440 -2749 8474 -2715
rect 8532 -2749 8566 -2715
rect 8624 -2749 8658 -2715
rect 8716 -2749 8750 -2715
rect 8808 -2749 8842 -2715
rect 8900 -2749 8934 -2715
rect 8992 -2749 9026 -2715
rect 9084 -2749 9118 -2715
rect 9176 -2749 9210 -2715
rect 9268 -2749 9302 -2715
rect 9360 -2749 9394 -2715
rect 9452 -2749 9486 -2715
rect 9544 -2749 9578 -2715
rect 9636 -2749 9670 -2715
rect 9728 -2749 9762 -2715
rect 9820 -2749 9854 -2715
rect 9912 -2749 9946 -2715
rect 10004 -2749 10038 -2715
rect 10096 -2749 10130 -2715
rect 10188 -2749 10222 -2715
rect 10280 -2749 10314 -2715
rect 10372 -2749 10406 -2715
rect 10464 -2749 10498 -2715
rect 10556 -2749 10590 -2715
rect 10648 -2749 10682 -2715
rect 10740 -2749 10774 -2715
rect 10832 -2749 10866 -2715
rect 10924 -2749 10958 -2715
rect 11016 -2749 11050 -2715
rect 11108 -2749 11142 -2715
rect 11200 -2749 11234 -2715
rect 11292 -2749 11326 -2715
rect 11384 -2749 11418 -2715
rect 11476 -2749 11510 -2715
rect 11568 -2749 11602 -2715
rect 11660 -2749 11694 -2715
rect 11752 -2749 11786 -2715
rect 11844 -2749 11878 -2715
rect 11936 -2749 11970 -2715
rect 12028 -2749 12062 -2715
rect 12120 -2749 12154 -2715
rect 12212 -2749 12246 -2715
rect 12304 -2749 12338 -2715
rect 12396 -2749 12430 -2715
rect 12488 -2749 12522 -2715
rect 12580 -2749 12614 -2715
rect 12672 -2749 12706 -2715
rect 12764 -2749 12798 -2715
rect 12856 -2749 12890 -2715
rect 12948 -2749 12982 -2715
rect 13040 -2749 13074 -2715
rect 13132 -2749 13166 -2715
rect 13224 -2749 13258 -2715
rect 13316 -2749 13350 -2715
rect 13408 -2749 13442 -2715
rect 13500 -2749 13534 -2715
rect 13592 -2749 13626 -2715
rect 13684 -2749 13718 -2715
rect 13776 -2749 13810 -2715
rect 13868 -2749 13902 -2715
rect 13960 -2749 13994 -2715
rect 14052 -2749 14086 -2715
rect 14144 -2749 14178 -2715
rect 14236 -2749 14270 -2715
rect 14328 -2749 14362 -2715
rect 14420 -2749 14454 -2715
rect 14512 -2749 14546 -2715
rect 14604 -2749 14638 -2715
rect 14696 -2749 14730 -2715
rect 14788 -2749 14822 -2715
rect 14880 -2749 14914 -2715
rect 14972 -2749 15006 -2715
rect 15064 -2749 15098 -2715
rect 15156 -2749 15190 -2715
rect 15248 -2749 15282 -2715
rect 15340 -2749 15374 -2715
rect 15432 -2749 15466 -2715
rect 15524 -2749 15558 -2715
rect 15616 -2749 15650 -2715
rect 15708 -2749 15742 -2715
rect 15800 -2749 15834 -2715
rect 15892 -2749 15926 -2715
rect 15984 -2749 16018 -2715
rect 16076 -2749 16110 -2715
rect 16168 -2749 16202 -2715
rect 16260 -2749 16294 -2715
rect 16352 -2749 16386 -2715
rect 16444 -2749 16478 -2715
rect 16536 -2749 16570 -2715
rect 16628 -2749 16662 -2715
rect -1960 -2981 -1954 -2952
rect -1954 -2981 -1926 -2952
rect -1960 -2986 -1926 -2981
rect -1783 -2949 -1749 -2915
rect 429 -3021 463 -2987
rect 1072 -2981 1086 -2952
rect 1086 -2981 1106 -2952
rect 1072 -2986 1106 -2981
rect 3016 -2987 3050 -2953
rect 3630 -2981 3662 -2953
rect 3662 -2981 3664 -2953
rect 3630 -2987 3664 -2981
rect 5590 -2987 5624 -2953
rect 6204 -2981 6238 -2953
rect 6204 -2987 6238 -2981
rect 8164 -2987 8198 -2953
rect 8778 -2981 8780 -2953
rect 8780 -2981 8812 -2953
rect 8778 -2987 8812 -2981
rect 10738 -2988 10772 -2954
rect 11384 -2981 11390 -2952
rect 11390 -2981 11418 -2952
rect 11384 -2986 11418 -2981
rect -2968 -3293 -2934 -3259
rect -2876 -3293 -2842 -3259
rect -2784 -3293 -2750 -3259
rect -2692 -3293 -2658 -3259
rect -2600 -3293 -2566 -3259
rect -2508 -3293 -2474 -3259
rect -2416 -3293 -2382 -3259
rect -2324 -3293 -2290 -3259
rect -2232 -3293 -2198 -3259
rect -2140 -3293 -2106 -3259
rect -2048 -3293 -2014 -3259
rect -1956 -3293 -1922 -3259
rect -1864 -3293 -1830 -3259
rect -1772 -3293 -1738 -3259
rect -1680 -3293 -1646 -3259
rect -1588 -3293 -1554 -3259
rect -1496 -3293 -1462 -3259
rect -1404 -3293 -1370 -3259
rect -1312 -3293 -1278 -3259
rect -1220 -3293 -1186 -3259
rect -1128 -3293 -1094 -3259
rect -1036 -3293 -1002 -3259
rect -944 -3293 -910 -3259
rect -852 -3293 -818 -3259
rect -760 -3293 -726 -3259
rect -668 -3293 -634 -3259
rect -576 -3293 -542 -3259
rect -484 -3293 -450 -3259
rect -392 -3293 -358 -3259
rect -300 -3293 -266 -3259
rect -208 -3293 -174 -3259
rect -116 -3293 -82 -3259
rect -24 -3293 10 -3259
rect 68 -3293 102 -3259
rect 160 -3293 194 -3259
rect 252 -3293 286 -3259
rect 344 -3293 378 -3259
rect 436 -3293 470 -3259
rect 528 -3293 562 -3259
rect 620 -3293 654 -3259
rect 712 -3293 746 -3259
rect 804 -3293 838 -3259
rect 896 -3293 930 -3259
rect 988 -3293 1022 -3259
rect 1080 -3293 1114 -3259
rect 1172 -3293 1206 -3259
rect 1264 -3293 1298 -3259
rect 1356 -3293 1390 -3259
rect 1448 -3293 1482 -3259
rect 1540 -3293 1574 -3259
rect 1632 -3293 1666 -3259
rect 1724 -3293 1758 -3259
rect 1816 -3293 1850 -3259
rect 1908 -3293 1942 -3259
rect 2000 -3293 2034 -3259
rect 2092 -3293 2126 -3259
rect 2184 -3293 2218 -3259
rect 2276 -3293 2310 -3259
rect 2368 -3293 2402 -3259
rect 2460 -3293 2494 -3259
rect 2552 -3293 2586 -3259
rect 2644 -3293 2678 -3259
rect 2736 -3293 2770 -3259
rect 2828 -3293 2862 -3259
rect 2920 -3293 2954 -3259
rect 3012 -3293 3046 -3259
rect 3104 -3293 3138 -3259
rect 3196 -3293 3230 -3259
rect 3288 -3293 3322 -3259
rect 3380 -3293 3414 -3259
rect 3472 -3293 3506 -3259
rect 3564 -3293 3598 -3259
rect 3656 -3293 3690 -3259
rect 3748 -3293 3782 -3259
rect 3840 -3293 3874 -3259
rect 3932 -3293 3966 -3259
rect 4024 -3293 4058 -3259
rect 4116 -3293 4150 -3259
rect 4208 -3293 4242 -3259
rect 4300 -3293 4334 -3259
rect 4392 -3293 4426 -3259
rect 4484 -3293 4518 -3259
rect 4576 -3293 4610 -3259
rect 4668 -3293 4702 -3259
rect 4760 -3293 4794 -3259
rect 4852 -3293 4886 -3259
rect 4944 -3293 4978 -3259
rect 5036 -3293 5070 -3259
rect 5128 -3293 5162 -3259
rect 5220 -3293 5254 -3259
rect 5312 -3293 5346 -3259
rect 5404 -3293 5438 -3259
rect 5496 -3293 5530 -3259
rect 5588 -3293 5622 -3259
rect 5680 -3293 5714 -3259
rect 5772 -3293 5806 -3259
rect 5864 -3293 5898 -3259
rect 5956 -3293 5990 -3259
rect 6048 -3293 6082 -3259
rect 6140 -3293 6174 -3259
rect 6232 -3293 6266 -3259
rect 6324 -3293 6358 -3259
rect 6416 -3293 6450 -3259
rect 6508 -3293 6542 -3259
rect 6600 -3293 6634 -3259
rect 6692 -3293 6726 -3259
rect 6784 -3293 6818 -3259
rect 6876 -3293 6910 -3259
rect 6968 -3293 7002 -3259
rect 7060 -3293 7094 -3259
rect 7152 -3293 7186 -3259
rect 7244 -3293 7278 -3259
rect 7336 -3293 7370 -3259
rect 7428 -3293 7462 -3259
rect 7520 -3293 7554 -3259
rect 7612 -3293 7646 -3259
rect 7704 -3293 7738 -3259
rect 7796 -3293 7830 -3259
rect 7888 -3293 7922 -3259
rect 7980 -3293 8014 -3259
rect 8072 -3293 8106 -3259
rect 8164 -3293 8198 -3259
rect 8256 -3293 8290 -3259
rect 8348 -3293 8382 -3259
rect 8440 -3293 8474 -3259
rect 8532 -3293 8566 -3259
rect 8624 -3293 8658 -3259
rect 8716 -3293 8750 -3259
rect 8808 -3293 8842 -3259
rect 8900 -3293 8934 -3259
rect 8992 -3293 9026 -3259
rect 9084 -3293 9118 -3259
rect 9176 -3293 9210 -3259
rect 9268 -3293 9302 -3259
rect 9360 -3293 9394 -3259
rect 9452 -3293 9486 -3259
rect 9544 -3293 9578 -3259
rect 9636 -3293 9670 -3259
rect 9728 -3293 9762 -3259
rect 9820 -3293 9854 -3259
rect 9912 -3293 9946 -3259
rect 10004 -3293 10038 -3259
rect 10096 -3293 10130 -3259
rect 10188 -3293 10222 -3259
rect 10280 -3293 10314 -3259
rect 10372 -3293 10406 -3259
rect 10464 -3293 10498 -3259
rect 10556 -3293 10590 -3259
rect 10648 -3293 10682 -3259
rect 10740 -3293 10774 -3259
rect 10832 -3293 10866 -3259
rect 10924 -3293 10958 -3259
rect 11016 -3293 11050 -3259
rect 11108 -3293 11142 -3259
rect 11200 -3293 11234 -3259
rect 11292 -3293 11326 -3259
rect 11384 -3293 11418 -3259
rect 11476 -3293 11510 -3259
rect 11568 -3293 11602 -3259
rect 11660 -3293 11694 -3259
rect 11752 -3293 11786 -3259
rect 11844 -3293 11878 -3259
rect 11936 -3293 11970 -3259
rect 12028 -3293 12062 -3259
rect 12120 -3293 12154 -3259
rect 12212 -3293 12246 -3259
rect 12304 -3293 12338 -3259
rect 12396 -3293 12430 -3259
rect 12488 -3293 12522 -3259
rect 12580 -3293 12614 -3259
rect 12672 -3293 12706 -3259
rect 12764 -3293 12798 -3259
rect 12856 -3293 12890 -3259
rect 12948 -3293 12982 -3259
rect 13040 -3293 13074 -3259
rect 13132 -3293 13166 -3259
rect 13224 -3293 13258 -3259
rect 13316 -3293 13350 -3259
rect 13408 -3293 13442 -3259
rect 13500 -3293 13534 -3259
rect 13592 -3293 13626 -3259
rect 13684 -3293 13718 -3259
rect 13776 -3293 13810 -3259
rect 13868 -3293 13902 -3259
rect 13960 -3293 13994 -3259
rect 14052 -3293 14086 -3259
rect 14144 -3293 14178 -3259
rect 14236 -3293 14270 -3259
rect 14328 -3293 14362 -3259
rect 14420 -3293 14454 -3259
rect 14512 -3293 14546 -3259
rect 14604 -3293 14638 -3259
rect 14696 -3293 14730 -3259
rect 14788 -3293 14822 -3259
rect 14880 -3293 14914 -3259
rect 14972 -3293 15006 -3259
rect 15064 -3293 15098 -3259
rect 15156 -3293 15190 -3259
rect 15248 -3293 15282 -3259
rect 15340 -3293 15374 -3259
rect 15432 -3293 15466 -3259
rect 15524 -3293 15558 -3259
rect 15616 -3293 15650 -3259
rect 15708 -3293 15742 -3259
rect 15800 -3293 15834 -3259
rect 15892 -3293 15926 -3259
rect 15984 -3293 16018 -3259
rect 16076 -3293 16110 -3259
rect 16168 -3293 16202 -3259
rect 16260 -3293 16294 -3259
rect 16352 -3293 16386 -3259
rect 16444 -3293 16478 -3259
rect 16536 -3293 16570 -3259
rect 16628 -3293 16662 -3259
rect 432 -3565 466 -3531
rect 1070 -3571 1104 -3568
rect 1070 -3602 1086 -3571
rect 1086 -3602 1104 -3571
rect 3016 -3599 3050 -3565
rect 3630 -3571 3664 -3565
rect 3630 -3599 3662 -3571
rect 3662 -3599 3664 -3571
rect 5590 -3599 5624 -3565
rect 6204 -3571 6238 -3565
rect 6204 -3599 6238 -3571
rect 8164 -3599 8198 -3565
rect 8778 -3571 8812 -3565
rect 8778 -3599 8780 -3571
rect 8780 -3599 8812 -3571
rect 10735 -3602 10769 -3568
rect 11383 -3571 11417 -3567
rect 11383 -3601 11390 -3571
rect 11390 -3601 11417 -3571
rect -2968 -3837 -2934 -3803
rect -2876 -3837 -2842 -3803
rect -2784 -3837 -2750 -3803
rect -2692 -3837 -2658 -3803
rect -2600 -3837 -2566 -3803
rect -2508 -3837 -2474 -3803
rect -2416 -3837 -2382 -3803
rect -2324 -3837 -2290 -3803
rect -2232 -3837 -2198 -3803
rect -2140 -3837 -2106 -3803
rect -2048 -3837 -2014 -3803
rect -1956 -3837 -1922 -3803
rect -1864 -3837 -1830 -3803
rect -1772 -3837 -1738 -3803
rect -1680 -3837 -1646 -3803
rect -1588 -3837 -1554 -3803
rect -1496 -3837 -1462 -3803
rect -1404 -3837 -1370 -3803
rect -1312 -3837 -1278 -3803
rect -1220 -3837 -1186 -3803
rect -1128 -3837 -1094 -3803
rect -1036 -3837 -1002 -3803
rect -944 -3837 -910 -3803
rect -852 -3837 -818 -3803
rect -760 -3837 -726 -3803
rect -668 -3837 -634 -3803
rect -576 -3837 -542 -3803
rect -484 -3837 -450 -3803
rect -392 -3837 -358 -3803
rect -300 -3837 -266 -3803
rect -208 -3837 -174 -3803
rect -116 -3837 -82 -3803
rect -24 -3837 10 -3803
rect 68 -3837 102 -3803
rect 160 -3837 194 -3803
rect 252 -3837 286 -3803
rect 344 -3837 378 -3803
rect 436 -3837 470 -3803
rect 528 -3837 562 -3803
rect 620 -3837 654 -3803
rect 712 -3837 746 -3803
rect 804 -3837 838 -3803
rect 896 -3837 930 -3803
rect 988 -3837 1022 -3803
rect 1080 -3837 1114 -3803
rect 1172 -3837 1206 -3803
rect 1264 -3837 1298 -3803
rect 1356 -3837 1390 -3803
rect 1448 -3837 1482 -3803
rect 1540 -3837 1574 -3803
rect 1632 -3837 1666 -3803
rect 1724 -3837 1758 -3803
rect 1816 -3837 1850 -3803
rect 1908 -3837 1942 -3803
rect 2000 -3837 2034 -3803
rect 2092 -3837 2126 -3803
rect 2184 -3837 2218 -3803
rect 2276 -3837 2310 -3803
rect 2368 -3837 2402 -3803
rect 2460 -3837 2494 -3803
rect 2552 -3837 2586 -3803
rect 2644 -3837 2678 -3803
rect 2736 -3837 2770 -3803
rect 2828 -3837 2862 -3803
rect 2920 -3837 2954 -3803
rect 3012 -3837 3046 -3803
rect 3104 -3837 3138 -3803
rect 3196 -3837 3230 -3803
rect 3288 -3837 3322 -3803
rect 3380 -3837 3414 -3803
rect 3472 -3837 3506 -3803
rect 3564 -3837 3598 -3803
rect 3656 -3837 3690 -3803
rect 3748 -3837 3782 -3803
rect 3840 -3837 3874 -3803
rect 3932 -3837 3966 -3803
rect 4024 -3837 4058 -3803
rect 4116 -3837 4150 -3803
rect 4208 -3837 4242 -3803
rect 4300 -3837 4334 -3803
rect 4392 -3837 4426 -3803
rect 4484 -3837 4518 -3803
rect 4576 -3837 4610 -3803
rect 4668 -3837 4702 -3803
rect 4760 -3837 4794 -3803
rect 4852 -3837 4886 -3803
rect 4944 -3837 4978 -3803
rect 5036 -3837 5070 -3803
rect 5128 -3837 5162 -3803
rect 5220 -3837 5254 -3803
rect 5312 -3837 5346 -3803
rect 5404 -3837 5438 -3803
rect 5496 -3837 5530 -3803
rect 5588 -3837 5622 -3803
rect 5680 -3837 5714 -3803
rect 5772 -3837 5806 -3803
rect 5864 -3837 5898 -3803
rect 5956 -3837 5990 -3803
rect 6048 -3837 6082 -3803
rect 6140 -3837 6174 -3803
rect 6232 -3837 6266 -3803
rect 6324 -3837 6358 -3803
rect 6416 -3837 6450 -3803
rect 6508 -3837 6542 -3803
rect 6600 -3837 6634 -3803
rect 6692 -3837 6726 -3803
rect 6784 -3837 6818 -3803
rect 6876 -3837 6910 -3803
rect 6968 -3837 7002 -3803
rect 7060 -3837 7094 -3803
rect 7152 -3837 7186 -3803
rect 7244 -3837 7278 -3803
rect 7336 -3837 7370 -3803
rect 7428 -3837 7462 -3803
rect 7520 -3837 7554 -3803
rect 7612 -3837 7646 -3803
rect 7704 -3837 7738 -3803
rect 7796 -3837 7830 -3803
rect 7888 -3837 7922 -3803
rect 7980 -3837 8014 -3803
rect 8072 -3837 8106 -3803
rect 8164 -3837 8198 -3803
rect 8256 -3837 8290 -3803
rect 8348 -3837 8382 -3803
rect 8440 -3837 8474 -3803
rect 8532 -3837 8566 -3803
rect 8624 -3837 8658 -3803
rect 8716 -3837 8750 -3803
rect 8808 -3837 8842 -3803
rect 8900 -3837 8934 -3803
rect 8992 -3837 9026 -3803
rect 9084 -3837 9118 -3803
rect 9176 -3837 9210 -3803
rect 9268 -3837 9302 -3803
rect 9360 -3837 9394 -3803
rect 9452 -3837 9486 -3803
rect 9544 -3837 9578 -3803
rect 9636 -3837 9670 -3803
rect 9728 -3837 9762 -3803
rect 9820 -3837 9854 -3803
rect 9912 -3837 9946 -3803
rect 10004 -3837 10038 -3803
rect 10096 -3837 10130 -3803
rect 10188 -3837 10222 -3803
rect 10280 -3837 10314 -3803
rect 10372 -3837 10406 -3803
rect 10464 -3837 10498 -3803
rect 10556 -3837 10590 -3803
rect 10648 -3837 10682 -3803
rect 10740 -3837 10774 -3803
rect 10832 -3837 10866 -3803
rect 10924 -3837 10958 -3803
rect 11016 -3837 11050 -3803
rect 11108 -3837 11142 -3803
rect 11200 -3837 11234 -3803
rect 11292 -3837 11326 -3803
rect 11384 -3837 11418 -3803
rect 11476 -3837 11510 -3803
rect 11568 -3837 11602 -3803
rect 11660 -3837 11694 -3803
rect 11752 -3837 11786 -3803
rect 11844 -3837 11878 -3803
rect 11936 -3837 11970 -3803
rect 12028 -3837 12062 -3803
rect 12120 -3837 12154 -3803
rect 12212 -3837 12246 -3803
rect 12304 -3837 12338 -3803
rect 12396 -3837 12430 -3803
rect 12488 -3837 12522 -3803
rect 12580 -3837 12614 -3803
rect 12672 -3837 12706 -3803
rect 12764 -3837 12798 -3803
rect 12856 -3837 12890 -3803
rect 12948 -3837 12982 -3803
rect 13040 -3837 13074 -3803
rect 13132 -3837 13166 -3803
rect 13224 -3837 13258 -3803
rect 13316 -3837 13350 -3803
rect 13408 -3837 13442 -3803
rect 13500 -3837 13534 -3803
rect 13592 -3837 13626 -3803
rect 13684 -3837 13718 -3803
rect 13776 -3837 13810 -3803
rect 13868 -3837 13902 -3803
rect 13960 -3837 13994 -3803
rect 14052 -3837 14086 -3803
rect 14144 -3837 14178 -3803
rect 14236 -3837 14270 -3803
rect 14328 -3837 14362 -3803
rect 14420 -3837 14454 -3803
rect 14512 -3837 14546 -3803
rect 14604 -3837 14638 -3803
rect 14696 -3837 14730 -3803
rect 14788 -3837 14822 -3803
rect 14880 -3837 14914 -3803
rect 14972 -3837 15006 -3803
rect 15064 -3837 15098 -3803
rect 15156 -3837 15190 -3803
rect 15248 -3837 15282 -3803
rect 15340 -3837 15374 -3803
rect 15432 -3837 15466 -3803
rect 15524 -3837 15558 -3803
rect 15616 -3837 15650 -3803
rect 15708 -3837 15742 -3803
rect 15800 -3837 15834 -3803
rect 15892 -3837 15926 -3803
rect 15984 -3837 16018 -3803
rect 16076 -3837 16110 -3803
rect 16168 -3837 16202 -3803
rect 16260 -3837 16294 -3803
rect 16352 -3837 16386 -3803
rect 16444 -3837 16478 -3803
rect 16536 -3837 16570 -3803
rect 16628 -3837 16662 -3803
rect 436 -4069 464 -4040
rect 464 -4069 470 -4040
rect 436 -4074 470 -4069
rect 1081 -4074 1115 -4040
rect 3041 -4069 3074 -4040
rect 3074 -4069 3075 -4040
rect 3041 -4074 3075 -4069
rect 3655 -4074 3689 -4040
rect 5615 -4069 5616 -4040
rect 5616 -4069 5649 -4040
rect 5615 -4074 5649 -4069
rect 6229 -4074 6263 -4040
rect 8189 -4069 8192 -4040
rect 8192 -4069 8223 -4040
rect 8189 -4074 8223 -4069
rect 8806 -4074 8840 -4040
rect 10763 -4069 10768 -4040
rect 10768 -4069 10797 -4040
rect 10763 -4074 10797 -4069
rect 11386 -4111 11420 -4077
rect 12480 -3999 12514 -3965
rect 13042 -4009 13076 -3975
rect 12480 -4071 12514 -4037
rect 12568 -4069 12574 -4039
rect 12574 -4069 12602 -4039
rect 12659 -4069 12676 -4039
rect 12676 -4069 12693 -4039
rect 12765 -4069 12778 -4039
rect 12778 -4069 12799 -4039
rect 12858 -4069 12880 -4041
rect 12880 -4069 12892 -4041
rect 12942 -4069 12948 -4041
rect 12948 -4069 12976 -4041
rect 12568 -4073 12602 -4069
rect 12659 -4073 12693 -4069
rect 12765 -4073 12799 -4069
rect 12858 -4075 12892 -4069
rect 12942 -4075 12976 -4069
rect 12480 -4145 12514 -4111
rect 13039 -4086 13073 -4052
rect 13685 -4035 13719 -4008
rect 13685 -4042 13692 -4035
rect 13692 -4042 13719 -4035
rect 15248 -4030 15282 -3996
rect 15341 -4030 15375 -3996
rect 15248 -4126 15282 -4092
rect 15340 -4126 15374 -4092
rect -2968 -4381 -2934 -4347
rect -2876 -4381 -2842 -4347
rect -2784 -4381 -2750 -4347
rect -2692 -4381 -2658 -4347
rect -2600 -4381 -2566 -4347
rect -2508 -4381 -2474 -4347
rect -2416 -4381 -2382 -4347
rect -2324 -4381 -2290 -4347
rect -2232 -4381 -2198 -4347
rect -2140 -4381 -2106 -4347
rect -2048 -4381 -2014 -4347
rect -1956 -4381 -1922 -4347
rect -1864 -4381 -1830 -4347
rect -1772 -4381 -1738 -4347
rect -1680 -4381 -1646 -4347
rect -1588 -4381 -1554 -4347
rect -1496 -4381 -1462 -4347
rect -1404 -4381 -1370 -4347
rect -1312 -4381 -1278 -4347
rect -1220 -4381 -1186 -4347
rect -1128 -4381 -1094 -4347
rect -1036 -4381 -1002 -4347
rect -944 -4381 -910 -4347
rect -852 -4381 -818 -4347
rect -760 -4381 -726 -4347
rect -668 -4381 -634 -4347
rect -576 -4381 -542 -4347
rect -484 -4381 -450 -4347
rect -392 -4381 -358 -4347
rect -300 -4381 -266 -4347
rect -208 -4381 -174 -4347
rect -116 -4381 -82 -4347
rect -24 -4381 10 -4347
rect 68 -4381 102 -4347
rect 160 -4381 194 -4347
rect 252 -4381 286 -4347
rect 344 -4381 378 -4347
rect 436 -4381 470 -4347
rect 528 -4381 562 -4347
rect 620 -4381 654 -4347
rect 712 -4381 746 -4347
rect 804 -4381 838 -4347
rect 896 -4381 930 -4347
rect 988 -4381 1022 -4347
rect 1080 -4381 1114 -4347
rect 1172 -4381 1206 -4347
rect 1264 -4381 1298 -4347
rect 1356 -4381 1390 -4347
rect 1448 -4381 1482 -4347
rect 1540 -4381 1574 -4347
rect 1632 -4381 1666 -4347
rect 1724 -4381 1758 -4347
rect 1816 -4381 1850 -4347
rect 1908 -4381 1942 -4347
rect 2000 -4381 2034 -4347
rect 2092 -4381 2126 -4347
rect 2184 -4381 2218 -4347
rect 2276 -4381 2310 -4347
rect 2368 -4381 2402 -4347
rect 2460 -4381 2494 -4347
rect 2552 -4381 2586 -4347
rect 2644 -4381 2678 -4347
rect 2736 -4381 2770 -4347
rect 2828 -4381 2862 -4347
rect 2920 -4381 2954 -4347
rect 3012 -4381 3046 -4347
rect 3104 -4381 3138 -4347
rect 3196 -4381 3230 -4347
rect 3288 -4381 3322 -4347
rect 3380 -4381 3414 -4347
rect 3472 -4381 3506 -4347
rect 3564 -4381 3598 -4347
rect 3656 -4381 3690 -4347
rect 3748 -4381 3782 -4347
rect 3840 -4381 3874 -4347
rect 3932 -4381 3966 -4347
rect 4024 -4381 4058 -4347
rect 4116 -4381 4150 -4347
rect 4208 -4381 4242 -4347
rect 4300 -4381 4334 -4347
rect 4392 -4381 4426 -4347
rect 4484 -4381 4518 -4347
rect 4576 -4381 4610 -4347
rect 4668 -4381 4702 -4347
rect 4760 -4381 4794 -4347
rect 4852 -4381 4886 -4347
rect 4944 -4381 4978 -4347
rect 5036 -4381 5070 -4347
rect 5128 -4381 5162 -4347
rect 5220 -4381 5254 -4347
rect 5312 -4381 5346 -4347
rect 5404 -4381 5438 -4347
rect 5496 -4381 5530 -4347
rect 5588 -4381 5622 -4347
rect 5680 -4381 5714 -4347
rect 5772 -4381 5806 -4347
rect 5864 -4381 5898 -4347
rect 5956 -4381 5990 -4347
rect 6048 -4381 6082 -4347
rect 6140 -4381 6174 -4347
rect 6232 -4381 6266 -4347
rect 6324 -4381 6358 -4347
rect 6416 -4381 6450 -4347
rect 6508 -4381 6542 -4347
rect 6600 -4381 6634 -4347
rect 6692 -4381 6726 -4347
rect 6784 -4381 6818 -4347
rect 6876 -4381 6910 -4347
rect 6968 -4381 7002 -4347
rect 7060 -4381 7094 -4347
rect 7152 -4381 7186 -4347
rect 7244 -4381 7278 -4347
rect 7336 -4381 7370 -4347
rect 7428 -4381 7462 -4347
rect 7520 -4381 7554 -4347
rect 7612 -4381 7646 -4347
rect 7704 -4381 7738 -4347
rect 7796 -4381 7830 -4347
rect 7888 -4381 7922 -4347
rect 7980 -4381 8014 -4347
rect 8072 -4381 8106 -4347
rect 8164 -4381 8198 -4347
rect 8256 -4381 8290 -4347
rect 8348 -4381 8382 -4347
rect 8440 -4381 8474 -4347
rect 8532 -4381 8566 -4347
rect 8624 -4381 8658 -4347
rect 8716 -4381 8750 -4347
rect 8808 -4381 8842 -4347
rect 8900 -4381 8934 -4347
rect 8992 -4381 9026 -4347
rect 9084 -4381 9118 -4347
rect 9176 -4381 9210 -4347
rect 9268 -4381 9302 -4347
rect 9360 -4381 9394 -4347
rect 9452 -4381 9486 -4347
rect 9544 -4381 9578 -4347
rect 9636 -4381 9670 -4347
rect 9728 -4381 9762 -4347
rect 9820 -4381 9854 -4347
rect 9912 -4381 9946 -4347
rect 10004 -4381 10038 -4347
rect 10096 -4381 10130 -4347
rect 10188 -4381 10222 -4347
rect 10280 -4381 10314 -4347
rect 10372 -4381 10406 -4347
rect 10464 -4381 10498 -4347
rect 10556 -4381 10590 -4347
rect 10648 -4381 10682 -4347
rect 10740 -4381 10774 -4347
rect 10832 -4381 10866 -4347
rect 10924 -4381 10958 -4347
rect 11016 -4381 11050 -4347
rect 11108 -4381 11142 -4347
rect 11200 -4381 11234 -4347
rect 11292 -4381 11326 -4347
rect 11384 -4381 11418 -4347
rect 11476 -4381 11510 -4347
rect 11568 -4381 11602 -4347
rect 11660 -4381 11694 -4347
rect 11752 -4381 11786 -4347
rect 11844 -4381 11878 -4347
rect 11936 -4381 11970 -4347
rect 12028 -4381 12062 -4347
rect 12120 -4381 12154 -4347
rect 12212 -4381 12246 -4347
rect 12304 -4381 12338 -4347
rect 12396 -4381 12430 -4347
rect 12488 -4381 12522 -4347
rect 12580 -4381 12614 -4347
rect 12672 -4381 12706 -4347
rect 12764 -4381 12798 -4347
rect 12856 -4381 12890 -4347
rect 12948 -4381 12982 -4347
rect 13040 -4381 13074 -4347
rect 13132 -4381 13166 -4347
rect 13224 -4381 13258 -4347
rect 13316 -4381 13350 -4347
rect 13408 -4381 13442 -4347
rect 13500 -4381 13534 -4347
rect 13592 -4381 13626 -4347
rect 13684 -4381 13718 -4347
rect 13776 -4381 13810 -4347
rect 13868 -4381 13902 -4347
rect 13960 -4381 13994 -4347
rect 14052 -4381 14086 -4347
rect 14144 -4381 14178 -4347
rect 14236 -4381 14270 -4347
rect 14328 -4381 14362 -4347
rect 14420 -4381 14454 -4347
rect 14512 -4381 14546 -4347
rect 14604 -4381 14638 -4347
rect 14696 -4381 14730 -4347
rect 14788 -4381 14822 -4347
rect 14880 -4381 14914 -4347
rect 14972 -4381 15006 -4347
rect 15064 -4381 15098 -4347
rect 15156 -4381 15190 -4347
rect 15248 -4381 15282 -4347
rect 15340 -4381 15374 -4347
rect 15432 -4381 15466 -4347
rect 15524 -4381 15558 -4347
rect 15616 -4381 15650 -4347
rect 15708 -4381 15742 -4347
rect 15800 -4381 15834 -4347
rect 15892 -4381 15926 -4347
rect 15984 -4381 16018 -4347
rect 16076 -4381 16110 -4347
rect 16168 -4381 16202 -4347
rect 16260 -4381 16294 -4347
rect 16352 -4381 16386 -4347
rect 16444 -4381 16478 -4347
rect 16536 -4381 16570 -4347
rect 16628 -4381 16662 -4347
rect -855 -4653 -821 -4619
rect -210 -4659 -176 -4656
rect -210 -4690 -202 -4659
rect -202 -4690 -176 -4659
rect 433 -4653 467 -4619
rect 1054 -4659 1088 -4652
rect 1054 -4686 1086 -4659
rect 1086 -4686 1088 -4659
rect 3014 -4686 3048 -4652
rect 3628 -4659 3662 -4652
rect 3628 -4686 3662 -4659
rect 5588 -4686 5622 -4652
rect 6202 -4659 6236 -4652
rect 6202 -4686 6204 -4659
rect 6204 -4686 6236 -4659
rect 8162 -4686 8196 -4652
rect 8776 -4659 8810 -4652
rect 8776 -4686 8780 -4659
rect 8780 -4686 8810 -4659
rect 10736 -4686 10770 -4652
rect 11384 -4659 11418 -4657
rect 11384 -4691 11390 -4659
rect 11390 -4691 11418 -4659
rect 15248 -4640 15282 -4606
rect 15341 -4640 15375 -4606
rect 13685 -4693 13692 -4686
rect 13692 -4693 13719 -4686
rect 13685 -4720 13719 -4693
rect 15248 -4736 15282 -4702
rect 15340 -4735 15374 -4701
rect -2968 -4925 -2934 -4891
rect -2876 -4925 -2842 -4891
rect -2784 -4925 -2750 -4891
rect -2692 -4925 -2658 -4891
rect -2600 -4925 -2566 -4891
rect -2508 -4925 -2474 -4891
rect -2416 -4925 -2382 -4891
rect -2324 -4925 -2290 -4891
rect -2232 -4925 -2198 -4891
rect -2140 -4925 -2106 -4891
rect -2048 -4925 -2014 -4891
rect -1956 -4925 -1922 -4891
rect -1864 -4925 -1830 -4891
rect -1772 -4925 -1738 -4891
rect -1680 -4925 -1646 -4891
rect -1588 -4925 -1554 -4891
rect -1496 -4925 -1462 -4891
rect -1404 -4925 -1370 -4891
rect -1312 -4925 -1278 -4891
rect -1220 -4925 -1186 -4891
rect -1128 -4925 -1094 -4891
rect -1036 -4925 -1002 -4891
rect -944 -4925 -910 -4891
rect -852 -4925 -818 -4891
rect -760 -4925 -726 -4891
rect -668 -4925 -634 -4891
rect -576 -4925 -542 -4891
rect -484 -4925 -450 -4891
rect -392 -4925 -358 -4891
rect -300 -4925 -266 -4891
rect -208 -4925 -174 -4891
rect -116 -4925 -82 -4891
rect -24 -4925 10 -4891
rect 68 -4925 102 -4891
rect 160 -4925 194 -4891
rect 252 -4925 286 -4891
rect 344 -4925 378 -4891
rect 436 -4925 470 -4891
rect 528 -4925 562 -4891
rect 620 -4925 654 -4891
rect 712 -4925 746 -4891
rect 804 -4925 838 -4891
rect 896 -4925 930 -4891
rect 988 -4925 1022 -4891
rect 1080 -4925 1114 -4891
rect 1172 -4925 1206 -4891
rect 1264 -4925 1298 -4891
rect 1356 -4925 1390 -4891
rect 1448 -4925 1482 -4891
rect 1540 -4925 1574 -4891
rect 1632 -4925 1666 -4891
rect 1724 -4925 1758 -4891
rect 1816 -4925 1850 -4891
rect 1908 -4925 1942 -4891
rect 2000 -4925 2034 -4891
rect 2092 -4925 2126 -4891
rect 2184 -4925 2218 -4891
rect 2276 -4925 2310 -4891
rect 2368 -4925 2402 -4891
rect 2460 -4925 2494 -4891
rect 2552 -4925 2586 -4891
rect 2644 -4925 2678 -4891
rect 2736 -4925 2770 -4891
rect 2828 -4925 2862 -4891
rect 2920 -4925 2954 -4891
rect 3012 -4925 3046 -4891
rect 3104 -4925 3138 -4891
rect 3196 -4925 3230 -4891
rect 3288 -4925 3322 -4891
rect 3380 -4925 3414 -4891
rect 3472 -4925 3506 -4891
rect 3564 -4925 3598 -4891
rect 3656 -4925 3690 -4891
rect 3748 -4925 3782 -4891
rect 3840 -4925 3874 -4891
rect 3932 -4925 3966 -4891
rect 4024 -4925 4058 -4891
rect 4116 -4925 4150 -4891
rect 4208 -4925 4242 -4891
rect 4300 -4925 4334 -4891
rect 4392 -4925 4426 -4891
rect 4484 -4925 4518 -4891
rect 4576 -4925 4610 -4891
rect 4668 -4925 4702 -4891
rect 4760 -4925 4794 -4891
rect 4852 -4925 4886 -4891
rect 4944 -4925 4978 -4891
rect 5036 -4925 5070 -4891
rect 5128 -4925 5162 -4891
rect 5220 -4925 5254 -4891
rect 5312 -4925 5346 -4891
rect 5404 -4925 5438 -4891
rect 5496 -4925 5530 -4891
rect 5588 -4925 5622 -4891
rect 5680 -4925 5714 -4891
rect 5772 -4925 5806 -4891
rect 5864 -4925 5898 -4891
rect 5956 -4925 5990 -4891
rect 6048 -4925 6082 -4891
rect 6140 -4925 6174 -4891
rect 6232 -4925 6266 -4891
rect 6324 -4925 6358 -4891
rect 6416 -4925 6450 -4891
rect 6508 -4925 6542 -4891
rect 6600 -4925 6634 -4891
rect 6692 -4925 6726 -4891
rect 6784 -4925 6818 -4891
rect 6876 -4925 6910 -4891
rect 6968 -4925 7002 -4891
rect 7060 -4925 7094 -4891
rect 7152 -4925 7186 -4891
rect 7244 -4925 7278 -4891
rect 7336 -4925 7370 -4891
rect 7428 -4925 7462 -4891
rect 7520 -4925 7554 -4891
rect 7612 -4925 7646 -4891
rect 7704 -4925 7738 -4891
rect 7796 -4925 7830 -4891
rect 7888 -4925 7922 -4891
rect 7980 -4925 8014 -4891
rect 8072 -4925 8106 -4891
rect 8164 -4925 8198 -4891
rect 8256 -4925 8290 -4891
rect 8348 -4925 8382 -4891
rect 8440 -4925 8474 -4891
rect 8532 -4925 8566 -4891
rect 8624 -4925 8658 -4891
rect 8716 -4925 8750 -4891
rect 8808 -4925 8842 -4891
rect 8900 -4925 8934 -4891
rect 8992 -4925 9026 -4891
rect 9084 -4925 9118 -4891
rect 9176 -4925 9210 -4891
rect 9268 -4925 9302 -4891
rect 9360 -4925 9394 -4891
rect 9452 -4925 9486 -4891
rect 9544 -4925 9578 -4891
rect 9636 -4925 9670 -4891
rect 9728 -4925 9762 -4891
rect 9820 -4925 9854 -4891
rect 9912 -4925 9946 -4891
rect 10004 -4925 10038 -4891
rect 10096 -4925 10130 -4891
rect 10188 -4925 10222 -4891
rect 10280 -4925 10314 -4891
rect 10372 -4925 10406 -4891
rect 10464 -4925 10498 -4891
rect 10556 -4925 10590 -4891
rect 10648 -4925 10682 -4891
rect 10740 -4925 10774 -4891
rect 10832 -4925 10866 -4891
rect 10924 -4925 10958 -4891
rect 11016 -4925 11050 -4891
rect 11108 -4925 11142 -4891
rect 11200 -4925 11234 -4891
rect 11292 -4925 11326 -4891
rect 11384 -4925 11418 -4891
rect 11476 -4925 11510 -4891
rect 11568 -4925 11602 -4891
rect 11660 -4925 11694 -4891
rect 11752 -4925 11786 -4891
rect 11844 -4925 11878 -4891
rect 11936 -4925 11970 -4891
rect 12028 -4925 12062 -4891
rect 12120 -4925 12154 -4891
rect 12212 -4925 12246 -4891
rect 12304 -4925 12338 -4891
rect 12396 -4925 12430 -4891
rect 12488 -4925 12522 -4891
rect 12580 -4925 12614 -4891
rect 12672 -4925 12706 -4891
rect 12764 -4925 12798 -4891
rect 12856 -4925 12890 -4891
rect 12948 -4925 12982 -4891
rect 13040 -4925 13074 -4891
rect 13132 -4925 13166 -4891
rect 13224 -4925 13258 -4891
rect 13316 -4925 13350 -4891
rect 13408 -4925 13442 -4891
rect 13500 -4925 13534 -4891
rect 13592 -4925 13626 -4891
rect 13684 -4925 13718 -4891
rect 13776 -4925 13810 -4891
rect 13868 -4925 13902 -4891
rect 13960 -4925 13994 -4891
rect 14052 -4925 14086 -4891
rect 14144 -4925 14178 -4891
rect 14236 -4925 14270 -4891
rect 14328 -4925 14362 -4891
rect 14420 -4925 14454 -4891
rect 14512 -4925 14546 -4891
rect 14604 -4925 14638 -4891
rect 14696 -4925 14730 -4891
rect 14788 -4925 14822 -4891
rect 14880 -4925 14914 -4891
rect 14972 -4925 15006 -4891
rect 15064 -4925 15098 -4891
rect 15156 -4925 15190 -4891
rect 15248 -4925 15282 -4891
rect 15340 -4925 15374 -4891
rect 15432 -4925 15466 -4891
rect 15524 -4925 15558 -4891
rect 15616 -4925 15650 -4891
rect 15708 -4925 15742 -4891
rect 15800 -4925 15834 -4891
rect 15892 -4925 15926 -4891
rect 15984 -4925 16018 -4891
rect 16076 -4925 16110 -4891
rect 16168 -4925 16202 -4891
rect 16260 -4925 16294 -4891
rect 16352 -4925 16386 -4891
rect 16444 -4925 16478 -4891
rect 16536 -4925 16570 -4891
rect 16628 -4925 16662 -4891
rect 436 -5157 464 -5128
rect 464 -5157 470 -5128
rect 436 -5162 470 -5157
rect 1082 -5163 1116 -5129
rect 3042 -5157 3074 -5129
rect 3074 -5157 3076 -5129
rect 3042 -5163 3076 -5157
rect 3656 -5163 3690 -5129
rect 5616 -5157 5650 -5129
rect 5616 -5163 5650 -5157
rect 6230 -5163 6264 -5129
rect 8190 -5157 8192 -5129
rect 8192 -5157 8224 -5129
rect 8190 -5163 8224 -5157
rect 8804 -5163 8838 -5129
rect 10764 -5157 10768 -5129
rect 10768 -5157 10798 -5129
rect 10764 -5163 10798 -5157
rect 11389 -5196 11423 -5162
rect 13038 -5095 13072 -5061
rect 12558 -5157 12574 -5126
rect 12574 -5157 12592 -5126
rect 12642 -5157 12676 -5126
rect 12739 -5157 12744 -5126
rect 12744 -5157 12773 -5126
rect 12836 -5157 12846 -5126
rect 12846 -5157 12870 -5126
rect 12942 -5157 12948 -5126
rect 12948 -5157 12976 -5126
rect 12558 -5160 12592 -5157
rect 12642 -5160 12676 -5157
rect 12739 -5160 12773 -5157
rect 12836 -5160 12870 -5157
rect 12942 -5160 12976 -5157
rect 13038 -5167 13072 -5133
rect 13684 -5123 13718 -5096
rect 13684 -5130 13692 -5123
rect 13692 -5130 13718 -5123
rect 15248 -5118 15282 -5084
rect 15341 -5118 15375 -5084
rect 15248 -5214 15282 -5180
rect 15340 -5213 15374 -5179
rect -2968 -5469 -2934 -5435
rect -2876 -5469 -2842 -5435
rect -2784 -5469 -2750 -5435
rect -2692 -5469 -2658 -5435
rect -2600 -5469 -2566 -5435
rect -2508 -5469 -2474 -5435
rect -2416 -5469 -2382 -5435
rect -2324 -5469 -2290 -5435
rect -2232 -5469 -2198 -5435
rect -2140 -5469 -2106 -5435
rect -2048 -5469 -2014 -5435
rect -1956 -5469 -1922 -5435
rect -1864 -5469 -1830 -5435
rect -1772 -5469 -1738 -5435
rect -1680 -5469 -1646 -5435
rect -1588 -5469 -1554 -5435
rect -1496 -5469 -1462 -5435
rect -1404 -5469 -1370 -5435
rect -1312 -5469 -1278 -5435
rect -1220 -5469 -1186 -5435
rect -1128 -5469 -1094 -5435
rect -1036 -5469 -1002 -5435
rect -944 -5469 -910 -5435
rect -852 -5469 -818 -5435
rect -760 -5469 -726 -5435
rect -668 -5469 -634 -5435
rect -576 -5469 -542 -5435
rect -484 -5469 -450 -5435
rect -392 -5469 -358 -5435
rect -300 -5469 -266 -5435
rect -208 -5469 -174 -5435
rect -116 -5469 -82 -5435
rect -24 -5469 10 -5435
rect 68 -5469 102 -5435
rect 160 -5469 194 -5435
rect 252 -5469 286 -5435
rect 344 -5469 378 -5435
rect 436 -5469 470 -5435
rect 528 -5469 562 -5435
rect 620 -5469 654 -5435
rect 712 -5469 746 -5435
rect 804 -5469 838 -5435
rect 896 -5469 930 -5435
rect 988 -5469 1022 -5435
rect 1080 -5469 1114 -5435
rect 1172 -5469 1206 -5435
rect 1264 -5469 1298 -5435
rect 1356 -5469 1390 -5435
rect 1448 -5469 1482 -5435
rect 1540 -5469 1574 -5435
rect 1632 -5469 1666 -5435
rect 1724 -5469 1758 -5435
rect 1816 -5469 1850 -5435
rect 1908 -5469 1942 -5435
rect 2000 -5469 2034 -5435
rect 2092 -5469 2126 -5435
rect 2184 -5469 2218 -5435
rect 2276 -5469 2310 -5435
rect 2368 -5469 2402 -5435
rect 2460 -5469 2494 -5435
rect 2552 -5469 2586 -5435
rect 2644 -5469 2678 -5435
rect 2736 -5469 2770 -5435
rect 2828 -5469 2862 -5435
rect 2920 -5469 2954 -5435
rect 3012 -5469 3046 -5435
rect 3104 -5469 3138 -5435
rect 3196 -5469 3230 -5435
rect 3288 -5469 3322 -5435
rect 3380 -5469 3414 -5435
rect 3472 -5469 3506 -5435
rect 3564 -5469 3598 -5435
rect 3656 -5469 3690 -5435
rect 3748 -5469 3782 -5435
rect 3840 -5469 3874 -5435
rect 3932 -5469 3966 -5435
rect 4024 -5469 4058 -5435
rect 4116 -5469 4150 -5435
rect 4208 -5469 4242 -5435
rect 4300 -5469 4334 -5435
rect 4392 -5469 4426 -5435
rect 4484 -5469 4518 -5435
rect 4576 -5469 4610 -5435
rect 4668 -5469 4702 -5435
rect 4760 -5469 4794 -5435
rect 4852 -5469 4886 -5435
rect 4944 -5469 4978 -5435
rect 5036 -5469 5070 -5435
rect 5128 -5469 5162 -5435
rect 5220 -5469 5254 -5435
rect 5312 -5469 5346 -5435
rect 5404 -5469 5438 -5435
rect 5496 -5469 5530 -5435
rect 5588 -5469 5622 -5435
rect 5680 -5469 5714 -5435
rect 5772 -5469 5806 -5435
rect 5864 -5469 5898 -5435
rect 5956 -5469 5990 -5435
rect 6048 -5469 6082 -5435
rect 6140 -5469 6174 -5435
rect 6232 -5469 6266 -5435
rect 6324 -5469 6358 -5435
rect 6416 -5469 6450 -5435
rect 6508 -5469 6542 -5435
rect 6600 -5469 6634 -5435
rect 6692 -5469 6726 -5435
rect 6784 -5469 6818 -5435
rect 6876 -5469 6910 -5435
rect 6968 -5469 7002 -5435
rect 7060 -5469 7094 -5435
rect 7152 -5469 7186 -5435
rect 7244 -5469 7278 -5435
rect 7336 -5469 7370 -5435
rect 7428 -5469 7462 -5435
rect 7520 -5469 7554 -5435
rect 7612 -5469 7646 -5435
rect 7704 -5469 7738 -5435
rect 7796 -5469 7830 -5435
rect 7888 -5469 7922 -5435
rect 7980 -5469 8014 -5435
rect 8072 -5469 8106 -5435
rect 8164 -5469 8198 -5435
rect 8256 -5469 8290 -5435
rect 8348 -5469 8382 -5435
rect 8440 -5469 8474 -5435
rect 8532 -5469 8566 -5435
rect 8624 -5469 8658 -5435
rect 8716 -5469 8750 -5435
rect 8808 -5469 8842 -5435
rect 8900 -5469 8934 -5435
rect 8992 -5469 9026 -5435
rect 9084 -5469 9118 -5435
rect 9176 -5469 9210 -5435
rect 9268 -5469 9302 -5435
rect 9360 -5469 9394 -5435
rect 9452 -5469 9486 -5435
rect 9544 -5469 9578 -5435
rect 9636 -5469 9670 -5435
rect 9728 -5469 9762 -5435
rect 9820 -5469 9854 -5435
rect 9912 -5469 9946 -5435
rect 10004 -5469 10038 -5435
rect 10096 -5469 10130 -5435
rect 10188 -5469 10222 -5435
rect 10280 -5469 10314 -5435
rect 10372 -5469 10406 -5435
rect 10464 -5469 10498 -5435
rect 10556 -5469 10590 -5435
rect 10648 -5469 10682 -5435
rect 10740 -5469 10774 -5435
rect 10832 -5469 10866 -5435
rect 10924 -5469 10958 -5435
rect 11016 -5469 11050 -5435
rect 11108 -5469 11142 -5435
rect 11200 -5469 11234 -5435
rect 11292 -5469 11326 -5435
rect 11384 -5469 11418 -5435
rect 11476 -5469 11510 -5435
rect 11568 -5469 11602 -5435
rect 11660 -5469 11694 -5435
rect 11752 -5469 11786 -5435
rect 11844 -5469 11878 -5435
rect 11936 -5469 11970 -5435
rect 12028 -5469 12062 -5435
rect 12120 -5469 12154 -5435
rect 12212 -5469 12246 -5435
rect 12304 -5469 12338 -5435
rect 12396 -5469 12430 -5435
rect 12488 -5469 12522 -5435
rect 12580 -5469 12614 -5435
rect 12672 -5469 12706 -5435
rect 12764 -5469 12798 -5435
rect 12856 -5469 12890 -5435
rect 12948 -5469 12982 -5435
rect 13040 -5469 13074 -5435
rect 13132 -5469 13166 -5435
rect 13224 -5469 13258 -5435
rect 13316 -5469 13350 -5435
rect 13408 -5469 13442 -5435
rect 13500 -5469 13534 -5435
rect 13592 -5469 13626 -5435
rect 13684 -5469 13718 -5435
rect 13776 -5469 13810 -5435
rect 13868 -5469 13902 -5435
rect 13960 -5469 13994 -5435
rect 14052 -5469 14086 -5435
rect 14144 -5469 14178 -5435
rect 14236 -5469 14270 -5435
rect 14328 -5469 14362 -5435
rect 14420 -5469 14454 -5435
rect 14512 -5469 14546 -5435
rect 14604 -5469 14638 -5435
rect 14696 -5469 14730 -5435
rect 14788 -5469 14822 -5435
rect 14880 -5469 14914 -5435
rect 14972 -5469 15006 -5435
rect 15064 -5469 15098 -5435
rect 15156 -5469 15190 -5435
rect 15248 -5469 15282 -5435
rect 15340 -5469 15374 -5435
rect 15432 -5469 15466 -5435
rect 15524 -5469 15558 -5435
rect 15616 -5469 15650 -5435
rect 15708 -5469 15742 -5435
rect 15800 -5469 15834 -5435
rect 15892 -5469 15926 -5435
rect 15984 -5469 16018 -5435
rect 16076 -5469 16110 -5435
rect 16168 -5469 16202 -5435
rect 16260 -5469 16294 -5435
rect 16352 -5469 16386 -5435
rect 16444 -5469 16478 -5435
rect 16536 -5469 16570 -5435
rect 16628 -5469 16662 -5435
rect 432 -5742 466 -5708
rect 1052 -5747 1086 -5743
rect 1052 -5777 1086 -5747
rect 3012 -5777 3046 -5743
rect 3626 -5747 3660 -5743
rect 3626 -5777 3628 -5747
rect 3628 -5777 3660 -5747
rect 5586 -5777 5620 -5743
rect 6200 -5747 6234 -5743
rect 6200 -5777 6204 -5747
rect 6204 -5777 6234 -5747
rect 8160 -5777 8194 -5743
rect 8774 -5747 8808 -5743
rect 8774 -5777 8780 -5747
rect 8780 -5777 8808 -5747
rect 10737 -5775 10771 -5741
rect 11369 -5747 11403 -5740
rect 11369 -5774 11390 -5747
rect 11390 -5774 11403 -5747
rect 15248 -5728 15282 -5694
rect 15341 -5728 15375 -5694
rect 13685 -5781 13692 -5772
rect 13692 -5781 13719 -5772
rect 13685 -5806 13719 -5781
rect 15248 -5824 15282 -5790
rect 15340 -5823 15374 -5789
rect -2968 -6013 -2934 -5979
rect -2876 -6013 -2842 -5979
rect -2784 -6013 -2750 -5979
rect -2692 -6013 -2658 -5979
rect -2600 -6013 -2566 -5979
rect -2508 -6013 -2474 -5979
rect -2416 -6013 -2382 -5979
rect -2324 -6013 -2290 -5979
rect -2232 -6013 -2198 -5979
rect -2140 -6013 -2106 -5979
rect -2048 -6013 -2014 -5979
rect -1956 -6013 -1922 -5979
rect -1864 -6013 -1830 -5979
rect -1772 -6013 -1738 -5979
rect -1680 -6013 -1646 -5979
rect -1588 -6013 -1554 -5979
rect -1496 -6013 -1462 -5979
rect -1404 -6013 -1370 -5979
rect -1312 -6013 -1278 -5979
rect -1220 -6013 -1186 -5979
rect -1128 -6013 -1094 -5979
rect -1036 -6013 -1002 -5979
rect -944 -6013 -910 -5979
rect -852 -6013 -818 -5979
rect -760 -6013 -726 -5979
rect -668 -6013 -634 -5979
rect -576 -6013 -542 -5979
rect -484 -6013 -450 -5979
rect -392 -6013 -358 -5979
rect -300 -6013 -266 -5979
rect -208 -6013 -174 -5979
rect -116 -6013 -82 -5979
rect -24 -6013 10 -5979
rect 68 -6013 102 -5979
rect 160 -6013 194 -5979
rect 252 -6013 286 -5979
rect 344 -6013 378 -5979
rect 436 -6013 470 -5979
rect 528 -6013 562 -5979
rect 620 -6013 654 -5979
rect 712 -6013 746 -5979
rect 804 -6013 838 -5979
rect 896 -6013 930 -5979
rect 988 -6013 1022 -5979
rect 1080 -6013 1114 -5979
rect 1172 -6013 1206 -5979
rect 1264 -6013 1298 -5979
rect 1356 -6013 1390 -5979
rect 1448 -6013 1482 -5979
rect 1540 -6013 1574 -5979
rect 1632 -6013 1666 -5979
rect 1724 -6013 1758 -5979
rect 1816 -6013 1850 -5979
rect 1908 -6013 1942 -5979
rect 2000 -6013 2034 -5979
rect 2092 -6013 2126 -5979
rect 2184 -6013 2218 -5979
rect 2276 -6013 2310 -5979
rect 2368 -6013 2402 -5979
rect 2460 -6013 2494 -5979
rect 2552 -6013 2586 -5979
rect 2644 -6013 2678 -5979
rect 2736 -6013 2770 -5979
rect 2828 -6013 2862 -5979
rect 2920 -6013 2954 -5979
rect 3012 -6013 3046 -5979
rect 3104 -6013 3138 -5979
rect 3196 -6013 3230 -5979
rect 3288 -6013 3322 -5979
rect 3380 -6013 3414 -5979
rect 3472 -6013 3506 -5979
rect 3564 -6013 3598 -5979
rect 3656 -6013 3690 -5979
rect 3748 -6013 3782 -5979
rect 3840 -6013 3874 -5979
rect 3932 -6013 3966 -5979
rect 4024 -6013 4058 -5979
rect 4116 -6013 4150 -5979
rect 4208 -6013 4242 -5979
rect 4300 -6013 4334 -5979
rect 4392 -6013 4426 -5979
rect 4484 -6013 4518 -5979
rect 4576 -6013 4610 -5979
rect 4668 -6013 4702 -5979
rect 4760 -6013 4794 -5979
rect 4852 -6013 4886 -5979
rect 4944 -6013 4978 -5979
rect 5036 -6013 5070 -5979
rect 5128 -6013 5162 -5979
rect 5220 -6013 5254 -5979
rect 5312 -6013 5346 -5979
rect 5404 -6013 5438 -5979
rect 5496 -6013 5530 -5979
rect 5588 -6013 5622 -5979
rect 5680 -6013 5714 -5979
rect 5772 -6013 5806 -5979
rect 5864 -6013 5898 -5979
rect 5956 -6013 5990 -5979
rect 6048 -6013 6082 -5979
rect 6140 -6013 6174 -5979
rect 6232 -6013 6266 -5979
rect 6324 -6013 6358 -5979
rect 6416 -6013 6450 -5979
rect 6508 -6013 6542 -5979
rect 6600 -6013 6634 -5979
rect 6692 -6013 6726 -5979
rect 6784 -6013 6818 -5979
rect 6876 -6013 6910 -5979
rect 6968 -6013 7002 -5979
rect 7060 -6013 7094 -5979
rect 7152 -6013 7186 -5979
rect 7244 -6013 7278 -5979
rect 7336 -6013 7370 -5979
rect 7428 -6013 7462 -5979
rect 7520 -6013 7554 -5979
rect 7612 -6013 7646 -5979
rect 7704 -6013 7738 -5979
rect 7796 -6013 7830 -5979
rect 7888 -6013 7922 -5979
rect 7980 -6013 8014 -5979
rect 8072 -6013 8106 -5979
rect 8164 -6013 8198 -5979
rect 8256 -6013 8290 -5979
rect 8348 -6013 8382 -5979
rect 8440 -6013 8474 -5979
rect 8532 -6013 8566 -5979
rect 8624 -6013 8658 -5979
rect 8716 -6013 8750 -5979
rect 8808 -6013 8842 -5979
rect 8900 -6013 8934 -5979
rect 8992 -6013 9026 -5979
rect 9084 -6013 9118 -5979
rect 9176 -6013 9210 -5979
rect 9268 -6013 9302 -5979
rect 9360 -6013 9394 -5979
rect 9452 -6013 9486 -5979
rect 9544 -6013 9578 -5979
rect 9636 -6013 9670 -5979
rect 9728 -6013 9762 -5979
rect 9820 -6013 9854 -5979
rect 9912 -6013 9946 -5979
rect 10004 -6013 10038 -5979
rect 10096 -6013 10130 -5979
rect 10188 -6013 10222 -5979
rect 10280 -6013 10314 -5979
rect 10372 -6013 10406 -5979
rect 10464 -6013 10498 -5979
rect 10556 -6013 10590 -5979
rect 10648 -6013 10682 -5979
rect 10740 -6013 10774 -5979
rect 10832 -6013 10866 -5979
rect 10924 -6013 10958 -5979
rect 11016 -6013 11050 -5979
rect 11108 -6013 11142 -5979
rect 11200 -6013 11234 -5979
rect 11292 -6013 11326 -5979
rect 11384 -6013 11418 -5979
rect 11476 -6013 11510 -5979
rect 11568 -6013 11602 -5979
rect 11660 -6013 11694 -5979
rect 11752 -6013 11786 -5979
rect 11844 -6013 11878 -5979
rect 11936 -6013 11970 -5979
rect 12028 -6013 12062 -5979
rect 12120 -6013 12154 -5979
rect 12212 -6013 12246 -5979
rect 12304 -6013 12338 -5979
rect 12396 -6013 12430 -5979
rect 12488 -6013 12522 -5979
rect 12580 -6013 12614 -5979
rect 12672 -6013 12706 -5979
rect 12764 -6013 12798 -5979
rect 12856 -6013 12890 -5979
rect 12948 -6013 12982 -5979
rect 13040 -6013 13074 -5979
rect 13132 -6013 13166 -5979
rect 13224 -6013 13258 -5979
rect 13316 -6013 13350 -5979
rect 13408 -6013 13442 -5979
rect 13500 -6013 13534 -5979
rect 13592 -6013 13626 -5979
rect 13684 -6013 13718 -5979
rect 13776 -6013 13810 -5979
rect 13868 -6013 13902 -5979
rect 13960 -6013 13994 -5979
rect 14052 -6013 14086 -5979
rect 14144 -6013 14178 -5979
rect 14236 -6013 14270 -5979
rect 14328 -6013 14362 -5979
rect 14420 -6013 14454 -5979
rect 14512 -6013 14546 -5979
rect 14604 -6013 14638 -5979
rect 14696 -6013 14730 -5979
rect 14788 -6013 14822 -5979
rect 14880 -6013 14914 -5979
rect 14972 -6013 15006 -5979
rect 15064 -6013 15098 -5979
rect 15156 -6013 15190 -5979
rect 15248 -6013 15282 -5979
rect 15340 -6013 15374 -5979
rect 15432 -6013 15466 -5979
rect 15524 -6013 15558 -5979
rect 15616 -6013 15650 -5979
rect 15708 -6013 15742 -5979
rect 15800 -6013 15834 -5979
rect 15892 -6013 15926 -5979
rect 15984 -6013 16018 -5979
rect 16076 -6013 16110 -5979
rect 16168 -6013 16202 -5979
rect 16260 -6013 16294 -5979
rect 16352 -6013 16386 -5979
rect 16444 -6013 16478 -5979
rect 16536 -6013 16570 -5979
rect 16628 -6013 16662 -5979
rect -848 -6140 -814 -6106
rect -769 -6123 -735 -6106
rect -769 -6140 -766 -6123
rect -766 -6140 -735 -6123
rect -932 -6245 -903 -6218
rect -903 -6245 -898 -6218
rect -932 -6252 -898 -6245
rect -760 -6245 -735 -6217
rect -735 -6245 -726 -6217
rect -760 -6251 -726 -6245
rect 434 -6207 468 -6173
rect -30 -6245 4 -6211
rect 106 -6245 140 -6211
rect 242 -6245 276 -6211
rect 1076 -6167 1110 -6133
rect 1076 -6211 1110 -6206
rect 1076 -6240 1082 -6211
rect 1082 -6240 1110 -6211
rect 1171 -6246 1205 -6212
rect 1263 -6246 1297 -6212
rect 2369 -6245 2396 -6217
rect 2396 -6245 2403 -6217
rect 2369 -6251 2403 -6245
rect 3015 -6250 3049 -6216
rect 6876 -6245 6904 -6216
rect 6904 -6245 6910 -6216
rect 6876 -6250 6910 -6245
rect 7522 -6250 7556 -6216
rect 8164 -6245 8192 -6215
rect 8192 -6245 8198 -6215
rect 8164 -6249 8198 -6245
rect 8811 -6251 8845 -6217
rect 9453 -6245 9480 -6217
rect 9480 -6245 9487 -6217
rect 9453 -6251 9487 -6245
rect 10099 -6252 10133 -6218
rect 10741 -6245 10749 -6217
rect 10749 -6245 10775 -6217
rect 10832 -6245 10864 -6217
rect 10864 -6245 10866 -6217
rect 10925 -6245 10948 -6216
rect 10948 -6245 10959 -6216
rect 11017 -6245 11032 -6216
rect 11032 -6245 11051 -6216
rect 10741 -6251 10775 -6245
rect 10832 -6251 10866 -6245
rect 10925 -6250 10959 -6245
rect 11017 -6250 11051 -6245
rect 11129 -6284 11163 -6250
rect 11250 -6245 11284 -6219
rect 11344 -6245 11368 -6219
rect 11368 -6245 11378 -6219
rect 11250 -6253 11284 -6245
rect 11344 -6253 11378 -6245
rect -2968 -6557 -2934 -6523
rect -2876 -6557 -2842 -6523
rect -2784 -6557 -2750 -6523
rect -2692 -6557 -2658 -6523
rect -2600 -6557 -2566 -6523
rect -2508 -6557 -2474 -6523
rect -2416 -6557 -2382 -6523
rect -2324 -6557 -2290 -6523
rect -2232 -6557 -2198 -6523
rect -2140 -6557 -2106 -6523
rect -2048 -6557 -2014 -6523
rect -1956 -6557 -1922 -6523
rect -1864 -6557 -1830 -6523
rect -1772 -6557 -1738 -6523
rect -1680 -6557 -1646 -6523
rect -1588 -6557 -1554 -6523
rect -1496 -6557 -1462 -6523
rect -1404 -6557 -1370 -6523
rect -1312 -6557 -1278 -6523
rect -1220 -6557 -1186 -6523
rect -1128 -6557 -1094 -6523
rect -1036 -6557 -1002 -6523
rect -944 -6557 -910 -6523
rect -852 -6557 -818 -6523
rect -760 -6557 -726 -6523
rect -668 -6557 -634 -6523
rect -576 -6557 -542 -6523
rect -484 -6557 -450 -6523
rect -392 -6557 -358 -6523
rect -300 -6557 -266 -6523
rect -208 -6557 -174 -6523
rect -116 -6557 -82 -6523
rect -24 -6557 10 -6523
rect 68 -6557 102 -6523
rect 160 -6557 194 -6523
rect 252 -6557 286 -6523
rect 344 -6557 378 -6523
rect 436 -6557 470 -6523
rect 528 -6557 562 -6523
rect 620 -6557 654 -6523
rect 712 -6557 746 -6523
rect 804 -6557 838 -6523
rect 896 -6557 930 -6523
rect 988 -6557 1022 -6523
rect 1080 -6557 1114 -6523
rect 1172 -6557 1206 -6523
rect 1264 -6557 1298 -6523
rect 1356 -6557 1390 -6523
rect 1448 -6557 1482 -6523
rect 1540 -6557 1574 -6523
rect 1632 -6557 1666 -6523
rect 1724 -6557 1758 -6523
rect 1816 -6557 1850 -6523
rect 1908 -6557 1942 -6523
rect 2000 -6557 2034 -6523
rect 2092 -6557 2126 -6523
rect 2184 -6557 2218 -6523
rect 2276 -6557 2310 -6523
rect 2368 -6557 2402 -6523
rect 2460 -6557 2494 -6523
rect 2552 -6557 2586 -6523
rect 2644 -6557 2678 -6523
rect 2736 -6557 2770 -6523
rect 2828 -6557 2862 -6523
rect 2920 -6557 2954 -6523
rect 3012 -6557 3046 -6523
rect 3104 -6557 3138 -6523
rect 3196 -6557 3230 -6523
rect 3288 -6557 3322 -6523
rect 3380 -6557 3414 -6523
rect 3472 -6557 3506 -6523
rect 3564 -6557 3598 -6523
rect 3656 -6557 3690 -6523
rect 3748 -6557 3782 -6523
rect 3840 -6557 3874 -6523
rect 3932 -6557 3966 -6523
rect 4024 -6557 4058 -6523
rect 4116 -6557 4150 -6523
rect 4208 -6557 4242 -6523
rect 4300 -6557 4334 -6523
rect 4392 -6557 4426 -6523
rect 4484 -6557 4518 -6523
rect 4576 -6557 4610 -6523
rect 4668 -6557 4702 -6523
rect 4760 -6557 4794 -6523
rect 4852 -6557 4886 -6523
rect 4944 -6557 4978 -6523
rect 5036 -6557 5070 -6523
rect 5128 -6557 5162 -6523
rect 5220 -6557 5254 -6523
rect 5312 -6557 5346 -6523
rect 5404 -6557 5438 -6523
rect 5496 -6557 5530 -6523
rect 5588 -6557 5622 -6523
rect 5680 -6557 5714 -6523
rect 5772 -6557 5806 -6523
rect 5864 -6557 5898 -6523
rect 5956 -6557 5990 -6523
rect 6048 -6557 6082 -6523
rect 6140 -6557 6174 -6523
rect 6232 -6557 6266 -6523
rect 6324 -6557 6358 -6523
rect 6416 -6557 6450 -6523
rect 6508 -6557 6542 -6523
rect 6600 -6557 6634 -6523
rect 6692 -6557 6726 -6523
rect 6784 -6557 6818 -6523
rect 6876 -6557 6910 -6523
rect 6968 -6557 7002 -6523
rect 7060 -6557 7094 -6523
rect 7152 -6557 7186 -6523
rect 7244 -6557 7278 -6523
rect 7336 -6557 7370 -6523
rect 7428 -6557 7462 -6523
rect 7520 -6557 7554 -6523
rect 7612 -6557 7646 -6523
rect 7704 -6557 7738 -6523
rect 7796 -6557 7830 -6523
rect 7888 -6557 7922 -6523
rect 7980 -6557 8014 -6523
rect 8072 -6557 8106 -6523
rect 8164 -6557 8198 -6523
rect 8256 -6557 8290 -6523
rect 8348 -6557 8382 -6523
rect 8440 -6557 8474 -6523
rect 8532 -6557 8566 -6523
rect 8624 -6557 8658 -6523
rect 8716 -6557 8750 -6523
rect 8808 -6557 8842 -6523
rect 8900 -6557 8934 -6523
rect 8992 -6557 9026 -6523
rect 9084 -6557 9118 -6523
rect 9176 -6557 9210 -6523
rect 9268 -6557 9302 -6523
rect 9360 -6557 9394 -6523
rect 9452 -6557 9486 -6523
rect 9544 -6557 9578 -6523
rect 9636 -6557 9670 -6523
rect 9728 -6557 9762 -6523
rect 9820 -6557 9854 -6523
rect 9912 -6557 9946 -6523
rect 10004 -6557 10038 -6523
rect 10096 -6557 10130 -6523
rect 10188 -6557 10222 -6523
rect 10280 -6557 10314 -6523
rect 10372 -6557 10406 -6523
rect 10464 -6557 10498 -6523
rect 10556 -6557 10590 -6523
rect 10648 -6557 10682 -6523
rect 10740 -6557 10774 -6523
rect 10832 -6557 10866 -6523
rect 10924 -6557 10958 -6523
rect 11016 -6557 11050 -6523
rect 11108 -6557 11142 -6523
rect 11200 -6557 11234 -6523
rect 11292 -6557 11326 -6523
rect 11384 -6557 11418 -6523
rect 11476 -6557 11510 -6523
rect 11568 -6557 11602 -6523
rect 11660 -6557 11694 -6523
rect 11752 -6557 11786 -6523
rect 11844 -6557 11878 -6523
rect 11936 -6557 11970 -6523
rect 12028 -6557 12062 -6523
rect 12120 -6557 12154 -6523
rect 12212 -6557 12246 -6523
rect 12304 -6557 12338 -6523
rect 12396 -6557 12430 -6523
rect 12488 -6557 12522 -6523
rect 12580 -6557 12614 -6523
rect 12672 -6557 12706 -6523
rect 12764 -6557 12798 -6523
rect 12856 -6557 12890 -6523
rect 12948 -6557 12982 -6523
rect 13040 -6557 13074 -6523
rect 13132 -6557 13166 -6523
rect 13224 -6557 13258 -6523
rect 13316 -6557 13350 -6523
rect 13408 -6557 13442 -6523
rect 13500 -6557 13534 -6523
rect 13592 -6557 13626 -6523
rect 13684 -6557 13718 -6523
rect 13776 -6557 13810 -6523
rect 13868 -6557 13902 -6523
rect 13960 -6557 13994 -6523
rect 14052 -6557 14086 -6523
rect 14144 -6557 14178 -6523
rect 14236 -6557 14270 -6523
rect 14328 -6557 14362 -6523
rect 14420 -6557 14454 -6523
rect 14512 -6557 14546 -6523
rect 14604 -6557 14638 -6523
rect 14696 -6557 14730 -6523
rect 14788 -6557 14822 -6523
rect 14880 -6557 14914 -6523
rect 14972 -6557 15006 -6523
rect 15064 -6557 15098 -6523
rect 15156 -6557 15190 -6523
rect 15248 -6557 15282 -6523
rect 15340 -6557 15374 -6523
rect 15432 -6557 15466 -6523
rect 15524 -6557 15558 -6523
rect 15616 -6557 15650 -6523
rect 15708 -6557 15742 -6523
rect 15800 -6557 15834 -6523
rect 15892 -6557 15926 -6523
rect 15984 -6557 16018 -6523
rect 16076 -6557 16110 -6523
rect 16168 -6557 16202 -6523
rect 16260 -6557 16294 -6523
rect 16352 -6557 16386 -6523
rect 16444 -6557 16478 -6523
rect 16536 -6557 16570 -6523
rect 16628 -6557 16662 -6523
rect -2503 -6727 -2469 -6693
rect -2599 -6835 -2565 -6830
rect -2599 -6864 -2597 -6835
rect -2597 -6864 -2565 -6835
rect -2424 -6795 -2390 -6761
rect -2343 -6916 -2309 -6882
rect -2083 -6719 -2049 -6693
rect -2083 -6727 -2081 -6719
rect -2081 -6727 -2049 -6719
rect -2186 -6795 -2152 -6761
rect -1769 -6727 -1735 -6693
rect -1682 -6795 -1648 -6761
rect -1233 -6988 -1199 -6960
rect -1233 -6994 -1199 -6988
rect -940 -6914 -906 -6880
rect -2968 -7101 -2934 -7067
rect -2876 -7101 -2842 -7067
rect -2784 -7101 -2750 -7067
rect -2692 -7101 -2658 -7067
rect -2600 -7101 -2566 -7067
rect -2508 -7101 -2474 -7067
rect -2416 -7101 -2382 -7067
rect -2324 -7101 -2290 -7067
rect -2232 -7101 -2198 -7067
rect -2140 -7101 -2106 -7067
rect -2048 -7101 -2014 -7067
rect -1956 -7101 -1922 -7067
rect -1864 -7101 -1830 -7067
rect -1772 -7101 -1738 -7067
rect -1680 -7101 -1646 -7067
rect -1588 -7101 -1554 -7067
rect -1496 -7101 -1462 -7067
rect -1404 -7101 -1370 -7067
rect -1312 -7101 -1278 -7067
rect -1220 -7101 -1186 -7067
rect -1128 -7101 -1094 -7067
rect -1036 -7101 -1002 -7067
rect -944 -7101 -910 -7067
rect -852 -7101 -818 -7067
rect -760 -7101 -726 -7067
rect -668 -7101 -634 -7067
rect -576 -7101 -542 -7067
rect -484 -7101 -450 -7067
rect -392 -7101 -358 -7067
rect -300 -7101 -266 -7067
rect -208 -7101 -174 -7067
rect -116 -7101 -82 -7067
rect -24 -7101 10 -7067
rect 68 -7101 102 -7067
rect 160 -7101 194 -7067
rect 252 -7101 286 -7067
rect 344 -7101 378 -7067
rect 436 -7101 470 -7067
rect 528 -7101 562 -7067
rect 620 -7101 654 -7067
rect 712 -7101 746 -7067
rect 804 -7101 838 -7067
rect 896 -7101 930 -7067
rect 988 -7101 1022 -7067
rect 1080 -7101 1114 -7067
rect 1172 -7101 1206 -7067
rect 1264 -7101 1298 -7067
rect 1356 -7101 1390 -7067
rect 1448 -7101 1482 -7067
rect 1540 -7101 1574 -7067
rect 1632 -7101 1666 -7067
rect 1724 -7101 1758 -7067
rect 1816 -7101 1850 -7067
rect 1908 -7101 1942 -7067
rect 2000 -7101 2034 -7067
rect 2092 -7101 2126 -7067
rect 2184 -7101 2218 -7067
rect 2276 -7101 2310 -7067
rect 2368 -7101 2402 -7067
rect 2460 -7101 2494 -7067
rect 2552 -7101 2586 -7067
rect 2644 -7101 2678 -7067
rect 2736 -7101 2770 -7067
rect 2828 -7101 2862 -7067
rect 2920 -7101 2954 -7067
rect 3012 -7101 3046 -7067
rect 3104 -7101 3138 -7067
rect 3196 -7101 3230 -7067
rect 3288 -7101 3322 -7067
rect 3380 -7101 3414 -7067
rect 3472 -7101 3506 -7067
rect 3564 -7101 3598 -7067
rect 3656 -7101 3690 -7067
rect 3748 -7101 3782 -7067
rect 3840 -7101 3874 -7067
rect 3932 -7101 3966 -7067
rect 4024 -7101 4058 -7067
rect 4116 -7101 4150 -7067
rect 4208 -7101 4242 -7067
rect 4300 -7101 4334 -7067
rect 4392 -7101 4426 -7067
rect 4484 -7101 4518 -7067
rect 4576 -7101 4610 -7067
rect 4668 -7101 4702 -7067
rect 4760 -7101 4794 -7067
rect 4852 -7101 4886 -7067
rect 4944 -7101 4978 -7067
rect 5036 -7101 5070 -7067
rect 5128 -7101 5162 -7067
rect 5220 -7101 5254 -7067
rect 5312 -7101 5346 -7067
rect 5404 -7101 5438 -7067
rect 5496 -7101 5530 -7067
rect 5588 -7101 5622 -7067
rect 5680 -7101 5714 -7067
rect 5772 -7101 5806 -7067
rect 5864 -7101 5898 -7067
rect 5956 -7101 5990 -7067
rect 6048 -7101 6082 -7067
rect 6140 -7101 6174 -7067
rect 6232 -7101 6266 -7067
rect 6324 -7101 6358 -7067
rect 6416 -7101 6450 -7067
rect 6508 -7101 6542 -7067
rect 6600 -7101 6634 -7067
rect 6692 -7101 6726 -7067
rect 6784 -7101 6818 -7067
rect 6876 -7101 6910 -7067
rect 6968 -7101 7002 -7067
rect 7060 -7101 7094 -7067
rect 7152 -7101 7186 -7067
rect 7244 -7101 7278 -7067
rect 7336 -7101 7370 -7067
rect 7428 -7101 7462 -7067
rect 7520 -7101 7554 -7067
rect 7612 -7101 7646 -7067
rect 7704 -7101 7738 -7067
rect 7796 -7101 7830 -7067
rect 7888 -7101 7922 -7067
rect 7980 -7101 8014 -7067
rect 8072 -7101 8106 -7067
rect 8164 -7101 8198 -7067
rect 8256 -7101 8290 -7067
rect 8348 -7101 8382 -7067
rect 8440 -7101 8474 -7067
rect 8532 -7101 8566 -7067
rect 8624 -7101 8658 -7067
rect 8716 -7101 8750 -7067
rect 8808 -7101 8842 -7067
rect 8900 -7101 8934 -7067
rect 8992 -7101 9026 -7067
rect 9084 -7101 9118 -7067
rect 9176 -7101 9210 -7067
rect 9268 -7101 9302 -7067
rect 9360 -7101 9394 -7067
rect 9452 -7101 9486 -7067
rect 9544 -7101 9578 -7067
rect 9636 -7101 9670 -7067
rect 9728 -7101 9762 -7067
rect 9820 -7101 9854 -7067
rect 9912 -7101 9946 -7067
rect 10004 -7101 10038 -7067
rect 10096 -7101 10130 -7067
rect 10188 -7101 10222 -7067
rect 10280 -7101 10314 -7067
rect 10372 -7101 10406 -7067
rect 10464 -7101 10498 -7067
rect 10556 -7101 10590 -7067
rect 10648 -7101 10682 -7067
rect 10740 -7101 10774 -7067
rect 10832 -7101 10866 -7067
rect 10924 -7101 10958 -7067
rect 11016 -7101 11050 -7067
rect 11108 -7101 11142 -7067
rect 11200 -7101 11234 -7067
rect 11292 -7101 11326 -7067
rect 11384 -7101 11418 -7067
rect 11476 -7101 11510 -7067
rect 11568 -7101 11602 -7067
rect 11660 -7101 11694 -7067
rect 11752 -7101 11786 -7067
rect 11844 -7101 11878 -7067
rect 11936 -7101 11970 -7067
rect 12028 -7101 12062 -7067
rect 12120 -7101 12154 -7067
rect 12212 -7101 12246 -7067
rect 12304 -7101 12338 -7067
rect 12396 -7101 12430 -7067
rect 12488 -7101 12522 -7067
rect 12580 -7101 12614 -7067
rect 12672 -7101 12706 -7067
rect 12764 -7101 12798 -7067
rect 12856 -7101 12890 -7067
rect 12948 -7101 12982 -7067
rect 13040 -7101 13074 -7067
rect 13132 -7101 13166 -7067
rect 13224 -7101 13258 -7067
rect 13316 -7101 13350 -7067
rect 13408 -7101 13442 -7067
rect 13500 -7101 13534 -7067
rect 13592 -7101 13626 -7067
rect 13684 -7101 13718 -7067
rect 13776 -7101 13810 -7067
rect 13868 -7101 13902 -7067
rect 13960 -7101 13994 -7067
rect 14052 -7101 14086 -7067
rect 14144 -7101 14178 -7067
rect 14236 -7101 14270 -7067
rect 14328 -7101 14362 -7067
rect 14420 -7101 14454 -7067
rect 14512 -7101 14546 -7067
rect 14604 -7101 14638 -7067
rect 14696 -7101 14730 -7067
rect 14788 -7101 14822 -7067
rect 14880 -7101 14914 -7067
rect 14972 -7101 15006 -7067
rect 15064 -7101 15098 -7067
rect 15156 -7101 15190 -7067
rect 15248 -7101 15282 -7067
rect 15340 -7101 15374 -7067
rect 15432 -7101 15466 -7067
rect 15524 -7101 15558 -7067
rect 15616 -7101 15650 -7067
rect 15708 -7101 15742 -7067
rect 15800 -7101 15834 -7067
rect 15892 -7101 15926 -7067
rect 15984 -7101 16018 -7067
rect 16076 -7101 16110 -7067
rect 16168 -7101 16202 -7067
rect 16260 -7101 16294 -7067
rect 16352 -7101 16386 -7067
rect 16444 -7101 16478 -7067
rect 16536 -7101 16570 -7067
rect 16628 -7101 16662 -7067
rect 2934 -7304 2968 -7270
rect 3111 -7225 3145 -7191
rect 3852 -7222 3886 -7188
rect 3747 -7333 3755 -7304
rect 3755 -7333 3781 -7304
rect 3747 -7338 3781 -7333
rect 3928 -7333 3957 -7305
rect 3957 -7333 3962 -7305
rect 3928 -7339 3962 -7333
rect 4955 -7238 4989 -7204
rect 4565 -7338 4599 -7304
rect 5036 -7340 5070 -7306
rect 5171 -7407 5205 -7373
rect 6245 -7214 6279 -7180
rect 6694 -7407 6728 -7373
rect 6781 -7475 6815 -7441
rect 7198 -7407 7232 -7373
rect 7095 -7449 7127 -7441
rect 7127 -7449 7129 -7441
rect 7095 -7475 7129 -7449
rect 7356 -7298 7390 -7264
rect 7436 -7407 7470 -7373
rect 7604 -7299 7638 -7290
rect 7604 -7324 7609 -7299
rect 7609 -7324 7638 -7299
rect 7605 -7398 7639 -7364
rect 7515 -7475 7549 -7441
rect -2968 -7645 -2934 -7611
rect -2876 -7645 -2842 -7611
rect -2784 -7645 -2750 -7611
rect -2692 -7645 -2658 -7611
rect -2600 -7645 -2566 -7611
rect -2508 -7645 -2474 -7611
rect -2416 -7645 -2382 -7611
rect -2324 -7645 -2290 -7611
rect -2232 -7645 -2198 -7611
rect -2140 -7645 -2106 -7611
rect -2048 -7645 -2014 -7611
rect -1956 -7645 -1922 -7611
rect -1864 -7645 -1830 -7611
rect -1772 -7645 -1738 -7611
rect -1680 -7645 -1646 -7611
rect -1588 -7645 -1554 -7611
rect -1496 -7645 -1462 -7611
rect -1404 -7645 -1370 -7611
rect -1312 -7645 -1278 -7611
rect -1220 -7645 -1186 -7611
rect -1128 -7645 -1094 -7611
rect -1036 -7645 -1002 -7611
rect -944 -7645 -910 -7611
rect -852 -7645 -818 -7611
rect -760 -7645 -726 -7611
rect -668 -7645 -634 -7611
rect -576 -7645 -542 -7611
rect -484 -7645 -450 -7611
rect -392 -7645 -358 -7611
rect -300 -7645 -266 -7611
rect -208 -7645 -174 -7611
rect -116 -7645 -82 -7611
rect -24 -7645 10 -7611
rect 68 -7645 102 -7611
rect 160 -7645 194 -7611
rect 252 -7645 286 -7611
rect 344 -7645 378 -7611
rect 436 -7645 470 -7611
rect 528 -7645 562 -7611
rect 620 -7645 654 -7611
rect 712 -7645 746 -7611
rect 804 -7645 838 -7611
rect 896 -7645 930 -7611
rect 988 -7645 1022 -7611
rect 1080 -7645 1114 -7611
rect 1172 -7645 1206 -7611
rect 1264 -7645 1298 -7611
rect 1356 -7645 1390 -7611
rect 1448 -7645 1482 -7611
rect 1540 -7645 1574 -7611
rect 1632 -7645 1666 -7611
rect 1724 -7645 1758 -7611
rect 1816 -7645 1850 -7611
rect 1908 -7645 1942 -7611
rect 2000 -7645 2034 -7611
rect 2092 -7645 2126 -7611
rect 2184 -7645 2218 -7611
rect 2276 -7645 2310 -7611
rect 2368 -7645 2402 -7611
rect 2460 -7645 2494 -7611
rect 2552 -7645 2586 -7611
rect 2644 -7645 2678 -7611
rect 2736 -7645 2770 -7611
rect 2828 -7645 2862 -7611
rect 2920 -7645 2954 -7611
rect 3012 -7645 3046 -7611
rect 3104 -7645 3138 -7611
rect 3196 -7645 3230 -7611
rect 3288 -7645 3322 -7611
rect 3380 -7645 3414 -7611
rect 3472 -7645 3506 -7611
rect 3564 -7645 3598 -7611
rect 3656 -7645 3690 -7611
rect 3748 -7645 3782 -7611
rect 3840 -7645 3874 -7611
rect 3932 -7645 3966 -7611
rect 4024 -7645 4058 -7611
rect 4116 -7645 4150 -7611
rect 4208 -7645 4242 -7611
rect 4300 -7645 4334 -7611
rect 4392 -7645 4426 -7611
rect 4484 -7645 4518 -7611
rect 4576 -7645 4610 -7611
rect 4668 -7645 4702 -7611
rect 4760 -7645 4794 -7611
rect 4852 -7645 4886 -7611
rect 4944 -7645 4978 -7611
rect 5036 -7645 5070 -7611
rect 5128 -7645 5162 -7611
rect 5220 -7645 5254 -7611
rect 5312 -7645 5346 -7611
rect 5404 -7645 5438 -7611
rect 5496 -7645 5530 -7611
rect 5588 -7645 5622 -7611
rect 5680 -7645 5714 -7611
rect 5772 -7645 5806 -7611
rect 5864 -7645 5898 -7611
rect 5956 -7645 5990 -7611
rect 6048 -7645 6082 -7611
rect 6140 -7645 6174 -7611
rect 6232 -7645 6266 -7611
rect 6324 -7645 6358 -7611
rect 6416 -7645 6450 -7611
rect 6508 -7645 6542 -7611
rect 6600 -7645 6634 -7611
rect 6692 -7645 6726 -7611
rect 6784 -7645 6818 -7611
rect 6876 -7645 6910 -7611
rect 6968 -7645 7002 -7611
rect 7060 -7645 7094 -7611
rect 7152 -7645 7186 -7611
rect 7244 -7645 7278 -7611
rect 7336 -7645 7370 -7611
rect 7428 -7645 7462 -7611
rect 7520 -7645 7554 -7611
rect 7612 -7645 7646 -7611
rect 7704 -7645 7738 -7611
rect 7796 -7645 7830 -7611
rect 7888 -7645 7922 -7611
rect 7980 -7645 8014 -7611
rect 8072 -7645 8106 -7611
rect 8164 -7645 8198 -7611
rect 8256 -7645 8290 -7611
rect 8348 -7645 8382 -7611
rect 8440 -7645 8474 -7611
rect 8532 -7645 8566 -7611
rect 8624 -7645 8658 -7611
rect 8716 -7645 8750 -7611
rect 8808 -7645 8842 -7611
rect 8900 -7645 8934 -7611
rect 8992 -7645 9026 -7611
rect 9084 -7645 9118 -7611
rect 9176 -7645 9210 -7611
rect 9268 -7645 9302 -7611
rect 9360 -7645 9394 -7611
rect 9452 -7645 9486 -7611
rect 9544 -7645 9578 -7611
rect 9636 -7645 9670 -7611
rect 9728 -7645 9762 -7611
rect 9820 -7645 9854 -7611
rect 9912 -7645 9946 -7611
rect 10004 -7645 10038 -7611
rect 10096 -7645 10130 -7611
rect 10188 -7645 10222 -7611
rect 10280 -7645 10314 -7611
rect 10372 -7645 10406 -7611
rect 10464 -7645 10498 -7611
rect 10556 -7645 10590 -7611
rect 10648 -7645 10682 -7611
rect 10740 -7645 10774 -7611
rect 10832 -7645 10866 -7611
rect 10924 -7645 10958 -7611
rect 11016 -7645 11050 -7611
rect 11108 -7645 11142 -7611
rect 11200 -7645 11234 -7611
rect 11292 -7645 11326 -7611
rect 11384 -7645 11418 -7611
rect 11476 -7645 11510 -7611
rect 11568 -7645 11602 -7611
rect 11660 -7645 11694 -7611
rect 11752 -7645 11786 -7611
rect 11844 -7645 11878 -7611
rect 11936 -7645 11970 -7611
rect 12028 -7645 12062 -7611
rect 12120 -7645 12154 -7611
rect 12212 -7645 12246 -7611
rect 12304 -7645 12338 -7611
rect 12396 -7645 12430 -7611
rect 12488 -7645 12522 -7611
rect 12580 -7645 12614 -7611
rect 12672 -7645 12706 -7611
rect 12764 -7645 12798 -7611
rect 12856 -7645 12890 -7611
rect 12948 -7645 12982 -7611
rect 13040 -7645 13074 -7611
rect 13132 -7645 13166 -7611
rect 13224 -7645 13258 -7611
rect 13316 -7645 13350 -7611
rect 13408 -7645 13442 -7611
rect 13500 -7645 13534 -7611
rect 13592 -7645 13626 -7611
rect 13684 -7645 13718 -7611
rect 13776 -7645 13810 -7611
rect 13868 -7645 13902 -7611
rect 13960 -7645 13994 -7611
rect 14052 -7645 14086 -7611
rect 14144 -7645 14178 -7611
rect 14236 -7645 14270 -7611
rect 14328 -7645 14362 -7611
rect 14420 -7645 14454 -7611
rect 14512 -7645 14546 -7611
rect 14604 -7645 14638 -7611
rect 14696 -7645 14730 -7611
rect 14788 -7645 14822 -7611
rect 14880 -7645 14914 -7611
rect 14972 -7645 15006 -7611
rect 15064 -7645 15098 -7611
rect 15156 -7645 15190 -7611
rect 15248 -7645 15282 -7611
rect 15340 -7645 15374 -7611
rect 15432 -7645 15466 -7611
rect 15524 -7645 15558 -7611
rect 15616 -7645 15650 -7611
rect 15708 -7645 15742 -7611
rect 15800 -7645 15834 -7611
rect 15892 -7645 15926 -7611
rect 15984 -7645 16018 -7611
rect 16076 -7645 16110 -7611
rect 16168 -7645 16202 -7611
rect 16260 -7645 16294 -7611
rect 16352 -7645 16386 -7611
rect 16444 -7645 16478 -7611
rect 16536 -7645 16570 -7611
rect 16628 -7645 16662 -7611
rect -937 -7923 -903 -7918
rect -937 -7952 -903 -7923
rect -762 -7923 -728 -7917
rect -762 -7951 -735 -7923
rect -735 -7951 -728 -7923
rect -30 -7957 4 -7923
rect 106 -7957 140 -7923
rect 242 -7957 276 -7923
rect 434 -7995 468 -7961
rect -848 -8062 -814 -8028
rect -769 -8045 -766 -8028
rect -766 -8045 -735 -8028
rect -769 -8062 -735 -8045
rect 1076 -7957 1082 -7928
rect 1082 -7957 1110 -7928
rect 1076 -7962 1110 -7957
rect 1076 -8035 1110 -8001
rect 1171 -7956 1205 -7922
rect 1263 -7956 1297 -7922
rect 2369 -7923 2403 -7917
rect 2369 -7951 2396 -7923
rect 2396 -7951 2403 -7923
rect 3015 -7952 3049 -7918
rect 6876 -7923 6910 -7918
rect 6876 -7952 6904 -7923
rect 6904 -7952 6910 -7923
rect 7522 -7952 7556 -7918
rect 8164 -7923 8198 -7919
rect 8164 -7953 8192 -7923
rect 8192 -7953 8198 -7923
rect 8811 -7951 8845 -7917
rect 9453 -7923 9487 -7917
rect 9453 -7951 9480 -7923
rect 9480 -7951 9487 -7923
rect 10099 -7950 10133 -7916
rect 10741 -7923 10775 -7917
rect 10832 -7923 10866 -7917
rect 10925 -7923 10959 -7918
rect 11017 -7923 11051 -7918
rect 10741 -7951 10749 -7923
rect 10749 -7951 10775 -7923
rect 10832 -7951 10864 -7923
rect 10864 -7951 10866 -7923
rect 10925 -7952 10948 -7923
rect 10948 -7952 10959 -7923
rect 11017 -7952 11032 -7923
rect 11032 -7952 11051 -7923
rect 11129 -7918 11163 -7884
rect 11250 -7923 11284 -7915
rect 11344 -7923 11378 -7915
rect 11250 -7949 11284 -7923
rect 11344 -7949 11368 -7923
rect 11368 -7949 11378 -7923
rect -2968 -8189 -2934 -8155
rect -2876 -8189 -2842 -8155
rect -2784 -8189 -2750 -8155
rect -2692 -8189 -2658 -8155
rect -2600 -8189 -2566 -8155
rect -2508 -8189 -2474 -8155
rect -2416 -8189 -2382 -8155
rect -2324 -8189 -2290 -8155
rect -2232 -8189 -2198 -8155
rect -2140 -8189 -2106 -8155
rect -2048 -8189 -2014 -8155
rect -1956 -8189 -1922 -8155
rect -1864 -8189 -1830 -8155
rect -1772 -8189 -1738 -8155
rect -1680 -8189 -1646 -8155
rect -1588 -8189 -1554 -8155
rect -1496 -8189 -1462 -8155
rect -1404 -8189 -1370 -8155
rect -1312 -8189 -1278 -8155
rect -1220 -8189 -1186 -8155
rect -1128 -8189 -1094 -8155
rect -1036 -8189 -1002 -8155
rect -944 -8189 -910 -8155
rect -852 -8189 -818 -8155
rect -760 -8189 -726 -8155
rect -668 -8189 -634 -8155
rect -576 -8189 -542 -8155
rect -484 -8189 -450 -8155
rect -392 -8189 -358 -8155
rect -300 -8189 -266 -8155
rect -208 -8189 -174 -8155
rect -116 -8189 -82 -8155
rect -24 -8189 10 -8155
rect 68 -8189 102 -8155
rect 160 -8189 194 -8155
rect 252 -8189 286 -8155
rect 344 -8189 378 -8155
rect 436 -8189 470 -8155
rect 528 -8189 562 -8155
rect 620 -8189 654 -8155
rect 712 -8189 746 -8155
rect 804 -8189 838 -8155
rect 896 -8189 930 -8155
rect 988 -8189 1022 -8155
rect 1080 -8189 1114 -8155
rect 1172 -8189 1206 -8155
rect 1264 -8189 1298 -8155
rect 1356 -8189 1390 -8155
rect 1448 -8189 1482 -8155
rect 1540 -8189 1574 -8155
rect 1632 -8189 1666 -8155
rect 1724 -8189 1758 -8155
rect 1816 -8189 1850 -8155
rect 1908 -8189 1942 -8155
rect 2000 -8189 2034 -8155
rect 2092 -8189 2126 -8155
rect 2184 -8189 2218 -8155
rect 2276 -8189 2310 -8155
rect 2368 -8189 2402 -8155
rect 2460 -8189 2494 -8155
rect 2552 -8189 2586 -8155
rect 2644 -8189 2678 -8155
rect 2736 -8189 2770 -8155
rect 2828 -8189 2862 -8155
rect 2920 -8189 2954 -8155
rect 3012 -8189 3046 -8155
rect 3104 -8189 3138 -8155
rect 3196 -8189 3230 -8155
rect 3288 -8189 3322 -8155
rect 3380 -8189 3414 -8155
rect 3472 -8189 3506 -8155
rect 3564 -8189 3598 -8155
rect 3656 -8189 3690 -8155
rect 3748 -8189 3782 -8155
rect 3840 -8189 3874 -8155
rect 3932 -8189 3966 -8155
rect 4024 -8189 4058 -8155
rect 4116 -8189 4150 -8155
rect 4208 -8189 4242 -8155
rect 4300 -8189 4334 -8155
rect 4392 -8189 4426 -8155
rect 4484 -8189 4518 -8155
rect 4576 -8189 4610 -8155
rect 4668 -8189 4702 -8155
rect 4760 -8189 4794 -8155
rect 4852 -8189 4886 -8155
rect 4944 -8189 4978 -8155
rect 5036 -8189 5070 -8155
rect 5128 -8189 5162 -8155
rect 5220 -8189 5254 -8155
rect 5312 -8189 5346 -8155
rect 5404 -8189 5438 -8155
rect 5496 -8189 5530 -8155
rect 5588 -8189 5622 -8155
rect 5680 -8189 5714 -8155
rect 5772 -8189 5806 -8155
rect 5864 -8189 5898 -8155
rect 5956 -8189 5990 -8155
rect 6048 -8189 6082 -8155
rect 6140 -8189 6174 -8155
rect 6232 -8189 6266 -8155
rect 6324 -8189 6358 -8155
rect 6416 -8189 6450 -8155
rect 6508 -8189 6542 -8155
rect 6600 -8189 6634 -8155
rect 6692 -8189 6726 -8155
rect 6784 -8189 6818 -8155
rect 6876 -8189 6910 -8155
rect 6968 -8189 7002 -8155
rect 7060 -8189 7094 -8155
rect 7152 -8189 7186 -8155
rect 7244 -8189 7278 -8155
rect 7336 -8189 7370 -8155
rect 7428 -8189 7462 -8155
rect 7520 -8189 7554 -8155
rect 7612 -8189 7646 -8155
rect 7704 -8189 7738 -8155
rect 7796 -8189 7830 -8155
rect 7888 -8189 7922 -8155
rect 7980 -8189 8014 -8155
rect 8072 -8189 8106 -8155
rect 8164 -8189 8198 -8155
rect 8256 -8189 8290 -8155
rect 8348 -8189 8382 -8155
rect 8440 -8189 8474 -8155
rect 8532 -8189 8566 -8155
rect 8624 -8189 8658 -8155
rect 8716 -8189 8750 -8155
rect 8808 -8189 8842 -8155
rect 8900 -8189 8934 -8155
rect 8992 -8189 9026 -8155
rect 9084 -8189 9118 -8155
rect 9176 -8189 9210 -8155
rect 9268 -8189 9302 -8155
rect 9360 -8189 9394 -8155
rect 9452 -8189 9486 -8155
rect 9544 -8189 9578 -8155
rect 9636 -8189 9670 -8155
rect 9728 -8189 9762 -8155
rect 9820 -8189 9854 -8155
rect 9912 -8189 9946 -8155
rect 10004 -8189 10038 -8155
rect 10096 -8189 10130 -8155
rect 10188 -8189 10222 -8155
rect 10280 -8189 10314 -8155
rect 10372 -8189 10406 -8155
rect 10464 -8189 10498 -8155
rect 10556 -8189 10590 -8155
rect 10648 -8189 10682 -8155
rect 10740 -8189 10774 -8155
rect 10832 -8189 10866 -8155
rect 10924 -8189 10958 -8155
rect 11016 -8189 11050 -8155
rect 11108 -8189 11142 -8155
rect 11200 -8189 11234 -8155
rect 11292 -8189 11326 -8155
rect 11384 -8189 11418 -8155
rect 11476 -8189 11510 -8155
rect 11568 -8189 11602 -8155
rect 11660 -8189 11694 -8155
rect 11752 -8189 11786 -8155
rect 11844 -8189 11878 -8155
rect 11936 -8189 11970 -8155
rect 12028 -8189 12062 -8155
rect 12120 -8189 12154 -8155
rect 12212 -8189 12246 -8155
rect 12304 -8189 12338 -8155
rect 12396 -8189 12430 -8155
rect 12488 -8189 12522 -8155
rect 12580 -8189 12614 -8155
rect 12672 -8189 12706 -8155
rect 12764 -8189 12798 -8155
rect 12856 -8189 12890 -8155
rect 12948 -8189 12982 -8155
rect 13040 -8189 13074 -8155
rect 13132 -8189 13166 -8155
rect 13224 -8189 13258 -8155
rect 13316 -8189 13350 -8155
rect 13408 -8189 13442 -8155
rect 13500 -8189 13534 -8155
rect 13592 -8189 13626 -8155
rect 13684 -8189 13718 -8155
rect 13776 -8189 13810 -8155
rect 13868 -8189 13902 -8155
rect 13960 -8189 13994 -8155
rect 14052 -8189 14086 -8155
rect 14144 -8189 14178 -8155
rect 14236 -8189 14270 -8155
rect 14328 -8189 14362 -8155
rect 14420 -8189 14454 -8155
rect 14512 -8189 14546 -8155
rect 14604 -8189 14638 -8155
rect 14696 -8189 14730 -8155
rect 14788 -8189 14822 -8155
rect 14880 -8189 14914 -8155
rect 14972 -8189 15006 -8155
rect 15064 -8189 15098 -8155
rect 15156 -8189 15190 -8155
rect 15248 -8189 15282 -8155
rect 15340 -8189 15374 -8155
rect 15432 -8189 15466 -8155
rect 15524 -8189 15558 -8155
rect 15616 -8189 15650 -8155
rect 15708 -8189 15742 -8155
rect 15800 -8189 15834 -8155
rect 15892 -8189 15926 -8155
rect 15984 -8189 16018 -8155
rect 16076 -8189 16110 -8155
rect 16168 -8189 16202 -8155
rect 16260 -8189 16294 -8155
rect 16352 -8189 16386 -8155
rect 16444 -8189 16478 -8155
rect 16536 -8189 16570 -8155
rect 16628 -8189 16662 -8155
rect 433 -8462 467 -8428
rect 1052 -8421 1086 -8391
rect 1052 -8425 1086 -8421
rect 3012 -8425 3046 -8391
rect 3626 -8421 3628 -8391
rect 3628 -8421 3660 -8391
rect 3626 -8425 3660 -8421
rect 5586 -8425 5620 -8391
rect 6200 -8421 6204 -8391
rect 6204 -8421 6234 -8391
rect 6200 -8425 6234 -8421
rect 8160 -8425 8194 -8391
rect 8774 -8421 8780 -8391
rect 8780 -8421 8808 -8391
rect 8774 -8425 8808 -8421
rect 10737 -8427 10771 -8393
rect 11369 -8421 11390 -8394
rect 11390 -8421 11403 -8394
rect 11369 -8428 11403 -8421
rect 13685 -8387 13719 -8362
rect 13685 -8396 13692 -8387
rect 13692 -8396 13719 -8387
rect 15248 -8378 15282 -8344
rect 15340 -8379 15374 -8345
rect 15248 -8474 15282 -8440
rect 15341 -8474 15375 -8440
rect -2968 -8733 -2934 -8699
rect -2876 -8733 -2842 -8699
rect -2784 -8733 -2750 -8699
rect -2692 -8733 -2658 -8699
rect -2600 -8733 -2566 -8699
rect -2508 -8733 -2474 -8699
rect -2416 -8733 -2382 -8699
rect -2324 -8733 -2290 -8699
rect -2232 -8733 -2198 -8699
rect -2140 -8733 -2106 -8699
rect -2048 -8733 -2014 -8699
rect -1956 -8733 -1922 -8699
rect -1864 -8733 -1830 -8699
rect -1772 -8733 -1738 -8699
rect -1680 -8733 -1646 -8699
rect -1588 -8733 -1554 -8699
rect -1496 -8733 -1462 -8699
rect -1404 -8733 -1370 -8699
rect -1312 -8733 -1278 -8699
rect -1220 -8733 -1186 -8699
rect -1128 -8733 -1094 -8699
rect -1036 -8733 -1002 -8699
rect -944 -8733 -910 -8699
rect -852 -8733 -818 -8699
rect -760 -8733 -726 -8699
rect -668 -8733 -634 -8699
rect -576 -8733 -542 -8699
rect -484 -8733 -450 -8699
rect -392 -8733 -358 -8699
rect -300 -8733 -266 -8699
rect -208 -8733 -174 -8699
rect -116 -8733 -82 -8699
rect -24 -8733 10 -8699
rect 68 -8733 102 -8699
rect 160 -8733 194 -8699
rect 252 -8733 286 -8699
rect 344 -8733 378 -8699
rect 436 -8733 470 -8699
rect 528 -8733 562 -8699
rect 620 -8733 654 -8699
rect 712 -8733 746 -8699
rect 804 -8733 838 -8699
rect 896 -8733 930 -8699
rect 988 -8733 1022 -8699
rect 1080 -8733 1114 -8699
rect 1172 -8733 1206 -8699
rect 1264 -8733 1298 -8699
rect 1356 -8733 1390 -8699
rect 1448 -8733 1482 -8699
rect 1540 -8733 1574 -8699
rect 1632 -8733 1666 -8699
rect 1724 -8733 1758 -8699
rect 1816 -8733 1850 -8699
rect 1908 -8733 1942 -8699
rect 2000 -8733 2034 -8699
rect 2092 -8733 2126 -8699
rect 2184 -8733 2218 -8699
rect 2276 -8733 2310 -8699
rect 2368 -8733 2402 -8699
rect 2460 -8733 2494 -8699
rect 2552 -8733 2586 -8699
rect 2644 -8733 2678 -8699
rect 2736 -8733 2770 -8699
rect 2828 -8733 2862 -8699
rect 2920 -8733 2954 -8699
rect 3012 -8733 3046 -8699
rect 3104 -8733 3138 -8699
rect 3196 -8733 3230 -8699
rect 3288 -8733 3322 -8699
rect 3380 -8733 3414 -8699
rect 3472 -8733 3506 -8699
rect 3564 -8733 3598 -8699
rect 3656 -8733 3690 -8699
rect 3748 -8733 3782 -8699
rect 3840 -8733 3874 -8699
rect 3932 -8733 3966 -8699
rect 4024 -8733 4058 -8699
rect 4116 -8733 4150 -8699
rect 4208 -8733 4242 -8699
rect 4300 -8733 4334 -8699
rect 4392 -8733 4426 -8699
rect 4484 -8733 4518 -8699
rect 4576 -8733 4610 -8699
rect 4668 -8733 4702 -8699
rect 4760 -8733 4794 -8699
rect 4852 -8733 4886 -8699
rect 4944 -8733 4978 -8699
rect 5036 -8733 5070 -8699
rect 5128 -8733 5162 -8699
rect 5220 -8733 5254 -8699
rect 5312 -8733 5346 -8699
rect 5404 -8733 5438 -8699
rect 5496 -8733 5530 -8699
rect 5588 -8733 5622 -8699
rect 5680 -8733 5714 -8699
rect 5772 -8733 5806 -8699
rect 5864 -8733 5898 -8699
rect 5956 -8733 5990 -8699
rect 6048 -8733 6082 -8699
rect 6140 -8733 6174 -8699
rect 6232 -8733 6266 -8699
rect 6324 -8733 6358 -8699
rect 6416 -8733 6450 -8699
rect 6508 -8733 6542 -8699
rect 6600 -8733 6634 -8699
rect 6692 -8733 6726 -8699
rect 6784 -8733 6818 -8699
rect 6876 -8733 6910 -8699
rect 6968 -8733 7002 -8699
rect 7060 -8733 7094 -8699
rect 7152 -8733 7186 -8699
rect 7244 -8733 7278 -8699
rect 7336 -8733 7370 -8699
rect 7428 -8733 7462 -8699
rect 7520 -8733 7554 -8699
rect 7612 -8733 7646 -8699
rect 7704 -8733 7738 -8699
rect 7796 -8733 7830 -8699
rect 7888 -8733 7922 -8699
rect 7980 -8733 8014 -8699
rect 8072 -8733 8106 -8699
rect 8164 -8733 8198 -8699
rect 8256 -8733 8290 -8699
rect 8348 -8733 8382 -8699
rect 8440 -8733 8474 -8699
rect 8532 -8733 8566 -8699
rect 8624 -8733 8658 -8699
rect 8716 -8733 8750 -8699
rect 8808 -8733 8842 -8699
rect 8900 -8733 8934 -8699
rect 8992 -8733 9026 -8699
rect 9084 -8733 9118 -8699
rect 9176 -8733 9210 -8699
rect 9268 -8733 9302 -8699
rect 9360 -8733 9394 -8699
rect 9452 -8733 9486 -8699
rect 9544 -8733 9578 -8699
rect 9636 -8733 9670 -8699
rect 9728 -8733 9762 -8699
rect 9820 -8733 9854 -8699
rect 9912 -8733 9946 -8699
rect 10004 -8733 10038 -8699
rect 10096 -8733 10130 -8699
rect 10188 -8733 10222 -8699
rect 10280 -8733 10314 -8699
rect 10372 -8733 10406 -8699
rect 10464 -8733 10498 -8699
rect 10556 -8733 10590 -8699
rect 10648 -8733 10682 -8699
rect 10740 -8733 10774 -8699
rect 10832 -8733 10866 -8699
rect 10924 -8733 10958 -8699
rect 11016 -8733 11050 -8699
rect 11108 -8733 11142 -8699
rect 11200 -8733 11234 -8699
rect 11292 -8733 11326 -8699
rect 11384 -8733 11418 -8699
rect 11476 -8733 11510 -8699
rect 11568 -8733 11602 -8699
rect 11660 -8733 11694 -8699
rect 11752 -8733 11786 -8699
rect 11844 -8733 11878 -8699
rect 11936 -8733 11970 -8699
rect 12028 -8733 12062 -8699
rect 12120 -8733 12154 -8699
rect 12212 -8733 12246 -8699
rect 12304 -8733 12338 -8699
rect 12396 -8733 12430 -8699
rect 12488 -8733 12522 -8699
rect 12580 -8733 12614 -8699
rect 12672 -8733 12706 -8699
rect 12764 -8733 12798 -8699
rect 12856 -8733 12890 -8699
rect 12948 -8733 12982 -8699
rect 13040 -8733 13074 -8699
rect 13132 -8733 13166 -8699
rect 13224 -8733 13258 -8699
rect 13316 -8733 13350 -8699
rect 13408 -8733 13442 -8699
rect 13500 -8733 13534 -8699
rect 13592 -8733 13626 -8699
rect 13684 -8733 13718 -8699
rect 13776 -8733 13810 -8699
rect 13868 -8733 13902 -8699
rect 13960 -8733 13994 -8699
rect 14052 -8733 14086 -8699
rect 14144 -8733 14178 -8699
rect 14236 -8733 14270 -8699
rect 14328 -8733 14362 -8699
rect 14420 -8733 14454 -8699
rect 14512 -8733 14546 -8699
rect 14604 -8733 14638 -8699
rect 14696 -8733 14730 -8699
rect 14788 -8733 14822 -8699
rect 14880 -8733 14914 -8699
rect 14972 -8733 15006 -8699
rect 15064 -8733 15098 -8699
rect 15156 -8733 15190 -8699
rect 15248 -8733 15282 -8699
rect 15340 -8733 15374 -8699
rect 15432 -8733 15466 -8699
rect 15524 -8733 15558 -8699
rect 15616 -8733 15650 -8699
rect 15708 -8733 15742 -8699
rect 15800 -8733 15834 -8699
rect 15892 -8733 15926 -8699
rect 15984 -8733 16018 -8699
rect 16076 -8733 16110 -8699
rect 16168 -8733 16202 -8699
rect 16260 -8733 16294 -8699
rect 16352 -8733 16386 -8699
rect 16444 -8733 16478 -8699
rect 16536 -8733 16570 -8699
rect 16628 -8733 16662 -8699
rect 432 -9011 466 -9008
rect 432 -9042 464 -9011
rect 464 -9042 466 -9011
rect 1082 -9039 1116 -9005
rect 3042 -9011 3076 -9005
rect 3042 -9039 3074 -9011
rect 3074 -9039 3076 -9011
rect 3656 -9039 3690 -9005
rect 5616 -9011 5650 -9005
rect 5616 -9039 5650 -9011
rect 6230 -9039 6264 -9005
rect 8190 -9011 8224 -9005
rect 8190 -9039 8192 -9011
rect 8192 -9039 8224 -9011
rect 8804 -9039 8838 -9005
rect 10764 -9011 10798 -9005
rect 10764 -9039 10768 -9011
rect 10768 -9039 10798 -9011
rect 11387 -9005 11421 -8971
rect 12558 -9011 12592 -9008
rect 12642 -9011 12676 -9008
rect 12739 -9011 12773 -9008
rect 12836 -9011 12870 -9008
rect 12942 -9011 12976 -9008
rect 12558 -9042 12574 -9011
rect 12574 -9042 12592 -9011
rect 12642 -9042 12676 -9011
rect 12739 -9042 12744 -9011
rect 12744 -9042 12773 -9011
rect 12836 -9042 12846 -9011
rect 12846 -9042 12870 -9011
rect 12942 -9042 12948 -9011
rect 12948 -9042 12976 -9011
rect 13038 -9035 13072 -9001
rect 13038 -9107 13072 -9073
rect 15248 -8988 15282 -8954
rect 15340 -8989 15374 -8955
rect 13684 -9045 13692 -9038
rect 13692 -9045 13718 -9038
rect 13684 -9072 13718 -9045
rect 15248 -9084 15282 -9050
rect 15341 -9084 15375 -9050
rect -2968 -9277 -2934 -9243
rect -2876 -9277 -2842 -9243
rect -2784 -9277 -2750 -9243
rect -2692 -9277 -2658 -9243
rect -2600 -9277 -2566 -9243
rect -2508 -9277 -2474 -9243
rect -2416 -9277 -2382 -9243
rect -2324 -9277 -2290 -9243
rect -2232 -9277 -2198 -9243
rect -2140 -9277 -2106 -9243
rect -2048 -9277 -2014 -9243
rect -1956 -9277 -1922 -9243
rect -1864 -9277 -1830 -9243
rect -1772 -9277 -1738 -9243
rect -1680 -9277 -1646 -9243
rect -1588 -9277 -1554 -9243
rect -1496 -9277 -1462 -9243
rect -1404 -9277 -1370 -9243
rect -1312 -9277 -1278 -9243
rect -1220 -9277 -1186 -9243
rect -1128 -9277 -1094 -9243
rect -1036 -9277 -1002 -9243
rect -944 -9277 -910 -9243
rect -852 -9277 -818 -9243
rect -760 -9277 -726 -9243
rect -668 -9277 -634 -9243
rect -576 -9277 -542 -9243
rect -484 -9277 -450 -9243
rect -392 -9277 -358 -9243
rect -300 -9277 -266 -9243
rect -208 -9277 -174 -9243
rect -116 -9277 -82 -9243
rect -24 -9277 10 -9243
rect 68 -9277 102 -9243
rect 160 -9277 194 -9243
rect 252 -9277 286 -9243
rect 344 -9277 378 -9243
rect 436 -9277 470 -9243
rect 528 -9277 562 -9243
rect 620 -9277 654 -9243
rect 712 -9277 746 -9243
rect 804 -9277 838 -9243
rect 896 -9277 930 -9243
rect 988 -9277 1022 -9243
rect 1080 -9277 1114 -9243
rect 1172 -9277 1206 -9243
rect 1264 -9277 1298 -9243
rect 1356 -9277 1390 -9243
rect 1448 -9277 1482 -9243
rect 1540 -9277 1574 -9243
rect 1632 -9277 1666 -9243
rect 1724 -9277 1758 -9243
rect 1816 -9277 1850 -9243
rect 1908 -9277 1942 -9243
rect 2000 -9277 2034 -9243
rect 2092 -9277 2126 -9243
rect 2184 -9277 2218 -9243
rect 2276 -9277 2310 -9243
rect 2368 -9277 2402 -9243
rect 2460 -9277 2494 -9243
rect 2552 -9277 2586 -9243
rect 2644 -9277 2678 -9243
rect 2736 -9277 2770 -9243
rect 2828 -9277 2862 -9243
rect 2920 -9277 2954 -9243
rect 3012 -9277 3046 -9243
rect 3104 -9277 3138 -9243
rect 3196 -9277 3230 -9243
rect 3288 -9277 3322 -9243
rect 3380 -9277 3414 -9243
rect 3472 -9277 3506 -9243
rect 3564 -9277 3598 -9243
rect 3656 -9277 3690 -9243
rect 3748 -9277 3782 -9243
rect 3840 -9277 3874 -9243
rect 3932 -9277 3966 -9243
rect 4024 -9277 4058 -9243
rect 4116 -9277 4150 -9243
rect 4208 -9277 4242 -9243
rect 4300 -9277 4334 -9243
rect 4392 -9277 4426 -9243
rect 4484 -9277 4518 -9243
rect 4576 -9277 4610 -9243
rect 4668 -9277 4702 -9243
rect 4760 -9277 4794 -9243
rect 4852 -9277 4886 -9243
rect 4944 -9277 4978 -9243
rect 5036 -9277 5070 -9243
rect 5128 -9277 5162 -9243
rect 5220 -9277 5254 -9243
rect 5312 -9277 5346 -9243
rect 5404 -9277 5438 -9243
rect 5496 -9277 5530 -9243
rect 5588 -9277 5622 -9243
rect 5680 -9277 5714 -9243
rect 5772 -9277 5806 -9243
rect 5864 -9277 5898 -9243
rect 5956 -9277 5990 -9243
rect 6048 -9277 6082 -9243
rect 6140 -9277 6174 -9243
rect 6232 -9277 6266 -9243
rect 6324 -9277 6358 -9243
rect 6416 -9277 6450 -9243
rect 6508 -9277 6542 -9243
rect 6600 -9277 6634 -9243
rect 6692 -9277 6726 -9243
rect 6784 -9277 6818 -9243
rect 6876 -9277 6910 -9243
rect 6968 -9277 7002 -9243
rect 7060 -9277 7094 -9243
rect 7152 -9277 7186 -9243
rect 7244 -9277 7278 -9243
rect 7336 -9277 7370 -9243
rect 7428 -9277 7462 -9243
rect 7520 -9277 7554 -9243
rect 7612 -9277 7646 -9243
rect 7704 -9277 7738 -9243
rect 7796 -9277 7830 -9243
rect 7888 -9277 7922 -9243
rect 7980 -9277 8014 -9243
rect 8072 -9277 8106 -9243
rect 8164 -9277 8198 -9243
rect 8256 -9277 8290 -9243
rect 8348 -9277 8382 -9243
rect 8440 -9277 8474 -9243
rect 8532 -9277 8566 -9243
rect 8624 -9277 8658 -9243
rect 8716 -9277 8750 -9243
rect 8808 -9277 8842 -9243
rect 8900 -9277 8934 -9243
rect 8992 -9277 9026 -9243
rect 9084 -9277 9118 -9243
rect 9176 -9277 9210 -9243
rect 9268 -9277 9302 -9243
rect 9360 -9277 9394 -9243
rect 9452 -9277 9486 -9243
rect 9544 -9277 9578 -9243
rect 9636 -9277 9670 -9243
rect 9728 -9277 9762 -9243
rect 9820 -9277 9854 -9243
rect 9912 -9277 9946 -9243
rect 10004 -9277 10038 -9243
rect 10096 -9277 10130 -9243
rect 10188 -9277 10222 -9243
rect 10280 -9277 10314 -9243
rect 10372 -9277 10406 -9243
rect 10464 -9277 10498 -9243
rect 10556 -9277 10590 -9243
rect 10648 -9277 10682 -9243
rect 10740 -9277 10774 -9243
rect 10832 -9277 10866 -9243
rect 10924 -9277 10958 -9243
rect 11016 -9277 11050 -9243
rect 11108 -9277 11142 -9243
rect 11200 -9277 11234 -9243
rect 11292 -9277 11326 -9243
rect 11384 -9277 11418 -9243
rect 11476 -9277 11510 -9243
rect 11568 -9277 11602 -9243
rect 11660 -9277 11694 -9243
rect 11752 -9277 11786 -9243
rect 11844 -9277 11878 -9243
rect 11936 -9277 11970 -9243
rect 12028 -9277 12062 -9243
rect 12120 -9277 12154 -9243
rect 12212 -9277 12246 -9243
rect 12304 -9277 12338 -9243
rect 12396 -9277 12430 -9243
rect 12488 -9277 12522 -9243
rect 12580 -9277 12614 -9243
rect 12672 -9277 12706 -9243
rect 12764 -9277 12798 -9243
rect 12856 -9277 12890 -9243
rect 12948 -9277 12982 -9243
rect 13040 -9277 13074 -9243
rect 13132 -9277 13166 -9243
rect 13224 -9277 13258 -9243
rect 13316 -9277 13350 -9243
rect 13408 -9277 13442 -9243
rect 13500 -9277 13534 -9243
rect 13592 -9277 13626 -9243
rect 13684 -9277 13718 -9243
rect 13776 -9277 13810 -9243
rect 13868 -9277 13902 -9243
rect 13960 -9277 13994 -9243
rect 14052 -9277 14086 -9243
rect 14144 -9277 14178 -9243
rect 14236 -9277 14270 -9243
rect 14328 -9277 14362 -9243
rect 14420 -9277 14454 -9243
rect 14512 -9277 14546 -9243
rect 14604 -9277 14638 -9243
rect 14696 -9277 14730 -9243
rect 14788 -9277 14822 -9243
rect 14880 -9277 14914 -9243
rect 14972 -9277 15006 -9243
rect 15064 -9277 15098 -9243
rect 15156 -9277 15190 -9243
rect 15248 -9277 15282 -9243
rect 15340 -9277 15374 -9243
rect 15432 -9277 15466 -9243
rect 15524 -9277 15558 -9243
rect 15616 -9277 15650 -9243
rect 15708 -9277 15742 -9243
rect 15800 -9277 15834 -9243
rect 15892 -9277 15926 -9243
rect 15984 -9277 16018 -9243
rect 16076 -9277 16110 -9243
rect 16168 -9277 16202 -9243
rect 16260 -9277 16294 -9243
rect 16352 -9277 16386 -9243
rect 16444 -9277 16478 -9243
rect 16536 -9277 16570 -9243
rect 16628 -9277 16662 -9243
rect -856 -9550 -822 -9516
rect -210 -9509 -202 -9481
rect -202 -9509 -176 -9481
rect -210 -9515 -176 -9509
rect 432 -9550 466 -9516
rect 1054 -9509 1086 -9482
rect 1086 -9509 1088 -9482
rect 1054 -9516 1088 -9509
rect 3014 -9516 3048 -9482
rect 3628 -9509 3662 -9482
rect 3628 -9516 3662 -9509
rect 5588 -9516 5622 -9482
rect 6202 -9509 6204 -9482
rect 6204 -9509 6236 -9482
rect 6202 -9516 6236 -9509
rect 8162 -9516 8196 -9482
rect 8776 -9509 8780 -9482
rect 8780 -9509 8810 -9482
rect 8776 -9516 8810 -9509
rect 10736 -9516 10770 -9482
rect 11386 -9509 11390 -9479
rect 11390 -9509 11420 -9479
rect 11386 -9513 11420 -9509
rect 13685 -9475 13719 -9448
rect 13685 -9482 13692 -9475
rect 13692 -9482 13719 -9475
rect 15248 -9466 15282 -9432
rect 15340 -9467 15374 -9433
rect 15248 -9562 15282 -9528
rect 15341 -9562 15375 -9528
rect -2968 -9821 -2934 -9787
rect -2876 -9821 -2842 -9787
rect -2784 -9821 -2750 -9787
rect -2692 -9821 -2658 -9787
rect -2600 -9821 -2566 -9787
rect -2508 -9821 -2474 -9787
rect -2416 -9821 -2382 -9787
rect -2324 -9821 -2290 -9787
rect -2232 -9821 -2198 -9787
rect -2140 -9821 -2106 -9787
rect -2048 -9821 -2014 -9787
rect -1956 -9821 -1922 -9787
rect -1864 -9821 -1830 -9787
rect -1772 -9821 -1738 -9787
rect -1680 -9821 -1646 -9787
rect -1588 -9821 -1554 -9787
rect -1496 -9821 -1462 -9787
rect -1404 -9821 -1370 -9787
rect -1312 -9821 -1278 -9787
rect -1220 -9821 -1186 -9787
rect -1128 -9821 -1094 -9787
rect -1036 -9821 -1002 -9787
rect -944 -9821 -910 -9787
rect -852 -9821 -818 -9787
rect -760 -9821 -726 -9787
rect -668 -9821 -634 -9787
rect -576 -9821 -542 -9787
rect -484 -9821 -450 -9787
rect -392 -9821 -358 -9787
rect -300 -9821 -266 -9787
rect -208 -9821 -174 -9787
rect -116 -9821 -82 -9787
rect -24 -9821 10 -9787
rect 68 -9821 102 -9787
rect 160 -9821 194 -9787
rect 252 -9821 286 -9787
rect 344 -9821 378 -9787
rect 436 -9821 470 -9787
rect 528 -9821 562 -9787
rect 620 -9821 654 -9787
rect 712 -9821 746 -9787
rect 804 -9821 838 -9787
rect 896 -9821 930 -9787
rect 988 -9821 1022 -9787
rect 1080 -9821 1114 -9787
rect 1172 -9821 1206 -9787
rect 1264 -9821 1298 -9787
rect 1356 -9821 1390 -9787
rect 1448 -9821 1482 -9787
rect 1540 -9821 1574 -9787
rect 1632 -9821 1666 -9787
rect 1724 -9821 1758 -9787
rect 1816 -9821 1850 -9787
rect 1908 -9821 1942 -9787
rect 2000 -9821 2034 -9787
rect 2092 -9821 2126 -9787
rect 2184 -9821 2218 -9787
rect 2276 -9821 2310 -9787
rect 2368 -9821 2402 -9787
rect 2460 -9821 2494 -9787
rect 2552 -9821 2586 -9787
rect 2644 -9821 2678 -9787
rect 2736 -9821 2770 -9787
rect 2828 -9821 2862 -9787
rect 2920 -9821 2954 -9787
rect 3012 -9821 3046 -9787
rect 3104 -9821 3138 -9787
rect 3196 -9821 3230 -9787
rect 3288 -9821 3322 -9787
rect 3380 -9821 3414 -9787
rect 3472 -9821 3506 -9787
rect 3564 -9821 3598 -9787
rect 3656 -9821 3690 -9787
rect 3748 -9821 3782 -9787
rect 3840 -9821 3874 -9787
rect 3932 -9821 3966 -9787
rect 4024 -9821 4058 -9787
rect 4116 -9821 4150 -9787
rect 4208 -9821 4242 -9787
rect 4300 -9821 4334 -9787
rect 4392 -9821 4426 -9787
rect 4484 -9821 4518 -9787
rect 4576 -9821 4610 -9787
rect 4668 -9821 4702 -9787
rect 4760 -9821 4794 -9787
rect 4852 -9821 4886 -9787
rect 4944 -9821 4978 -9787
rect 5036 -9821 5070 -9787
rect 5128 -9821 5162 -9787
rect 5220 -9821 5254 -9787
rect 5312 -9821 5346 -9787
rect 5404 -9821 5438 -9787
rect 5496 -9821 5530 -9787
rect 5588 -9821 5622 -9787
rect 5680 -9821 5714 -9787
rect 5772 -9821 5806 -9787
rect 5864 -9821 5898 -9787
rect 5956 -9821 5990 -9787
rect 6048 -9821 6082 -9787
rect 6140 -9821 6174 -9787
rect 6232 -9821 6266 -9787
rect 6324 -9821 6358 -9787
rect 6416 -9821 6450 -9787
rect 6508 -9821 6542 -9787
rect 6600 -9821 6634 -9787
rect 6692 -9821 6726 -9787
rect 6784 -9821 6818 -9787
rect 6876 -9821 6910 -9787
rect 6968 -9821 7002 -9787
rect 7060 -9821 7094 -9787
rect 7152 -9821 7186 -9787
rect 7244 -9821 7278 -9787
rect 7336 -9821 7370 -9787
rect 7428 -9821 7462 -9787
rect 7520 -9821 7554 -9787
rect 7612 -9821 7646 -9787
rect 7704 -9821 7738 -9787
rect 7796 -9821 7830 -9787
rect 7888 -9821 7922 -9787
rect 7980 -9821 8014 -9787
rect 8072 -9821 8106 -9787
rect 8164 -9821 8198 -9787
rect 8256 -9821 8290 -9787
rect 8348 -9821 8382 -9787
rect 8440 -9821 8474 -9787
rect 8532 -9821 8566 -9787
rect 8624 -9821 8658 -9787
rect 8716 -9821 8750 -9787
rect 8808 -9821 8842 -9787
rect 8900 -9821 8934 -9787
rect 8992 -9821 9026 -9787
rect 9084 -9821 9118 -9787
rect 9176 -9821 9210 -9787
rect 9268 -9821 9302 -9787
rect 9360 -9821 9394 -9787
rect 9452 -9821 9486 -9787
rect 9544 -9821 9578 -9787
rect 9636 -9821 9670 -9787
rect 9728 -9821 9762 -9787
rect 9820 -9821 9854 -9787
rect 9912 -9821 9946 -9787
rect 10004 -9821 10038 -9787
rect 10096 -9821 10130 -9787
rect 10188 -9821 10222 -9787
rect 10280 -9821 10314 -9787
rect 10372 -9821 10406 -9787
rect 10464 -9821 10498 -9787
rect 10556 -9821 10590 -9787
rect 10648 -9821 10682 -9787
rect 10740 -9821 10774 -9787
rect 10832 -9821 10866 -9787
rect 10924 -9821 10958 -9787
rect 11016 -9821 11050 -9787
rect 11108 -9821 11142 -9787
rect 11200 -9821 11234 -9787
rect 11292 -9821 11326 -9787
rect 11384 -9821 11418 -9787
rect 11476 -9821 11510 -9787
rect 11568 -9821 11602 -9787
rect 11660 -9821 11694 -9787
rect 11752 -9821 11786 -9787
rect 11844 -9821 11878 -9787
rect 11936 -9821 11970 -9787
rect 12028 -9821 12062 -9787
rect 12120 -9821 12154 -9787
rect 12212 -9821 12246 -9787
rect 12304 -9821 12338 -9787
rect 12396 -9821 12430 -9787
rect 12488 -9821 12522 -9787
rect 12580 -9821 12614 -9787
rect 12672 -9821 12706 -9787
rect 12764 -9821 12798 -9787
rect 12856 -9821 12890 -9787
rect 12948 -9821 12982 -9787
rect 13040 -9821 13074 -9787
rect 13132 -9821 13166 -9787
rect 13224 -9821 13258 -9787
rect 13316 -9821 13350 -9787
rect 13408 -9821 13442 -9787
rect 13500 -9821 13534 -9787
rect 13592 -9821 13626 -9787
rect 13684 -9821 13718 -9787
rect 13776 -9821 13810 -9787
rect 13868 -9821 13902 -9787
rect 13960 -9821 13994 -9787
rect 14052 -9821 14086 -9787
rect 14144 -9821 14178 -9787
rect 14236 -9821 14270 -9787
rect 14328 -9821 14362 -9787
rect 14420 -9821 14454 -9787
rect 14512 -9821 14546 -9787
rect 14604 -9821 14638 -9787
rect 14696 -9821 14730 -9787
rect 14788 -9821 14822 -9787
rect 14880 -9821 14914 -9787
rect 14972 -9821 15006 -9787
rect 15064 -9821 15098 -9787
rect 15156 -9821 15190 -9787
rect 15248 -9821 15282 -9787
rect 15340 -9821 15374 -9787
rect 15432 -9821 15466 -9787
rect 15524 -9821 15558 -9787
rect 15616 -9821 15650 -9787
rect 15708 -9821 15742 -9787
rect 15800 -9821 15834 -9787
rect 15892 -9821 15926 -9787
rect 15984 -9821 16018 -9787
rect 16076 -9821 16110 -9787
rect 16168 -9821 16202 -9787
rect 16260 -9821 16294 -9787
rect 16352 -9821 16386 -9787
rect 16444 -9821 16478 -9787
rect 16536 -9821 16570 -9787
rect 16628 -9821 16662 -9787
rect 436 -10099 470 -10096
rect 436 -10130 464 -10099
rect 464 -10130 470 -10099
rect 1081 -10128 1115 -10094
rect 3041 -10099 3075 -10094
rect 3041 -10128 3074 -10099
rect 3074 -10128 3075 -10099
rect 3655 -10128 3689 -10094
rect 5615 -10099 5649 -10094
rect 5615 -10128 5616 -10099
rect 5616 -10128 5649 -10099
rect 6229 -10128 6263 -10094
rect 8189 -10099 8223 -10094
rect 8189 -10128 8192 -10099
rect 8192 -10128 8223 -10099
rect 8806 -10128 8840 -10094
rect 10763 -10099 10797 -10094
rect 10763 -10128 10768 -10099
rect 10768 -10128 10797 -10099
rect 11386 -10095 11420 -10061
rect 12480 -10057 12514 -10023
rect 12480 -10131 12514 -10097
rect 12568 -10099 12602 -10095
rect 12659 -10099 12693 -10095
rect 12765 -10099 12799 -10095
rect 12858 -10099 12892 -10093
rect 12942 -10099 12976 -10093
rect 12568 -10129 12574 -10099
rect 12574 -10129 12602 -10099
rect 12659 -10129 12676 -10099
rect 12676 -10129 12693 -10099
rect 12765 -10129 12778 -10099
rect 12778 -10129 12799 -10099
rect 12858 -10127 12880 -10099
rect 12880 -10127 12892 -10099
rect 12942 -10127 12948 -10099
rect 12948 -10127 12976 -10099
rect 13039 -10116 13073 -10082
rect 12480 -10203 12514 -10169
rect 13042 -10193 13076 -10159
rect 15248 -10076 15282 -10042
rect 15340 -10076 15374 -10042
rect 13685 -10133 13692 -10126
rect 13692 -10133 13719 -10126
rect 13685 -10160 13719 -10133
rect 15248 -10172 15282 -10138
rect 15341 -10172 15375 -10138
rect -2968 -10365 -2934 -10331
rect -2876 -10365 -2842 -10331
rect -2784 -10365 -2750 -10331
rect -2692 -10365 -2658 -10331
rect -2600 -10365 -2566 -10331
rect -2508 -10365 -2474 -10331
rect -2416 -10365 -2382 -10331
rect -2324 -10365 -2290 -10331
rect -2232 -10365 -2198 -10331
rect -2140 -10365 -2106 -10331
rect -2048 -10365 -2014 -10331
rect -1956 -10365 -1922 -10331
rect -1864 -10365 -1830 -10331
rect -1772 -10365 -1738 -10331
rect -1680 -10365 -1646 -10331
rect -1588 -10365 -1554 -10331
rect -1496 -10365 -1462 -10331
rect -1404 -10365 -1370 -10331
rect -1312 -10365 -1278 -10331
rect -1220 -10365 -1186 -10331
rect -1128 -10365 -1094 -10331
rect -1036 -10365 -1002 -10331
rect -944 -10365 -910 -10331
rect -852 -10365 -818 -10331
rect -760 -10365 -726 -10331
rect -668 -10365 -634 -10331
rect -576 -10365 -542 -10331
rect -484 -10365 -450 -10331
rect -392 -10365 -358 -10331
rect -300 -10365 -266 -10331
rect -208 -10365 -174 -10331
rect -116 -10365 -82 -10331
rect -24 -10365 10 -10331
rect 68 -10365 102 -10331
rect 160 -10365 194 -10331
rect 252 -10365 286 -10331
rect 344 -10365 378 -10331
rect 436 -10365 470 -10331
rect 528 -10365 562 -10331
rect 620 -10365 654 -10331
rect 712 -10365 746 -10331
rect 804 -10365 838 -10331
rect 896 -10365 930 -10331
rect 988 -10365 1022 -10331
rect 1080 -10365 1114 -10331
rect 1172 -10365 1206 -10331
rect 1264 -10365 1298 -10331
rect 1356 -10365 1390 -10331
rect 1448 -10365 1482 -10331
rect 1540 -10365 1574 -10331
rect 1632 -10365 1666 -10331
rect 1724 -10365 1758 -10331
rect 1816 -10365 1850 -10331
rect 1908 -10365 1942 -10331
rect 2000 -10365 2034 -10331
rect 2092 -10365 2126 -10331
rect 2184 -10365 2218 -10331
rect 2276 -10365 2310 -10331
rect 2368 -10365 2402 -10331
rect 2460 -10365 2494 -10331
rect 2552 -10365 2586 -10331
rect 2644 -10365 2678 -10331
rect 2736 -10365 2770 -10331
rect 2828 -10365 2862 -10331
rect 2920 -10365 2954 -10331
rect 3012 -10365 3046 -10331
rect 3104 -10365 3138 -10331
rect 3196 -10365 3230 -10331
rect 3288 -10365 3322 -10331
rect 3380 -10365 3414 -10331
rect 3472 -10365 3506 -10331
rect 3564 -10365 3598 -10331
rect 3656 -10365 3690 -10331
rect 3748 -10365 3782 -10331
rect 3840 -10365 3874 -10331
rect 3932 -10365 3966 -10331
rect 4024 -10365 4058 -10331
rect 4116 -10365 4150 -10331
rect 4208 -10365 4242 -10331
rect 4300 -10365 4334 -10331
rect 4392 -10365 4426 -10331
rect 4484 -10365 4518 -10331
rect 4576 -10365 4610 -10331
rect 4668 -10365 4702 -10331
rect 4760 -10365 4794 -10331
rect 4852 -10365 4886 -10331
rect 4944 -10365 4978 -10331
rect 5036 -10365 5070 -10331
rect 5128 -10365 5162 -10331
rect 5220 -10365 5254 -10331
rect 5312 -10365 5346 -10331
rect 5404 -10365 5438 -10331
rect 5496 -10365 5530 -10331
rect 5588 -10365 5622 -10331
rect 5680 -10365 5714 -10331
rect 5772 -10365 5806 -10331
rect 5864 -10365 5898 -10331
rect 5956 -10365 5990 -10331
rect 6048 -10365 6082 -10331
rect 6140 -10365 6174 -10331
rect 6232 -10365 6266 -10331
rect 6324 -10365 6358 -10331
rect 6416 -10365 6450 -10331
rect 6508 -10365 6542 -10331
rect 6600 -10365 6634 -10331
rect 6692 -10365 6726 -10331
rect 6784 -10365 6818 -10331
rect 6876 -10365 6910 -10331
rect 6968 -10365 7002 -10331
rect 7060 -10365 7094 -10331
rect 7152 -10365 7186 -10331
rect 7244 -10365 7278 -10331
rect 7336 -10365 7370 -10331
rect 7428 -10365 7462 -10331
rect 7520 -10365 7554 -10331
rect 7612 -10365 7646 -10331
rect 7704 -10365 7738 -10331
rect 7796 -10365 7830 -10331
rect 7888 -10365 7922 -10331
rect 7980 -10365 8014 -10331
rect 8072 -10365 8106 -10331
rect 8164 -10365 8198 -10331
rect 8256 -10365 8290 -10331
rect 8348 -10365 8382 -10331
rect 8440 -10365 8474 -10331
rect 8532 -10365 8566 -10331
rect 8624 -10365 8658 -10331
rect 8716 -10365 8750 -10331
rect 8808 -10365 8842 -10331
rect 8900 -10365 8934 -10331
rect 8992 -10365 9026 -10331
rect 9084 -10365 9118 -10331
rect 9176 -10365 9210 -10331
rect 9268 -10365 9302 -10331
rect 9360 -10365 9394 -10331
rect 9452 -10365 9486 -10331
rect 9544 -10365 9578 -10331
rect 9636 -10365 9670 -10331
rect 9728 -10365 9762 -10331
rect 9820 -10365 9854 -10331
rect 9912 -10365 9946 -10331
rect 10004 -10365 10038 -10331
rect 10096 -10365 10130 -10331
rect 10188 -10365 10222 -10331
rect 10280 -10365 10314 -10331
rect 10372 -10365 10406 -10331
rect 10464 -10365 10498 -10331
rect 10556 -10365 10590 -10331
rect 10648 -10365 10682 -10331
rect 10740 -10365 10774 -10331
rect 10832 -10365 10866 -10331
rect 10924 -10365 10958 -10331
rect 11016 -10365 11050 -10331
rect 11108 -10365 11142 -10331
rect 11200 -10365 11234 -10331
rect 11292 -10365 11326 -10331
rect 11384 -10365 11418 -10331
rect 11476 -10365 11510 -10331
rect 11568 -10365 11602 -10331
rect 11660 -10365 11694 -10331
rect 11752 -10365 11786 -10331
rect 11844 -10365 11878 -10331
rect 11936 -10365 11970 -10331
rect 12028 -10365 12062 -10331
rect 12120 -10365 12154 -10331
rect 12212 -10365 12246 -10331
rect 12304 -10365 12338 -10331
rect 12396 -10365 12430 -10331
rect 12488 -10365 12522 -10331
rect 12580 -10365 12614 -10331
rect 12672 -10365 12706 -10331
rect 12764 -10365 12798 -10331
rect 12856 -10365 12890 -10331
rect 12948 -10365 12982 -10331
rect 13040 -10365 13074 -10331
rect 13132 -10365 13166 -10331
rect 13224 -10365 13258 -10331
rect 13316 -10365 13350 -10331
rect 13408 -10365 13442 -10331
rect 13500 -10365 13534 -10331
rect 13592 -10365 13626 -10331
rect 13684 -10365 13718 -10331
rect 13776 -10365 13810 -10331
rect 13868 -10365 13902 -10331
rect 13960 -10365 13994 -10331
rect 14052 -10365 14086 -10331
rect 14144 -10365 14178 -10331
rect 14236 -10365 14270 -10331
rect 14328 -10365 14362 -10331
rect 14420 -10365 14454 -10331
rect 14512 -10365 14546 -10331
rect 14604 -10365 14638 -10331
rect 14696 -10365 14730 -10331
rect 14788 -10365 14822 -10331
rect 14880 -10365 14914 -10331
rect 14972 -10365 15006 -10331
rect 15064 -10365 15098 -10331
rect 15156 -10365 15190 -10331
rect 15248 -10365 15282 -10331
rect 15340 -10365 15374 -10331
rect 15432 -10365 15466 -10331
rect 15524 -10365 15558 -10331
rect 15616 -10365 15650 -10331
rect 15708 -10365 15742 -10331
rect 15800 -10365 15834 -10331
rect 15892 -10365 15926 -10331
rect 15984 -10365 16018 -10331
rect 16076 -10365 16110 -10331
rect 16168 -10365 16202 -10331
rect 16260 -10365 16294 -10331
rect 16352 -10365 16386 -10331
rect 16444 -10365 16478 -10331
rect 16536 -10365 16570 -10331
rect 16628 -10365 16662 -10331
rect -1961 -10533 -1927 -10499
rect -1813 -10568 -1779 -10534
rect 429 -10637 463 -10603
rect 1072 -10597 1086 -10568
rect 1086 -10597 1106 -10568
rect 1072 -10602 1106 -10597
rect 3016 -10603 3050 -10569
rect 3630 -10597 3662 -10569
rect 3662 -10597 3664 -10569
rect 3630 -10603 3664 -10597
rect 5590 -10603 5624 -10569
rect 6204 -10597 6238 -10569
rect 6204 -10603 6238 -10597
rect 8164 -10603 8198 -10569
rect 8778 -10597 8780 -10569
rect 8780 -10597 8812 -10569
rect 8778 -10603 8812 -10597
rect 10738 -10604 10772 -10570
rect 11384 -10597 11390 -10568
rect 11390 -10597 11418 -10568
rect 11384 -10602 11418 -10597
rect -2968 -10909 -2934 -10875
rect -2876 -10909 -2842 -10875
rect -2784 -10909 -2750 -10875
rect -2692 -10909 -2658 -10875
rect -2600 -10909 -2566 -10875
rect -2508 -10909 -2474 -10875
rect -2416 -10909 -2382 -10875
rect -2324 -10909 -2290 -10875
rect -2232 -10909 -2198 -10875
rect -2140 -10909 -2106 -10875
rect -2048 -10909 -2014 -10875
rect -1956 -10909 -1922 -10875
rect -1864 -10909 -1830 -10875
rect -1772 -10909 -1738 -10875
rect -1680 -10909 -1646 -10875
rect -1588 -10909 -1554 -10875
rect -1496 -10909 -1462 -10875
rect -1404 -10909 -1370 -10875
rect -1312 -10909 -1278 -10875
rect -1220 -10909 -1186 -10875
rect -1128 -10909 -1094 -10875
rect -1036 -10909 -1002 -10875
rect -944 -10909 -910 -10875
rect -852 -10909 -818 -10875
rect -760 -10909 -726 -10875
rect -668 -10909 -634 -10875
rect -576 -10909 -542 -10875
rect -484 -10909 -450 -10875
rect -392 -10909 -358 -10875
rect -300 -10909 -266 -10875
rect -208 -10909 -174 -10875
rect -116 -10909 -82 -10875
rect -24 -10909 10 -10875
rect 68 -10909 102 -10875
rect 160 -10909 194 -10875
rect 252 -10909 286 -10875
rect 344 -10909 378 -10875
rect 436 -10909 470 -10875
rect 528 -10909 562 -10875
rect 620 -10909 654 -10875
rect 712 -10909 746 -10875
rect 804 -10909 838 -10875
rect 896 -10909 930 -10875
rect 988 -10909 1022 -10875
rect 1080 -10909 1114 -10875
rect 1172 -10909 1206 -10875
rect 1264 -10909 1298 -10875
rect 1356 -10909 1390 -10875
rect 1448 -10909 1482 -10875
rect 1540 -10909 1574 -10875
rect 1632 -10909 1666 -10875
rect 1724 -10909 1758 -10875
rect 1816 -10909 1850 -10875
rect 1908 -10909 1942 -10875
rect 2000 -10909 2034 -10875
rect 2092 -10909 2126 -10875
rect 2184 -10909 2218 -10875
rect 2276 -10909 2310 -10875
rect 2368 -10909 2402 -10875
rect 2460 -10909 2494 -10875
rect 2552 -10909 2586 -10875
rect 2644 -10909 2678 -10875
rect 2736 -10909 2770 -10875
rect 2828 -10909 2862 -10875
rect 2920 -10909 2954 -10875
rect 3012 -10909 3046 -10875
rect 3104 -10909 3138 -10875
rect 3196 -10909 3230 -10875
rect 3288 -10909 3322 -10875
rect 3380 -10909 3414 -10875
rect 3472 -10909 3506 -10875
rect 3564 -10909 3598 -10875
rect 3656 -10909 3690 -10875
rect 3748 -10909 3782 -10875
rect 3840 -10909 3874 -10875
rect 3932 -10909 3966 -10875
rect 4024 -10909 4058 -10875
rect 4116 -10909 4150 -10875
rect 4208 -10909 4242 -10875
rect 4300 -10909 4334 -10875
rect 4392 -10909 4426 -10875
rect 4484 -10909 4518 -10875
rect 4576 -10909 4610 -10875
rect 4668 -10909 4702 -10875
rect 4760 -10909 4794 -10875
rect 4852 -10909 4886 -10875
rect 4944 -10909 4978 -10875
rect 5036 -10909 5070 -10875
rect 5128 -10909 5162 -10875
rect 5220 -10909 5254 -10875
rect 5312 -10909 5346 -10875
rect 5404 -10909 5438 -10875
rect 5496 -10909 5530 -10875
rect 5588 -10909 5622 -10875
rect 5680 -10909 5714 -10875
rect 5772 -10909 5806 -10875
rect 5864 -10909 5898 -10875
rect 5956 -10909 5990 -10875
rect 6048 -10909 6082 -10875
rect 6140 -10909 6174 -10875
rect 6232 -10909 6266 -10875
rect 6324 -10909 6358 -10875
rect 6416 -10909 6450 -10875
rect 6508 -10909 6542 -10875
rect 6600 -10909 6634 -10875
rect 6692 -10909 6726 -10875
rect 6784 -10909 6818 -10875
rect 6876 -10909 6910 -10875
rect 6968 -10909 7002 -10875
rect 7060 -10909 7094 -10875
rect 7152 -10909 7186 -10875
rect 7244 -10909 7278 -10875
rect 7336 -10909 7370 -10875
rect 7428 -10909 7462 -10875
rect 7520 -10909 7554 -10875
rect 7612 -10909 7646 -10875
rect 7704 -10909 7738 -10875
rect 7796 -10909 7830 -10875
rect 7888 -10909 7922 -10875
rect 7980 -10909 8014 -10875
rect 8072 -10909 8106 -10875
rect 8164 -10909 8198 -10875
rect 8256 -10909 8290 -10875
rect 8348 -10909 8382 -10875
rect 8440 -10909 8474 -10875
rect 8532 -10909 8566 -10875
rect 8624 -10909 8658 -10875
rect 8716 -10909 8750 -10875
rect 8808 -10909 8842 -10875
rect 8900 -10909 8934 -10875
rect 8992 -10909 9026 -10875
rect 9084 -10909 9118 -10875
rect 9176 -10909 9210 -10875
rect 9268 -10909 9302 -10875
rect 9360 -10909 9394 -10875
rect 9452 -10909 9486 -10875
rect 9544 -10909 9578 -10875
rect 9636 -10909 9670 -10875
rect 9728 -10909 9762 -10875
rect 9820 -10909 9854 -10875
rect 9912 -10909 9946 -10875
rect 10004 -10909 10038 -10875
rect 10096 -10909 10130 -10875
rect 10188 -10909 10222 -10875
rect 10280 -10909 10314 -10875
rect 10372 -10909 10406 -10875
rect 10464 -10909 10498 -10875
rect 10556 -10909 10590 -10875
rect 10648 -10909 10682 -10875
rect 10740 -10909 10774 -10875
rect 10832 -10909 10866 -10875
rect 10924 -10909 10958 -10875
rect 11016 -10909 11050 -10875
rect 11108 -10909 11142 -10875
rect 11200 -10909 11234 -10875
rect 11292 -10909 11326 -10875
rect 11384 -10909 11418 -10875
rect 11476 -10909 11510 -10875
rect 11568 -10909 11602 -10875
rect 11660 -10909 11694 -10875
rect 11752 -10909 11786 -10875
rect 11844 -10909 11878 -10875
rect 11936 -10909 11970 -10875
rect 12028 -10909 12062 -10875
rect 12120 -10909 12154 -10875
rect 12212 -10909 12246 -10875
rect 12304 -10909 12338 -10875
rect 12396 -10909 12430 -10875
rect 12488 -10909 12522 -10875
rect 12580 -10909 12614 -10875
rect 12672 -10909 12706 -10875
rect 12764 -10909 12798 -10875
rect 12856 -10909 12890 -10875
rect 12948 -10909 12982 -10875
rect 13040 -10909 13074 -10875
rect 13132 -10909 13166 -10875
rect 13224 -10909 13258 -10875
rect 13316 -10909 13350 -10875
rect 13408 -10909 13442 -10875
rect 13500 -10909 13534 -10875
rect 13592 -10909 13626 -10875
rect 13684 -10909 13718 -10875
rect 13776 -10909 13810 -10875
rect 13868 -10909 13902 -10875
rect 13960 -10909 13994 -10875
rect 14052 -10909 14086 -10875
rect 14144 -10909 14178 -10875
rect 14236 -10909 14270 -10875
rect 14328 -10909 14362 -10875
rect 14420 -10909 14454 -10875
rect 14512 -10909 14546 -10875
rect 14604 -10909 14638 -10875
rect 14696 -10909 14730 -10875
rect 14788 -10909 14822 -10875
rect 14880 -10909 14914 -10875
rect 14972 -10909 15006 -10875
rect 15064 -10909 15098 -10875
rect 15156 -10909 15190 -10875
rect 15248 -10909 15282 -10875
rect 15340 -10909 15374 -10875
rect 15432 -10909 15466 -10875
rect 15524 -10909 15558 -10875
rect 15616 -10909 15650 -10875
rect 15708 -10909 15742 -10875
rect 15800 -10909 15834 -10875
rect 15892 -10909 15926 -10875
rect 15984 -10909 16018 -10875
rect 16076 -10909 16110 -10875
rect 16168 -10909 16202 -10875
rect 16260 -10909 16294 -10875
rect 16352 -10909 16386 -10875
rect 16444 -10909 16478 -10875
rect 16536 -10909 16570 -10875
rect 16628 -10909 16662 -10875
rect 432 -11181 466 -11147
rect 1070 -11187 1104 -11184
rect 1070 -11218 1086 -11187
rect 1086 -11218 1104 -11187
rect 3016 -11215 3050 -11181
rect 3630 -11187 3664 -11181
rect 3630 -11215 3662 -11187
rect 3662 -11215 3664 -11187
rect 5590 -11215 5624 -11181
rect 6204 -11187 6238 -11181
rect 6204 -11215 6238 -11187
rect 8164 -11215 8198 -11181
rect 8778 -11187 8812 -11181
rect 8778 -11215 8780 -11187
rect 8780 -11215 8812 -11187
rect 10735 -11218 10769 -11184
rect 11383 -11187 11417 -11183
rect 11383 -11217 11390 -11187
rect 11390 -11217 11417 -11187
rect -2968 -11453 -2934 -11419
rect -2876 -11453 -2842 -11419
rect -2784 -11453 -2750 -11419
rect -2692 -11453 -2658 -11419
rect -2600 -11453 -2566 -11419
rect -2508 -11453 -2474 -11419
rect -2416 -11453 -2382 -11419
rect -2324 -11453 -2290 -11419
rect -2232 -11453 -2198 -11419
rect -2140 -11453 -2106 -11419
rect -2048 -11453 -2014 -11419
rect -1956 -11453 -1922 -11419
rect -1864 -11453 -1830 -11419
rect -1772 -11453 -1738 -11419
rect -1680 -11453 -1646 -11419
rect -1588 -11453 -1554 -11419
rect -1496 -11453 -1462 -11419
rect -1404 -11453 -1370 -11419
rect -1312 -11453 -1278 -11419
rect -1220 -11453 -1186 -11419
rect -1128 -11453 -1094 -11419
rect -1036 -11453 -1002 -11419
rect -944 -11453 -910 -11419
rect -852 -11453 -818 -11419
rect -760 -11453 -726 -11419
rect -668 -11453 -634 -11419
rect -576 -11453 -542 -11419
rect -484 -11453 -450 -11419
rect -392 -11453 -358 -11419
rect -300 -11453 -266 -11419
rect -208 -11453 -174 -11419
rect -116 -11453 -82 -11419
rect -24 -11453 10 -11419
rect 68 -11453 102 -11419
rect 160 -11453 194 -11419
rect 252 -11453 286 -11419
rect 344 -11453 378 -11419
rect 436 -11453 470 -11419
rect 528 -11453 562 -11419
rect 620 -11453 654 -11419
rect 712 -11453 746 -11419
rect 804 -11453 838 -11419
rect 896 -11453 930 -11419
rect 988 -11453 1022 -11419
rect 1080 -11453 1114 -11419
rect 1172 -11453 1206 -11419
rect 1264 -11453 1298 -11419
rect 1356 -11453 1390 -11419
rect 1448 -11453 1482 -11419
rect 1540 -11453 1574 -11419
rect 1632 -11453 1666 -11419
rect 1724 -11453 1758 -11419
rect 1816 -11453 1850 -11419
rect 1908 -11453 1942 -11419
rect 2000 -11453 2034 -11419
rect 2092 -11453 2126 -11419
rect 2184 -11453 2218 -11419
rect 2276 -11453 2310 -11419
rect 2368 -11453 2402 -11419
rect 2460 -11453 2494 -11419
rect 2552 -11453 2586 -11419
rect 2644 -11453 2678 -11419
rect 2736 -11453 2770 -11419
rect 2828 -11453 2862 -11419
rect 2920 -11453 2954 -11419
rect 3012 -11453 3046 -11419
rect 3104 -11453 3138 -11419
rect 3196 -11453 3230 -11419
rect 3288 -11453 3322 -11419
rect 3380 -11453 3414 -11419
rect 3472 -11453 3506 -11419
rect 3564 -11453 3598 -11419
rect 3656 -11453 3690 -11419
rect 3748 -11453 3782 -11419
rect 3840 -11453 3874 -11419
rect 3932 -11453 3966 -11419
rect 4024 -11453 4058 -11419
rect 4116 -11453 4150 -11419
rect 4208 -11453 4242 -11419
rect 4300 -11453 4334 -11419
rect 4392 -11453 4426 -11419
rect 4484 -11453 4518 -11419
rect 4576 -11453 4610 -11419
rect 4668 -11453 4702 -11419
rect 4760 -11453 4794 -11419
rect 4852 -11453 4886 -11419
rect 4944 -11453 4978 -11419
rect 5036 -11453 5070 -11419
rect 5128 -11453 5162 -11419
rect 5220 -11453 5254 -11419
rect 5312 -11453 5346 -11419
rect 5404 -11453 5438 -11419
rect 5496 -11453 5530 -11419
rect 5588 -11453 5622 -11419
rect 5680 -11453 5714 -11419
rect 5772 -11453 5806 -11419
rect 5864 -11453 5898 -11419
rect 5956 -11453 5990 -11419
rect 6048 -11453 6082 -11419
rect 6140 -11453 6174 -11419
rect 6232 -11453 6266 -11419
rect 6324 -11453 6358 -11419
rect 6416 -11453 6450 -11419
rect 6508 -11453 6542 -11419
rect 6600 -11453 6634 -11419
rect 6692 -11453 6726 -11419
rect 6784 -11453 6818 -11419
rect 6876 -11453 6910 -11419
rect 6968 -11453 7002 -11419
rect 7060 -11453 7094 -11419
rect 7152 -11453 7186 -11419
rect 7244 -11453 7278 -11419
rect 7336 -11453 7370 -11419
rect 7428 -11453 7462 -11419
rect 7520 -11453 7554 -11419
rect 7612 -11453 7646 -11419
rect 7704 -11453 7738 -11419
rect 7796 -11453 7830 -11419
rect 7888 -11453 7922 -11419
rect 7980 -11453 8014 -11419
rect 8072 -11453 8106 -11419
rect 8164 -11453 8198 -11419
rect 8256 -11453 8290 -11419
rect 8348 -11453 8382 -11419
rect 8440 -11453 8474 -11419
rect 8532 -11453 8566 -11419
rect 8624 -11453 8658 -11419
rect 8716 -11453 8750 -11419
rect 8808 -11453 8842 -11419
rect 8900 -11453 8934 -11419
rect 8992 -11453 9026 -11419
rect 9084 -11453 9118 -11419
rect 9176 -11453 9210 -11419
rect 9268 -11453 9302 -11419
rect 9360 -11453 9394 -11419
rect 9452 -11453 9486 -11419
rect 9544 -11453 9578 -11419
rect 9636 -11453 9670 -11419
rect 9728 -11453 9762 -11419
rect 9820 -11453 9854 -11419
rect 9912 -11453 9946 -11419
rect 10004 -11453 10038 -11419
rect 10096 -11453 10130 -11419
rect 10188 -11453 10222 -11419
rect 10280 -11453 10314 -11419
rect 10372 -11453 10406 -11419
rect 10464 -11453 10498 -11419
rect 10556 -11453 10590 -11419
rect 10648 -11453 10682 -11419
rect 10740 -11453 10774 -11419
rect 10832 -11453 10866 -11419
rect 10924 -11453 10958 -11419
rect 11016 -11453 11050 -11419
rect 11108 -11453 11142 -11419
rect 11200 -11453 11234 -11419
rect 11292 -11453 11326 -11419
rect 11384 -11453 11418 -11419
rect 11476 -11453 11510 -11419
rect 11568 -11453 11602 -11419
rect 11660 -11453 11694 -11419
rect 11752 -11453 11786 -11419
rect 11844 -11453 11878 -11419
rect 11936 -11453 11970 -11419
rect 12028 -11453 12062 -11419
rect 12120 -11453 12154 -11419
rect 12212 -11453 12246 -11419
rect 12304 -11453 12338 -11419
rect 12396 -11453 12430 -11419
rect 12488 -11453 12522 -11419
rect 12580 -11453 12614 -11419
rect 12672 -11453 12706 -11419
rect 12764 -11453 12798 -11419
rect 12856 -11453 12890 -11419
rect 12948 -11453 12982 -11419
rect 13040 -11453 13074 -11419
rect 13132 -11453 13166 -11419
rect 13224 -11453 13258 -11419
rect 13316 -11453 13350 -11419
rect 13408 -11453 13442 -11419
rect 13500 -11453 13534 -11419
rect 13592 -11453 13626 -11419
rect 13684 -11453 13718 -11419
rect 13776 -11453 13810 -11419
rect 13868 -11453 13902 -11419
rect 13960 -11453 13994 -11419
rect 14052 -11453 14086 -11419
rect 14144 -11453 14178 -11419
rect 14236 -11453 14270 -11419
rect 14328 -11453 14362 -11419
rect 14420 -11453 14454 -11419
rect 14512 -11453 14546 -11419
rect 14604 -11453 14638 -11419
rect 14696 -11453 14730 -11419
rect 14788 -11453 14822 -11419
rect 14880 -11453 14914 -11419
rect 14972 -11453 15006 -11419
rect 15064 -11453 15098 -11419
rect 15156 -11453 15190 -11419
rect 15248 -11453 15282 -11419
rect 15340 -11453 15374 -11419
rect 15432 -11453 15466 -11419
rect 15524 -11453 15558 -11419
rect 15616 -11453 15650 -11419
rect 15708 -11453 15742 -11419
rect 15800 -11453 15834 -11419
rect 15892 -11453 15926 -11419
rect 15984 -11453 16018 -11419
rect 16076 -11453 16110 -11419
rect 16168 -11453 16202 -11419
rect 16260 -11453 16294 -11419
rect 16352 -11453 16386 -11419
rect 16444 -11453 16478 -11419
rect 16536 -11453 16570 -11419
rect 16628 -11453 16662 -11419
rect 436 -11685 464 -11656
rect 464 -11685 470 -11656
rect 436 -11690 470 -11685
rect 1081 -11690 1115 -11656
rect 3041 -11685 3074 -11656
rect 3074 -11685 3075 -11656
rect 3041 -11690 3075 -11685
rect 3655 -11690 3689 -11656
rect 5615 -11685 5616 -11656
rect 5616 -11685 5649 -11656
rect 5615 -11690 5649 -11685
rect 6229 -11690 6263 -11656
rect 8189 -11685 8192 -11656
rect 8192 -11685 8223 -11656
rect 8189 -11690 8223 -11685
rect 8806 -11690 8840 -11656
rect 10763 -11685 10768 -11656
rect 10768 -11685 10797 -11656
rect 10763 -11690 10797 -11685
rect 11386 -11727 11420 -11693
rect 12480 -11615 12514 -11581
rect 13042 -11625 13076 -11591
rect 12480 -11687 12514 -11653
rect 12568 -11685 12574 -11655
rect 12574 -11685 12602 -11655
rect 12659 -11685 12676 -11655
rect 12676 -11685 12693 -11655
rect 12765 -11685 12778 -11655
rect 12778 -11685 12799 -11655
rect 12858 -11685 12880 -11657
rect 12880 -11685 12892 -11657
rect 12942 -11685 12948 -11657
rect 12948 -11685 12976 -11657
rect 12568 -11689 12602 -11685
rect 12659 -11689 12693 -11685
rect 12765 -11689 12799 -11685
rect 12858 -11691 12892 -11685
rect 12942 -11691 12976 -11685
rect 12480 -11761 12514 -11727
rect 13039 -11702 13073 -11668
rect 13685 -11651 13719 -11624
rect 13685 -11658 13692 -11651
rect 13692 -11658 13719 -11651
rect 15248 -11646 15282 -11612
rect 15341 -11646 15375 -11612
rect 15248 -11742 15282 -11708
rect 15340 -11742 15374 -11708
rect -2968 -11997 -2934 -11963
rect -2876 -11997 -2842 -11963
rect -2784 -11997 -2750 -11963
rect -2692 -11997 -2658 -11963
rect -2600 -11997 -2566 -11963
rect -2508 -11997 -2474 -11963
rect -2416 -11997 -2382 -11963
rect -2324 -11997 -2290 -11963
rect -2232 -11997 -2198 -11963
rect -2140 -11997 -2106 -11963
rect -2048 -11997 -2014 -11963
rect -1956 -11997 -1922 -11963
rect -1864 -11997 -1830 -11963
rect -1772 -11997 -1738 -11963
rect -1680 -11997 -1646 -11963
rect -1588 -11997 -1554 -11963
rect -1496 -11997 -1462 -11963
rect -1404 -11997 -1370 -11963
rect -1312 -11997 -1278 -11963
rect -1220 -11997 -1186 -11963
rect -1128 -11997 -1094 -11963
rect -1036 -11997 -1002 -11963
rect -944 -11997 -910 -11963
rect -852 -11997 -818 -11963
rect -760 -11997 -726 -11963
rect -668 -11997 -634 -11963
rect -576 -11997 -542 -11963
rect -484 -11997 -450 -11963
rect -392 -11997 -358 -11963
rect -300 -11997 -266 -11963
rect -208 -11997 -174 -11963
rect -116 -11997 -82 -11963
rect -24 -11997 10 -11963
rect 68 -11997 102 -11963
rect 160 -11997 194 -11963
rect 252 -11997 286 -11963
rect 344 -11997 378 -11963
rect 436 -11997 470 -11963
rect 528 -11997 562 -11963
rect 620 -11997 654 -11963
rect 712 -11997 746 -11963
rect 804 -11997 838 -11963
rect 896 -11997 930 -11963
rect 988 -11997 1022 -11963
rect 1080 -11997 1114 -11963
rect 1172 -11997 1206 -11963
rect 1264 -11997 1298 -11963
rect 1356 -11997 1390 -11963
rect 1448 -11997 1482 -11963
rect 1540 -11997 1574 -11963
rect 1632 -11997 1666 -11963
rect 1724 -11997 1758 -11963
rect 1816 -11997 1850 -11963
rect 1908 -11997 1942 -11963
rect 2000 -11997 2034 -11963
rect 2092 -11997 2126 -11963
rect 2184 -11997 2218 -11963
rect 2276 -11997 2310 -11963
rect 2368 -11997 2402 -11963
rect 2460 -11997 2494 -11963
rect 2552 -11997 2586 -11963
rect 2644 -11997 2678 -11963
rect 2736 -11997 2770 -11963
rect 2828 -11997 2862 -11963
rect 2920 -11997 2954 -11963
rect 3012 -11997 3046 -11963
rect 3104 -11997 3138 -11963
rect 3196 -11997 3230 -11963
rect 3288 -11997 3322 -11963
rect 3380 -11997 3414 -11963
rect 3472 -11997 3506 -11963
rect 3564 -11997 3598 -11963
rect 3656 -11997 3690 -11963
rect 3748 -11997 3782 -11963
rect 3840 -11997 3874 -11963
rect 3932 -11997 3966 -11963
rect 4024 -11997 4058 -11963
rect 4116 -11997 4150 -11963
rect 4208 -11997 4242 -11963
rect 4300 -11997 4334 -11963
rect 4392 -11997 4426 -11963
rect 4484 -11997 4518 -11963
rect 4576 -11997 4610 -11963
rect 4668 -11997 4702 -11963
rect 4760 -11997 4794 -11963
rect 4852 -11997 4886 -11963
rect 4944 -11997 4978 -11963
rect 5036 -11997 5070 -11963
rect 5128 -11997 5162 -11963
rect 5220 -11997 5254 -11963
rect 5312 -11997 5346 -11963
rect 5404 -11997 5438 -11963
rect 5496 -11997 5530 -11963
rect 5588 -11997 5622 -11963
rect 5680 -11997 5714 -11963
rect 5772 -11997 5806 -11963
rect 5864 -11997 5898 -11963
rect 5956 -11997 5990 -11963
rect 6048 -11997 6082 -11963
rect 6140 -11997 6174 -11963
rect 6232 -11997 6266 -11963
rect 6324 -11997 6358 -11963
rect 6416 -11997 6450 -11963
rect 6508 -11997 6542 -11963
rect 6600 -11997 6634 -11963
rect 6692 -11997 6726 -11963
rect 6784 -11997 6818 -11963
rect 6876 -11997 6910 -11963
rect 6968 -11997 7002 -11963
rect 7060 -11997 7094 -11963
rect 7152 -11997 7186 -11963
rect 7244 -11997 7278 -11963
rect 7336 -11997 7370 -11963
rect 7428 -11997 7462 -11963
rect 7520 -11997 7554 -11963
rect 7612 -11997 7646 -11963
rect 7704 -11997 7738 -11963
rect 7796 -11997 7830 -11963
rect 7888 -11997 7922 -11963
rect 7980 -11997 8014 -11963
rect 8072 -11997 8106 -11963
rect 8164 -11997 8198 -11963
rect 8256 -11997 8290 -11963
rect 8348 -11997 8382 -11963
rect 8440 -11997 8474 -11963
rect 8532 -11997 8566 -11963
rect 8624 -11997 8658 -11963
rect 8716 -11997 8750 -11963
rect 8808 -11997 8842 -11963
rect 8900 -11997 8934 -11963
rect 8992 -11997 9026 -11963
rect 9084 -11997 9118 -11963
rect 9176 -11997 9210 -11963
rect 9268 -11997 9302 -11963
rect 9360 -11997 9394 -11963
rect 9452 -11997 9486 -11963
rect 9544 -11997 9578 -11963
rect 9636 -11997 9670 -11963
rect 9728 -11997 9762 -11963
rect 9820 -11997 9854 -11963
rect 9912 -11997 9946 -11963
rect 10004 -11997 10038 -11963
rect 10096 -11997 10130 -11963
rect 10188 -11997 10222 -11963
rect 10280 -11997 10314 -11963
rect 10372 -11997 10406 -11963
rect 10464 -11997 10498 -11963
rect 10556 -11997 10590 -11963
rect 10648 -11997 10682 -11963
rect 10740 -11997 10774 -11963
rect 10832 -11997 10866 -11963
rect 10924 -11997 10958 -11963
rect 11016 -11997 11050 -11963
rect 11108 -11997 11142 -11963
rect 11200 -11997 11234 -11963
rect 11292 -11997 11326 -11963
rect 11384 -11997 11418 -11963
rect 11476 -11997 11510 -11963
rect 11568 -11997 11602 -11963
rect 11660 -11997 11694 -11963
rect 11752 -11997 11786 -11963
rect 11844 -11997 11878 -11963
rect 11936 -11997 11970 -11963
rect 12028 -11997 12062 -11963
rect 12120 -11997 12154 -11963
rect 12212 -11997 12246 -11963
rect 12304 -11997 12338 -11963
rect 12396 -11997 12430 -11963
rect 12488 -11997 12522 -11963
rect 12580 -11997 12614 -11963
rect 12672 -11997 12706 -11963
rect 12764 -11997 12798 -11963
rect 12856 -11997 12890 -11963
rect 12948 -11997 12982 -11963
rect 13040 -11997 13074 -11963
rect 13132 -11997 13166 -11963
rect 13224 -11997 13258 -11963
rect 13316 -11997 13350 -11963
rect 13408 -11997 13442 -11963
rect 13500 -11997 13534 -11963
rect 13592 -11997 13626 -11963
rect 13684 -11997 13718 -11963
rect 13776 -11997 13810 -11963
rect 13868 -11997 13902 -11963
rect 13960 -11997 13994 -11963
rect 14052 -11997 14086 -11963
rect 14144 -11997 14178 -11963
rect 14236 -11997 14270 -11963
rect 14328 -11997 14362 -11963
rect 14420 -11997 14454 -11963
rect 14512 -11997 14546 -11963
rect 14604 -11997 14638 -11963
rect 14696 -11997 14730 -11963
rect 14788 -11997 14822 -11963
rect 14880 -11997 14914 -11963
rect 14972 -11997 15006 -11963
rect 15064 -11997 15098 -11963
rect 15156 -11997 15190 -11963
rect 15248 -11997 15282 -11963
rect 15340 -11997 15374 -11963
rect 15432 -11997 15466 -11963
rect 15524 -11997 15558 -11963
rect 15616 -11997 15650 -11963
rect 15708 -11997 15742 -11963
rect 15800 -11997 15834 -11963
rect 15892 -11997 15926 -11963
rect 15984 -11997 16018 -11963
rect 16076 -11997 16110 -11963
rect 16168 -11997 16202 -11963
rect 16260 -11997 16294 -11963
rect 16352 -11997 16386 -11963
rect 16444 -11997 16478 -11963
rect 16536 -11997 16570 -11963
rect 16628 -11997 16662 -11963
rect -855 -12269 -821 -12235
rect -210 -12275 -176 -12272
rect -210 -12306 -202 -12275
rect -202 -12306 -176 -12275
rect 433 -12269 467 -12235
rect 1054 -12275 1088 -12268
rect 1054 -12302 1086 -12275
rect 1086 -12302 1088 -12275
rect 3014 -12302 3048 -12268
rect 3628 -12275 3662 -12268
rect 3628 -12302 3662 -12275
rect 5588 -12302 5622 -12268
rect 6202 -12275 6236 -12268
rect 6202 -12302 6204 -12275
rect 6204 -12302 6236 -12275
rect 8162 -12302 8196 -12268
rect 8776 -12275 8810 -12268
rect 8776 -12302 8780 -12275
rect 8780 -12302 8810 -12275
rect 10736 -12302 10770 -12268
rect 11384 -12275 11418 -12273
rect 11384 -12307 11390 -12275
rect 11390 -12307 11418 -12275
rect 15248 -12256 15282 -12222
rect 15341 -12256 15375 -12222
rect 13685 -12309 13692 -12302
rect 13692 -12309 13719 -12302
rect 13685 -12336 13719 -12309
rect 15248 -12352 15282 -12318
rect 15340 -12351 15374 -12317
rect -2968 -12541 -2934 -12507
rect -2876 -12541 -2842 -12507
rect -2784 -12541 -2750 -12507
rect -2692 -12541 -2658 -12507
rect -2600 -12541 -2566 -12507
rect -2508 -12541 -2474 -12507
rect -2416 -12541 -2382 -12507
rect -2324 -12541 -2290 -12507
rect -2232 -12541 -2198 -12507
rect -2140 -12541 -2106 -12507
rect -2048 -12541 -2014 -12507
rect -1956 -12541 -1922 -12507
rect -1864 -12541 -1830 -12507
rect -1772 -12541 -1738 -12507
rect -1680 -12541 -1646 -12507
rect -1588 -12541 -1554 -12507
rect -1496 -12541 -1462 -12507
rect -1404 -12541 -1370 -12507
rect -1312 -12541 -1278 -12507
rect -1220 -12541 -1186 -12507
rect -1128 -12541 -1094 -12507
rect -1036 -12541 -1002 -12507
rect -944 -12541 -910 -12507
rect -852 -12541 -818 -12507
rect -760 -12541 -726 -12507
rect -668 -12541 -634 -12507
rect -576 -12541 -542 -12507
rect -484 -12541 -450 -12507
rect -392 -12541 -358 -12507
rect -300 -12541 -266 -12507
rect -208 -12541 -174 -12507
rect -116 -12541 -82 -12507
rect -24 -12541 10 -12507
rect 68 -12541 102 -12507
rect 160 -12541 194 -12507
rect 252 -12541 286 -12507
rect 344 -12541 378 -12507
rect 436 -12541 470 -12507
rect 528 -12541 562 -12507
rect 620 -12541 654 -12507
rect 712 -12541 746 -12507
rect 804 -12541 838 -12507
rect 896 -12541 930 -12507
rect 988 -12541 1022 -12507
rect 1080 -12541 1114 -12507
rect 1172 -12541 1206 -12507
rect 1264 -12541 1298 -12507
rect 1356 -12541 1390 -12507
rect 1448 -12541 1482 -12507
rect 1540 -12541 1574 -12507
rect 1632 -12541 1666 -12507
rect 1724 -12541 1758 -12507
rect 1816 -12541 1850 -12507
rect 1908 -12541 1942 -12507
rect 2000 -12541 2034 -12507
rect 2092 -12541 2126 -12507
rect 2184 -12541 2218 -12507
rect 2276 -12541 2310 -12507
rect 2368 -12541 2402 -12507
rect 2460 -12541 2494 -12507
rect 2552 -12541 2586 -12507
rect 2644 -12541 2678 -12507
rect 2736 -12541 2770 -12507
rect 2828 -12541 2862 -12507
rect 2920 -12541 2954 -12507
rect 3012 -12541 3046 -12507
rect 3104 -12541 3138 -12507
rect 3196 -12541 3230 -12507
rect 3288 -12541 3322 -12507
rect 3380 -12541 3414 -12507
rect 3472 -12541 3506 -12507
rect 3564 -12541 3598 -12507
rect 3656 -12541 3690 -12507
rect 3748 -12541 3782 -12507
rect 3840 -12541 3874 -12507
rect 3932 -12541 3966 -12507
rect 4024 -12541 4058 -12507
rect 4116 -12541 4150 -12507
rect 4208 -12541 4242 -12507
rect 4300 -12541 4334 -12507
rect 4392 -12541 4426 -12507
rect 4484 -12541 4518 -12507
rect 4576 -12541 4610 -12507
rect 4668 -12541 4702 -12507
rect 4760 -12541 4794 -12507
rect 4852 -12541 4886 -12507
rect 4944 -12541 4978 -12507
rect 5036 -12541 5070 -12507
rect 5128 -12541 5162 -12507
rect 5220 -12541 5254 -12507
rect 5312 -12541 5346 -12507
rect 5404 -12541 5438 -12507
rect 5496 -12541 5530 -12507
rect 5588 -12541 5622 -12507
rect 5680 -12541 5714 -12507
rect 5772 -12541 5806 -12507
rect 5864 -12541 5898 -12507
rect 5956 -12541 5990 -12507
rect 6048 -12541 6082 -12507
rect 6140 -12541 6174 -12507
rect 6232 -12541 6266 -12507
rect 6324 -12541 6358 -12507
rect 6416 -12541 6450 -12507
rect 6508 -12541 6542 -12507
rect 6600 -12541 6634 -12507
rect 6692 -12541 6726 -12507
rect 6784 -12541 6818 -12507
rect 6876 -12541 6910 -12507
rect 6968 -12541 7002 -12507
rect 7060 -12541 7094 -12507
rect 7152 -12541 7186 -12507
rect 7244 -12541 7278 -12507
rect 7336 -12541 7370 -12507
rect 7428 -12541 7462 -12507
rect 7520 -12541 7554 -12507
rect 7612 -12541 7646 -12507
rect 7704 -12541 7738 -12507
rect 7796 -12541 7830 -12507
rect 7888 -12541 7922 -12507
rect 7980 -12541 8014 -12507
rect 8072 -12541 8106 -12507
rect 8164 -12541 8198 -12507
rect 8256 -12541 8290 -12507
rect 8348 -12541 8382 -12507
rect 8440 -12541 8474 -12507
rect 8532 -12541 8566 -12507
rect 8624 -12541 8658 -12507
rect 8716 -12541 8750 -12507
rect 8808 -12541 8842 -12507
rect 8900 -12541 8934 -12507
rect 8992 -12541 9026 -12507
rect 9084 -12541 9118 -12507
rect 9176 -12541 9210 -12507
rect 9268 -12541 9302 -12507
rect 9360 -12541 9394 -12507
rect 9452 -12541 9486 -12507
rect 9544 -12541 9578 -12507
rect 9636 -12541 9670 -12507
rect 9728 -12541 9762 -12507
rect 9820 -12541 9854 -12507
rect 9912 -12541 9946 -12507
rect 10004 -12541 10038 -12507
rect 10096 -12541 10130 -12507
rect 10188 -12541 10222 -12507
rect 10280 -12541 10314 -12507
rect 10372 -12541 10406 -12507
rect 10464 -12541 10498 -12507
rect 10556 -12541 10590 -12507
rect 10648 -12541 10682 -12507
rect 10740 -12541 10774 -12507
rect 10832 -12541 10866 -12507
rect 10924 -12541 10958 -12507
rect 11016 -12541 11050 -12507
rect 11108 -12541 11142 -12507
rect 11200 -12541 11234 -12507
rect 11292 -12541 11326 -12507
rect 11384 -12541 11418 -12507
rect 11476 -12541 11510 -12507
rect 11568 -12541 11602 -12507
rect 11660 -12541 11694 -12507
rect 11752 -12541 11786 -12507
rect 11844 -12541 11878 -12507
rect 11936 -12541 11970 -12507
rect 12028 -12541 12062 -12507
rect 12120 -12541 12154 -12507
rect 12212 -12541 12246 -12507
rect 12304 -12541 12338 -12507
rect 12396 -12541 12430 -12507
rect 12488 -12541 12522 -12507
rect 12580 -12541 12614 -12507
rect 12672 -12541 12706 -12507
rect 12764 -12541 12798 -12507
rect 12856 -12541 12890 -12507
rect 12948 -12541 12982 -12507
rect 13040 -12541 13074 -12507
rect 13132 -12541 13166 -12507
rect 13224 -12541 13258 -12507
rect 13316 -12541 13350 -12507
rect 13408 -12541 13442 -12507
rect 13500 -12541 13534 -12507
rect 13592 -12541 13626 -12507
rect 13684 -12541 13718 -12507
rect 13776 -12541 13810 -12507
rect 13868 -12541 13902 -12507
rect 13960 -12541 13994 -12507
rect 14052 -12541 14086 -12507
rect 14144 -12541 14178 -12507
rect 14236 -12541 14270 -12507
rect 14328 -12541 14362 -12507
rect 14420 -12541 14454 -12507
rect 14512 -12541 14546 -12507
rect 14604 -12541 14638 -12507
rect 14696 -12541 14730 -12507
rect 14788 -12541 14822 -12507
rect 14880 -12541 14914 -12507
rect 14972 -12541 15006 -12507
rect 15064 -12541 15098 -12507
rect 15156 -12541 15190 -12507
rect 15248 -12541 15282 -12507
rect 15340 -12541 15374 -12507
rect 15432 -12541 15466 -12507
rect 15524 -12541 15558 -12507
rect 15616 -12541 15650 -12507
rect 15708 -12541 15742 -12507
rect 15800 -12541 15834 -12507
rect 15892 -12541 15926 -12507
rect 15984 -12541 16018 -12507
rect 16076 -12541 16110 -12507
rect 16168 -12541 16202 -12507
rect 16260 -12541 16294 -12507
rect 16352 -12541 16386 -12507
rect 16444 -12541 16478 -12507
rect 16536 -12541 16570 -12507
rect 16628 -12541 16662 -12507
rect 436 -12773 464 -12744
rect 464 -12773 470 -12744
rect 436 -12778 470 -12773
rect 1082 -12779 1116 -12745
rect 3042 -12773 3074 -12745
rect 3074 -12773 3076 -12745
rect 3042 -12779 3076 -12773
rect 3656 -12779 3690 -12745
rect 5616 -12773 5650 -12745
rect 5616 -12779 5650 -12773
rect 6230 -12779 6264 -12745
rect 8190 -12773 8192 -12745
rect 8192 -12773 8224 -12745
rect 8190 -12779 8224 -12773
rect 8804 -12779 8838 -12745
rect 10764 -12773 10768 -12745
rect 10768 -12773 10798 -12745
rect 10764 -12779 10798 -12773
rect 11389 -12812 11423 -12778
rect 13038 -12711 13072 -12677
rect 12558 -12773 12574 -12742
rect 12574 -12773 12592 -12742
rect 12642 -12773 12676 -12742
rect 12739 -12773 12744 -12742
rect 12744 -12773 12773 -12742
rect 12836 -12773 12846 -12742
rect 12846 -12773 12870 -12742
rect 12942 -12773 12948 -12742
rect 12948 -12773 12976 -12742
rect 12558 -12776 12592 -12773
rect 12642 -12776 12676 -12773
rect 12739 -12776 12773 -12773
rect 12836 -12776 12870 -12773
rect 12942 -12776 12976 -12773
rect 13038 -12783 13072 -12749
rect 13684 -12739 13718 -12712
rect 13684 -12746 13692 -12739
rect 13692 -12746 13718 -12739
rect 15248 -12734 15282 -12700
rect 15341 -12734 15375 -12700
rect 15248 -12830 15282 -12796
rect 15340 -12829 15374 -12795
rect -2968 -13085 -2934 -13051
rect -2876 -13085 -2842 -13051
rect -2784 -13085 -2750 -13051
rect -2692 -13085 -2658 -13051
rect -2600 -13085 -2566 -13051
rect -2508 -13085 -2474 -13051
rect -2416 -13085 -2382 -13051
rect -2324 -13085 -2290 -13051
rect -2232 -13085 -2198 -13051
rect -2140 -13085 -2106 -13051
rect -2048 -13085 -2014 -13051
rect -1956 -13085 -1922 -13051
rect -1864 -13085 -1830 -13051
rect -1772 -13085 -1738 -13051
rect -1680 -13085 -1646 -13051
rect -1588 -13085 -1554 -13051
rect -1496 -13085 -1462 -13051
rect -1404 -13085 -1370 -13051
rect -1312 -13085 -1278 -13051
rect -1220 -13085 -1186 -13051
rect -1128 -13085 -1094 -13051
rect -1036 -13085 -1002 -13051
rect -944 -13085 -910 -13051
rect -852 -13085 -818 -13051
rect -760 -13085 -726 -13051
rect -668 -13085 -634 -13051
rect -576 -13085 -542 -13051
rect -484 -13085 -450 -13051
rect -392 -13085 -358 -13051
rect -300 -13085 -266 -13051
rect -208 -13085 -174 -13051
rect -116 -13085 -82 -13051
rect -24 -13085 10 -13051
rect 68 -13085 102 -13051
rect 160 -13085 194 -13051
rect 252 -13085 286 -13051
rect 344 -13085 378 -13051
rect 436 -13085 470 -13051
rect 528 -13085 562 -13051
rect 620 -13085 654 -13051
rect 712 -13085 746 -13051
rect 804 -13085 838 -13051
rect 896 -13085 930 -13051
rect 988 -13085 1022 -13051
rect 1080 -13085 1114 -13051
rect 1172 -13085 1206 -13051
rect 1264 -13085 1298 -13051
rect 1356 -13085 1390 -13051
rect 1448 -13085 1482 -13051
rect 1540 -13085 1574 -13051
rect 1632 -13085 1666 -13051
rect 1724 -13085 1758 -13051
rect 1816 -13085 1850 -13051
rect 1908 -13085 1942 -13051
rect 2000 -13085 2034 -13051
rect 2092 -13085 2126 -13051
rect 2184 -13085 2218 -13051
rect 2276 -13085 2310 -13051
rect 2368 -13085 2402 -13051
rect 2460 -13085 2494 -13051
rect 2552 -13085 2586 -13051
rect 2644 -13085 2678 -13051
rect 2736 -13085 2770 -13051
rect 2828 -13085 2862 -13051
rect 2920 -13085 2954 -13051
rect 3012 -13085 3046 -13051
rect 3104 -13085 3138 -13051
rect 3196 -13085 3230 -13051
rect 3288 -13085 3322 -13051
rect 3380 -13085 3414 -13051
rect 3472 -13085 3506 -13051
rect 3564 -13085 3598 -13051
rect 3656 -13085 3690 -13051
rect 3748 -13085 3782 -13051
rect 3840 -13085 3874 -13051
rect 3932 -13085 3966 -13051
rect 4024 -13085 4058 -13051
rect 4116 -13085 4150 -13051
rect 4208 -13085 4242 -13051
rect 4300 -13085 4334 -13051
rect 4392 -13085 4426 -13051
rect 4484 -13085 4518 -13051
rect 4576 -13085 4610 -13051
rect 4668 -13085 4702 -13051
rect 4760 -13085 4794 -13051
rect 4852 -13085 4886 -13051
rect 4944 -13085 4978 -13051
rect 5036 -13085 5070 -13051
rect 5128 -13085 5162 -13051
rect 5220 -13085 5254 -13051
rect 5312 -13085 5346 -13051
rect 5404 -13085 5438 -13051
rect 5496 -13085 5530 -13051
rect 5588 -13085 5622 -13051
rect 5680 -13085 5714 -13051
rect 5772 -13085 5806 -13051
rect 5864 -13085 5898 -13051
rect 5956 -13085 5990 -13051
rect 6048 -13085 6082 -13051
rect 6140 -13085 6174 -13051
rect 6232 -13085 6266 -13051
rect 6324 -13085 6358 -13051
rect 6416 -13085 6450 -13051
rect 6508 -13085 6542 -13051
rect 6600 -13085 6634 -13051
rect 6692 -13085 6726 -13051
rect 6784 -13085 6818 -13051
rect 6876 -13085 6910 -13051
rect 6968 -13085 7002 -13051
rect 7060 -13085 7094 -13051
rect 7152 -13085 7186 -13051
rect 7244 -13085 7278 -13051
rect 7336 -13085 7370 -13051
rect 7428 -13085 7462 -13051
rect 7520 -13085 7554 -13051
rect 7612 -13085 7646 -13051
rect 7704 -13085 7738 -13051
rect 7796 -13085 7830 -13051
rect 7888 -13085 7922 -13051
rect 7980 -13085 8014 -13051
rect 8072 -13085 8106 -13051
rect 8164 -13085 8198 -13051
rect 8256 -13085 8290 -13051
rect 8348 -13085 8382 -13051
rect 8440 -13085 8474 -13051
rect 8532 -13085 8566 -13051
rect 8624 -13085 8658 -13051
rect 8716 -13085 8750 -13051
rect 8808 -13085 8842 -13051
rect 8900 -13085 8934 -13051
rect 8992 -13085 9026 -13051
rect 9084 -13085 9118 -13051
rect 9176 -13085 9210 -13051
rect 9268 -13085 9302 -13051
rect 9360 -13085 9394 -13051
rect 9452 -13085 9486 -13051
rect 9544 -13085 9578 -13051
rect 9636 -13085 9670 -13051
rect 9728 -13085 9762 -13051
rect 9820 -13085 9854 -13051
rect 9912 -13085 9946 -13051
rect 10004 -13085 10038 -13051
rect 10096 -13085 10130 -13051
rect 10188 -13085 10222 -13051
rect 10280 -13085 10314 -13051
rect 10372 -13085 10406 -13051
rect 10464 -13085 10498 -13051
rect 10556 -13085 10590 -13051
rect 10648 -13085 10682 -13051
rect 10740 -13085 10774 -13051
rect 10832 -13085 10866 -13051
rect 10924 -13085 10958 -13051
rect 11016 -13085 11050 -13051
rect 11108 -13085 11142 -13051
rect 11200 -13085 11234 -13051
rect 11292 -13085 11326 -13051
rect 11384 -13085 11418 -13051
rect 11476 -13085 11510 -13051
rect 11568 -13085 11602 -13051
rect 11660 -13085 11694 -13051
rect 11752 -13085 11786 -13051
rect 11844 -13085 11878 -13051
rect 11936 -13085 11970 -13051
rect 12028 -13085 12062 -13051
rect 12120 -13085 12154 -13051
rect 12212 -13085 12246 -13051
rect 12304 -13085 12338 -13051
rect 12396 -13085 12430 -13051
rect 12488 -13085 12522 -13051
rect 12580 -13085 12614 -13051
rect 12672 -13085 12706 -13051
rect 12764 -13085 12798 -13051
rect 12856 -13085 12890 -13051
rect 12948 -13085 12982 -13051
rect 13040 -13085 13074 -13051
rect 13132 -13085 13166 -13051
rect 13224 -13085 13258 -13051
rect 13316 -13085 13350 -13051
rect 13408 -13085 13442 -13051
rect 13500 -13085 13534 -13051
rect 13592 -13085 13626 -13051
rect 13684 -13085 13718 -13051
rect 13776 -13085 13810 -13051
rect 13868 -13085 13902 -13051
rect 13960 -13085 13994 -13051
rect 14052 -13085 14086 -13051
rect 14144 -13085 14178 -13051
rect 14236 -13085 14270 -13051
rect 14328 -13085 14362 -13051
rect 14420 -13085 14454 -13051
rect 14512 -13085 14546 -13051
rect 14604 -13085 14638 -13051
rect 14696 -13085 14730 -13051
rect 14788 -13085 14822 -13051
rect 14880 -13085 14914 -13051
rect 14972 -13085 15006 -13051
rect 15064 -13085 15098 -13051
rect 15156 -13085 15190 -13051
rect 15248 -13085 15282 -13051
rect 15340 -13085 15374 -13051
rect 15432 -13085 15466 -13051
rect 15524 -13085 15558 -13051
rect 15616 -13085 15650 -13051
rect 15708 -13085 15742 -13051
rect 15800 -13085 15834 -13051
rect 15892 -13085 15926 -13051
rect 15984 -13085 16018 -13051
rect 16076 -13085 16110 -13051
rect 16168 -13085 16202 -13051
rect 16260 -13085 16294 -13051
rect 16352 -13085 16386 -13051
rect 16444 -13085 16478 -13051
rect 16536 -13085 16570 -13051
rect 16628 -13085 16662 -13051
rect 432 -13358 466 -13324
rect 1052 -13363 1086 -13359
rect 1052 -13393 1086 -13363
rect 3012 -13393 3046 -13359
rect 3626 -13363 3660 -13359
rect 3626 -13393 3628 -13363
rect 3628 -13393 3660 -13363
rect 5586 -13393 5620 -13359
rect 6200 -13363 6234 -13359
rect 6200 -13393 6204 -13363
rect 6204 -13393 6234 -13363
rect 8160 -13393 8194 -13359
rect 8774 -13363 8808 -13359
rect 8774 -13393 8780 -13363
rect 8780 -13393 8808 -13363
rect 10737 -13391 10771 -13357
rect 11369 -13363 11403 -13356
rect 11369 -13390 11390 -13363
rect 11390 -13390 11403 -13363
rect 15248 -13344 15282 -13310
rect 15341 -13344 15375 -13310
rect 13685 -13397 13692 -13388
rect 13692 -13397 13719 -13388
rect 13685 -13422 13719 -13397
rect 15248 -13440 15282 -13406
rect 15340 -13439 15374 -13405
rect -2968 -13629 -2934 -13595
rect -2876 -13629 -2842 -13595
rect -2784 -13629 -2750 -13595
rect -2692 -13629 -2658 -13595
rect -2600 -13629 -2566 -13595
rect -2508 -13629 -2474 -13595
rect -2416 -13629 -2382 -13595
rect -2324 -13629 -2290 -13595
rect -2232 -13629 -2198 -13595
rect -2140 -13629 -2106 -13595
rect -2048 -13629 -2014 -13595
rect -1956 -13629 -1922 -13595
rect -1864 -13629 -1830 -13595
rect -1772 -13629 -1738 -13595
rect -1680 -13629 -1646 -13595
rect -1588 -13629 -1554 -13595
rect -1496 -13629 -1462 -13595
rect -1404 -13629 -1370 -13595
rect -1312 -13629 -1278 -13595
rect -1220 -13629 -1186 -13595
rect -1128 -13629 -1094 -13595
rect -1036 -13629 -1002 -13595
rect -944 -13629 -910 -13595
rect -852 -13629 -818 -13595
rect -760 -13629 -726 -13595
rect -668 -13629 -634 -13595
rect -576 -13629 -542 -13595
rect -484 -13629 -450 -13595
rect -392 -13629 -358 -13595
rect -300 -13629 -266 -13595
rect -208 -13629 -174 -13595
rect -116 -13629 -82 -13595
rect -24 -13629 10 -13595
rect 68 -13629 102 -13595
rect 160 -13629 194 -13595
rect 252 -13629 286 -13595
rect 344 -13629 378 -13595
rect 436 -13629 470 -13595
rect 528 -13629 562 -13595
rect 620 -13629 654 -13595
rect 712 -13629 746 -13595
rect 804 -13629 838 -13595
rect 896 -13629 930 -13595
rect 988 -13629 1022 -13595
rect 1080 -13629 1114 -13595
rect 1172 -13629 1206 -13595
rect 1264 -13629 1298 -13595
rect 1356 -13629 1390 -13595
rect 1448 -13629 1482 -13595
rect 1540 -13629 1574 -13595
rect 1632 -13629 1666 -13595
rect 1724 -13629 1758 -13595
rect 1816 -13629 1850 -13595
rect 1908 -13629 1942 -13595
rect 2000 -13629 2034 -13595
rect 2092 -13629 2126 -13595
rect 2184 -13629 2218 -13595
rect 2276 -13629 2310 -13595
rect 2368 -13629 2402 -13595
rect 2460 -13629 2494 -13595
rect 2552 -13629 2586 -13595
rect 2644 -13629 2678 -13595
rect 2736 -13629 2770 -13595
rect 2828 -13629 2862 -13595
rect 2920 -13629 2954 -13595
rect 3012 -13629 3046 -13595
rect 3104 -13629 3138 -13595
rect 3196 -13629 3230 -13595
rect 3288 -13629 3322 -13595
rect 3380 -13629 3414 -13595
rect 3472 -13629 3506 -13595
rect 3564 -13629 3598 -13595
rect 3656 -13629 3690 -13595
rect 3748 -13629 3782 -13595
rect 3840 -13629 3874 -13595
rect 3932 -13629 3966 -13595
rect 4024 -13629 4058 -13595
rect 4116 -13629 4150 -13595
rect 4208 -13629 4242 -13595
rect 4300 -13629 4334 -13595
rect 4392 -13629 4426 -13595
rect 4484 -13629 4518 -13595
rect 4576 -13629 4610 -13595
rect 4668 -13629 4702 -13595
rect 4760 -13629 4794 -13595
rect 4852 -13629 4886 -13595
rect 4944 -13629 4978 -13595
rect 5036 -13629 5070 -13595
rect 5128 -13629 5162 -13595
rect 5220 -13629 5254 -13595
rect 5312 -13629 5346 -13595
rect 5404 -13629 5438 -13595
rect 5496 -13629 5530 -13595
rect 5588 -13629 5622 -13595
rect 5680 -13629 5714 -13595
rect 5772 -13629 5806 -13595
rect 5864 -13629 5898 -13595
rect 5956 -13629 5990 -13595
rect 6048 -13629 6082 -13595
rect 6140 -13629 6174 -13595
rect 6232 -13629 6266 -13595
rect 6324 -13629 6358 -13595
rect 6416 -13629 6450 -13595
rect 6508 -13629 6542 -13595
rect 6600 -13629 6634 -13595
rect 6692 -13629 6726 -13595
rect 6784 -13629 6818 -13595
rect 6876 -13629 6910 -13595
rect 6968 -13629 7002 -13595
rect 7060 -13629 7094 -13595
rect 7152 -13629 7186 -13595
rect 7244 -13629 7278 -13595
rect 7336 -13629 7370 -13595
rect 7428 -13629 7462 -13595
rect 7520 -13629 7554 -13595
rect 7612 -13629 7646 -13595
rect 7704 -13629 7738 -13595
rect 7796 -13629 7830 -13595
rect 7888 -13629 7922 -13595
rect 7980 -13629 8014 -13595
rect 8072 -13629 8106 -13595
rect 8164 -13629 8198 -13595
rect 8256 -13629 8290 -13595
rect 8348 -13629 8382 -13595
rect 8440 -13629 8474 -13595
rect 8532 -13629 8566 -13595
rect 8624 -13629 8658 -13595
rect 8716 -13629 8750 -13595
rect 8808 -13629 8842 -13595
rect 8900 -13629 8934 -13595
rect 8992 -13629 9026 -13595
rect 9084 -13629 9118 -13595
rect 9176 -13629 9210 -13595
rect 9268 -13629 9302 -13595
rect 9360 -13629 9394 -13595
rect 9452 -13629 9486 -13595
rect 9544 -13629 9578 -13595
rect 9636 -13629 9670 -13595
rect 9728 -13629 9762 -13595
rect 9820 -13629 9854 -13595
rect 9912 -13629 9946 -13595
rect 10004 -13629 10038 -13595
rect 10096 -13629 10130 -13595
rect 10188 -13629 10222 -13595
rect 10280 -13629 10314 -13595
rect 10372 -13629 10406 -13595
rect 10464 -13629 10498 -13595
rect 10556 -13629 10590 -13595
rect 10648 -13629 10682 -13595
rect 10740 -13629 10774 -13595
rect 10832 -13629 10866 -13595
rect 10924 -13629 10958 -13595
rect 11016 -13629 11050 -13595
rect 11108 -13629 11142 -13595
rect 11200 -13629 11234 -13595
rect 11292 -13629 11326 -13595
rect 11384 -13629 11418 -13595
rect 11476 -13629 11510 -13595
rect 11568 -13629 11602 -13595
rect 11660 -13629 11694 -13595
rect 11752 -13629 11786 -13595
rect 11844 -13629 11878 -13595
rect 11936 -13629 11970 -13595
rect 12028 -13629 12062 -13595
rect 12120 -13629 12154 -13595
rect 12212 -13629 12246 -13595
rect 12304 -13629 12338 -13595
rect 12396 -13629 12430 -13595
rect 12488 -13629 12522 -13595
rect 12580 -13629 12614 -13595
rect 12672 -13629 12706 -13595
rect 12764 -13629 12798 -13595
rect 12856 -13629 12890 -13595
rect 12948 -13629 12982 -13595
rect 13040 -13629 13074 -13595
rect 13132 -13629 13166 -13595
rect 13224 -13629 13258 -13595
rect 13316 -13629 13350 -13595
rect 13408 -13629 13442 -13595
rect 13500 -13629 13534 -13595
rect 13592 -13629 13626 -13595
rect 13684 -13629 13718 -13595
rect 13776 -13629 13810 -13595
rect 13868 -13629 13902 -13595
rect 13960 -13629 13994 -13595
rect 14052 -13629 14086 -13595
rect 14144 -13629 14178 -13595
rect 14236 -13629 14270 -13595
rect 14328 -13629 14362 -13595
rect 14420 -13629 14454 -13595
rect 14512 -13629 14546 -13595
rect 14604 -13629 14638 -13595
rect 14696 -13629 14730 -13595
rect 14788 -13629 14822 -13595
rect 14880 -13629 14914 -13595
rect 14972 -13629 15006 -13595
rect 15064 -13629 15098 -13595
rect 15156 -13629 15190 -13595
rect 15248 -13629 15282 -13595
rect 15340 -13629 15374 -13595
rect 15432 -13629 15466 -13595
rect 15524 -13629 15558 -13595
rect 15616 -13629 15650 -13595
rect 15708 -13629 15742 -13595
rect 15800 -13629 15834 -13595
rect 15892 -13629 15926 -13595
rect 15984 -13629 16018 -13595
rect 16076 -13629 16110 -13595
rect 16168 -13629 16202 -13595
rect 16260 -13629 16294 -13595
rect 16352 -13629 16386 -13595
rect 16444 -13629 16478 -13595
rect 16536 -13629 16570 -13595
rect 16628 -13629 16662 -13595
rect -848 -13756 -814 -13722
rect -769 -13739 -735 -13722
rect -769 -13756 -766 -13739
rect -766 -13756 -735 -13739
rect -932 -13861 -903 -13834
rect -903 -13861 -898 -13834
rect -932 -13868 -898 -13861
rect -764 -13861 -735 -13835
rect -735 -13861 -730 -13835
rect -764 -13869 -730 -13861
rect 434 -13823 468 -13789
rect -30 -13861 4 -13827
rect 106 -13861 140 -13827
rect 242 -13861 276 -13827
rect 1076 -13783 1110 -13749
rect 1076 -13827 1110 -13822
rect 1076 -13856 1082 -13827
rect 1082 -13856 1110 -13827
rect 1171 -13862 1205 -13828
rect 1263 -13862 1297 -13828
rect 2369 -13861 2396 -13833
rect 2396 -13861 2403 -13833
rect 2369 -13867 2403 -13861
rect 3015 -13866 3049 -13832
rect 6876 -13861 6904 -13832
rect 6904 -13861 6910 -13832
rect 6876 -13866 6910 -13861
rect 7522 -13866 7556 -13832
rect 8164 -13861 8192 -13831
rect 8192 -13861 8198 -13831
rect 8164 -13865 8198 -13861
rect 8811 -13867 8845 -13833
rect 9453 -13861 9480 -13833
rect 9480 -13861 9487 -13833
rect 9453 -13867 9487 -13861
rect 10099 -13868 10133 -13834
rect 10741 -13861 10749 -13833
rect 10749 -13861 10775 -13833
rect 10832 -13861 10864 -13833
rect 10864 -13861 10866 -13833
rect 10925 -13861 10948 -13832
rect 10948 -13861 10959 -13832
rect 11017 -13861 11032 -13832
rect 11032 -13861 11051 -13832
rect 10741 -13867 10775 -13861
rect 10832 -13867 10866 -13861
rect 10925 -13866 10959 -13861
rect 11017 -13866 11051 -13861
rect 11129 -13900 11163 -13866
rect 11250 -13861 11284 -13835
rect 11344 -13861 11368 -13835
rect 11368 -13861 11378 -13835
rect 11250 -13869 11284 -13861
rect 11344 -13869 11378 -13861
rect -2968 -14173 -2934 -14139
rect -2876 -14173 -2842 -14139
rect -2784 -14173 -2750 -14139
rect -2692 -14173 -2658 -14139
rect -2600 -14173 -2566 -14139
rect -2508 -14173 -2474 -14139
rect -2416 -14173 -2382 -14139
rect -2324 -14173 -2290 -14139
rect -2232 -14173 -2198 -14139
rect -2140 -14173 -2106 -14139
rect -2048 -14173 -2014 -14139
rect -1956 -14173 -1922 -14139
rect -1864 -14173 -1830 -14139
rect -1772 -14173 -1738 -14139
rect -1680 -14173 -1646 -14139
rect -1588 -14173 -1554 -14139
rect -1496 -14173 -1462 -14139
rect -1404 -14173 -1370 -14139
rect -1312 -14173 -1278 -14139
rect -1220 -14173 -1186 -14139
rect -1128 -14173 -1094 -14139
rect -1036 -14173 -1002 -14139
rect -944 -14173 -910 -14139
rect -852 -14173 -818 -14139
rect -760 -14173 -726 -14139
rect -668 -14173 -634 -14139
rect -576 -14173 -542 -14139
rect -484 -14173 -450 -14139
rect -392 -14173 -358 -14139
rect -300 -14173 -266 -14139
rect -208 -14173 -174 -14139
rect -116 -14173 -82 -14139
rect -24 -14173 10 -14139
rect 68 -14173 102 -14139
rect 160 -14173 194 -14139
rect 252 -14173 286 -14139
rect 344 -14173 378 -14139
rect 436 -14173 470 -14139
rect 528 -14173 562 -14139
rect 620 -14173 654 -14139
rect 712 -14173 746 -14139
rect 804 -14173 838 -14139
rect 896 -14173 930 -14139
rect 988 -14173 1022 -14139
rect 1080 -14173 1114 -14139
rect 1172 -14173 1206 -14139
rect 1264 -14173 1298 -14139
rect 1356 -14173 1390 -14139
rect 1448 -14173 1482 -14139
rect 1540 -14173 1574 -14139
rect 1632 -14173 1666 -14139
rect 1724 -14173 1758 -14139
rect 1816 -14173 1850 -14139
rect 1908 -14173 1942 -14139
rect 2000 -14173 2034 -14139
rect 2092 -14173 2126 -14139
rect 2184 -14173 2218 -14139
rect 2276 -14173 2310 -14139
rect 2368 -14173 2402 -14139
rect 2460 -14173 2494 -14139
rect 2552 -14173 2586 -14139
rect 2644 -14173 2678 -14139
rect 2736 -14173 2770 -14139
rect 2828 -14173 2862 -14139
rect 2920 -14173 2954 -14139
rect 3012 -14173 3046 -14139
rect 3104 -14173 3138 -14139
rect 3196 -14173 3230 -14139
rect 3288 -14173 3322 -14139
rect 3380 -14173 3414 -14139
rect 3472 -14173 3506 -14139
rect 3564 -14173 3598 -14139
rect 3656 -14173 3690 -14139
rect 3748 -14173 3782 -14139
rect 3840 -14173 3874 -14139
rect 3932 -14173 3966 -14139
rect 4024 -14173 4058 -14139
rect 4116 -14173 4150 -14139
rect 4208 -14173 4242 -14139
rect 4300 -14173 4334 -14139
rect 4392 -14173 4426 -14139
rect 4484 -14173 4518 -14139
rect 4576 -14173 4610 -14139
rect 4668 -14173 4702 -14139
rect 4760 -14173 4794 -14139
rect 4852 -14173 4886 -14139
rect 4944 -14173 4978 -14139
rect 5036 -14173 5070 -14139
rect 5128 -14173 5162 -14139
rect 5220 -14173 5254 -14139
rect 5312 -14173 5346 -14139
rect 5404 -14173 5438 -14139
rect 5496 -14173 5530 -14139
rect 5588 -14173 5622 -14139
rect 5680 -14173 5714 -14139
rect 5772 -14173 5806 -14139
rect 5864 -14173 5898 -14139
rect 5956 -14173 5990 -14139
rect 6048 -14173 6082 -14139
rect 6140 -14173 6174 -14139
rect 6232 -14173 6266 -14139
rect 6324 -14173 6358 -14139
rect 6416 -14173 6450 -14139
rect 6508 -14173 6542 -14139
rect 6600 -14173 6634 -14139
rect 6692 -14173 6726 -14139
rect 6784 -14173 6818 -14139
rect 6876 -14173 6910 -14139
rect 6968 -14173 7002 -14139
rect 7060 -14173 7094 -14139
rect 7152 -14173 7186 -14139
rect 7244 -14173 7278 -14139
rect 7336 -14173 7370 -14139
rect 7428 -14173 7462 -14139
rect 7520 -14173 7554 -14139
rect 7612 -14173 7646 -14139
rect 7704 -14173 7738 -14139
rect 7796 -14173 7830 -14139
rect 7888 -14173 7922 -14139
rect 7980 -14173 8014 -14139
rect 8072 -14173 8106 -14139
rect 8164 -14173 8198 -14139
rect 8256 -14173 8290 -14139
rect 8348 -14173 8382 -14139
rect 8440 -14173 8474 -14139
rect 8532 -14173 8566 -14139
rect 8624 -14173 8658 -14139
rect 8716 -14173 8750 -14139
rect 8808 -14173 8842 -14139
rect 8900 -14173 8934 -14139
rect 8992 -14173 9026 -14139
rect 9084 -14173 9118 -14139
rect 9176 -14173 9210 -14139
rect 9268 -14173 9302 -14139
rect 9360 -14173 9394 -14139
rect 9452 -14173 9486 -14139
rect 9544 -14173 9578 -14139
rect 9636 -14173 9670 -14139
rect 9728 -14173 9762 -14139
rect 9820 -14173 9854 -14139
rect 9912 -14173 9946 -14139
rect 10004 -14173 10038 -14139
rect 10096 -14173 10130 -14139
rect 10188 -14173 10222 -14139
rect 10280 -14173 10314 -14139
rect 10372 -14173 10406 -14139
rect 10464 -14173 10498 -14139
rect 10556 -14173 10590 -14139
rect 10648 -14173 10682 -14139
rect 10740 -14173 10774 -14139
rect 10832 -14173 10866 -14139
rect 10924 -14173 10958 -14139
rect 11016 -14173 11050 -14139
rect 11108 -14173 11142 -14139
rect 11200 -14173 11234 -14139
rect 11292 -14173 11326 -14139
rect 11384 -14173 11418 -14139
rect 11476 -14173 11510 -14139
rect 11568 -14173 11602 -14139
rect 11660 -14173 11694 -14139
rect 11752 -14173 11786 -14139
rect 11844 -14173 11878 -14139
rect 11936 -14173 11970 -14139
rect 12028 -14173 12062 -14139
rect 12120 -14173 12154 -14139
rect 12212 -14173 12246 -14139
rect 12304 -14173 12338 -14139
rect 12396 -14173 12430 -14139
rect 12488 -14173 12522 -14139
rect 12580 -14173 12614 -14139
rect 12672 -14173 12706 -14139
rect 12764 -14173 12798 -14139
rect 12856 -14173 12890 -14139
rect 12948 -14173 12982 -14139
rect 13040 -14173 13074 -14139
rect 13132 -14173 13166 -14139
rect 13224 -14173 13258 -14139
rect 13316 -14173 13350 -14139
rect 13408 -14173 13442 -14139
rect 13500 -14173 13534 -14139
rect 13592 -14173 13626 -14139
rect 13684 -14173 13718 -14139
rect 13776 -14173 13810 -14139
rect 13868 -14173 13902 -14139
rect 13960 -14173 13994 -14139
rect 14052 -14173 14086 -14139
rect 14144 -14173 14178 -14139
rect 14236 -14173 14270 -14139
rect 14328 -14173 14362 -14139
rect 14420 -14173 14454 -14139
rect 14512 -14173 14546 -14139
rect 14604 -14173 14638 -14139
rect 14696 -14173 14730 -14139
rect 14788 -14173 14822 -14139
rect 14880 -14173 14914 -14139
rect 14972 -14173 15006 -14139
rect 15064 -14173 15098 -14139
rect 15156 -14173 15190 -14139
rect 15248 -14173 15282 -14139
rect 15340 -14173 15374 -14139
rect 15432 -14173 15466 -14139
rect 15524 -14173 15558 -14139
rect 15616 -14173 15650 -14139
rect 15708 -14173 15742 -14139
rect 15800 -14173 15834 -14139
rect 15892 -14173 15926 -14139
rect 15984 -14173 16018 -14139
rect 16076 -14173 16110 -14139
rect 16168 -14173 16202 -14139
rect 16260 -14173 16294 -14139
rect 16352 -14173 16386 -14139
rect 16444 -14173 16478 -14139
rect 16536 -14173 16570 -14139
rect 16628 -14173 16662 -14139
<< metal1 >>
rect -3193 5 16946 36
rect -3193 -29 -2968 5
rect -2934 -29 -2876 5
rect -2842 -29 -2784 5
rect -2750 -29 -2692 5
rect -2658 -29 -2600 5
rect -2566 -29 -2508 5
rect -2474 -29 -2416 5
rect -2382 -29 -2324 5
rect -2290 -29 -2232 5
rect -2198 -29 -2140 5
rect -2106 -29 -2048 5
rect -2014 -29 -1956 5
rect -1922 -29 -1864 5
rect -1830 -29 -1772 5
rect -1738 -29 -1680 5
rect -1646 -29 -1588 5
rect -1554 -29 -1496 5
rect -1462 -29 -1404 5
rect -1370 -29 -1312 5
rect -1278 -29 -1220 5
rect -1186 -29 -1128 5
rect -1094 -29 -1036 5
rect -1002 -29 -944 5
rect -910 -29 -852 5
rect -818 -29 -760 5
rect -726 -29 -668 5
rect -634 -29 -576 5
rect -542 -29 -484 5
rect -450 -29 -392 5
rect -358 -29 -300 5
rect -266 -29 -208 5
rect -174 -29 -116 5
rect -82 -29 -24 5
rect 10 -29 68 5
rect 102 -29 160 5
rect 194 -29 252 5
rect 286 -29 344 5
rect 378 -29 436 5
rect 470 -29 528 5
rect 562 -29 620 5
rect 654 -29 712 5
rect 746 -29 804 5
rect 838 -29 896 5
rect 930 -29 988 5
rect 1022 -29 1080 5
rect 1114 -29 1172 5
rect 1206 -29 1264 5
rect 1298 -29 1356 5
rect 1390 -29 1448 5
rect 1482 -29 1540 5
rect 1574 -29 1632 5
rect 1666 -29 1724 5
rect 1758 -29 1816 5
rect 1850 -29 1908 5
rect 1942 -29 2000 5
rect 2034 -29 2092 5
rect 2126 -29 2184 5
rect 2218 -29 2276 5
rect 2310 -29 2368 5
rect 2402 -29 2460 5
rect 2494 -29 2552 5
rect 2586 -29 2644 5
rect 2678 -29 2736 5
rect 2770 -29 2828 5
rect 2862 -29 2920 5
rect 2954 -29 3012 5
rect 3046 -29 3104 5
rect 3138 -29 3196 5
rect 3230 -29 3288 5
rect 3322 -29 3380 5
rect 3414 -29 3472 5
rect 3506 -29 3564 5
rect 3598 -29 3656 5
rect 3690 -29 3748 5
rect 3782 -29 3840 5
rect 3874 -29 3932 5
rect 3966 -29 4024 5
rect 4058 -29 4116 5
rect 4150 -29 4208 5
rect 4242 -29 4300 5
rect 4334 -29 4392 5
rect 4426 -29 4484 5
rect 4518 -29 4576 5
rect 4610 -29 4668 5
rect 4702 -29 4760 5
rect 4794 -29 4852 5
rect 4886 -29 4944 5
rect 4978 -29 5036 5
rect 5070 -29 5128 5
rect 5162 -29 5220 5
rect 5254 -29 5312 5
rect 5346 -29 5404 5
rect 5438 -29 5496 5
rect 5530 -29 5588 5
rect 5622 -29 5680 5
rect 5714 -29 5772 5
rect 5806 -29 5864 5
rect 5898 -29 5956 5
rect 5990 -29 6048 5
rect 6082 -29 6140 5
rect 6174 -29 6232 5
rect 6266 -29 6324 5
rect 6358 -29 6416 5
rect 6450 -29 6508 5
rect 6542 -29 6600 5
rect 6634 -29 6692 5
rect 6726 -29 6784 5
rect 6818 -29 6876 5
rect 6910 -29 6968 5
rect 7002 -29 7060 5
rect 7094 -29 7152 5
rect 7186 -29 7244 5
rect 7278 -29 7336 5
rect 7370 -29 7428 5
rect 7462 -29 7520 5
rect 7554 -29 7612 5
rect 7646 -29 7704 5
rect 7738 -29 7796 5
rect 7830 -29 7888 5
rect 7922 -29 7980 5
rect 8014 -29 8072 5
rect 8106 -29 8164 5
rect 8198 -29 8256 5
rect 8290 -29 8348 5
rect 8382 -29 8440 5
rect 8474 -29 8532 5
rect 8566 -29 8624 5
rect 8658 -29 8716 5
rect 8750 -29 8808 5
rect 8842 -29 8900 5
rect 8934 -29 8992 5
rect 9026 -29 9084 5
rect 9118 -29 9176 5
rect 9210 -29 9268 5
rect 9302 -29 9360 5
rect 9394 -29 9452 5
rect 9486 -29 9544 5
rect 9578 -29 9636 5
rect 9670 -29 9728 5
rect 9762 -29 9820 5
rect 9854 -29 9912 5
rect 9946 -29 10004 5
rect 10038 -29 10096 5
rect 10130 -29 10188 5
rect 10222 -29 10280 5
rect 10314 -29 10372 5
rect 10406 -29 10464 5
rect 10498 -29 10556 5
rect 10590 -29 10648 5
rect 10682 -29 10740 5
rect 10774 -29 10832 5
rect 10866 -29 10924 5
rect 10958 -29 11016 5
rect 11050 -29 11108 5
rect 11142 -29 11200 5
rect 11234 -29 11292 5
rect 11326 -29 11384 5
rect 11418 -29 11476 5
rect 11510 -29 11568 5
rect 11602 -29 11660 5
rect 11694 -29 11752 5
rect 11786 -29 11844 5
rect 11878 -29 11936 5
rect 11970 -29 12028 5
rect 12062 -29 12120 5
rect 12154 -29 12212 5
rect 12246 -29 12304 5
rect 12338 -29 12396 5
rect 12430 -29 12488 5
rect 12522 -29 12580 5
rect 12614 -29 12672 5
rect 12706 -29 12764 5
rect 12798 -29 12856 5
rect 12890 -29 12948 5
rect 12982 -29 13040 5
rect 13074 -29 13132 5
rect 13166 -29 13224 5
rect 13258 -29 13316 5
rect 13350 -29 13408 5
rect 13442 -29 13500 5
rect 13534 -29 13592 5
rect 13626 -29 13684 5
rect 13718 -29 13776 5
rect 13810 -29 13868 5
rect 13902 -29 13960 5
rect 13994 -29 14052 5
rect 14086 -29 14144 5
rect 14178 -29 14236 5
rect 14270 -29 14328 5
rect 14362 -29 14420 5
rect 14454 -29 14512 5
rect 14546 -29 14604 5
rect 14638 -29 14696 5
rect 14730 -29 14788 5
rect 14822 -29 14880 5
rect 14914 -29 14972 5
rect 15006 -29 15064 5
rect 15098 -29 15156 5
rect 15190 -29 15248 5
rect 15282 -29 15340 5
rect 15374 -29 15432 5
rect 15466 -29 15524 5
rect 15558 -29 15616 5
rect 15650 -29 15708 5
rect 15742 -29 15800 5
rect 15834 -29 15892 5
rect 15926 -29 15984 5
rect 16018 -29 16076 5
rect 16110 -29 16168 5
rect 16202 -29 16260 5
rect 16294 -29 16352 5
rect 16386 -29 16444 5
rect 16478 -29 16536 5
rect 16570 -29 16628 5
rect 16662 -29 16946 5
rect -3193 -60 16946 -29
rect 308 -212 11419 -127
rect -1802 -343 -1792 -291
rect -1740 -294 -1730 -291
rect -1740 -301 -896 -294
rect -1740 -335 -943 -301
rect -909 -335 -896 -301
rect -1740 -342 -896 -335
rect -781 -342 -771 -290
rect -719 -342 -709 -290
rect 308 -298 387 -212
rect 1153 -284 1310 -283
rect -57 -307 389 -298
rect -57 -341 -30 -307
rect 4 -341 106 -307
rect 140 -341 242 -307
rect 276 -341 389 -307
rect -1740 -343 -1730 -342
rect -57 -346 389 -341
rect -57 -347 16 -346
rect 94 -347 152 -346
rect 227 -347 389 -346
rect 418 -312 1122 -294
rect 418 -325 1076 -312
rect 418 -345 982 -325
rect -57 -403 12 -347
rect 418 -379 434 -345
rect 468 -377 982 -345
rect 1034 -346 1076 -325
rect 1110 -346 1122 -312
rect 1034 -377 1122 -346
rect 468 -379 1122 -377
rect 418 -385 1122 -379
rect -862 -412 13 -403
rect 418 -405 1076 -385
rect 418 -409 485 -405
rect -862 -446 -848 -412
rect -814 -446 -769 -412
rect -735 -446 13 -412
rect -862 -452 13 -446
rect 1064 -419 1076 -405
rect 1110 -419 1122 -385
rect 1153 -301 2449 -284
rect 1153 -306 2369 -301
rect 1153 -340 1171 -306
rect 1205 -340 1263 -306
rect 1297 -335 2369 -306
rect 2403 -335 2449 -301
rect 1297 -340 2449 -335
rect 1153 -346 2449 -340
rect 2994 -302 6963 -282
rect 2994 -336 3015 -302
rect 3049 -336 6876 -302
rect 6910 -336 6963 -302
rect 1153 -406 1310 -346
rect 2994 -353 6963 -336
rect 7509 -302 8255 -281
rect 7509 -336 7522 -302
rect 7556 -303 8255 -302
rect 7556 -336 8164 -303
rect 7509 -337 8164 -336
rect 8198 -337 8255 -303
rect 7509 -355 8255 -337
rect 8799 -301 9545 -283
rect 8799 -335 8811 -301
rect 8845 -335 9453 -301
rect 9487 -335 9545 -301
rect 8799 -354 9545 -335
rect 10086 -296 11058 -278
rect 10086 -300 11063 -296
rect 10086 -334 10099 -300
rect 10133 -301 11063 -300
rect 10133 -334 10741 -301
rect 10086 -335 10741 -334
rect 10775 -335 10832 -301
rect 10866 -302 11063 -301
rect 10866 -335 10925 -302
rect 10086 -336 10925 -335
rect 10959 -336 11017 -302
rect 11051 -336 11063 -302
rect 11110 -311 11120 -259
rect 11172 -311 11182 -259
rect 11233 -299 11418 -212
rect 10086 -342 11063 -336
rect 11233 -333 11250 -299
rect 11284 -333 11344 -299
rect 11378 -333 11418 -299
rect 11233 -341 11418 -333
rect 10086 -348 11058 -342
rect 1064 -474 1122 -419
rect 1070 -478 1116 -474
rect -3193 -539 16946 -508
rect -3193 -573 -2968 -539
rect -2934 -573 -2876 -539
rect -2842 -573 -2784 -539
rect -2750 -573 -2692 -539
rect -2658 -573 -2600 -539
rect -2566 -573 -2508 -539
rect -2474 -573 -2416 -539
rect -2382 -573 -2324 -539
rect -2290 -573 -2232 -539
rect -2198 -573 -2140 -539
rect -2106 -573 -2048 -539
rect -2014 -573 -1956 -539
rect -1922 -573 -1864 -539
rect -1830 -573 -1772 -539
rect -1738 -573 -1680 -539
rect -1646 -573 -1588 -539
rect -1554 -573 -1496 -539
rect -1462 -573 -1404 -539
rect -1370 -573 -1312 -539
rect -1278 -573 -1220 -539
rect -1186 -573 -1128 -539
rect -1094 -573 -1036 -539
rect -1002 -573 -944 -539
rect -910 -573 -852 -539
rect -818 -573 -760 -539
rect -726 -573 -668 -539
rect -634 -573 -576 -539
rect -542 -573 -484 -539
rect -450 -573 -392 -539
rect -358 -573 -300 -539
rect -266 -573 -208 -539
rect -174 -573 -116 -539
rect -82 -573 -24 -539
rect 10 -573 68 -539
rect 102 -573 160 -539
rect 194 -573 252 -539
rect 286 -573 344 -539
rect 378 -573 436 -539
rect 470 -573 528 -539
rect 562 -573 620 -539
rect 654 -573 712 -539
rect 746 -573 804 -539
rect 838 -573 896 -539
rect 930 -573 988 -539
rect 1022 -573 1080 -539
rect 1114 -573 1172 -539
rect 1206 -573 1264 -539
rect 1298 -573 1356 -539
rect 1390 -573 1448 -539
rect 1482 -573 1540 -539
rect 1574 -573 1632 -539
rect 1666 -573 1724 -539
rect 1758 -573 1816 -539
rect 1850 -573 1908 -539
rect 1942 -573 2000 -539
rect 2034 -573 2092 -539
rect 2126 -573 2184 -539
rect 2218 -573 2276 -539
rect 2310 -573 2368 -539
rect 2402 -573 2460 -539
rect 2494 -573 2552 -539
rect 2586 -573 2644 -539
rect 2678 -573 2736 -539
rect 2770 -573 2828 -539
rect 2862 -573 2920 -539
rect 2954 -573 3012 -539
rect 3046 -573 3104 -539
rect 3138 -573 3196 -539
rect 3230 -573 3288 -539
rect 3322 -573 3380 -539
rect 3414 -573 3472 -539
rect 3506 -573 3564 -539
rect 3598 -573 3656 -539
rect 3690 -573 3748 -539
rect 3782 -573 3840 -539
rect 3874 -573 3932 -539
rect 3966 -573 4024 -539
rect 4058 -573 4116 -539
rect 4150 -573 4208 -539
rect 4242 -573 4300 -539
rect 4334 -573 4392 -539
rect 4426 -573 4484 -539
rect 4518 -573 4576 -539
rect 4610 -573 4668 -539
rect 4702 -573 4760 -539
rect 4794 -573 4852 -539
rect 4886 -573 4944 -539
rect 4978 -573 5036 -539
rect 5070 -573 5128 -539
rect 5162 -573 5220 -539
rect 5254 -573 5312 -539
rect 5346 -573 5404 -539
rect 5438 -573 5496 -539
rect 5530 -573 5588 -539
rect 5622 -573 5680 -539
rect 5714 -573 5772 -539
rect 5806 -573 5864 -539
rect 5898 -573 5956 -539
rect 5990 -573 6048 -539
rect 6082 -573 6140 -539
rect 6174 -573 6232 -539
rect 6266 -573 6324 -539
rect 6358 -573 6416 -539
rect 6450 -573 6508 -539
rect 6542 -573 6600 -539
rect 6634 -573 6692 -539
rect 6726 -573 6784 -539
rect 6818 -573 6876 -539
rect 6910 -573 6968 -539
rect 7002 -573 7060 -539
rect 7094 -573 7152 -539
rect 7186 -573 7244 -539
rect 7278 -573 7336 -539
rect 7370 -573 7428 -539
rect 7462 -573 7520 -539
rect 7554 -573 7612 -539
rect 7646 -573 7704 -539
rect 7738 -573 7796 -539
rect 7830 -573 7888 -539
rect 7922 -573 7980 -539
rect 8014 -573 8072 -539
rect 8106 -573 8164 -539
rect 8198 -573 8256 -539
rect 8290 -573 8348 -539
rect 8382 -573 8440 -539
rect 8474 -573 8532 -539
rect 8566 -573 8624 -539
rect 8658 -573 8716 -539
rect 8750 -573 8808 -539
rect 8842 -573 8900 -539
rect 8934 -573 8992 -539
rect 9026 -573 9084 -539
rect 9118 -573 9176 -539
rect 9210 -573 9268 -539
rect 9302 -573 9360 -539
rect 9394 -573 9452 -539
rect 9486 -573 9544 -539
rect 9578 -573 9636 -539
rect 9670 -573 9728 -539
rect 9762 -573 9820 -539
rect 9854 -573 9912 -539
rect 9946 -573 10004 -539
rect 10038 -573 10096 -539
rect 10130 -573 10188 -539
rect 10222 -573 10280 -539
rect 10314 -573 10372 -539
rect 10406 -573 10464 -539
rect 10498 -573 10556 -539
rect 10590 -573 10648 -539
rect 10682 -573 10740 -539
rect 10774 -573 10832 -539
rect 10866 -573 10924 -539
rect 10958 -573 11016 -539
rect 11050 -573 11108 -539
rect 11142 -573 11200 -539
rect 11234 -573 11292 -539
rect 11326 -573 11384 -539
rect 11418 -573 11476 -539
rect 11510 -573 11568 -539
rect 11602 -573 11660 -539
rect 11694 -573 11752 -539
rect 11786 -573 11844 -539
rect 11878 -573 11936 -539
rect 11970 -573 12028 -539
rect 12062 -573 12120 -539
rect 12154 -573 12212 -539
rect 12246 -573 12304 -539
rect 12338 -573 12396 -539
rect 12430 -573 12488 -539
rect 12522 -573 12580 -539
rect 12614 -573 12672 -539
rect 12706 -573 12764 -539
rect 12798 -573 12856 -539
rect 12890 -573 12948 -539
rect 12982 -573 13040 -539
rect 13074 -573 13132 -539
rect 13166 -573 13224 -539
rect 13258 -573 13316 -539
rect 13350 -573 13408 -539
rect 13442 -573 13500 -539
rect 13534 -573 13592 -539
rect 13626 -573 13684 -539
rect 13718 -573 13776 -539
rect 13810 -573 13868 -539
rect 13902 -573 13960 -539
rect 13994 -573 14052 -539
rect 14086 -573 14144 -539
rect 14178 -573 14236 -539
rect 14270 -573 14328 -539
rect 14362 -573 14420 -539
rect 14454 -573 14512 -539
rect 14546 -573 14604 -539
rect 14638 -573 14696 -539
rect 14730 -573 14788 -539
rect 14822 -573 14880 -539
rect 14914 -573 14972 -539
rect 15006 -573 15064 -539
rect 15098 -573 15156 -539
rect 15190 -573 15248 -539
rect 15282 -573 15340 -539
rect 15374 -573 15432 -539
rect 15466 -573 15524 -539
rect 15558 -573 15616 -539
rect 15650 -573 15708 -539
rect 15742 -573 15800 -539
rect 15834 -573 15892 -539
rect 15926 -573 15984 -539
rect 16018 -573 16076 -539
rect 16110 -573 16168 -539
rect 16202 -573 16260 -539
rect 16294 -573 16352 -539
rect 16386 -573 16444 -539
rect 16478 -573 16536 -539
rect 16570 -573 16628 -539
rect 16662 -573 16946 -539
rect -3193 -604 16946 -573
rect 13669 -681 13738 -679
rect 966 -733 982 -681
rect 1034 -682 13738 -681
rect 1034 -733 12753 -682
rect 966 -734 12753 -733
rect 12805 -734 13738 -682
rect 966 -736 13738 -734
rect 13669 -746 13738 -736
rect 1040 -770 1098 -769
rect 3000 -770 3058 -769
rect 1040 -775 3058 -770
rect 413 -854 423 -802
rect 475 -854 485 -802
rect 1040 -809 1052 -775
rect 1086 -809 3012 -775
rect 3046 -809 3058 -775
rect 1040 -814 3058 -809
rect 1040 -815 1098 -814
rect 3000 -815 3058 -814
rect 3614 -770 3672 -769
rect 5574 -770 5632 -769
rect 3614 -775 5632 -770
rect 3614 -809 3626 -775
rect 3660 -809 5586 -775
rect 5620 -809 5632 -775
rect 3614 -814 5632 -809
rect 3614 -815 3672 -814
rect 5574 -815 5632 -814
rect 6188 -770 6246 -769
rect 8148 -770 8206 -769
rect 6188 -775 8206 -770
rect 6188 -809 6200 -775
rect 6234 -809 8160 -775
rect 8194 -809 8206 -775
rect 6188 -814 8206 -809
rect 6188 -815 6246 -814
rect 8148 -815 8206 -814
rect 8762 -770 8820 -769
rect 8762 -771 10131 -770
rect 8762 -775 10783 -771
rect 8762 -809 8774 -775
rect 8808 -777 10783 -775
rect 8808 -809 10737 -777
rect 8762 -811 10737 -809
rect 10771 -811 10783 -777
rect 8762 -814 10783 -811
rect 8762 -815 8820 -814
rect 10129 -815 10783 -814
rect 10725 -817 10783 -815
rect 11338 -778 11430 -771
rect 11338 -812 11369 -778
rect 11403 -812 11430 -778
rect 11338 -828 11430 -812
rect 13669 -780 13685 -746
rect 13719 -780 13738 -746
rect 13669 -823 13738 -780
rect 15236 -728 15294 -722
rect 15328 -728 15386 -723
rect 15236 -762 15248 -728
rect 15282 -729 15394 -728
rect 15282 -762 15340 -729
rect 15236 -763 15340 -762
rect 15374 -763 15394 -729
rect 15236 -808 15394 -763
rect 15236 -824 16946 -808
rect 11338 -883 12463 -828
rect 11339 -887 12463 -883
rect 12522 -887 12532 -828
rect 15236 -858 15248 -824
rect 15282 -858 15341 -824
rect 15375 -848 16946 -824
rect 15375 -858 15394 -848
rect 15236 -864 15294 -858
rect 15329 -864 15387 -858
rect -3193 -1083 16946 -1052
rect -3193 -1117 -2968 -1083
rect -2934 -1117 -2876 -1083
rect -2842 -1117 -2784 -1083
rect -2750 -1117 -2692 -1083
rect -2658 -1117 -2600 -1083
rect -2566 -1117 -2508 -1083
rect -2474 -1117 -2416 -1083
rect -2382 -1117 -2324 -1083
rect -2290 -1117 -2232 -1083
rect -2198 -1117 -2140 -1083
rect -2106 -1117 -2048 -1083
rect -2014 -1117 -1956 -1083
rect -1922 -1117 -1864 -1083
rect -1830 -1117 -1772 -1083
rect -1738 -1117 -1680 -1083
rect -1646 -1117 -1588 -1083
rect -1554 -1117 -1496 -1083
rect -1462 -1117 -1404 -1083
rect -1370 -1117 -1312 -1083
rect -1278 -1117 -1220 -1083
rect -1186 -1117 -1128 -1083
rect -1094 -1117 -1036 -1083
rect -1002 -1117 -944 -1083
rect -910 -1117 -852 -1083
rect -818 -1117 -760 -1083
rect -726 -1117 -668 -1083
rect -634 -1117 -576 -1083
rect -542 -1117 -484 -1083
rect -450 -1117 -392 -1083
rect -358 -1117 -300 -1083
rect -266 -1117 -208 -1083
rect -174 -1117 -116 -1083
rect -82 -1117 -24 -1083
rect 10 -1117 68 -1083
rect 102 -1117 160 -1083
rect 194 -1117 252 -1083
rect 286 -1117 344 -1083
rect 378 -1117 436 -1083
rect 470 -1117 528 -1083
rect 562 -1117 620 -1083
rect 654 -1117 712 -1083
rect 746 -1117 804 -1083
rect 838 -1117 896 -1083
rect 930 -1117 988 -1083
rect 1022 -1117 1080 -1083
rect 1114 -1117 1172 -1083
rect 1206 -1117 1264 -1083
rect 1298 -1117 1356 -1083
rect 1390 -1117 1448 -1083
rect 1482 -1117 1540 -1083
rect 1574 -1117 1632 -1083
rect 1666 -1117 1724 -1083
rect 1758 -1117 1816 -1083
rect 1850 -1117 1908 -1083
rect 1942 -1117 2000 -1083
rect 2034 -1117 2092 -1083
rect 2126 -1117 2184 -1083
rect 2218 -1117 2276 -1083
rect 2310 -1117 2368 -1083
rect 2402 -1117 2460 -1083
rect 2494 -1117 2552 -1083
rect 2586 -1117 2644 -1083
rect 2678 -1117 2736 -1083
rect 2770 -1117 2828 -1083
rect 2862 -1117 2920 -1083
rect 2954 -1117 3012 -1083
rect 3046 -1117 3104 -1083
rect 3138 -1117 3196 -1083
rect 3230 -1117 3288 -1083
rect 3322 -1117 3380 -1083
rect 3414 -1117 3472 -1083
rect 3506 -1117 3564 -1083
rect 3598 -1117 3656 -1083
rect 3690 -1117 3748 -1083
rect 3782 -1117 3840 -1083
rect 3874 -1117 3932 -1083
rect 3966 -1117 4024 -1083
rect 4058 -1117 4116 -1083
rect 4150 -1117 4208 -1083
rect 4242 -1117 4300 -1083
rect 4334 -1117 4392 -1083
rect 4426 -1117 4484 -1083
rect 4518 -1117 4576 -1083
rect 4610 -1117 4668 -1083
rect 4702 -1117 4760 -1083
rect 4794 -1117 4852 -1083
rect 4886 -1117 4944 -1083
rect 4978 -1117 5036 -1083
rect 5070 -1117 5128 -1083
rect 5162 -1117 5220 -1083
rect 5254 -1117 5312 -1083
rect 5346 -1117 5404 -1083
rect 5438 -1117 5496 -1083
rect 5530 -1117 5588 -1083
rect 5622 -1117 5680 -1083
rect 5714 -1117 5772 -1083
rect 5806 -1117 5864 -1083
rect 5898 -1117 5956 -1083
rect 5990 -1117 6048 -1083
rect 6082 -1117 6140 -1083
rect 6174 -1117 6232 -1083
rect 6266 -1117 6324 -1083
rect 6358 -1117 6416 -1083
rect 6450 -1117 6508 -1083
rect 6542 -1117 6600 -1083
rect 6634 -1117 6692 -1083
rect 6726 -1117 6784 -1083
rect 6818 -1117 6876 -1083
rect 6910 -1117 6968 -1083
rect 7002 -1117 7060 -1083
rect 7094 -1117 7152 -1083
rect 7186 -1117 7244 -1083
rect 7278 -1117 7336 -1083
rect 7370 -1117 7428 -1083
rect 7462 -1117 7520 -1083
rect 7554 -1117 7612 -1083
rect 7646 -1117 7704 -1083
rect 7738 -1117 7796 -1083
rect 7830 -1117 7888 -1083
rect 7922 -1117 7980 -1083
rect 8014 -1117 8072 -1083
rect 8106 -1117 8164 -1083
rect 8198 -1117 8256 -1083
rect 8290 -1117 8348 -1083
rect 8382 -1117 8440 -1083
rect 8474 -1117 8532 -1083
rect 8566 -1117 8624 -1083
rect 8658 -1117 8716 -1083
rect 8750 -1117 8808 -1083
rect 8842 -1117 8900 -1083
rect 8934 -1117 8992 -1083
rect 9026 -1117 9084 -1083
rect 9118 -1117 9176 -1083
rect 9210 -1117 9268 -1083
rect 9302 -1117 9360 -1083
rect 9394 -1117 9452 -1083
rect 9486 -1117 9544 -1083
rect 9578 -1117 9636 -1083
rect 9670 -1117 9728 -1083
rect 9762 -1117 9820 -1083
rect 9854 -1117 9912 -1083
rect 9946 -1117 10004 -1083
rect 10038 -1117 10096 -1083
rect 10130 -1117 10188 -1083
rect 10222 -1117 10280 -1083
rect 10314 -1117 10372 -1083
rect 10406 -1117 10464 -1083
rect 10498 -1117 10556 -1083
rect 10590 -1117 10648 -1083
rect 10682 -1117 10740 -1083
rect 10774 -1117 10832 -1083
rect 10866 -1117 10924 -1083
rect 10958 -1117 11016 -1083
rect 11050 -1117 11108 -1083
rect 11142 -1117 11200 -1083
rect 11234 -1117 11292 -1083
rect 11326 -1117 11384 -1083
rect 11418 -1117 11476 -1083
rect 11510 -1117 11568 -1083
rect 11602 -1117 11660 -1083
rect 11694 -1117 11752 -1083
rect 11786 -1117 11844 -1083
rect 11878 -1117 11936 -1083
rect 11970 -1117 12028 -1083
rect 12062 -1117 12120 -1083
rect 12154 -1117 12212 -1083
rect 12246 -1117 12304 -1083
rect 12338 -1117 12396 -1083
rect 12430 -1117 12488 -1083
rect 12522 -1117 12580 -1083
rect 12614 -1117 12672 -1083
rect 12706 -1117 12764 -1083
rect 12798 -1117 12856 -1083
rect 12890 -1117 12948 -1083
rect 12982 -1117 13040 -1083
rect 13074 -1117 13132 -1083
rect 13166 -1117 13224 -1083
rect 13258 -1117 13316 -1083
rect 13350 -1117 13408 -1083
rect 13442 -1117 13500 -1083
rect 13534 -1117 13592 -1083
rect 13626 -1117 13684 -1083
rect 13718 -1117 13776 -1083
rect 13810 -1117 13868 -1083
rect 13902 -1117 13960 -1083
rect 13994 -1117 14052 -1083
rect 14086 -1117 14144 -1083
rect 14178 -1117 14236 -1083
rect 14270 -1117 14328 -1083
rect 14362 -1117 14420 -1083
rect 14454 -1117 14512 -1083
rect 14546 -1117 14604 -1083
rect 14638 -1117 14696 -1083
rect 14730 -1117 14788 -1083
rect 14822 -1117 14880 -1083
rect 14914 -1117 14972 -1083
rect 15006 -1117 15064 -1083
rect 15098 -1117 15156 -1083
rect 15190 -1117 15248 -1083
rect 15282 -1117 15340 -1083
rect 15374 -1117 15432 -1083
rect 15466 -1117 15524 -1083
rect 15558 -1117 15616 -1083
rect 15650 -1117 15708 -1083
rect 15742 -1117 15800 -1083
rect 15834 -1117 15892 -1083
rect 15926 -1117 15984 -1083
rect 16018 -1117 16076 -1083
rect 16110 -1117 16168 -1083
rect 16202 -1117 16260 -1083
rect 16294 -1117 16352 -1083
rect 16386 -1117 16444 -1083
rect 16478 -1117 16536 -1083
rect 16570 -1117 16628 -1083
rect 16662 -1117 16946 -1083
rect -3193 -1148 16946 -1117
rect 7161 -1232 11181 -1231
rect 7161 -1235 11118 -1232
rect 7155 -1287 7165 -1235
rect 7217 -1284 11118 -1235
rect 11170 -1284 11181 -1232
rect 7217 -1287 11181 -1284
rect 7161 -1293 11181 -1287
rect 15236 -1338 15294 -1332
rect 15328 -1338 15386 -1333
rect 413 -1435 423 -1383
rect 475 -1435 485 -1383
rect 1070 -1384 1128 -1383
rect 3030 -1384 3088 -1383
rect 1070 -1389 3088 -1384
rect 1070 -1423 1082 -1389
rect 1116 -1423 3042 -1389
rect 3076 -1423 3088 -1389
rect 1070 -1428 3088 -1423
rect 1070 -1429 1128 -1428
rect 3030 -1429 3088 -1428
rect 3644 -1384 3702 -1383
rect 5604 -1384 5662 -1383
rect 3644 -1389 5662 -1384
rect 3644 -1423 3656 -1389
rect 3690 -1423 5616 -1389
rect 5650 -1423 5662 -1389
rect 3644 -1428 5662 -1423
rect 3644 -1429 3702 -1428
rect 5604 -1429 5662 -1428
rect 6218 -1384 6276 -1383
rect 8178 -1384 8236 -1383
rect 6218 -1389 8236 -1384
rect 6218 -1423 6230 -1389
rect 6264 -1423 8190 -1389
rect 8224 -1423 8236 -1389
rect 6218 -1428 8236 -1423
rect 6218 -1429 6276 -1428
rect 8178 -1429 8236 -1428
rect 8792 -1384 8850 -1383
rect 10752 -1384 10810 -1383
rect 8792 -1389 10810 -1384
rect 8792 -1423 8804 -1389
rect 8838 -1423 10764 -1389
rect 10798 -1423 10810 -1389
rect 11368 -1397 11378 -1345
rect 11430 -1397 11440 -1345
rect 15236 -1372 15248 -1338
rect 15282 -1339 15394 -1338
rect 15282 -1372 15340 -1339
rect 15236 -1373 15340 -1372
rect 15374 -1352 15394 -1339
rect 15374 -1373 16946 -1352
rect 13026 -1380 13084 -1379
rect 12548 -1386 12752 -1382
rect 12546 -1392 12752 -1386
rect 12804 -1392 12992 -1382
rect 8792 -1428 10810 -1423
rect 8792 -1429 8850 -1428
rect 10752 -1429 10810 -1428
rect 12546 -1426 12558 -1392
rect 12592 -1426 12642 -1392
rect 12676 -1426 12739 -1392
rect 12804 -1426 12836 -1392
rect 12870 -1426 12942 -1392
rect 12976 -1426 12992 -1392
rect 12546 -1432 12752 -1426
rect 12548 -1434 12752 -1432
rect 12804 -1434 12992 -1426
rect 12548 -1435 12992 -1434
rect 13026 -1385 13737 -1380
rect 13026 -1419 13038 -1385
rect 13072 -1419 13737 -1385
rect 13026 -1422 13737 -1419
rect 13026 -1456 13684 -1422
rect 13718 -1456 13737 -1422
rect 13026 -1457 13737 -1456
rect 13026 -1491 13038 -1457
rect 13072 -1490 13737 -1457
rect 15236 -1392 16946 -1373
rect 15236 -1434 15394 -1392
rect 15236 -1468 15248 -1434
rect 15282 -1468 15341 -1434
rect 15375 -1468 15394 -1434
rect 15236 -1474 15294 -1468
rect 15329 -1474 15387 -1468
rect 13072 -1491 13084 -1490
rect 13026 -1498 13084 -1491
rect -3193 -1627 16946 -1596
rect -3193 -1661 -2968 -1627
rect -2934 -1661 -2876 -1627
rect -2842 -1661 -2784 -1627
rect -2750 -1661 -2692 -1627
rect -2658 -1661 -2600 -1627
rect -2566 -1661 -2508 -1627
rect -2474 -1661 -2416 -1627
rect -2382 -1661 -2324 -1627
rect -2290 -1661 -2232 -1627
rect -2198 -1661 -2140 -1627
rect -2106 -1661 -2048 -1627
rect -2014 -1661 -1956 -1627
rect -1922 -1661 -1864 -1627
rect -1830 -1661 -1772 -1627
rect -1738 -1661 -1680 -1627
rect -1646 -1661 -1588 -1627
rect -1554 -1661 -1496 -1627
rect -1462 -1661 -1404 -1627
rect -1370 -1661 -1312 -1627
rect -1278 -1661 -1220 -1627
rect -1186 -1661 -1128 -1627
rect -1094 -1661 -1036 -1627
rect -1002 -1661 -944 -1627
rect -910 -1661 -852 -1627
rect -818 -1661 -760 -1627
rect -726 -1661 -668 -1627
rect -634 -1661 -576 -1627
rect -542 -1661 -484 -1627
rect -450 -1661 -392 -1627
rect -358 -1661 -300 -1627
rect -266 -1661 -208 -1627
rect -174 -1661 -116 -1627
rect -82 -1661 -24 -1627
rect 10 -1661 68 -1627
rect 102 -1661 160 -1627
rect 194 -1661 252 -1627
rect 286 -1661 344 -1627
rect 378 -1661 436 -1627
rect 470 -1661 528 -1627
rect 562 -1661 620 -1627
rect 654 -1661 712 -1627
rect 746 -1661 804 -1627
rect 838 -1661 896 -1627
rect 930 -1661 988 -1627
rect 1022 -1661 1080 -1627
rect 1114 -1661 1172 -1627
rect 1206 -1661 1264 -1627
rect 1298 -1661 1356 -1627
rect 1390 -1661 1448 -1627
rect 1482 -1661 1540 -1627
rect 1574 -1661 1632 -1627
rect 1666 -1661 1724 -1627
rect 1758 -1661 1816 -1627
rect 1850 -1661 1908 -1627
rect 1942 -1661 2000 -1627
rect 2034 -1661 2092 -1627
rect 2126 -1661 2184 -1627
rect 2218 -1661 2276 -1627
rect 2310 -1661 2368 -1627
rect 2402 -1661 2460 -1627
rect 2494 -1661 2552 -1627
rect 2586 -1661 2644 -1627
rect 2678 -1661 2736 -1627
rect 2770 -1661 2828 -1627
rect 2862 -1661 2920 -1627
rect 2954 -1661 3012 -1627
rect 3046 -1661 3104 -1627
rect 3138 -1661 3196 -1627
rect 3230 -1661 3288 -1627
rect 3322 -1661 3380 -1627
rect 3414 -1661 3472 -1627
rect 3506 -1661 3564 -1627
rect 3598 -1661 3656 -1627
rect 3690 -1661 3748 -1627
rect 3782 -1661 3840 -1627
rect 3874 -1661 3932 -1627
rect 3966 -1661 4024 -1627
rect 4058 -1661 4116 -1627
rect 4150 -1661 4208 -1627
rect 4242 -1661 4300 -1627
rect 4334 -1661 4392 -1627
rect 4426 -1661 4484 -1627
rect 4518 -1661 4576 -1627
rect 4610 -1661 4668 -1627
rect 4702 -1661 4760 -1627
rect 4794 -1661 4852 -1627
rect 4886 -1661 4944 -1627
rect 4978 -1661 5036 -1627
rect 5070 -1661 5128 -1627
rect 5162 -1661 5220 -1627
rect 5254 -1661 5312 -1627
rect 5346 -1661 5404 -1627
rect 5438 -1661 5496 -1627
rect 5530 -1661 5588 -1627
rect 5622 -1661 5680 -1627
rect 5714 -1661 5772 -1627
rect 5806 -1661 5864 -1627
rect 5898 -1661 5956 -1627
rect 5990 -1661 6048 -1627
rect 6082 -1661 6140 -1627
rect 6174 -1661 6232 -1627
rect 6266 -1661 6324 -1627
rect 6358 -1661 6416 -1627
rect 6450 -1661 6508 -1627
rect 6542 -1661 6600 -1627
rect 6634 -1661 6692 -1627
rect 6726 -1661 6784 -1627
rect 6818 -1661 6876 -1627
rect 6910 -1661 6968 -1627
rect 7002 -1661 7060 -1627
rect 7094 -1661 7152 -1627
rect 7186 -1661 7244 -1627
rect 7278 -1661 7336 -1627
rect 7370 -1661 7428 -1627
rect 7462 -1661 7520 -1627
rect 7554 -1661 7612 -1627
rect 7646 -1661 7704 -1627
rect 7738 -1661 7796 -1627
rect 7830 -1661 7888 -1627
rect 7922 -1661 7980 -1627
rect 8014 -1661 8072 -1627
rect 8106 -1661 8164 -1627
rect 8198 -1661 8256 -1627
rect 8290 -1661 8348 -1627
rect 8382 -1661 8440 -1627
rect 8474 -1661 8532 -1627
rect 8566 -1661 8624 -1627
rect 8658 -1661 8716 -1627
rect 8750 -1661 8808 -1627
rect 8842 -1661 8900 -1627
rect 8934 -1661 8992 -1627
rect 9026 -1661 9084 -1627
rect 9118 -1661 9176 -1627
rect 9210 -1661 9268 -1627
rect 9302 -1661 9360 -1627
rect 9394 -1661 9452 -1627
rect 9486 -1661 9544 -1627
rect 9578 -1661 9636 -1627
rect 9670 -1661 9728 -1627
rect 9762 -1661 9820 -1627
rect 9854 -1661 9912 -1627
rect 9946 -1661 10004 -1627
rect 10038 -1661 10096 -1627
rect 10130 -1661 10188 -1627
rect 10222 -1661 10280 -1627
rect 10314 -1661 10372 -1627
rect 10406 -1661 10464 -1627
rect 10498 -1661 10556 -1627
rect 10590 -1661 10648 -1627
rect 10682 -1661 10740 -1627
rect 10774 -1661 10832 -1627
rect 10866 -1661 10924 -1627
rect 10958 -1661 11016 -1627
rect 11050 -1661 11108 -1627
rect 11142 -1661 11200 -1627
rect 11234 -1661 11292 -1627
rect 11326 -1661 11384 -1627
rect 11418 -1661 11476 -1627
rect 11510 -1661 11568 -1627
rect 11602 -1661 11660 -1627
rect 11694 -1661 11752 -1627
rect 11786 -1661 11844 -1627
rect 11878 -1661 11936 -1627
rect 11970 -1661 12028 -1627
rect 12062 -1661 12120 -1627
rect 12154 -1661 12212 -1627
rect 12246 -1661 12304 -1627
rect 12338 -1661 12396 -1627
rect 12430 -1661 12488 -1627
rect 12522 -1661 12580 -1627
rect 12614 -1661 12672 -1627
rect 12706 -1661 12764 -1627
rect 12798 -1661 12856 -1627
rect 12890 -1661 12948 -1627
rect 12982 -1661 13040 -1627
rect 13074 -1661 13132 -1627
rect 13166 -1661 13224 -1627
rect 13258 -1661 13316 -1627
rect 13350 -1661 13408 -1627
rect 13442 -1661 13500 -1627
rect 13534 -1661 13592 -1627
rect 13626 -1661 13684 -1627
rect 13718 -1661 13776 -1627
rect 13810 -1661 13868 -1627
rect 13902 -1661 13960 -1627
rect 13994 -1661 14052 -1627
rect 14086 -1661 14144 -1627
rect 14178 -1661 14236 -1627
rect 14270 -1661 14328 -1627
rect 14362 -1661 14420 -1627
rect 14454 -1661 14512 -1627
rect 14546 -1661 14604 -1627
rect 14638 -1661 14696 -1627
rect 14730 -1661 14788 -1627
rect 14822 -1661 14880 -1627
rect 14914 -1661 14972 -1627
rect 15006 -1661 15064 -1627
rect 15098 -1661 15156 -1627
rect 15190 -1661 15248 -1627
rect 15282 -1661 15340 -1627
rect 15374 -1661 15432 -1627
rect 15466 -1661 15524 -1627
rect 15558 -1661 15616 -1627
rect 15650 -1661 15708 -1627
rect 15742 -1661 15800 -1627
rect 15834 -1661 15892 -1627
rect 15926 -1661 15984 -1627
rect 16018 -1661 16076 -1627
rect 16110 -1661 16168 -1627
rect 16202 -1661 16260 -1627
rect 16294 -1661 16352 -1627
rect 16386 -1661 16444 -1627
rect 16478 -1661 16536 -1627
rect 16570 -1661 16628 -1627
rect 16662 -1661 16946 -1627
rect -3193 -1692 16946 -1661
rect 13671 -1762 13735 -1761
rect 7153 -1763 13735 -1762
rect 7153 -1815 7163 -1763
rect 7215 -1766 13735 -1763
rect 7215 -1815 12756 -1766
rect 7153 -1816 12756 -1815
rect 12746 -1818 12756 -1816
rect 12808 -1816 13735 -1766
rect 12808 -1818 12818 -1816
rect 13671 -1832 13735 -1816
rect -952 -1943 -942 -1891
rect -890 -1893 -880 -1891
rect -890 -1900 -809 -1893
rect -890 -1934 -856 -1900
rect -822 -1934 -809 -1900
rect -227 -1906 -217 -1854
rect -165 -1906 -155 -1854
rect 1042 -1861 1100 -1860
rect 3002 -1861 3060 -1860
rect 1042 -1866 3060 -1861
rect -890 -1941 -809 -1934
rect -890 -1943 -880 -1941
rect 413 -1942 423 -1890
rect 475 -1942 485 -1890
rect 1042 -1900 1054 -1866
rect 1088 -1900 3014 -1866
rect 3048 -1900 3060 -1866
rect 1042 -1905 3060 -1900
rect 1042 -1906 1100 -1905
rect 3002 -1906 3060 -1905
rect 3616 -1861 3674 -1860
rect 5576 -1861 5634 -1860
rect 3616 -1866 5634 -1861
rect 3616 -1900 3628 -1866
rect 3662 -1900 5588 -1866
rect 5622 -1900 5634 -1866
rect 3616 -1905 5634 -1900
rect 3616 -1906 3674 -1905
rect 5576 -1906 5634 -1905
rect 6190 -1861 6248 -1860
rect 8150 -1861 8208 -1860
rect 6190 -1866 8208 -1861
rect 6190 -1900 6202 -1866
rect 6236 -1900 8162 -1866
rect 8196 -1900 8208 -1866
rect 6190 -1905 8208 -1900
rect 6190 -1906 6248 -1905
rect 8150 -1906 8208 -1905
rect 8764 -1861 8822 -1860
rect 10724 -1861 10782 -1860
rect 8764 -1866 10782 -1861
rect 8764 -1900 8776 -1866
rect 8810 -1900 10736 -1866
rect 10770 -1900 10782 -1866
rect 8764 -1905 10782 -1900
rect 8764 -1906 8822 -1905
rect 10724 -1906 10782 -1905
rect 11365 -1908 11375 -1856
rect 11427 -1908 11437 -1856
rect 13671 -1866 13685 -1832
rect 13719 -1866 13735 -1832
rect 13671 -1910 13735 -1866
rect 15236 -1816 15294 -1810
rect 15328 -1816 15386 -1811
rect 15236 -1850 15248 -1816
rect 15282 -1817 15394 -1816
rect 15282 -1850 15340 -1817
rect 15236 -1851 15340 -1850
rect 15374 -1851 15394 -1817
rect 15236 -1896 15394 -1851
rect 15236 -1912 16946 -1896
rect 15236 -1946 15248 -1912
rect 15282 -1946 15341 -1912
rect 15375 -1936 16946 -1912
rect 15375 -1946 15394 -1936
rect 15236 -1952 15294 -1946
rect 15329 -1952 15387 -1946
rect -3193 -2171 16946 -2140
rect -3193 -2205 -2968 -2171
rect -2934 -2205 -2876 -2171
rect -2842 -2205 -2784 -2171
rect -2750 -2205 -2692 -2171
rect -2658 -2205 -2600 -2171
rect -2566 -2205 -2508 -2171
rect -2474 -2205 -2416 -2171
rect -2382 -2205 -2324 -2171
rect -2290 -2205 -2232 -2171
rect -2198 -2205 -2140 -2171
rect -2106 -2205 -2048 -2171
rect -2014 -2205 -1956 -2171
rect -1922 -2205 -1864 -2171
rect -1830 -2205 -1772 -2171
rect -1738 -2205 -1680 -2171
rect -1646 -2205 -1588 -2171
rect -1554 -2205 -1496 -2171
rect -1462 -2205 -1404 -2171
rect -1370 -2205 -1312 -2171
rect -1278 -2205 -1220 -2171
rect -1186 -2205 -1128 -2171
rect -1094 -2205 -1036 -2171
rect -1002 -2205 -944 -2171
rect -910 -2205 -852 -2171
rect -818 -2205 -760 -2171
rect -726 -2205 -668 -2171
rect -634 -2205 -576 -2171
rect -542 -2205 -484 -2171
rect -450 -2205 -392 -2171
rect -358 -2205 -300 -2171
rect -266 -2205 -208 -2171
rect -174 -2205 -116 -2171
rect -82 -2205 -24 -2171
rect 10 -2205 68 -2171
rect 102 -2205 160 -2171
rect 194 -2205 252 -2171
rect 286 -2205 344 -2171
rect 378 -2205 436 -2171
rect 470 -2205 528 -2171
rect 562 -2205 620 -2171
rect 654 -2205 712 -2171
rect 746 -2205 804 -2171
rect 838 -2205 896 -2171
rect 930 -2205 988 -2171
rect 1022 -2205 1080 -2171
rect 1114 -2205 1172 -2171
rect 1206 -2205 1264 -2171
rect 1298 -2205 1356 -2171
rect 1390 -2205 1448 -2171
rect 1482 -2205 1540 -2171
rect 1574 -2205 1632 -2171
rect 1666 -2205 1724 -2171
rect 1758 -2205 1816 -2171
rect 1850 -2205 1908 -2171
rect 1942 -2205 2000 -2171
rect 2034 -2205 2092 -2171
rect 2126 -2205 2184 -2171
rect 2218 -2205 2276 -2171
rect 2310 -2205 2368 -2171
rect 2402 -2205 2460 -2171
rect 2494 -2205 2552 -2171
rect 2586 -2205 2644 -2171
rect 2678 -2205 2736 -2171
rect 2770 -2205 2828 -2171
rect 2862 -2205 2920 -2171
rect 2954 -2205 3012 -2171
rect 3046 -2205 3104 -2171
rect 3138 -2205 3196 -2171
rect 3230 -2205 3288 -2171
rect 3322 -2205 3380 -2171
rect 3414 -2205 3472 -2171
rect 3506 -2205 3564 -2171
rect 3598 -2205 3656 -2171
rect 3690 -2205 3748 -2171
rect 3782 -2205 3840 -2171
rect 3874 -2205 3932 -2171
rect 3966 -2205 4024 -2171
rect 4058 -2205 4116 -2171
rect 4150 -2205 4208 -2171
rect 4242 -2205 4300 -2171
rect 4334 -2205 4392 -2171
rect 4426 -2205 4484 -2171
rect 4518 -2205 4576 -2171
rect 4610 -2205 4668 -2171
rect 4702 -2205 4760 -2171
rect 4794 -2205 4852 -2171
rect 4886 -2205 4944 -2171
rect 4978 -2205 5036 -2171
rect 5070 -2205 5128 -2171
rect 5162 -2205 5220 -2171
rect 5254 -2205 5312 -2171
rect 5346 -2205 5404 -2171
rect 5438 -2205 5496 -2171
rect 5530 -2205 5588 -2171
rect 5622 -2205 5680 -2171
rect 5714 -2205 5772 -2171
rect 5806 -2205 5864 -2171
rect 5898 -2205 5956 -2171
rect 5990 -2205 6048 -2171
rect 6082 -2205 6140 -2171
rect 6174 -2205 6232 -2171
rect 6266 -2205 6324 -2171
rect 6358 -2205 6416 -2171
rect 6450 -2205 6508 -2171
rect 6542 -2205 6600 -2171
rect 6634 -2205 6692 -2171
rect 6726 -2205 6784 -2171
rect 6818 -2205 6876 -2171
rect 6910 -2205 6968 -2171
rect 7002 -2205 7060 -2171
rect 7094 -2205 7152 -2171
rect 7186 -2205 7244 -2171
rect 7278 -2205 7336 -2171
rect 7370 -2205 7428 -2171
rect 7462 -2205 7520 -2171
rect 7554 -2205 7612 -2171
rect 7646 -2205 7704 -2171
rect 7738 -2205 7796 -2171
rect 7830 -2205 7888 -2171
rect 7922 -2205 7980 -2171
rect 8014 -2205 8072 -2171
rect 8106 -2205 8164 -2171
rect 8198 -2205 8256 -2171
rect 8290 -2205 8348 -2171
rect 8382 -2205 8440 -2171
rect 8474 -2205 8532 -2171
rect 8566 -2205 8624 -2171
rect 8658 -2205 8716 -2171
rect 8750 -2205 8808 -2171
rect 8842 -2205 8900 -2171
rect 8934 -2205 8992 -2171
rect 9026 -2205 9084 -2171
rect 9118 -2205 9176 -2171
rect 9210 -2205 9268 -2171
rect 9302 -2205 9360 -2171
rect 9394 -2205 9452 -2171
rect 9486 -2205 9544 -2171
rect 9578 -2205 9636 -2171
rect 9670 -2205 9728 -2171
rect 9762 -2205 9820 -2171
rect 9854 -2205 9912 -2171
rect 9946 -2205 10004 -2171
rect 10038 -2205 10096 -2171
rect 10130 -2205 10188 -2171
rect 10222 -2205 10280 -2171
rect 10314 -2205 10372 -2171
rect 10406 -2205 10464 -2171
rect 10498 -2205 10556 -2171
rect 10590 -2205 10648 -2171
rect 10682 -2205 10740 -2171
rect 10774 -2205 10832 -2171
rect 10866 -2205 10924 -2171
rect 10958 -2205 11016 -2171
rect 11050 -2205 11108 -2171
rect 11142 -2205 11200 -2171
rect 11234 -2205 11292 -2171
rect 11326 -2205 11384 -2171
rect 11418 -2205 11476 -2171
rect 11510 -2205 11568 -2171
rect 11602 -2205 11660 -2171
rect 11694 -2205 11752 -2171
rect 11786 -2205 11844 -2171
rect 11878 -2205 11936 -2171
rect 11970 -2205 12028 -2171
rect 12062 -2205 12120 -2171
rect 12154 -2205 12212 -2171
rect 12246 -2205 12304 -2171
rect 12338 -2205 12396 -2171
rect 12430 -2205 12488 -2171
rect 12522 -2205 12580 -2171
rect 12614 -2205 12672 -2171
rect 12706 -2205 12764 -2171
rect 12798 -2205 12856 -2171
rect 12890 -2205 12948 -2171
rect 12982 -2205 13040 -2171
rect 13074 -2205 13132 -2171
rect 13166 -2205 13224 -2171
rect 13258 -2205 13316 -2171
rect 13350 -2205 13408 -2171
rect 13442 -2205 13500 -2171
rect 13534 -2205 13592 -2171
rect 13626 -2205 13684 -2171
rect 13718 -2205 13776 -2171
rect 13810 -2205 13868 -2171
rect 13902 -2205 13960 -2171
rect 13994 -2205 14052 -2171
rect 14086 -2205 14144 -2171
rect 14178 -2205 14236 -2171
rect 14270 -2205 14328 -2171
rect 14362 -2205 14420 -2171
rect 14454 -2205 14512 -2171
rect 14546 -2205 14604 -2171
rect 14638 -2205 14696 -2171
rect 14730 -2205 14788 -2171
rect 14822 -2205 14880 -2171
rect 14914 -2205 14972 -2171
rect 15006 -2205 15064 -2171
rect 15098 -2205 15156 -2171
rect 15190 -2205 15248 -2171
rect 15282 -2205 15340 -2171
rect 15374 -2205 15432 -2171
rect 15466 -2205 15524 -2171
rect 15558 -2205 15616 -2171
rect 15650 -2205 15708 -2171
rect 15742 -2205 15800 -2171
rect 15834 -2205 15892 -2171
rect 15926 -2205 15984 -2171
rect 16018 -2205 16076 -2171
rect 16110 -2205 16168 -2171
rect 16202 -2205 16260 -2171
rect 16294 -2205 16352 -2171
rect 16386 -2205 16444 -2171
rect 16478 -2205 16536 -2171
rect 16570 -2205 16628 -2171
rect 16662 -2205 16946 -2171
rect -3193 -2236 16946 -2205
rect 12467 -2407 12520 -2375
rect 12467 -2414 12480 -2407
rect 12514 -2414 12520 -2407
rect 418 -2521 428 -2469
rect 480 -2521 490 -2469
rect 1069 -2473 1127 -2472
rect 3029 -2473 3087 -2472
rect 1069 -2478 3087 -2473
rect 1069 -2512 1081 -2478
rect 1115 -2512 3041 -2478
rect 3075 -2512 3087 -2478
rect 1069 -2517 3087 -2512
rect 1069 -2518 1127 -2517
rect 3029 -2518 3087 -2517
rect 3643 -2473 3701 -2472
rect 5603 -2473 5661 -2472
rect 3643 -2478 5661 -2473
rect 3643 -2512 3655 -2478
rect 3689 -2512 5615 -2478
rect 5649 -2512 5661 -2478
rect 3643 -2517 5661 -2512
rect 3643 -2518 3701 -2517
rect 5603 -2518 5661 -2517
rect 6217 -2473 6275 -2472
rect 8177 -2473 8235 -2472
rect 6217 -2478 8235 -2473
rect 6217 -2512 6229 -2478
rect 6263 -2512 8189 -2478
rect 8223 -2512 8235 -2478
rect 6217 -2517 8235 -2512
rect 6217 -2518 6275 -2517
rect 8177 -2518 8235 -2517
rect 8791 -2473 8849 -2472
rect 10751 -2473 10809 -2472
rect 8791 -2478 10809 -2473
rect 8791 -2512 8806 -2478
rect 8840 -2512 10763 -2478
rect 10797 -2512 10809 -2478
rect 11368 -2488 11378 -2436
rect 11430 -2488 11440 -2436
rect 12456 -2466 12466 -2414
rect 12518 -2466 12520 -2414
rect 15236 -2426 15294 -2420
rect 15328 -2426 15386 -2420
rect 13027 -2461 13085 -2460
rect 12467 -2481 12520 -2466
rect 13023 -2466 13738 -2461
rect 12846 -2472 12991 -2471
rect 8791 -2517 10809 -2512
rect 8791 -2518 8849 -2517
rect 10751 -2518 10809 -2517
rect 12467 -2515 12480 -2481
rect 12514 -2515 12520 -2481
rect 12467 -2528 12520 -2515
rect 12548 -2479 12755 -2472
rect 12807 -2477 12993 -2472
rect 12548 -2513 12568 -2479
rect 12602 -2513 12659 -2479
rect 12693 -2513 12755 -2479
rect 12807 -2511 12858 -2477
rect 12892 -2511 12942 -2477
rect 12976 -2511 12993 -2477
rect 12548 -2521 12755 -2513
rect 12745 -2524 12755 -2521
rect 12807 -2521 12993 -2511
rect 13023 -2500 13039 -2466
rect 13073 -2500 13738 -2466
rect 13916 -2485 13926 -2433
rect 13978 -2440 13988 -2433
rect 15236 -2440 15248 -2426
rect 13978 -2460 15248 -2440
rect 15282 -2460 15340 -2426
rect 15374 -2440 15394 -2426
rect 15374 -2460 16946 -2440
rect 13978 -2480 16946 -2460
rect 13978 -2485 13988 -2480
rect 13023 -2510 13738 -2500
rect 12807 -2524 12817 -2521
rect 12456 -2580 12466 -2528
rect 12518 -2580 12520 -2528
rect 12467 -2587 12480 -2580
rect 12514 -2587 12520 -2580
rect 13023 -2543 13685 -2510
rect 13023 -2577 13042 -2543
rect 13076 -2544 13685 -2543
rect 13719 -2544 13738 -2510
rect 13076 -2577 13738 -2544
rect 15236 -2522 15394 -2480
rect 15236 -2556 15248 -2522
rect 15282 -2556 15341 -2522
rect 15375 -2556 15394 -2522
rect 15236 -2562 15294 -2556
rect 15329 -2562 15387 -2556
rect 13023 -2584 13738 -2577
rect 12467 -2612 12520 -2587
rect -3193 -2715 16946 -2684
rect -3193 -2749 -2968 -2715
rect -2934 -2749 -2876 -2715
rect -2842 -2749 -2784 -2715
rect -2750 -2749 -2692 -2715
rect -2658 -2749 -2600 -2715
rect -2566 -2749 -2508 -2715
rect -2474 -2749 -2416 -2715
rect -2382 -2749 -2324 -2715
rect -2290 -2749 -2232 -2715
rect -2198 -2749 -2140 -2715
rect -2106 -2749 -2048 -2715
rect -2014 -2749 -1956 -2715
rect -1922 -2749 -1864 -2715
rect -1830 -2749 -1772 -2715
rect -1738 -2749 -1680 -2715
rect -1646 -2749 -1588 -2715
rect -1554 -2749 -1496 -2715
rect -1462 -2749 -1404 -2715
rect -1370 -2749 -1312 -2715
rect -1278 -2749 -1220 -2715
rect -1186 -2749 -1128 -2715
rect -1094 -2749 -1036 -2715
rect -1002 -2749 -944 -2715
rect -910 -2749 -852 -2715
rect -818 -2749 -760 -2715
rect -726 -2749 -668 -2715
rect -634 -2749 -576 -2715
rect -542 -2749 -484 -2715
rect -450 -2749 -392 -2715
rect -358 -2749 -300 -2715
rect -266 -2749 -208 -2715
rect -174 -2749 -116 -2715
rect -82 -2749 -24 -2715
rect 10 -2749 68 -2715
rect 102 -2749 160 -2715
rect 194 -2749 252 -2715
rect 286 -2749 344 -2715
rect 378 -2749 436 -2715
rect 470 -2749 528 -2715
rect 562 -2749 620 -2715
rect 654 -2749 712 -2715
rect 746 -2749 804 -2715
rect 838 -2749 896 -2715
rect 930 -2749 988 -2715
rect 1022 -2749 1080 -2715
rect 1114 -2749 1172 -2715
rect 1206 -2749 1264 -2715
rect 1298 -2749 1356 -2715
rect 1390 -2749 1448 -2715
rect 1482 -2749 1540 -2715
rect 1574 -2749 1632 -2715
rect 1666 -2749 1724 -2715
rect 1758 -2749 1816 -2715
rect 1850 -2749 1908 -2715
rect 1942 -2749 2000 -2715
rect 2034 -2749 2092 -2715
rect 2126 -2749 2184 -2715
rect 2218 -2749 2276 -2715
rect 2310 -2749 2368 -2715
rect 2402 -2749 2460 -2715
rect 2494 -2749 2552 -2715
rect 2586 -2749 2644 -2715
rect 2678 -2749 2736 -2715
rect 2770 -2749 2828 -2715
rect 2862 -2749 2920 -2715
rect 2954 -2749 3012 -2715
rect 3046 -2749 3104 -2715
rect 3138 -2749 3196 -2715
rect 3230 -2749 3288 -2715
rect 3322 -2749 3380 -2715
rect 3414 -2749 3472 -2715
rect 3506 -2749 3564 -2715
rect 3598 -2749 3656 -2715
rect 3690 -2749 3748 -2715
rect 3782 -2749 3840 -2715
rect 3874 -2749 3932 -2715
rect 3966 -2749 4024 -2715
rect 4058 -2749 4116 -2715
rect 4150 -2749 4208 -2715
rect 4242 -2749 4300 -2715
rect 4334 -2749 4392 -2715
rect 4426 -2749 4484 -2715
rect 4518 -2749 4576 -2715
rect 4610 -2749 4668 -2715
rect 4702 -2749 4760 -2715
rect 4794 -2749 4852 -2715
rect 4886 -2749 4944 -2715
rect 4978 -2749 5036 -2715
rect 5070 -2749 5128 -2715
rect 5162 -2749 5220 -2715
rect 5254 -2749 5312 -2715
rect 5346 -2749 5404 -2715
rect 5438 -2749 5496 -2715
rect 5530 -2749 5588 -2715
rect 5622 -2749 5680 -2715
rect 5714 -2749 5772 -2715
rect 5806 -2749 5864 -2715
rect 5898 -2749 5956 -2715
rect 5990 -2749 6048 -2715
rect 6082 -2749 6140 -2715
rect 6174 -2749 6232 -2715
rect 6266 -2749 6324 -2715
rect 6358 -2749 6416 -2715
rect 6450 -2749 6508 -2715
rect 6542 -2749 6600 -2715
rect 6634 -2749 6692 -2715
rect 6726 -2749 6784 -2715
rect 6818 -2749 6876 -2715
rect 6910 -2749 6968 -2715
rect 7002 -2749 7060 -2715
rect 7094 -2749 7152 -2715
rect 7186 -2749 7244 -2715
rect 7278 -2749 7336 -2715
rect 7370 -2749 7428 -2715
rect 7462 -2749 7520 -2715
rect 7554 -2749 7612 -2715
rect 7646 -2749 7704 -2715
rect 7738 -2749 7796 -2715
rect 7830 -2749 7888 -2715
rect 7922 -2749 7980 -2715
rect 8014 -2749 8072 -2715
rect 8106 -2749 8164 -2715
rect 8198 -2749 8256 -2715
rect 8290 -2749 8348 -2715
rect 8382 -2749 8440 -2715
rect 8474 -2749 8532 -2715
rect 8566 -2749 8624 -2715
rect 8658 -2749 8716 -2715
rect 8750 -2749 8808 -2715
rect 8842 -2749 8900 -2715
rect 8934 -2749 8992 -2715
rect 9026 -2749 9084 -2715
rect 9118 -2749 9176 -2715
rect 9210 -2749 9268 -2715
rect 9302 -2749 9360 -2715
rect 9394 -2749 9452 -2715
rect 9486 -2749 9544 -2715
rect 9578 -2749 9636 -2715
rect 9670 -2749 9728 -2715
rect 9762 -2749 9820 -2715
rect 9854 -2749 9912 -2715
rect 9946 -2749 10004 -2715
rect 10038 -2749 10096 -2715
rect 10130 -2749 10188 -2715
rect 10222 -2749 10280 -2715
rect 10314 -2749 10372 -2715
rect 10406 -2749 10464 -2715
rect 10498 -2749 10556 -2715
rect 10590 -2749 10648 -2715
rect 10682 -2749 10740 -2715
rect 10774 -2749 10832 -2715
rect 10866 -2749 10924 -2715
rect 10958 -2749 11016 -2715
rect 11050 -2749 11108 -2715
rect 11142 -2749 11200 -2715
rect 11234 -2749 11292 -2715
rect 11326 -2749 11384 -2715
rect 11418 -2749 11476 -2715
rect 11510 -2749 11568 -2715
rect 11602 -2749 11660 -2715
rect 11694 -2749 11752 -2715
rect 11786 -2749 11844 -2715
rect 11878 -2749 11936 -2715
rect 11970 -2749 12028 -2715
rect 12062 -2749 12120 -2715
rect 12154 -2749 12212 -2715
rect 12246 -2749 12304 -2715
rect 12338 -2749 12396 -2715
rect 12430 -2749 12488 -2715
rect 12522 -2749 12580 -2715
rect 12614 -2749 12672 -2715
rect 12706 -2749 12764 -2715
rect 12798 -2749 12856 -2715
rect 12890 -2749 12948 -2715
rect 12982 -2749 13040 -2715
rect 13074 -2749 13132 -2715
rect 13166 -2749 13224 -2715
rect 13258 -2749 13316 -2715
rect 13350 -2749 13408 -2715
rect 13442 -2749 13500 -2715
rect 13534 -2749 13592 -2715
rect 13626 -2749 13684 -2715
rect 13718 -2749 13776 -2715
rect 13810 -2749 13868 -2715
rect 13902 -2749 13960 -2715
rect 13994 -2749 14052 -2715
rect 14086 -2749 14144 -2715
rect 14178 -2749 14236 -2715
rect 14270 -2749 14328 -2715
rect 14362 -2749 14420 -2715
rect 14454 -2749 14512 -2715
rect 14546 -2749 14604 -2715
rect 14638 -2749 14696 -2715
rect 14730 -2749 14788 -2715
rect 14822 -2749 14880 -2715
rect 14914 -2749 14972 -2715
rect 15006 -2749 15064 -2715
rect 15098 -2749 15156 -2715
rect 15190 -2749 15248 -2715
rect 15282 -2749 15340 -2715
rect 15374 -2749 15432 -2715
rect 15466 -2749 15524 -2715
rect 15558 -2749 15616 -2715
rect 15650 -2749 15708 -2715
rect 15742 -2749 15800 -2715
rect 15834 -2749 15892 -2715
rect 15926 -2749 15984 -2715
rect 16018 -2749 16076 -2715
rect 16110 -2749 16168 -2715
rect 16202 -2749 16260 -2715
rect 16294 -2749 16352 -2715
rect 16386 -2749 16444 -2715
rect 16478 -2749 16536 -2715
rect 16570 -2749 16628 -2715
rect 16662 -2749 16946 -2715
rect -3193 -2780 16946 -2749
rect -1978 -2996 -1968 -2944
rect -1916 -2996 -1906 -2944
rect -1802 -2958 -1792 -2906
rect -1740 -2958 -1730 -2906
rect 1035 -2952 3062 -2946
rect -225 -2981 479 -2979
rect -231 -3033 -221 -2981
rect -169 -2987 479 -2981
rect -169 -3021 429 -2987
rect 463 -3021 479 -2987
rect 1035 -2986 1072 -2952
rect 1106 -2953 3062 -2952
rect 1106 -2986 3016 -2953
rect 1035 -2987 3016 -2986
rect 3050 -2987 3062 -2953
rect 1035 -2993 3062 -2987
rect 3618 -2948 3676 -2947
rect 5578 -2948 5636 -2947
rect 3618 -2953 5636 -2948
rect 3618 -2987 3630 -2953
rect 3664 -2987 5590 -2953
rect 5624 -2987 5636 -2953
rect 3618 -2992 5636 -2987
rect 3618 -2993 3676 -2992
rect 5578 -2993 5636 -2992
rect 6192 -2948 6250 -2947
rect 8152 -2948 8210 -2947
rect 6192 -2953 8210 -2948
rect 6192 -2987 6204 -2953
rect 6238 -2987 8164 -2953
rect 8198 -2987 8210 -2953
rect 6192 -2992 8210 -2987
rect 6192 -2993 6250 -2992
rect 8152 -2993 8210 -2992
rect 8766 -2948 8824 -2947
rect 8766 -2953 10784 -2948
rect 8766 -2987 8778 -2953
rect 8812 -2954 10784 -2953
rect 8812 -2987 10738 -2954
rect 8766 -2988 10738 -2987
rect 10772 -2988 10784 -2954
rect 8766 -2994 10784 -2988
rect 11366 -2995 11376 -2943
rect 11428 -2995 11438 -2943
rect -169 -3033 479 -3021
rect -1968 -3059 -1201 -3058
rect -1968 -3062 -1272 -3059
rect -1978 -3114 -1968 -3062
rect -1916 -3114 -1272 -3062
rect -1968 -3118 -1272 -3114
rect -1213 -3118 -1201 -3059
rect -1968 -3119 -1201 -3118
rect -3193 -3259 16946 -3228
rect -3193 -3293 -2968 -3259
rect -2934 -3293 -2876 -3259
rect -2842 -3293 -2784 -3259
rect -2750 -3293 -2692 -3259
rect -2658 -3293 -2600 -3259
rect -2566 -3293 -2508 -3259
rect -2474 -3293 -2416 -3259
rect -2382 -3293 -2324 -3259
rect -2290 -3293 -2232 -3259
rect -2198 -3293 -2140 -3259
rect -2106 -3293 -2048 -3259
rect -2014 -3293 -1956 -3259
rect -1922 -3293 -1864 -3259
rect -1830 -3293 -1772 -3259
rect -1738 -3293 -1680 -3259
rect -1646 -3293 -1588 -3259
rect -1554 -3293 -1496 -3259
rect -1462 -3293 -1404 -3259
rect -1370 -3293 -1312 -3259
rect -1278 -3293 -1220 -3259
rect -1186 -3293 -1128 -3259
rect -1094 -3293 -1036 -3259
rect -1002 -3293 -944 -3259
rect -910 -3293 -852 -3259
rect -818 -3293 -760 -3259
rect -726 -3293 -668 -3259
rect -634 -3293 -576 -3259
rect -542 -3293 -484 -3259
rect -450 -3293 -392 -3259
rect -358 -3293 -300 -3259
rect -266 -3293 -208 -3259
rect -174 -3293 -116 -3259
rect -82 -3293 -24 -3259
rect 10 -3293 68 -3259
rect 102 -3293 160 -3259
rect 194 -3293 252 -3259
rect 286 -3293 344 -3259
rect 378 -3293 436 -3259
rect 470 -3293 528 -3259
rect 562 -3293 620 -3259
rect 654 -3293 712 -3259
rect 746 -3293 804 -3259
rect 838 -3293 896 -3259
rect 930 -3293 988 -3259
rect 1022 -3293 1080 -3259
rect 1114 -3293 1172 -3259
rect 1206 -3293 1264 -3259
rect 1298 -3293 1356 -3259
rect 1390 -3293 1448 -3259
rect 1482 -3293 1540 -3259
rect 1574 -3293 1632 -3259
rect 1666 -3293 1724 -3259
rect 1758 -3293 1816 -3259
rect 1850 -3293 1908 -3259
rect 1942 -3293 2000 -3259
rect 2034 -3293 2092 -3259
rect 2126 -3293 2184 -3259
rect 2218 -3293 2276 -3259
rect 2310 -3293 2368 -3259
rect 2402 -3293 2460 -3259
rect 2494 -3293 2552 -3259
rect 2586 -3293 2644 -3259
rect 2678 -3293 2736 -3259
rect 2770 -3293 2828 -3259
rect 2862 -3293 2920 -3259
rect 2954 -3293 3012 -3259
rect 3046 -3293 3104 -3259
rect 3138 -3293 3196 -3259
rect 3230 -3293 3288 -3259
rect 3322 -3293 3380 -3259
rect 3414 -3293 3472 -3259
rect 3506 -3293 3564 -3259
rect 3598 -3293 3656 -3259
rect 3690 -3293 3748 -3259
rect 3782 -3293 3840 -3259
rect 3874 -3293 3932 -3259
rect 3966 -3293 4024 -3259
rect 4058 -3293 4116 -3259
rect 4150 -3293 4208 -3259
rect 4242 -3293 4300 -3259
rect 4334 -3293 4392 -3259
rect 4426 -3293 4484 -3259
rect 4518 -3293 4576 -3259
rect 4610 -3293 4668 -3259
rect 4702 -3293 4760 -3259
rect 4794 -3293 4852 -3259
rect 4886 -3293 4944 -3259
rect 4978 -3293 5036 -3259
rect 5070 -3293 5128 -3259
rect 5162 -3293 5220 -3259
rect 5254 -3293 5312 -3259
rect 5346 -3293 5404 -3259
rect 5438 -3293 5496 -3259
rect 5530 -3293 5588 -3259
rect 5622 -3293 5680 -3259
rect 5714 -3293 5772 -3259
rect 5806 -3293 5864 -3259
rect 5898 -3293 5956 -3259
rect 5990 -3293 6048 -3259
rect 6082 -3293 6140 -3259
rect 6174 -3293 6232 -3259
rect 6266 -3293 6324 -3259
rect 6358 -3293 6416 -3259
rect 6450 -3293 6508 -3259
rect 6542 -3293 6600 -3259
rect 6634 -3293 6692 -3259
rect 6726 -3293 6784 -3259
rect 6818 -3293 6876 -3259
rect 6910 -3293 6968 -3259
rect 7002 -3293 7060 -3259
rect 7094 -3293 7152 -3259
rect 7186 -3293 7244 -3259
rect 7278 -3293 7336 -3259
rect 7370 -3293 7428 -3259
rect 7462 -3293 7520 -3259
rect 7554 -3293 7612 -3259
rect 7646 -3293 7704 -3259
rect 7738 -3293 7796 -3259
rect 7830 -3293 7888 -3259
rect 7922 -3293 7980 -3259
rect 8014 -3293 8072 -3259
rect 8106 -3293 8164 -3259
rect 8198 -3293 8256 -3259
rect 8290 -3293 8348 -3259
rect 8382 -3293 8440 -3259
rect 8474 -3293 8532 -3259
rect 8566 -3293 8624 -3259
rect 8658 -3293 8716 -3259
rect 8750 -3293 8808 -3259
rect 8842 -3293 8900 -3259
rect 8934 -3293 8992 -3259
rect 9026 -3293 9084 -3259
rect 9118 -3293 9176 -3259
rect 9210 -3293 9268 -3259
rect 9302 -3293 9360 -3259
rect 9394 -3293 9452 -3259
rect 9486 -3293 9544 -3259
rect 9578 -3293 9636 -3259
rect 9670 -3293 9728 -3259
rect 9762 -3293 9820 -3259
rect 9854 -3293 9912 -3259
rect 9946 -3293 10004 -3259
rect 10038 -3293 10096 -3259
rect 10130 -3293 10188 -3259
rect 10222 -3293 10280 -3259
rect 10314 -3293 10372 -3259
rect 10406 -3293 10464 -3259
rect 10498 -3293 10556 -3259
rect 10590 -3293 10648 -3259
rect 10682 -3293 10740 -3259
rect 10774 -3293 10832 -3259
rect 10866 -3293 10924 -3259
rect 10958 -3293 11016 -3259
rect 11050 -3293 11108 -3259
rect 11142 -3293 11200 -3259
rect 11234 -3293 11292 -3259
rect 11326 -3293 11384 -3259
rect 11418 -3293 11476 -3259
rect 11510 -3293 11568 -3259
rect 11602 -3293 11660 -3259
rect 11694 -3293 11752 -3259
rect 11786 -3293 11844 -3259
rect 11878 -3293 11936 -3259
rect 11970 -3293 12028 -3259
rect 12062 -3293 12120 -3259
rect 12154 -3293 12212 -3259
rect 12246 -3293 12304 -3259
rect 12338 -3293 12396 -3259
rect 12430 -3293 12488 -3259
rect 12522 -3293 12580 -3259
rect 12614 -3293 12672 -3259
rect 12706 -3293 12764 -3259
rect 12798 -3293 12856 -3259
rect 12890 -3293 12948 -3259
rect 12982 -3293 13040 -3259
rect 13074 -3293 13132 -3259
rect 13166 -3293 13224 -3259
rect 13258 -3293 13316 -3259
rect 13350 -3293 13408 -3259
rect 13442 -3293 13500 -3259
rect 13534 -3293 13592 -3259
rect 13626 -3293 13684 -3259
rect 13718 -3293 13776 -3259
rect 13810 -3293 13868 -3259
rect 13902 -3293 13960 -3259
rect 13994 -3293 14052 -3259
rect 14086 -3293 14144 -3259
rect 14178 -3293 14236 -3259
rect 14270 -3293 14328 -3259
rect 14362 -3293 14420 -3259
rect 14454 -3293 14512 -3259
rect 14546 -3293 14604 -3259
rect 14638 -3293 14696 -3259
rect 14730 -3293 14788 -3259
rect 14822 -3293 14880 -3259
rect 14914 -3293 14972 -3259
rect 15006 -3293 15064 -3259
rect 15098 -3293 15156 -3259
rect 15190 -3293 15248 -3259
rect 15282 -3293 15340 -3259
rect 15374 -3293 15432 -3259
rect 15466 -3293 15524 -3259
rect 15558 -3293 15616 -3259
rect 15650 -3293 15708 -3259
rect 15742 -3293 15800 -3259
rect 15834 -3293 15892 -3259
rect 15926 -3293 15984 -3259
rect 16018 -3293 16076 -3259
rect 16110 -3293 16168 -3259
rect 16202 -3293 16260 -3259
rect 16294 -3293 16352 -3259
rect 16386 -3293 16444 -3259
rect 16478 -3293 16536 -3259
rect 16570 -3293 16628 -3259
rect 16662 -3293 16946 -3259
rect -3193 -3324 16946 -3293
rect 105 -3573 115 -3521
rect 167 -3523 177 -3521
rect 167 -3531 481 -3523
rect 167 -3565 432 -3531
rect 466 -3565 481 -3531
rect 167 -3572 481 -3565
rect 1033 -3565 3062 -3559
rect 1033 -3568 3016 -3565
rect 167 -3573 177 -3572
rect 1033 -3602 1070 -3568
rect 1104 -3599 3016 -3568
rect 3050 -3599 3062 -3565
rect 1104 -3602 3062 -3599
rect 1033 -3610 3062 -3602
rect 3618 -3560 3676 -3559
rect 5578 -3560 5636 -3559
rect 3618 -3565 5636 -3560
rect 3618 -3599 3630 -3565
rect 3664 -3599 5590 -3565
rect 5624 -3599 5636 -3565
rect 3618 -3604 5636 -3599
rect 3618 -3605 3676 -3604
rect 5578 -3605 5636 -3604
rect 6192 -3560 6250 -3559
rect 8152 -3560 8210 -3559
rect 6192 -3565 8210 -3560
rect 6192 -3599 6204 -3565
rect 6238 -3599 8164 -3565
rect 8198 -3599 8210 -3565
rect 6192 -3604 8210 -3599
rect 6192 -3605 6250 -3604
rect 8152 -3605 8210 -3604
rect 8766 -3565 10783 -3557
rect 8766 -3599 8778 -3565
rect 8812 -3568 10783 -3565
rect 8812 -3599 10735 -3568
rect 8766 -3602 10735 -3599
rect 10769 -3602 10783 -3568
rect 8766 -3607 10783 -3602
rect 10723 -3608 10781 -3607
rect 11363 -3609 11373 -3557
rect 11425 -3609 11435 -3557
rect -3193 -3803 16946 -3772
rect -3193 -3837 -2968 -3803
rect -2934 -3837 -2876 -3803
rect -2842 -3837 -2784 -3803
rect -2750 -3837 -2692 -3803
rect -2658 -3837 -2600 -3803
rect -2566 -3837 -2508 -3803
rect -2474 -3837 -2416 -3803
rect -2382 -3837 -2324 -3803
rect -2290 -3837 -2232 -3803
rect -2198 -3837 -2140 -3803
rect -2106 -3837 -2048 -3803
rect -2014 -3837 -1956 -3803
rect -1922 -3837 -1864 -3803
rect -1830 -3837 -1772 -3803
rect -1738 -3837 -1680 -3803
rect -1646 -3837 -1588 -3803
rect -1554 -3837 -1496 -3803
rect -1462 -3837 -1404 -3803
rect -1370 -3837 -1312 -3803
rect -1278 -3837 -1220 -3803
rect -1186 -3837 -1128 -3803
rect -1094 -3837 -1036 -3803
rect -1002 -3837 -944 -3803
rect -910 -3837 -852 -3803
rect -818 -3837 -760 -3803
rect -726 -3837 -668 -3803
rect -634 -3837 -576 -3803
rect -542 -3837 -484 -3803
rect -450 -3837 -392 -3803
rect -358 -3837 -300 -3803
rect -266 -3837 -208 -3803
rect -174 -3837 -116 -3803
rect -82 -3837 -24 -3803
rect 10 -3837 68 -3803
rect 102 -3837 160 -3803
rect 194 -3837 252 -3803
rect 286 -3837 344 -3803
rect 378 -3837 436 -3803
rect 470 -3837 528 -3803
rect 562 -3837 620 -3803
rect 654 -3837 712 -3803
rect 746 -3837 804 -3803
rect 838 -3837 896 -3803
rect 930 -3837 988 -3803
rect 1022 -3837 1080 -3803
rect 1114 -3837 1172 -3803
rect 1206 -3837 1264 -3803
rect 1298 -3837 1356 -3803
rect 1390 -3837 1448 -3803
rect 1482 -3837 1540 -3803
rect 1574 -3837 1632 -3803
rect 1666 -3837 1724 -3803
rect 1758 -3837 1816 -3803
rect 1850 -3837 1908 -3803
rect 1942 -3837 2000 -3803
rect 2034 -3837 2092 -3803
rect 2126 -3837 2184 -3803
rect 2218 -3837 2276 -3803
rect 2310 -3837 2368 -3803
rect 2402 -3837 2460 -3803
rect 2494 -3837 2552 -3803
rect 2586 -3837 2644 -3803
rect 2678 -3837 2736 -3803
rect 2770 -3837 2828 -3803
rect 2862 -3837 2920 -3803
rect 2954 -3837 3012 -3803
rect 3046 -3837 3104 -3803
rect 3138 -3837 3196 -3803
rect 3230 -3837 3288 -3803
rect 3322 -3837 3380 -3803
rect 3414 -3837 3472 -3803
rect 3506 -3837 3564 -3803
rect 3598 -3837 3656 -3803
rect 3690 -3837 3748 -3803
rect 3782 -3837 3840 -3803
rect 3874 -3837 3932 -3803
rect 3966 -3837 4024 -3803
rect 4058 -3837 4116 -3803
rect 4150 -3837 4208 -3803
rect 4242 -3837 4300 -3803
rect 4334 -3837 4392 -3803
rect 4426 -3837 4484 -3803
rect 4518 -3837 4576 -3803
rect 4610 -3837 4668 -3803
rect 4702 -3837 4760 -3803
rect 4794 -3837 4852 -3803
rect 4886 -3837 4944 -3803
rect 4978 -3837 5036 -3803
rect 5070 -3837 5128 -3803
rect 5162 -3837 5220 -3803
rect 5254 -3837 5312 -3803
rect 5346 -3837 5404 -3803
rect 5438 -3837 5496 -3803
rect 5530 -3837 5588 -3803
rect 5622 -3837 5680 -3803
rect 5714 -3837 5772 -3803
rect 5806 -3837 5864 -3803
rect 5898 -3837 5956 -3803
rect 5990 -3837 6048 -3803
rect 6082 -3837 6140 -3803
rect 6174 -3837 6232 -3803
rect 6266 -3837 6324 -3803
rect 6358 -3837 6416 -3803
rect 6450 -3837 6508 -3803
rect 6542 -3837 6600 -3803
rect 6634 -3837 6692 -3803
rect 6726 -3837 6784 -3803
rect 6818 -3837 6876 -3803
rect 6910 -3837 6968 -3803
rect 7002 -3837 7060 -3803
rect 7094 -3837 7152 -3803
rect 7186 -3837 7244 -3803
rect 7278 -3837 7336 -3803
rect 7370 -3837 7428 -3803
rect 7462 -3837 7520 -3803
rect 7554 -3837 7612 -3803
rect 7646 -3837 7704 -3803
rect 7738 -3837 7796 -3803
rect 7830 -3837 7888 -3803
rect 7922 -3837 7980 -3803
rect 8014 -3837 8072 -3803
rect 8106 -3837 8164 -3803
rect 8198 -3837 8256 -3803
rect 8290 -3837 8348 -3803
rect 8382 -3837 8440 -3803
rect 8474 -3837 8532 -3803
rect 8566 -3837 8624 -3803
rect 8658 -3837 8716 -3803
rect 8750 -3837 8808 -3803
rect 8842 -3837 8900 -3803
rect 8934 -3837 8992 -3803
rect 9026 -3837 9084 -3803
rect 9118 -3837 9176 -3803
rect 9210 -3837 9268 -3803
rect 9302 -3837 9360 -3803
rect 9394 -3837 9452 -3803
rect 9486 -3837 9544 -3803
rect 9578 -3837 9636 -3803
rect 9670 -3837 9728 -3803
rect 9762 -3837 9820 -3803
rect 9854 -3837 9912 -3803
rect 9946 -3837 10004 -3803
rect 10038 -3837 10096 -3803
rect 10130 -3837 10188 -3803
rect 10222 -3837 10280 -3803
rect 10314 -3837 10372 -3803
rect 10406 -3837 10464 -3803
rect 10498 -3837 10556 -3803
rect 10590 -3837 10648 -3803
rect 10682 -3837 10740 -3803
rect 10774 -3837 10832 -3803
rect 10866 -3837 10924 -3803
rect 10958 -3837 11016 -3803
rect 11050 -3837 11108 -3803
rect 11142 -3837 11200 -3803
rect 11234 -3837 11292 -3803
rect 11326 -3837 11384 -3803
rect 11418 -3837 11476 -3803
rect 11510 -3837 11568 -3803
rect 11602 -3837 11660 -3803
rect 11694 -3837 11752 -3803
rect 11786 -3837 11844 -3803
rect 11878 -3837 11936 -3803
rect 11970 -3837 12028 -3803
rect 12062 -3837 12120 -3803
rect 12154 -3837 12212 -3803
rect 12246 -3837 12304 -3803
rect 12338 -3837 12396 -3803
rect 12430 -3837 12488 -3803
rect 12522 -3837 12580 -3803
rect 12614 -3837 12672 -3803
rect 12706 -3837 12764 -3803
rect 12798 -3837 12856 -3803
rect 12890 -3837 12948 -3803
rect 12982 -3837 13040 -3803
rect 13074 -3837 13132 -3803
rect 13166 -3837 13224 -3803
rect 13258 -3837 13316 -3803
rect 13350 -3837 13408 -3803
rect 13442 -3837 13500 -3803
rect 13534 -3837 13592 -3803
rect 13626 -3837 13684 -3803
rect 13718 -3837 13776 -3803
rect 13810 -3837 13868 -3803
rect 13902 -3837 13960 -3803
rect 13994 -3837 14052 -3803
rect 14086 -3837 14144 -3803
rect 14178 -3837 14236 -3803
rect 14270 -3837 14328 -3803
rect 14362 -3837 14420 -3803
rect 14454 -3837 14512 -3803
rect 14546 -3837 14604 -3803
rect 14638 -3837 14696 -3803
rect 14730 -3837 14788 -3803
rect 14822 -3837 14880 -3803
rect 14914 -3837 14972 -3803
rect 15006 -3837 15064 -3803
rect 15098 -3837 15156 -3803
rect 15190 -3837 15248 -3803
rect 15282 -3837 15340 -3803
rect 15374 -3837 15432 -3803
rect 15466 -3837 15524 -3803
rect 15558 -3837 15616 -3803
rect 15650 -3837 15708 -3803
rect 15742 -3837 15800 -3803
rect 15834 -3837 15892 -3803
rect 15926 -3837 15984 -3803
rect 16018 -3837 16076 -3803
rect 16110 -3837 16168 -3803
rect 16202 -3837 16260 -3803
rect 16294 -3837 16352 -3803
rect 16386 -3837 16444 -3803
rect 16478 -3837 16536 -3803
rect 16570 -3837 16628 -3803
rect 16662 -3837 16946 -3803
rect -3193 -3868 16946 -3837
rect 12467 -3965 12520 -3940
rect 12467 -3972 12480 -3965
rect 12514 -3972 12520 -3965
rect 12456 -4024 12466 -3972
rect 12518 -4024 12520 -3972
rect 417 -4083 427 -4031
rect 479 -4083 489 -4031
rect 1069 -4035 1127 -4034
rect 3029 -4035 3087 -4034
rect 1069 -4040 3087 -4035
rect 1069 -4074 1081 -4040
rect 1115 -4074 3041 -4040
rect 3075 -4074 3087 -4040
rect 1069 -4079 3087 -4074
rect 1069 -4080 1127 -4079
rect 3029 -4080 3087 -4079
rect 3643 -4035 3701 -4034
rect 5603 -4035 5661 -4034
rect 3643 -4040 5661 -4035
rect 3643 -4074 3655 -4040
rect 3689 -4074 5615 -4040
rect 5649 -4074 5661 -4040
rect 3643 -4079 5661 -4074
rect 3643 -4080 3701 -4079
rect 5603 -4080 5661 -4079
rect 6217 -4035 6275 -4034
rect 8177 -4035 8235 -4034
rect 6217 -4040 8235 -4035
rect 6217 -4074 6229 -4040
rect 6263 -4074 8189 -4040
rect 8223 -4074 8235 -4040
rect 6217 -4079 8235 -4074
rect 6217 -4080 6275 -4079
rect 8177 -4080 8235 -4079
rect 8791 -4035 8849 -4034
rect 10751 -4035 10809 -4034
rect 8791 -4040 10809 -4035
rect 8791 -4074 8806 -4040
rect 8840 -4074 10763 -4040
rect 10797 -4074 10809 -4040
rect 12467 -4037 12520 -4024
rect 13023 -3975 13738 -3968
rect 13023 -4009 13042 -3975
rect 13076 -4008 13738 -3975
rect 13076 -4009 13685 -4008
rect 12745 -4031 12755 -4028
rect 8791 -4079 10809 -4074
rect 8791 -4080 8849 -4079
rect 10751 -4080 10809 -4079
rect 11367 -4119 11377 -4067
rect 11429 -4119 11439 -4067
rect 12467 -4071 12480 -4037
rect 12514 -4071 12520 -4037
rect 12467 -4086 12520 -4071
rect 12548 -4039 12755 -4031
rect 12807 -4031 12817 -4028
rect 12548 -4073 12568 -4039
rect 12602 -4073 12659 -4039
rect 12693 -4073 12755 -4039
rect 12807 -4041 12993 -4031
rect 12548 -4080 12755 -4073
rect 12807 -4075 12858 -4041
rect 12892 -4075 12942 -4041
rect 12976 -4075 12993 -4041
rect 12807 -4080 12993 -4075
rect 13023 -4042 13685 -4009
rect 13719 -4042 13738 -4008
rect 13023 -4052 13738 -4042
rect 12846 -4081 12991 -4080
rect 12456 -4138 12466 -4086
rect 12518 -4138 12520 -4086
rect 13023 -4086 13039 -4052
rect 13073 -4086 13738 -4052
rect 15236 -3996 15294 -3990
rect 15329 -3996 15387 -3990
rect 15236 -4030 15248 -3996
rect 15282 -4030 15341 -3996
rect 15375 -4030 15394 -3996
rect 13023 -4091 13738 -4086
rect 13027 -4092 13085 -4091
rect 14618 -4118 14628 -4064
rect 14682 -4072 14692 -4064
rect 15236 -4072 15394 -4030
rect 14682 -4092 16946 -4072
rect 14682 -4112 15248 -4092
rect 14682 -4118 14692 -4112
rect 15236 -4126 15248 -4112
rect 15282 -4126 15340 -4092
rect 15374 -4112 16946 -4092
rect 15374 -4126 15394 -4112
rect 15236 -4132 15294 -4126
rect 15328 -4132 15386 -4126
rect 12467 -4145 12480 -4138
rect 12514 -4145 12520 -4138
rect 12467 -4177 12520 -4145
rect -3193 -4347 16946 -4316
rect -3193 -4381 -2968 -4347
rect -2934 -4381 -2876 -4347
rect -2842 -4381 -2784 -4347
rect -2750 -4381 -2692 -4347
rect -2658 -4381 -2600 -4347
rect -2566 -4381 -2508 -4347
rect -2474 -4381 -2416 -4347
rect -2382 -4381 -2324 -4347
rect -2290 -4381 -2232 -4347
rect -2198 -4381 -2140 -4347
rect -2106 -4381 -2048 -4347
rect -2014 -4381 -1956 -4347
rect -1922 -4381 -1864 -4347
rect -1830 -4381 -1772 -4347
rect -1738 -4381 -1680 -4347
rect -1646 -4381 -1588 -4347
rect -1554 -4381 -1496 -4347
rect -1462 -4381 -1404 -4347
rect -1370 -4381 -1312 -4347
rect -1278 -4381 -1220 -4347
rect -1186 -4381 -1128 -4347
rect -1094 -4381 -1036 -4347
rect -1002 -4381 -944 -4347
rect -910 -4381 -852 -4347
rect -818 -4381 -760 -4347
rect -726 -4381 -668 -4347
rect -634 -4381 -576 -4347
rect -542 -4381 -484 -4347
rect -450 -4381 -392 -4347
rect -358 -4381 -300 -4347
rect -266 -4381 -208 -4347
rect -174 -4381 -116 -4347
rect -82 -4381 -24 -4347
rect 10 -4381 68 -4347
rect 102 -4381 160 -4347
rect 194 -4381 252 -4347
rect 286 -4381 344 -4347
rect 378 -4381 436 -4347
rect 470 -4381 528 -4347
rect 562 -4381 620 -4347
rect 654 -4381 712 -4347
rect 746 -4381 804 -4347
rect 838 -4381 896 -4347
rect 930 -4381 988 -4347
rect 1022 -4381 1080 -4347
rect 1114 -4381 1172 -4347
rect 1206 -4381 1264 -4347
rect 1298 -4381 1356 -4347
rect 1390 -4381 1448 -4347
rect 1482 -4381 1540 -4347
rect 1574 -4381 1632 -4347
rect 1666 -4381 1724 -4347
rect 1758 -4381 1816 -4347
rect 1850 -4381 1908 -4347
rect 1942 -4381 2000 -4347
rect 2034 -4381 2092 -4347
rect 2126 -4381 2184 -4347
rect 2218 -4381 2276 -4347
rect 2310 -4381 2368 -4347
rect 2402 -4381 2460 -4347
rect 2494 -4381 2552 -4347
rect 2586 -4381 2644 -4347
rect 2678 -4381 2736 -4347
rect 2770 -4381 2828 -4347
rect 2862 -4381 2920 -4347
rect 2954 -4381 3012 -4347
rect 3046 -4381 3104 -4347
rect 3138 -4381 3196 -4347
rect 3230 -4381 3288 -4347
rect 3322 -4381 3380 -4347
rect 3414 -4381 3472 -4347
rect 3506 -4381 3564 -4347
rect 3598 -4381 3656 -4347
rect 3690 -4381 3748 -4347
rect 3782 -4381 3840 -4347
rect 3874 -4381 3932 -4347
rect 3966 -4381 4024 -4347
rect 4058 -4381 4116 -4347
rect 4150 -4381 4208 -4347
rect 4242 -4381 4300 -4347
rect 4334 -4381 4392 -4347
rect 4426 -4381 4484 -4347
rect 4518 -4381 4576 -4347
rect 4610 -4381 4668 -4347
rect 4702 -4381 4760 -4347
rect 4794 -4381 4852 -4347
rect 4886 -4381 4944 -4347
rect 4978 -4381 5036 -4347
rect 5070 -4381 5128 -4347
rect 5162 -4381 5220 -4347
rect 5254 -4381 5312 -4347
rect 5346 -4381 5404 -4347
rect 5438 -4381 5496 -4347
rect 5530 -4381 5588 -4347
rect 5622 -4381 5680 -4347
rect 5714 -4381 5772 -4347
rect 5806 -4381 5864 -4347
rect 5898 -4381 5956 -4347
rect 5990 -4381 6048 -4347
rect 6082 -4381 6140 -4347
rect 6174 -4381 6232 -4347
rect 6266 -4381 6324 -4347
rect 6358 -4381 6416 -4347
rect 6450 -4381 6508 -4347
rect 6542 -4381 6600 -4347
rect 6634 -4381 6692 -4347
rect 6726 -4381 6784 -4347
rect 6818 -4381 6876 -4347
rect 6910 -4381 6968 -4347
rect 7002 -4381 7060 -4347
rect 7094 -4381 7152 -4347
rect 7186 -4381 7244 -4347
rect 7278 -4381 7336 -4347
rect 7370 -4381 7428 -4347
rect 7462 -4381 7520 -4347
rect 7554 -4381 7612 -4347
rect 7646 -4381 7704 -4347
rect 7738 -4381 7796 -4347
rect 7830 -4381 7888 -4347
rect 7922 -4381 7980 -4347
rect 8014 -4381 8072 -4347
rect 8106 -4381 8164 -4347
rect 8198 -4381 8256 -4347
rect 8290 -4381 8348 -4347
rect 8382 -4381 8440 -4347
rect 8474 -4381 8532 -4347
rect 8566 -4381 8624 -4347
rect 8658 -4381 8716 -4347
rect 8750 -4381 8808 -4347
rect 8842 -4381 8900 -4347
rect 8934 -4381 8992 -4347
rect 9026 -4381 9084 -4347
rect 9118 -4381 9176 -4347
rect 9210 -4381 9268 -4347
rect 9302 -4381 9360 -4347
rect 9394 -4381 9452 -4347
rect 9486 -4381 9544 -4347
rect 9578 -4381 9636 -4347
rect 9670 -4381 9728 -4347
rect 9762 -4381 9820 -4347
rect 9854 -4381 9912 -4347
rect 9946 -4381 10004 -4347
rect 10038 -4381 10096 -4347
rect 10130 -4381 10188 -4347
rect 10222 -4381 10280 -4347
rect 10314 -4381 10372 -4347
rect 10406 -4381 10464 -4347
rect 10498 -4381 10556 -4347
rect 10590 -4381 10648 -4347
rect 10682 -4381 10740 -4347
rect 10774 -4381 10832 -4347
rect 10866 -4381 10924 -4347
rect 10958 -4381 11016 -4347
rect 11050 -4381 11108 -4347
rect 11142 -4381 11200 -4347
rect 11234 -4381 11292 -4347
rect 11326 -4381 11384 -4347
rect 11418 -4381 11476 -4347
rect 11510 -4381 11568 -4347
rect 11602 -4381 11660 -4347
rect 11694 -4381 11752 -4347
rect 11786 -4381 11844 -4347
rect 11878 -4381 11936 -4347
rect 11970 -4381 12028 -4347
rect 12062 -4381 12120 -4347
rect 12154 -4381 12212 -4347
rect 12246 -4381 12304 -4347
rect 12338 -4381 12396 -4347
rect 12430 -4381 12488 -4347
rect 12522 -4381 12580 -4347
rect 12614 -4381 12672 -4347
rect 12706 -4381 12764 -4347
rect 12798 -4381 12856 -4347
rect 12890 -4381 12948 -4347
rect 12982 -4381 13040 -4347
rect 13074 -4381 13132 -4347
rect 13166 -4381 13224 -4347
rect 13258 -4381 13316 -4347
rect 13350 -4381 13408 -4347
rect 13442 -4381 13500 -4347
rect 13534 -4381 13592 -4347
rect 13626 -4381 13684 -4347
rect 13718 -4381 13776 -4347
rect 13810 -4381 13868 -4347
rect 13902 -4381 13960 -4347
rect 13994 -4381 14052 -4347
rect 14086 -4381 14144 -4347
rect 14178 -4381 14236 -4347
rect 14270 -4381 14328 -4347
rect 14362 -4381 14420 -4347
rect 14454 -4381 14512 -4347
rect 14546 -4381 14604 -4347
rect 14638 -4381 14696 -4347
rect 14730 -4381 14788 -4347
rect 14822 -4381 14880 -4347
rect 14914 -4381 14972 -4347
rect 15006 -4381 15064 -4347
rect 15098 -4381 15156 -4347
rect 15190 -4381 15248 -4347
rect 15282 -4381 15340 -4347
rect 15374 -4381 15432 -4347
rect 15466 -4381 15524 -4347
rect 15558 -4381 15616 -4347
rect 15650 -4381 15708 -4347
rect 15742 -4381 15800 -4347
rect 15834 -4381 15892 -4347
rect 15926 -4381 15984 -4347
rect 16018 -4381 16076 -4347
rect 16110 -4381 16168 -4347
rect 16202 -4381 16260 -4347
rect 16294 -4381 16352 -4347
rect 16386 -4381 16444 -4347
rect 16478 -4381 16536 -4347
rect 16570 -4381 16628 -4347
rect 16662 -4381 16946 -4347
rect -3193 -4412 16946 -4381
rect 15236 -4606 15294 -4600
rect 15329 -4606 15387 -4600
rect -866 -4613 -771 -4608
rect -867 -4619 -771 -4613
rect -867 -4653 -855 -4619
rect -821 -4653 -771 -4619
rect -867 -4659 -771 -4653
rect -866 -4663 -771 -4659
rect -716 -4663 -706 -4608
rect 105 -4647 115 -4643
rect -866 -4666 -706 -4663
rect -253 -4656 115 -4647
rect -253 -4690 -210 -4656
rect -176 -4690 115 -4656
rect -253 -4693 115 -4690
rect -222 -4696 -164 -4693
rect 105 -4695 115 -4693
rect 167 -4695 177 -4643
rect 414 -4662 424 -4610
rect 476 -4662 486 -4610
rect 15236 -4640 15248 -4606
rect 15282 -4640 15341 -4606
rect 15375 -4616 15394 -4606
rect 15375 -4640 16946 -4616
rect 1042 -4647 1100 -4646
rect 3002 -4647 3060 -4646
rect 1042 -4652 3060 -4647
rect 1042 -4686 1054 -4652
rect 1088 -4686 3014 -4652
rect 3048 -4686 3060 -4652
rect 1042 -4691 3060 -4686
rect 1042 -4692 1100 -4691
rect 3002 -4692 3060 -4691
rect 3616 -4647 3674 -4646
rect 5576 -4647 5634 -4646
rect 3616 -4652 5634 -4647
rect 3616 -4686 3628 -4652
rect 3662 -4686 5588 -4652
rect 5622 -4686 5634 -4652
rect 3616 -4691 5634 -4686
rect 3616 -4692 3674 -4691
rect 5576 -4692 5634 -4691
rect 6190 -4647 6248 -4646
rect 8150 -4647 8208 -4646
rect 6190 -4652 8208 -4647
rect 6190 -4686 6202 -4652
rect 6236 -4686 8162 -4652
rect 8196 -4686 8208 -4652
rect 6190 -4691 8208 -4686
rect 6190 -4692 6248 -4691
rect 8150 -4692 8208 -4691
rect 8764 -4647 8822 -4646
rect 10724 -4647 10782 -4646
rect 8764 -4652 10782 -4647
rect 8764 -4686 8776 -4652
rect 8810 -4686 10736 -4652
rect 10770 -4686 10782 -4652
rect 8764 -4691 10782 -4686
rect 8764 -4692 8822 -4691
rect 10724 -4692 10782 -4691
rect 11365 -4697 11375 -4645
rect 11427 -4697 11437 -4645
rect 13671 -4686 13735 -4642
rect 13671 -4720 13685 -4686
rect 13719 -4720 13735 -4686
rect 12746 -4736 12756 -4734
rect 7153 -4737 12756 -4736
rect 7153 -4789 7163 -4737
rect 7215 -4786 12756 -4737
rect 12808 -4736 12818 -4734
rect 13671 -4736 13735 -4720
rect 12808 -4786 13735 -4736
rect 15236 -4656 16946 -4640
rect 15236 -4701 15394 -4656
rect 15236 -4702 15340 -4701
rect 15236 -4736 15248 -4702
rect 15282 -4735 15340 -4702
rect 15374 -4735 15394 -4701
rect 15282 -4736 15394 -4735
rect 15236 -4742 15294 -4736
rect 15328 -4741 15386 -4736
rect 7215 -4789 13735 -4786
rect 7153 -4790 13735 -4789
rect 13671 -4791 13735 -4790
rect -3193 -4891 16946 -4860
rect -3193 -4925 -2968 -4891
rect -2934 -4925 -2876 -4891
rect -2842 -4925 -2784 -4891
rect -2750 -4925 -2692 -4891
rect -2658 -4925 -2600 -4891
rect -2566 -4925 -2508 -4891
rect -2474 -4925 -2416 -4891
rect -2382 -4925 -2324 -4891
rect -2290 -4925 -2232 -4891
rect -2198 -4925 -2140 -4891
rect -2106 -4925 -2048 -4891
rect -2014 -4925 -1956 -4891
rect -1922 -4925 -1864 -4891
rect -1830 -4925 -1772 -4891
rect -1738 -4925 -1680 -4891
rect -1646 -4925 -1588 -4891
rect -1554 -4925 -1496 -4891
rect -1462 -4925 -1404 -4891
rect -1370 -4925 -1312 -4891
rect -1278 -4925 -1220 -4891
rect -1186 -4925 -1128 -4891
rect -1094 -4925 -1036 -4891
rect -1002 -4925 -944 -4891
rect -910 -4925 -852 -4891
rect -818 -4925 -760 -4891
rect -726 -4925 -668 -4891
rect -634 -4925 -576 -4891
rect -542 -4925 -484 -4891
rect -450 -4925 -392 -4891
rect -358 -4925 -300 -4891
rect -266 -4925 -208 -4891
rect -174 -4925 -116 -4891
rect -82 -4925 -24 -4891
rect 10 -4925 68 -4891
rect 102 -4925 160 -4891
rect 194 -4925 252 -4891
rect 286 -4925 344 -4891
rect 378 -4925 436 -4891
rect 470 -4925 528 -4891
rect 562 -4925 620 -4891
rect 654 -4925 712 -4891
rect 746 -4925 804 -4891
rect 838 -4925 896 -4891
rect 930 -4925 988 -4891
rect 1022 -4925 1080 -4891
rect 1114 -4925 1172 -4891
rect 1206 -4925 1264 -4891
rect 1298 -4925 1356 -4891
rect 1390 -4925 1448 -4891
rect 1482 -4925 1540 -4891
rect 1574 -4925 1632 -4891
rect 1666 -4925 1724 -4891
rect 1758 -4925 1816 -4891
rect 1850 -4925 1908 -4891
rect 1942 -4925 2000 -4891
rect 2034 -4925 2092 -4891
rect 2126 -4925 2184 -4891
rect 2218 -4925 2276 -4891
rect 2310 -4925 2368 -4891
rect 2402 -4925 2460 -4891
rect 2494 -4925 2552 -4891
rect 2586 -4925 2644 -4891
rect 2678 -4925 2736 -4891
rect 2770 -4925 2828 -4891
rect 2862 -4925 2920 -4891
rect 2954 -4925 3012 -4891
rect 3046 -4925 3104 -4891
rect 3138 -4925 3196 -4891
rect 3230 -4925 3288 -4891
rect 3322 -4925 3380 -4891
rect 3414 -4925 3472 -4891
rect 3506 -4925 3564 -4891
rect 3598 -4925 3656 -4891
rect 3690 -4925 3748 -4891
rect 3782 -4925 3840 -4891
rect 3874 -4925 3932 -4891
rect 3966 -4925 4024 -4891
rect 4058 -4925 4116 -4891
rect 4150 -4925 4208 -4891
rect 4242 -4925 4300 -4891
rect 4334 -4925 4392 -4891
rect 4426 -4925 4484 -4891
rect 4518 -4925 4576 -4891
rect 4610 -4925 4668 -4891
rect 4702 -4925 4760 -4891
rect 4794 -4925 4852 -4891
rect 4886 -4925 4944 -4891
rect 4978 -4925 5036 -4891
rect 5070 -4925 5128 -4891
rect 5162 -4925 5220 -4891
rect 5254 -4925 5312 -4891
rect 5346 -4925 5404 -4891
rect 5438 -4925 5496 -4891
rect 5530 -4925 5588 -4891
rect 5622 -4925 5680 -4891
rect 5714 -4925 5772 -4891
rect 5806 -4925 5864 -4891
rect 5898 -4925 5956 -4891
rect 5990 -4925 6048 -4891
rect 6082 -4925 6140 -4891
rect 6174 -4925 6232 -4891
rect 6266 -4925 6324 -4891
rect 6358 -4925 6416 -4891
rect 6450 -4925 6508 -4891
rect 6542 -4925 6600 -4891
rect 6634 -4925 6692 -4891
rect 6726 -4925 6784 -4891
rect 6818 -4925 6876 -4891
rect 6910 -4925 6968 -4891
rect 7002 -4925 7060 -4891
rect 7094 -4925 7152 -4891
rect 7186 -4925 7244 -4891
rect 7278 -4925 7336 -4891
rect 7370 -4925 7428 -4891
rect 7462 -4925 7520 -4891
rect 7554 -4925 7612 -4891
rect 7646 -4925 7704 -4891
rect 7738 -4925 7796 -4891
rect 7830 -4925 7888 -4891
rect 7922 -4925 7980 -4891
rect 8014 -4925 8072 -4891
rect 8106 -4925 8164 -4891
rect 8198 -4925 8256 -4891
rect 8290 -4925 8348 -4891
rect 8382 -4925 8440 -4891
rect 8474 -4925 8532 -4891
rect 8566 -4925 8624 -4891
rect 8658 -4925 8716 -4891
rect 8750 -4925 8808 -4891
rect 8842 -4925 8900 -4891
rect 8934 -4925 8992 -4891
rect 9026 -4925 9084 -4891
rect 9118 -4925 9176 -4891
rect 9210 -4925 9268 -4891
rect 9302 -4925 9360 -4891
rect 9394 -4925 9452 -4891
rect 9486 -4925 9544 -4891
rect 9578 -4925 9636 -4891
rect 9670 -4925 9728 -4891
rect 9762 -4925 9820 -4891
rect 9854 -4925 9912 -4891
rect 9946 -4925 10004 -4891
rect 10038 -4925 10096 -4891
rect 10130 -4925 10188 -4891
rect 10222 -4925 10280 -4891
rect 10314 -4925 10372 -4891
rect 10406 -4925 10464 -4891
rect 10498 -4925 10556 -4891
rect 10590 -4925 10648 -4891
rect 10682 -4925 10740 -4891
rect 10774 -4925 10832 -4891
rect 10866 -4925 10924 -4891
rect 10958 -4925 11016 -4891
rect 11050 -4925 11108 -4891
rect 11142 -4925 11200 -4891
rect 11234 -4925 11292 -4891
rect 11326 -4925 11384 -4891
rect 11418 -4925 11476 -4891
rect 11510 -4925 11568 -4891
rect 11602 -4925 11660 -4891
rect 11694 -4925 11752 -4891
rect 11786 -4925 11844 -4891
rect 11878 -4925 11936 -4891
rect 11970 -4925 12028 -4891
rect 12062 -4925 12120 -4891
rect 12154 -4925 12212 -4891
rect 12246 -4925 12304 -4891
rect 12338 -4925 12396 -4891
rect 12430 -4925 12488 -4891
rect 12522 -4925 12580 -4891
rect 12614 -4925 12672 -4891
rect 12706 -4925 12764 -4891
rect 12798 -4925 12856 -4891
rect 12890 -4925 12948 -4891
rect 12982 -4925 13040 -4891
rect 13074 -4925 13132 -4891
rect 13166 -4925 13224 -4891
rect 13258 -4925 13316 -4891
rect 13350 -4925 13408 -4891
rect 13442 -4925 13500 -4891
rect 13534 -4925 13592 -4891
rect 13626 -4925 13684 -4891
rect 13718 -4925 13776 -4891
rect 13810 -4925 13868 -4891
rect 13902 -4925 13960 -4891
rect 13994 -4925 14052 -4891
rect 14086 -4925 14144 -4891
rect 14178 -4925 14236 -4891
rect 14270 -4925 14328 -4891
rect 14362 -4925 14420 -4891
rect 14454 -4925 14512 -4891
rect 14546 -4925 14604 -4891
rect 14638 -4925 14696 -4891
rect 14730 -4925 14788 -4891
rect 14822 -4925 14880 -4891
rect 14914 -4925 14972 -4891
rect 15006 -4925 15064 -4891
rect 15098 -4925 15156 -4891
rect 15190 -4925 15248 -4891
rect 15282 -4925 15340 -4891
rect 15374 -4925 15432 -4891
rect 15466 -4925 15524 -4891
rect 15558 -4925 15616 -4891
rect 15650 -4925 15708 -4891
rect 15742 -4925 15800 -4891
rect 15834 -4925 15892 -4891
rect 15926 -4925 15984 -4891
rect 16018 -4925 16076 -4891
rect 16110 -4925 16168 -4891
rect 16202 -4925 16260 -4891
rect 16294 -4925 16352 -4891
rect 16386 -4925 16444 -4891
rect 16478 -4925 16536 -4891
rect 16570 -4925 16628 -4891
rect 16662 -4925 16946 -4891
rect -3193 -4956 16946 -4925
rect 13026 -5061 13084 -5054
rect 13026 -5095 13038 -5061
rect 13072 -5062 13084 -5061
rect 13072 -5095 13737 -5062
rect 13026 -5096 13737 -5095
rect 12548 -5118 12992 -5117
rect 12548 -5120 12752 -5118
rect 417 -5172 427 -5120
rect 479 -5172 489 -5120
rect 1070 -5124 1128 -5123
rect 3030 -5124 3088 -5123
rect 1070 -5129 3088 -5124
rect 1070 -5163 1082 -5129
rect 1116 -5163 3042 -5129
rect 3076 -5163 3088 -5129
rect 1070 -5168 3088 -5163
rect 1070 -5169 1128 -5168
rect 3030 -5169 3088 -5168
rect 3644 -5124 3702 -5123
rect 5604 -5124 5662 -5123
rect 3644 -5129 5662 -5124
rect 3644 -5163 3656 -5129
rect 3690 -5163 5616 -5129
rect 5650 -5163 5662 -5129
rect 3644 -5168 5662 -5163
rect 3644 -5169 3702 -5168
rect 5604 -5169 5662 -5168
rect 6218 -5124 6276 -5123
rect 8178 -5124 8236 -5123
rect 6218 -5129 8236 -5124
rect 6218 -5163 6230 -5129
rect 6264 -5163 8190 -5129
rect 8224 -5163 8236 -5129
rect 6218 -5168 8236 -5163
rect 6218 -5169 6276 -5168
rect 8178 -5169 8236 -5168
rect 8792 -5124 8850 -5123
rect 10752 -5124 10810 -5123
rect 8792 -5129 10810 -5124
rect 8792 -5163 8804 -5129
rect 8838 -5163 10764 -5129
rect 10798 -5163 10810 -5129
rect 12546 -5126 12752 -5120
rect 12804 -5126 12992 -5118
rect 8792 -5168 10810 -5163
rect 8792 -5169 8850 -5168
rect 10752 -5169 10810 -5168
rect 11370 -5204 11380 -5152
rect 11432 -5204 11442 -5152
rect 12546 -5160 12558 -5126
rect 12592 -5160 12642 -5126
rect 12676 -5160 12739 -5126
rect 12804 -5160 12836 -5126
rect 12870 -5160 12942 -5126
rect 12976 -5160 12992 -5126
rect 12546 -5166 12752 -5160
rect 12548 -5170 12752 -5166
rect 12804 -5170 12992 -5160
rect 13026 -5130 13684 -5096
rect 13718 -5130 13737 -5096
rect 13026 -5133 13737 -5130
rect 13026 -5167 13038 -5133
rect 13072 -5167 13737 -5133
rect 13026 -5172 13737 -5167
rect 15236 -5084 15294 -5078
rect 15329 -5084 15387 -5078
rect 15236 -5118 15248 -5084
rect 15282 -5118 15341 -5084
rect 15375 -5118 15394 -5084
rect 15236 -5160 15394 -5118
rect 13026 -5173 13084 -5172
rect 15236 -5179 16946 -5160
rect 15236 -5180 15340 -5179
rect 15236 -5214 15248 -5180
rect 15282 -5213 15340 -5180
rect 15374 -5200 16946 -5179
rect 15374 -5213 15394 -5200
rect 15282 -5214 15394 -5213
rect 15236 -5220 15294 -5214
rect 15328 -5219 15386 -5214
rect 7161 -5265 11181 -5259
rect 7155 -5317 7165 -5265
rect 7217 -5268 11181 -5265
rect 7217 -5317 11118 -5268
rect 7161 -5320 11118 -5317
rect 11170 -5320 11181 -5268
rect 7161 -5321 11181 -5320
rect -3193 -5435 16946 -5404
rect -3193 -5469 -2968 -5435
rect -2934 -5469 -2876 -5435
rect -2842 -5469 -2784 -5435
rect -2750 -5469 -2692 -5435
rect -2658 -5469 -2600 -5435
rect -2566 -5469 -2508 -5435
rect -2474 -5469 -2416 -5435
rect -2382 -5469 -2324 -5435
rect -2290 -5469 -2232 -5435
rect -2198 -5469 -2140 -5435
rect -2106 -5469 -2048 -5435
rect -2014 -5469 -1956 -5435
rect -1922 -5469 -1864 -5435
rect -1830 -5469 -1772 -5435
rect -1738 -5469 -1680 -5435
rect -1646 -5469 -1588 -5435
rect -1554 -5469 -1496 -5435
rect -1462 -5469 -1404 -5435
rect -1370 -5469 -1312 -5435
rect -1278 -5469 -1220 -5435
rect -1186 -5469 -1128 -5435
rect -1094 -5469 -1036 -5435
rect -1002 -5469 -944 -5435
rect -910 -5469 -852 -5435
rect -818 -5469 -760 -5435
rect -726 -5469 -668 -5435
rect -634 -5469 -576 -5435
rect -542 -5469 -484 -5435
rect -450 -5469 -392 -5435
rect -358 -5469 -300 -5435
rect -266 -5469 -208 -5435
rect -174 -5469 -116 -5435
rect -82 -5469 -24 -5435
rect 10 -5469 68 -5435
rect 102 -5469 160 -5435
rect 194 -5469 252 -5435
rect 286 -5469 344 -5435
rect 378 -5469 436 -5435
rect 470 -5469 528 -5435
rect 562 -5469 620 -5435
rect 654 -5469 712 -5435
rect 746 -5469 804 -5435
rect 838 -5469 896 -5435
rect 930 -5469 988 -5435
rect 1022 -5469 1080 -5435
rect 1114 -5469 1172 -5435
rect 1206 -5469 1264 -5435
rect 1298 -5469 1356 -5435
rect 1390 -5469 1448 -5435
rect 1482 -5469 1540 -5435
rect 1574 -5469 1632 -5435
rect 1666 -5469 1724 -5435
rect 1758 -5469 1816 -5435
rect 1850 -5469 1908 -5435
rect 1942 -5469 2000 -5435
rect 2034 -5469 2092 -5435
rect 2126 -5469 2184 -5435
rect 2218 -5469 2276 -5435
rect 2310 -5469 2368 -5435
rect 2402 -5469 2460 -5435
rect 2494 -5469 2552 -5435
rect 2586 -5469 2644 -5435
rect 2678 -5469 2736 -5435
rect 2770 -5469 2828 -5435
rect 2862 -5469 2920 -5435
rect 2954 -5469 3012 -5435
rect 3046 -5469 3104 -5435
rect 3138 -5469 3196 -5435
rect 3230 -5469 3288 -5435
rect 3322 -5469 3380 -5435
rect 3414 -5469 3472 -5435
rect 3506 -5469 3564 -5435
rect 3598 -5469 3656 -5435
rect 3690 -5469 3748 -5435
rect 3782 -5469 3840 -5435
rect 3874 -5469 3932 -5435
rect 3966 -5469 4024 -5435
rect 4058 -5469 4116 -5435
rect 4150 -5469 4208 -5435
rect 4242 -5469 4300 -5435
rect 4334 -5469 4392 -5435
rect 4426 -5469 4484 -5435
rect 4518 -5469 4576 -5435
rect 4610 -5469 4668 -5435
rect 4702 -5469 4760 -5435
rect 4794 -5469 4852 -5435
rect 4886 -5469 4944 -5435
rect 4978 -5469 5036 -5435
rect 5070 -5469 5128 -5435
rect 5162 -5469 5220 -5435
rect 5254 -5469 5312 -5435
rect 5346 -5469 5404 -5435
rect 5438 -5469 5496 -5435
rect 5530 -5469 5588 -5435
rect 5622 -5469 5680 -5435
rect 5714 -5469 5772 -5435
rect 5806 -5469 5864 -5435
rect 5898 -5469 5956 -5435
rect 5990 -5469 6048 -5435
rect 6082 -5469 6140 -5435
rect 6174 -5469 6232 -5435
rect 6266 -5469 6324 -5435
rect 6358 -5469 6416 -5435
rect 6450 -5469 6508 -5435
rect 6542 -5469 6600 -5435
rect 6634 -5469 6692 -5435
rect 6726 -5469 6784 -5435
rect 6818 -5469 6876 -5435
rect 6910 -5469 6968 -5435
rect 7002 -5469 7060 -5435
rect 7094 -5469 7152 -5435
rect 7186 -5469 7244 -5435
rect 7278 -5469 7336 -5435
rect 7370 -5469 7428 -5435
rect 7462 -5469 7520 -5435
rect 7554 -5469 7612 -5435
rect 7646 -5469 7704 -5435
rect 7738 -5469 7796 -5435
rect 7830 -5469 7888 -5435
rect 7922 -5469 7980 -5435
rect 8014 -5469 8072 -5435
rect 8106 -5469 8164 -5435
rect 8198 -5469 8256 -5435
rect 8290 -5469 8348 -5435
rect 8382 -5469 8440 -5435
rect 8474 -5469 8532 -5435
rect 8566 -5469 8624 -5435
rect 8658 -5469 8716 -5435
rect 8750 -5469 8808 -5435
rect 8842 -5469 8900 -5435
rect 8934 -5469 8992 -5435
rect 9026 -5469 9084 -5435
rect 9118 -5469 9176 -5435
rect 9210 -5469 9268 -5435
rect 9302 -5469 9360 -5435
rect 9394 -5469 9452 -5435
rect 9486 -5469 9544 -5435
rect 9578 -5469 9636 -5435
rect 9670 -5469 9728 -5435
rect 9762 -5469 9820 -5435
rect 9854 -5469 9912 -5435
rect 9946 -5469 10004 -5435
rect 10038 -5469 10096 -5435
rect 10130 -5469 10188 -5435
rect 10222 -5469 10280 -5435
rect 10314 -5469 10372 -5435
rect 10406 -5469 10464 -5435
rect 10498 -5469 10556 -5435
rect 10590 -5469 10648 -5435
rect 10682 -5469 10740 -5435
rect 10774 -5469 10832 -5435
rect 10866 -5469 10924 -5435
rect 10958 -5469 11016 -5435
rect 11050 -5469 11108 -5435
rect 11142 -5469 11200 -5435
rect 11234 -5469 11292 -5435
rect 11326 -5469 11384 -5435
rect 11418 -5469 11476 -5435
rect 11510 -5469 11568 -5435
rect 11602 -5469 11660 -5435
rect 11694 -5469 11752 -5435
rect 11786 -5469 11844 -5435
rect 11878 -5469 11936 -5435
rect 11970 -5469 12028 -5435
rect 12062 -5469 12120 -5435
rect 12154 -5469 12212 -5435
rect 12246 -5469 12304 -5435
rect 12338 -5469 12396 -5435
rect 12430 -5469 12488 -5435
rect 12522 -5469 12580 -5435
rect 12614 -5469 12672 -5435
rect 12706 -5469 12764 -5435
rect 12798 -5469 12856 -5435
rect 12890 -5469 12948 -5435
rect 12982 -5469 13040 -5435
rect 13074 -5469 13132 -5435
rect 13166 -5469 13224 -5435
rect 13258 -5469 13316 -5435
rect 13350 -5469 13408 -5435
rect 13442 -5469 13500 -5435
rect 13534 -5469 13592 -5435
rect 13626 -5469 13684 -5435
rect 13718 -5469 13776 -5435
rect 13810 -5469 13868 -5435
rect 13902 -5469 13960 -5435
rect 13994 -5469 14052 -5435
rect 14086 -5469 14144 -5435
rect 14178 -5469 14236 -5435
rect 14270 -5469 14328 -5435
rect 14362 -5469 14420 -5435
rect 14454 -5469 14512 -5435
rect 14546 -5469 14604 -5435
rect 14638 -5469 14696 -5435
rect 14730 -5469 14788 -5435
rect 14822 -5469 14880 -5435
rect 14914 -5469 14972 -5435
rect 15006 -5469 15064 -5435
rect 15098 -5469 15156 -5435
rect 15190 -5469 15248 -5435
rect 15282 -5469 15340 -5435
rect 15374 -5469 15432 -5435
rect 15466 -5469 15524 -5435
rect 15558 -5469 15616 -5435
rect 15650 -5469 15708 -5435
rect 15742 -5469 15800 -5435
rect 15834 -5469 15892 -5435
rect 15926 -5469 15984 -5435
rect 16018 -5469 16076 -5435
rect 16110 -5469 16168 -5435
rect 16202 -5469 16260 -5435
rect 16294 -5469 16352 -5435
rect 16386 -5469 16444 -5435
rect 16478 -5469 16536 -5435
rect 16570 -5469 16628 -5435
rect 16662 -5469 16946 -5435
rect -3193 -5500 16946 -5469
rect 11339 -5669 12463 -5665
rect 11338 -5699 12463 -5669
rect 412 -5751 422 -5699
rect 474 -5751 484 -5699
rect 11338 -5724 11586 -5699
rect 12030 -5724 12463 -5699
rect 12522 -5724 12532 -5665
rect 15236 -5694 15294 -5688
rect 15329 -5694 15387 -5688
rect 10725 -5737 10783 -5735
rect 1040 -5738 1098 -5737
rect 3000 -5738 3058 -5737
rect 1040 -5743 3058 -5738
rect 1040 -5777 1052 -5743
rect 1086 -5777 3012 -5743
rect 3046 -5777 3058 -5743
rect 1040 -5782 3058 -5777
rect 1040 -5783 1098 -5782
rect 3000 -5783 3058 -5782
rect 3614 -5738 3672 -5737
rect 5574 -5738 5632 -5737
rect 3614 -5743 5632 -5738
rect 3614 -5777 3626 -5743
rect 3660 -5777 5586 -5743
rect 5620 -5777 5632 -5743
rect 3614 -5782 5632 -5777
rect 3614 -5783 3672 -5782
rect 5574 -5783 5632 -5782
rect 6188 -5738 6246 -5737
rect 8148 -5738 8206 -5737
rect 6188 -5743 8206 -5738
rect 6188 -5777 6200 -5743
rect 6234 -5777 8160 -5743
rect 8194 -5777 8206 -5743
rect 6188 -5782 8206 -5777
rect 6188 -5783 6246 -5782
rect 8148 -5783 8206 -5782
rect 8762 -5738 8820 -5737
rect 10133 -5738 10783 -5737
rect 8762 -5741 10783 -5738
rect 8762 -5743 10737 -5741
rect 8762 -5777 8774 -5743
rect 8808 -5775 10737 -5743
rect 10771 -5775 10783 -5741
rect 8808 -5777 10783 -5775
rect 8762 -5781 10783 -5777
rect 11338 -5740 11430 -5724
rect 15236 -5728 15248 -5694
rect 15282 -5728 15341 -5694
rect 15375 -5704 15394 -5694
rect 15375 -5728 16946 -5704
rect 11338 -5774 11369 -5740
rect 11403 -5774 11430 -5740
rect 11338 -5781 11430 -5774
rect 13669 -5772 13738 -5729
rect 8762 -5782 10231 -5781
rect 8762 -5783 8820 -5782
rect 13669 -5806 13685 -5772
rect 13719 -5806 13738 -5772
rect 13669 -5816 13738 -5806
rect 966 -5818 13738 -5816
rect 966 -5819 12753 -5818
rect 966 -5871 982 -5819
rect 1034 -5870 12753 -5819
rect 12805 -5870 13738 -5818
rect 15236 -5744 16946 -5728
rect 15236 -5789 15394 -5744
rect 15236 -5790 15340 -5789
rect 15236 -5824 15248 -5790
rect 15282 -5823 15340 -5790
rect 15374 -5823 15394 -5789
rect 15282 -5824 15394 -5823
rect 15236 -5830 15294 -5824
rect 15328 -5829 15386 -5824
rect 1034 -5871 13738 -5870
rect 13669 -5873 13738 -5871
rect -3193 -5979 16946 -5948
rect -3193 -6013 -2968 -5979
rect -2934 -6013 -2876 -5979
rect -2842 -6013 -2784 -5979
rect -2750 -6013 -2692 -5979
rect -2658 -6013 -2600 -5979
rect -2566 -6013 -2508 -5979
rect -2474 -6013 -2416 -5979
rect -2382 -6013 -2324 -5979
rect -2290 -6013 -2232 -5979
rect -2198 -6013 -2140 -5979
rect -2106 -6013 -2048 -5979
rect -2014 -6013 -1956 -5979
rect -1922 -6013 -1864 -5979
rect -1830 -6013 -1772 -5979
rect -1738 -6013 -1680 -5979
rect -1646 -6013 -1588 -5979
rect -1554 -6013 -1496 -5979
rect -1462 -6013 -1404 -5979
rect -1370 -6013 -1312 -5979
rect -1278 -6013 -1220 -5979
rect -1186 -6013 -1128 -5979
rect -1094 -6013 -1036 -5979
rect -1002 -6013 -944 -5979
rect -910 -6013 -852 -5979
rect -818 -6013 -760 -5979
rect -726 -6013 -668 -5979
rect -634 -6013 -576 -5979
rect -542 -6013 -484 -5979
rect -450 -6013 -392 -5979
rect -358 -6013 -300 -5979
rect -266 -6013 -208 -5979
rect -174 -6013 -116 -5979
rect -82 -6013 -24 -5979
rect 10 -6013 68 -5979
rect 102 -6013 160 -5979
rect 194 -6013 252 -5979
rect 286 -6013 344 -5979
rect 378 -6013 436 -5979
rect 470 -6013 528 -5979
rect 562 -6013 620 -5979
rect 654 -6013 712 -5979
rect 746 -6013 804 -5979
rect 838 -6013 896 -5979
rect 930 -6013 988 -5979
rect 1022 -6013 1080 -5979
rect 1114 -6013 1172 -5979
rect 1206 -6013 1264 -5979
rect 1298 -6013 1356 -5979
rect 1390 -6013 1448 -5979
rect 1482 -6013 1540 -5979
rect 1574 -6013 1632 -5979
rect 1666 -6013 1724 -5979
rect 1758 -6013 1816 -5979
rect 1850 -6013 1908 -5979
rect 1942 -6013 2000 -5979
rect 2034 -6013 2092 -5979
rect 2126 -6013 2184 -5979
rect 2218 -6013 2276 -5979
rect 2310 -6013 2368 -5979
rect 2402 -6013 2460 -5979
rect 2494 -6013 2552 -5979
rect 2586 -6013 2644 -5979
rect 2678 -6013 2736 -5979
rect 2770 -6013 2828 -5979
rect 2862 -6013 2920 -5979
rect 2954 -6013 3012 -5979
rect 3046 -6013 3104 -5979
rect 3138 -6013 3196 -5979
rect 3230 -6013 3288 -5979
rect 3322 -6013 3380 -5979
rect 3414 -6013 3472 -5979
rect 3506 -6013 3564 -5979
rect 3598 -6013 3656 -5979
rect 3690 -6013 3748 -5979
rect 3782 -6013 3840 -5979
rect 3874 -6013 3932 -5979
rect 3966 -6013 4024 -5979
rect 4058 -6013 4116 -5979
rect 4150 -6013 4208 -5979
rect 4242 -6013 4300 -5979
rect 4334 -6013 4392 -5979
rect 4426 -6013 4484 -5979
rect 4518 -6013 4576 -5979
rect 4610 -6013 4668 -5979
rect 4702 -6013 4760 -5979
rect 4794 -6013 4852 -5979
rect 4886 -6013 4944 -5979
rect 4978 -6013 5036 -5979
rect 5070 -6013 5128 -5979
rect 5162 -6013 5220 -5979
rect 5254 -6013 5312 -5979
rect 5346 -6013 5404 -5979
rect 5438 -6013 5496 -5979
rect 5530 -6013 5588 -5979
rect 5622 -6013 5680 -5979
rect 5714 -6013 5772 -5979
rect 5806 -6013 5864 -5979
rect 5898 -6013 5956 -5979
rect 5990 -6013 6048 -5979
rect 6082 -6013 6140 -5979
rect 6174 -6013 6232 -5979
rect 6266 -6013 6324 -5979
rect 6358 -6013 6416 -5979
rect 6450 -6013 6508 -5979
rect 6542 -6013 6600 -5979
rect 6634 -6013 6692 -5979
rect 6726 -6013 6784 -5979
rect 6818 -6013 6876 -5979
rect 6910 -6013 6968 -5979
rect 7002 -6013 7060 -5979
rect 7094 -6013 7152 -5979
rect 7186 -6013 7244 -5979
rect 7278 -6013 7336 -5979
rect 7370 -6013 7428 -5979
rect 7462 -6013 7520 -5979
rect 7554 -6013 7612 -5979
rect 7646 -6013 7704 -5979
rect 7738 -6013 7796 -5979
rect 7830 -6013 7888 -5979
rect 7922 -6013 7980 -5979
rect 8014 -6013 8072 -5979
rect 8106 -6013 8164 -5979
rect 8198 -6013 8256 -5979
rect 8290 -6013 8348 -5979
rect 8382 -6013 8440 -5979
rect 8474 -6013 8532 -5979
rect 8566 -6013 8624 -5979
rect 8658 -6013 8716 -5979
rect 8750 -6013 8808 -5979
rect 8842 -6013 8900 -5979
rect 8934 -6013 8992 -5979
rect 9026 -6013 9084 -5979
rect 9118 -6013 9176 -5979
rect 9210 -6013 9268 -5979
rect 9302 -6013 9360 -5979
rect 9394 -6013 9452 -5979
rect 9486 -6013 9544 -5979
rect 9578 -6013 9636 -5979
rect 9670 -6013 9728 -5979
rect 9762 -6013 9820 -5979
rect 9854 -6013 9912 -5979
rect 9946 -6013 10004 -5979
rect 10038 -6013 10096 -5979
rect 10130 -6013 10188 -5979
rect 10222 -6013 10280 -5979
rect 10314 -6013 10372 -5979
rect 10406 -6013 10464 -5979
rect 10498 -6013 10556 -5979
rect 10590 -6013 10648 -5979
rect 10682 -6013 10740 -5979
rect 10774 -6013 10832 -5979
rect 10866 -6013 10924 -5979
rect 10958 -6013 11016 -5979
rect 11050 -6013 11108 -5979
rect 11142 -6013 11200 -5979
rect 11234 -6013 11292 -5979
rect 11326 -6013 11384 -5979
rect 11418 -6013 11476 -5979
rect 11510 -6013 11568 -5979
rect 11602 -6013 11660 -5979
rect 11694 -6013 11752 -5979
rect 11786 -6013 11844 -5979
rect 11878 -6013 11936 -5979
rect 11970 -6013 12028 -5979
rect 12062 -6013 12120 -5979
rect 12154 -6013 12212 -5979
rect 12246 -6013 12304 -5979
rect 12338 -6013 12396 -5979
rect 12430 -6013 12488 -5979
rect 12522 -6013 12580 -5979
rect 12614 -6013 12672 -5979
rect 12706 -6013 12764 -5979
rect 12798 -6013 12856 -5979
rect 12890 -6013 12948 -5979
rect 12982 -6013 13040 -5979
rect 13074 -6013 13132 -5979
rect 13166 -6013 13224 -5979
rect 13258 -6013 13316 -5979
rect 13350 -6013 13408 -5979
rect 13442 -6013 13500 -5979
rect 13534 -6013 13592 -5979
rect 13626 -6013 13684 -5979
rect 13718 -6013 13776 -5979
rect 13810 -6013 13868 -5979
rect 13902 -6013 13960 -5979
rect 13994 -6013 14052 -5979
rect 14086 -6013 14144 -5979
rect 14178 -6013 14236 -5979
rect 14270 -6013 14328 -5979
rect 14362 -6013 14420 -5979
rect 14454 -6013 14512 -5979
rect 14546 -6013 14604 -5979
rect 14638 -6013 14696 -5979
rect 14730 -6013 14788 -5979
rect 14822 -6013 14880 -5979
rect 14914 -6013 14972 -5979
rect 15006 -6013 15064 -5979
rect 15098 -6013 15156 -5979
rect 15190 -6013 15248 -5979
rect 15282 -6013 15340 -5979
rect 15374 -6013 15432 -5979
rect 15466 -6013 15524 -5979
rect 15558 -6013 15616 -5979
rect 15650 -6013 15708 -5979
rect 15742 -6013 15800 -5979
rect 15834 -6013 15892 -5979
rect 15926 -6013 15984 -5979
rect 16018 -6013 16076 -5979
rect 16110 -6013 16168 -5979
rect 16202 -6013 16260 -5979
rect 16294 -6013 16352 -5979
rect 16386 -6013 16444 -5979
rect 16478 -6013 16536 -5979
rect 16570 -6013 16628 -5979
rect 16662 -6013 16946 -5979
rect -3193 -6044 16946 -6013
rect 1070 -6078 1116 -6074
rect -862 -6106 13 -6100
rect -862 -6140 -848 -6106
rect -814 -6140 -769 -6106
rect -735 -6140 13 -6106
rect -862 -6149 13 -6140
rect 1064 -6133 1122 -6078
rect 418 -6147 485 -6143
rect 1064 -6147 1076 -6133
rect -57 -6205 12 -6149
rect 418 -6167 1076 -6147
rect 1110 -6167 1122 -6133
rect 418 -6173 1122 -6167
rect -57 -6206 16 -6205
rect 94 -6206 152 -6205
rect 227 -6206 389 -6205
rect -954 -6263 -944 -6207
rect -886 -6263 -876 -6207
rect -782 -6263 -772 -6207
rect -714 -6263 -704 -6207
rect -57 -6211 389 -6206
rect -57 -6245 -30 -6211
rect 4 -6245 106 -6211
rect 140 -6245 242 -6211
rect 276 -6245 389 -6211
rect -57 -6254 389 -6245
rect 418 -6207 434 -6173
rect 468 -6175 1122 -6173
rect 468 -6207 982 -6175
rect 418 -6227 982 -6207
rect 1034 -6206 1122 -6175
rect 1034 -6227 1076 -6206
rect 418 -6240 1076 -6227
rect 1110 -6240 1122 -6206
rect 308 -6340 387 -6254
rect 418 -6258 1122 -6240
rect 1153 -6206 1310 -6146
rect 1153 -6212 2449 -6206
rect 1153 -6246 1171 -6212
rect 1205 -6246 1263 -6212
rect 1297 -6217 2449 -6212
rect 1297 -6246 2369 -6217
rect 1153 -6251 2369 -6246
rect 2403 -6251 2449 -6217
rect 1153 -6268 2449 -6251
rect 2994 -6216 6963 -6199
rect 2994 -6250 3015 -6216
rect 3049 -6250 6876 -6216
rect 6910 -6250 6963 -6216
rect 1153 -6269 1310 -6268
rect 2994 -6270 6963 -6250
rect 7509 -6215 8255 -6197
rect 7509 -6216 8164 -6215
rect 7509 -6250 7522 -6216
rect 7556 -6249 8164 -6216
rect 8198 -6249 8255 -6215
rect 7556 -6250 8255 -6249
rect 7509 -6271 8255 -6250
rect 8799 -6217 9545 -6198
rect 8799 -6251 8811 -6217
rect 8845 -6251 9453 -6217
rect 9487 -6251 9545 -6217
rect 8799 -6269 9545 -6251
rect 10086 -6210 11058 -6204
rect 10086 -6216 11063 -6210
rect 10086 -6217 10925 -6216
rect 10086 -6218 10741 -6217
rect 10086 -6252 10099 -6218
rect 10133 -6251 10741 -6218
rect 10775 -6251 10832 -6217
rect 10866 -6250 10925 -6217
rect 10959 -6250 11017 -6216
rect 11051 -6250 11063 -6216
rect 11233 -6219 11418 -6211
rect 10866 -6251 11063 -6250
rect 10133 -6252 11063 -6251
rect 10086 -6256 11063 -6252
rect 10086 -6274 11058 -6256
rect 11110 -6293 11120 -6241
rect 11172 -6293 11182 -6241
rect 11233 -6253 11250 -6219
rect 11284 -6253 11344 -6219
rect 11378 -6253 11418 -6219
rect 11233 -6340 11418 -6253
rect 14617 -6274 14627 -6219
rect 14682 -6226 14692 -6219
rect 15824 -6226 15834 -6219
rect 14682 -6266 15834 -6226
rect 14682 -6274 14692 -6266
rect 15824 -6274 15834 -6266
rect 15889 -6274 15899 -6219
rect -1281 -6409 -1271 -6353
rect -1213 -6356 -1203 -6353
rect -1213 -6409 -768 -6356
rect -715 -6409 -705 -6356
rect -1267 -6410 -705 -6409
rect 308 -6425 11419 -6340
rect -3193 -6523 16946 -6492
rect -3193 -6557 -2968 -6523
rect -2934 -6557 -2876 -6523
rect -2842 -6557 -2784 -6523
rect -2750 -6557 -2692 -6523
rect -2658 -6557 -2600 -6523
rect -2566 -6557 -2508 -6523
rect -2474 -6557 -2416 -6523
rect -2382 -6557 -2324 -6523
rect -2290 -6557 -2232 -6523
rect -2198 -6557 -2140 -6523
rect -2106 -6557 -2048 -6523
rect -2014 -6557 -1956 -6523
rect -1922 -6557 -1864 -6523
rect -1830 -6557 -1772 -6523
rect -1738 -6557 -1680 -6523
rect -1646 -6557 -1588 -6523
rect -1554 -6557 -1496 -6523
rect -1462 -6557 -1404 -6523
rect -1370 -6557 -1312 -6523
rect -1278 -6557 -1220 -6523
rect -1186 -6557 -1128 -6523
rect -1094 -6557 -1036 -6523
rect -1002 -6557 -944 -6523
rect -910 -6557 -852 -6523
rect -818 -6557 -760 -6523
rect -726 -6557 -668 -6523
rect -634 -6557 -576 -6523
rect -542 -6557 -484 -6523
rect -450 -6557 -392 -6523
rect -358 -6557 -300 -6523
rect -266 -6557 -208 -6523
rect -174 -6557 -116 -6523
rect -82 -6557 -24 -6523
rect 10 -6557 68 -6523
rect 102 -6557 160 -6523
rect 194 -6557 252 -6523
rect 286 -6557 344 -6523
rect 378 -6557 436 -6523
rect 470 -6557 528 -6523
rect 562 -6557 620 -6523
rect 654 -6557 712 -6523
rect 746 -6557 804 -6523
rect 838 -6557 896 -6523
rect 930 -6557 988 -6523
rect 1022 -6557 1080 -6523
rect 1114 -6557 1172 -6523
rect 1206 -6557 1264 -6523
rect 1298 -6557 1356 -6523
rect 1390 -6557 1448 -6523
rect 1482 -6557 1540 -6523
rect 1574 -6557 1632 -6523
rect 1666 -6557 1724 -6523
rect 1758 -6557 1816 -6523
rect 1850 -6557 1908 -6523
rect 1942 -6557 2000 -6523
rect 2034 -6557 2092 -6523
rect 2126 -6557 2184 -6523
rect 2218 -6557 2276 -6523
rect 2310 -6557 2368 -6523
rect 2402 -6557 2460 -6523
rect 2494 -6557 2552 -6523
rect 2586 -6557 2644 -6523
rect 2678 -6557 2736 -6523
rect 2770 -6557 2828 -6523
rect 2862 -6557 2920 -6523
rect 2954 -6557 3012 -6523
rect 3046 -6557 3104 -6523
rect 3138 -6557 3196 -6523
rect 3230 -6557 3288 -6523
rect 3322 -6557 3380 -6523
rect 3414 -6557 3472 -6523
rect 3506 -6557 3564 -6523
rect 3598 -6557 3656 -6523
rect 3690 -6557 3748 -6523
rect 3782 -6557 3840 -6523
rect 3874 -6557 3932 -6523
rect 3966 -6557 4024 -6523
rect 4058 -6557 4116 -6523
rect 4150 -6557 4208 -6523
rect 4242 -6557 4300 -6523
rect 4334 -6557 4392 -6523
rect 4426 -6557 4484 -6523
rect 4518 -6557 4576 -6523
rect 4610 -6557 4668 -6523
rect 4702 -6557 4760 -6523
rect 4794 -6557 4852 -6523
rect 4886 -6557 4944 -6523
rect 4978 -6557 5036 -6523
rect 5070 -6557 5128 -6523
rect 5162 -6557 5220 -6523
rect 5254 -6557 5312 -6523
rect 5346 -6557 5404 -6523
rect 5438 -6557 5496 -6523
rect 5530 -6557 5588 -6523
rect 5622 -6557 5680 -6523
rect 5714 -6557 5772 -6523
rect 5806 -6557 5864 -6523
rect 5898 -6557 5956 -6523
rect 5990 -6557 6048 -6523
rect 6082 -6557 6140 -6523
rect 6174 -6557 6232 -6523
rect 6266 -6557 6324 -6523
rect 6358 -6557 6416 -6523
rect 6450 -6557 6508 -6523
rect 6542 -6557 6600 -6523
rect 6634 -6557 6692 -6523
rect 6726 -6557 6784 -6523
rect 6818 -6557 6876 -6523
rect 6910 -6557 6968 -6523
rect 7002 -6557 7060 -6523
rect 7094 -6557 7152 -6523
rect 7186 -6557 7244 -6523
rect 7278 -6557 7336 -6523
rect 7370 -6557 7428 -6523
rect 7462 -6557 7520 -6523
rect 7554 -6557 7612 -6523
rect 7646 -6557 7704 -6523
rect 7738 -6557 7796 -6523
rect 7830 -6557 7888 -6523
rect 7922 -6557 7980 -6523
rect 8014 -6557 8072 -6523
rect 8106 -6557 8164 -6523
rect 8198 -6557 8256 -6523
rect 8290 -6557 8348 -6523
rect 8382 -6557 8440 -6523
rect 8474 -6557 8532 -6523
rect 8566 -6557 8624 -6523
rect 8658 -6557 8716 -6523
rect 8750 -6557 8808 -6523
rect 8842 -6557 8900 -6523
rect 8934 -6557 8992 -6523
rect 9026 -6557 9084 -6523
rect 9118 -6557 9176 -6523
rect 9210 -6557 9268 -6523
rect 9302 -6557 9360 -6523
rect 9394 -6557 9452 -6523
rect 9486 -6557 9544 -6523
rect 9578 -6557 9636 -6523
rect 9670 -6557 9728 -6523
rect 9762 -6557 9820 -6523
rect 9854 -6557 9912 -6523
rect 9946 -6557 10004 -6523
rect 10038 -6557 10096 -6523
rect 10130 -6557 10188 -6523
rect 10222 -6557 10280 -6523
rect 10314 -6557 10372 -6523
rect 10406 -6557 10464 -6523
rect 10498 -6557 10556 -6523
rect 10590 -6557 10648 -6523
rect 10682 -6557 10740 -6523
rect 10774 -6557 10832 -6523
rect 10866 -6557 10924 -6523
rect 10958 -6557 11016 -6523
rect 11050 -6557 11108 -6523
rect 11142 -6557 11200 -6523
rect 11234 -6557 11292 -6523
rect 11326 -6557 11384 -6523
rect 11418 -6557 11476 -6523
rect 11510 -6557 11568 -6523
rect 11602 -6557 11660 -6523
rect 11694 -6557 11752 -6523
rect 11786 -6557 11844 -6523
rect 11878 -6557 11936 -6523
rect 11970 -6557 12028 -6523
rect 12062 -6557 12120 -6523
rect 12154 -6557 12212 -6523
rect 12246 -6557 12304 -6523
rect 12338 -6557 12396 -6523
rect 12430 -6557 12488 -6523
rect 12522 -6557 12580 -6523
rect 12614 -6557 12672 -6523
rect 12706 -6557 12764 -6523
rect 12798 -6557 12856 -6523
rect 12890 -6557 12948 -6523
rect 12982 -6557 13040 -6523
rect 13074 -6557 13132 -6523
rect 13166 -6557 13224 -6523
rect 13258 -6557 13316 -6523
rect 13350 -6557 13408 -6523
rect 13442 -6557 13500 -6523
rect 13534 -6557 13592 -6523
rect 13626 -6557 13684 -6523
rect 13718 -6557 13776 -6523
rect 13810 -6557 13868 -6523
rect 13902 -6557 13960 -6523
rect 13994 -6557 14052 -6523
rect 14086 -6557 14144 -6523
rect 14178 -6557 14236 -6523
rect 14270 -6557 14328 -6523
rect 14362 -6557 14420 -6523
rect 14454 -6557 14512 -6523
rect 14546 -6557 14604 -6523
rect 14638 -6557 14696 -6523
rect 14730 -6557 14788 -6523
rect 14822 -6557 14880 -6523
rect 14914 -6557 14972 -6523
rect 15006 -6557 15064 -6523
rect 15098 -6557 15156 -6523
rect 15190 -6557 15248 -6523
rect 15282 -6557 15340 -6523
rect 15374 -6557 15432 -6523
rect 15466 -6557 15524 -6523
rect 15558 -6557 15616 -6523
rect 15650 -6557 15708 -6523
rect 15742 -6557 15800 -6523
rect 15834 -6557 15892 -6523
rect 15926 -6557 15984 -6523
rect 16018 -6557 16076 -6523
rect 16110 -6557 16168 -6523
rect 16202 -6557 16260 -6523
rect 16294 -6557 16352 -6523
rect 16386 -6557 16444 -6523
rect 16478 -6557 16536 -6523
rect 16570 -6557 16628 -6523
rect 16662 -6557 16946 -6523
rect -3193 -6588 16946 -6557
rect -787 -6671 7349 -6670
rect -2515 -6693 -2457 -6687
rect -2515 -6727 -2503 -6693
rect -2469 -6696 -2457 -6693
rect -2095 -6693 -2037 -6687
rect -2095 -6696 -2083 -6693
rect -2469 -6724 -2083 -6696
rect -2469 -6727 -2457 -6724
rect -2515 -6733 -2457 -6727
rect -2095 -6727 -2083 -6724
rect -2049 -6696 -2037 -6693
rect -1781 -6693 -1723 -6687
rect -1781 -6696 -1769 -6693
rect -2049 -6724 -1769 -6696
rect -2049 -6727 -2037 -6724
rect -2095 -6733 -2037 -6727
rect -1781 -6727 -1769 -6724
rect -1735 -6727 -1723 -6693
rect -1781 -6733 -1723 -6727
rect -787 -6727 -772 -6671
rect -714 -6726 7349 -6671
rect 7407 -6726 7417 -6670
rect -714 -6727 7403 -6726
rect -787 -6728 7403 -6727
rect -2436 -6761 -2378 -6755
rect -2436 -6795 -2424 -6761
rect -2390 -6764 -2378 -6761
rect -2198 -6761 -2140 -6755
rect -2198 -6764 -2186 -6761
rect -2390 -6792 -2186 -6764
rect -2390 -6795 -2378 -6792
rect -2436 -6801 -2378 -6795
rect -2198 -6795 -2186 -6792
rect -2152 -6764 -2140 -6761
rect -1694 -6761 -1636 -6755
rect -1694 -6764 -1682 -6761
rect -2152 -6792 -1682 -6764
rect -2152 -6795 -2140 -6792
rect -2198 -6801 -2140 -6795
rect -1694 -6795 -1682 -6792
rect -1648 -6795 -1636 -6761
rect -1694 -6801 -1636 -6795
rect -2617 -6824 -2607 -6821
rect -3193 -6870 -2607 -6824
rect -2617 -6873 -2607 -6870
rect -2554 -6873 -2544 -6821
rect 5018 -6840 5028 -6786
rect 5082 -6840 13925 -6786
rect 13979 -6840 13989 -6786
rect -2356 -6875 -2299 -6868
rect -952 -6875 -894 -6874
rect -2356 -6880 -894 -6875
rect -2356 -6882 -940 -6880
rect -2356 -6916 -2343 -6882
rect -2309 -6914 -940 -6882
rect -906 -6914 -894 -6880
rect -2309 -6916 -894 -6914
rect -2356 -6917 -894 -6916
rect -2356 -6923 -2299 -6917
rect -952 -6920 -894 -6917
rect -1978 -7003 -1968 -6951
rect -1915 -6954 -1908 -6951
rect -1915 -6960 -1183 -6954
rect -415 -6958 -405 -6899
rect -346 -6958 3736 -6899
rect 3795 -6958 3805 -6899
rect -1915 -6994 -1233 -6960
rect -1199 -6994 -1183 -6960
rect 4934 -6977 4945 -6923
rect 4999 -6977 15832 -6923
rect 15886 -6977 15896 -6923
rect -1915 -7000 -1183 -6994
rect -1915 -7003 -1908 -7000
rect -3193 -7067 16946 -7036
rect -3193 -7101 -2968 -7067
rect -2934 -7101 -2876 -7067
rect -2842 -7101 -2784 -7067
rect -2750 -7101 -2692 -7067
rect -2658 -7101 -2600 -7067
rect -2566 -7101 -2508 -7067
rect -2474 -7101 -2416 -7067
rect -2382 -7101 -2324 -7067
rect -2290 -7101 -2232 -7067
rect -2198 -7101 -2140 -7067
rect -2106 -7101 -2048 -7067
rect -2014 -7101 -1956 -7067
rect -1922 -7101 -1864 -7067
rect -1830 -7101 -1772 -7067
rect -1738 -7101 -1680 -7067
rect -1646 -7101 -1588 -7067
rect -1554 -7101 -1496 -7067
rect -1462 -7101 -1404 -7067
rect -1370 -7101 -1312 -7067
rect -1278 -7101 -1220 -7067
rect -1186 -7101 -1128 -7067
rect -1094 -7101 -1036 -7067
rect -1002 -7101 -944 -7067
rect -910 -7101 -852 -7067
rect -818 -7101 -760 -7067
rect -726 -7101 -668 -7067
rect -634 -7101 -576 -7067
rect -542 -7101 -484 -7067
rect -450 -7101 -392 -7067
rect -358 -7101 -300 -7067
rect -266 -7101 -208 -7067
rect -174 -7101 -116 -7067
rect -82 -7101 -24 -7067
rect 10 -7101 68 -7067
rect 102 -7101 160 -7067
rect 194 -7101 252 -7067
rect 286 -7101 344 -7067
rect 378 -7101 436 -7067
rect 470 -7101 528 -7067
rect 562 -7101 620 -7067
rect 654 -7101 712 -7067
rect 746 -7101 804 -7067
rect 838 -7101 896 -7067
rect 930 -7101 988 -7067
rect 1022 -7101 1080 -7067
rect 1114 -7101 1172 -7067
rect 1206 -7101 1264 -7067
rect 1298 -7101 1356 -7067
rect 1390 -7101 1448 -7067
rect 1482 -7101 1540 -7067
rect 1574 -7101 1632 -7067
rect 1666 -7101 1724 -7067
rect 1758 -7101 1816 -7067
rect 1850 -7101 1908 -7067
rect 1942 -7101 2000 -7067
rect 2034 -7101 2092 -7067
rect 2126 -7101 2184 -7067
rect 2218 -7101 2276 -7067
rect 2310 -7101 2368 -7067
rect 2402 -7101 2460 -7067
rect 2494 -7101 2552 -7067
rect 2586 -7101 2644 -7067
rect 2678 -7101 2736 -7067
rect 2770 -7101 2828 -7067
rect 2862 -7101 2920 -7067
rect 2954 -7101 3012 -7067
rect 3046 -7101 3104 -7067
rect 3138 -7101 3196 -7067
rect 3230 -7101 3288 -7067
rect 3322 -7101 3380 -7067
rect 3414 -7101 3472 -7067
rect 3506 -7101 3564 -7067
rect 3598 -7101 3656 -7067
rect 3690 -7101 3748 -7067
rect 3782 -7101 3840 -7067
rect 3874 -7101 3932 -7067
rect 3966 -7101 4024 -7067
rect 4058 -7101 4116 -7067
rect 4150 -7101 4208 -7067
rect 4242 -7101 4300 -7067
rect 4334 -7101 4392 -7067
rect 4426 -7101 4484 -7067
rect 4518 -7101 4576 -7067
rect 4610 -7101 4668 -7067
rect 4702 -7101 4760 -7067
rect 4794 -7101 4852 -7067
rect 4886 -7101 4944 -7067
rect 4978 -7101 5036 -7067
rect 5070 -7101 5128 -7067
rect 5162 -7101 5220 -7067
rect 5254 -7101 5312 -7067
rect 5346 -7101 5404 -7067
rect 5438 -7101 5496 -7067
rect 5530 -7101 5588 -7067
rect 5622 -7101 5680 -7067
rect 5714 -7101 5772 -7067
rect 5806 -7101 5864 -7067
rect 5898 -7101 5956 -7067
rect 5990 -7101 6048 -7067
rect 6082 -7101 6140 -7067
rect 6174 -7101 6232 -7067
rect 6266 -7101 6324 -7067
rect 6358 -7101 6416 -7067
rect 6450 -7101 6508 -7067
rect 6542 -7101 6600 -7067
rect 6634 -7101 6692 -7067
rect 6726 -7101 6784 -7067
rect 6818 -7101 6876 -7067
rect 6910 -7101 6968 -7067
rect 7002 -7101 7060 -7067
rect 7094 -7101 7152 -7067
rect 7186 -7101 7244 -7067
rect 7278 -7101 7336 -7067
rect 7370 -7101 7428 -7067
rect 7462 -7101 7520 -7067
rect 7554 -7101 7612 -7067
rect 7646 -7101 7704 -7067
rect 7738 -7101 7796 -7067
rect 7830 -7101 7888 -7067
rect 7922 -7101 7980 -7067
rect 8014 -7101 8072 -7067
rect 8106 -7101 8164 -7067
rect 8198 -7101 8256 -7067
rect 8290 -7101 8348 -7067
rect 8382 -7101 8440 -7067
rect 8474 -7101 8532 -7067
rect 8566 -7101 8624 -7067
rect 8658 -7101 8716 -7067
rect 8750 -7101 8808 -7067
rect 8842 -7101 8900 -7067
rect 8934 -7101 8992 -7067
rect 9026 -7101 9084 -7067
rect 9118 -7101 9176 -7067
rect 9210 -7101 9268 -7067
rect 9302 -7101 9360 -7067
rect 9394 -7101 9452 -7067
rect 9486 -7101 9544 -7067
rect 9578 -7101 9636 -7067
rect 9670 -7101 9728 -7067
rect 9762 -7101 9820 -7067
rect 9854 -7101 9912 -7067
rect 9946 -7101 10004 -7067
rect 10038 -7101 10096 -7067
rect 10130 -7101 10188 -7067
rect 10222 -7101 10280 -7067
rect 10314 -7101 10372 -7067
rect 10406 -7101 10464 -7067
rect 10498 -7101 10556 -7067
rect 10590 -7101 10648 -7067
rect 10682 -7101 10740 -7067
rect 10774 -7101 10832 -7067
rect 10866 -7101 10924 -7067
rect 10958 -7101 11016 -7067
rect 11050 -7101 11108 -7067
rect 11142 -7101 11200 -7067
rect 11234 -7101 11292 -7067
rect 11326 -7101 11384 -7067
rect 11418 -7101 11476 -7067
rect 11510 -7101 11568 -7067
rect 11602 -7101 11660 -7067
rect 11694 -7101 11752 -7067
rect 11786 -7101 11844 -7067
rect 11878 -7101 11936 -7067
rect 11970 -7101 12028 -7067
rect 12062 -7101 12120 -7067
rect 12154 -7101 12212 -7067
rect 12246 -7101 12304 -7067
rect 12338 -7101 12396 -7067
rect 12430 -7101 12488 -7067
rect 12522 -7101 12580 -7067
rect 12614 -7101 12672 -7067
rect 12706 -7101 12764 -7067
rect 12798 -7101 12856 -7067
rect 12890 -7101 12948 -7067
rect 12982 -7101 13040 -7067
rect 13074 -7101 13132 -7067
rect 13166 -7101 13224 -7067
rect 13258 -7101 13316 -7067
rect 13350 -7101 13408 -7067
rect 13442 -7101 13500 -7067
rect 13534 -7101 13592 -7067
rect 13626 -7101 13684 -7067
rect 13718 -7101 13776 -7067
rect 13810 -7101 13868 -7067
rect 13902 -7101 13960 -7067
rect 13994 -7101 14052 -7067
rect 14086 -7101 14144 -7067
rect 14178 -7101 14236 -7067
rect 14270 -7101 14328 -7067
rect 14362 -7101 14420 -7067
rect 14454 -7101 14512 -7067
rect 14546 -7101 14604 -7067
rect 14638 -7101 14696 -7067
rect 14730 -7101 14788 -7067
rect 14822 -7101 14880 -7067
rect 14914 -7101 14972 -7067
rect 15006 -7101 15064 -7067
rect 15098 -7101 15156 -7067
rect 15190 -7101 15248 -7067
rect 15282 -7101 15340 -7067
rect 15374 -7101 15432 -7067
rect 15466 -7101 15524 -7067
rect 15558 -7101 15616 -7067
rect 15650 -7101 15708 -7067
rect 15742 -7101 15800 -7067
rect 15834 -7101 15892 -7067
rect 15926 -7101 15984 -7067
rect 16018 -7101 16076 -7067
rect 16110 -7101 16168 -7067
rect 16202 -7101 16260 -7067
rect 16294 -7101 16352 -7067
rect 16386 -7101 16444 -7067
rect 16478 -7101 16536 -7067
rect 16570 -7101 16628 -7067
rect 16662 -7101 16946 -7067
rect -3193 -7132 16946 -7101
rect 5736 -7180 6293 -7173
rect 3840 -7185 3898 -7182
rect 3099 -7188 3898 -7185
rect 3099 -7191 3852 -7188
rect 3099 -7225 3111 -7191
rect 3145 -7222 3852 -7191
rect 3886 -7222 3898 -7188
rect 3145 -7225 3898 -7222
rect 3099 -7228 3898 -7225
rect 3099 -7230 3872 -7228
rect 3099 -7231 3157 -7230
rect 4935 -7249 4945 -7195
rect 4999 -7249 5009 -7195
rect 5736 -7214 6245 -7180
rect 6279 -7214 6293 -7180
rect 5736 -7220 6293 -7214
rect 2724 -7317 2736 -7258
rect 2795 -7270 2991 -7258
rect 2795 -7304 2934 -7270
rect 2968 -7304 2991 -7270
rect 2795 -7317 2991 -7304
rect 2724 -7318 2991 -7317
rect 3726 -7351 3736 -7292
rect 3795 -7351 3805 -7292
rect 4553 -7299 4611 -7298
rect 3906 -7304 4611 -7299
rect 3906 -7305 4565 -7304
rect 3906 -7339 3928 -7305
rect 3962 -7338 4565 -7305
rect 4599 -7338 4611 -7304
rect 3962 -7339 4611 -7338
rect 3906 -7344 4611 -7339
rect 5028 -7299 5082 -7290
rect 3906 -7348 4599 -7344
rect 5028 -7372 5082 -7353
rect 5736 -7367 5783 -7220
rect 7339 -7310 7349 -7254
rect 7407 -7310 7417 -7254
rect 7582 -7267 16044 -7265
rect 7582 -7290 15971 -7267
rect 7582 -7324 7604 -7290
rect 7638 -7324 15971 -7290
rect 7582 -7326 15971 -7324
rect 16030 -7326 16044 -7267
rect 7582 -7330 16044 -7326
rect 7582 -7364 7661 -7330
rect 5131 -7373 5783 -7367
rect 5131 -7407 5171 -7373
rect 5205 -7407 5783 -7373
rect 5131 -7414 5783 -7407
rect 6682 -7373 6740 -7367
rect 6682 -7407 6694 -7373
rect 6728 -7376 6740 -7373
rect 7186 -7373 7244 -7367
rect 7186 -7376 7198 -7373
rect 6728 -7404 7198 -7376
rect 6728 -7407 6740 -7404
rect 6682 -7413 6740 -7407
rect 7186 -7407 7198 -7404
rect 7232 -7376 7244 -7373
rect 7424 -7373 7482 -7367
rect 7424 -7376 7436 -7373
rect 7232 -7404 7436 -7376
rect 7232 -7407 7244 -7404
rect 7186 -7413 7244 -7407
rect 7424 -7407 7436 -7404
rect 7470 -7407 7482 -7373
rect 7424 -7413 7482 -7407
rect 7582 -7398 7605 -7364
rect 7639 -7398 7661 -7364
rect 7582 -7408 7661 -7398
rect -631 -7498 -620 -7439
rect -561 -7498 2736 -7439
rect 2795 -7498 2805 -7439
rect 6769 -7441 6827 -7435
rect 6769 -7475 6781 -7441
rect 6815 -7444 6827 -7441
rect 7083 -7441 7141 -7435
rect 7083 -7444 7095 -7441
rect 6815 -7472 7095 -7444
rect 6815 -7475 6827 -7472
rect 6769 -7481 6827 -7475
rect 7083 -7475 7095 -7472
rect 7129 -7444 7141 -7441
rect 7503 -7441 7561 -7435
rect 7503 -7444 7515 -7441
rect 7129 -7472 7515 -7444
rect 7129 -7475 7141 -7472
rect 7083 -7481 7141 -7475
rect 7503 -7475 7515 -7472
rect 7549 -7475 7561 -7441
rect 7503 -7481 7561 -7475
rect -3193 -7611 16946 -7580
rect -3193 -7645 -2968 -7611
rect -2934 -7645 -2876 -7611
rect -2842 -7645 -2784 -7611
rect -2750 -7645 -2692 -7611
rect -2658 -7645 -2600 -7611
rect -2566 -7645 -2508 -7611
rect -2474 -7645 -2416 -7611
rect -2382 -7645 -2324 -7611
rect -2290 -7645 -2232 -7611
rect -2198 -7645 -2140 -7611
rect -2106 -7645 -2048 -7611
rect -2014 -7645 -1956 -7611
rect -1922 -7645 -1864 -7611
rect -1830 -7645 -1772 -7611
rect -1738 -7645 -1680 -7611
rect -1646 -7645 -1588 -7611
rect -1554 -7645 -1496 -7611
rect -1462 -7645 -1404 -7611
rect -1370 -7645 -1312 -7611
rect -1278 -7645 -1220 -7611
rect -1186 -7645 -1128 -7611
rect -1094 -7645 -1036 -7611
rect -1002 -7645 -944 -7611
rect -910 -7645 -852 -7611
rect -818 -7645 -760 -7611
rect -726 -7645 -668 -7611
rect -634 -7645 -576 -7611
rect -542 -7645 -484 -7611
rect -450 -7645 -392 -7611
rect -358 -7645 -300 -7611
rect -266 -7645 -208 -7611
rect -174 -7645 -116 -7611
rect -82 -7645 -24 -7611
rect 10 -7645 68 -7611
rect 102 -7645 160 -7611
rect 194 -7645 252 -7611
rect 286 -7645 344 -7611
rect 378 -7645 436 -7611
rect 470 -7645 528 -7611
rect 562 -7645 620 -7611
rect 654 -7645 712 -7611
rect 746 -7645 804 -7611
rect 838 -7645 896 -7611
rect 930 -7645 988 -7611
rect 1022 -7645 1080 -7611
rect 1114 -7645 1172 -7611
rect 1206 -7645 1264 -7611
rect 1298 -7645 1356 -7611
rect 1390 -7645 1448 -7611
rect 1482 -7645 1540 -7611
rect 1574 -7645 1632 -7611
rect 1666 -7645 1724 -7611
rect 1758 -7645 1816 -7611
rect 1850 -7645 1908 -7611
rect 1942 -7645 2000 -7611
rect 2034 -7645 2092 -7611
rect 2126 -7645 2184 -7611
rect 2218 -7645 2276 -7611
rect 2310 -7645 2368 -7611
rect 2402 -7645 2460 -7611
rect 2494 -7645 2552 -7611
rect 2586 -7645 2644 -7611
rect 2678 -7645 2736 -7611
rect 2770 -7645 2828 -7611
rect 2862 -7645 2920 -7611
rect 2954 -7645 3012 -7611
rect 3046 -7645 3104 -7611
rect 3138 -7645 3196 -7611
rect 3230 -7645 3288 -7611
rect 3322 -7645 3380 -7611
rect 3414 -7645 3472 -7611
rect 3506 -7645 3564 -7611
rect 3598 -7645 3656 -7611
rect 3690 -7645 3748 -7611
rect 3782 -7645 3840 -7611
rect 3874 -7645 3932 -7611
rect 3966 -7645 4024 -7611
rect 4058 -7645 4116 -7611
rect 4150 -7645 4208 -7611
rect 4242 -7645 4300 -7611
rect 4334 -7645 4392 -7611
rect 4426 -7645 4484 -7611
rect 4518 -7645 4576 -7611
rect 4610 -7645 4668 -7611
rect 4702 -7645 4760 -7611
rect 4794 -7645 4852 -7611
rect 4886 -7645 4944 -7611
rect 4978 -7645 5036 -7611
rect 5070 -7645 5128 -7611
rect 5162 -7645 5220 -7611
rect 5254 -7645 5312 -7611
rect 5346 -7645 5404 -7611
rect 5438 -7645 5496 -7611
rect 5530 -7645 5588 -7611
rect 5622 -7645 5680 -7611
rect 5714 -7645 5772 -7611
rect 5806 -7645 5864 -7611
rect 5898 -7645 5956 -7611
rect 5990 -7645 6048 -7611
rect 6082 -7645 6140 -7611
rect 6174 -7645 6232 -7611
rect 6266 -7645 6324 -7611
rect 6358 -7645 6416 -7611
rect 6450 -7645 6508 -7611
rect 6542 -7645 6600 -7611
rect 6634 -7645 6692 -7611
rect 6726 -7645 6784 -7611
rect 6818 -7645 6876 -7611
rect 6910 -7645 6968 -7611
rect 7002 -7645 7060 -7611
rect 7094 -7645 7152 -7611
rect 7186 -7645 7244 -7611
rect 7278 -7645 7336 -7611
rect 7370 -7645 7428 -7611
rect 7462 -7645 7520 -7611
rect 7554 -7645 7612 -7611
rect 7646 -7645 7704 -7611
rect 7738 -7645 7796 -7611
rect 7830 -7645 7888 -7611
rect 7922 -7645 7980 -7611
rect 8014 -7645 8072 -7611
rect 8106 -7645 8164 -7611
rect 8198 -7645 8256 -7611
rect 8290 -7645 8348 -7611
rect 8382 -7645 8440 -7611
rect 8474 -7645 8532 -7611
rect 8566 -7645 8624 -7611
rect 8658 -7645 8716 -7611
rect 8750 -7645 8808 -7611
rect 8842 -7645 8900 -7611
rect 8934 -7645 8992 -7611
rect 9026 -7645 9084 -7611
rect 9118 -7645 9176 -7611
rect 9210 -7645 9268 -7611
rect 9302 -7645 9360 -7611
rect 9394 -7645 9452 -7611
rect 9486 -7645 9544 -7611
rect 9578 -7645 9636 -7611
rect 9670 -7645 9728 -7611
rect 9762 -7645 9820 -7611
rect 9854 -7645 9912 -7611
rect 9946 -7645 10004 -7611
rect 10038 -7645 10096 -7611
rect 10130 -7645 10188 -7611
rect 10222 -7645 10280 -7611
rect 10314 -7645 10372 -7611
rect 10406 -7645 10464 -7611
rect 10498 -7645 10556 -7611
rect 10590 -7645 10648 -7611
rect 10682 -7645 10740 -7611
rect 10774 -7645 10832 -7611
rect 10866 -7645 10924 -7611
rect 10958 -7645 11016 -7611
rect 11050 -7645 11108 -7611
rect 11142 -7645 11200 -7611
rect 11234 -7645 11292 -7611
rect 11326 -7645 11384 -7611
rect 11418 -7645 11476 -7611
rect 11510 -7645 11568 -7611
rect 11602 -7645 11660 -7611
rect 11694 -7645 11752 -7611
rect 11786 -7645 11844 -7611
rect 11878 -7645 11936 -7611
rect 11970 -7645 12028 -7611
rect 12062 -7645 12120 -7611
rect 12154 -7645 12212 -7611
rect 12246 -7645 12304 -7611
rect 12338 -7645 12396 -7611
rect 12430 -7645 12488 -7611
rect 12522 -7645 12580 -7611
rect 12614 -7645 12672 -7611
rect 12706 -7645 12764 -7611
rect 12798 -7645 12856 -7611
rect 12890 -7645 12948 -7611
rect 12982 -7645 13040 -7611
rect 13074 -7645 13132 -7611
rect 13166 -7645 13224 -7611
rect 13258 -7645 13316 -7611
rect 13350 -7645 13408 -7611
rect 13442 -7645 13500 -7611
rect 13534 -7645 13592 -7611
rect 13626 -7645 13684 -7611
rect 13718 -7645 13776 -7611
rect 13810 -7645 13868 -7611
rect 13902 -7645 13960 -7611
rect 13994 -7645 14052 -7611
rect 14086 -7645 14144 -7611
rect 14178 -7645 14236 -7611
rect 14270 -7645 14328 -7611
rect 14362 -7645 14420 -7611
rect 14454 -7645 14512 -7611
rect 14546 -7645 14604 -7611
rect 14638 -7645 14696 -7611
rect 14730 -7645 14788 -7611
rect 14822 -7645 14880 -7611
rect 14914 -7645 14972 -7611
rect 15006 -7645 15064 -7611
rect 15098 -7645 15156 -7611
rect 15190 -7645 15248 -7611
rect 15282 -7645 15340 -7611
rect 15374 -7645 15432 -7611
rect 15466 -7645 15524 -7611
rect 15558 -7645 15616 -7611
rect 15650 -7645 15708 -7611
rect 15742 -7645 15800 -7611
rect 15834 -7645 15892 -7611
rect 15926 -7645 15984 -7611
rect 16018 -7645 16076 -7611
rect 16110 -7645 16168 -7611
rect 16202 -7645 16260 -7611
rect 16294 -7645 16352 -7611
rect 16386 -7645 16444 -7611
rect 16478 -7645 16536 -7611
rect 16570 -7645 16628 -7611
rect 16662 -7645 16946 -7611
rect -3193 -7676 16946 -7645
rect 308 -7828 11419 -7743
rect -629 -7906 -619 -7902
rect -1978 -7960 -1968 -7908
rect -1915 -7911 -1905 -7908
rect -1915 -7918 -889 -7911
rect -1915 -7952 -937 -7918
rect -903 -7952 -889 -7918
rect -1915 -7958 -889 -7952
rect -781 -7917 -619 -7906
rect -781 -7951 -762 -7917
rect -728 -7951 -619 -7917
rect -781 -7957 -619 -7951
rect -781 -7958 -709 -7957
rect -1915 -7960 -1905 -7958
rect -629 -7961 -619 -7957
rect -560 -7961 -550 -7902
rect 308 -7914 387 -7828
rect 1153 -7900 1310 -7899
rect -57 -7923 389 -7914
rect -57 -7957 -30 -7923
rect 4 -7957 106 -7923
rect 140 -7957 242 -7923
rect 276 -7957 389 -7923
rect -57 -7962 389 -7957
rect -57 -7963 16 -7962
rect 94 -7963 152 -7962
rect 227 -7963 389 -7962
rect 418 -7928 1122 -7910
rect 418 -7941 1076 -7928
rect 418 -7961 982 -7941
rect -57 -8019 12 -7963
rect 418 -7995 434 -7961
rect 468 -7993 982 -7961
rect 1034 -7962 1076 -7941
rect 1110 -7962 1122 -7928
rect 1034 -7993 1122 -7962
rect 468 -7995 1122 -7993
rect 418 -8001 1122 -7995
rect -862 -8028 13 -8019
rect 418 -8021 1076 -8001
rect 418 -8025 485 -8021
rect -862 -8062 -848 -8028
rect -814 -8062 -769 -8028
rect -735 -8062 13 -8028
rect -862 -8068 13 -8062
rect 1064 -8035 1076 -8021
rect 1110 -8035 1122 -8001
rect 1153 -7917 2449 -7900
rect 1153 -7922 2369 -7917
rect 1153 -7956 1171 -7922
rect 1205 -7956 1263 -7922
rect 1297 -7951 2369 -7922
rect 2403 -7951 2449 -7917
rect 1297 -7956 2449 -7951
rect 1153 -7962 2449 -7956
rect 2994 -7918 6963 -7898
rect 2994 -7952 3015 -7918
rect 3049 -7952 6876 -7918
rect 6910 -7952 6963 -7918
rect 1153 -8022 1310 -7962
rect 2994 -7969 6963 -7952
rect 7509 -7918 8255 -7897
rect 7509 -7952 7522 -7918
rect 7556 -7919 8255 -7918
rect 7556 -7952 8164 -7919
rect 7509 -7953 8164 -7952
rect 8198 -7953 8255 -7919
rect 7509 -7971 8255 -7953
rect 8799 -7917 9545 -7899
rect 8799 -7951 8811 -7917
rect 8845 -7951 9453 -7917
rect 9487 -7951 9545 -7917
rect 8799 -7970 9545 -7951
rect 10086 -7912 11058 -7894
rect 10086 -7916 11063 -7912
rect 10086 -7950 10099 -7916
rect 10133 -7917 11063 -7916
rect 10133 -7950 10741 -7917
rect 10086 -7951 10741 -7950
rect 10775 -7951 10832 -7917
rect 10866 -7918 11063 -7917
rect 10866 -7951 10925 -7918
rect 10086 -7952 10925 -7951
rect 10959 -7952 11017 -7918
rect 11051 -7952 11063 -7918
rect 11110 -7927 11120 -7875
rect 11172 -7927 11182 -7875
rect 11233 -7915 11418 -7828
rect 10086 -7958 11063 -7952
rect 11233 -7949 11250 -7915
rect 11284 -7949 11344 -7915
rect 11378 -7949 11418 -7915
rect 11233 -7957 11418 -7949
rect 10086 -7964 11058 -7958
rect 1064 -8090 1122 -8035
rect 1070 -8094 1116 -8090
rect -3193 -8155 16946 -8124
rect -3193 -8189 -2968 -8155
rect -2934 -8189 -2876 -8155
rect -2842 -8189 -2784 -8155
rect -2750 -8189 -2692 -8155
rect -2658 -8189 -2600 -8155
rect -2566 -8189 -2508 -8155
rect -2474 -8189 -2416 -8155
rect -2382 -8189 -2324 -8155
rect -2290 -8189 -2232 -8155
rect -2198 -8189 -2140 -8155
rect -2106 -8189 -2048 -8155
rect -2014 -8189 -1956 -8155
rect -1922 -8189 -1864 -8155
rect -1830 -8189 -1772 -8155
rect -1738 -8189 -1680 -8155
rect -1646 -8189 -1588 -8155
rect -1554 -8189 -1496 -8155
rect -1462 -8189 -1404 -8155
rect -1370 -8189 -1312 -8155
rect -1278 -8189 -1220 -8155
rect -1186 -8189 -1128 -8155
rect -1094 -8189 -1036 -8155
rect -1002 -8189 -944 -8155
rect -910 -8189 -852 -8155
rect -818 -8189 -760 -8155
rect -726 -8189 -668 -8155
rect -634 -8189 -576 -8155
rect -542 -8189 -484 -8155
rect -450 -8189 -392 -8155
rect -358 -8189 -300 -8155
rect -266 -8189 -208 -8155
rect -174 -8189 -116 -8155
rect -82 -8189 -24 -8155
rect 10 -8189 68 -8155
rect 102 -8189 160 -8155
rect 194 -8189 252 -8155
rect 286 -8189 344 -8155
rect 378 -8189 436 -8155
rect 470 -8189 528 -8155
rect 562 -8189 620 -8155
rect 654 -8189 712 -8155
rect 746 -8189 804 -8155
rect 838 -8189 896 -8155
rect 930 -8189 988 -8155
rect 1022 -8189 1080 -8155
rect 1114 -8189 1172 -8155
rect 1206 -8189 1264 -8155
rect 1298 -8189 1356 -8155
rect 1390 -8189 1448 -8155
rect 1482 -8189 1540 -8155
rect 1574 -8189 1632 -8155
rect 1666 -8189 1724 -8155
rect 1758 -8189 1816 -8155
rect 1850 -8189 1908 -8155
rect 1942 -8189 2000 -8155
rect 2034 -8189 2092 -8155
rect 2126 -8189 2184 -8155
rect 2218 -8189 2276 -8155
rect 2310 -8189 2368 -8155
rect 2402 -8189 2460 -8155
rect 2494 -8189 2552 -8155
rect 2586 -8189 2644 -8155
rect 2678 -8189 2736 -8155
rect 2770 -8189 2828 -8155
rect 2862 -8189 2920 -8155
rect 2954 -8189 3012 -8155
rect 3046 -8189 3104 -8155
rect 3138 -8189 3196 -8155
rect 3230 -8189 3288 -8155
rect 3322 -8189 3380 -8155
rect 3414 -8189 3472 -8155
rect 3506 -8189 3564 -8155
rect 3598 -8189 3656 -8155
rect 3690 -8189 3748 -8155
rect 3782 -8189 3840 -8155
rect 3874 -8189 3932 -8155
rect 3966 -8189 4024 -8155
rect 4058 -8189 4116 -8155
rect 4150 -8189 4208 -8155
rect 4242 -8189 4300 -8155
rect 4334 -8189 4392 -8155
rect 4426 -8189 4484 -8155
rect 4518 -8189 4576 -8155
rect 4610 -8189 4668 -8155
rect 4702 -8189 4760 -8155
rect 4794 -8189 4852 -8155
rect 4886 -8189 4944 -8155
rect 4978 -8189 5036 -8155
rect 5070 -8189 5128 -8155
rect 5162 -8189 5220 -8155
rect 5254 -8189 5312 -8155
rect 5346 -8189 5404 -8155
rect 5438 -8189 5496 -8155
rect 5530 -8189 5588 -8155
rect 5622 -8189 5680 -8155
rect 5714 -8189 5772 -8155
rect 5806 -8189 5864 -8155
rect 5898 -8189 5956 -8155
rect 5990 -8189 6048 -8155
rect 6082 -8189 6140 -8155
rect 6174 -8189 6232 -8155
rect 6266 -8189 6324 -8155
rect 6358 -8189 6416 -8155
rect 6450 -8189 6508 -8155
rect 6542 -8189 6600 -8155
rect 6634 -8189 6692 -8155
rect 6726 -8189 6784 -8155
rect 6818 -8189 6876 -8155
rect 6910 -8189 6968 -8155
rect 7002 -8189 7060 -8155
rect 7094 -8189 7152 -8155
rect 7186 -8189 7244 -8155
rect 7278 -8189 7336 -8155
rect 7370 -8189 7428 -8155
rect 7462 -8189 7520 -8155
rect 7554 -8189 7612 -8155
rect 7646 -8189 7704 -8155
rect 7738 -8189 7796 -8155
rect 7830 -8189 7888 -8155
rect 7922 -8189 7980 -8155
rect 8014 -8189 8072 -8155
rect 8106 -8189 8164 -8155
rect 8198 -8189 8256 -8155
rect 8290 -8189 8348 -8155
rect 8382 -8189 8440 -8155
rect 8474 -8189 8532 -8155
rect 8566 -8189 8624 -8155
rect 8658 -8189 8716 -8155
rect 8750 -8189 8808 -8155
rect 8842 -8189 8900 -8155
rect 8934 -8189 8992 -8155
rect 9026 -8189 9084 -8155
rect 9118 -8189 9176 -8155
rect 9210 -8189 9268 -8155
rect 9302 -8189 9360 -8155
rect 9394 -8189 9452 -8155
rect 9486 -8189 9544 -8155
rect 9578 -8189 9636 -8155
rect 9670 -8189 9728 -8155
rect 9762 -8189 9820 -8155
rect 9854 -8189 9912 -8155
rect 9946 -8189 10004 -8155
rect 10038 -8189 10096 -8155
rect 10130 -8189 10188 -8155
rect 10222 -8189 10280 -8155
rect 10314 -8189 10372 -8155
rect 10406 -8189 10464 -8155
rect 10498 -8189 10556 -8155
rect 10590 -8189 10648 -8155
rect 10682 -8189 10740 -8155
rect 10774 -8189 10832 -8155
rect 10866 -8189 10924 -8155
rect 10958 -8189 11016 -8155
rect 11050 -8189 11108 -8155
rect 11142 -8189 11200 -8155
rect 11234 -8189 11292 -8155
rect 11326 -8189 11384 -8155
rect 11418 -8189 11476 -8155
rect 11510 -8189 11568 -8155
rect 11602 -8189 11660 -8155
rect 11694 -8189 11752 -8155
rect 11786 -8189 11844 -8155
rect 11878 -8189 11936 -8155
rect 11970 -8189 12028 -8155
rect 12062 -8189 12120 -8155
rect 12154 -8189 12212 -8155
rect 12246 -8189 12304 -8155
rect 12338 -8189 12396 -8155
rect 12430 -8189 12488 -8155
rect 12522 -8189 12580 -8155
rect 12614 -8189 12672 -8155
rect 12706 -8189 12764 -8155
rect 12798 -8189 12856 -8155
rect 12890 -8189 12948 -8155
rect 12982 -8189 13040 -8155
rect 13074 -8189 13132 -8155
rect 13166 -8189 13224 -8155
rect 13258 -8189 13316 -8155
rect 13350 -8189 13408 -8155
rect 13442 -8189 13500 -8155
rect 13534 -8189 13592 -8155
rect 13626 -8189 13684 -8155
rect 13718 -8189 13776 -8155
rect 13810 -8189 13868 -8155
rect 13902 -8189 13960 -8155
rect 13994 -8189 14052 -8155
rect 14086 -8189 14144 -8155
rect 14178 -8189 14236 -8155
rect 14270 -8189 14328 -8155
rect 14362 -8189 14420 -8155
rect 14454 -8189 14512 -8155
rect 14546 -8189 14604 -8155
rect 14638 -8189 14696 -8155
rect 14730 -8189 14788 -8155
rect 14822 -8189 14880 -8155
rect 14914 -8189 14972 -8155
rect 15006 -8189 15064 -8155
rect 15098 -8189 15156 -8155
rect 15190 -8189 15248 -8155
rect 15282 -8189 15340 -8155
rect 15374 -8189 15432 -8155
rect 15466 -8189 15524 -8155
rect 15558 -8189 15616 -8155
rect 15650 -8189 15708 -8155
rect 15742 -8189 15800 -8155
rect 15834 -8189 15892 -8155
rect 15926 -8189 15984 -8155
rect 16018 -8189 16076 -8155
rect 16110 -8189 16168 -8155
rect 16202 -8189 16260 -8155
rect 16294 -8189 16352 -8155
rect 16386 -8189 16444 -8155
rect 16478 -8189 16536 -8155
rect 16570 -8189 16628 -8155
rect 16662 -8189 16946 -8155
rect -3193 -8220 16946 -8189
rect 13669 -8297 13738 -8295
rect 966 -8349 982 -8297
rect 1034 -8298 13738 -8297
rect 1034 -8349 12753 -8298
rect 966 -8350 12753 -8349
rect 12805 -8350 13738 -8298
rect 966 -8352 13738 -8350
rect 13669 -8362 13738 -8352
rect 1040 -8386 1098 -8385
rect 3000 -8386 3058 -8385
rect 1040 -8391 3058 -8386
rect 413 -8470 423 -8418
rect 475 -8470 485 -8418
rect 1040 -8425 1052 -8391
rect 1086 -8425 3012 -8391
rect 3046 -8425 3058 -8391
rect 1040 -8430 3058 -8425
rect 1040 -8431 1098 -8430
rect 3000 -8431 3058 -8430
rect 3614 -8386 3672 -8385
rect 5574 -8386 5632 -8385
rect 3614 -8391 5632 -8386
rect 3614 -8425 3626 -8391
rect 3660 -8425 5586 -8391
rect 5620 -8425 5632 -8391
rect 3614 -8430 5632 -8425
rect 3614 -8431 3672 -8430
rect 5574 -8431 5632 -8430
rect 6188 -8386 6246 -8385
rect 8148 -8386 8206 -8385
rect 6188 -8391 8206 -8386
rect 6188 -8425 6200 -8391
rect 6234 -8425 8160 -8391
rect 8194 -8425 8206 -8391
rect 6188 -8430 8206 -8425
rect 6188 -8431 6246 -8430
rect 8148 -8431 8206 -8430
rect 8762 -8386 8820 -8385
rect 8762 -8387 10320 -8386
rect 8762 -8391 10783 -8387
rect 8762 -8425 8774 -8391
rect 8808 -8393 10783 -8391
rect 8808 -8425 10737 -8393
rect 8762 -8427 10737 -8425
rect 10771 -8427 10783 -8393
rect 8762 -8430 10783 -8427
rect 8762 -8431 8820 -8430
rect 10131 -8431 10783 -8430
rect 10725 -8433 10783 -8431
rect 11338 -8394 11430 -8387
rect 11338 -8428 11369 -8394
rect 11403 -8428 11430 -8394
rect 11338 -8444 11430 -8428
rect 13669 -8396 13685 -8362
rect 13719 -8396 13738 -8362
rect 13669 -8439 13738 -8396
rect 15236 -8344 15294 -8338
rect 15328 -8344 15386 -8339
rect 15236 -8378 15248 -8344
rect 15282 -8345 15394 -8344
rect 15282 -8378 15340 -8345
rect 15236 -8379 15340 -8378
rect 15374 -8379 15394 -8345
rect 15236 -8424 15394 -8379
rect 15962 -8424 15972 -8416
rect 15236 -8440 15972 -8424
rect 11338 -8499 12463 -8444
rect 11339 -8503 12463 -8499
rect 12522 -8503 12532 -8444
rect 15236 -8474 15248 -8440
rect 15282 -8474 15341 -8440
rect 15375 -8464 15972 -8440
rect 15375 -8474 15394 -8464
rect 15236 -8480 15294 -8474
rect 15329 -8480 15387 -8474
rect 15962 -8475 15972 -8464
rect 16031 -8424 16041 -8416
rect 16031 -8464 16946 -8424
rect 16031 -8475 16041 -8464
rect -3193 -8699 16946 -8668
rect -3193 -8733 -2968 -8699
rect -2934 -8733 -2876 -8699
rect -2842 -8733 -2784 -8699
rect -2750 -8733 -2692 -8699
rect -2658 -8733 -2600 -8699
rect -2566 -8733 -2508 -8699
rect -2474 -8733 -2416 -8699
rect -2382 -8733 -2324 -8699
rect -2290 -8733 -2232 -8699
rect -2198 -8733 -2140 -8699
rect -2106 -8733 -2048 -8699
rect -2014 -8733 -1956 -8699
rect -1922 -8733 -1864 -8699
rect -1830 -8733 -1772 -8699
rect -1738 -8733 -1680 -8699
rect -1646 -8733 -1588 -8699
rect -1554 -8733 -1496 -8699
rect -1462 -8733 -1404 -8699
rect -1370 -8733 -1312 -8699
rect -1278 -8733 -1220 -8699
rect -1186 -8733 -1128 -8699
rect -1094 -8733 -1036 -8699
rect -1002 -8733 -944 -8699
rect -910 -8733 -852 -8699
rect -818 -8733 -760 -8699
rect -726 -8733 -668 -8699
rect -634 -8733 -576 -8699
rect -542 -8733 -484 -8699
rect -450 -8733 -392 -8699
rect -358 -8733 -300 -8699
rect -266 -8733 -208 -8699
rect -174 -8733 -116 -8699
rect -82 -8733 -24 -8699
rect 10 -8733 68 -8699
rect 102 -8733 160 -8699
rect 194 -8733 252 -8699
rect 286 -8733 344 -8699
rect 378 -8733 436 -8699
rect 470 -8733 528 -8699
rect 562 -8733 620 -8699
rect 654 -8733 712 -8699
rect 746 -8733 804 -8699
rect 838 -8733 896 -8699
rect 930 -8733 988 -8699
rect 1022 -8733 1080 -8699
rect 1114 -8733 1172 -8699
rect 1206 -8733 1264 -8699
rect 1298 -8733 1356 -8699
rect 1390 -8733 1448 -8699
rect 1482 -8733 1540 -8699
rect 1574 -8733 1632 -8699
rect 1666 -8733 1724 -8699
rect 1758 -8733 1816 -8699
rect 1850 -8733 1908 -8699
rect 1942 -8733 2000 -8699
rect 2034 -8733 2092 -8699
rect 2126 -8733 2184 -8699
rect 2218 -8733 2276 -8699
rect 2310 -8733 2368 -8699
rect 2402 -8733 2460 -8699
rect 2494 -8733 2552 -8699
rect 2586 -8733 2644 -8699
rect 2678 -8733 2736 -8699
rect 2770 -8733 2828 -8699
rect 2862 -8733 2920 -8699
rect 2954 -8733 3012 -8699
rect 3046 -8733 3104 -8699
rect 3138 -8733 3196 -8699
rect 3230 -8733 3288 -8699
rect 3322 -8733 3380 -8699
rect 3414 -8733 3472 -8699
rect 3506 -8733 3564 -8699
rect 3598 -8733 3656 -8699
rect 3690 -8733 3748 -8699
rect 3782 -8733 3840 -8699
rect 3874 -8733 3932 -8699
rect 3966 -8733 4024 -8699
rect 4058 -8733 4116 -8699
rect 4150 -8733 4208 -8699
rect 4242 -8733 4300 -8699
rect 4334 -8733 4392 -8699
rect 4426 -8733 4484 -8699
rect 4518 -8733 4576 -8699
rect 4610 -8733 4668 -8699
rect 4702 -8733 4760 -8699
rect 4794 -8733 4852 -8699
rect 4886 -8733 4944 -8699
rect 4978 -8733 5036 -8699
rect 5070 -8733 5128 -8699
rect 5162 -8733 5220 -8699
rect 5254 -8733 5312 -8699
rect 5346 -8733 5404 -8699
rect 5438 -8733 5496 -8699
rect 5530 -8733 5588 -8699
rect 5622 -8733 5680 -8699
rect 5714 -8733 5772 -8699
rect 5806 -8733 5864 -8699
rect 5898 -8733 5956 -8699
rect 5990 -8733 6048 -8699
rect 6082 -8733 6140 -8699
rect 6174 -8733 6232 -8699
rect 6266 -8733 6324 -8699
rect 6358 -8733 6416 -8699
rect 6450 -8733 6508 -8699
rect 6542 -8733 6600 -8699
rect 6634 -8733 6692 -8699
rect 6726 -8733 6784 -8699
rect 6818 -8733 6876 -8699
rect 6910 -8733 6968 -8699
rect 7002 -8733 7060 -8699
rect 7094 -8733 7152 -8699
rect 7186 -8733 7244 -8699
rect 7278 -8733 7336 -8699
rect 7370 -8733 7428 -8699
rect 7462 -8733 7520 -8699
rect 7554 -8733 7612 -8699
rect 7646 -8733 7704 -8699
rect 7738 -8733 7796 -8699
rect 7830 -8733 7888 -8699
rect 7922 -8733 7980 -8699
rect 8014 -8733 8072 -8699
rect 8106 -8733 8164 -8699
rect 8198 -8733 8256 -8699
rect 8290 -8733 8348 -8699
rect 8382 -8733 8440 -8699
rect 8474 -8733 8532 -8699
rect 8566 -8733 8624 -8699
rect 8658 -8733 8716 -8699
rect 8750 -8733 8808 -8699
rect 8842 -8733 8900 -8699
rect 8934 -8733 8992 -8699
rect 9026 -8733 9084 -8699
rect 9118 -8733 9176 -8699
rect 9210 -8733 9268 -8699
rect 9302 -8733 9360 -8699
rect 9394 -8733 9452 -8699
rect 9486 -8733 9544 -8699
rect 9578 -8733 9636 -8699
rect 9670 -8733 9728 -8699
rect 9762 -8733 9820 -8699
rect 9854 -8733 9912 -8699
rect 9946 -8733 10004 -8699
rect 10038 -8733 10096 -8699
rect 10130 -8733 10188 -8699
rect 10222 -8733 10280 -8699
rect 10314 -8733 10372 -8699
rect 10406 -8733 10464 -8699
rect 10498 -8733 10556 -8699
rect 10590 -8733 10648 -8699
rect 10682 -8733 10740 -8699
rect 10774 -8733 10832 -8699
rect 10866 -8733 10924 -8699
rect 10958 -8733 11016 -8699
rect 11050 -8733 11108 -8699
rect 11142 -8733 11200 -8699
rect 11234 -8733 11292 -8699
rect 11326 -8733 11384 -8699
rect 11418 -8733 11476 -8699
rect 11510 -8733 11568 -8699
rect 11602 -8733 11660 -8699
rect 11694 -8733 11752 -8699
rect 11786 -8733 11844 -8699
rect 11878 -8733 11936 -8699
rect 11970 -8733 12028 -8699
rect 12062 -8733 12120 -8699
rect 12154 -8733 12212 -8699
rect 12246 -8733 12304 -8699
rect 12338 -8733 12396 -8699
rect 12430 -8733 12488 -8699
rect 12522 -8733 12580 -8699
rect 12614 -8733 12672 -8699
rect 12706 -8733 12764 -8699
rect 12798 -8733 12856 -8699
rect 12890 -8733 12948 -8699
rect 12982 -8733 13040 -8699
rect 13074 -8733 13132 -8699
rect 13166 -8733 13224 -8699
rect 13258 -8733 13316 -8699
rect 13350 -8733 13408 -8699
rect 13442 -8733 13500 -8699
rect 13534 -8733 13592 -8699
rect 13626 -8733 13684 -8699
rect 13718 -8733 13776 -8699
rect 13810 -8733 13868 -8699
rect 13902 -8733 13960 -8699
rect 13994 -8733 14052 -8699
rect 14086 -8733 14144 -8699
rect 14178 -8733 14236 -8699
rect 14270 -8733 14328 -8699
rect 14362 -8733 14420 -8699
rect 14454 -8733 14512 -8699
rect 14546 -8733 14604 -8699
rect 14638 -8733 14696 -8699
rect 14730 -8733 14788 -8699
rect 14822 -8733 14880 -8699
rect 14914 -8733 14972 -8699
rect 15006 -8733 15064 -8699
rect 15098 -8733 15156 -8699
rect 15190 -8733 15248 -8699
rect 15282 -8733 15340 -8699
rect 15374 -8733 15432 -8699
rect 15466 -8733 15524 -8699
rect 15558 -8733 15616 -8699
rect 15650 -8733 15708 -8699
rect 15742 -8733 15800 -8699
rect 15834 -8733 15892 -8699
rect 15926 -8733 15984 -8699
rect 16018 -8733 16076 -8699
rect 16110 -8733 16168 -8699
rect 16202 -8733 16260 -8699
rect 16294 -8733 16352 -8699
rect 16386 -8733 16444 -8699
rect 16478 -8733 16536 -8699
rect 16570 -8733 16628 -8699
rect 16662 -8733 16946 -8699
rect -3193 -8764 16946 -8733
rect 7161 -8848 11181 -8847
rect 7161 -8851 11118 -8848
rect 7155 -8903 7165 -8851
rect 7217 -8900 11118 -8851
rect 11170 -8900 11181 -8848
rect 7217 -8903 11181 -8900
rect 7161 -8909 11181 -8903
rect 15236 -8954 15294 -8948
rect 15328 -8954 15386 -8949
rect 413 -9051 423 -8999
rect 475 -9051 485 -8999
rect 1070 -9000 1128 -8999
rect 3030 -9000 3088 -8999
rect 1070 -9005 3088 -9000
rect 1070 -9039 1082 -9005
rect 1116 -9039 3042 -9005
rect 3076 -9039 3088 -9005
rect 1070 -9044 3088 -9039
rect 1070 -9045 1128 -9044
rect 3030 -9045 3088 -9044
rect 3644 -9000 3702 -8999
rect 5604 -9000 5662 -8999
rect 3644 -9005 5662 -9000
rect 3644 -9039 3656 -9005
rect 3690 -9039 5616 -9005
rect 5650 -9039 5662 -9005
rect 3644 -9044 5662 -9039
rect 3644 -9045 3702 -9044
rect 5604 -9045 5662 -9044
rect 6218 -9000 6276 -8999
rect 8178 -9000 8236 -8999
rect 6218 -9005 8236 -9000
rect 6218 -9039 6230 -9005
rect 6264 -9039 8190 -9005
rect 8224 -9039 8236 -9005
rect 6218 -9044 8236 -9039
rect 6218 -9045 6276 -9044
rect 8178 -9045 8236 -9044
rect 8792 -9000 8850 -8999
rect 10752 -9000 10810 -8999
rect 8792 -9005 10810 -9000
rect 8792 -9039 8804 -9005
rect 8838 -9039 10764 -9005
rect 10798 -9039 10810 -9005
rect 11368 -9013 11378 -8961
rect 11430 -9013 11440 -8961
rect 15236 -8988 15248 -8954
rect 15282 -8955 15394 -8954
rect 15282 -8988 15340 -8955
rect 15236 -8989 15340 -8988
rect 15374 -8968 15394 -8955
rect 15374 -8989 16946 -8968
rect 13026 -8996 13084 -8995
rect 12548 -9002 12752 -8998
rect 12546 -9008 12752 -9002
rect 12804 -9008 12992 -8998
rect 8792 -9044 10810 -9039
rect 8792 -9045 8850 -9044
rect 10752 -9045 10810 -9044
rect 12546 -9042 12558 -9008
rect 12592 -9042 12642 -9008
rect 12676 -9042 12739 -9008
rect 12804 -9042 12836 -9008
rect 12870 -9042 12942 -9008
rect 12976 -9042 12992 -9008
rect 12546 -9048 12752 -9042
rect 12548 -9050 12752 -9048
rect 12804 -9050 12992 -9042
rect 12548 -9051 12992 -9050
rect 13026 -9001 13737 -8996
rect 13026 -9035 13038 -9001
rect 13072 -9035 13737 -9001
rect 13026 -9038 13737 -9035
rect 13026 -9072 13684 -9038
rect 13718 -9072 13737 -9038
rect 13026 -9073 13737 -9072
rect 13026 -9107 13038 -9073
rect 13072 -9106 13737 -9073
rect 15236 -9008 16946 -8989
rect 15236 -9050 15394 -9008
rect 15236 -9084 15248 -9050
rect 15282 -9084 15341 -9050
rect 15375 -9084 15394 -9050
rect 15236 -9090 15294 -9084
rect 15329 -9090 15387 -9084
rect 13072 -9107 13084 -9106
rect 13026 -9114 13084 -9107
rect -3193 -9243 16946 -9212
rect -3193 -9277 -2968 -9243
rect -2934 -9277 -2876 -9243
rect -2842 -9277 -2784 -9243
rect -2750 -9277 -2692 -9243
rect -2658 -9277 -2600 -9243
rect -2566 -9277 -2508 -9243
rect -2474 -9277 -2416 -9243
rect -2382 -9277 -2324 -9243
rect -2290 -9277 -2232 -9243
rect -2198 -9277 -2140 -9243
rect -2106 -9277 -2048 -9243
rect -2014 -9277 -1956 -9243
rect -1922 -9277 -1864 -9243
rect -1830 -9277 -1772 -9243
rect -1738 -9277 -1680 -9243
rect -1646 -9277 -1588 -9243
rect -1554 -9277 -1496 -9243
rect -1462 -9277 -1404 -9243
rect -1370 -9277 -1312 -9243
rect -1278 -9277 -1220 -9243
rect -1186 -9277 -1128 -9243
rect -1094 -9277 -1036 -9243
rect -1002 -9277 -944 -9243
rect -910 -9277 -852 -9243
rect -818 -9277 -760 -9243
rect -726 -9277 -668 -9243
rect -634 -9277 -576 -9243
rect -542 -9277 -484 -9243
rect -450 -9277 -392 -9243
rect -358 -9277 -300 -9243
rect -266 -9277 -208 -9243
rect -174 -9277 -116 -9243
rect -82 -9277 -24 -9243
rect 10 -9277 68 -9243
rect 102 -9277 160 -9243
rect 194 -9277 252 -9243
rect 286 -9277 344 -9243
rect 378 -9277 436 -9243
rect 470 -9277 528 -9243
rect 562 -9277 620 -9243
rect 654 -9277 712 -9243
rect 746 -9277 804 -9243
rect 838 -9277 896 -9243
rect 930 -9277 988 -9243
rect 1022 -9277 1080 -9243
rect 1114 -9277 1172 -9243
rect 1206 -9277 1264 -9243
rect 1298 -9277 1356 -9243
rect 1390 -9277 1448 -9243
rect 1482 -9277 1540 -9243
rect 1574 -9277 1632 -9243
rect 1666 -9277 1724 -9243
rect 1758 -9277 1816 -9243
rect 1850 -9277 1908 -9243
rect 1942 -9277 2000 -9243
rect 2034 -9277 2092 -9243
rect 2126 -9277 2184 -9243
rect 2218 -9277 2276 -9243
rect 2310 -9277 2368 -9243
rect 2402 -9277 2460 -9243
rect 2494 -9277 2552 -9243
rect 2586 -9277 2644 -9243
rect 2678 -9277 2736 -9243
rect 2770 -9277 2828 -9243
rect 2862 -9277 2920 -9243
rect 2954 -9277 3012 -9243
rect 3046 -9277 3104 -9243
rect 3138 -9277 3196 -9243
rect 3230 -9277 3288 -9243
rect 3322 -9277 3380 -9243
rect 3414 -9277 3472 -9243
rect 3506 -9277 3564 -9243
rect 3598 -9277 3656 -9243
rect 3690 -9277 3748 -9243
rect 3782 -9277 3840 -9243
rect 3874 -9277 3932 -9243
rect 3966 -9277 4024 -9243
rect 4058 -9277 4116 -9243
rect 4150 -9277 4208 -9243
rect 4242 -9277 4300 -9243
rect 4334 -9277 4392 -9243
rect 4426 -9277 4484 -9243
rect 4518 -9277 4576 -9243
rect 4610 -9277 4668 -9243
rect 4702 -9277 4760 -9243
rect 4794 -9277 4852 -9243
rect 4886 -9277 4944 -9243
rect 4978 -9277 5036 -9243
rect 5070 -9277 5128 -9243
rect 5162 -9277 5220 -9243
rect 5254 -9277 5312 -9243
rect 5346 -9277 5404 -9243
rect 5438 -9277 5496 -9243
rect 5530 -9277 5588 -9243
rect 5622 -9277 5680 -9243
rect 5714 -9277 5772 -9243
rect 5806 -9277 5864 -9243
rect 5898 -9277 5956 -9243
rect 5990 -9277 6048 -9243
rect 6082 -9277 6140 -9243
rect 6174 -9277 6232 -9243
rect 6266 -9277 6324 -9243
rect 6358 -9277 6416 -9243
rect 6450 -9277 6508 -9243
rect 6542 -9277 6600 -9243
rect 6634 -9277 6692 -9243
rect 6726 -9277 6784 -9243
rect 6818 -9277 6876 -9243
rect 6910 -9277 6968 -9243
rect 7002 -9277 7060 -9243
rect 7094 -9277 7152 -9243
rect 7186 -9277 7244 -9243
rect 7278 -9277 7336 -9243
rect 7370 -9277 7428 -9243
rect 7462 -9277 7520 -9243
rect 7554 -9277 7612 -9243
rect 7646 -9277 7704 -9243
rect 7738 -9277 7796 -9243
rect 7830 -9277 7888 -9243
rect 7922 -9277 7980 -9243
rect 8014 -9277 8072 -9243
rect 8106 -9277 8164 -9243
rect 8198 -9277 8256 -9243
rect 8290 -9277 8348 -9243
rect 8382 -9277 8440 -9243
rect 8474 -9277 8532 -9243
rect 8566 -9277 8624 -9243
rect 8658 -9277 8716 -9243
rect 8750 -9277 8808 -9243
rect 8842 -9277 8900 -9243
rect 8934 -9277 8992 -9243
rect 9026 -9277 9084 -9243
rect 9118 -9277 9176 -9243
rect 9210 -9277 9268 -9243
rect 9302 -9277 9360 -9243
rect 9394 -9277 9452 -9243
rect 9486 -9277 9544 -9243
rect 9578 -9277 9636 -9243
rect 9670 -9277 9728 -9243
rect 9762 -9277 9820 -9243
rect 9854 -9277 9912 -9243
rect 9946 -9277 10004 -9243
rect 10038 -9277 10096 -9243
rect 10130 -9277 10188 -9243
rect 10222 -9277 10280 -9243
rect 10314 -9277 10372 -9243
rect 10406 -9277 10464 -9243
rect 10498 -9277 10556 -9243
rect 10590 -9277 10648 -9243
rect 10682 -9277 10740 -9243
rect 10774 -9277 10832 -9243
rect 10866 -9277 10924 -9243
rect 10958 -9277 11016 -9243
rect 11050 -9277 11108 -9243
rect 11142 -9277 11200 -9243
rect 11234 -9277 11292 -9243
rect 11326 -9277 11384 -9243
rect 11418 -9277 11476 -9243
rect 11510 -9277 11568 -9243
rect 11602 -9277 11660 -9243
rect 11694 -9277 11752 -9243
rect 11786 -9277 11844 -9243
rect 11878 -9277 11936 -9243
rect 11970 -9277 12028 -9243
rect 12062 -9277 12120 -9243
rect 12154 -9277 12212 -9243
rect 12246 -9277 12304 -9243
rect 12338 -9277 12396 -9243
rect 12430 -9277 12488 -9243
rect 12522 -9277 12580 -9243
rect 12614 -9277 12672 -9243
rect 12706 -9277 12764 -9243
rect 12798 -9277 12856 -9243
rect 12890 -9277 12948 -9243
rect 12982 -9277 13040 -9243
rect 13074 -9277 13132 -9243
rect 13166 -9277 13224 -9243
rect 13258 -9277 13316 -9243
rect 13350 -9277 13408 -9243
rect 13442 -9277 13500 -9243
rect 13534 -9277 13592 -9243
rect 13626 -9277 13684 -9243
rect 13718 -9277 13776 -9243
rect 13810 -9277 13868 -9243
rect 13902 -9277 13960 -9243
rect 13994 -9277 14052 -9243
rect 14086 -9277 14144 -9243
rect 14178 -9277 14236 -9243
rect 14270 -9277 14328 -9243
rect 14362 -9277 14420 -9243
rect 14454 -9277 14512 -9243
rect 14546 -9277 14604 -9243
rect 14638 -9277 14696 -9243
rect 14730 -9277 14788 -9243
rect 14822 -9277 14880 -9243
rect 14914 -9277 14972 -9243
rect 15006 -9277 15064 -9243
rect 15098 -9277 15156 -9243
rect 15190 -9277 15248 -9243
rect 15282 -9277 15340 -9243
rect 15374 -9277 15432 -9243
rect 15466 -9277 15524 -9243
rect 15558 -9277 15616 -9243
rect 15650 -9277 15708 -9243
rect 15742 -9277 15800 -9243
rect 15834 -9277 15892 -9243
rect 15926 -9277 15984 -9243
rect 16018 -9277 16076 -9243
rect 16110 -9277 16168 -9243
rect 16202 -9277 16260 -9243
rect 16294 -9277 16352 -9243
rect 16386 -9277 16444 -9243
rect 16478 -9277 16536 -9243
rect 16570 -9277 16628 -9243
rect 16662 -9277 16946 -9243
rect -3193 -9308 16946 -9277
rect 13671 -9378 13735 -9377
rect 7153 -9379 13735 -9378
rect 7153 -9431 7163 -9379
rect 7215 -9382 13735 -9379
rect 7215 -9431 12756 -9382
rect 7153 -9432 12756 -9431
rect 12746 -9434 12756 -9432
rect 12808 -9432 13735 -9382
rect 12808 -9434 12818 -9432
rect 13671 -9448 13735 -9432
rect -952 -9559 -942 -9507
rect -890 -9509 -880 -9507
rect -890 -9516 -809 -9509
rect -890 -9550 -856 -9516
rect -822 -9550 -809 -9516
rect -227 -9522 -217 -9470
rect -165 -9522 -155 -9470
rect 1042 -9477 1100 -9476
rect 3002 -9477 3060 -9476
rect 1042 -9482 3060 -9477
rect -890 -9557 -809 -9550
rect -890 -9559 -880 -9557
rect 413 -9558 423 -9506
rect 475 -9558 485 -9506
rect 1042 -9516 1054 -9482
rect 1088 -9516 3014 -9482
rect 3048 -9516 3060 -9482
rect 1042 -9521 3060 -9516
rect 1042 -9522 1100 -9521
rect 3002 -9522 3060 -9521
rect 3616 -9477 3674 -9476
rect 5576 -9477 5634 -9476
rect 3616 -9482 5634 -9477
rect 3616 -9516 3628 -9482
rect 3662 -9516 5588 -9482
rect 5622 -9516 5634 -9482
rect 3616 -9521 5634 -9516
rect 3616 -9522 3674 -9521
rect 5576 -9522 5634 -9521
rect 6190 -9477 6248 -9476
rect 8150 -9477 8208 -9476
rect 6190 -9482 8208 -9477
rect 6190 -9516 6202 -9482
rect 6236 -9516 8162 -9482
rect 8196 -9516 8208 -9482
rect 6190 -9521 8208 -9516
rect 6190 -9522 6248 -9521
rect 8150 -9522 8208 -9521
rect 8764 -9477 8822 -9476
rect 10724 -9477 10782 -9476
rect 8764 -9482 10782 -9477
rect 8764 -9516 8776 -9482
rect 8810 -9516 10736 -9482
rect 10770 -9516 10782 -9482
rect 8764 -9521 10782 -9516
rect 8764 -9522 8822 -9521
rect 10724 -9522 10782 -9521
rect 11365 -9524 11375 -9472
rect 11427 -9524 11437 -9472
rect 13671 -9482 13685 -9448
rect 13719 -9482 13735 -9448
rect 13671 -9526 13735 -9482
rect 15236 -9432 15294 -9426
rect 15328 -9432 15386 -9427
rect 15236 -9466 15248 -9432
rect 15282 -9433 15394 -9432
rect 15282 -9466 15340 -9433
rect 15236 -9467 15340 -9466
rect 15374 -9467 15394 -9433
rect 15236 -9512 15394 -9467
rect 15236 -9528 16946 -9512
rect 15236 -9562 15248 -9528
rect 15282 -9562 15341 -9528
rect 15375 -9552 16946 -9528
rect 15375 -9562 15394 -9552
rect 15236 -9568 15294 -9562
rect 15329 -9568 15387 -9562
rect -3193 -9787 16946 -9756
rect -3193 -9821 -2968 -9787
rect -2934 -9821 -2876 -9787
rect -2842 -9821 -2784 -9787
rect -2750 -9821 -2692 -9787
rect -2658 -9821 -2600 -9787
rect -2566 -9821 -2508 -9787
rect -2474 -9821 -2416 -9787
rect -2382 -9821 -2324 -9787
rect -2290 -9821 -2232 -9787
rect -2198 -9821 -2140 -9787
rect -2106 -9821 -2048 -9787
rect -2014 -9821 -1956 -9787
rect -1922 -9821 -1864 -9787
rect -1830 -9821 -1772 -9787
rect -1738 -9821 -1680 -9787
rect -1646 -9821 -1588 -9787
rect -1554 -9821 -1496 -9787
rect -1462 -9821 -1404 -9787
rect -1370 -9821 -1312 -9787
rect -1278 -9821 -1220 -9787
rect -1186 -9821 -1128 -9787
rect -1094 -9821 -1036 -9787
rect -1002 -9821 -944 -9787
rect -910 -9821 -852 -9787
rect -818 -9821 -760 -9787
rect -726 -9821 -668 -9787
rect -634 -9821 -576 -9787
rect -542 -9821 -484 -9787
rect -450 -9821 -392 -9787
rect -358 -9821 -300 -9787
rect -266 -9821 -208 -9787
rect -174 -9821 -116 -9787
rect -82 -9821 -24 -9787
rect 10 -9821 68 -9787
rect 102 -9821 160 -9787
rect 194 -9821 252 -9787
rect 286 -9821 344 -9787
rect 378 -9821 436 -9787
rect 470 -9821 528 -9787
rect 562 -9821 620 -9787
rect 654 -9821 712 -9787
rect 746 -9821 804 -9787
rect 838 -9821 896 -9787
rect 930 -9821 988 -9787
rect 1022 -9821 1080 -9787
rect 1114 -9821 1172 -9787
rect 1206 -9821 1264 -9787
rect 1298 -9821 1356 -9787
rect 1390 -9821 1448 -9787
rect 1482 -9821 1540 -9787
rect 1574 -9821 1632 -9787
rect 1666 -9821 1724 -9787
rect 1758 -9821 1816 -9787
rect 1850 -9821 1908 -9787
rect 1942 -9821 2000 -9787
rect 2034 -9821 2092 -9787
rect 2126 -9821 2184 -9787
rect 2218 -9821 2276 -9787
rect 2310 -9821 2368 -9787
rect 2402 -9821 2460 -9787
rect 2494 -9821 2552 -9787
rect 2586 -9821 2644 -9787
rect 2678 -9821 2736 -9787
rect 2770 -9821 2828 -9787
rect 2862 -9821 2920 -9787
rect 2954 -9821 3012 -9787
rect 3046 -9821 3104 -9787
rect 3138 -9821 3196 -9787
rect 3230 -9821 3288 -9787
rect 3322 -9821 3380 -9787
rect 3414 -9821 3472 -9787
rect 3506 -9821 3564 -9787
rect 3598 -9821 3656 -9787
rect 3690 -9821 3748 -9787
rect 3782 -9821 3840 -9787
rect 3874 -9821 3932 -9787
rect 3966 -9821 4024 -9787
rect 4058 -9821 4116 -9787
rect 4150 -9821 4208 -9787
rect 4242 -9821 4300 -9787
rect 4334 -9821 4392 -9787
rect 4426 -9821 4484 -9787
rect 4518 -9821 4576 -9787
rect 4610 -9821 4668 -9787
rect 4702 -9821 4760 -9787
rect 4794 -9821 4852 -9787
rect 4886 -9821 4944 -9787
rect 4978 -9821 5036 -9787
rect 5070 -9821 5128 -9787
rect 5162 -9821 5220 -9787
rect 5254 -9821 5312 -9787
rect 5346 -9821 5404 -9787
rect 5438 -9821 5496 -9787
rect 5530 -9821 5588 -9787
rect 5622 -9821 5680 -9787
rect 5714 -9821 5772 -9787
rect 5806 -9821 5864 -9787
rect 5898 -9821 5956 -9787
rect 5990 -9821 6048 -9787
rect 6082 -9821 6140 -9787
rect 6174 -9821 6232 -9787
rect 6266 -9821 6324 -9787
rect 6358 -9821 6416 -9787
rect 6450 -9821 6508 -9787
rect 6542 -9821 6600 -9787
rect 6634 -9821 6692 -9787
rect 6726 -9821 6784 -9787
rect 6818 -9821 6876 -9787
rect 6910 -9821 6968 -9787
rect 7002 -9821 7060 -9787
rect 7094 -9821 7152 -9787
rect 7186 -9821 7244 -9787
rect 7278 -9821 7336 -9787
rect 7370 -9821 7428 -9787
rect 7462 -9821 7520 -9787
rect 7554 -9821 7612 -9787
rect 7646 -9821 7704 -9787
rect 7738 -9821 7796 -9787
rect 7830 -9821 7888 -9787
rect 7922 -9821 7980 -9787
rect 8014 -9821 8072 -9787
rect 8106 -9821 8164 -9787
rect 8198 -9821 8256 -9787
rect 8290 -9821 8348 -9787
rect 8382 -9821 8440 -9787
rect 8474 -9821 8532 -9787
rect 8566 -9821 8624 -9787
rect 8658 -9821 8716 -9787
rect 8750 -9821 8808 -9787
rect 8842 -9821 8900 -9787
rect 8934 -9821 8992 -9787
rect 9026 -9821 9084 -9787
rect 9118 -9821 9176 -9787
rect 9210 -9821 9268 -9787
rect 9302 -9821 9360 -9787
rect 9394 -9821 9452 -9787
rect 9486 -9821 9544 -9787
rect 9578 -9821 9636 -9787
rect 9670 -9821 9728 -9787
rect 9762 -9821 9820 -9787
rect 9854 -9821 9912 -9787
rect 9946 -9821 10004 -9787
rect 10038 -9821 10096 -9787
rect 10130 -9821 10188 -9787
rect 10222 -9821 10280 -9787
rect 10314 -9821 10372 -9787
rect 10406 -9821 10464 -9787
rect 10498 -9821 10556 -9787
rect 10590 -9821 10648 -9787
rect 10682 -9821 10740 -9787
rect 10774 -9821 10832 -9787
rect 10866 -9821 10924 -9787
rect 10958 -9821 11016 -9787
rect 11050 -9821 11108 -9787
rect 11142 -9821 11200 -9787
rect 11234 -9821 11292 -9787
rect 11326 -9821 11384 -9787
rect 11418 -9821 11476 -9787
rect 11510 -9821 11568 -9787
rect 11602 -9821 11660 -9787
rect 11694 -9821 11752 -9787
rect 11786 -9821 11844 -9787
rect 11878 -9821 11936 -9787
rect 11970 -9821 12028 -9787
rect 12062 -9821 12120 -9787
rect 12154 -9821 12212 -9787
rect 12246 -9821 12304 -9787
rect 12338 -9821 12396 -9787
rect 12430 -9821 12488 -9787
rect 12522 -9821 12580 -9787
rect 12614 -9821 12672 -9787
rect 12706 -9821 12764 -9787
rect 12798 -9821 12856 -9787
rect 12890 -9821 12948 -9787
rect 12982 -9821 13040 -9787
rect 13074 -9821 13132 -9787
rect 13166 -9821 13224 -9787
rect 13258 -9821 13316 -9787
rect 13350 -9821 13408 -9787
rect 13442 -9821 13500 -9787
rect 13534 -9821 13592 -9787
rect 13626 -9821 13684 -9787
rect 13718 -9821 13776 -9787
rect 13810 -9821 13868 -9787
rect 13902 -9821 13960 -9787
rect 13994 -9821 14052 -9787
rect 14086 -9821 14144 -9787
rect 14178 -9821 14236 -9787
rect 14270 -9821 14328 -9787
rect 14362 -9821 14420 -9787
rect 14454 -9821 14512 -9787
rect 14546 -9821 14604 -9787
rect 14638 -9821 14696 -9787
rect 14730 -9821 14788 -9787
rect 14822 -9821 14880 -9787
rect 14914 -9821 14972 -9787
rect 15006 -9821 15064 -9787
rect 15098 -9821 15156 -9787
rect 15190 -9821 15248 -9787
rect 15282 -9821 15340 -9787
rect 15374 -9821 15432 -9787
rect 15466 -9821 15524 -9787
rect 15558 -9821 15616 -9787
rect 15650 -9821 15708 -9787
rect 15742 -9821 15800 -9787
rect 15834 -9821 15892 -9787
rect 15926 -9821 15984 -9787
rect 16018 -9821 16076 -9787
rect 16110 -9821 16168 -9787
rect 16202 -9821 16260 -9787
rect 16294 -9821 16352 -9787
rect 16386 -9821 16444 -9787
rect 16478 -9821 16536 -9787
rect 16570 -9821 16628 -9787
rect 16662 -9821 16946 -9787
rect -3193 -9852 16946 -9821
rect 12467 -10023 12520 -9991
rect 12467 -10030 12480 -10023
rect 12514 -10030 12520 -10023
rect 418 -10137 428 -10085
rect 480 -10137 490 -10085
rect 1069 -10089 1127 -10088
rect 3029 -10089 3087 -10088
rect 1069 -10094 3087 -10089
rect 1069 -10128 1081 -10094
rect 1115 -10128 3041 -10094
rect 3075 -10128 3087 -10094
rect 1069 -10133 3087 -10128
rect 1069 -10134 1127 -10133
rect 3029 -10134 3087 -10133
rect 3643 -10089 3701 -10088
rect 5603 -10089 5661 -10088
rect 3643 -10094 5661 -10089
rect 3643 -10128 3655 -10094
rect 3689 -10128 5615 -10094
rect 5649 -10128 5661 -10094
rect 3643 -10133 5661 -10128
rect 3643 -10134 3701 -10133
rect 5603 -10134 5661 -10133
rect 6217 -10089 6275 -10088
rect 8177 -10089 8235 -10088
rect 6217 -10094 8235 -10089
rect 6217 -10128 6229 -10094
rect 6263 -10128 8189 -10094
rect 8223 -10128 8235 -10094
rect 6217 -10133 8235 -10128
rect 6217 -10134 6275 -10133
rect 8177 -10134 8235 -10133
rect 8791 -10089 8849 -10088
rect 10751 -10089 10809 -10088
rect 8791 -10094 10809 -10089
rect 8791 -10128 8806 -10094
rect 8840 -10128 10763 -10094
rect 10797 -10128 10809 -10094
rect 11368 -10104 11378 -10052
rect 11430 -10104 11440 -10052
rect 12456 -10082 12466 -10030
rect 12518 -10082 12520 -10030
rect 15236 -10042 15294 -10036
rect 15328 -10042 15386 -10036
rect 15236 -10076 15248 -10042
rect 15282 -10076 15340 -10042
rect 15374 -10056 15394 -10042
rect 15374 -10076 16946 -10056
rect 13027 -10077 13085 -10076
rect 12467 -10097 12520 -10082
rect 13023 -10082 13738 -10077
rect 12846 -10088 12991 -10087
rect 8791 -10133 10809 -10128
rect 8791 -10134 8849 -10133
rect 10751 -10134 10809 -10133
rect 12467 -10131 12480 -10097
rect 12514 -10131 12520 -10097
rect 12467 -10144 12520 -10131
rect 12548 -10095 12755 -10088
rect 12807 -10093 12993 -10088
rect 12548 -10129 12568 -10095
rect 12602 -10129 12659 -10095
rect 12693 -10129 12755 -10095
rect 12807 -10127 12858 -10093
rect 12892 -10127 12942 -10093
rect 12976 -10127 12993 -10093
rect 12548 -10137 12755 -10129
rect 12745 -10140 12755 -10137
rect 12807 -10137 12993 -10127
rect 13023 -10116 13039 -10082
rect 13073 -10116 13738 -10082
rect 13023 -10126 13738 -10116
rect 12807 -10140 12817 -10137
rect 12456 -10196 12466 -10144
rect 12518 -10196 12520 -10144
rect 12467 -10203 12480 -10196
rect 12514 -10203 12520 -10196
rect 13023 -10159 13685 -10126
rect 13023 -10193 13042 -10159
rect 13076 -10160 13685 -10159
rect 13719 -10160 13738 -10126
rect 13076 -10193 13738 -10160
rect 15236 -10096 16946 -10076
rect 15236 -10138 15394 -10096
rect 15236 -10172 15248 -10138
rect 15282 -10172 15341 -10138
rect 15375 -10172 15394 -10138
rect 15236 -10178 15294 -10172
rect 15329 -10178 15387 -10172
rect 13023 -10200 13738 -10193
rect 12467 -10228 12520 -10203
rect -3193 -10331 16946 -10300
rect -3193 -10365 -2968 -10331
rect -2934 -10365 -2876 -10331
rect -2842 -10365 -2784 -10331
rect -2750 -10365 -2692 -10331
rect -2658 -10365 -2600 -10331
rect -2566 -10365 -2508 -10331
rect -2474 -10365 -2416 -10331
rect -2382 -10365 -2324 -10331
rect -2290 -10365 -2232 -10331
rect -2198 -10365 -2140 -10331
rect -2106 -10365 -2048 -10331
rect -2014 -10365 -1956 -10331
rect -1922 -10365 -1864 -10331
rect -1830 -10365 -1772 -10331
rect -1738 -10365 -1680 -10331
rect -1646 -10365 -1588 -10331
rect -1554 -10365 -1496 -10331
rect -1462 -10365 -1404 -10331
rect -1370 -10365 -1312 -10331
rect -1278 -10365 -1220 -10331
rect -1186 -10365 -1128 -10331
rect -1094 -10365 -1036 -10331
rect -1002 -10365 -944 -10331
rect -910 -10365 -852 -10331
rect -818 -10365 -760 -10331
rect -726 -10365 -668 -10331
rect -634 -10365 -576 -10331
rect -542 -10365 -484 -10331
rect -450 -10365 -392 -10331
rect -358 -10365 -300 -10331
rect -266 -10365 -208 -10331
rect -174 -10365 -116 -10331
rect -82 -10365 -24 -10331
rect 10 -10365 68 -10331
rect 102 -10365 160 -10331
rect 194 -10365 252 -10331
rect 286 -10365 344 -10331
rect 378 -10365 436 -10331
rect 470 -10365 528 -10331
rect 562 -10365 620 -10331
rect 654 -10365 712 -10331
rect 746 -10365 804 -10331
rect 838 -10365 896 -10331
rect 930 -10365 988 -10331
rect 1022 -10365 1080 -10331
rect 1114 -10365 1172 -10331
rect 1206 -10365 1264 -10331
rect 1298 -10365 1356 -10331
rect 1390 -10365 1448 -10331
rect 1482 -10365 1540 -10331
rect 1574 -10365 1632 -10331
rect 1666 -10365 1724 -10331
rect 1758 -10365 1816 -10331
rect 1850 -10365 1908 -10331
rect 1942 -10365 2000 -10331
rect 2034 -10365 2092 -10331
rect 2126 -10365 2184 -10331
rect 2218 -10365 2276 -10331
rect 2310 -10365 2368 -10331
rect 2402 -10365 2460 -10331
rect 2494 -10365 2552 -10331
rect 2586 -10365 2644 -10331
rect 2678 -10365 2736 -10331
rect 2770 -10365 2828 -10331
rect 2862 -10365 2920 -10331
rect 2954 -10365 3012 -10331
rect 3046 -10365 3104 -10331
rect 3138 -10365 3196 -10331
rect 3230 -10365 3288 -10331
rect 3322 -10365 3380 -10331
rect 3414 -10365 3472 -10331
rect 3506 -10365 3564 -10331
rect 3598 -10365 3656 -10331
rect 3690 -10365 3748 -10331
rect 3782 -10365 3840 -10331
rect 3874 -10365 3932 -10331
rect 3966 -10365 4024 -10331
rect 4058 -10365 4116 -10331
rect 4150 -10365 4208 -10331
rect 4242 -10365 4300 -10331
rect 4334 -10365 4392 -10331
rect 4426 -10365 4484 -10331
rect 4518 -10365 4576 -10331
rect 4610 -10365 4668 -10331
rect 4702 -10365 4760 -10331
rect 4794 -10365 4852 -10331
rect 4886 -10365 4944 -10331
rect 4978 -10365 5036 -10331
rect 5070 -10365 5128 -10331
rect 5162 -10365 5220 -10331
rect 5254 -10365 5312 -10331
rect 5346 -10365 5404 -10331
rect 5438 -10365 5496 -10331
rect 5530 -10365 5588 -10331
rect 5622 -10365 5680 -10331
rect 5714 -10365 5772 -10331
rect 5806 -10365 5864 -10331
rect 5898 -10365 5956 -10331
rect 5990 -10365 6048 -10331
rect 6082 -10365 6140 -10331
rect 6174 -10365 6232 -10331
rect 6266 -10365 6324 -10331
rect 6358 -10365 6416 -10331
rect 6450 -10365 6508 -10331
rect 6542 -10365 6600 -10331
rect 6634 -10365 6692 -10331
rect 6726 -10365 6784 -10331
rect 6818 -10365 6876 -10331
rect 6910 -10365 6968 -10331
rect 7002 -10365 7060 -10331
rect 7094 -10365 7152 -10331
rect 7186 -10365 7244 -10331
rect 7278 -10365 7336 -10331
rect 7370 -10365 7428 -10331
rect 7462 -10365 7520 -10331
rect 7554 -10365 7612 -10331
rect 7646 -10365 7704 -10331
rect 7738 -10365 7796 -10331
rect 7830 -10365 7888 -10331
rect 7922 -10365 7980 -10331
rect 8014 -10365 8072 -10331
rect 8106 -10365 8164 -10331
rect 8198 -10365 8256 -10331
rect 8290 -10365 8348 -10331
rect 8382 -10365 8440 -10331
rect 8474 -10365 8532 -10331
rect 8566 -10365 8624 -10331
rect 8658 -10365 8716 -10331
rect 8750 -10365 8808 -10331
rect 8842 -10365 8900 -10331
rect 8934 -10365 8992 -10331
rect 9026 -10365 9084 -10331
rect 9118 -10365 9176 -10331
rect 9210 -10365 9268 -10331
rect 9302 -10365 9360 -10331
rect 9394 -10365 9452 -10331
rect 9486 -10365 9544 -10331
rect 9578 -10365 9636 -10331
rect 9670 -10365 9728 -10331
rect 9762 -10365 9820 -10331
rect 9854 -10365 9912 -10331
rect 9946 -10365 10004 -10331
rect 10038 -10365 10096 -10331
rect 10130 -10365 10188 -10331
rect 10222 -10365 10280 -10331
rect 10314 -10365 10372 -10331
rect 10406 -10365 10464 -10331
rect 10498 -10365 10556 -10331
rect 10590 -10365 10648 -10331
rect 10682 -10365 10740 -10331
rect 10774 -10365 10832 -10331
rect 10866 -10365 10924 -10331
rect 10958 -10365 11016 -10331
rect 11050 -10365 11108 -10331
rect 11142 -10365 11200 -10331
rect 11234 -10365 11292 -10331
rect 11326 -10365 11384 -10331
rect 11418 -10365 11476 -10331
rect 11510 -10365 11568 -10331
rect 11602 -10365 11660 -10331
rect 11694 -10365 11752 -10331
rect 11786 -10365 11844 -10331
rect 11878 -10365 11936 -10331
rect 11970 -10365 12028 -10331
rect 12062 -10365 12120 -10331
rect 12154 -10365 12212 -10331
rect 12246 -10365 12304 -10331
rect 12338 -10365 12396 -10331
rect 12430 -10365 12488 -10331
rect 12522 -10365 12580 -10331
rect 12614 -10365 12672 -10331
rect 12706 -10365 12764 -10331
rect 12798 -10365 12856 -10331
rect 12890 -10365 12948 -10331
rect 12982 -10365 13040 -10331
rect 13074 -10365 13132 -10331
rect 13166 -10365 13224 -10331
rect 13258 -10365 13316 -10331
rect 13350 -10365 13408 -10331
rect 13442 -10365 13500 -10331
rect 13534 -10365 13592 -10331
rect 13626 -10365 13684 -10331
rect 13718 -10365 13776 -10331
rect 13810 -10365 13868 -10331
rect 13902 -10365 13960 -10331
rect 13994 -10365 14052 -10331
rect 14086 -10365 14144 -10331
rect 14178 -10365 14236 -10331
rect 14270 -10365 14328 -10331
rect 14362 -10365 14420 -10331
rect 14454 -10365 14512 -10331
rect 14546 -10365 14604 -10331
rect 14638 -10365 14696 -10331
rect 14730 -10365 14788 -10331
rect 14822 -10365 14880 -10331
rect 14914 -10365 14972 -10331
rect 15006 -10365 15064 -10331
rect 15098 -10365 15156 -10331
rect 15190 -10365 15248 -10331
rect 15282 -10365 15340 -10331
rect 15374 -10365 15432 -10331
rect 15466 -10365 15524 -10331
rect 15558 -10365 15616 -10331
rect 15650 -10365 15708 -10331
rect 15742 -10365 15800 -10331
rect 15834 -10365 15892 -10331
rect 15926 -10365 15984 -10331
rect 16018 -10365 16076 -10331
rect 16110 -10365 16168 -10331
rect 16202 -10365 16260 -10331
rect 16294 -10365 16352 -10331
rect 16386 -10365 16444 -10331
rect 16478 -10365 16536 -10331
rect 16570 -10365 16628 -10331
rect 16662 -10365 16946 -10331
rect -3193 -10396 16946 -10365
rect -2617 -10490 -1969 -10489
rect -2617 -10543 -2607 -10490
rect -2554 -10543 -1969 -10490
rect -1915 -10543 -1905 -10489
rect -1833 -10579 -1823 -10525
rect -1769 -10579 -1759 -10525
rect 1035 -10568 1699 -10562
rect 3004 -10564 3062 -10563
rect -225 -10597 479 -10595
rect -231 -10649 -221 -10597
rect -169 -10603 479 -10597
rect -169 -10637 429 -10603
rect 463 -10637 479 -10603
rect 1035 -10602 1072 -10568
rect 1106 -10602 1699 -10568
rect 1035 -10609 1699 -10602
rect 2401 -10569 3062 -10564
rect 2401 -10603 3016 -10569
rect 3050 -10603 3062 -10569
rect 2401 -10608 3062 -10603
rect 3004 -10609 3062 -10608
rect 3618 -10564 3676 -10563
rect 5578 -10564 5636 -10563
rect 3618 -10569 5636 -10564
rect 3618 -10603 3630 -10569
rect 3664 -10603 5590 -10569
rect 5624 -10603 5636 -10569
rect 3618 -10608 5636 -10603
rect 3618 -10609 3676 -10608
rect 5578 -10609 5636 -10608
rect 6192 -10564 6250 -10563
rect 8152 -10564 8210 -10563
rect 6192 -10569 8210 -10564
rect 6192 -10603 6204 -10569
rect 6238 -10603 8164 -10569
rect 8198 -10603 8210 -10569
rect 6192 -10608 8210 -10603
rect 6192 -10609 6250 -10608
rect 8152 -10609 8210 -10608
rect 8766 -10564 8824 -10563
rect 10145 -10564 10783 -10562
rect 8766 -10569 10784 -10564
rect 8766 -10603 8778 -10569
rect 8812 -10570 10784 -10569
rect 8812 -10603 10738 -10570
rect 8766 -10604 10738 -10603
rect 10772 -10604 10784 -10570
rect 8766 -10608 10784 -10604
rect 8766 -10609 8824 -10608
rect 10145 -10610 10784 -10608
rect 10145 -10614 10783 -10610
rect 11366 -10611 11376 -10559
rect 11428 -10611 11438 -10559
rect -169 -10649 479 -10637
rect -3193 -10875 16946 -10844
rect -3193 -10909 -2968 -10875
rect -2934 -10909 -2876 -10875
rect -2842 -10909 -2784 -10875
rect -2750 -10909 -2692 -10875
rect -2658 -10909 -2600 -10875
rect -2566 -10909 -2508 -10875
rect -2474 -10909 -2416 -10875
rect -2382 -10909 -2324 -10875
rect -2290 -10909 -2232 -10875
rect -2198 -10909 -2140 -10875
rect -2106 -10909 -2048 -10875
rect -2014 -10909 -1956 -10875
rect -1922 -10909 -1864 -10875
rect -1830 -10909 -1772 -10875
rect -1738 -10909 -1680 -10875
rect -1646 -10909 -1588 -10875
rect -1554 -10909 -1496 -10875
rect -1462 -10909 -1404 -10875
rect -1370 -10909 -1312 -10875
rect -1278 -10909 -1220 -10875
rect -1186 -10909 -1128 -10875
rect -1094 -10909 -1036 -10875
rect -1002 -10909 -944 -10875
rect -910 -10909 -852 -10875
rect -818 -10909 -760 -10875
rect -726 -10909 -668 -10875
rect -634 -10909 -576 -10875
rect -542 -10909 -484 -10875
rect -450 -10909 -392 -10875
rect -358 -10909 -300 -10875
rect -266 -10909 -208 -10875
rect -174 -10909 -116 -10875
rect -82 -10909 -24 -10875
rect 10 -10909 68 -10875
rect 102 -10909 160 -10875
rect 194 -10909 252 -10875
rect 286 -10909 344 -10875
rect 378 -10909 436 -10875
rect 470 -10909 528 -10875
rect 562 -10909 620 -10875
rect 654 -10909 712 -10875
rect 746 -10909 804 -10875
rect 838 -10909 896 -10875
rect 930 -10909 988 -10875
rect 1022 -10909 1080 -10875
rect 1114 -10909 1172 -10875
rect 1206 -10909 1264 -10875
rect 1298 -10909 1356 -10875
rect 1390 -10909 1448 -10875
rect 1482 -10909 1540 -10875
rect 1574 -10909 1632 -10875
rect 1666 -10909 1724 -10875
rect 1758 -10909 1816 -10875
rect 1850 -10909 1908 -10875
rect 1942 -10909 2000 -10875
rect 2034 -10909 2092 -10875
rect 2126 -10909 2184 -10875
rect 2218 -10909 2276 -10875
rect 2310 -10909 2368 -10875
rect 2402 -10909 2460 -10875
rect 2494 -10909 2552 -10875
rect 2586 -10909 2644 -10875
rect 2678 -10909 2736 -10875
rect 2770 -10909 2828 -10875
rect 2862 -10909 2920 -10875
rect 2954 -10909 3012 -10875
rect 3046 -10909 3104 -10875
rect 3138 -10909 3196 -10875
rect 3230 -10909 3288 -10875
rect 3322 -10909 3380 -10875
rect 3414 -10909 3472 -10875
rect 3506 -10909 3564 -10875
rect 3598 -10909 3656 -10875
rect 3690 -10909 3748 -10875
rect 3782 -10909 3840 -10875
rect 3874 -10909 3932 -10875
rect 3966 -10909 4024 -10875
rect 4058 -10909 4116 -10875
rect 4150 -10909 4208 -10875
rect 4242 -10909 4300 -10875
rect 4334 -10909 4392 -10875
rect 4426 -10909 4484 -10875
rect 4518 -10909 4576 -10875
rect 4610 -10909 4668 -10875
rect 4702 -10909 4760 -10875
rect 4794 -10909 4852 -10875
rect 4886 -10909 4944 -10875
rect 4978 -10909 5036 -10875
rect 5070 -10909 5128 -10875
rect 5162 -10909 5220 -10875
rect 5254 -10909 5312 -10875
rect 5346 -10909 5404 -10875
rect 5438 -10909 5496 -10875
rect 5530 -10909 5588 -10875
rect 5622 -10909 5680 -10875
rect 5714 -10909 5772 -10875
rect 5806 -10909 5864 -10875
rect 5898 -10909 5956 -10875
rect 5990 -10909 6048 -10875
rect 6082 -10909 6140 -10875
rect 6174 -10909 6232 -10875
rect 6266 -10909 6324 -10875
rect 6358 -10909 6416 -10875
rect 6450 -10909 6508 -10875
rect 6542 -10909 6600 -10875
rect 6634 -10909 6692 -10875
rect 6726 -10909 6784 -10875
rect 6818 -10909 6876 -10875
rect 6910 -10909 6968 -10875
rect 7002 -10909 7060 -10875
rect 7094 -10909 7152 -10875
rect 7186 -10909 7244 -10875
rect 7278 -10909 7336 -10875
rect 7370 -10909 7428 -10875
rect 7462 -10909 7520 -10875
rect 7554 -10909 7612 -10875
rect 7646 -10909 7704 -10875
rect 7738 -10909 7796 -10875
rect 7830 -10909 7888 -10875
rect 7922 -10909 7980 -10875
rect 8014 -10909 8072 -10875
rect 8106 -10909 8164 -10875
rect 8198 -10909 8256 -10875
rect 8290 -10909 8348 -10875
rect 8382 -10909 8440 -10875
rect 8474 -10909 8532 -10875
rect 8566 -10909 8624 -10875
rect 8658 -10909 8716 -10875
rect 8750 -10909 8808 -10875
rect 8842 -10909 8900 -10875
rect 8934 -10909 8992 -10875
rect 9026 -10909 9084 -10875
rect 9118 -10909 9176 -10875
rect 9210 -10909 9268 -10875
rect 9302 -10909 9360 -10875
rect 9394 -10909 9452 -10875
rect 9486 -10909 9544 -10875
rect 9578 -10909 9636 -10875
rect 9670 -10909 9728 -10875
rect 9762 -10909 9820 -10875
rect 9854 -10909 9912 -10875
rect 9946 -10909 10004 -10875
rect 10038 -10909 10096 -10875
rect 10130 -10909 10188 -10875
rect 10222 -10909 10280 -10875
rect 10314 -10909 10372 -10875
rect 10406 -10909 10464 -10875
rect 10498 -10909 10556 -10875
rect 10590 -10909 10648 -10875
rect 10682 -10909 10740 -10875
rect 10774 -10909 10832 -10875
rect 10866 -10909 10924 -10875
rect 10958 -10909 11016 -10875
rect 11050 -10909 11108 -10875
rect 11142 -10909 11200 -10875
rect 11234 -10909 11292 -10875
rect 11326 -10909 11384 -10875
rect 11418 -10909 11476 -10875
rect 11510 -10909 11568 -10875
rect 11602 -10909 11660 -10875
rect 11694 -10909 11752 -10875
rect 11786 -10909 11844 -10875
rect 11878 -10909 11936 -10875
rect 11970 -10909 12028 -10875
rect 12062 -10909 12120 -10875
rect 12154 -10909 12212 -10875
rect 12246 -10909 12304 -10875
rect 12338 -10909 12396 -10875
rect 12430 -10909 12488 -10875
rect 12522 -10909 12580 -10875
rect 12614 -10909 12672 -10875
rect 12706 -10909 12764 -10875
rect 12798 -10909 12856 -10875
rect 12890 -10909 12948 -10875
rect 12982 -10909 13040 -10875
rect 13074 -10909 13132 -10875
rect 13166 -10909 13224 -10875
rect 13258 -10909 13316 -10875
rect 13350 -10909 13408 -10875
rect 13442 -10909 13500 -10875
rect 13534 -10909 13592 -10875
rect 13626 -10909 13684 -10875
rect 13718 -10909 13776 -10875
rect 13810 -10909 13868 -10875
rect 13902 -10909 13960 -10875
rect 13994 -10909 14052 -10875
rect 14086 -10909 14144 -10875
rect 14178 -10909 14236 -10875
rect 14270 -10909 14328 -10875
rect 14362 -10909 14420 -10875
rect 14454 -10909 14512 -10875
rect 14546 -10909 14604 -10875
rect 14638 -10909 14696 -10875
rect 14730 -10909 14788 -10875
rect 14822 -10909 14880 -10875
rect 14914 -10909 14972 -10875
rect 15006 -10909 15064 -10875
rect 15098 -10909 15156 -10875
rect 15190 -10909 15248 -10875
rect 15282 -10909 15340 -10875
rect 15374 -10909 15432 -10875
rect 15466 -10909 15524 -10875
rect 15558 -10909 15616 -10875
rect 15650 -10909 15708 -10875
rect 15742 -10909 15800 -10875
rect 15834 -10909 15892 -10875
rect 15926 -10909 15984 -10875
rect 16018 -10909 16076 -10875
rect 16110 -10909 16168 -10875
rect 16202 -10909 16260 -10875
rect 16294 -10909 16352 -10875
rect 16386 -10909 16444 -10875
rect 16478 -10909 16536 -10875
rect 16570 -10909 16628 -10875
rect 16662 -10909 16946 -10875
rect -3193 -10940 16946 -10909
rect 105 -11189 115 -11137
rect 167 -11139 177 -11137
rect 167 -11147 481 -11139
rect 167 -11181 432 -11147
rect 466 -11181 481 -11147
rect 3004 -11176 3062 -11175
rect 2409 -11177 3062 -11176
rect 167 -11188 481 -11181
rect 1033 -11181 3062 -11177
rect 1033 -11184 3016 -11181
rect 167 -11189 177 -11188
rect 1033 -11218 1070 -11184
rect 1104 -11215 3016 -11184
rect 3050 -11215 3062 -11181
rect 1104 -11218 3062 -11215
rect 1033 -11220 3062 -11218
rect 1033 -11226 2499 -11220
rect 3004 -11221 3062 -11220
rect 3618 -11176 3676 -11175
rect 5578 -11176 5636 -11175
rect 3618 -11181 5636 -11176
rect 3618 -11215 3630 -11181
rect 3664 -11215 5590 -11181
rect 5624 -11215 5636 -11181
rect 3618 -11220 5636 -11215
rect 3618 -11221 3676 -11220
rect 5578 -11221 5636 -11220
rect 6192 -11176 6250 -11175
rect 8152 -11176 8210 -11175
rect 6192 -11181 8210 -11176
rect 6192 -11215 6204 -11181
rect 6238 -11215 8164 -11181
rect 8198 -11215 8210 -11181
rect 6192 -11220 8210 -11215
rect 6192 -11221 6250 -11220
rect 8152 -11221 8210 -11220
rect 8766 -11176 8824 -11175
rect 10147 -11176 10783 -11173
rect 8766 -11181 10783 -11176
rect 8766 -11215 8778 -11181
rect 8812 -11184 10783 -11181
rect 8812 -11215 10735 -11184
rect 8766 -11218 10735 -11215
rect 10769 -11218 10783 -11184
rect 8766 -11220 10783 -11218
rect 8766 -11221 8824 -11220
rect 10147 -11223 10783 -11220
rect 10723 -11224 10781 -11223
rect 11363 -11225 11373 -11173
rect 11425 -11225 11435 -11173
rect -3193 -11419 16946 -11388
rect -3193 -11453 -2968 -11419
rect -2934 -11453 -2876 -11419
rect -2842 -11453 -2784 -11419
rect -2750 -11453 -2692 -11419
rect -2658 -11453 -2600 -11419
rect -2566 -11453 -2508 -11419
rect -2474 -11453 -2416 -11419
rect -2382 -11453 -2324 -11419
rect -2290 -11453 -2232 -11419
rect -2198 -11453 -2140 -11419
rect -2106 -11453 -2048 -11419
rect -2014 -11453 -1956 -11419
rect -1922 -11453 -1864 -11419
rect -1830 -11453 -1772 -11419
rect -1738 -11453 -1680 -11419
rect -1646 -11453 -1588 -11419
rect -1554 -11453 -1496 -11419
rect -1462 -11453 -1404 -11419
rect -1370 -11453 -1312 -11419
rect -1278 -11453 -1220 -11419
rect -1186 -11453 -1128 -11419
rect -1094 -11453 -1036 -11419
rect -1002 -11453 -944 -11419
rect -910 -11453 -852 -11419
rect -818 -11453 -760 -11419
rect -726 -11453 -668 -11419
rect -634 -11453 -576 -11419
rect -542 -11453 -484 -11419
rect -450 -11453 -392 -11419
rect -358 -11453 -300 -11419
rect -266 -11453 -208 -11419
rect -174 -11453 -116 -11419
rect -82 -11453 -24 -11419
rect 10 -11453 68 -11419
rect 102 -11453 160 -11419
rect 194 -11453 252 -11419
rect 286 -11453 344 -11419
rect 378 -11453 436 -11419
rect 470 -11453 528 -11419
rect 562 -11453 620 -11419
rect 654 -11453 712 -11419
rect 746 -11453 804 -11419
rect 838 -11453 896 -11419
rect 930 -11453 988 -11419
rect 1022 -11453 1080 -11419
rect 1114 -11453 1172 -11419
rect 1206 -11453 1264 -11419
rect 1298 -11453 1356 -11419
rect 1390 -11453 1448 -11419
rect 1482 -11453 1540 -11419
rect 1574 -11453 1632 -11419
rect 1666 -11453 1724 -11419
rect 1758 -11453 1816 -11419
rect 1850 -11453 1908 -11419
rect 1942 -11453 2000 -11419
rect 2034 -11453 2092 -11419
rect 2126 -11453 2184 -11419
rect 2218 -11453 2276 -11419
rect 2310 -11453 2368 -11419
rect 2402 -11453 2460 -11419
rect 2494 -11453 2552 -11419
rect 2586 -11453 2644 -11419
rect 2678 -11453 2736 -11419
rect 2770 -11453 2828 -11419
rect 2862 -11453 2920 -11419
rect 2954 -11453 3012 -11419
rect 3046 -11453 3104 -11419
rect 3138 -11453 3196 -11419
rect 3230 -11453 3288 -11419
rect 3322 -11453 3380 -11419
rect 3414 -11453 3472 -11419
rect 3506 -11453 3564 -11419
rect 3598 -11453 3656 -11419
rect 3690 -11453 3748 -11419
rect 3782 -11453 3840 -11419
rect 3874 -11453 3932 -11419
rect 3966 -11453 4024 -11419
rect 4058 -11453 4116 -11419
rect 4150 -11453 4208 -11419
rect 4242 -11453 4300 -11419
rect 4334 -11453 4392 -11419
rect 4426 -11453 4484 -11419
rect 4518 -11453 4576 -11419
rect 4610 -11453 4668 -11419
rect 4702 -11453 4760 -11419
rect 4794 -11453 4852 -11419
rect 4886 -11453 4944 -11419
rect 4978 -11453 5036 -11419
rect 5070 -11453 5128 -11419
rect 5162 -11453 5220 -11419
rect 5254 -11453 5312 -11419
rect 5346 -11453 5404 -11419
rect 5438 -11453 5496 -11419
rect 5530 -11453 5588 -11419
rect 5622 -11453 5680 -11419
rect 5714 -11453 5772 -11419
rect 5806 -11453 5864 -11419
rect 5898 -11453 5956 -11419
rect 5990 -11453 6048 -11419
rect 6082 -11453 6140 -11419
rect 6174 -11453 6232 -11419
rect 6266 -11453 6324 -11419
rect 6358 -11453 6416 -11419
rect 6450 -11453 6508 -11419
rect 6542 -11453 6600 -11419
rect 6634 -11453 6692 -11419
rect 6726 -11453 6784 -11419
rect 6818 -11453 6876 -11419
rect 6910 -11453 6968 -11419
rect 7002 -11453 7060 -11419
rect 7094 -11453 7152 -11419
rect 7186 -11453 7244 -11419
rect 7278 -11453 7336 -11419
rect 7370 -11453 7428 -11419
rect 7462 -11453 7520 -11419
rect 7554 -11453 7612 -11419
rect 7646 -11453 7704 -11419
rect 7738 -11453 7796 -11419
rect 7830 -11453 7888 -11419
rect 7922 -11453 7980 -11419
rect 8014 -11453 8072 -11419
rect 8106 -11453 8164 -11419
rect 8198 -11453 8256 -11419
rect 8290 -11453 8348 -11419
rect 8382 -11453 8440 -11419
rect 8474 -11453 8532 -11419
rect 8566 -11453 8624 -11419
rect 8658 -11453 8716 -11419
rect 8750 -11453 8808 -11419
rect 8842 -11453 8900 -11419
rect 8934 -11453 8992 -11419
rect 9026 -11453 9084 -11419
rect 9118 -11453 9176 -11419
rect 9210 -11453 9268 -11419
rect 9302 -11453 9360 -11419
rect 9394 -11453 9452 -11419
rect 9486 -11453 9544 -11419
rect 9578 -11453 9636 -11419
rect 9670 -11453 9728 -11419
rect 9762 -11453 9820 -11419
rect 9854 -11453 9912 -11419
rect 9946 -11453 10004 -11419
rect 10038 -11453 10096 -11419
rect 10130 -11453 10188 -11419
rect 10222 -11453 10280 -11419
rect 10314 -11453 10372 -11419
rect 10406 -11453 10464 -11419
rect 10498 -11453 10556 -11419
rect 10590 -11453 10648 -11419
rect 10682 -11453 10740 -11419
rect 10774 -11453 10832 -11419
rect 10866 -11453 10924 -11419
rect 10958 -11453 11016 -11419
rect 11050 -11453 11108 -11419
rect 11142 -11453 11200 -11419
rect 11234 -11453 11292 -11419
rect 11326 -11453 11384 -11419
rect 11418 -11453 11476 -11419
rect 11510 -11453 11568 -11419
rect 11602 -11453 11660 -11419
rect 11694 -11453 11752 -11419
rect 11786 -11453 11844 -11419
rect 11878 -11453 11936 -11419
rect 11970 -11453 12028 -11419
rect 12062 -11453 12120 -11419
rect 12154 -11453 12212 -11419
rect 12246 -11453 12304 -11419
rect 12338 -11453 12396 -11419
rect 12430 -11453 12488 -11419
rect 12522 -11453 12580 -11419
rect 12614 -11453 12672 -11419
rect 12706 -11453 12764 -11419
rect 12798 -11453 12856 -11419
rect 12890 -11453 12948 -11419
rect 12982 -11453 13040 -11419
rect 13074 -11453 13132 -11419
rect 13166 -11453 13224 -11419
rect 13258 -11453 13316 -11419
rect 13350 -11453 13408 -11419
rect 13442 -11453 13500 -11419
rect 13534 -11453 13592 -11419
rect 13626 -11453 13684 -11419
rect 13718 -11453 13776 -11419
rect 13810 -11453 13868 -11419
rect 13902 -11453 13960 -11419
rect 13994 -11453 14052 -11419
rect 14086 -11453 14144 -11419
rect 14178 -11453 14236 -11419
rect 14270 -11453 14328 -11419
rect 14362 -11453 14420 -11419
rect 14454 -11453 14512 -11419
rect 14546 -11453 14604 -11419
rect 14638 -11453 14696 -11419
rect 14730 -11453 14788 -11419
rect 14822 -11453 14880 -11419
rect 14914 -11453 14972 -11419
rect 15006 -11453 15064 -11419
rect 15098 -11453 15156 -11419
rect 15190 -11453 15248 -11419
rect 15282 -11453 15340 -11419
rect 15374 -11453 15432 -11419
rect 15466 -11453 15524 -11419
rect 15558 -11453 15616 -11419
rect 15650 -11453 15708 -11419
rect 15742 -11453 15800 -11419
rect 15834 -11453 15892 -11419
rect 15926 -11453 15984 -11419
rect 16018 -11453 16076 -11419
rect 16110 -11453 16168 -11419
rect 16202 -11453 16260 -11419
rect 16294 -11453 16352 -11419
rect 16386 -11453 16444 -11419
rect 16478 -11453 16536 -11419
rect 16570 -11453 16628 -11419
rect 16662 -11453 16946 -11419
rect -3193 -11484 16946 -11453
rect 12467 -11581 12520 -11556
rect 12467 -11588 12480 -11581
rect 12514 -11588 12520 -11581
rect 12456 -11640 12466 -11588
rect 12518 -11640 12520 -11588
rect 417 -11699 427 -11647
rect 479 -11699 489 -11647
rect 1069 -11651 1127 -11650
rect 3029 -11651 3087 -11650
rect 1069 -11656 3087 -11651
rect 1069 -11690 1081 -11656
rect 1115 -11690 3041 -11656
rect 3075 -11690 3087 -11656
rect 1069 -11695 3087 -11690
rect 1069 -11696 1127 -11695
rect 3029 -11696 3087 -11695
rect 3643 -11651 3701 -11650
rect 5603 -11651 5661 -11650
rect 3643 -11656 5661 -11651
rect 3643 -11690 3655 -11656
rect 3689 -11690 5615 -11656
rect 5649 -11690 5661 -11656
rect 3643 -11695 5661 -11690
rect 3643 -11696 3701 -11695
rect 5603 -11696 5661 -11695
rect 6217 -11651 6275 -11650
rect 8177 -11651 8235 -11650
rect 6217 -11656 8235 -11651
rect 6217 -11690 6229 -11656
rect 6263 -11690 8189 -11656
rect 8223 -11690 8235 -11656
rect 6217 -11695 8235 -11690
rect 6217 -11696 6275 -11695
rect 8177 -11696 8235 -11695
rect 8791 -11651 8849 -11650
rect 10751 -11651 10809 -11650
rect 8791 -11656 10809 -11651
rect 8791 -11690 8806 -11656
rect 8840 -11690 10763 -11656
rect 10797 -11690 10809 -11656
rect 12467 -11653 12520 -11640
rect 13023 -11591 13738 -11584
rect 13023 -11625 13042 -11591
rect 13076 -11624 13738 -11591
rect 13076 -11625 13685 -11624
rect 12745 -11647 12755 -11644
rect 8791 -11695 10809 -11690
rect 8791 -11696 8849 -11695
rect 10751 -11696 10809 -11695
rect 11367 -11735 11377 -11683
rect 11429 -11735 11439 -11683
rect 12467 -11687 12480 -11653
rect 12514 -11687 12520 -11653
rect 12467 -11702 12520 -11687
rect 12548 -11655 12755 -11647
rect 12807 -11647 12817 -11644
rect 12548 -11689 12568 -11655
rect 12602 -11689 12659 -11655
rect 12693 -11689 12755 -11655
rect 12807 -11657 12993 -11647
rect 12548 -11696 12755 -11689
rect 12807 -11691 12858 -11657
rect 12892 -11691 12942 -11657
rect 12976 -11691 12993 -11657
rect 12807 -11696 12993 -11691
rect 13023 -11658 13685 -11625
rect 13719 -11658 13738 -11624
rect 13023 -11668 13738 -11658
rect 12846 -11697 12991 -11696
rect 12456 -11754 12466 -11702
rect 12518 -11754 12520 -11702
rect 13023 -11702 13039 -11668
rect 13073 -11702 13738 -11668
rect 13023 -11707 13738 -11702
rect 15236 -11612 15294 -11606
rect 15329 -11612 15387 -11606
rect 15236 -11646 15248 -11612
rect 15282 -11646 15341 -11612
rect 15375 -11646 15394 -11612
rect 15236 -11688 15394 -11646
rect 13027 -11708 13085 -11707
rect 15236 -11708 16946 -11688
rect 15236 -11742 15248 -11708
rect 15282 -11742 15340 -11708
rect 15374 -11728 16946 -11708
rect 15374 -11742 15394 -11728
rect 15236 -11748 15294 -11742
rect 15328 -11748 15386 -11742
rect 12467 -11761 12480 -11754
rect 12514 -11761 12520 -11754
rect 12467 -11793 12520 -11761
rect -3193 -11963 16946 -11932
rect -3193 -11997 -2968 -11963
rect -2934 -11997 -2876 -11963
rect -2842 -11997 -2784 -11963
rect -2750 -11997 -2692 -11963
rect -2658 -11997 -2600 -11963
rect -2566 -11997 -2508 -11963
rect -2474 -11997 -2416 -11963
rect -2382 -11997 -2324 -11963
rect -2290 -11997 -2232 -11963
rect -2198 -11997 -2140 -11963
rect -2106 -11997 -2048 -11963
rect -2014 -11997 -1956 -11963
rect -1922 -11997 -1864 -11963
rect -1830 -11997 -1772 -11963
rect -1738 -11997 -1680 -11963
rect -1646 -11997 -1588 -11963
rect -1554 -11997 -1496 -11963
rect -1462 -11997 -1404 -11963
rect -1370 -11997 -1312 -11963
rect -1278 -11997 -1220 -11963
rect -1186 -11997 -1128 -11963
rect -1094 -11997 -1036 -11963
rect -1002 -11997 -944 -11963
rect -910 -11997 -852 -11963
rect -818 -11997 -760 -11963
rect -726 -11997 -668 -11963
rect -634 -11997 -576 -11963
rect -542 -11997 -484 -11963
rect -450 -11997 -392 -11963
rect -358 -11997 -300 -11963
rect -266 -11997 -208 -11963
rect -174 -11997 -116 -11963
rect -82 -11997 -24 -11963
rect 10 -11997 68 -11963
rect 102 -11997 160 -11963
rect 194 -11997 252 -11963
rect 286 -11997 344 -11963
rect 378 -11997 436 -11963
rect 470 -11997 528 -11963
rect 562 -11997 620 -11963
rect 654 -11997 712 -11963
rect 746 -11997 804 -11963
rect 838 -11997 896 -11963
rect 930 -11997 988 -11963
rect 1022 -11997 1080 -11963
rect 1114 -11997 1172 -11963
rect 1206 -11997 1264 -11963
rect 1298 -11997 1356 -11963
rect 1390 -11997 1448 -11963
rect 1482 -11997 1540 -11963
rect 1574 -11997 1632 -11963
rect 1666 -11997 1724 -11963
rect 1758 -11997 1816 -11963
rect 1850 -11997 1908 -11963
rect 1942 -11997 2000 -11963
rect 2034 -11997 2092 -11963
rect 2126 -11997 2184 -11963
rect 2218 -11997 2276 -11963
rect 2310 -11997 2368 -11963
rect 2402 -11997 2460 -11963
rect 2494 -11997 2552 -11963
rect 2586 -11997 2644 -11963
rect 2678 -11997 2736 -11963
rect 2770 -11997 2828 -11963
rect 2862 -11997 2920 -11963
rect 2954 -11997 3012 -11963
rect 3046 -11997 3104 -11963
rect 3138 -11997 3196 -11963
rect 3230 -11997 3288 -11963
rect 3322 -11997 3380 -11963
rect 3414 -11997 3472 -11963
rect 3506 -11997 3564 -11963
rect 3598 -11997 3656 -11963
rect 3690 -11997 3748 -11963
rect 3782 -11997 3840 -11963
rect 3874 -11997 3932 -11963
rect 3966 -11997 4024 -11963
rect 4058 -11997 4116 -11963
rect 4150 -11997 4208 -11963
rect 4242 -11997 4300 -11963
rect 4334 -11997 4392 -11963
rect 4426 -11997 4484 -11963
rect 4518 -11997 4576 -11963
rect 4610 -11997 4668 -11963
rect 4702 -11997 4760 -11963
rect 4794 -11997 4852 -11963
rect 4886 -11997 4944 -11963
rect 4978 -11997 5036 -11963
rect 5070 -11997 5128 -11963
rect 5162 -11997 5220 -11963
rect 5254 -11997 5312 -11963
rect 5346 -11997 5404 -11963
rect 5438 -11997 5496 -11963
rect 5530 -11997 5588 -11963
rect 5622 -11997 5680 -11963
rect 5714 -11997 5772 -11963
rect 5806 -11997 5864 -11963
rect 5898 -11997 5956 -11963
rect 5990 -11997 6048 -11963
rect 6082 -11997 6140 -11963
rect 6174 -11997 6232 -11963
rect 6266 -11997 6324 -11963
rect 6358 -11997 6416 -11963
rect 6450 -11997 6508 -11963
rect 6542 -11997 6600 -11963
rect 6634 -11997 6692 -11963
rect 6726 -11997 6784 -11963
rect 6818 -11997 6876 -11963
rect 6910 -11997 6968 -11963
rect 7002 -11997 7060 -11963
rect 7094 -11997 7152 -11963
rect 7186 -11997 7244 -11963
rect 7278 -11997 7336 -11963
rect 7370 -11997 7428 -11963
rect 7462 -11997 7520 -11963
rect 7554 -11997 7612 -11963
rect 7646 -11997 7704 -11963
rect 7738 -11997 7796 -11963
rect 7830 -11997 7888 -11963
rect 7922 -11997 7980 -11963
rect 8014 -11997 8072 -11963
rect 8106 -11997 8164 -11963
rect 8198 -11997 8256 -11963
rect 8290 -11997 8348 -11963
rect 8382 -11997 8440 -11963
rect 8474 -11997 8532 -11963
rect 8566 -11997 8624 -11963
rect 8658 -11997 8716 -11963
rect 8750 -11997 8808 -11963
rect 8842 -11997 8900 -11963
rect 8934 -11997 8992 -11963
rect 9026 -11997 9084 -11963
rect 9118 -11997 9176 -11963
rect 9210 -11997 9268 -11963
rect 9302 -11997 9360 -11963
rect 9394 -11997 9452 -11963
rect 9486 -11997 9544 -11963
rect 9578 -11997 9636 -11963
rect 9670 -11997 9728 -11963
rect 9762 -11997 9820 -11963
rect 9854 -11997 9912 -11963
rect 9946 -11997 10004 -11963
rect 10038 -11997 10096 -11963
rect 10130 -11997 10188 -11963
rect 10222 -11997 10280 -11963
rect 10314 -11997 10372 -11963
rect 10406 -11997 10464 -11963
rect 10498 -11997 10556 -11963
rect 10590 -11997 10648 -11963
rect 10682 -11997 10740 -11963
rect 10774 -11997 10832 -11963
rect 10866 -11997 10924 -11963
rect 10958 -11997 11016 -11963
rect 11050 -11997 11108 -11963
rect 11142 -11997 11200 -11963
rect 11234 -11997 11292 -11963
rect 11326 -11997 11384 -11963
rect 11418 -11997 11476 -11963
rect 11510 -11997 11568 -11963
rect 11602 -11997 11660 -11963
rect 11694 -11997 11752 -11963
rect 11786 -11997 11844 -11963
rect 11878 -11997 11936 -11963
rect 11970 -11997 12028 -11963
rect 12062 -11997 12120 -11963
rect 12154 -11997 12212 -11963
rect 12246 -11997 12304 -11963
rect 12338 -11997 12396 -11963
rect 12430 -11997 12488 -11963
rect 12522 -11997 12580 -11963
rect 12614 -11997 12672 -11963
rect 12706 -11997 12764 -11963
rect 12798 -11997 12856 -11963
rect 12890 -11997 12948 -11963
rect 12982 -11997 13040 -11963
rect 13074 -11997 13132 -11963
rect 13166 -11997 13224 -11963
rect 13258 -11997 13316 -11963
rect 13350 -11997 13408 -11963
rect 13442 -11997 13500 -11963
rect 13534 -11997 13592 -11963
rect 13626 -11997 13684 -11963
rect 13718 -11997 13776 -11963
rect 13810 -11997 13868 -11963
rect 13902 -11997 13960 -11963
rect 13994 -11997 14052 -11963
rect 14086 -11997 14144 -11963
rect 14178 -11997 14236 -11963
rect 14270 -11997 14328 -11963
rect 14362 -11997 14420 -11963
rect 14454 -11997 14512 -11963
rect 14546 -11997 14604 -11963
rect 14638 -11997 14696 -11963
rect 14730 -11997 14788 -11963
rect 14822 -11997 14880 -11963
rect 14914 -11997 14972 -11963
rect 15006 -11997 15064 -11963
rect 15098 -11997 15156 -11963
rect 15190 -11997 15248 -11963
rect 15282 -11997 15340 -11963
rect 15374 -11997 15432 -11963
rect 15466 -11997 15524 -11963
rect 15558 -11997 15616 -11963
rect 15650 -11997 15708 -11963
rect 15742 -11997 15800 -11963
rect 15834 -11997 15892 -11963
rect 15926 -11997 15984 -11963
rect 16018 -11997 16076 -11963
rect 16110 -11997 16168 -11963
rect 16202 -11997 16260 -11963
rect 16294 -11997 16352 -11963
rect 16386 -11997 16444 -11963
rect 16478 -11997 16536 -11963
rect 16570 -11997 16628 -11963
rect 16662 -11997 16946 -11963
rect -3193 -12028 16946 -11997
rect 15236 -12222 15294 -12216
rect 15329 -12222 15387 -12216
rect -866 -12229 -404 -12224
rect -867 -12235 -404 -12229
rect -867 -12269 -855 -12235
rect -821 -12269 -404 -12235
rect -867 -12275 -404 -12269
rect -866 -12282 -404 -12275
rect -346 -12282 -336 -12224
rect 105 -12263 115 -12259
rect -253 -12272 115 -12263
rect -253 -12306 -210 -12272
rect -176 -12306 115 -12272
rect -253 -12309 115 -12306
rect -222 -12312 -164 -12309
rect 105 -12311 115 -12309
rect 167 -12311 177 -12259
rect 414 -12278 424 -12226
rect 476 -12278 486 -12226
rect 15236 -12256 15248 -12222
rect 15282 -12256 15341 -12222
rect 15375 -12232 15394 -12222
rect 15375 -12256 16946 -12232
rect 1042 -12263 1100 -12262
rect 3002 -12263 3060 -12262
rect 1042 -12268 3060 -12263
rect 1042 -12302 1054 -12268
rect 1088 -12302 3014 -12268
rect 3048 -12302 3060 -12268
rect 1042 -12307 3060 -12302
rect 1042 -12308 1100 -12307
rect 3002 -12308 3060 -12307
rect 3616 -12263 3674 -12262
rect 5576 -12263 5634 -12262
rect 3616 -12268 5634 -12263
rect 3616 -12302 3628 -12268
rect 3662 -12302 5588 -12268
rect 5622 -12302 5634 -12268
rect 3616 -12307 5634 -12302
rect 3616 -12308 3674 -12307
rect 5576 -12308 5634 -12307
rect 6190 -12263 6248 -12262
rect 8150 -12263 8208 -12262
rect 6190 -12268 8208 -12263
rect 6190 -12302 6202 -12268
rect 6236 -12302 8162 -12268
rect 8196 -12302 8208 -12268
rect 6190 -12307 8208 -12302
rect 6190 -12308 6248 -12307
rect 8150 -12308 8208 -12307
rect 8764 -12263 8822 -12262
rect 10724 -12263 10782 -12262
rect 8764 -12268 10782 -12263
rect 8764 -12302 8776 -12268
rect 8810 -12302 10736 -12268
rect 10770 -12302 10782 -12268
rect 8764 -12307 10782 -12302
rect 8764 -12308 8822 -12307
rect 10724 -12308 10782 -12307
rect 11365 -12313 11375 -12261
rect 11427 -12313 11437 -12261
rect 13671 -12302 13735 -12258
rect 13671 -12336 13685 -12302
rect 13719 -12336 13735 -12302
rect 12746 -12352 12756 -12350
rect 7153 -12353 12756 -12352
rect 7153 -12405 7163 -12353
rect 7215 -12402 12756 -12353
rect 12808 -12352 12818 -12350
rect 13671 -12352 13735 -12336
rect 12808 -12402 13735 -12352
rect 15236 -12272 16946 -12256
rect 15236 -12317 15394 -12272
rect 15236 -12318 15340 -12317
rect 15236 -12352 15248 -12318
rect 15282 -12351 15340 -12318
rect 15374 -12351 15394 -12317
rect 15282 -12352 15394 -12351
rect 15236 -12358 15294 -12352
rect 15328 -12357 15386 -12352
rect 7215 -12405 13735 -12402
rect 7153 -12406 13735 -12405
rect 13671 -12407 13735 -12406
rect -3193 -12507 16946 -12476
rect -3193 -12541 -2968 -12507
rect -2934 -12541 -2876 -12507
rect -2842 -12541 -2784 -12507
rect -2750 -12541 -2692 -12507
rect -2658 -12541 -2600 -12507
rect -2566 -12541 -2508 -12507
rect -2474 -12541 -2416 -12507
rect -2382 -12541 -2324 -12507
rect -2290 -12541 -2232 -12507
rect -2198 -12541 -2140 -12507
rect -2106 -12541 -2048 -12507
rect -2014 -12541 -1956 -12507
rect -1922 -12541 -1864 -12507
rect -1830 -12541 -1772 -12507
rect -1738 -12541 -1680 -12507
rect -1646 -12541 -1588 -12507
rect -1554 -12541 -1496 -12507
rect -1462 -12541 -1404 -12507
rect -1370 -12541 -1312 -12507
rect -1278 -12541 -1220 -12507
rect -1186 -12541 -1128 -12507
rect -1094 -12541 -1036 -12507
rect -1002 -12541 -944 -12507
rect -910 -12541 -852 -12507
rect -818 -12541 -760 -12507
rect -726 -12541 -668 -12507
rect -634 -12541 -576 -12507
rect -542 -12541 -484 -12507
rect -450 -12541 -392 -12507
rect -358 -12541 -300 -12507
rect -266 -12541 -208 -12507
rect -174 -12541 -116 -12507
rect -82 -12541 -24 -12507
rect 10 -12541 68 -12507
rect 102 -12541 160 -12507
rect 194 -12541 252 -12507
rect 286 -12541 344 -12507
rect 378 -12541 436 -12507
rect 470 -12541 528 -12507
rect 562 -12541 620 -12507
rect 654 -12541 712 -12507
rect 746 -12541 804 -12507
rect 838 -12541 896 -12507
rect 930 -12541 988 -12507
rect 1022 -12541 1080 -12507
rect 1114 -12541 1172 -12507
rect 1206 -12541 1264 -12507
rect 1298 -12541 1356 -12507
rect 1390 -12541 1448 -12507
rect 1482 -12541 1540 -12507
rect 1574 -12541 1632 -12507
rect 1666 -12541 1724 -12507
rect 1758 -12541 1816 -12507
rect 1850 -12541 1908 -12507
rect 1942 -12541 2000 -12507
rect 2034 -12541 2092 -12507
rect 2126 -12541 2184 -12507
rect 2218 -12541 2276 -12507
rect 2310 -12541 2368 -12507
rect 2402 -12541 2460 -12507
rect 2494 -12541 2552 -12507
rect 2586 -12541 2644 -12507
rect 2678 -12541 2736 -12507
rect 2770 -12541 2828 -12507
rect 2862 -12541 2920 -12507
rect 2954 -12541 3012 -12507
rect 3046 -12541 3104 -12507
rect 3138 -12541 3196 -12507
rect 3230 -12541 3288 -12507
rect 3322 -12541 3380 -12507
rect 3414 -12541 3472 -12507
rect 3506 -12541 3564 -12507
rect 3598 -12541 3656 -12507
rect 3690 -12541 3748 -12507
rect 3782 -12541 3840 -12507
rect 3874 -12541 3932 -12507
rect 3966 -12541 4024 -12507
rect 4058 -12541 4116 -12507
rect 4150 -12541 4208 -12507
rect 4242 -12541 4300 -12507
rect 4334 -12541 4392 -12507
rect 4426 -12541 4484 -12507
rect 4518 -12541 4576 -12507
rect 4610 -12541 4668 -12507
rect 4702 -12541 4760 -12507
rect 4794 -12541 4852 -12507
rect 4886 -12541 4944 -12507
rect 4978 -12541 5036 -12507
rect 5070 -12541 5128 -12507
rect 5162 -12541 5220 -12507
rect 5254 -12541 5312 -12507
rect 5346 -12541 5404 -12507
rect 5438 -12541 5496 -12507
rect 5530 -12541 5588 -12507
rect 5622 -12541 5680 -12507
rect 5714 -12541 5772 -12507
rect 5806 -12541 5864 -12507
rect 5898 -12541 5956 -12507
rect 5990 -12541 6048 -12507
rect 6082 -12541 6140 -12507
rect 6174 -12541 6232 -12507
rect 6266 -12541 6324 -12507
rect 6358 -12541 6416 -12507
rect 6450 -12541 6508 -12507
rect 6542 -12541 6600 -12507
rect 6634 -12541 6692 -12507
rect 6726 -12541 6784 -12507
rect 6818 -12541 6876 -12507
rect 6910 -12541 6968 -12507
rect 7002 -12541 7060 -12507
rect 7094 -12541 7152 -12507
rect 7186 -12541 7244 -12507
rect 7278 -12541 7336 -12507
rect 7370 -12541 7428 -12507
rect 7462 -12541 7520 -12507
rect 7554 -12541 7612 -12507
rect 7646 -12541 7704 -12507
rect 7738 -12541 7796 -12507
rect 7830 -12541 7888 -12507
rect 7922 -12541 7980 -12507
rect 8014 -12541 8072 -12507
rect 8106 -12541 8164 -12507
rect 8198 -12541 8256 -12507
rect 8290 -12541 8348 -12507
rect 8382 -12541 8440 -12507
rect 8474 -12541 8532 -12507
rect 8566 -12541 8624 -12507
rect 8658 -12541 8716 -12507
rect 8750 -12541 8808 -12507
rect 8842 -12541 8900 -12507
rect 8934 -12541 8992 -12507
rect 9026 -12541 9084 -12507
rect 9118 -12541 9176 -12507
rect 9210 -12541 9268 -12507
rect 9302 -12541 9360 -12507
rect 9394 -12541 9452 -12507
rect 9486 -12541 9544 -12507
rect 9578 -12541 9636 -12507
rect 9670 -12541 9728 -12507
rect 9762 -12541 9820 -12507
rect 9854 -12541 9912 -12507
rect 9946 -12541 10004 -12507
rect 10038 -12541 10096 -12507
rect 10130 -12541 10188 -12507
rect 10222 -12541 10280 -12507
rect 10314 -12541 10372 -12507
rect 10406 -12541 10464 -12507
rect 10498 -12541 10556 -12507
rect 10590 -12541 10648 -12507
rect 10682 -12541 10740 -12507
rect 10774 -12541 10832 -12507
rect 10866 -12541 10924 -12507
rect 10958 -12541 11016 -12507
rect 11050 -12541 11108 -12507
rect 11142 -12541 11200 -12507
rect 11234 -12541 11292 -12507
rect 11326 -12541 11384 -12507
rect 11418 -12541 11476 -12507
rect 11510 -12541 11568 -12507
rect 11602 -12541 11660 -12507
rect 11694 -12541 11752 -12507
rect 11786 -12541 11844 -12507
rect 11878 -12541 11936 -12507
rect 11970 -12541 12028 -12507
rect 12062 -12541 12120 -12507
rect 12154 -12541 12212 -12507
rect 12246 -12541 12304 -12507
rect 12338 -12541 12396 -12507
rect 12430 -12541 12488 -12507
rect 12522 -12541 12580 -12507
rect 12614 -12541 12672 -12507
rect 12706 -12541 12764 -12507
rect 12798 -12541 12856 -12507
rect 12890 -12541 12948 -12507
rect 12982 -12541 13040 -12507
rect 13074 -12541 13132 -12507
rect 13166 -12541 13224 -12507
rect 13258 -12541 13316 -12507
rect 13350 -12541 13408 -12507
rect 13442 -12541 13500 -12507
rect 13534 -12541 13592 -12507
rect 13626 -12541 13684 -12507
rect 13718 -12541 13776 -12507
rect 13810 -12541 13868 -12507
rect 13902 -12541 13960 -12507
rect 13994 -12541 14052 -12507
rect 14086 -12541 14144 -12507
rect 14178 -12541 14236 -12507
rect 14270 -12541 14328 -12507
rect 14362 -12541 14420 -12507
rect 14454 -12541 14512 -12507
rect 14546 -12541 14604 -12507
rect 14638 -12541 14696 -12507
rect 14730 -12541 14788 -12507
rect 14822 -12541 14880 -12507
rect 14914 -12541 14972 -12507
rect 15006 -12541 15064 -12507
rect 15098 -12541 15156 -12507
rect 15190 -12541 15248 -12507
rect 15282 -12541 15340 -12507
rect 15374 -12541 15432 -12507
rect 15466 -12541 15524 -12507
rect 15558 -12541 15616 -12507
rect 15650 -12541 15708 -12507
rect 15742 -12541 15800 -12507
rect 15834 -12541 15892 -12507
rect 15926 -12541 15984 -12507
rect 16018 -12541 16076 -12507
rect 16110 -12541 16168 -12507
rect 16202 -12541 16260 -12507
rect 16294 -12541 16352 -12507
rect 16386 -12541 16444 -12507
rect 16478 -12541 16536 -12507
rect 16570 -12541 16628 -12507
rect 16662 -12541 16946 -12507
rect -3193 -12572 16946 -12541
rect 13026 -12677 13084 -12670
rect 13026 -12711 13038 -12677
rect 13072 -12678 13084 -12677
rect 13072 -12711 13737 -12678
rect 13026 -12712 13737 -12711
rect 12548 -12734 12992 -12733
rect 12548 -12736 12752 -12734
rect 417 -12788 427 -12736
rect 479 -12788 489 -12736
rect 1070 -12740 1128 -12739
rect 3030 -12740 3088 -12739
rect 1070 -12745 3088 -12740
rect 1070 -12779 1082 -12745
rect 1116 -12779 3042 -12745
rect 3076 -12779 3088 -12745
rect 1070 -12784 3088 -12779
rect 1070 -12785 1128 -12784
rect 3030 -12785 3088 -12784
rect 3644 -12740 3702 -12739
rect 5604 -12740 5662 -12739
rect 3644 -12745 5662 -12740
rect 3644 -12779 3656 -12745
rect 3690 -12779 5616 -12745
rect 5650 -12779 5662 -12745
rect 3644 -12784 5662 -12779
rect 3644 -12785 3702 -12784
rect 5604 -12785 5662 -12784
rect 6218 -12740 6276 -12739
rect 8178 -12740 8236 -12739
rect 6218 -12745 8236 -12740
rect 6218 -12779 6230 -12745
rect 6264 -12779 8190 -12745
rect 8224 -12779 8236 -12745
rect 6218 -12784 8236 -12779
rect 6218 -12785 6276 -12784
rect 8178 -12785 8236 -12784
rect 8792 -12740 8850 -12739
rect 10752 -12740 10810 -12739
rect 8792 -12745 10810 -12740
rect 8792 -12779 8804 -12745
rect 8838 -12779 10764 -12745
rect 10798 -12779 10810 -12745
rect 12546 -12742 12752 -12736
rect 12804 -12742 12992 -12734
rect 8792 -12784 10810 -12779
rect 8792 -12785 8850 -12784
rect 10752 -12785 10810 -12784
rect 11370 -12820 11380 -12768
rect 11432 -12820 11442 -12768
rect 12546 -12776 12558 -12742
rect 12592 -12776 12642 -12742
rect 12676 -12776 12739 -12742
rect 12804 -12776 12836 -12742
rect 12870 -12776 12942 -12742
rect 12976 -12776 12992 -12742
rect 12546 -12782 12752 -12776
rect 12548 -12786 12752 -12782
rect 12804 -12786 12992 -12776
rect 13026 -12746 13684 -12712
rect 13718 -12746 13737 -12712
rect 13026 -12749 13737 -12746
rect 13026 -12783 13038 -12749
rect 13072 -12783 13737 -12749
rect 13026 -12788 13737 -12783
rect 15236 -12700 15294 -12694
rect 15329 -12700 15387 -12694
rect 15236 -12734 15248 -12700
rect 15282 -12734 15341 -12700
rect 15375 -12734 15394 -12700
rect 15236 -12776 15394 -12734
rect 13026 -12789 13084 -12788
rect 15236 -12795 16946 -12776
rect 15236 -12796 15340 -12795
rect 15236 -12830 15248 -12796
rect 15282 -12829 15340 -12796
rect 15374 -12816 16946 -12795
rect 15374 -12829 15394 -12816
rect 15282 -12830 15394 -12829
rect 15236 -12836 15294 -12830
rect 15328 -12835 15386 -12830
rect 7161 -12881 11181 -12875
rect 7155 -12933 7165 -12881
rect 7217 -12884 11181 -12881
rect 7217 -12933 11118 -12884
rect 7161 -12936 11118 -12933
rect 11170 -12936 11181 -12884
rect 7161 -12937 11181 -12936
rect -3193 -13051 16946 -13020
rect -3193 -13085 -2968 -13051
rect -2934 -13085 -2876 -13051
rect -2842 -13085 -2784 -13051
rect -2750 -13085 -2692 -13051
rect -2658 -13085 -2600 -13051
rect -2566 -13085 -2508 -13051
rect -2474 -13085 -2416 -13051
rect -2382 -13085 -2324 -13051
rect -2290 -13085 -2232 -13051
rect -2198 -13085 -2140 -13051
rect -2106 -13085 -2048 -13051
rect -2014 -13085 -1956 -13051
rect -1922 -13085 -1864 -13051
rect -1830 -13085 -1772 -13051
rect -1738 -13085 -1680 -13051
rect -1646 -13085 -1588 -13051
rect -1554 -13085 -1496 -13051
rect -1462 -13085 -1404 -13051
rect -1370 -13085 -1312 -13051
rect -1278 -13085 -1220 -13051
rect -1186 -13085 -1128 -13051
rect -1094 -13085 -1036 -13051
rect -1002 -13085 -944 -13051
rect -910 -13085 -852 -13051
rect -818 -13085 -760 -13051
rect -726 -13085 -668 -13051
rect -634 -13085 -576 -13051
rect -542 -13085 -484 -13051
rect -450 -13085 -392 -13051
rect -358 -13085 -300 -13051
rect -266 -13085 -208 -13051
rect -174 -13085 -116 -13051
rect -82 -13085 -24 -13051
rect 10 -13085 68 -13051
rect 102 -13085 160 -13051
rect 194 -13085 252 -13051
rect 286 -13085 344 -13051
rect 378 -13085 436 -13051
rect 470 -13085 528 -13051
rect 562 -13085 620 -13051
rect 654 -13085 712 -13051
rect 746 -13085 804 -13051
rect 838 -13085 896 -13051
rect 930 -13085 988 -13051
rect 1022 -13085 1080 -13051
rect 1114 -13085 1172 -13051
rect 1206 -13085 1264 -13051
rect 1298 -13085 1356 -13051
rect 1390 -13085 1448 -13051
rect 1482 -13085 1540 -13051
rect 1574 -13085 1632 -13051
rect 1666 -13085 1724 -13051
rect 1758 -13085 1816 -13051
rect 1850 -13085 1908 -13051
rect 1942 -13085 2000 -13051
rect 2034 -13085 2092 -13051
rect 2126 -13085 2184 -13051
rect 2218 -13085 2276 -13051
rect 2310 -13085 2368 -13051
rect 2402 -13085 2460 -13051
rect 2494 -13085 2552 -13051
rect 2586 -13085 2644 -13051
rect 2678 -13085 2736 -13051
rect 2770 -13085 2828 -13051
rect 2862 -13085 2920 -13051
rect 2954 -13085 3012 -13051
rect 3046 -13085 3104 -13051
rect 3138 -13085 3196 -13051
rect 3230 -13085 3288 -13051
rect 3322 -13085 3380 -13051
rect 3414 -13085 3472 -13051
rect 3506 -13085 3564 -13051
rect 3598 -13085 3656 -13051
rect 3690 -13085 3748 -13051
rect 3782 -13085 3840 -13051
rect 3874 -13085 3932 -13051
rect 3966 -13085 4024 -13051
rect 4058 -13085 4116 -13051
rect 4150 -13085 4208 -13051
rect 4242 -13085 4300 -13051
rect 4334 -13085 4392 -13051
rect 4426 -13085 4484 -13051
rect 4518 -13085 4576 -13051
rect 4610 -13085 4668 -13051
rect 4702 -13085 4760 -13051
rect 4794 -13085 4852 -13051
rect 4886 -13085 4944 -13051
rect 4978 -13085 5036 -13051
rect 5070 -13085 5128 -13051
rect 5162 -13085 5220 -13051
rect 5254 -13085 5312 -13051
rect 5346 -13085 5404 -13051
rect 5438 -13085 5496 -13051
rect 5530 -13085 5588 -13051
rect 5622 -13085 5680 -13051
rect 5714 -13085 5772 -13051
rect 5806 -13085 5864 -13051
rect 5898 -13085 5956 -13051
rect 5990 -13085 6048 -13051
rect 6082 -13085 6140 -13051
rect 6174 -13085 6232 -13051
rect 6266 -13085 6324 -13051
rect 6358 -13085 6416 -13051
rect 6450 -13085 6508 -13051
rect 6542 -13085 6600 -13051
rect 6634 -13085 6692 -13051
rect 6726 -13085 6784 -13051
rect 6818 -13085 6876 -13051
rect 6910 -13085 6968 -13051
rect 7002 -13085 7060 -13051
rect 7094 -13085 7152 -13051
rect 7186 -13085 7244 -13051
rect 7278 -13085 7336 -13051
rect 7370 -13085 7428 -13051
rect 7462 -13085 7520 -13051
rect 7554 -13085 7612 -13051
rect 7646 -13085 7704 -13051
rect 7738 -13085 7796 -13051
rect 7830 -13085 7888 -13051
rect 7922 -13085 7980 -13051
rect 8014 -13085 8072 -13051
rect 8106 -13085 8164 -13051
rect 8198 -13085 8256 -13051
rect 8290 -13085 8348 -13051
rect 8382 -13085 8440 -13051
rect 8474 -13085 8532 -13051
rect 8566 -13085 8624 -13051
rect 8658 -13085 8716 -13051
rect 8750 -13085 8808 -13051
rect 8842 -13085 8900 -13051
rect 8934 -13085 8992 -13051
rect 9026 -13085 9084 -13051
rect 9118 -13085 9176 -13051
rect 9210 -13085 9268 -13051
rect 9302 -13085 9360 -13051
rect 9394 -13085 9452 -13051
rect 9486 -13085 9544 -13051
rect 9578 -13085 9636 -13051
rect 9670 -13085 9728 -13051
rect 9762 -13085 9820 -13051
rect 9854 -13085 9912 -13051
rect 9946 -13085 10004 -13051
rect 10038 -13085 10096 -13051
rect 10130 -13085 10188 -13051
rect 10222 -13085 10280 -13051
rect 10314 -13085 10372 -13051
rect 10406 -13085 10464 -13051
rect 10498 -13085 10556 -13051
rect 10590 -13085 10648 -13051
rect 10682 -13085 10740 -13051
rect 10774 -13085 10832 -13051
rect 10866 -13085 10924 -13051
rect 10958 -13085 11016 -13051
rect 11050 -13085 11108 -13051
rect 11142 -13085 11200 -13051
rect 11234 -13085 11292 -13051
rect 11326 -13085 11384 -13051
rect 11418 -13085 11476 -13051
rect 11510 -13085 11568 -13051
rect 11602 -13085 11660 -13051
rect 11694 -13085 11752 -13051
rect 11786 -13085 11844 -13051
rect 11878 -13085 11936 -13051
rect 11970 -13085 12028 -13051
rect 12062 -13085 12120 -13051
rect 12154 -13085 12212 -13051
rect 12246 -13085 12304 -13051
rect 12338 -13085 12396 -13051
rect 12430 -13085 12488 -13051
rect 12522 -13085 12580 -13051
rect 12614 -13085 12672 -13051
rect 12706 -13085 12764 -13051
rect 12798 -13085 12856 -13051
rect 12890 -13085 12948 -13051
rect 12982 -13085 13040 -13051
rect 13074 -13085 13132 -13051
rect 13166 -13085 13224 -13051
rect 13258 -13085 13316 -13051
rect 13350 -13085 13408 -13051
rect 13442 -13085 13500 -13051
rect 13534 -13085 13592 -13051
rect 13626 -13085 13684 -13051
rect 13718 -13085 13776 -13051
rect 13810 -13085 13868 -13051
rect 13902 -13085 13960 -13051
rect 13994 -13085 14052 -13051
rect 14086 -13085 14144 -13051
rect 14178 -13085 14236 -13051
rect 14270 -13085 14328 -13051
rect 14362 -13085 14420 -13051
rect 14454 -13085 14512 -13051
rect 14546 -13085 14604 -13051
rect 14638 -13085 14696 -13051
rect 14730 -13085 14788 -13051
rect 14822 -13085 14880 -13051
rect 14914 -13085 14972 -13051
rect 15006 -13085 15064 -13051
rect 15098 -13085 15156 -13051
rect 15190 -13085 15248 -13051
rect 15282 -13085 15340 -13051
rect 15374 -13085 15432 -13051
rect 15466 -13085 15524 -13051
rect 15558 -13085 15616 -13051
rect 15650 -13085 15708 -13051
rect 15742 -13085 15800 -13051
rect 15834 -13085 15892 -13051
rect 15926 -13085 15984 -13051
rect 16018 -13085 16076 -13051
rect 16110 -13085 16168 -13051
rect 16202 -13085 16260 -13051
rect 16294 -13085 16352 -13051
rect 16386 -13085 16444 -13051
rect 16478 -13085 16536 -13051
rect 16570 -13085 16628 -13051
rect 16662 -13085 16946 -13051
rect -3193 -13116 16946 -13085
rect 11339 -13285 12463 -13281
rect 412 -13367 422 -13315
rect 474 -13367 484 -13315
rect 11338 -13340 12463 -13285
rect 12522 -13340 12532 -13281
rect 15236 -13310 15294 -13304
rect 15329 -13310 15387 -13304
rect 10725 -13353 10783 -13351
rect 1040 -13354 1098 -13353
rect 3000 -13354 3058 -13353
rect 1040 -13359 3058 -13354
rect 1040 -13393 1052 -13359
rect 1086 -13393 3012 -13359
rect 3046 -13393 3058 -13359
rect 1040 -13398 3058 -13393
rect 1040 -13399 1098 -13398
rect 3000 -13399 3058 -13398
rect 3614 -13354 3672 -13353
rect 5574 -13354 5632 -13353
rect 3614 -13359 5632 -13354
rect 3614 -13393 3626 -13359
rect 3660 -13393 5586 -13359
rect 5620 -13393 5632 -13359
rect 3614 -13398 5632 -13393
rect 3614 -13399 3672 -13398
rect 5574 -13399 5632 -13398
rect 6188 -13354 6246 -13353
rect 8148 -13354 8206 -13353
rect 6188 -13359 8206 -13354
rect 6188 -13393 6200 -13359
rect 6234 -13393 8160 -13359
rect 8194 -13393 8206 -13359
rect 6188 -13398 8206 -13393
rect 6188 -13399 6246 -13398
rect 8148 -13399 8206 -13398
rect 8762 -13354 8820 -13353
rect 10139 -13354 10783 -13353
rect 8762 -13357 10783 -13354
rect 8762 -13359 10737 -13357
rect 8762 -13393 8774 -13359
rect 8808 -13391 10737 -13359
rect 10771 -13391 10783 -13357
rect 8808 -13393 10783 -13391
rect 8762 -13397 10783 -13393
rect 11338 -13356 11430 -13340
rect 15236 -13344 15248 -13310
rect 15282 -13344 15341 -13310
rect 15375 -13320 15394 -13310
rect 15375 -13344 16946 -13320
rect 11338 -13390 11369 -13356
rect 11403 -13390 11430 -13356
rect 11338 -13397 11430 -13390
rect 13669 -13388 13738 -13345
rect 8762 -13398 10273 -13397
rect 8762 -13399 8820 -13398
rect 13669 -13422 13685 -13388
rect 13719 -13422 13738 -13388
rect 13669 -13432 13738 -13422
rect 966 -13434 13738 -13432
rect 966 -13435 12753 -13434
rect 966 -13487 982 -13435
rect 1034 -13486 12753 -13435
rect 12805 -13486 13738 -13434
rect 15236 -13360 16946 -13344
rect 15236 -13405 15394 -13360
rect 15236 -13406 15340 -13405
rect 15236 -13440 15248 -13406
rect 15282 -13439 15340 -13406
rect 15374 -13439 15394 -13405
rect 15282 -13440 15394 -13439
rect 15236 -13446 15294 -13440
rect 15328 -13445 15386 -13440
rect 1034 -13487 13738 -13486
rect 13669 -13489 13738 -13487
rect -3193 -13595 16946 -13564
rect -3193 -13629 -2968 -13595
rect -2934 -13629 -2876 -13595
rect -2842 -13629 -2784 -13595
rect -2750 -13629 -2692 -13595
rect -2658 -13629 -2600 -13595
rect -2566 -13629 -2508 -13595
rect -2474 -13629 -2416 -13595
rect -2382 -13629 -2324 -13595
rect -2290 -13629 -2232 -13595
rect -2198 -13629 -2140 -13595
rect -2106 -13629 -2048 -13595
rect -2014 -13629 -1956 -13595
rect -1922 -13629 -1864 -13595
rect -1830 -13629 -1772 -13595
rect -1738 -13629 -1680 -13595
rect -1646 -13629 -1588 -13595
rect -1554 -13629 -1496 -13595
rect -1462 -13629 -1404 -13595
rect -1370 -13629 -1312 -13595
rect -1278 -13629 -1220 -13595
rect -1186 -13629 -1128 -13595
rect -1094 -13629 -1036 -13595
rect -1002 -13629 -944 -13595
rect -910 -13629 -852 -13595
rect -818 -13629 -760 -13595
rect -726 -13629 -668 -13595
rect -634 -13629 -576 -13595
rect -542 -13629 -484 -13595
rect -450 -13629 -392 -13595
rect -358 -13629 -300 -13595
rect -266 -13629 -208 -13595
rect -174 -13629 -116 -13595
rect -82 -13629 -24 -13595
rect 10 -13629 68 -13595
rect 102 -13629 160 -13595
rect 194 -13629 252 -13595
rect 286 -13629 344 -13595
rect 378 -13629 436 -13595
rect 470 -13629 528 -13595
rect 562 -13629 620 -13595
rect 654 -13629 712 -13595
rect 746 -13629 804 -13595
rect 838 -13629 896 -13595
rect 930 -13629 988 -13595
rect 1022 -13629 1080 -13595
rect 1114 -13629 1172 -13595
rect 1206 -13629 1264 -13595
rect 1298 -13629 1356 -13595
rect 1390 -13629 1448 -13595
rect 1482 -13629 1540 -13595
rect 1574 -13629 1632 -13595
rect 1666 -13629 1724 -13595
rect 1758 -13629 1816 -13595
rect 1850 -13629 1908 -13595
rect 1942 -13629 2000 -13595
rect 2034 -13629 2092 -13595
rect 2126 -13629 2184 -13595
rect 2218 -13629 2276 -13595
rect 2310 -13629 2368 -13595
rect 2402 -13629 2460 -13595
rect 2494 -13629 2552 -13595
rect 2586 -13629 2644 -13595
rect 2678 -13629 2736 -13595
rect 2770 -13629 2828 -13595
rect 2862 -13629 2920 -13595
rect 2954 -13629 3012 -13595
rect 3046 -13629 3104 -13595
rect 3138 -13629 3196 -13595
rect 3230 -13629 3288 -13595
rect 3322 -13629 3380 -13595
rect 3414 -13629 3472 -13595
rect 3506 -13629 3564 -13595
rect 3598 -13629 3656 -13595
rect 3690 -13629 3748 -13595
rect 3782 -13629 3840 -13595
rect 3874 -13629 3932 -13595
rect 3966 -13629 4024 -13595
rect 4058 -13629 4116 -13595
rect 4150 -13629 4208 -13595
rect 4242 -13629 4300 -13595
rect 4334 -13629 4392 -13595
rect 4426 -13629 4484 -13595
rect 4518 -13629 4576 -13595
rect 4610 -13629 4668 -13595
rect 4702 -13629 4760 -13595
rect 4794 -13629 4852 -13595
rect 4886 -13629 4944 -13595
rect 4978 -13629 5036 -13595
rect 5070 -13629 5128 -13595
rect 5162 -13629 5220 -13595
rect 5254 -13629 5312 -13595
rect 5346 -13629 5404 -13595
rect 5438 -13629 5496 -13595
rect 5530 -13629 5588 -13595
rect 5622 -13629 5680 -13595
rect 5714 -13629 5772 -13595
rect 5806 -13629 5864 -13595
rect 5898 -13629 5956 -13595
rect 5990 -13629 6048 -13595
rect 6082 -13629 6140 -13595
rect 6174 -13629 6232 -13595
rect 6266 -13629 6324 -13595
rect 6358 -13629 6416 -13595
rect 6450 -13629 6508 -13595
rect 6542 -13629 6600 -13595
rect 6634 -13629 6692 -13595
rect 6726 -13629 6784 -13595
rect 6818 -13629 6876 -13595
rect 6910 -13629 6968 -13595
rect 7002 -13629 7060 -13595
rect 7094 -13629 7152 -13595
rect 7186 -13629 7244 -13595
rect 7278 -13629 7336 -13595
rect 7370 -13629 7428 -13595
rect 7462 -13629 7520 -13595
rect 7554 -13629 7612 -13595
rect 7646 -13629 7704 -13595
rect 7738 -13629 7796 -13595
rect 7830 -13629 7888 -13595
rect 7922 -13629 7980 -13595
rect 8014 -13629 8072 -13595
rect 8106 -13629 8164 -13595
rect 8198 -13629 8256 -13595
rect 8290 -13629 8348 -13595
rect 8382 -13629 8440 -13595
rect 8474 -13629 8532 -13595
rect 8566 -13629 8624 -13595
rect 8658 -13629 8716 -13595
rect 8750 -13629 8808 -13595
rect 8842 -13629 8900 -13595
rect 8934 -13629 8992 -13595
rect 9026 -13629 9084 -13595
rect 9118 -13629 9176 -13595
rect 9210 -13629 9268 -13595
rect 9302 -13629 9360 -13595
rect 9394 -13629 9452 -13595
rect 9486 -13629 9544 -13595
rect 9578 -13629 9636 -13595
rect 9670 -13629 9728 -13595
rect 9762 -13629 9820 -13595
rect 9854 -13629 9912 -13595
rect 9946 -13629 10004 -13595
rect 10038 -13629 10096 -13595
rect 10130 -13629 10188 -13595
rect 10222 -13629 10280 -13595
rect 10314 -13629 10372 -13595
rect 10406 -13629 10464 -13595
rect 10498 -13629 10556 -13595
rect 10590 -13629 10648 -13595
rect 10682 -13629 10740 -13595
rect 10774 -13629 10832 -13595
rect 10866 -13629 10924 -13595
rect 10958 -13629 11016 -13595
rect 11050 -13629 11108 -13595
rect 11142 -13629 11200 -13595
rect 11234 -13629 11292 -13595
rect 11326 -13629 11384 -13595
rect 11418 -13629 11476 -13595
rect 11510 -13629 11568 -13595
rect 11602 -13629 11660 -13595
rect 11694 -13629 11752 -13595
rect 11786 -13629 11844 -13595
rect 11878 -13629 11936 -13595
rect 11970 -13629 12028 -13595
rect 12062 -13629 12120 -13595
rect 12154 -13629 12212 -13595
rect 12246 -13629 12304 -13595
rect 12338 -13629 12396 -13595
rect 12430 -13629 12488 -13595
rect 12522 -13629 12580 -13595
rect 12614 -13629 12672 -13595
rect 12706 -13629 12764 -13595
rect 12798 -13629 12856 -13595
rect 12890 -13629 12948 -13595
rect 12982 -13629 13040 -13595
rect 13074 -13629 13132 -13595
rect 13166 -13629 13224 -13595
rect 13258 -13629 13316 -13595
rect 13350 -13629 13408 -13595
rect 13442 -13629 13500 -13595
rect 13534 -13629 13592 -13595
rect 13626 -13629 13684 -13595
rect 13718 -13629 13776 -13595
rect 13810 -13629 13868 -13595
rect 13902 -13629 13960 -13595
rect 13994 -13629 14052 -13595
rect 14086 -13629 14144 -13595
rect 14178 -13629 14236 -13595
rect 14270 -13629 14328 -13595
rect 14362 -13629 14420 -13595
rect 14454 -13629 14512 -13595
rect 14546 -13629 14604 -13595
rect 14638 -13629 14696 -13595
rect 14730 -13629 14788 -13595
rect 14822 -13629 14880 -13595
rect 14914 -13629 14972 -13595
rect 15006 -13629 15064 -13595
rect 15098 -13629 15156 -13595
rect 15190 -13629 15248 -13595
rect 15282 -13629 15340 -13595
rect 15374 -13629 15432 -13595
rect 15466 -13629 15524 -13595
rect 15558 -13629 15616 -13595
rect 15650 -13629 15708 -13595
rect 15742 -13629 15800 -13595
rect 15834 -13629 15892 -13595
rect 15926 -13629 15984 -13595
rect 16018 -13629 16076 -13595
rect 16110 -13629 16168 -13595
rect 16202 -13629 16260 -13595
rect 16294 -13629 16352 -13595
rect 16386 -13629 16444 -13595
rect 16478 -13629 16536 -13595
rect 16570 -13629 16628 -13595
rect 16662 -13629 16946 -13595
rect -3193 -13660 16946 -13629
rect 1070 -13694 1116 -13690
rect -862 -13722 13 -13716
rect -862 -13756 -848 -13722
rect -814 -13756 -769 -13722
rect -735 -13756 13 -13722
rect -862 -13765 13 -13756
rect 1064 -13749 1122 -13694
rect 418 -13763 485 -13759
rect 1064 -13763 1076 -13749
rect -57 -13821 12 -13765
rect 418 -13783 1076 -13763
rect 1110 -13783 1122 -13749
rect 418 -13789 1122 -13783
rect -57 -13822 16 -13821
rect 94 -13822 152 -13821
rect 227 -13822 389 -13821
rect -954 -13879 -944 -13823
rect -886 -13879 -876 -13823
rect -778 -13829 -723 -13826
rect -57 -13827 389 -13822
rect -778 -13835 -718 -13829
rect -778 -13869 -764 -13835
rect -730 -13869 -718 -13835
rect -778 -13875 -718 -13869
rect -57 -13861 -30 -13827
rect 4 -13861 106 -13827
rect 140 -13861 242 -13827
rect 276 -13861 389 -13827
rect -57 -13870 389 -13861
rect 418 -13823 434 -13789
rect 468 -13791 1122 -13789
rect 468 -13823 982 -13791
rect 418 -13843 982 -13823
rect 1034 -13822 1122 -13791
rect 1034 -13843 1076 -13822
rect 418 -13856 1076 -13843
rect 1110 -13856 1122 -13822
rect -778 -13916 -723 -13875
rect -1834 -13971 -1824 -13916
rect -1769 -13971 -723 -13916
rect 308 -13956 387 -13870
rect 418 -13874 1122 -13856
rect 1153 -13822 1310 -13762
rect 1153 -13828 2449 -13822
rect 1153 -13862 1171 -13828
rect 1205 -13862 1263 -13828
rect 1297 -13833 2449 -13828
rect 1297 -13862 2369 -13833
rect 1153 -13867 2369 -13862
rect 2403 -13867 2449 -13833
rect 1153 -13884 2449 -13867
rect 2994 -13832 6963 -13815
rect 2994 -13866 3015 -13832
rect 3049 -13866 6876 -13832
rect 6910 -13866 6963 -13832
rect 1153 -13885 1310 -13884
rect 2994 -13886 6963 -13866
rect 7509 -13831 8255 -13813
rect 7509 -13832 8164 -13831
rect 7509 -13866 7522 -13832
rect 7556 -13865 8164 -13832
rect 8198 -13865 8255 -13831
rect 7556 -13866 8255 -13865
rect 7509 -13887 8255 -13866
rect 8799 -13833 9545 -13814
rect 8799 -13867 8811 -13833
rect 8845 -13867 9453 -13833
rect 9487 -13867 9545 -13833
rect 8799 -13885 9545 -13867
rect 10086 -13826 11058 -13820
rect 10086 -13832 11063 -13826
rect 10086 -13833 10925 -13832
rect 10086 -13834 10741 -13833
rect 10086 -13868 10099 -13834
rect 10133 -13867 10741 -13834
rect 10775 -13867 10832 -13833
rect 10866 -13866 10925 -13833
rect 10959 -13866 11017 -13832
rect 11051 -13866 11063 -13832
rect 11233 -13835 11418 -13827
rect 10866 -13867 11063 -13866
rect 10133 -13868 11063 -13867
rect 10086 -13872 11063 -13868
rect 10086 -13890 11058 -13872
rect 11110 -13909 11120 -13857
rect 11172 -13909 11182 -13857
rect 11233 -13869 11250 -13835
rect 11284 -13869 11344 -13835
rect 11378 -13869 11418 -13835
rect 11233 -13956 11418 -13869
rect 308 -13992 11419 -13956
rect -3193 -14139 16946 -14108
rect -3193 -14173 -2968 -14139
rect -2934 -14173 -2876 -14139
rect -2842 -14173 -2784 -14139
rect -2750 -14173 -2692 -14139
rect -2658 -14173 -2600 -14139
rect -2566 -14173 -2508 -14139
rect -2474 -14173 -2416 -14139
rect -2382 -14173 -2324 -14139
rect -2290 -14173 -2232 -14139
rect -2198 -14173 -2140 -14139
rect -2106 -14173 -2048 -14139
rect -2014 -14173 -1956 -14139
rect -1922 -14173 -1864 -14139
rect -1830 -14173 -1772 -14139
rect -1738 -14173 -1680 -14139
rect -1646 -14173 -1588 -14139
rect -1554 -14173 -1496 -14139
rect -1462 -14173 -1404 -14139
rect -1370 -14173 -1312 -14139
rect -1278 -14173 -1220 -14139
rect -1186 -14173 -1128 -14139
rect -1094 -14173 -1036 -14139
rect -1002 -14173 -944 -14139
rect -910 -14173 -852 -14139
rect -818 -14173 -760 -14139
rect -726 -14173 -668 -14139
rect -634 -14173 -576 -14139
rect -542 -14173 -484 -14139
rect -450 -14173 -392 -14139
rect -358 -14173 -300 -14139
rect -266 -14173 -208 -14139
rect -174 -14173 -116 -14139
rect -82 -14173 -24 -14139
rect 10 -14173 68 -14139
rect 102 -14173 160 -14139
rect 194 -14173 252 -14139
rect 286 -14173 344 -14139
rect 378 -14173 436 -14139
rect 470 -14173 528 -14139
rect 562 -14173 620 -14139
rect 654 -14173 712 -14139
rect 746 -14173 804 -14139
rect 838 -14173 896 -14139
rect 930 -14173 988 -14139
rect 1022 -14173 1080 -14139
rect 1114 -14173 1172 -14139
rect 1206 -14173 1264 -14139
rect 1298 -14173 1356 -14139
rect 1390 -14173 1448 -14139
rect 1482 -14173 1540 -14139
rect 1574 -14173 1632 -14139
rect 1666 -14173 1724 -14139
rect 1758 -14173 1816 -14139
rect 1850 -14173 1908 -14139
rect 1942 -14173 2000 -14139
rect 2034 -14173 2092 -14139
rect 2126 -14173 2184 -14139
rect 2218 -14173 2276 -14139
rect 2310 -14173 2368 -14139
rect 2402 -14173 2460 -14139
rect 2494 -14173 2552 -14139
rect 2586 -14173 2644 -14139
rect 2678 -14173 2736 -14139
rect 2770 -14173 2828 -14139
rect 2862 -14173 2920 -14139
rect 2954 -14173 3012 -14139
rect 3046 -14173 3104 -14139
rect 3138 -14173 3196 -14139
rect 3230 -14173 3288 -14139
rect 3322 -14173 3380 -14139
rect 3414 -14173 3472 -14139
rect 3506 -14173 3564 -14139
rect 3598 -14173 3656 -14139
rect 3690 -14173 3748 -14139
rect 3782 -14173 3840 -14139
rect 3874 -14173 3932 -14139
rect 3966 -14173 4024 -14139
rect 4058 -14173 4116 -14139
rect 4150 -14173 4208 -14139
rect 4242 -14173 4300 -14139
rect 4334 -14173 4392 -14139
rect 4426 -14173 4484 -14139
rect 4518 -14173 4576 -14139
rect 4610 -14173 4668 -14139
rect 4702 -14173 4760 -14139
rect 4794 -14173 4852 -14139
rect 4886 -14173 4944 -14139
rect 4978 -14173 5036 -14139
rect 5070 -14173 5128 -14139
rect 5162 -14173 5220 -14139
rect 5254 -14173 5312 -14139
rect 5346 -14173 5404 -14139
rect 5438 -14173 5496 -14139
rect 5530 -14173 5588 -14139
rect 5622 -14173 5680 -14139
rect 5714 -14173 5772 -14139
rect 5806 -14173 5864 -14139
rect 5898 -14173 5956 -14139
rect 5990 -14173 6048 -14139
rect 6082 -14173 6140 -14139
rect 6174 -14173 6232 -14139
rect 6266 -14173 6324 -14139
rect 6358 -14173 6416 -14139
rect 6450 -14173 6508 -14139
rect 6542 -14173 6600 -14139
rect 6634 -14173 6692 -14139
rect 6726 -14173 6784 -14139
rect 6818 -14173 6876 -14139
rect 6910 -14173 6968 -14139
rect 7002 -14173 7060 -14139
rect 7094 -14173 7152 -14139
rect 7186 -14173 7244 -14139
rect 7278 -14173 7336 -14139
rect 7370 -14173 7428 -14139
rect 7462 -14173 7520 -14139
rect 7554 -14173 7612 -14139
rect 7646 -14173 7704 -14139
rect 7738 -14173 7796 -14139
rect 7830 -14173 7888 -14139
rect 7922 -14173 7980 -14139
rect 8014 -14173 8072 -14139
rect 8106 -14173 8164 -14139
rect 8198 -14173 8256 -14139
rect 8290 -14173 8348 -14139
rect 8382 -14173 8440 -14139
rect 8474 -14173 8532 -14139
rect 8566 -14173 8624 -14139
rect 8658 -14173 8716 -14139
rect 8750 -14173 8808 -14139
rect 8842 -14173 8900 -14139
rect 8934 -14173 8992 -14139
rect 9026 -14173 9084 -14139
rect 9118 -14173 9176 -14139
rect 9210 -14173 9268 -14139
rect 9302 -14173 9360 -14139
rect 9394 -14173 9452 -14139
rect 9486 -14173 9544 -14139
rect 9578 -14173 9636 -14139
rect 9670 -14173 9728 -14139
rect 9762 -14173 9820 -14139
rect 9854 -14173 9912 -14139
rect 9946 -14173 10004 -14139
rect 10038 -14173 10096 -14139
rect 10130 -14173 10188 -14139
rect 10222 -14173 10280 -14139
rect 10314 -14173 10372 -14139
rect 10406 -14173 10464 -14139
rect 10498 -14173 10556 -14139
rect 10590 -14173 10648 -14139
rect 10682 -14173 10740 -14139
rect 10774 -14173 10832 -14139
rect 10866 -14173 10924 -14139
rect 10958 -14173 11016 -14139
rect 11050 -14173 11108 -14139
rect 11142 -14173 11200 -14139
rect 11234 -14173 11292 -14139
rect 11326 -14173 11384 -14139
rect 11418 -14173 11476 -14139
rect 11510 -14173 11568 -14139
rect 11602 -14173 11660 -14139
rect 11694 -14173 11752 -14139
rect 11786 -14173 11844 -14139
rect 11878 -14173 11936 -14139
rect 11970 -14173 12028 -14139
rect 12062 -14173 12120 -14139
rect 12154 -14173 12212 -14139
rect 12246 -14173 12304 -14139
rect 12338 -14173 12396 -14139
rect 12430 -14173 12488 -14139
rect 12522 -14173 12580 -14139
rect 12614 -14173 12672 -14139
rect 12706 -14173 12764 -14139
rect 12798 -14173 12856 -14139
rect 12890 -14173 12948 -14139
rect 12982 -14173 13040 -14139
rect 13074 -14173 13132 -14139
rect 13166 -14173 13224 -14139
rect 13258 -14173 13316 -14139
rect 13350 -14173 13408 -14139
rect 13442 -14173 13500 -14139
rect 13534 -14173 13592 -14139
rect 13626 -14173 13684 -14139
rect 13718 -14173 13776 -14139
rect 13810 -14173 13868 -14139
rect 13902 -14173 13960 -14139
rect 13994 -14173 14052 -14139
rect 14086 -14173 14144 -14139
rect 14178 -14173 14236 -14139
rect 14270 -14173 14328 -14139
rect 14362 -14173 14420 -14139
rect 14454 -14173 14512 -14139
rect 14546 -14173 14604 -14139
rect 14638 -14173 14696 -14139
rect 14730 -14173 14788 -14139
rect 14822 -14173 14880 -14139
rect 14914 -14173 14972 -14139
rect 15006 -14173 15064 -14139
rect 15098 -14173 15156 -14139
rect 15190 -14173 15248 -14139
rect 15282 -14173 15340 -14139
rect 15374 -14173 15432 -14139
rect 15466 -14173 15524 -14139
rect 15558 -14173 15616 -14139
rect 15650 -14173 15708 -14139
rect 15742 -14173 15800 -14139
rect 15834 -14173 15892 -14139
rect 15926 -14173 15984 -14139
rect 16018 -14173 16076 -14139
rect 16110 -14173 16168 -14139
rect 16202 -14173 16260 -14139
rect 16294 -14173 16352 -14139
rect 16386 -14173 16444 -14139
rect 16478 -14173 16536 -14139
rect 16570 -14173 16628 -14139
rect 16662 -14173 16946 -14139
rect -3193 -14204 16946 -14173
<< via1 >>
rect -1792 -343 -1740 -291
rect -771 -301 -719 -290
rect -771 -335 -762 -301
rect -762 -335 -728 -301
rect -728 -335 -719 -301
rect -771 -342 -719 -335
rect 982 -377 1034 -325
rect 11120 -268 11172 -259
rect 11120 -302 11129 -268
rect 11129 -302 11163 -268
rect 11163 -302 11172 -268
rect 11120 -311 11172 -302
rect 982 -733 1034 -681
rect 12753 -734 12805 -682
rect 423 -812 475 -802
rect 423 -846 433 -812
rect 433 -846 467 -812
rect 467 -846 475 -812
rect 423 -854 475 -846
rect 12463 -887 12522 -828
rect 7165 -1287 7217 -1235
rect 11118 -1284 11170 -1232
rect 423 -1392 475 -1383
rect 423 -1426 432 -1392
rect 432 -1426 466 -1392
rect 466 -1426 475 -1392
rect 423 -1435 475 -1426
rect 11378 -1355 11430 -1345
rect 11378 -1389 11387 -1355
rect 11387 -1389 11421 -1355
rect 11421 -1389 11430 -1355
rect 11378 -1397 11430 -1389
rect 12752 -1392 12804 -1382
rect 12752 -1426 12773 -1392
rect 12773 -1426 12804 -1392
rect 12752 -1434 12804 -1426
rect 7163 -1815 7215 -1763
rect 12756 -1818 12808 -1766
rect -942 -1943 -890 -1891
rect -217 -1865 -165 -1854
rect -217 -1899 -210 -1865
rect -210 -1899 -176 -1865
rect -176 -1899 -165 -1865
rect -217 -1906 -165 -1899
rect 423 -1900 475 -1890
rect 423 -1934 432 -1900
rect 432 -1934 466 -1900
rect 466 -1934 475 -1900
rect 423 -1942 475 -1934
rect 11375 -1863 11427 -1856
rect 11375 -1897 11386 -1863
rect 11386 -1897 11420 -1863
rect 11420 -1897 11427 -1863
rect 11375 -1908 11427 -1897
rect 428 -2480 480 -2469
rect 428 -2514 436 -2480
rect 436 -2514 470 -2480
rect 470 -2514 480 -2480
rect 428 -2521 480 -2514
rect 11378 -2445 11430 -2436
rect 11378 -2479 11386 -2445
rect 11386 -2479 11420 -2445
rect 11420 -2479 11430 -2445
rect 11378 -2488 11430 -2479
rect 12466 -2441 12480 -2414
rect 12480 -2441 12514 -2414
rect 12514 -2441 12518 -2414
rect 12466 -2466 12518 -2441
rect 12755 -2479 12807 -2472
rect 12755 -2513 12765 -2479
rect 12765 -2513 12799 -2479
rect 12799 -2513 12807 -2479
rect 12755 -2524 12807 -2513
rect 13926 -2485 13978 -2433
rect 12466 -2553 12518 -2528
rect 12466 -2580 12480 -2553
rect 12480 -2580 12514 -2553
rect 12514 -2580 12518 -2553
rect -1968 -2952 -1916 -2944
rect -1968 -2986 -1960 -2952
rect -1960 -2986 -1926 -2952
rect -1926 -2986 -1916 -2952
rect -1968 -2996 -1916 -2986
rect -1792 -2915 -1740 -2906
rect -1792 -2949 -1783 -2915
rect -1783 -2949 -1749 -2915
rect -1749 -2949 -1740 -2915
rect -1792 -2958 -1740 -2949
rect -221 -3033 -169 -2981
rect 11376 -2952 11428 -2943
rect 11376 -2986 11384 -2952
rect 11384 -2986 11418 -2952
rect 11418 -2986 11428 -2952
rect 11376 -2995 11428 -2986
rect -1968 -3114 -1916 -3062
rect -1272 -3118 -1213 -3059
rect 115 -3573 167 -3521
rect 11373 -3567 11425 -3557
rect 11373 -3601 11383 -3567
rect 11383 -3601 11417 -3567
rect 11417 -3601 11425 -3567
rect 11373 -3609 11425 -3601
rect 12466 -3999 12480 -3972
rect 12480 -3999 12514 -3972
rect 12514 -3999 12518 -3972
rect 12466 -4024 12518 -3999
rect 427 -4040 479 -4031
rect 427 -4074 436 -4040
rect 436 -4074 470 -4040
rect 470 -4074 479 -4040
rect 427 -4083 479 -4074
rect 11377 -4077 11429 -4067
rect 11377 -4111 11386 -4077
rect 11386 -4111 11420 -4077
rect 11420 -4111 11429 -4077
rect 11377 -4119 11429 -4111
rect 12755 -4039 12807 -4028
rect 12755 -4073 12765 -4039
rect 12765 -4073 12799 -4039
rect 12799 -4073 12807 -4039
rect 12755 -4080 12807 -4073
rect 12466 -4111 12518 -4086
rect 12466 -4138 12480 -4111
rect 12480 -4138 12514 -4111
rect 12514 -4138 12518 -4111
rect 14628 -4118 14682 -4064
rect -771 -4663 -716 -4608
rect 115 -4695 167 -4643
rect 424 -4619 476 -4610
rect 424 -4653 433 -4619
rect 433 -4653 467 -4619
rect 467 -4653 476 -4619
rect 424 -4662 476 -4653
rect 11375 -4657 11427 -4645
rect 11375 -4691 11384 -4657
rect 11384 -4691 11418 -4657
rect 11418 -4691 11427 -4657
rect 11375 -4697 11427 -4691
rect 7163 -4789 7215 -4737
rect 12756 -4786 12808 -4734
rect 427 -5128 479 -5120
rect 427 -5162 436 -5128
rect 436 -5162 470 -5128
rect 470 -5162 479 -5128
rect 427 -5172 479 -5162
rect 12752 -5126 12804 -5118
rect 11380 -5162 11432 -5152
rect 11380 -5196 11389 -5162
rect 11389 -5196 11423 -5162
rect 11423 -5196 11432 -5162
rect 11380 -5204 11432 -5196
rect 12752 -5160 12773 -5126
rect 12773 -5160 12804 -5126
rect 12752 -5170 12804 -5160
rect 7165 -5317 7217 -5265
rect 11118 -5320 11170 -5268
rect 422 -5708 474 -5699
rect 422 -5742 432 -5708
rect 432 -5742 466 -5708
rect 466 -5742 474 -5708
rect 422 -5751 474 -5742
rect 12463 -5724 12522 -5665
rect 982 -5871 1034 -5819
rect 12753 -5870 12805 -5818
rect -944 -6218 -886 -6207
rect -944 -6252 -932 -6218
rect -932 -6252 -898 -6218
rect -898 -6252 -886 -6218
rect -944 -6263 -886 -6252
rect -772 -6217 -714 -6207
rect -772 -6251 -760 -6217
rect -760 -6251 -726 -6217
rect -726 -6251 -714 -6217
rect -772 -6263 -714 -6251
rect 982 -6227 1034 -6175
rect 11120 -6250 11172 -6241
rect 11120 -6284 11129 -6250
rect 11129 -6284 11163 -6250
rect 11163 -6284 11172 -6250
rect 11120 -6293 11172 -6284
rect 14627 -6274 14682 -6219
rect 15834 -6274 15889 -6219
rect -1271 -6409 -1213 -6353
rect -768 -6409 -715 -6356
rect -772 -6727 -714 -6671
rect 7349 -6726 7407 -6670
rect -2607 -6830 -2554 -6821
rect -2607 -6864 -2599 -6830
rect -2599 -6864 -2565 -6830
rect -2565 -6864 -2554 -6830
rect -2607 -6873 -2554 -6864
rect 5028 -6840 5082 -6786
rect 13925 -6840 13979 -6786
rect -1968 -7003 -1915 -6951
rect -405 -6958 -346 -6899
rect 3736 -6958 3795 -6899
rect 4945 -6977 4999 -6923
rect 15832 -6977 15886 -6923
rect 4945 -7204 4999 -7195
rect 4945 -7238 4955 -7204
rect 4955 -7238 4989 -7204
rect 4989 -7238 4999 -7204
rect 4945 -7249 4999 -7238
rect 2736 -7317 2795 -7258
rect 3736 -7304 3795 -7292
rect 3736 -7338 3747 -7304
rect 3747 -7338 3781 -7304
rect 3781 -7338 3795 -7304
rect 3736 -7351 3795 -7338
rect 5028 -7306 5082 -7299
rect 5028 -7340 5036 -7306
rect 5036 -7340 5070 -7306
rect 5070 -7340 5082 -7306
rect 5028 -7353 5082 -7340
rect 7349 -7264 7407 -7254
rect 7349 -7298 7356 -7264
rect 7356 -7298 7390 -7264
rect 7390 -7298 7407 -7264
rect 7349 -7310 7407 -7298
rect 15971 -7326 16030 -7267
rect -620 -7498 -561 -7439
rect 2736 -7498 2795 -7439
rect -1968 -7960 -1915 -7908
rect -619 -7961 -560 -7902
rect 982 -7993 1034 -7941
rect 11120 -7884 11172 -7875
rect 11120 -7918 11129 -7884
rect 11129 -7918 11163 -7884
rect 11163 -7918 11172 -7884
rect 11120 -7927 11172 -7918
rect 982 -8349 1034 -8297
rect 12753 -8350 12805 -8298
rect 423 -8428 475 -8418
rect 423 -8462 433 -8428
rect 433 -8462 467 -8428
rect 467 -8462 475 -8428
rect 423 -8470 475 -8462
rect 12463 -8503 12522 -8444
rect 15972 -8475 16031 -8416
rect 7165 -8903 7217 -8851
rect 11118 -8900 11170 -8848
rect 423 -9008 475 -8999
rect 423 -9042 432 -9008
rect 432 -9042 466 -9008
rect 466 -9042 475 -9008
rect 423 -9051 475 -9042
rect 11378 -8971 11430 -8961
rect 11378 -9005 11387 -8971
rect 11387 -9005 11421 -8971
rect 11421 -9005 11430 -8971
rect 11378 -9013 11430 -9005
rect 12752 -9008 12804 -8998
rect 12752 -9042 12773 -9008
rect 12773 -9042 12804 -9008
rect 12752 -9050 12804 -9042
rect 7163 -9431 7215 -9379
rect 12756 -9434 12808 -9382
rect -942 -9559 -890 -9507
rect -217 -9481 -165 -9470
rect -217 -9515 -210 -9481
rect -210 -9515 -176 -9481
rect -176 -9515 -165 -9481
rect -217 -9522 -165 -9515
rect 423 -9516 475 -9506
rect 423 -9550 432 -9516
rect 432 -9550 466 -9516
rect 466 -9550 475 -9516
rect 423 -9558 475 -9550
rect 11375 -9479 11427 -9472
rect 11375 -9513 11386 -9479
rect 11386 -9513 11420 -9479
rect 11420 -9513 11427 -9479
rect 11375 -9524 11427 -9513
rect 428 -10096 480 -10085
rect 428 -10130 436 -10096
rect 436 -10130 470 -10096
rect 470 -10130 480 -10096
rect 428 -10137 480 -10130
rect 11378 -10061 11430 -10052
rect 11378 -10095 11386 -10061
rect 11386 -10095 11420 -10061
rect 11420 -10095 11430 -10061
rect 11378 -10104 11430 -10095
rect 12466 -10057 12480 -10030
rect 12480 -10057 12514 -10030
rect 12514 -10057 12518 -10030
rect 12466 -10082 12518 -10057
rect 12755 -10095 12807 -10088
rect 12755 -10129 12765 -10095
rect 12765 -10129 12799 -10095
rect 12799 -10129 12807 -10095
rect 12755 -10140 12807 -10129
rect 12466 -10169 12518 -10144
rect 12466 -10196 12480 -10169
rect 12480 -10196 12514 -10169
rect 12514 -10196 12518 -10169
rect -2607 -10543 -2554 -10490
rect -1969 -10499 -1915 -10489
rect -1969 -10533 -1961 -10499
rect -1961 -10533 -1927 -10499
rect -1927 -10533 -1915 -10499
rect -1969 -10543 -1915 -10533
rect -1823 -10534 -1769 -10525
rect -1823 -10568 -1813 -10534
rect -1813 -10568 -1779 -10534
rect -1779 -10568 -1769 -10534
rect -1823 -10579 -1769 -10568
rect -221 -10649 -169 -10597
rect 11376 -10568 11428 -10559
rect 11376 -10602 11384 -10568
rect 11384 -10602 11418 -10568
rect 11418 -10602 11428 -10568
rect 11376 -10611 11428 -10602
rect 115 -11189 167 -11137
rect 11373 -11183 11425 -11173
rect 11373 -11217 11383 -11183
rect 11383 -11217 11417 -11183
rect 11417 -11217 11425 -11183
rect 11373 -11225 11425 -11217
rect 12466 -11615 12480 -11588
rect 12480 -11615 12514 -11588
rect 12514 -11615 12518 -11588
rect 12466 -11640 12518 -11615
rect 427 -11656 479 -11647
rect 427 -11690 436 -11656
rect 436 -11690 470 -11656
rect 470 -11690 479 -11656
rect 427 -11699 479 -11690
rect 11377 -11693 11429 -11683
rect 11377 -11727 11386 -11693
rect 11386 -11727 11420 -11693
rect 11420 -11727 11429 -11693
rect 11377 -11735 11429 -11727
rect 12755 -11655 12807 -11644
rect 12755 -11689 12765 -11655
rect 12765 -11689 12799 -11655
rect 12799 -11689 12807 -11655
rect 12755 -11696 12807 -11689
rect 12466 -11727 12518 -11702
rect 12466 -11754 12480 -11727
rect 12480 -11754 12514 -11727
rect 12514 -11754 12518 -11727
rect -404 -12282 -346 -12224
rect 115 -12311 167 -12259
rect 424 -12235 476 -12226
rect 424 -12269 433 -12235
rect 433 -12269 467 -12235
rect 467 -12269 476 -12235
rect 424 -12278 476 -12269
rect 11375 -12273 11427 -12261
rect 11375 -12307 11384 -12273
rect 11384 -12307 11418 -12273
rect 11418 -12307 11427 -12273
rect 11375 -12313 11427 -12307
rect 7163 -12405 7215 -12353
rect 12756 -12402 12808 -12350
rect 427 -12744 479 -12736
rect 427 -12778 436 -12744
rect 436 -12778 470 -12744
rect 470 -12778 479 -12744
rect 427 -12788 479 -12778
rect 12752 -12742 12804 -12734
rect 11380 -12778 11432 -12768
rect 11380 -12812 11389 -12778
rect 11389 -12812 11423 -12778
rect 11423 -12812 11432 -12778
rect 11380 -12820 11432 -12812
rect 12752 -12776 12773 -12742
rect 12773 -12776 12804 -12742
rect 12752 -12786 12804 -12776
rect 7165 -12933 7217 -12881
rect 11118 -12936 11170 -12884
rect 422 -13324 474 -13315
rect 422 -13358 432 -13324
rect 432 -13358 466 -13324
rect 466 -13358 474 -13324
rect 422 -13367 474 -13358
rect 12463 -13340 12522 -13281
rect 982 -13487 1034 -13435
rect 12753 -13486 12805 -13434
rect -944 -13834 -886 -13823
rect -944 -13868 -932 -13834
rect -932 -13868 -898 -13834
rect -898 -13868 -886 -13834
rect -944 -13879 -886 -13868
rect 982 -13843 1034 -13791
rect -1824 -13971 -1769 -13916
rect 11120 -13866 11172 -13857
rect 11120 -13900 11129 -13866
rect 11129 -13900 11163 -13866
rect 11163 -13900 11172 -13866
rect 11120 -13909 11172 -13900
<< metal2 >>
rect 11110 -259 11178 -243
rect -1792 -291 -1740 -280
rect -1792 -2906 -1740 -343
rect -771 -290 -716 -279
rect -719 -342 -716 -290
rect 11110 -311 11120 -259
rect 11172 -311 11178 -259
rect -1968 -2944 -1915 -2933
rect -1916 -2996 -1915 -2944
rect -1792 -2988 -1740 -2958
rect -944 -1891 -886 -1879
rect -944 -1943 -942 -1891
rect -890 -1943 -886 -1891
rect -1968 -3062 -1915 -2996
rect -1916 -3114 -1915 -3062
rect -2607 -6821 -2554 -6811
rect -2607 -10490 -2554 -6873
rect -1968 -6951 -1915 -3114
rect -1272 -3059 -1213 -3049
rect -1272 -6353 -1213 -3118
rect -944 -6207 -886 -1943
rect -771 -4608 -716 -342
rect 979 -325 1039 -314
rect 979 -377 982 -325
rect 1034 -377 1039 -325
rect 979 -681 1039 -377
rect 979 -733 982 -681
rect 1034 -733 1039 -681
rect 979 -743 1039 -733
rect 423 -802 475 -792
rect 423 -1383 475 -854
rect 423 -1445 475 -1435
rect 7154 -1235 7223 -1225
rect 7154 -1287 7165 -1235
rect 7217 -1287 7223 -1235
rect 7154 -1763 7223 -1287
rect 11110 -1232 11178 -311
rect 12751 -682 12806 -671
rect 12751 -734 12753 -682
rect 12805 -734 12806 -682
rect 11110 -1284 11118 -1232
rect 11170 -1284 11178 -1232
rect 11110 -1294 11178 -1284
rect 12463 -828 12522 -818
rect 7154 -1815 7163 -1763
rect 7215 -1815 7223 -1763
rect 7154 -1821 7223 -1815
rect 11372 -1345 11434 -1332
rect 11372 -1397 11378 -1345
rect 11430 -1397 11434 -1345
rect 7163 -1825 7215 -1821
rect -217 -1854 -165 -1844
rect -227 -1906 -217 -1860
rect 11372 -1856 11434 -1397
rect -165 -1906 -164 -1860
rect 427 -1880 476 -1879
rect -227 -2981 -164 -1906
rect 423 -1890 476 -1880
rect 475 -1942 476 -1890
rect 11372 -1908 11375 -1856
rect 11427 -1908 11434 -1856
rect 11372 -1921 11434 -1908
rect 423 -1952 476 -1942
rect 427 -2459 476 -1952
rect 12463 -2414 12522 -887
rect 12751 -1382 12806 -734
rect 12751 -1434 12752 -1382
rect 12804 -1434 12806 -1382
rect 12751 -1435 12806 -1434
rect 12752 -1444 12804 -1435
rect 11374 -2436 11433 -2423
rect 427 -2469 480 -2459
rect 427 -2521 428 -2469
rect 427 -2531 480 -2521
rect 11374 -2488 11378 -2436
rect 11430 -2488 11433 -2436
rect 427 -2533 476 -2531
rect -227 -3033 -221 -2981
rect -169 -3033 -164 -2981
rect 11374 -2943 11433 -2488
rect 12463 -2466 12466 -2414
rect 12518 -2466 12522 -2414
rect 12463 -2528 12522 -2466
rect 12463 -2580 12466 -2528
rect 12518 -2580 12522 -2528
rect 12753 -1766 12812 -1753
rect 12753 -1818 12756 -1766
rect 12808 -1818 12812 -1766
rect 12753 -2472 12812 -1818
rect 12753 -2524 12755 -2472
rect 12807 -2524 12812 -2472
rect 12753 -2538 12812 -2524
rect 13925 -2433 13979 -2422
rect 13925 -2485 13926 -2433
rect 13978 -2485 13979 -2433
rect 12463 -2593 12522 -2580
rect 11374 -2995 11376 -2943
rect 11428 -2995 11433 -2943
rect 11374 -3008 11433 -2995
rect -227 -3048 -164 -3033
rect -771 -4673 -716 -4663
rect 113 -3521 170 -3507
rect 113 -3573 115 -3521
rect 167 -3573 170 -3521
rect 11375 -3547 11426 -3545
rect 113 -4643 170 -3573
rect 11373 -3557 11426 -3547
rect 11425 -3609 11426 -3557
rect 11373 -3619 11426 -3609
rect 425 -4031 480 -4018
rect 425 -4083 427 -4031
rect 479 -4083 480 -4031
rect 425 -4600 480 -4083
rect 11375 -4057 11426 -3619
rect 12463 -3972 12522 -3959
rect 12463 -4024 12466 -3972
rect 12518 -4024 12522 -3972
rect 11375 -4067 11429 -4057
rect 11375 -4119 11377 -4067
rect 11375 -4129 11429 -4119
rect 12463 -4086 12522 -4024
rect 11375 -4132 11426 -4129
rect 113 -4695 115 -4643
rect 167 -4695 170 -4643
rect 424 -4610 480 -4600
rect 476 -4662 480 -4610
rect 12463 -4138 12466 -4086
rect 12518 -4138 12522 -4086
rect 424 -4672 480 -4662
rect 425 -4675 480 -4672
rect 11373 -4645 11435 -4633
rect 113 -4701 170 -4695
rect 11373 -4697 11375 -4645
rect 11427 -4697 11435 -4645
rect 115 -4705 167 -4701
rect 7163 -4731 7215 -4727
rect 7154 -4737 7223 -4731
rect 7154 -4789 7163 -4737
rect 7215 -4789 7223 -4737
rect 424 -5110 476 -5107
rect 424 -5120 479 -5110
rect 424 -5172 427 -5120
rect 424 -5182 479 -5172
rect 424 -5689 476 -5182
rect 7154 -5265 7223 -4789
rect 11373 -5152 11435 -4697
rect 11373 -5204 11380 -5152
rect 11432 -5204 11435 -5152
rect 11373 -5217 11435 -5204
rect 7154 -5317 7165 -5265
rect 7217 -5317 7223 -5265
rect 7154 -5327 7223 -5317
rect 11110 -5268 11178 -5258
rect 11110 -5320 11118 -5268
rect 11170 -5320 11178 -5268
rect 422 -5699 476 -5689
rect 474 -5751 476 -5699
rect 422 -5761 476 -5751
rect 424 -5764 476 -5761
rect 979 -5819 1039 -5809
rect 979 -5871 982 -5819
rect 1034 -5871 1039 -5819
rect 979 -6175 1039 -5871
rect -944 -6273 -886 -6263
rect -773 -6207 -712 -6194
rect -773 -6263 -772 -6207
rect -714 -6263 -712 -6207
rect 979 -6227 982 -6175
rect 1034 -6227 1039 -6175
rect 979 -6238 1039 -6227
rect -1272 -6409 -1271 -6353
rect -1272 -6420 -1213 -6409
rect -773 -6356 -712 -6263
rect 11110 -6241 11178 -5320
rect 12463 -5665 12522 -4138
rect 12753 -4028 12812 -4014
rect 12753 -4080 12755 -4028
rect 12807 -4080 12812 -4028
rect 12753 -4734 12812 -4080
rect 12753 -4786 12756 -4734
rect 12808 -4786 12812 -4734
rect 12753 -4799 12812 -4786
rect 12752 -5117 12804 -5108
rect 12463 -5734 12522 -5724
rect 12751 -5118 12806 -5117
rect 12751 -5170 12752 -5118
rect 12804 -5170 12806 -5118
rect 12751 -5818 12806 -5170
rect 12751 -5870 12753 -5818
rect 12805 -5870 12806 -5818
rect 12751 -5881 12806 -5870
rect 11110 -6293 11120 -6241
rect 11172 -6293 11178 -6241
rect 11110 -6309 11178 -6293
rect -773 -6409 -768 -6356
rect -715 -6409 -712 -6356
rect -773 -6671 -712 -6409
rect -773 -6709 -772 -6671
rect -714 -6709 -712 -6671
rect 7345 -6670 7409 -6658
rect -772 -6737 -714 -6727
rect 7345 -6726 7349 -6670
rect 7407 -6726 7409 -6670
rect 5028 -6786 5082 -6776
rect -1968 -7010 -1915 -7003
rect -405 -6899 -346 -6889
rect -620 -7439 -561 -7429
rect -561 -7498 -559 -7460
rect -2607 -10553 -2554 -10543
rect -1969 -7908 -1915 -7898
rect -1969 -7960 -1968 -7908
rect -1969 -10489 -1915 -7960
rect -620 -7902 -559 -7498
rect -620 -7961 -619 -7902
rect -560 -7961 -559 -7902
rect -620 -7973 -559 -7961
rect -944 -9507 -886 -9495
rect -944 -9559 -942 -9507
rect -890 -9559 -886 -9507
rect -1969 -10556 -1915 -10543
rect -1824 -10525 -1769 -10514
rect -1824 -10579 -1823 -10525
rect -1824 -13916 -1769 -10579
rect -944 -13823 -886 -9559
rect -405 -12224 -346 -6958
rect 3736 -6899 3795 -6889
rect 2736 -7255 2795 -7248
rect 2735 -7258 2796 -7255
rect 2735 -7317 2736 -7258
rect 2795 -7317 2796 -7258
rect 2735 -7439 2796 -7317
rect 3736 -7292 3795 -6958
rect 4945 -6923 4999 -6905
rect 4945 -7195 4999 -6977
rect 4945 -7259 4999 -7249
rect 3736 -7361 3795 -7351
rect 5028 -7299 5082 -6840
rect 7345 -7254 7409 -6726
rect 13925 -6786 13979 -2485
rect 14627 -4064 14682 -4053
rect 14627 -4118 14628 -4064
rect 14627 -6219 14682 -4118
rect 14627 -6284 14682 -6274
rect 15829 -6219 15892 -6206
rect 15829 -6274 15834 -6219
rect 15889 -6274 15892 -6219
rect 13925 -6850 13979 -6840
rect 15829 -6923 15892 -6274
rect 15829 -6977 15832 -6923
rect 15886 -6977 15892 -6923
rect 15829 -6991 15892 -6977
rect 7345 -7310 7349 -7254
rect 7407 -7310 7409 -7254
rect 15971 -7262 16030 -7257
rect 7345 -7339 7409 -7310
rect 15968 -7267 16033 -7262
rect 15968 -7326 15971 -7267
rect 16030 -7326 16033 -7267
rect 5028 -7363 5082 -7353
rect 2735 -7498 2736 -7439
rect 2795 -7498 2796 -7439
rect 2735 -7508 2796 -7498
rect 11110 -7875 11178 -7859
rect 11110 -7927 11120 -7875
rect 11172 -7927 11178 -7875
rect 979 -7941 1039 -7930
rect 979 -7993 982 -7941
rect 1034 -7993 1039 -7941
rect 979 -8297 1039 -7993
rect 979 -8349 982 -8297
rect 1034 -8349 1039 -8297
rect 979 -8359 1039 -8349
rect 423 -8418 475 -8408
rect 423 -8999 475 -8470
rect 423 -9061 475 -9051
rect 7154 -8851 7223 -8841
rect 7154 -8903 7165 -8851
rect 7217 -8903 7223 -8851
rect 7154 -9379 7223 -8903
rect 11110 -8848 11178 -7927
rect 12751 -8298 12806 -8287
rect 12751 -8350 12753 -8298
rect 12805 -8350 12806 -8298
rect 11110 -8900 11118 -8848
rect 11170 -8900 11178 -8848
rect 11110 -8910 11178 -8900
rect 12463 -8444 12522 -8434
rect 7154 -9431 7163 -9379
rect 7215 -9431 7223 -9379
rect 7154 -9437 7223 -9431
rect 11372 -8961 11434 -8948
rect 11372 -9013 11378 -8961
rect 11430 -9013 11434 -8961
rect 7163 -9441 7215 -9437
rect -217 -9470 -165 -9460
rect -227 -9522 -217 -9476
rect 11372 -9472 11434 -9013
rect -165 -9522 -164 -9476
rect 427 -9496 476 -9495
rect -227 -10597 -164 -9522
rect 423 -9506 476 -9496
rect 475 -9558 476 -9506
rect 11372 -9524 11375 -9472
rect 11427 -9524 11434 -9472
rect 11372 -9537 11434 -9524
rect 423 -9568 476 -9558
rect 427 -10075 476 -9568
rect 12463 -10030 12522 -8503
rect 12751 -8998 12806 -8350
rect 15968 -8416 16033 -7326
rect 15968 -8475 15972 -8416
rect 16031 -8475 16033 -8416
rect 15968 -8489 16033 -8475
rect 12751 -9050 12752 -8998
rect 12804 -9050 12806 -8998
rect 12751 -9051 12806 -9050
rect 12752 -9060 12804 -9051
rect 11374 -10052 11433 -10039
rect 427 -10085 480 -10075
rect 427 -10137 428 -10085
rect 427 -10147 480 -10137
rect 11374 -10104 11378 -10052
rect 11430 -10104 11433 -10052
rect 427 -10149 476 -10147
rect -227 -10649 -221 -10597
rect -169 -10649 -164 -10597
rect 11374 -10559 11433 -10104
rect 12463 -10082 12466 -10030
rect 12518 -10082 12522 -10030
rect 12463 -10144 12522 -10082
rect 12463 -10196 12466 -10144
rect 12518 -10196 12522 -10144
rect 12753 -9382 12812 -9369
rect 12753 -9434 12756 -9382
rect 12808 -9434 12812 -9382
rect 12753 -10088 12812 -9434
rect 12753 -10140 12755 -10088
rect 12807 -10140 12812 -10088
rect 12753 -10154 12812 -10140
rect 12463 -10209 12522 -10196
rect 11374 -10611 11376 -10559
rect 11428 -10611 11433 -10559
rect 11374 -10624 11433 -10611
rect -227 -10664 -164 -10649
rect -405 -12282 -404 -12224
rect -405 -12293 -346 -12282
rect 113 -11137 170 -11123
rect 113 -11189 115 -11137
rect 167 -11189 170 -11137
rect 11375 -11163 11426 -11161
rect 113 -12259 170 -11189
rect 11373 -11173 11426 -11163
rect 11425 -11225 11426 -11173
rect 11373 -11235 11426 -11225
rect 425 -11647 480 -11634
rect 425 -11699 427 -11647
rect 479 -11699 480 -11647
rect 425 -12216 480 -11699
rect 11375 -11673 11426 -11235
rect 12463 -11588 12522 -11575
rect 12463 -11640 12466 -11588
rect 12518 -11640 12522 -11588
rect 11375 -11683 11429 -11673
rect 11375 -11735 11377 -11683
rect 11375 -11745 11429 -11735
rect 12463 -11702 12522 -11640
rect 11375 -11748 11426 -11745
rect 113 -12311 115 -12259
rect 167 -12311 170 -12259
rect 424 -12226 480 -12216
rect 476 -12278 480 -12226
rect 12463 -11754 12466 -11702
rect 12518 -11754 12522 -11702
rect 424 -12288 480 -12278
rect 425 -12291 480 -12288
rect 11373 -12261 11435 -12249
rect 113 -12317 170 -12311
rect 11373 -12313 11375 -12261
rect 11427 -12313 11435 -12261
rect 115 -12321 167 -12317
rect 7163 -12347 7215 -12343
rect 7154 -12353 7223 -12347
rect 7154 -12405 7163 -12353
rect 7215 -12405 7223 -12353
rect 424 -12726 476 -12723
rect 424 -12736 479 -12726
rect 424 -12788 427 -12736
rect 424 -12798 479 -12788
rect 424 -13305 476 -12798
rect 7154 -12881 7223 -12405
rect 11373 -12768 11435 -12313
rect 11373 -12820 11380 -12768
rect 11432 -12820 11435 -12768
rect 11373 -12833 11435 -12820
rect 7154 -12933 7165 -12881
rect 7217 -12933 7223 -12881
rect 7154 -12943 7223 -12933
rect 11110 -12884 11178 -12874
rect 11110 -12936 11118 -12884
rect 11170 -12936 11178 -12884
rect 422 -13315 476 -13305
rect 474 -13367 476 -13315
rect 422 -13377 476 -13367
rect 424 -13380 476 -13377
rect 979 -13435 1039 -13425
rect 979 -13487 982 -13435
rect 1034 -13487 1039 -13435
rect 979 -13791 1039 -13487
rect 979 -13843 982 -13791
rect 1034 -13843 1039 -13791
rect 979 -13854 1039 -13843
rect -944 -13889 -886 -13879
rect 11110 -13857 11178 -12936
rect 12463 -13281 12522 -11754
rect 12753 -11644 12812 -11630
rect 12753 -11696 12755 -11644
rect 12807 -11696 12812 -11644
rect 12753 -12350 12812 -11696
rect 12753 -12402 12756 -12350
rect 12808 -12402 12812 -12350
rect 12753 -12415 12812 -12402
rect 12752 -12733 12804 -12724
rect 12463 -13350 12522 -13340
rect 12751 -12734 12806 -12733
rect 12751 -12786 12752 -12734
rect 12804 -12786 12806 -12734
rect 12751 -13434 12806 -12786
rect 12751 -13486 12753 -13434
rect 12805 -13486 12806 -13434
rect 12751 -13497 12806 -13486
rect 11110 -13909 11120 -13857
rect 11172 -13909 11178 -13857
rect 11110 -13925 11178 -13909
rect -1824 -13981 -1769 -13971
<< labels >>
flabel metal1 -3181 -14 -3181 -14 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -1102 -3181 -1102 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -2190 -3181 -2190 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -3278 -3181 -3278 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -4366 -3181 -4366 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -5454 -3181 -5454 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -6542 -3181 -6542 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -7630 -3181 -7630 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -8718 -3181 -8718 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -9806 -3181 -9806 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -10894 -3181 -10894 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -11982 -3181 -11982 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -13070 -3181 -13070 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -14158 -3181 -14158 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 -3181 -555 -3181 -555 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -1643 -3181 -1643 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -2731 -3181 -2731 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -3819 -3181 -3819 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -4907 -3181 -4907 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -5995 -3181 -5995 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -7083 -3181 -7083 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -8171 -3181 -8171 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -9259 -3181 -9259 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -10347 -3181 -10347 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -11435 -3181 -11435 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -12523 -3181 -12523 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -13611 -3181 -13611 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -12 16932 -12 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -1100 16932 -1100 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -2188 16932 -2188 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -3276 16932 -3276 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -4364 16932 -4364 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -5452 16932 -5452 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -6540 16932 -6540 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -7628 16932 -7628 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -8716 16932 -8716 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -9804 16932 -9804 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -10892 16932 -10892 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -11980 16932 -11980 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -13068 16932 -13068 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -14156 16932 -14156 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel metal1 16932 -556 16932 -556 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -1644 16932 -1644 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -2732 16932 -2732 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -3820 16932 -3820 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -4908 16932 -4908 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -5996 16932 -5996 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -7084 16932 -7084 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -8172 16932 -8172 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -9260 16932 -9260 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -10348 16932 -10348 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -11436 16932 -11436 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -12524 16932 -12524 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 16932 -13612 16932 -13612 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
flabel metal1 -3181 -6847 -3181 -6847 1 FreeSans 400 0 0 0 clk
port 1 n
flabel metal1 16932 -828 16932 -828 1 FreeSans 400 0 0 0 B
port 17 n
flabel metal1 16932 -1372 16932 -1372 1 FreeSans 400 0 0 0 B_b
port 16 n
flabel metal1 16932 -1916 16932 -1916 1 FreeSans 400 0 0 0 Bd
port 15 n
flabel metal1 16932 -2460 16932 -2460 1 FreeSans 400 0 0 0 Bd_b
port 14 n
flabel metal1 16932 -4092 16932 -4092 1 FreeSans 400 0 0 0 Ad_b
port 10 n
flabel metal1 16932 -4636 16932 -4636 1 FreeSans 400 0 0 0 Ad
port 11 n
flabel metal1 16932 -5180 16932 -5180 1 FreeSans 400 0 0 0 A_b
port 12 n
flabel metal1 16932 -5724 16932 -5724 1 FreeSans 400 0 0 0 A
port 13 n
flabel metal1 16932 -8444 16932 -8444 1 FreeSans 400 0 0 0 p2
port 5 n
flabel metal1 16932 -8988 16932 -8988 1 FreeSans 400 0 0 0 p2_b
port 4 n
flabel metal1 16932 -9532 16932 -9532 1 FreeSans 400 0 0 0 p2d
port 3 n
flabel metal1 16932 -10076 16932 -10076 1 FreeSans 400 0 0 0 p2d_b
port 2 n
flabel metal1 16932 -11708 16932 -11708 1 FreeSans 400 0 0 0 p1d_b
port 6 n
flabel metal1 16932 -12252 16932 -12252 1 FreeSans 400 0 0 0 p1d
port 7 n
flabel metal1 16932 -12796 16932 -12796 1 FreeSans 400 0 0 0 p1_b
port 8 n
flabel metal1 16932 -13340 16932 -13340 1 FreeSans 400 0 0 0 p1
port 9 n
flabel metal1 -2239 -13088 -2186 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_555/VPWR
flabel metal1 -2240 -13630 -2189 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_555/VGND
rlabel comment -2261 -13612 -2261 -13612 4 sky130_fd_sc_hd__tapvpwrvgnd_1_555/tapvpwrvgnd_1
rlabel metal1 -2261 -13660 -2169 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_555/VGND
rlabel metal1 -2261 -13116 -2169 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_555/VPWR
flabel metal1 -2244 -14165 -2191 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_554/VPWR
flabel metal1 -2241 -13632 -2190 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_554/VGND
rlabel comment -2169 -13612 -2169 -13612 8 sky130_fd_sc_hd__tapvpwrvgnd_1_554/tapvpwrvgnd_1
rlabel metal1 -2261 -13660 -2169 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_554/VGND
rlabel metal1 -2261 -14204 -2169 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_554/VPWR
flabel metal1 -2968 -13085 -2934 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_90/VPWR
flabel metal1 -2968 -13629 -2934 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_90/VGND
flabel nwell -2968 -13085 -2934 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_90/VPB
flabel pwell -2968 -13629 -2934 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_90/VNB
rlabel comment -2997 -13612 -2997 -13612 4 sky130_fd_sc_hd__decap_8_90/decap_8
rlabel metal1 -2997 -13660 -2261 -13564 1 sky130_fd_sc_hd__decap_8_90/VGND
rlabel metal1 -2997 -13116 -2261 -13020 1 sky130_fd_sc_hd__decap_8_90/VPWR
flabel metal1 -2324 -14173 -2290 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_89/VPWR
flabel metal1 -2324 -13629 -2290 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_89/VGND
flabel nwell -2324 -14173 -2290 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_89/VPB
flabel pwell -2324 -13629 -2290 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_89/VNB
rlabel comment -2261 -13612 -2261 -13612 8 sky130_fd_sc_hd__decap_8_89/decap_8
rlabel metal1 -2997 -13660 -2261 -13564 5 sky130_fd_sc_hd__decap_8_89/VGND
rlabel metal1 -2997 -14204 -2261 -14108 5 sky130_fd_sc_hd__decap_8_89/VPWR
flabel metal1 -2135 -13622 -2112 -13603 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_38/VGND
flabel metal1 -2135 -13077 -2115 -13060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_38/VPWR
flabel nwell -2134 -13082 -2109 -13056 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_38/VPB
flabel pwell -2134 -13624 -2112 -13600 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_38/VNB
rlabel comment -2169 -13612 -2169 -13612 4 sky130_fd_sc_hd__fill_4_38/fill_4
rlabel metal1 -2169 -13660 -1801 -13564 1 sky130_fd_sc_hd__fill_4_38/VGND
rlabel metal1 -2169 -13116 -1801 -13020 1 sky130_fd_sc_hd__fill_4_38/VPWR
flabel metal1 -1858 -13621 -1835 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_37/VGND
flabel metal1 -1855 -14164 -1835 -14147 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_37/VPWR
flabel nwell -1861 -14168 -1836 -14142 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_37/VPB
flabel pwell -1858 -13624 -1836 -13600 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_37/VNB
rlabel comment -1801 -13612 -1801 -13612 8 sky130_fd_sc_hd__fill_4_37/fill_4
rlabel metal1 -2169 -13660 -1801 -13564 5 sky130_fd_sc_hd__fill_4_37/VGND
rlabel metal1 -2169 -14204 -1801 -14108 5 sky130_fd_sc_hd__fill_4_37/VPWR
flabel metal1 -1781 -13626 -1728 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_29/VGND
flabel metal1 -1780 -13082 -1728 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_29/VPWR
flabel nwell -1773 -13077 -1739 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_29/VPB
flabel pwell -1770 -13622 -1738 -13600 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_29/VNB
rlabel comment -1801 -13612 -1801 -13612 4 sky130_fd_sc_hd__fill_2_29/fill_2
rlabel metal1 -1801 -13660 -1617 -13564 1 sky130_fd_sc_hd__fill_2_29/VGND
rlabel metal1 -1801 -13116 -1617 -13020 1 sky130_fd_sc_hd__fill_2_29/VPWR
flabel metal1 -1690 -13630 -1637 -13598 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_28/VGND
flabel metal1 -1690 -14173 -1638 -14142 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_28/VPWR
flabel nwell -1679 -14165 -1645 -14147 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_28/VPB
flabel pwell -1680 -13624 -1648 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_28/VNB
rlabel comment -1617 -13612 -1617 -13612 8 sky130_fd_sc_hd__fill_2_28/fill_2
rlabel metal1 -1801 -13660 -1617 -13564 5 sky130_fd_sc_hd__fill_2_28/VGND
rlabel metal1 -1801 -14204 -1617 -14108 5 sky130_fd_sc_hd__fill_2_28/VPWR
flabel metal1 -1597 -13630 -1544 -13598 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_2/VGND
flabel metal1 -1596 -14173 -1544 -14142 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_2/VPWR
flabel nwell -1589 -14165 -1555 -14147 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_2/VPB
flabel pwell -1586 -13624 -1554 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_2/VNB
rlabel comment -1617 -13612 -1617 -13612 2 sky130_fd_sc_hd__fill_2_2/fill_2
rlabel metal1 -1617 -13660 -1433 -13564 5 sky130_fd_sc_hd__fill_2_2/VGND
rlabel metal1 -1617 -14204 -1433 -14108 5 sky130_fd_sc_hd__fill_2_2/VPWR
flabel metal1 -944 -13085 -910 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_23/VPWR
flabel metal1 -944 -13629 -910 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_23/VGND
flabel nwell -944 -13085 -910 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_23/VPB
flabel pwell -944 -13629 -910 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_23/VNB
rlabel comment -881 -13612 -881 -13612 6 sky130_fd_sc_hd__decap_8_23/decap_8
rlabel metal1 -1617 -13660 -881 -13564 1 sky130_fd_sc_hd__decap_8_23/VGND
rlabel metal1 -1617 -13116 -881 -13020 1 sky130_fd_sc_hd__decap_8_23/VPWR
flabel metal1 -1404 -13629 -1370 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_126/VGND
flabel metal1 -1404 -14173 -1370 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_126/VPWR
flabel nwell -1404 -14173 -1370 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_126/VPB
flabel pwell -1404 -13629 -1370 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_126/VNB
rlabel comment -1433 -13612 -1433 -13612 2 sky130_fd_sc_hd__decap_4_126/decap_4
rlabel metal1 -1433 -13660 -1065 -13564 5 sky130_fd_sc_hd__decap_4_126/VGND
rlabel metal1 -1433 -14204 -1065 -14108 5 sky130_fd_sc_hd__decap_4_126/VPWR
flabel metal1 -1043 -14165 -990 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_257/VPWR
flabel metal1 -1044 -13632 -993 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_257/VGND
rlabel comment -1065 -13612 -1065 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_257/tapvpwrvgnd_1
rlabel metal1 -1065 -13660 -973 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_257/VGND
rlabel metal1 -1065 -14204 -973 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_257/VPWR
flabel metal1 -675 -14165 -622 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_256/VPWR
flabel metal1 -676 -13632 -625 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_256/VGND
rlabel comment -697 -13612 -697 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_256/tapvpwrvgnd_1
rlabel metal1 -697 -13660 -605 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_256/VGND
rlabel metal1 -697 -14204 -605 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_256/VPWR
flabel locali -853 -13731 -819 -13697 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/Y
flabel locali -853 -13799 -819 -13765 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/Y
flabel locali -853 -13867 -819 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/Y
flabel locali -945 -13867 -911 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/B
flabel locali -761 -13867 -727 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/A
flabel nwell -945 -14173 -911 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VPB
flabel pwell -945 -13629 -911 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VNB
flabel metal1 -945 -13629 -911 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VGND
flabel metal1 -945 -14173 -911 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VPWR
rlabel comment -973 -13612 -973 -13612 2 sky130_fd_sc_hd__nand2_1_2/nand2_1
rlabel metal1 -973 -13660 -697 -13564 5 sky130_fd_sc_hd__nand2_1_2/VGND
rlabel metal1 -973 -14204 -697 -14108 5 sky130_fd_sc_hd__nand2_1_2/VPWR
flabel metal1 -208 -13085 -174 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_24/VPWR
flabel metal1 -208 -13629 -174 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_24/VGND
flabel nwell -208 -13085 -174 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_24/VPB
flabel pwell -208 -13629 -174 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_24/VNB
rlabel comment -145 -13612 -145 -13612 6 sky130_fd_sc_hd__decap_8_24/decap_8
rlabel metal1 -881 -13660 -145 -13564 1 sky130_fd_sc_hd__decap_8_24/VGND
rlabel metal1 -881 -13116 -145 -13020 1 sky130_fd_sc_hd__decap_8_24/VPWR
flabel metal1 -576 -13629 -542 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_128/VGND
flabel metal1 -576 -14173 -542 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_128/VPWR
flabel nwell -576 -14173 -542 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_128/VPB
flabel pwell -576 -13629 -542 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_128/VNB
rlabel comment -605 -13612 -605 -13612 2 sky130_fd_sc_hd__decap_4_128/decap_4
rlabel metal1 -605 -13660 -237 -13564 5 sky130_fd_sc_hd__decap_4_128/VGND
rlabel metal1 -605 -14204 -237 -14108 5 sky130_fd_sc_hd__decap_4_128/VPWR
flabel metal1 -128 -13088 -75 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_277/VPWR
flabel metal1 -125 -13630 -74 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_277/VGND
rlabel comment -53 -13612 -53 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_277/tapvpwrvgnd_1
rlabel metal1 -145 -13660 -53 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_277/VGND
rlabel metal1 -145 -13116 -53 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_277/VPWR
flabel metal1 332 -13088 385 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_276/VPWR
flabel metal1 335 -13630 386 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_276/VGND
rlabel comment 407 -13612 407 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_276/tapvpwrvgnd_1
rlabel metal1 315 -13660 407 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_276/VGND
rlabel metal1 315 -13116 407 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_276/VPWR
flabel metal1 521 -14165 574 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_255/VPWR
flabel metal1 520 -13632 571 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_255/VGND
rlabel comment 499 -13612 499 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_255/tapvpwrvgnd_1
rlabel metal1 499 -13660 591 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_255/VGND
rlabel metal1 499 -14204 591 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_255/VPWR
flabel metal1 -215 -14165 -162 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_254/VPWR
flabel metal1 -216 -13632 -165 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_254/VGND
rlabel comment -237 -13612 -237 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_254/tapvpwrvgnd_1
rlabel metal1 -237 -13660 -145 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_254/VGND
rlabel metal1 -237 -14204 -145 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_254/VPWR
flabel metal1 252 -13629 286 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_137/VGND
flabel metal1 252 -13085 286 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_137/VPWR
flabel nwell 252 -13085 286 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_137/VPB
flabel pwell 252 -13629 286 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_137/VNB
rlabel comment 315 -13612 315 -13612 6 sky130_fd_sc_hd__decap_4_137/decap_4
rlabel metal1 -53 -13660 315 -13564 1 sky130_fd_sc_hd__decap_4_137/VGND
rlabel metal1 -53 -13116 315 -13020 1 sky130_fd_sc_hd__decap_4_137/VPWR
flabel locali 68 -13867 102 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/A
flabel locali 160 -13867 194 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/A
flabel locali 436 -13799 470 -13765 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/Y
flabel locali -24 -13867 10 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/A
flabel locali 436 -13935 470 -13901 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/Y
flabel locali 344 -13867 378 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/A
flabel locali 252 -13867 286 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/A
flabel locali 436 -13867 470 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_6/Y
flabel pwell -116 -13629 -82 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_6/VNB
flabel nwell -116 -14173 -82 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_6/VPB
flabel metal1 -116 -14173 -82 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_6/VPWR
flabel metal1 -116 -13629 -82 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_6/VGND
rlabel comment -145 -13612 -145 -13612 2 sky130_fd_sc_hd__clkinv_4_6/clkinv_4
rlabel metal1 -145 -13660 499 -13564 5 sky130_fd_sc_hd__clkinv_4_6/VGND
rlabel metal1 -145 -14204 499 -14108 5 sky130_fd_sc_hd__clkinv_4_6/VPWR
flabel locali 1079 -13391 1113 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/A
flabel locali 433 -13187 467 -13153 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/X
flabel locali 433 -13255 467 -13221 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/X
flabel locali 433 -13323 467 -13289 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/X
flabel locali 433 -13391 467 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/X
flabel locali 433 -13459 467 -13425 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/X
flabel locali 433 -13527 467 -13493 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/X
flabel pwell 1079 -13629 1113 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/VNB
flabel nwell 1079 -13085 1113 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/VPB
flabel metal1 1079 -13629 1113 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/VGND
flabel metal1 1079 -13085 1113 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_104/VPWR
rlabel comment 1143 -13612 1143 -13612 6 sky130_fd_sc_hd__clkdlybuf4s50_1_104/clkdlybuf4s50_1
rlabel metal1 407 -13660 1143 -13564 1 sky130_fd_sc_hd__clkdlybuf4s50_1_104/VGND
rlabel metal1 407 -13116 1143 -13020 1 sky130_fd_sc_hd__clkdlybuf4s50_1_104/VPWR
flabel metal1 620 -13629 654 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_127/VGND
flabel metal1 620 -14173 654 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_127/VPWR
flabel nwell 620 -14173 654 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_127/VPB
flabel pwell 620 -13629 654 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_127/VNB
rlabel comment 591 -13612 591 -13612 2 sky130_fd_sc_hd__decap_4_127/decap_4
rlabel metal1 591 -13660 959 -13564 5 sky130_fd_sc_hd__decap_4_127/VGND
rlabel metal1 591 -14204 959 -14108 5 sky130_fd_sc_hd__decap_4_127/VPWR
flabel metal1 1160 -13088 1213 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_280/VPWR
flabel metal1 1163 -13630 1214 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_280/VGND
rlabel comment 1235 -13612 1235 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_280/tapvpwrvgnd_1
rlabel metal1 1143 -13660 1235 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_280/VGND
rlabel metal1 1143 -13116 1235 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_280/VPWR
flabel metal1 1620 -13088 1673 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_279/VPWR
flabel metal1 1623 -13630 1674 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_279/VGND
rlabel comment 1695 -13612 1695 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_279/tapvpwrvgnd_1
rlabel metal1 1603 -13660 1695 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_279/VGND
rlabel metal1 1603 -13116 1695 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_279/VPWR
flabel metal1 1349 -14165 1402 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_259/VPWR
flabel metal1 1348 -13632 1399 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_259/VGND
rlabel comment 1327 -13612 1327 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_259/tapvpwrvgnd_1
rlabel metal1 1327 -13660 1419 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_259/VGND
rlabel metal1 1327 -14204 1419 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_259/VPWR
flabel metal1 981 -14165 1034 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_258/VPWR
flabel metal1 980 -13632 1031 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_258/VGND
rlabel comment 959 -13612 959 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_258/tapvpwrvgnd_1
rlabel metal1 959 -13660 1051 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_258/VGND
rlabel metal1 959 -14204 1051 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_258/VPWR
flabel metal1 1540 -13629 1574 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_139/VGND
flabel metal1 1540 -13085 1574 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_139/VPWR
flabel nwell 1540 -13085 1574 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_139/VPB
flabel pwell 1540 -13629 1574 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_139/VNB
rlabel comment 1603 -13612 1603 -13612 6 sky130_fd_sc_hd__decap_4_139/decap_4
rlabel metal1 1235 -13660 1603 -13564 1 sky130_fd_sc_hd__decap_4_139/VGND
rlabel metal1 1235 -13116 1603 -13020 1 sky130_fd_sc_hd__decap_4_139/VPWR
flabel metal1 1448 -13629 1482 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_129/VGND
flabel metal1 1448 -14173 1482 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_129/VPWR
flabel nwell 1448 -14173 1482 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_129/VPB
flabel pwell 1448 -13629 1482 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_129/VNB
rlabel comment 1419 -13612 1419 -13612 2 sky130_fd_sc_hd__decap_4_129/decap_4
rlabel metal1 1419 -13660 1787 -13564 5 sky130_fd_sc_hd__decap_4_129/VGND
rlabel metal1 1419 -14204 1787 -14108 5 sky130_fd_sc_hd__decap_4_129/VPWR
flabel locali 1264 -13799 1298 -13765 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/Y
flabel locali 1264 -13867 1298 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/Y
flabel locali 1172 -13935 1206 -13901 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/Y
flabel locali 1172 -13867 1206 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/Y
flabel locali 1172 -13799 1206 -13765 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/Y
flabel locali 1080 -13731 1114 -13697 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/A
flabel locali 1080 -13799 1114 -13765 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/A
flabel locali 1080 -13867 1114 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_2/A
flabel nwell 1080 -14173 1114 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_2/VPB
flabel pwell 1080 -13629 1114 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_2/VNB
flabel metal1 1080 -13629 1114 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_2/VGND
flabel metal1 1080 -14173 1114 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_2/VPWR
rlabel comment 1051 -13612 1051 -13612 2 sky130_fd_sc_hd__clkinv_1_2/clkinv_1
rlabel metal1 1051 -13660 1327 -13564 5 sky130_fd_sc_hd__clkinv_1_2/VGND
rlabel metal1 1051 -14204 1327 -14108 5 sky130_fd_sc_hd__clkinv_1_2/VPWR
flabel metal1 2448 -13088 2501 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_278/VPWR
flabel metal1 2451 -13630 2502 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_278/VGND
rlabel comment 2523 -13612 2523 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_278/tapvpwrvgnd_1
rlabel metal1 2431 -13660 2523 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_278/VGND
rlabel metal1 2431 -13116 2523 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_278/VPWR
flabel metal1 2269 -14165 2322 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_261/VPWR
flabel metal1 2268 -13632 2319 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_261/VGND
rlabel comment 2247 -13612 2247 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_261/tapvpwrvgnd_1
rlabel metal1 2247 -13660 2339 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_261/VGND
rlabel metal1 2247 -14204 2339 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_261/VPWR
flabel metal1 1809 -14165 1862 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_260/VPWR
flabel metal1 1808 -13632 1859 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_260/VGND
rlabel comment 1787 -13612 1787 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_260/tapvpwrvgnd_1
rlabel metal1 1787 -13660 1879 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_260/VGND
rlabel metal1 1787 -14204 1879 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_260/VPWR
flabel metal1 1724 -13085 1758 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_140/VPWR
flabel metal1 1724 -13629 1758 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_140/VGND
flabel nwell 1724 -13085 1758 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_140/VPB
flabel pwell 1724 -13629 1758 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_140/VNB
rlabel comment 1695 -13612 1695 -13612 4 sky130_fd_sc_hd__decap_8_140/decap_8
rlabel metal1 1695 -13660 2431 -13564 1 sky130_fd_sc_hd__decap_8_140/VGND
rlabel metal1 1695 -13116 2431 -13020 1 sky130_fd_sc_hd__decap_8_140/VPWR
flabel metal1 1908 -13629 1942 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_130/VGND
flabel metal1 1908 -14173 1942 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_130/VPWR
flabel nwell 1908 -14173 1942 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_130/VPB
flabel pwell 1908 -13629 1942 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_130/VNB
rlabel comment 1879 -13612 1879 -13612 2 sky130_fd_sc_hd__decap_4_130/decap_4
rlabel metal1 1879 -13660 2247 -13564 5 sky130_fd_sc_hd__decap_4_130/VGND
rlabel metal1 1879 -14204 2247 -14108 5 sky130_fd_sc_hd__decap_4_130/VPWR
flabel locali 2369 -13867 2403 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A
flabel locali 3015 -14071 3049 -14037 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/X
flabel locali 3015 -14003 3049 -13969 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/X
flabel locali 3015 -13935 3049 -13901 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/X
flabel locali 3015 -13867 3049 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/X
flabel locali 3015 -13799 3049 -13765 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/X
flabel locali 3015 -13731 3049 -13697 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/X
flabel pwell 2369 -13629 2403 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/VNB
flabel nwell 2369 -14173 2403 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/VPB
flabel metal1 2369 -13629 2403 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/VGND
flabel metal1 2369 -14173 2403 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_100/VPWR
rlabel comment 2339 -13612 2339 -13612 2 sky130_fd_sc_hd__clkdlybuf4s50_1_100/clkdlybuf4s50_1
rlabel metal1 2339 -13660 3075 -13564 5 sky130_fd_sc_hd__clkdlybuf4s50_1_100/VGND
rlabel metal1 2339 -14204 3075 -14108 5 sky130_fd_sc_hd__clkdlybuf4s50_1_100/VPWR
flabel metal1 2828 -13629 2862 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_138/VGND
flabel metal1 2828 -13085 2862 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_138/VPWR
flabel nwell 2828 -13085 2862 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_138/VPB
flabel pwell 2828 -13629 2862 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_138/VNB
rlabel comment 2891 -13612 2891 -13612 6 sky130_fd_sc_hd__decap_4_138/decap_4
rlabel metal1 2523 -13660 2891 -13564 1 sky130_fd_sc_hd__decap_4_138/VGND
rlabel metal1 2523 -13116 2891 -13020 1 sky130_fd_sc_hd__decap_4_138/VPWR
flabel metal1 2908 -13088 2961 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_283/VPWR
flabel metal1 2911 -13630 2962 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_283/VGND
rlabel comment 2983 -13612 2983 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_283/tapvpwrvgnd_1
rlabel metal1 2891 -13660 2983 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_283/VGND
rlabel metal1 2891 -13116 2983 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_283/VPWR
flabel metal1 3097 -14165 3150 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_263/VPWR
flabel metal1 3096 -13632 3147 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_263/VGND
rlabel comment 3075 -13612 3075 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_263/tapvpwrvgnd_1
rlabel metal1 3075 -13660 3167 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_263/VGND
rlabel metal1 3075 -14204 3167 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_263/VPWR
flabel metal1 3557 -14165 3610 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_262/VPWR
flabel metal1 3556 -13632 3607 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_262/VGND
rlabel comment 3535 -13612 3535 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_262/tapvpwrvgnd_1
rlabel metal1 3535 -13660 3627 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_262/VGND
rlabel metal1 3535 -14204 3627 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_262/VPWR
flabel metal1 3662 -13622 3694 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_18/VGND
flabel metal1 3656 -14167 3694 -14135 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_18/VPWR
flabel nwell 3647 -14165 3704 -14134 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_18/VPB
flabel pwell 3653 -13622 3697 -13588 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_18/VNB
rlabel comment 3627 -13612 3627 -13612 2 sky130_fd_sc_hd__fill_8_18/fill_8
rlabel metal1 3627 -13660 4363 -13564 5 sky130_fd_sc_hd__fill_8_18/VGND
rlabel metal1 3627 -14204 4363 -14108 5 sky130_fd_sc_hd__fill_8_18/VPWR
flabel metal1 3196 -13629 3230 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_131/VGND
flabel metal1 3196 -14173 3230 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_131/VPWR
flabel nwell 3196 -14173 3230 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_131/VPB
flabel pwell 3196 -13629 3230 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_131/VNB
rlabel comment 3167 -13612 3167 -13612 2 sky130_fd_sc_hd__decap_4_131/decap_4
rlabel metal1 3167 -13660 3535 -13564 5 sky130_fd_sc_hd__decap_4_131/VGND
rlabel metal1 3167 -14204 3535 -14108 5 sky130_fd_sc_hd__decap_4_131/VPWR
flabel locali 3655 -13391 3689 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/A
flabel locali 3009 -13187 3043 -13153 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
flabel locali 3009 -13255 3043 -13221 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
flabel locali 3009 -13323 3043 -13289 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
flabel locali 3009 -13391 3043 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
flabel locali 3009 -13459 3043 -13425 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
flabel locali 3009 -13527 3043 -13493 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
flabel pwell 3655 -13629 3689 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/VNB
flabel nwell 3655 -13085 3689 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/VPB
flabel metal1 3655 -13629 3689 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/VGND
flabel metal1 3655 -13085 3689 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_107/VPWR
rlabel comment 3719 -13612 3719 -13612 6 sky130_fd_sc_hd__clkdlybuf4s50_1_107/clkdlybuf4s50_1
rlabel metal1 2983 -13660 3719 -13564 1 sky130_fd_sc_hd__clkdlybuf4s50_1_107/VGND
rlabel metal1 2983 -13116 3719 -13020 1 sky130_fd_sc_hd__clkdlybuf4s50_1_107/VPWR
flabel metal1 4196 -13088 4249 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_282/VPWR
flabel metal1 4199 -13630 4250 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_282/VGND
rlabel comment 4271 -13612 4271 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_282/tapvpwrvgnd_1
rlabel metal1 4179 -13660 4271 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_282/VGND
rlabel metal1 4179 -13116 4271 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_282/VPWR
flabel metal1 3736 -13088 3789 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_281/VPWR
flabel metal1 3739 -13630 3790 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_281/VGND
rlabel comment 3811 -13612 3811 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_281/tapvpwrvgnd_1
rlabel metal1 3719 -13660 3811 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_281/VGND
rlabel metal1 3719 -13116 3811 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_281/VPWR
flabel metal1 4300 -13085 4334 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_142/VPWR
flabel metal1 4300 -13629 4334 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_142/VGND
flabel nwell 4300 -13085 4334 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_142/VPB
flabel pwell 4300 -13629 4334 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_142/VNB
rlabel comment 4271 -13612 4271 -13612 4 sky130_fd_sc_hd__decap_8_142/decap_8
rlabel metal1 4271 -13660 5007 -13564 1 sky130_fd_sc_hd__decap_8_142/VGND
rlabel metal1 4271 -13116 5007 -13020 1 sky130_fd_sc_hd__decap_8_142/VPWR
flabel metal1 4116 -13629 4150 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_140/VGND
flabel metal1 4116 -13085 4150 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_140/VPWR
flabel nwell 4116 -13085 4150 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_140/VPB
flabel pwell 4116 -13629 4150 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_140/VNB
rlabel comment 4179 -13612 4179 -13612 6 sky130_fd_sc_hd__decap_4_140/decap_4
rlabel metal1 3811 -13660 4179 -13564 1 sky130_fd_sc_hd__decap_4_140/VGND
rlabel metal1 3811 -13116 4179 -13020 1 sky130_fd_sc_hd__decap_4_140/VPWR
flabel metal1 4392 -13629 4426 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_18/VGND
flabel metal1 4392 -14173 4426 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_18/VPWR
flabel nwell 4392 -14173 4426 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_18/VPB
flabel pwell 4392 -13629 4426 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_18/VNB
rlabel comment 4363 -13612 4363 -13612 2 sky130_fd_sc_hd__decap_12_18/decap_12
rlabel metal1 4363 -13660 5467 -13564 5 sky130_fd_sc_hd__decap_12_18/VGND
rlabel metal1 4363 -14204 5467 -14108 5 sky130_fd_sc_hd__decap_12_18/VPWR
flabel metal1 5024 -13088 5077 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_286/VPWR
flabel metal1 5027 -13630 5078 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_286/VGND
rlabel comment 5099 -13612 5099 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_286/tapvpwrvgnd_1
rlabel metal1 5007 -13660 5099 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_286/VGND
rlabel metal1 5007 -13116 5099 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_286/VPWR
flabel metal1 5484 -13088 5537 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_285/VPWR
flabel metal1 5487 -13630 5538 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_285/VGND
rlabel comment 5559 -13612 5559 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_285/tapvpwrvgnd_1
rlabel metal1 5467 -13660 5559 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_285/VGND
rlabel metal1 5467 -13116 5559 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_285/VPWR
flabel metal1 5501 -13621 5524 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_8/VGND
flabel metal1 5501 -14164 5521 -14147 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_8/VPWR
flabel nwell 5502 -14168 5527 -14142 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_8/VPB
flabel pwell 5502 -13624 5524 -13600 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_8/VNB
rlabel comment 5467 -13612 5467 -13612 2 sky130_fd_sc_hd__fill_4_8/fill_4
rlabel metal1 5467 -13660 5835 -13564 5 sky130_fd_sc_hd__fill_4_8/VGND
rlabel metal1 5467 -14204 5835 -14108 5 sky130_fd_sc_hd__fill_4_8/VPWR
flabel metal1 5404 -13629 5438 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_142/VGND
flabel metal1 5404 -13085 5438 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_142/VPWR
flabel nwell 5404 -13085 5438 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_142/VPB
flabel pwell 5404 -13629 5438 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_142/VNB
rlabel comment 5467 -13612 5467 -13612 6 sky130_fd_sc_hd__decap_4_142/decap_4
rlabel metal1 5099 -13660 5467 -13564 1 sky130_fd_sc_hd__decap_4_142/VGND
rlabel metal1 5099 -13116 5467 -13020 1 sky130_fd_sc_hd__decap_4_142/VPWR
flabel metal1 6312 -13088 6365 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_284/VPWR
flabel metal1 6315 -13630 6366 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_284/VGND
rlabel comment 6387 -13612 6387 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_284/tapvpwrvgnd_1
rlabel metal1 6295 -13660 6387 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_284/VGND
rlabel metal1 6295 -13116 6387 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_284/VPWR
flabel metal1 6317 -14165 6370 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_264/VPWR
flabel metal1 6316 -13632 6367 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_264/VGND
rlabel comment 6295 -13612 6295 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_264/tapvpwrvgnd_1
rlabel metal1 6295 -13660 6387 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_264/VGND
rlabel metal1 6295 -14204 6387 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_264/VPWR
flabel metal1 5961 -13621 5984 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_9/VGND
flabel metal1 5961 -14164 5981 -14147 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_9/VPWR
flabel nwell 5962 -14168 5987 -14142 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_9/VPB
flabel pwell 5962 -13624 5984 -13600 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_9/VNB
rlabel comment 5927 -13612 5927 -13612 2 sky130_fd_sc_hd__fill_4_9/fill_4
rlabel metal1 5927 -13660 6295 -13564 5 sky130_fd_sc_hd__fill_4_9/VGND
rlabel metal1 5927 -14204 6295 -14108 5 sky130_fd_sc_hd__fill_4_9/VPWR
flabel metal1 5857 -14169 5893 -14139 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_36/VPWR
flabel metal1 5857 -13628 5893 -13599 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_36/VGND
flabel nwell 5866 -14163 5886 -14146 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_36/VPB
flabel pwell 5863 -13623 5887 -13601 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_36/VNB
rlabel comment 5835 -13612 5835 -13612 2 sky130_fd_sc_hd__fill_1_36/fill_1
rlabel metal1 5835 -13660 5927 -13564 5 sky130_fd_sc_hd__fill_1_36/VGND
rlabel metal1 5835 -14204 5927 -14108 5 sky130_fd_sc_hd__fill_1_36/VPWR
flabel locali 6231 -13391 6265 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/A
flabel locali 5585 -13187 5619 -13153 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X
flabel locali 5585 -13255 5619 -13221 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X
flabel locali 5585 -13323 5619 -13289 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X
flabel locali 5585 -13391 5619 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X
flabel locali 5585 -13459 5619 -13425 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X
flabel locali 5585 -13527 5619 -13493 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X
flabel pwell 6231 -13629 6265 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/VNB
flabel nwell 6231 -13085 6265 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/VPB
flabel metal1 6231 -13629 6265 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/VGND
flabel metal1 6231 -13085 6265 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_108/VPWR
rlabel comment 6295 -13612 6295 -13612 6 sky130_fd_sc_hd__clkdlybuf4s50_1_108/clkdlybuf4s50_1
rlabel metal1 5559 -13660 6295 -13564 1 sky130_fd_sc_hd__clkdlybuf4s50_1_108/VGND
rlabel metal1 5559 -13116 6295 -13020 1 sky130_fd_sc_hd__clkdlybuf4s50_1_108/VPWR
flabel metal1 6692 -13629 6726 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_141/VGND
flabel metal1 6692 -13085 6726 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_141/VPWR
flabel nwell 6692 -13085 6726 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_141/VPB
flabel pwell 6692 -13629 6726 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_141/VNB
rlabel comment 6755 -13612 6755 -13612 6 sky130_fd_sc_hd__decap_4_141/decap_4
rlabel metal1 6387 -13660 6755 -13564 1 sky130_fd_sc_hd__decap_4_141/VGND
rlabel metal1 6387 -13116 6755 -13020 1 sky130_fd_sc_hd__decap_4_141/VPWR
flabel metal1 6416 -13629 6450 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_132/VGND
flabel metal1 6416 -14173 6450 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_132/VPWR
flabel nwell 6416 -14173 6450 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_132/VPB
flabel pwell 6416 -13629 6450 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_132/VNB
rlabel comment 6387 -13612 6387 -13612 2 sky130_fd_sc_hd__decap_4_132/decap_4
rlabel metal1 6387 -13660 6755 -13564 5 sky130_fd_sc_hd__decap_4_132/VGND
rlabel metal1 6387 -14204 6755 -14108 5 sky130_fd_sc_hd__decap_4_132/VPWR
flabel metal1 6772 -13088 6825 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_289/VPWR
flabel metal1 6775 -13630 6826 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_289/VGND
rlabel comment 6847 -13612 6847 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_289/tapvpwrvgnd_1
rlabel metal1 6755 -13660 6847 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_289/VGND
rlabel metal1 6755 -13116 6847 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_289/VPWR
flabel metal1 6777 -14165 6830 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_265/VPWR
flabel metal1 6776 -13632 6827 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_265/VGND
rlabel comment 6755 -13612 6755 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_265/tapvpwrvgnd_1
rlabel metal1 6755 -13660 6847 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_265/VGND
rlabel metal1 6755 -14204 6847 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_265/VPWR
flabel metal1 6876 -13085 6910 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_152/VPWR
flabel metal1 6876 -13629 6910 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_152/VGND
flabel nwell 6876 -13085 6910 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_152/VPB
flabel pwell 6876 -13629 6910 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_152/VNB
rlabel comment 6847 -13612 6847 -13612 4 sky130_fd_sc_hd__decap_8_152/decap_8
rlabel metal1 6847 -13660 7583 -13564 1 sky130_fd_sc_hd__decap_8_152/VGND
rlabel metal1 6847 -13116 7583 -13020 1 sky130_fd_sc_hd__decap_8_152/VPWR
flabel locali 6877 -13867 6911 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A
flabel locali 7523 -14071 7557 -14037 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/X
flabel locali 7523 -14003 7557 -13969 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/X
flabel locali 7523 -13935 7557 -13901 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/X
flabel locali 7523 -13867 7557 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/X
flabel locali 7523 -13799 7557 -13765 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/X
flabel locali 7523 -13731 7557 -13697 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/X
flabel pwell 6877 -13629 6911 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/VNB
flabel nwell 6877 -14173 6911 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/VPB
flabel metal1 6877 -13629 6911 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/VGND
flabel metal1 6877 -14173 6911 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_101/VPWR
rlabel comment 6847 -13612 6847 -13612 2 sky130_fd_sc_hd__clkdlybuf4s50_1_101/clkdlybuf4s50_1
rlabel metal1 6847 -13660 7583 -13564 5 sky130_fd_sc_hd__clkdlybuf4s50_1_101/VGND
rlabel metal1 6847 -14204 7583 -14108 5 sky130_fd_sc_hd__clkdlybuf4s50_1_101/VPWR
flabel metal1 8060 -13088 8113 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_288/VPWR
flabel metal1 8063 -13630 8114 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_288/VGND
rlabel comment 8135 -13612 8135 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_288/tapvpwrvgnd_1
rlabel metal1 8043 -13660 8135 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_288/VGND
rlabel metal1 8043 -13116 8135 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_288/VPWR
flabel metal1 7600 -13088 7653 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_287/VPWR
flabel metal1 7603 -13630 7654 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_287/VGND
rlabel comment 7675 -13612 7675 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_287/tapvpwrvgnd_1
rlabel metal1 7583 -13660 7675 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_287/VGND
rlabel metal1 7583 -13116 7675 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_287/VPWR
flabel metal1 7605 -14165 7658 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_267/VPWR
flabel metal1 7604 -13632 7655 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_267/VGND
rlabel comment 7583 -13612 7583 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_267/tapvpwrvgnd_1
rlabel metal1 7583 -13660 7675 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_267/VGND
rlabel metal1 7583 -14204 7675 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_267/VPWR
flabel metal1 8065 -14165 8118 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_266/VPWR
flabel metal1 8064 -13632 8115 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_266/VGND
rlabel comment 8043 -13612 8043 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_266/tapvpwrvgnd_1
rlabel metal1 8043 -13660 8135 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_266/VGND
rlabel metal1 8043 -14204 8135 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_266/VPWR
flabel metal1 7980 -13629 8014 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_143/VGND
flabel metal1 7980 -13085 8014 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_143/VPWR
flabel nwell 7980 -13085 8014 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_143/VPB
flabel pwell 7980 -13629 8014 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_143/VNB
rlabel comment 8043 -13612 8043 -13612 6 sky130_fd_sc_hd__decap_4_143/decap_4
rlabel metal1 7675 -13660 8043 -13564 1 sky130_fd_sc_hd__decap_4_143/VGND
rlabel metal1 7675 -13116 8043 -13020 1 sky130_fd_sc_hd__decap_4_143/VPWR
flabel metal1 7704 -13629 7738 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_133/VGND
flabel metal1 7704 -14173 7738 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_133/VPWR
flabel nwell 7704 -14173 7738 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_133/VPB
flabel pwell 7704 -13629 7738 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_133/VNB
rlabel comment 7675 -13612 7675 -13612 2 sky130_fd_sc_hd__decap_4_133/decap_4
rlabel metal1 7675 -13660 8043 -13564 5 sky130_fd_sc_hd__decap_4_133/VGND
rlabel metal1 7675 -14204 8043 -14108 5 sky130_fd_sc_hd__decap_4_133/VPWR
flabel locali 8807 -13391 8841 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/A
flabel locali 8161 -13187 8195 -13153 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X
flabel locali 8161 -13255 8195 -13221 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X
flabel locali 8161 -13323 8195 -13289 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X
flabel locali 8161 -13391 8195 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X
flabel locali 8161 -13459 8195 -13425 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X
flabel locali 8161 -13527 8195 -13493 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X
flabel pwell 8807 -13629 8841 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/VNB
flabel nwell 8807 -13085 8841 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/VPB
flabel metal1 8807 -13629 8841 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/VGND
flabel metal1 8807 -13085 8841 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_109/VPWR
rlabel comment 8871 -13612 8871 -13612 6 sky130_fd_sc_hd__clkdlybuf4s50_1_109/clkdlybuf4s50_1
rlabel metal1 8135 -13660 8871 -13564 1 sky130_fd_sc_hd__clkdlybuf4s50_1_109/VGND
rlabel metal1 8135 -13116 8871 -13020 1 sky130_fd_sc_hd__clkdlybuf4s50_1_109/VPWR
flabel locali 8165 -13867 8199 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A
flabel locali 8811 -14071 8845 -14037 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/X
flabel locali 8811 -14003 8845 -13969 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/X
flabel locali 8811 -13935 8845 -13901 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/X
flabel locali 8811 -13867 8845 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/X
flabel locali 8811 -13799 8845 -13765 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/X
flabel locali 8811 -13731 8845 -13697 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/X
flabel pwell 8165 -13629 8199 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/VNB
flabel nwell 8165 -14173 8199 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/VPB
flabel metal1 8165 -13629 8199 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/VGND
flabel metal1 8165 -14173 8199 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_102/VPWR
rlabel comment 8135 -13612 8135 -13612 2 sky130_fd_sc_hd__clkdlybuf4s50_1_102/clkdlybuf4s50_1
rlabel metal1 8135 -13660 8871 -13564 5 sky130_fd_sc_hd__clkdlybuf4s50_1_102/VGND
rlabel metal1 8135 -14204 8871 -14108 5 sky130_fd_sc_hd__clkdlybuf4s50_1_102/VPWR
flabel metal1 8888 -13088 8941 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_292/VPWR
flabel metal1 8891 -13630 8942 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_292/VGND
rlabel comment 8963 -13612 8963 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_292/tapvpwrvgnd_1
rlabel metal1 8871 -13660 8963 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_292/VGND
rlabel metal1 8871 -13116 8963 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_292/VPWR
flabel metal1 8893 -14165 8946 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_268/VPWR
flabel metal1 8892 -13632 8943 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_268/VGND
rlabel comment 8871 -13612 8871 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_268/tapvpwrvgnd_1
rlabel metal1 8871 -13660 8963 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_268/VGND
rlabel metal1 8871 -14204 8963 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_268/VPWR
flabel metal1 9268 -13629 9302 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_144/VGND
flabel metal1 9268 -13085 9302 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_144/VPWR
flabel nwell 9268 -13085 9302 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_144/VPB
flabel pwell 9268 -13629 9302 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_144/VNB
rlabel comment 9331 -13612 9331 -13612 6 sky130_fd_sc_hd__decap_4_144/decap_4
rlabel metal1 8963 -13660 9331 -13564 1 sky130_fd_sc_hd__decap_4_144/VGND
rlabel metal1 8963 -13116 9331 -13020 1 sky130_fd_sc_hd__decap_4_144/VPWR
flabel metal1 8992 -13629 9026 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_134/VGND
flabel metal1 8992 -14173 9026 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_134/VPWR
flabel nwell 8992 -14173 9026 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_134/VPB
flabel pwell 8992 -13629 9026 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_134/VNB
rlabel comment 8963 -13612 8963 -13612 2 sky130_fd_sc_hd__decap_4_134/decap_4
rlabel metal1 8963 -13660 9331 -13564 5 sky130_fd_sc_hd__decap_4_134/VGND
rlabel metal1 8963 -14204 9331 -14108 5 sky130_fd_sc_hd__decap_4_134/VPWR
flabel metal1 9348 -13088 9401 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_291/VPWR
flabel metal1 9351 -13630 9402 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_291/VGND
rlabel comment 9423 -13612 9423 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_291/tapvpwrvgnd_1
rlabel metal1 9331 -13660 9423 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_291/VGND
rlabel metal1 9331 -13116 9423 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_291/VPWR
flabel metal1 9353 -14165 9406 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_269/VPWR
flabel metal1 9352 -13632 9403 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_269/VGND
rlabel comment 9331 -13612 9331 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_269/tapvpwrvgnd_1
rlabel metal1 9331 -13660 9423 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_269/VGND
rlabel metal1 9331 -14204 9423 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_269/VPWR
flabel metal1 9452 -13085 9486 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_161/VPWR
flabel metal1 9452 -13629 9486 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_161/VGND
flabel nwell 9452 -13085 9486 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_161/VPB
flabel pwell 9452 -13629 9486 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_161/VNB
rlabel comment 9423 -13612 9423 -13612 4 sky130_fd_sc_hd__decap_8_161/decap_8
rlabel metal1 9423 -13660 10159 -13564 1 sky130_fd_sc_hd__decap_8_161/VGND
rlabel metal1 9423 -13116 10159 -13020 1 sky130_fd_sc_hd__decap_8_161/VPWR
flabel locali 9453 -13867 9487 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A
flabel locali 10099 -14071 10133 -14037 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/X
flabel locali 10099 -14003 10133 -13969 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/X
flabel locali 10099 -13935 10133 -13901 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/X
flabel locali 10099 -13867 10133 -13833 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/X
flabel locali 10099 -13799 10133 -13765 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/X
flabel locali 10099 -13731 10133 -13697 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/X
flabel pwell 9453 -13629 9487 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/VNB
flabel nwell 9453 -14173 9487 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/VPB
flabel metal1 9453 -13629 9487 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/VGND
flabel metal1 9453 -14173 9487 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_103/VPWR
rlabel comment 9423 -13612 9423 -13612 2 sky130_fd_sc_hd__clkdlybuf4s50_1_103/clkdlybuf4s50_1
rlabel metal1 9423 -13660 10159 -13564 5 sky130_fd_sc_hd__clkdlybuf4s50_1_103/VGND
rlabel metal1 9423 -14204 10159 -14108 5 sky130_fd_sc_hd__clkdlybuf4s50_1_103/VPWR
flabel metal1 10176 -13088 10229 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_290/VPWR
flabel metal1 10179 -13630 10230 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_290/VGND
rlabel comment 10251 -13612 10251 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_290/tapvpwrvgnd_1
rlabel metal1 10159 -13660 10251 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_290/VGND
rlabel metal1 10159 -13116 10251 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_290/VPWR
flabel metal1 10181 -14165 10234 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_270/VPWR
flabel metal1 10180 -13632 10231 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_270/VGND
rlabel comment 10159 -13612 10159 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_270/tapvpwrvgnd_1
rlabel metal1 10159 -13660 10251 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_270/VGND
rlabel metal1 10159 -14204 10251 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_270/VPWR
flabel metal1 10285 -13085 10321 -13055 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_37/VPWR
flabel metal1 10285 -13625 10321 -13596 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_37/VGND
flabel nwell 10292 -13078 10312 -13061 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_37/VPB
flabel pwell 10291 -13623 10315 -13601 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_37/VNB
rlabel comment 10343 -13612 10343 -13612 6 sky130_fd_sc_hd__fill_1_37/fill_1
rlabel metal1 10251 -13660 10343 -13564 1 sky130_fd_sc_hd__fill_1_37/VGND
rlabel metal1 10251 -13116 10343 -13020 1 sky130_fd_sc_hd__fill_1_37/VPWR
flabel metal1 10648 -13629 10682 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_146/VGND
flabel metal1 10648 -13085 10682 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_146/VPWR
flabel nwell 10648 -13085 10682 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_146/VPB
flabel pwell 10648 -13629 10682 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_146/VNB
rlabel comment 10711 -13612 10711 -13612 6 sky130_fd_sc_hd__decap_4_146/decap_4
rlabel metal1 10343 -13660 10711 -13564 1 sky130_fd_sc_hd__decap_4_146/VGND
rlabel metal1 10343 -13116 10711 -13020 1 sky130_fd_sc_hd__decap_4_146/VPWR
flabel metal1 10280 -13629 10314 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_135/VGND
flabel metal1 10280 -14173 10314 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_135/VPWR
flabel nwell 10280 -14173 10314 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_135/VPB
flabel pwell 10280 -13629 10314 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_135/VNB
rlabel comment 10251 -13612 10251 -13612 2 sky130_fd_sc_hd__decap_4_135/decap_4
rlabel metal1 10251 -13660 10619 -13564 5 sky130_fd_sc_hd__decap_4_135/VGND
rlabel metal1 10251 -14204 10619 -14108 5 sky130_fd_sc_hd__decap_4_135/VPWR
flabel metal1 10641 -14165 10694 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_272/VPWR
flabel metal1 10640 -13632 10691 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_272/VGND
rlabel comment 10619 -13612 10619 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_272/tapvpwrvgnd_1
rlabel metal1 10619 -13660 10711 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_272/VGND
rlabel metal1 10619 -14204 10711 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_272/VPWR
flabel locali 11109 -13867 11143 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/Y
flabel locali 11109 -13935 11143 -13901 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/Y
flabel locali 11385 -13867 11419 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/A
flabel locali 11293 -13867 11327 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/A
flabel locali 11017 -13867 11051 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/B
flabel locali 10925 -13867 10959 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/B
flabel locali 10741 -13867 10775 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/B
flabel locali 10833 -13867 10867 -13833 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_2/B
flabel nwell 10741 -14173 10775 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_2/VPB
flabel pwell 10741 -13629 10775 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_2/VNB
flabel metal1 10741 -13629 10775 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_2/VGND
flabel metal1 10741 -14173 10775 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_2/VPWR
rlabel comment 10711 -13612 10711 -13612 2 sky130_fd_sc_hd__nand2_4_2/nand2_4
rlabel metal1 10711 -13660 11539 -13564 5 sky130_fd_sc_hd__nand2_4_2/VGND
rlabel metal1 10711 -14204 11539 -14108 5 sky130_fd_sc_hd__nand2_4_2/VPWR
flabel metal1 10653 -13085 10689 -13055 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_39/VPWR
flabel metal1 10653 -13625 10689 -13596 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_39/VGND
flabel nwell 10660 -13078 10680 -13061 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_39/VPB
flabel pwell 10659 -13623 10683 -13601 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_39/VNB
rlabel comment 10711 -13612 10711 -13612 6 sky130_fd_sc_hd__fill_1_39/fill_1
rlabel metal1 10619 -13660 10711 -13564 1 sky130_fd_sc_hd__fill_1_39/VGND
rlabel metal1 10619 -13116 10711 -13020 1 sky130_fd_sc_hd__fill_1_39/VPWR
flabel locali 11383 -13391 11417 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/A
flabel locali 10737 -13187 10771 -13153 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
flabel locali 10737 -13255 10771 -13221 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
flabel locali 10737 -13323 10771 -13289 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
flabel locali 10737 -13391 10771 -13357 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
flabel locali 10737 -13459 10771 -13425 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
flabel locali 10737 -13527 10771 -13493 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
flabel pwell 11383 -13629 11417 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/VNB
flabel nwell 11383 -13085 11417 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/VPB
flabel metal1 11383 -13629 11417 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/VGND
flabel metal1 11383 -13085 11417 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_112/VPWR
rlabel comment 11447 -13612 11447 -13612 6 sky130_fd_sc_hd__clkdlybuf4s50_1_112/clkdlybuf4s50_1
rlabel metal1 10711 -13660 11447 -13564 1 sky130_fd_sc_hd__clkdlybuf4s50_1_112/VGND
rlabel metal1 10711 -13116 11447 -13020 1 sky130_fd_sc_hd__clkdlybuf4s50_1_112/VPWR
flabel metal1 11464 -13088 11517 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_293/VPWR
flabel metal1 11467 -13630 11518 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_293/VGND
rlabel comment 11539 -13612 11539 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_293/tapvpwrvgnd_1
rlabel metal1 11447 -13660 11539 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_293/VGND
rlabel metal1 11447 -13116 11539 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_293/VPWR
flabel metal1 11561 -14165 11614 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_271/VPWR
flabel metal1 11560 -13632 11611 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_271/VGND
rlabel comment 11539 -13612 11539 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_271/tapvpwrvgnd_1
rlabel metal1 11539 -13660 11631 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_271/VGND
rlabel metal1 11539 -14204 11631 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_271/VPWR
flabel metal1 12668 -13632 12700 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_21/VGND
flabel metal1 12668 -13089 12706 -13057 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_21/VPWR
flabel nwell 12658 -13090 12715 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_21/VPB
flabel pwell 12665 -13636 12709 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_21/VNB
rlabel comment 12735 -13612 12735 -13612 6 sky130_fd_sc_hd__fill_8_21/fill_8
rlabel metal1 11999 -13660 12735 -13564 1 sky130_fd_sc_hd__fill_8_21/VGND
rlabel metal1 11999 -13116 12735 -13020 1 sky130_fd_sc_hd__fill_8_21/VPWR
flabel metal1 12034 -13622 12066 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_19/VGND
flabel metal1 12028 -14167 12066 -14135 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_19/VPWR
flabel nwell 12019 -14165 12076 -14134 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_19/VPB
flabel pwell 12025 -13622 12069 -13588 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_19/VNB
rlabel comment 11999 -13612 11999 -13612 2 sky130_fd_sc_hd__fill_8_19/fill_8
rlabel metal1 11999 -13660 12735 -13564 5 sky130_fd_sc_hd__fill_8_19/VGND
rlabel metal1 11999 -14204 12735 -14108 5 sky130_fd_sc_hd__fill_8_19/VPWR
flabel metal1 11573 -13085 11609 -13055 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_38/VPWR
flabel metal1 11573 -13625 11609 -13596 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_38/VGND
flabel nwell 11580 -13078 11600 -13061 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_38/VPB
flabel pwell 11579 -13623 11603 -13601 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_38/VNB
rlabel comment 11631 -13612 11631 -13612 6 sky130_fd_sc_hd__fill_1_38/fill_1
rlabel metal1 11539 -13660 11631 -13564 1 sky130_fd_sc_hd__fill_1_38/VGND
rlabel metal1 11539 -13116 11631 -13020 1 sky130_fd_sc_hd__fill_1_38/VPWR
flabel metal1 11936 -13629 11970 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_145/VGND
flabel metal1 11936 -13085 11970 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_145/VPWR
flabel nwell 11936 -13085 11970 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_145/VPB
flabel pwell 11936 -13629 11970 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_145/VNB
rlabel comment 11999 -13612 11999 -13612 6 sky130_fd_sc_hd__decap_4_145/decap_4
rlabel metal1 11631 -13660 11999 -13564 1 sky130_fd_sc_hd__decap_4_145/VGND
rlabel metal1 11631 -13116 11999 -13020 1 sky130_fd_sc_hd__decap_4_145/VPWR
flabel metal1 11660 -13629 11694 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_136/VGND
flabel metal1 11660 -14173 11694 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_136/VPWR
flabel nwell 11660 -14173 11694 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_136/VPB
flabel pwell 11660 -13629 11694 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_136/VNB
rlabel comment 11631 -13612 11631 -13612 2 sky130_fd_sc_hd__decap_4_136/decap_4
rlabel metal1 11631 -13660 11999 -13564 5 sky130_fd_sc_hd__decap_4_136/VGND
rlabel metal1 11631 -14204 11999 -14108 5 sky130_fd_sc_hd__decap_4_136/VPWR
flabel locali 15248 -13323 15282 -13289 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/X
flabel locali 15340 -13323 15374 -13289 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/X
flabel locali 15340 -13391 15374 -13357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/X
flabel locali 15248 -13391 15282 -13357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/X
flabel locali 15248 -13459 15282 -13425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/X
flabel locali 15340 -13459 15374 -13425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/X
flabel locali 13684 -13459 13718 -13425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/A
flabel locali 13684 -13391 13718 -13357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/A
flabel pwell 13684 -13629 13718 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/VNB
flabel pwell 13701 -13612 13701 -13612 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/VNB
flabel nwell 13684 -13085 13718 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/VPB
flabel nwell 13701 -13068 13701 -13068 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/VPB
flabel metal1 13684 -13629 13718 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/VGND
flabel metal1 13684 -13085 13718 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_8/VPWR
rlabel comment 13655 -13612 13655 -13612 4 sky130_fd_sc_hd__clkbuf_16_8/clkbuf_16
rlabel metal1 13655 -13660 15495 -13564 1 sky130_fd_sc_hd__clkbuf_16_8/VGND
rlabel metal1 13655 -13116 15495 -13020 1 sky130_fd_sc_hd__clkbuf_16_8/VPWR
flabel metal1 13592 -13629 13626 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_19/VGND
flabel metal1 13592 -14173 13626 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_19/VPWR
flabel nwell 13592 -14173 13626 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_19/VPB
flabel pwell 13592 -13629 13626 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_19/VNB
rlabel comment 13563 -13612 13563 -13612 2 sky130_fd_sc_hd__decap_12_19/decap_12
rlabel metal1 13563 -13660 14667 -13564 5 sky130_fd_sc_hd__decap_12_19/VGND
rlabel metal1 13563 -14204 14667 -14108 5 sky130_fd_sc_hd__decap_12_19/VPWR
flabel metal1 13505 -13085 13541 -13055 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_40/VPWR
flabel metal1 13505 -13625 13541 -13596 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_40/VGND
flabel nwell 13512 -13078 13532 -13061 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_40/VPB
flabel pwell 13511 -13623 13535 -13601 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_40/VNB
rlabel comment 13563 -13612 13563 -13612 6 sky130_fd_sc_hd__fill_1_40/fill_1
rlabel metal1 13471 -13660 13563 -13564 1 sky130_fd_sc_hd__fill_1_40/VGND
rlabel metal1 13471 -13116 13563 -13020 1 sky130_fd_sc_hd__fill_1_40/VPWR
flabel metal1 12770 -13622 12802 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_20/VGND
flabel metal1 12764 -14167 12802 -14135 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_20/VPWR
flabel nwell 12755 -14165 12812 -14134 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_20/VPB
flabel pwell 12761 -13622 12805 -13588 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_20/VNB
rlabel comment 12735 -13612 12735 -13612 2 sky130_fd_sc_hd__fill_8_20/fill_8
rlabel metal1 12735 -13660 13471 -13564 5 sky130_fd_sc_hd__fill_8_20/VGND
rlabel metal1 12735 -14204 13471 -14108 5 sky130_fd_sc_hd__fill_8_20/VPWR
flabel metal1 13404 -13632 13436 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_22/VGND
flabel metal1 13404 -13089 13442 -13057 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_22/VPWR
flabel nwell 13394 -13090 13451 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_22/VPB
flabel pwell 13401 -13636 13445 -13602 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_22/VNB
rlabel comment 13471 -13612 13471 -13612 6 sky130_fd_sc_hd__fill_8_22/fill_8
rlabel metal1 12735 -13660 13471 -13564 1 sky130_fd_sc_hd__fill_8_22/VGND
rlabel metal1 12735 -13116 13471 -13020 1 sky130_fd_sc_hd__fill_8_22/VPWR
flabel metal1 13493 -14165 13546 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_273/VPWR
flabel metal1 13492 -13632 13543 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_273/VGND
rlabel comment 13471 -13612 13471 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_273/tapvpwrvgnd_1
rlabel metal1 13471 -13660 13563 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_273/VGND
rlabel metal1 13471 -14204 13563 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_273/VPWR
flabel metal1 13580 -13088 13633 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_294/VPWR
flabel metal1 13583 -13630 13634 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_294/VGND
rlabel comment 13655 -13612 13655 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_294/tapvpwrvgnd_1
rlabel metal1 13563 -13660 13655 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_294/VGND
rlabel metal1 13563 -13116 13655 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_294/VPWR
flabel metal1 15984 -14173 16018 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_22/VPWR
flabel metal1 15984 -13629 16018 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_22/VGND
flabel nwell 15984 -14173 16018 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_22/VPB
flabel pwell 15984 -13629 16018 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_22/VNB
rlabel comment 15955 -13612 15955 -13612 2 sky130_fd_sc_hd__decap_8_22/decap_8
rlabel metal1 15955 -13660 16691 -13564 5 sky130_fd_sc_hd__decap_8_22/VGND
rlabel metal1 15955 -14204 16691 -14108 5 sky130_fd_sc_hd__decap_8_22/VPWR
flabel metal1 14788 -13629 14822 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_20/VGND
flabel metal1 14788 -14173 14822 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_20/VPWR
flabel nwell 14788 -14173 14822 -14139 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_20/VPB
flabel pwell 14788 -13629 14822 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_20/VNB
rlabel comment 14759 -13612 14759 -13612 2 sky130_fd_sc_hd__decap_12_20/decap_12
rlabel metal1 14759 -13660 15863 -13564 5 sky130_fd_sc_hd__decap_12_20/VGND
rlabel metal1 14759 -14204 15863 -14108 5 sky130_fd_sc_hd__decap_12_20/VPWR
flabel metal1 16628 -13629 16662 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_21/VGND
flabel metal1 16628 -13085 16662 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_21/VPWR
flabel nwell 16628 -13085 16662 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_21/VPB
flabel pwell 16628 -13629 16662 -13595 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_21/VNB
rlabel comment 16691 -13612 16691 -13612 6 sky130_fd_sc_hd__decap_12_21/decap_12
rlabel metal1 15587 -13660 16691 -13564 1 sky130_fd_sc_hd__decap_12_21/VGND
rlabel metal1 15587 -13116 16691 -13020 1 sky130_fd_sc_hd__decap_12_21/VPWR
flabel metal1 14689 -14165 14742 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_274/VPWR
flabel metal1 14688 -13632 14739 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_274/VGND
rlabel comment 14667 -13612 14667 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_274/tapvpwrvgnd_1
rlabel metal1 14667 -13660 14759 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_274/VGND
rlabel metal1 14667 -14204 14759 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_274/VPWR
flabel metal1 15885 -14165 15938 -14136 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_275/VPWR
flabel metal1 15884 -13632 15935 -13594 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_275/VGND
rlabel comment 15863 -13612 15863 -13612 2 sky130_fd_sc_hd__tapvpwrvgnd_1_275/tapvpwrvgnd_1
rlabel metal1 15863 -13660 15955 -13564 5 sky130_fd_sc_hd__tapvpwrvgnd_1_275/VGND
rlabel metal1 15863 -14204 15955 -14108 5 sky130_fd_sc_hd__tapvpwrvgnd_1_275/VPWR
flabel metal1 15512 -13088 15565 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_295/VPWR
flabel metal1 15515 -13630 15566 -13592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_295/VGND
rlabel comment 15587 -13612 15587 -13612 6 sky130_fd_sc_hd__tapvpwrvgnd_1_295/tapvpwrvgnd_1
rlabel metal1 15495 -13660 15587 -13564 1 sky130_fd_sc_hd__tapvpwrvgnd_1_295/VGND
rlabel metal1 15495 -13116 15587 -13020 1 sky130_fd_sc_hd__tapvpwrvgnd_1_295/VPWR
flabel metal1 -1588 -13085 -1554 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_25/VPWR
flabel metal1 -1588 -12541 -1554 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_25/VGND
flabel nwell -1588 -13085 -1554 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_25/VPB
flabel pwell -1588 -12541 -1554 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_25/VNB
rlabel comment -1617 -12524 -1617 -12524 2 sky130_fd_sc_hd__decap_8_25/decap_8
rlabel metal1 -1617 -12572 -881 -12476 5 sky130_fd_sc_hd__decap_8_25/VGND
rlabel metal1 -1617 -13116 -881 -13020 5 sky130_fd_sc_hd__decap_8_25/VPWR
flabel metal1 -2324 -13085 -2290 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_88/VPWR
flabel metal1 -2324 -12541 -2290 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_88/VGND
flabel nwell -2324 -13085 -2290 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_88/VPB
flabel pwell -2324 -12541 -2290 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_88/VNB
rlabel comment -2261 -12524 -2261 -12524 8 sky130_fd_sc_hd__decap_8_88/decap_8
rlabel metal1 -2997 -12572 -2261 -12476 5 sky130_fd_sc_hd__decap_8_88/VGND
rlabel metal1 -2997 -13116 -2261 -13020 5 sky130_fd_sc_hd__decap_8_88/VPWR
flabel metal1 -1690 -12542 -1637 -12510 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_27/VGND
flabel metal1 -1690 -13085 -1638 -13054 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_27/VPWR
flabel nwell -1679 -13077 -1645 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_27/VPB
flabel pwell -1680 -12536 -1648 -12514 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_27/VNB
rlabel comment -1617 -12524 -1617 -12524 8 sky130_fd_sc_hd__fill_2_27/fill_2
rlabel metal1 -1801 -12572 -1617 -12476 5 sky130_fd_sc_hd__fill_2_27/VGND
rlabel metal1 -1801 -13116 -1617 -13020 5 sky130_fd_sc_hd__fill_2_27/VPWR
flabel metal1 -1858 -12533 -1835 -12514 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_35/VGND
flabel metal1 -1855 -13076 -1835 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_35/VPWR
flabel nwell -1861 -13080 -1836 -13054 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_35/VPB
flabel pwell -1858 -12536 -1836 -12512 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_35/VNB
rlabel comment -1801 -12524 -1801 -12524 8 sky130_fd_sc_hd__fill_4_35/fill_4
rlabel metal1 -2169 -12572 -1801 -12476 5 sky130_fd_sc_hd__fill_4_35/VGND
rlabel metal1 -2169 -13116 -1801 -13020 5 sky130_fd_sc_hd__fill_4_35/VPWR
flabel metal1 -2244 -13077 -2191 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_553/VPWR
flabel metal1 -2241 -12544 -2190 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_553/VGND
rlabel comment -2169 -12524 -2169 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_553/tapvpwrvgnd_1
rlabel metal1 -2261 -12572 -2169 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_553/VGND
rlabel metal1 -2261 -13116 -2169 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_553/VPWR
flabel locali 437 -12779 471 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A
flabel locali 1083 -12983 1117 -12949 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/X
flabel locali 1083 -12915 1117 -12881 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/X
flabel locali 1083 -12847 1117 -12813 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/X
flabel locali 1083 -12779 1117 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/X
flabel locali 1083 -12711 1117 -12677 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/X
flabel locali 1083 -12643 1117 -12609 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/X
flabel pwell 437 -12541 471 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/VNB
flabel nwell 437 -13085 471 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/VPB
flabel metal1 437 -12541 471 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/VGND
flabel metal1 437 -13085 471 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_113/VPWR
rlabel comment 407 -12524 407 -12524 2 sky130_fd_sc_hd__clkdlybuf4s50_1_113/clkdlybuf4s50_1
rlabel metal1 407 -12572 1143 -12476 5 sky130_fd_sc_hd__clkdlybuf4s50_1_113/VGND
rlabel metal1 407 -13116 1143 -13020 5 sky130_fd_sc_hd__clkdlybuf4s50_1_113/VPWR
flabel metal1 252 -12541 286 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_147/VGND
flabel metal1 252 -13085 286 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_147/VPWR
flabel nwell 252 -13085 286 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_147/VPB
flabel pwell 252 -12541 286 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_147/VNB
rlabel comment 315 -12524 315 -12524 8 sky130_fd_sc_hd__decap_4_147/decap_4
rlabel metal1 -53 -12572 315 -12476 5 sky130_fd_sc_hd__decap_4_147/VGND
rlabel metal1 -53 -13116 315 -13020 5 sky130_fd_sc_hd__decap_4_147/VPWR
flabel metal1 -852 -13085 -818 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_26/VPWR
flabel metal1 -852 -12541 -818 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_26/VGND
flabel nwell -852 -13085 -818 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_26/VPB
flabel pwell -852 -12541 -818 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_26/VNB
rlabel comment -881 -12524 -881 -12524 2 sky130_fd_sc_hd__decap_8_26/decap_8
rlabel metal1 -881 -12572 -145 -12476 5 sky130_fd_sc_hd__decap_8_26/VGND
rlabel metal1 -881 -13116 -145 -13020 5 sky130_fd_sc_hd__decap_8_26/VPWR
flabel metal1 332 -13077 385 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_296/VPWR
flabel metal1 335 -12544 386 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_296/VGND
rlabel comment 407 -12524 407 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_296/tapvpwrvgnd_1
rlabel metal1 315 -12572 407 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_296/VGND
rlabel metal1 315 -13116 407 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_296/VPWR
flabel metal1 -128 -13077 -75 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_297/VPWR
flabel metal1 -125 -12544 -74 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_297/VGND
rlabel comment -53 -12524 -53 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_297/tapvpwrvgnd_1
rlabel metal1 -145 -12572 -53 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_297/VGND
rlabel metal1 -145 -13116 -53 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_297/VPWR
flabel metal1 2828 -12541 2862 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_148/VGND
flabel metal1 2828 -13085 2862 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_148/VPWR
flabel nwell 2828 -13085 2862 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_148/VPB
flabel pwell 2828 -12541 2862 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_148/VNB
rlabel comment 2891 -12524 2891 -12524 8 sky130_fd_sc_hd__decap_4_148/decap_4
rlabel metal1 2523 -12572 2891 -12476 5 sky130_fd_sc_hd__decap_4_148/VGND
rlabel metal1 2523 -13116 2891 -13020 5 sky130_fd_sc_hd__decap_4_148/VPWR
flabel metal1 1540 -12541 1574 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_149/VGND
flabel metal1 1540 -13085 1574 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_149/VPWR
flabel nwell 1540 -13085 1574 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_149/VPB
flabel pwell 1540 -12541 1574 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_149/VNB
rlabel comment 1603 -12524 1603 -12524 8 sky130_fd_sc_hd__decap_4_149/decap_4
rlabel metal1 1235 -12572 1603 -12476 5 sky130_fd_sc_hd__decap_4_149/VGND
rlabel metal1 1235 -13116 1603 -13020 5 sky130_fd_sc_hd__decap_4_149/VPWR
flabel metal1 2368 -13085 2402 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_139/VPWR
flabel metal1 2368 -12541 2402 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_139/VGND
flabel nwell 2368 -13085 2402 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_139/VPB
flabel pwell 2368 -12541 2402 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_139/VNB
rlabel comment 2431 -12524 2431 -12524 8 sky130_fd_sc_hd__decap_8_139/decap_8
rlabel metal1 1695 -12572 2431 -12476 5 sky130_fd_sc_hd__decap_8_139/VGND
rlabel metal1 1695 -13116 2431 -13020 5 sky130_fd_sc_hd__decap_8_139/VPWR
flabel metal1 2448 -13077 2501 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_298/VPWR
flabel metal1 2451 -12544 2502 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_298/VGND
rlabel comment 2523 -12524 2523 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_298/tapvpwrvgnd_1
rlabel metal1 2431 -12572 2523 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_298/VGND
rlabel metal1 2431 -13116 2523 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_298/VPWR
flabel metal1 1620 -13077 1673 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_299/VPWR
flabel metal1 1623 -12544 1674 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_299/VGND
rlabel comment 1695 -12524 1695 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_299/tapvpwrvgnd_1
rlabel metal1 1603 -12572 1695 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_299/VGND
rlabel metal1 1603 -13116 1695 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_299/VPWR
flabel metal1 1160 -13077 1213 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_300/VPWR
flabel metal1 1163 -12544 1214 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_300/VGND
rlabel comment 1235 -12524 1235 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_300/tapvpwrvgnd_1
rlabel metal1 1143 -12572 1235 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_300/VGND
rlabel metal1 1143 -13116 1235 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_300/VPWR
flabel locali 3013 -12779 3047 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A
flabel locali 3659 -12983 3693 -12949 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X
flabel locali 3659 -12915 3693 -12881 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X
flabel locali 3659 -12847 3693 -12813 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X
flabel locali 3659 -12779 3693 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X
flabel locali 3659 -12711 3693 -12677 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X
flabel locali 3659 -12643 3693 -12609 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X
flabel pwell 3013 -12541 3047 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/VNB
flabel nwell 3013 -13085 3047 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/VPB
flabel metal1 3013 -12541 3047 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/VGND
flabel metal1 3013 -13085 3047 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_116/VPWR
rlabel comment 2983 -12524 2983 -12524 2 sky130_fd_sc_hd__clkdlybuf4s50_1_116/clkdlybuf4s50_1
rlabel metal1 2983 -12572 3719 -12476 5 sky130_fd_sc_hd__clkdlybuf4s50_1_116/VGND
rlabel metal1 2983 -13116 3719 -13020 5 sky130_fd_sc_hd__clkdlybuf4s50_1_116/VPWR
flabel metal1 4116 -12541 4150 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_150/VGND
flabel metal1 4116 -13085 4150 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_150/VPWR
flabel nwell 4116 -13085 4150 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_150/VPB
flabel pwell 4116 -12541 4150 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_150/VNB
rlabel comment 4179 -12524 4179 -12524 8 sky130_fd_sc_hd__decap_4_150/decap_4
rlabel metal1 3811 -12572 4179 -12476 5 sky130_fd_sc_hd__decap_4_150/VGND
rlabel metal1 3811 -13116 4179 -13020 5 sky130_fd_sc_hd__decap_4_150/VPWR
flabel metal1 4944 -13085 4978 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_141/VPWR
flabel metal1 4944 -12541 4978 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_141/VGND
flabel nwell 4944 -13085 4978 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_141/VPB
flabel pwell 4944 -12541 4978 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_141/VNB
rlabel comment 5007 -12524 5007 -12524 8 sky130_fd_sc_hd__decap_8_141/decap_8
rlabel metal1 4271 -12572 5007 -12476 5 sky130_fd_sc_hd__decap_8_141/VGND
rlabel metal1 4271 -13116 5007 -13020 5 sky130_fd_sc_hd__decap_8_141/VPWR
flabel metal1 3736 -13077 3789 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_301/VPWR
flabel metal1 3739 -12544 3790 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_301/VGND
rlabel comment 3811 -12524 3811 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_301/tapvpwrvgnd_1
rlabel metal1 3719 -12572 3811 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_301/VGND
rlabel metal1 3719 -13116 3811 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_301/VPWR
flabel metal1 4196 -13077 4249 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_302/VPWR
flabel metal1 4199 -12544 4250 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_302/VGND
rlabel comment 4271 -12524 4271 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_302/tapvpwrvgnd_1
rlabel metal1 4179 -12572 4271 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_302/VGND
rlabel metal1 4179 -13116 4271 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_302/VPWR
flabel metal1 2908 -13077 2961 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_303/VPWR
flabel metal1 2911 -12544 2962 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_303/VGND
rlabel comment 2983 -12524 2983 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_303/tapvpwrvgnd_1
rlabel metal1 2891 -12572 2983 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_303/VGND
rlabel metal1 2891 -13116 2983 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_303/VPWR
flabel locali 5589 -12779 5623 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A
flabel locali 6235 -12983 6269 -12949 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/X
flabel locali 6235 -12915 6269 -12881 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/X
flabel locali 6235 -12847 6269 -12813 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/X
flabel locali 6235 -12779 6269 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/X
flabel locali 6235 -12711 6269 -12677 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/X
flabel locali 6235 -12643 6269 -12609 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/X
flabel pwell 5589 -12541 5623 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/VNB
flabel nwell 5589 -13085 5623 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/VPB
flabel metal1 5589 -12541 5623 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/VGND
flabel metal1 5589 -13085 5623 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_117/VPWR
rlabel comment 5559 -12524 5559 -12524 2 sky130_fd_sc_hd__clkdlybuf4s50_1_117/clkdlybuf4s50_1
rlabel metal1 5559 -12572 6295 -12476 5 sky130_fd_sc_hd__clkdlybuf4s50_1_117/VGND
rlabel metal1 5559 -13116 6295 -13020 5 sky130_fd_sc_hd__clkdlybuf4s50_1_117/VPWR
flabel metal1 6692 -12541 6726 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_151/VGND
flabel metal1 6692 -13085 6726 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_151/VPWR
flabel nwell 6692 -13085 6726 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_151/VPB
flabel pwell 6692 -12541 6726 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_151/VNB
rlabel comment 6755 -12524 6755 -12524 8 sky130_fd_sc_hd__decap_4_151/decap_4
rlabel metal1 6387 -12572 6755 -12476 5 sky130_fd_sc_hd__decap_4_151/VGND
rlabel metal1 6387 -13116 6755 -13020 5 sky130_fd_sc_hd__decap_4_151/VPWR
flabel metal1 5404 -12541 5438 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_152/VGND
flabel metal1 5404 -13085 5438 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_152/VPWR
flabel nwell 5404 -13085 5438 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_152/VPB
flabel pwell 5404 -12541 5438 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_152/VNB
rlabel comment 5467 -12524 5467 -12524 8 sky130_fd_sc_hd__decap_4_152/decap_4
rlabel metal1 5099 -12572 5467 -12476 5 sky130_fd_sc_hd__decap_4_152/VGND
rlabel metal1 5099 -13116 5467 -13020 5 sky130_fd_sc_hd__decap_4_152/VPWR
flabel metal1 6312 -13077 6365 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_304/VPWR
flabel metal1 6315 -12544 6366 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_304/VGND
rlabel comment 6387 -12524 6387 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_304/tapvpwrvgnd_1
rlabel metal1 6295 -12572 6387 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_304/VGND
rlabel metal1 6295 -13116 6387 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_304/VPWR
flabel metal1 5484 -13077 5537 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_305/VPWR
flabel metal1 5487 -12544 5538 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_305/VGND
rlabel comment 5559 -12524 5559 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_305/tapvpwrvgnd_1
rlabel metal1 5467 -12572 5559 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_305/VGND
rlabel metal1 5467 -13116 5559 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_305/VPWR
flabel metal1 5024 -13077 5077 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_306/VPWR
flabel metal1 5027 -12544 5078 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_306/VGND
rlabel comment 5099 -12524 5099 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_306/tapvpwrvgnd_1
rlabel metal1 5007 -12572 5099 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_306/VGND
rlabel metal1 5007 -13116 5099 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_306/VPWR
flabel locali 8165 -12779 8199 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A
flabel locali 8811 -12983 8845 -12949 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/X
flabel locali 8811 -12915 8845 -12881 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/X
flabel locali 8811 -12847 8845 -12813 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/X
flabel locali 8811 -12779 8845 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/X
flabel locali 8811 -12711 8845 -12677 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/X
flabel locali 8811 -12643 8845 -12609 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/X
flabel pwell 8165 -12541 8199 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/VNB
flabel nwell 8165 -13085 8199 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/VPB
flabel metal1 8165 -12541 8199 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/VGND
flabel metal1 8165 -13085 8199 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_118/VPWR
rlabel comment 8135 -12524 8135 -12524 2 sky130_fd_sc_hd__clkdlybuf4s50_1_118/clkdlybuf4s50_1
rlabel metal1 8135 -12572 8871 -12476 5 sky130_fd_sc_hd__clkdlybuf4s50_1_118/VGND
rlabel metal1 8135 -13116 8871 -13020 5 sky130_fd_sc_hd__clkdlybuf4s50_1_118/VPWR
flabel metal1 7980 -12541 8014 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_153/VGND
flabel metal1 7980 -13085 8014 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_153/VPWR
flabel nwell 7980 -13085 8014 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_153/VPB
flabel pwell 7980 -12541 8014 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_153/VNB
rlabel comment 8043 -12524 8043 -12524 8 sky130_fd_sc_hd__decap_4_153/decap_4
rlabel metal1 7675 -12572 8043 -12476 5 sky130_fd_sc_hd__decap_4_153/VGND
rlabel metal1 7675 -13116 8043 -13020 5 sky130_fd_sc_hd__decap_4_153/VPWR
flabel metal1 7520 -13085 7554 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_151/VPWR
flabel metal1 7520 -12541 7554 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_151/VGND
flabel nwell 7520 -13085 7554 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_151/VPB
flabel pwell 7520 -12541 7554 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_151/VNB
rlabel comment 7583 -12524 7583 -12524 8 sky130_fd_sc_hd__decap_8_151/decap_8
rlabel metal1 6847 -12572 7583 -12476 5 sky130_fd_sc_hd__decap_8_151/VGND
rlabel metal1 6847 -13116 7583 -13020 5 sky130_fd_sc_hd__decap_8_151/VPWR
flabel metal1 7600 -13077 7653 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_307/VPWR
flabel metal1 7603 -12544 7654 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_307/VGND
rlabel comment 7675 -12524 7675 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_307/tapvpwrvgnd_1
rlabel metal1 7583 -12572 7675 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_307/VGND
rlabel metal1 7583 -13116 7675 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_307/VPWR
flabel metal1 8060 -13077 8113 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_308/VPWR
flabel metal1 8063 -12544 8114 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_308/VGND
rlabel comment 8135 -12524 8135 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_308/tapvpwrvgnd_1
rlabel metal1 8043 -12572 8135 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_308/VGND
rlabel metal1 8043 -13116 8135 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_308/VPWR
flabel metal1 6772 -13077 6825 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_309/VPWR
flabel metal1 6775 -12544 6826 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_309/VGND
rlabel comment 6847 -12524 6847 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_309/tapvpwrvgnd_1
rlabel metal1 6755 -12572 6847 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_309/VGND
rlabel metal1 6755 -13116 6847 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_309/VPWR
flabel metal1 9268 -12541 9302 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_154/VGND
flabel metal1 9268 -13085 9302 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_154/VPWR
flabel nwell 9268 -13085 9302 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_154/VPB
flabel pwell 9268 -12541 9302 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_154/VNB
rlabel comment 9331 -12524 9331 -12524 8 sky130_fd_sc_hd__decap_4_154/decap_4
rlabel metal1 8963 -12572 9331 -12476 5 sky130_fd_sc_hd__decap_4_154/VGND
rlabel metal1 8963 -13116 9331 -13020 5 sky130_fd_sc_hd__decap_4_154/VPWR
flabel metal1 10648 -12541 10682 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_156/VGND
flabel metal1 10648 -13085 10682 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_156/VPWR
flabel nwell 10648 -13085 10682 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_156/VPB
flabel pwell 10648 -12541 10682 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_156/VNB
rlabel comment 10711 -12524 10711 -12524 8 sky130_fd_sc_hd__decap_4_156/decap_4
rlabel metal1 10343 -12572 10711 -12476 5 sky130_fd_sc_hd__decap_4_156/VGND
rlabel metal1 10343 -13116 10711 -13020 5 sky130_fd_sc_hd__decap_4_156/VPWR
flabel metal1 10096 -13085 10130 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_162/VPWR
flabel metal1 10096 -12541 10130 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_162/VGND
flabel nwell 10096 -13085 10130 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_162/VPB
flabel pwell 10096 -12541 10130 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_162/VNB
rlabel comment 10159 -12524 10159 -12524 8 sky130_fd_sc_hd__decap_8_162/decap_8
rlabel metal1 9423 -12572 10159 -12476 5 sky130_fd_sc_hd__decap_8_162/VGND
rlabel metal1 9423 -13116 10159 -13020 5 sky130_fd_sc_hd__decap_8_162/VPWR
flabel metal1 10285 -13081 10321 -13051 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_41/VPWR
flabel metal1 10285 -12540 10321 -12511 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_41/VGND
flabel nwell 10292 -13075 10312 -13058 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_41/VPB
flabel pwell 10291 -12535 10315 -12513 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_41/VNB
rlabel comment 10343 -12524 10343 -12524 8 sky130_fd_sc_hd__fill_1_41/fill_1
rlabel metal1 10251 -12572 10343 -12476 5 sky130_fd_sc_hd__fill_1_41/VGND
rlabel metal1 10251 -13116 10343 -13020 5 sky130_fd_sc_hd__fill_1_41/VPWR
flabel metal1 10176 -13077 10229 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_310/VPWR
flabel metal1 10179 -12544 10230 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_310/VGND
rlabel comment 10251 -12524 10251 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_310/tapvpwrvgnd_1
rlabel metal1 10159 -12572 10251 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_310/VGND
rlabel metal1 10159 -13116 10251 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_310/VPWR
flabel metal1 9348 -13077 9401 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_311/VPWR
flabel metal1 9351 -12544 9402 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_311/VGND
rlabel comment 9423 -12524 9423 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_311/tapvpwrvgnd_1
rlabel metal1 9331 -12572 9423 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_311/VGND
rlabel metal1 9331 -13116 9423 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_311/VPWR
flabel metal1 8888 -13077 8941 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_312/VPWR
flabel metal1 8891 -12544 8942 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_312/VGND
rlabel comment 8963 -12524 8963 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_312/tapvpwrvgnd_1
rlabel metal1 8871 -12572 8963 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_312/VGND
rlabel metal1 8871 -13116 8963 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_312/VPWR
flabel locali 10741 -12779 10775 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A
flabel locali 11387 -12983 11421 -12949 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/X
flabel locali 11387 -12915 11421 -12881 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/X
flabel locali 11387 -12847 11421 -12813 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/X
flabel locali 11387 -12779 11421 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/X
flabel locali 11387 -12711 11421 -12677 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/X
flabel locali 11387 -12643 11421 -12609 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/X
flabel pwell 10741 -12541 10775 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/VNB
flabel nwell 10741 -13085 10775 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/VPB
flabel metal1 10741 -12541 10775 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/VGND
flabel metal1 10741 -13085 10775 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_121/VPWR
rlabel comment 10711 -12524 10711 -12524 2 sky130_fd_sc_hd__clkdlybuf4s50_1_121/clkdlybuf4s50_1
rlabel metal1 10711 -12572 11447 -12476 5 sky130_fd_sc_hd__clkdlybuf4s50_1_121/VGND
rlabel metal1 10711 -13116 11447 -13020 5 sky130_fd_sc_hd__clkdlybuf4s50_1_121/VPWR
flabel metal1 11936 -12541 11970 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_155/VGND
flabel metal1 11936 -13085 11970 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_155/VPWR
flabel nwell 11936 -13085 11970 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_155/VPB
flabel pwell 11936 -12541 11970 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_155/VNB
rlabel comment 11999 -12524 11999 -12524 8 sky130_fd_sc_hd__decap_4_155/decap_4
rlabel metal1 11631 -12572 11999 -12476 5 sky130_fd_sc_hd__decap_4_155/VGND
rlabel metal1 11631 -13116 11999 -13020 5 sky130_fd_sc_hd__decap_4_155/VPWR
flabel metal1 11573 -13081 11609 -13051 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_42/VPWR
flabel metal1 11573 -12540 11609 -12511 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_42/VGND
flabel nwell 11580 -13075 11600 -13058 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_42/VPB
flabel pwell 11579 -12535 11603 -12513 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_42/VNB
rlabel comment 11631 -12524 11631 -12524 8 sky130_fd_sc_hd__fill_1_42/fill_1
rlabel metal1 11539 -12572 11631 -12476 5 sky130_fd_sc_hd__fill_1_42/VGND
rlabel metal1 11539 -13116 11631 -13020 5 sky130_fd_sc_hd__fill_1_42/VPWR
flabel metal1 10653 -13081 10689 -13051 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_43/VPWR
flabel metal1 10653 -12540 10689 -12511 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_43/VGND
flabel nwell 10660 -13075 10680 -13058 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_43/VPB
flabel pwell 10659 -12535 10683 -12513 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_43/VNB
rlabel comment 10711 -12524 10711 -12524 8 sky130_fd_sc_hd__fill_1_43/fill_1
rlabel metal1 10619 -12572 10711 -12476 5 sky130_fd_sc_hd__fill_1_43/VGND
rlabel metal1 10619 -13116 10711 -13020 5 sky130_fd_sc_hd__fill_1_43/VPWR
flabel metal1 12033 -12533 12056 -12514 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_10/VGND
flabel metal1 12033 -13076 12053 -13059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_10/VPWR
flabel nwell 12034 -13080 12059 -13054 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_10/VPB
flabel pwell 12034 -12536 12056 -12512 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_10/VNB
rlabel comment 11999 -12524 11999 -12524 2 sky130_fd_sc_hd__fill_4_10/fill_4
rlabel metal1 11999 -12572 12367 -12476 5 sky130_fd_sc_hd__fill_4_10/VGND
rlabel metal1 11999 -13116 12367 -13020 5 sky130_fd_sc_hd__fill_4_10/VPWR
flabel metal1 11464 -13077 11517 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_313/VPWR
flabel metal1 11467 -12544 11518 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_313/VGND
rlabel comment 11539 -12524 11539 -12524 8 sky130_fd_sc_hd__tapvpwrvgnd_1_313/tapvpwrvgnd_1
rlabel metal1 11447 -12572 11539 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_313/VGND
rlabel metal1 11447 -13116 11539 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_313/VPWR
flabel locali 15248 -12847 15282 -12813 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/X
flabel locali 15340 -12847 15374 -12813 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/X
flabel locali 15340 -12779 15374 -12745 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/X
flabel locali 15248 -12779 15282 -12745 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/X
flabel locali 15248 -12711 15282 -12677 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/X
flabel locali 15340 -12711 15374 -12677 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/X
flabel locali 13684 -12711 13718 -12677 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/A
flabel locali 13684 -12779 13718 -12745 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/A
flabel pwell 13684 -12541 13718 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/VNB
flabel pwell 13701 -12524 13701 -12524 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/VNB
flabel nwell 13684 -13085 13718 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/VPB
flabel nwell 13701 -13068 13701 -13068 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/VPB
flabel metal1 13684 -12541 13718 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/VGND
flabel metal1 13684 -13085 13718 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_9/VPWR
rlabel comment 13655 -12524 13655 -12524 2 sky130_fd_sc_hd__clkbuf_16_9/clkbuf_16
rlabel metal1 13655 -12572 15495 -12476 5 sky130_fd_sc_hd__clkbuf_16_9/VGND
rlabel metal1 13655 -13116 15495 -13020 5 sky130_fd_sc_hd__clkbuf_16_9/VPWR
flabel locali 12672 -12779 12706 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/A
flabel locali 12764 -12779 12798 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/A
flabel locali 13040 -12711 13074 -12677 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/Y
flabel locali 12580 -12779 12614 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/A
flabel locali 13040 -12847 13074 -12813 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/Y
flabel locali 12948 -12779 12982 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/A
flabel locali 12856 -12779 12890 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/A
flabel locali 13040 -12779 13074 -12745 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_7/Y
flabel pwell 12488 -12541 12522 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_7/VNB
flabel nwell 12488 -13085 12522 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_7/VPB
flabel metal1 12488 -13085 12522 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_7/VPWR
flabel metal1 12488 -12541 12522 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_7/VGND
rlabel comment 12459 -12524 12459 -12524 2 sky130_fd_sc_hd__clkinv_4_7/clkinv_4
rlabel metal1 12459 -12572 13103 -12476 5 sky130_fd_sc_hd__clkinv_4_7/VGND
rlabel metal1 12459 -13116 13103 -13020 5 sky130_fd_sc_hd__clkinv_4_7/VPWR
flabel metal1 13224 -12541 13258 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_157/VGND
flabel metal1 13224 -13085 13258 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_157/VPWR
flabel nwell 13224 -13085 13258 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_157/VPB
flabel pwell 13224 -12541 13258 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_157/VNB
rlabel comment 13195 -12524 13195 -12524 2 sky130_fd_sc_hd__decap_4_157/decap_4
rlabel metal1 13195 -12572 13563 -12476 5 sky130_fd_sc_hd__decap_4_157/VGND
rlabel metal1 13195 -13116 13563 -13020 5 sky130_fd_sc_hd__decap_4_157/VPWR
flabel metal1 13585 -13077 13638 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_314/VPWR
flabel metal1 13584 -12544 13635 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_314/VGND
rlabel comment 13563 -12524 13563 -12524 2 sky130_fd_sc_hd__tapvpwrvgnd_1_314/tapvpwrvgnd_1
rlabel metal1 13563 -12572 13655 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_314/VGND
rlabel metal1 13563 -13116 13655 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_314/VPWR
flabel metal1 13125 -13077 13178 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_315/VPWR
flabel metal1 13124 -12544 13175 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_315/VGND
rlabel comment 13103 -12524 13103 -12524 2 sky130_fd_sc_hd__tapvpwrvgnd_1_315/tapvpwrvgnd_1
rlabel metal1 13103 -12572 13195 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_315/VGND
rlabel metal1 13103 -13116 13195 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_315/VPWR
flabel metal1 12389 -13077 12442 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_316/VPWR
flabel metal1 12388 -12544 12439 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_316/VGND
rlabel comment 12367 -12524 12367 -12524 2 sky130_fd_sc_hd__tapvpwrvgnd_1_316/tapvpwrvgnd_1
rlabel metal1 12367 -12572 12459 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_316/VGND
rlabel metal1 12367 -13116 12459 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_316/VPWR
flabel metal1 15616 -12541 15650 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_22/VGND
flabel metal1 15616 -13085 15650 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_22/VPWR
flabel nwell 15616 -13085 15650 -13051 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_22/VPB
flabel pwell 15616 -12541 15650 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_22/VNB
rlabel comment 15587 -12524 15587 -12524 2 sky130_fd_sc_hd__decap_12_22/decap_12
rlabel metal1 15587 -12572 16691 -12476 5 sky130_fd_sc_hd__decap_12_22/VGND
rlabel metal1 15587 -13116 16691 -13020 5 sky130_fd_sc_hd__decap_12_22/VPWR
flabel metal1 15517 -13077 15570 -13048 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_317/VPWR
flabel metal1 15516 -12544 15567 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_317/VGND
rlabel comment 15495 -12524 15495 -12524 2 sky130_fd_sc_hd__tapvpwrvgnd_1_317/tapvpwrvgnd_1
rlabel metal1 15495 -12572 15587 -12476 5 sky130_fd_sc_hd__tapvpwrvgnd_1_317/VGND
rlabel metal1 15495 -13116 15587 -13020 5 sky130_fd_sc_hd__tapvpwrvgnd_1_317/VPWR
flabel metal1 -944 -11997 -910 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_27/VPWR
flabel metal1 -944 -12541 -910 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_27/VGND
flabel nwell -944 -11997 -910 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_27/VPB
flabel pwell -944 -12541 -910 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_27/VNB
rlabel comment -881 -12524 -881 -12524 6 sky130_fd_sc_hd__decap_8_27/decap_8
rlabel metal1 -1617 -12572 -881 -12476 1 sky130_fd_sc_hd__decap_8_27/VGND
rlabel metal1 -1617 -12028 -881 -11932 1 sky130_fd_sc_hd__decap_8_27/VPWR
flabel metal1 -2968 -11997 -2934 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_87/VPWR
flabel metal1 -2968 -12541 -2934 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_87/VGND
flabel nwell -2968 -11997 -2934 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_87/VPB
flabel pwell -2968 -12541 -2934 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_87/VNB
rlabel comment -2997 -12524 -2997 -12524 4 sky130_fd_sc_hd__decap_8_87/decap_8
rlabel metal1 -2997 -12572 -2261 -12476 1 sky130_fd_sc_hd__decap_8_87/VGND
rlabel metal1 -2997 -12028 -2261 -11932 1 sky130_fd_sc_hd__decap_8_87/VPWR
flabel metal1 -1781 -12538 -1728 -12506 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_26/VGND
flabel metal1 -1780 -11994 -1728 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_26/VPWR
flabel nwell -1773 -11989 -1739 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_26/VPB
flabel pwell -1770 -12534 -1738 -12512 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_26/VNB
rlabel comment -1801 -12524 -1801 -12524 4 sky130_fd_sc_hd__fill_2_26/fill_2
rlabel metal1 -1801 -12572 -1617 -12476 1 sky130_fd_sc_hd__fill_2_26/VGND
rlabel metal1 -1801 -12028 -1617 -11932 1 sky130_fd_sc_hd__fill_2_26/VPWR
flabel metal1 -2135 -12534 -2112 -12515 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_36/VGND
flabel metal1 -2135 -11989 -2115 -11972 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_36/VPWR
flabel nwell -2134 -11994 -2109 -11968 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_36/VPB
flabel pwell -2134 -12536 -2112 -12512 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_36/VNB
rlabel comment -2169 -12524 -2169 -12524 4 sky130_fd_sc_hd__fill_4_36/fill_4
rlabel metal1 -2169 -12572 -1801 -12476 1 sky130_fd_sc_hd__fill_4_36/VGND
rlabel metal1 -2169 -12028 -1801 -11932 1 sky130_fd_sc_hd__fill_4_36/VPWR
flabel metal1 -2239 -12000 -2186 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_552/VPWR
flabel metal1 -2240 -12542 -2189 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_552/VGND
rlabel comment -2261 -12524 -2261 -12524 4 sky130_fd_sc_hd__tapvpwrvgnd_1_552/tapvpwrvgnd_1
rlabel metal1 -2261 -12572 -2169 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_552/VGND
rlabel metal1 -2261 -12028 -2169 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_552/VPWR
flabel locali -209 -12303 -175 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/A
flabel locali -855 -12099 -821 -12065 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/X
flabel locali -855 -12167 -821 -12133 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/X
flabel locali -855 -12235 -821 -12201 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/X
flabel locali -855 -12303 -821 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/X
flabel locali -855 -12371 -821 -12337 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/X
flabel locali -855 -12439 -821 -12405 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/X
flabel pwell -209 -12541 -175 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/VNB
flabel nwell -209 -11997 -175 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/VPB
flabel metal1 -209 -12541 -175 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/VGND
flabel metal1 -209 -11997 -175 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_122/VPWR
rlabel comment -145 -12524 -145 -12524 6 sky130_fd_sc_hd__clkdlybuf4s50_1_122/clkdlybuf4s50_1
rlabel metal1 -881 -12572 -145 -12476 1 sky130_fd_sc_hd__clkdlybuf4s50_1_122/VGND
rlabel metal1 -881 -12028 -145 -11932 1 sky130_fd_sc_hd__clkdlybuf4s50_1_122/VPWR
flabel locali 1079 -12303 1113 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/A
flabel locali 433 -12099 467 -12065 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/X
flabel locali 433 -12167 467 -12133 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/X
flabel locali 433 -12235 467 -12201 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/X
flabel locali 433 -12303 467 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/X
flabel locali 433 -12371 467 -12337 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/X
flabel locali 433 -12439 467 -12405 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/X
flabel pwell 1079 -12541 1113 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/VNB
flabel nwell 1079 -11997 1113 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/VPB
flabel metal1 1079 -12541 1113 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/VGND
flabel metal1 1079 -11997 1113 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_123/VPWR
rlabel comment 1143 -12524 1143 -12524 6 sky130_fd_sc_hd__clkdlybuf4s50_1_123/clkdlybuf4s50_1
rlabel metal1 407 -12572 1143 -12476 1 sky130_fd_sc_hd__clkdlybuf4s50_1_123/VGND
rlabel metal1 407 -12028 1143 -11932 1 sky130_fd_sc_hd__clkdlybuf4s50_1_123/VPWR
flabel metal1 252 -12541 286 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_158/VGND
flabel metal1 252 -11997 286 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_158/VPWR
flabel nwell 252 -11997 286 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_158/VPB
flabel pwell 252 -12541 286 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_158/VNB
rlabel comment 315 -12524 315 -12524 6 sky130_fd_sc_hd__decap_4_158/decap_4
rlabel metal1 -53 -12572 315 -12476 1 sky130_fd_sc_hd__decap_4_158/VGND
rlabel metal1 -53 -12028 315 -11932 1 sky130_fd_sc_hd__decap_4_158/VPWR
flabel metal1 -128 -12000 -75 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_318/VPWR
flabel metal1 -125 -12542 -74 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_318/VGND
rlabel comment -53 -12524 -53 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_318/tapvpwrvgnd_1
rlabel metal1 -145 -12572 -53 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_318/VGND
rlabel metal1 -145 -12028 -53 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_318/VPWR
flabel metal1 332 -12000 385 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_319/VPWR
flabel metal1 335 -12542 386 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_319/VGND
rlabel comment 407 -12524 407 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_319/tapvpwrvgnd_1
rlabel metal1 315 -12572 407 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_319/VGND
rlabel metal1 315 -12028 407 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_319/VPWR
flabel metal1 1540 -12541 1574 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_159/VGND
flabel metal1 1540 -11997 1574 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_159/VPWR
flabel nwell 1540 -11997 1574 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_159/VPB
flabel pwell 1540 -12541 1574 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_159/VNB
rlabel comment 1603 -12524 1603 -12524 6 sky130_fd_sc_hd__decap_4_159/decap_4
rlabel metal1 1235 -12572 1603 -12476 1 sky130_fd_sc_hd__decap_4_159/VGND
rlabel metal1 1235 -12028 1603 -11932 1 sky130_fd_sc_hd__decap_4_159/VPWR
flabel metal1 2828 -12541 2862 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_160/VGND
flabel metal1 2828 -11997 2862 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_160/VPWR
flabel nwell 2828 -11997 2862 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_160/VPB
flabel pwell 2828 -12541 2862 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_160/VNB
rlabel comment 2891 -12524 2891 -12524 6 sky130_fd_sc_hd__decap_4_160/decap_4
rlabel metal1 2523 -12572 2891 -12476 1 sky130_fd_sc_hd__decap_4_160/VGND
rlabel metal1 2523 -12028 2891 -11932 1 sky130_fd_sc_hd__decap_4_160/VPWR
flabel metal1 1724 -11997 1758 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_138/VPWR
flabel metal1 1724 -12541 1758 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_138/VGND
flabel nwell 1724 -11997 1758 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_138/VPB
flabel pwell 1724 -12541 1758 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_138/VNB
rlabel comment 1695 -12524 1695 -12524 4 sky130_fd_sc_hd__decap_8_138/decap_8
rlabel metal1 1695 -12572 2431 -12476 1 sky130_fd_sc_hd__decap_8_138/VGND
rlabel metal1 1695 -12028 2431 -11932 1 sky130_fd_sc_hd__decap_8_138/VPWR
flabel metal1 1160 -12000 1213 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_320/VPWR
flabel metal1 1163 -12542 1214 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_320/VGND
rlabel comment 1235 -12524 1235 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_320/tapvpwrvgnd_1
rlabel metal1 1143 -12572 1235 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_320/VGND
rlabel metal1 1143 -12028 1235 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_320/VPWR
flabel metal1 1620 -12000 1673 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_321/VPWR
flabel metal1 1623 -12542 1674 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_321/VGND
rlabel comment 1695 -12524 1695 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_321/tapvpwrvgnd_1
rlabel metal1 1603 -12572 1695 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_321/VGND
rlabel metal1 1603 -12028 1695 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_321/VPWR
flabel metal1 2448 -12000 2501 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_322/VPWR
flabel metal1 2451 -12542 2502 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_322/VGND
rlabel comment 2523 -12524 2523 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_322/tapvpwrvgnd_1
rlabel metal1 2431 -12572 2523 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_322/VGND
rlabel metal1 2431 -12028 2523 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_322/VPWR
flabel locali 3655 -12303 3689 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/A
flabel locali 3009 -12099 3043 -12065 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X
flabel locali 3009 -12167 3043 -12133 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X
flabel locali 3009 -12235 3043 -12201 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X
flabel locali 3009 -12303 3043 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X
flabel locali 3009 -12371 3043 -12337 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X
flabel locali 3009 -12439 3043 -12405 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X
flabel pwell 3655 -12541 3689 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/VNB
flabel nwell 3655 -11997 3689 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/VPB
flabel metal1 3655 -12541 3689 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/VGND
flabel metal1 3655 -11997 3689 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_125/VPWR
rlabel comment 3719 -12524 3719 -12524 6 sky130_fd_sc_hd__clkdlybuf4s50_1_125/clkdlybuf4s50_1
rlabel metal1 2983 -12572 3719 -12476 1 sky130_fd_sc_hd__clkdlybuf4s50_1_125/VGND
rlabel metal1 2983 -12028 3719 -11932 1 sky130_fd_sc_hd__clkdlybuf4s50_1_125/VPWR
flabel metal1 4116 -12541 4150 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_161/VGND
flabel metal1 4116 -11997 4150 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_161/VPWR
flabel nwell 4116 -11997 4150 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_161/VPB
flabel pwell 4116 -12541 4150 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_161/VNB
rlabel comment 4179 -12524 4179 -12524 6 sky130_fd_sc_hd__decap_4_161/decap_4
rlabel metal1 3811 -12572 4179 -12476 1 sky130_fd_sc_hd__decap_4_161/VGND
rlabel metal1 3811 -12028 4179 -11932 1 sky130_fd_sc_hd__decap_4_161/VPWR
flabel metal1 4300 -11997 4334 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_144/VPWR
flabel metal1 4300 -12541 4334 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_144/VGND
flabel nwell 4300 -11997 4334 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_144/VPB
flabel pwell 4300 -12541 4334 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_144/VNB
rlabel comment 4271 -12524 4271 -12524 4 sky130_fd_sc_hd__decap_8_144/decap_8
rlabel metal1 4271 -12572 5007 -12476 1 sky130_fd_sc_hd__decap_8_144/VGND
rlabel metal1 4271 -12028 5007 -11932 1 sky130_fd_sc_hd__decap_8_144/VPWR
flabel metal1 2908 -12000 2961 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_323/VPWR
flabel metal1 2911 -12542 2962 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_323/VGND
rlabel comment 2983 -12524 2983 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_323/tapvpwrvgnd_1
rlabel metal1 2891 -12572 2983 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_323/VGND
rlabel metal1 2891 -12028 2983 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_323/VPWR
flabel metal1 4196 -12000 4249 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_324/VPWR
flabel metal1 4199 -12542 4250 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_324/VGND
rlabel comment 4271 -12524 4271 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_324/tapvpwrvgnd_1
rlabel metal1 4179 -12572 4271 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_324/VGND
rlabel metal1 4179 -12028 4271 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_324/VPWR
flabel metal1 3736 -12000 3789 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_325/VPWR
flabel metal1 3739 -12542 3790 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_325/VGND
rlabel comment 3811 -12524 3811 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_325/tapvpwrvgnd_1
rlabel metal1 3719 -12572 3811 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_325/VGND
rlabel metal1 3719 -12028 3811 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_325/VPWR
flabel locali 6231 -12303 6265 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/A
flabel locali 5585 -12099 5619 -12065 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X
flabel locali 5585 -12167 5619 -12133 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X
flabel locali 5585 -12235 5619 -12201 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X
flabel locali 5585 -12303 5619 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X
flabel locali 5585 -12371 5619 -12337 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X
flabel locali 5585 -12439 5619 -12405 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X
flabel pwell 6231 -12541 6265 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/VNB
flabel nwell 6231 -11997 6265 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/VPB
flabel metal1 6231 -12541 6265 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/VGND
flabel metal1 6231 -11997 6265 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_127/VPWR
rlabel comment 6295 -12524 6295 -12524 6 sky130_fd_sc_hd__clkdlybuf4s50_1_127/clkdlybuf4s50_1
rlabel metal1 5559 -12572 6295 -12476 1 sky130_fd_sc_hd__clkdlybuf4s50_1_127/VGND
rlabel metal1 5559 -12028 6295 -11932 1 sky130_fd_sc_hd__clkdlybuf4s50_1_127/VPWR
flabel metal1 5404 -12541 5438 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_162/VGND
flabel metal1 5404 -11997 5438 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_162/VPWR
flabel nwell 5404 -11997 5438 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_162/VPB
flabel pwell 5404 -12541 5438 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_162/VNB
rlabel comment 5467 -12524 5467 -12524 6 sky130_fd_sc_hd__decap_4_162/decap_4
rlabel metal1 5099 -12572 5467 -12476 1 sky130_fd_sc_hd__decap_4_162/VGND
rlabel metal1 5099 -12028 5467 -11932 1 sky130_fd_sc_hd__decap_4_162/VPWR
flabel metal1 6692 -12541 6726 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_163/VGND
flabel metal1 6692 -11997 6726 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_163/VPWR
flabel nwell 6692 -11997 6726 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_163/VPB
flabel pwell 6692 -12541 6726 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_163/VNB
rlabel comment 6755 -12524 6755 -12524 6 sky130_fd_sc_hd__decap_4_163/decap_4
rlabel metal1 6387 -12572 6755 -12476 1 sky130_fd_sc_hd__decap_4_163/VGND
rlabel metal1 6387 -12028 6755 -11932 1 sky130_fd_sc_hd__decap_4_163/VPWR
flabel metal1 5024 -12000 5077 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_326/VPWR
flabel metal1 5027 -12542 5078 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_326/VGND
rlabel comment 5099 -12524 5099 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_326/tapvpwrvgnd_1
rlabel metal1 5007 -12572 5099 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_326/VGND
rlabel metal1 5007 -12028 5099 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_326/VPWR
flabel metal1 5484 -12000 5537 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_327/VPWR
flabel metal1 5487 -12542 5538 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_327/VGND
rlabel comment 5559 -12524 5559 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_327/tapvpwrvgnd_1
rlabel metal1 5467 -12572 5559 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_327/VGND
rlabel metal1 5467 -12028 5559 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_327/VPWR
flabel metal1 6312 -12000 6365 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_328/VPWR
flabel metal1 6315 -12542 6366 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_328/VGND
rlabel comment 6387 -12524 6387 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_328/tapvpwrvgnd_1
rlabel metal1 6295 -12572 6387 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_328/VGND
rlabel metal1 6295 -12028 6387 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_328/VPWR
flabel locali 8807 -12303 8841 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/A
flabel locali 8161 -12099 8195 -12065 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X
flabel locali 8161 -12167 8195 -12133 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X
flabel locali 8161 -12235 8195 -12201 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X
flabel locali 8161 -12303 8195 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X
flabel locali 8161 -12371 8195 -12337 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X
flabel locali 8161 -12439 8195 -12405 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X
flabel pwell 8807 -12541 8841 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/VNB
flabel nwell 8807 -11997 8841 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/VPB
flabel metal1 8807 -12541 8841 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/VGND
flabel metal1 8807 -11997 8841 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_129/VPWR
rlabel comment 8871 -12524 8871 -12524 6 sky130_fd_sc_hd__clkdlybuf4s50_1_129/clkdlybuf4s50_1
rlabel metal1 8135 -12572 8871 -12476 1 sky130_fd_sc_hd__clkdlybuf4s50_1_129/VGND
rlabel metal1 8135 -12028 8871 -11932 1 sky130_fd_sc_hd__clkdlybuf4s50_1_129/VPWR
flabel metal1 7980 -12541 8014 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_164/VGND
flabel metal1 7980 -11997 8014 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_164/VPWR
flabel nwell 7980 -11997 8014 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_164/VPB
flabel pwell 7980 -12541 8014 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_164/VNB
rlabel comment 8043 -12524 8043 -12524 6 sky130_fd_sc_hd__decap_4_164/decap_4
rlabel metal1 7675 -12572 8043 -12476 1 sky130_fd_sc_hd__decap_4_164/VGND
rlabel metal1 7675 -12028 8043 -11932 1 sky130_fd_sc_hd__decap_4_164/VPWR
flabel metal1 6876 -11997 6910 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_154/VPWR
flabel metal1 6876 -12541 6910 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_154/VGND
flabel nwell 6876 -11997 6910 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_154/VPB
flabel pwell 6876 -12541 6910 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_154/VNB
rlabel comment 6847 -12524 6847 -12524 4 sky130_fd_sc_hd__decap_8_154/decap_8
rlabel metal1 6847 -12572 7583 -12476 1 sky130_fd_sc_hd__decap_8_154/VGND
rlabel metal1 6847 -12028 7583 -11932 1 sky130_fd_sc_hd__decap_8_154/VPWR
flabel metal1 6772 -12000 6825 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_329/VPWR
flabel metal1 6775 -12542 6826 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_329/VGND
rlabel comment 6847 -12524 6847 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_329/tapvpwrvgnd_1
rlabel metal1 6755 -12572 6847 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_329/VGND
rlabel metal1 6755 -12028 6847 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_329/VPWR
flabel metal1 8060 -12000 8113 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_330/VPWR
flabel metal1 8063 -12542 8114 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_330/VGND
rlabel comment 8135 -12524 8135 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_330/tapvpwrvgnd_1
rlabel metal1 8043 -12572 8135 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_330/VGND
rlabel metal1 8043 -12028 8135 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_330/VPWR
flabel metal1 7600 -12000 7653 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_331/VPWR
flabel metal1 7603 -12542 7654 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_331/VGND
rlabel comment 7675 -12524 7675 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_331/tapvpwrvgnd_1
rlabel metal1 7583 -12572 7675 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_331/VGND
rlabel metal1 7583 -12028 7675 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_331/VPWR
flabel metal1 9268 -12541 9302 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_165/VGND
flabel metal1 9268 -11997 9302 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_165/VPWR
flabel nwell 9268 -11997 9302 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_165/VPB
flabel pwell 9268 -12541 9302 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_165/VNB
rlabel comment 9331 -12524 9331 -12524 6 sky130_fd_sc_hd__decap_4_165/decap_4
rlabel metal1 8963 -12572 9331 -12476 1 sky130_fd_sc_hd__decap_4_165/VGND
rlabel metal1 8963 -12028 9331 -11932 1 sky130_fd_sc_hd__decap_4_165/VPWR
flabel metal1 10648 -12541 10682 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_166/VGND
flabel metal1 10648 -11997 10682 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_166/VPWR
flabel nwell 10648 -11997 10682 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_166/VPB
flabel pwell 10648 -12541 10682 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_166/VNB
rlabel comment 10711 -12524 10711 -12524 6 sky130_fd_sc_hd__decap_4_166/decap_4
rlabel metal1 10343 -12572 10711 -12476 1 sky130_fd_sc_hd__decap_4_166/VGND
rlabel metal1 10343 -12028 10711 -11932 1 sky130_fd_sc_hd__decap_4_166/VPWR
flabel metal1 9452 -11997 9486 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_163/VPWR
flabel metal1 9452 -12541 9486 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_163/VGND
flabel nwell 9452 -11997 9486 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_163/VPB
flabel pwell 9452 -12541 9486 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_163/VNB
rlabel comment 9423 -12524 9423 -12524 4 sky130_fd_sc_hd__decap_8_163/decap_8
rlabel metal1 9423 -12572 10159 -12476 1 sky130_fd_sc_hd__decap_8_163/VGND
rlabel metal1 9423 -12028 10159 -11932 1 sky130_fd_sc_hd__decap_8_163/VPWR
flabel metal1 10285 -11997 10321 -11967 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_44/VPWR
flabel metal1 10285 -12537 10321 -12508 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_44/VGND
flabel nwell 10292 -11990 10312 -11973 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_44/VPB
flabel pwell 10291 -12535 10315 -12513 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_44/VNB
rlabel comment 10343 -12524 10343 -12524 6 sky130_fd_sc_hd__fill_1_44/fill_1
rlabel metal1 10251 -12572 10343 -12476 1 sky130_fd_sc_hd__fill_1_44/VGND
rlabel metal1 10251 -12028 10343 -11932 1 sky130_fd_sc_hd__fill_1_44/VPWR
flabel metal1 8888 -12000 8941 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_332/VPWR
flabel metal1 8891 -12542 8942 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_332/VGND
rlabel comment 8963 -12524 8963 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_332/tapvpwrvgnd_1
rlabel metal1 8871 -12572 8963 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_332/VGND
rlabel metal1 8871 -12028 8963 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_332/VPWR
flabel metal1 9348 -12000 9401 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_333/VPWR
flabel metal1 9351 -12542 9402 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_333/VGND
rlabel comment 9423 -12524 9423 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_333/tapvpwrvgnd_1
rlabel metal1 9331 -12572 9423 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_333/VGND
rlabel metal1 9331 -12028 9423 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_333/VPWR
flabel metal1 10176 -12000 10229 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_334/VPWR
flabel metal1 10179 -12542 10230 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_334/VGND
rlabel comment 10251 -12524 10251 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_334/tapvpwrvgnd_1
rlabel metal1 10159 -12572 10251 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_334/VGND
rlabel metal1 10159 -12028 10251 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_334/VPWR
flabel locali 11383 -12303 11417 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A
flabel locali 10737 -12099 10771 -12065 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
flabel locali 10737 -12167 10771 -12133 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
flabel locali 10737 -12235 10771 -12201 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
flabel locali 10737 -12303 10771 -12269 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
flabel locali 10737 -12371 10771 -12337 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
flabel locali 10737 -12439 10771 -12405 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
flabel pwell 11383 -12541 11417 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/VNB
flabel nwell 11383 -11997 11417 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/VPB
flabel metal1 11383 -12541 11417 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/VGND
flabel metal1 11383 -11997 11417 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_131/VPWR
rlabel comment 11447 -12524 11447 -12524 6 sky130_fd_sc_hd__clkdlybuf4s50_1_131/clkdlybuf4s50_1
rlabel metal1 10711 -12572 11447 -12476 1 sky130_fd_sc_hd__clkdlybuf4s50_1_131/VGND
rlabel metal1 10711 -12028 11447 -11932 1 sky130_fd_sc_hd__clkdlybuf4s50_1_131/VPWR
flabel metal1 11936 -12541 11970 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_167/VGND
flabel metal1 11936 -11997 11970 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_167/VPWR
flabel nwell 11936 -11997 11970 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_167/VPB
flabel pwell 11936 -12541 11970 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_167/VNB
rlabel comment 11999 -12524 11999 -12524 6 sky130_fd_sc_hd__decap_4_167/decap_4
rlabel metal1 11631 -12572 11999 -12476 1 sky130_fd_sc_hd__decap_4_167/VGND
rlabel metal1 11631 -12028 11999 -11932 1 sky130_fd_sc_hd__decap_4_167/VPWR
flabel metal1 10653 -11997 10689 -11967 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_45/VPWR
flabel metal1 10653 -12537 10689 -12508 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_45/VGND
flabel nwell 10660 -11990 10680 -11973 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_45/VPB
flabel pwell 10659 -12535 10683 -12513 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_45/VNB
rlabel comment 10711 -12524 10711 -12524 6 sky130_fd_sc_hd__fill_1_45/fill_1
rlabel metal1 10619 -12572 10711 -12476 1 sky130_fd_sc_hd__fill_1_45/VGND
rlabel metal1 10619 -12028 10711 -11932 1 sky130_fd_sc_hd__fill_1_45/VPWR
flabel metal1 11573 -11997 11609 -11967 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_46/VPWR
flabel metal1 11573 -12537 11609 -12508 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_46/VGND
flabel nwell 11580 -11990 11600 -11973 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_46/VPB
flabel pwell 11579 -12535 11603 -12513 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_46/VNB
rlabel comment 11631 -12524 11631 -12524 6 sky130_fd_sc_hd__fill_1_46/fill_1
rlabel metal1 11539 -12572 11631 -12476 1 sky130_fd_sc_hd__fill_1_46/VGND
rlabel metal1 11539 -12028 11631 -11932 1 sky130_fd_sc_hd__fill_1_46/VPWR
flabel metal1 12668 -12544 12700 -12514 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_23/VGND
flabel metal1 12668 -12001 12706 -11969 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_23/VPWR
flabel nwell 12658 -12002 12715 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_23/VPB
flabel pwell 12665 -12548 12709 -12514 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_23/VNB
rlabel comment 12735 -12524 12735 -12524 6 sky130_fd_sc_hd__fill_8_23/fill_8
rlabel metal1 11999 -12572 12735 -12476 1 sky130_fd_sc_hd__fill_8_23/VGND
rlabel metal1 11999 -12028 12735 -11932 1 sky130_fd_sc_hd__fill_8_23/VPWR
flabel metal1 11464 -12000 11517 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_335/VPWR
flabel metal1 11467 -12542 11518 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_335/VGND
rlabel comment 11539 -12524 11539 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_335/tapvpwrvgnd_1
rlabel metal1 11447 -12572 11539 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_335/VGND
rlabel metal1 11447 -12028 11539 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_335/VPWR
flabel locali 15248 -12235 15282 -12201 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/X
flabel locali 15340 -12235 15374 -12201 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/X
flabel locali 15340 -12303 15374 -12269 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/X
flabel locali 15248 -12303 15282 -12269 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/X
flabel locali 15248 -12371 15282 -12337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/X
flabel locali 15340 -12371 15374 -12337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/X
flabel locali 13684 -12371 13718 -12337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/A
flabel locali 13684 -12303 13718 -12269 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/A
flabel pwell 13684 -12541 13718 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/VNB
flabel pwell 13701 -12524 13701 -12524 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/VNB
flabel nwell 13684 -11997 13718 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/VPB
flabel nwell 13701 -11980 13701 -11980 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/VPB
flabel metal1 13684 -12541 13718 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/VGND
flabel metal1 13684 -11997 13718 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_10/VPWR
rlabel comment 13655 -12524 13655 -12524 4 sky130_fd_sc_hd__clkbuf_16_10/clkbuf_16
rlabel metal1 13655 -12572 15495 -12476 1 sky130_fd_sc_hd__clkbuf_16_10/VGND
rlabel metal1 13655 -12028 15495 -11932 1 sky130_fd_sc_hd__clkbuf_16_10/VPWR
flabel metal1 13505 -11997 13541 -11967 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_47/VPWR
flabel metal1 13505 -12537 13541 -12508 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_47/VGND
flabel nwell 13512 -11990 13532 -11973 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_47/VPB
flabel pwell 13511 -12535 13535 -12513 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_47/VNB
rlabel comment 13563 -12524 13563 -12524 6 sky130_fd_sc_hd__fill_1_47/fill_1
rlabel metal1 13471 -12572 13563 -12476 1 sky130_fd_sc_hd__fill_1_47/VGND
rlabel metal1 13471 -12028 13563 -11932 1 sky130_fd_sc_hd__fill_1_47/VPWR
flabel metal1 13404 -12544 13436 -12514 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_24/VGND
flabel metal1 13404 -12001 13442 -11969 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_24/VPWR
flabel nwell 13394 -12002 13451 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_24/VPB
flabel pwell 13401 -12548 13445 -12514 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_24/VNB
rlabel comment 13471 -12524 13471 -12524 6 sky130_fd_sc_hd__fill_8_24/fill_8
rlabel metal1 12735 -12572 13471 -12476 1 sky130_fd_sc_hd__fill_8_24/VGND
rlabel metal1 12735 -12028 13471 -11932 1 sky130_fd_sc_hd__fill_8_24/VPWR
flabel metal1 13580 -12000 13633 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_336/VPWR
flabel metal1 13583 -12542 13634 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_336/VGND
rlabel comment 13655 -12524 13655 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_336/tapvpwrvgnd_1
rlabel metal1 13563 -12572 13655 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_336/VGND
rlabel metal1 13563 -12028 13655 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_336/VPWR
flabel metal1 16628 -12541 16662 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_23/VGND
flabel metal1 16628 -11997 16662 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_23/VPWR
flabel nwell 16628 -11997 16662 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_23/VPB
flabel pwell 16628 -12541 16662 -12507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_23/VNB
rlabel comment 16691 -12524 16691 -12524 6 sky130_fd_sc_hd__decap_12_23/decap_12
rlabel metal1 15587 -12572 16691 -12476 1 sky130_fd_sc_hd__decap_12_23/VGND
rlabel metal1 15587 -12028 16691 -11932 1 sky130_fd_sc_hd__decap_12_23/VPWR
flabel metal1 15512 -12000 15565 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_337/VPWR
flabel metal1 15515 -12542 15566 -12504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_337/VGND
rlabel comment 15587 -12524 15587 -12524 6 sky130_fd_sc_hd__tapvpwrvgnd_1_337/tapvpwrvgnd_1
rlabel metal1 15495 -12572 15587 -12476 1 sky130_fd_sc_hd__tapvpwrvgnd_1_337/VGND
rlabel metal1 15495 -12028 15587 -11932 1 sky130_fd_sc_hd__tapvpwrvgnd_1_337/VPWR
flabel metal1 -1588 -11997 -1554 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_28/VPWR
flabel metal1 -1588 -11453 -1554 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_28/VGND
flabel nwell -1588 -11997 -1554 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_28/VPB
flabel pwell -1588 -11453 -1554 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_28/VNB
rlabel comment -1617 -11436 -1617 -11436 2 sky130_fd_sc_hd__decap_8_28/decap_8
rlabel metal1 -1617 -11484 -881 -11388 5 sky130_fd_sc_hd__decap_8_28/VGND
rlabel metal1 -1617 -12028 -881 -11932 5 sky130_fd_sc_hd__decap_8_28/VPWR
flabel metal1 -2324 -11997 -2290 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_86/VPWR
flabel metal1 -2324 -11453 -2290 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_86/VGND
flabel nwell -2324 -11997 -2290 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_86/VPB
flabel pwell -2324 -11453 -2290 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_86/VNB
rlabel comment -2261 -11436 -2261 -11436 8 sky130_fd_sc_hd__decap_8_86/decap_8
rlabel metal1 -2997 -11484 -2261 -11388 5 sky130_fd_sc_hd__decap_8_86/VGND
rlabel metal1 -2997 -12028 -2261 -11932 5 sky130_fd_sc_hd__decap_8_86/VPWR
flabel metal1 -1690 -11454 -1637 -11422 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_25/VGND
flabel metal1 -1690 -11997 -1638 -11966 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_25/VPWR
flabel nwell -1679 -11989 -1645 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_25/VPB
flabel pwell -1680 -11448 -1648 -11426 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_25/VNB
rlabel comment -1617 -11436 -1617 -11436 8 sky130_fd_sc_hd__fill_2_25/fill_2
rlabel metal1 -1801 -11484 -1617 -11388 5 sky130_fd_sc_hd__fill_2_25/VGND
rlabel metal1 -1801 -12028 -1617 -11932 5 sky130_fd_sc_hd__fill_2_25/VPWR
flabel metal1 -1858 -11445 -1835 -11426 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_34/VGND
flabel metal1 -1855 -11988 -1835 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_34/VPWR
flabel nwell -1861 -11992 -1836 -11966 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_34/VPB
flabel pwell -1858 -11448 -1836 -11424 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_34/VNB
rlabel comment -1801 -11436 -1801 -11436 8 sky130_fd_sc_hd__fill_4_34/fill_4
rlabel metal1 -2169 -11484 -1801 -11388 5 sky130_fd_sc_hd__fill_4_34/VGND
rlabel metal1 -2169 -12028 -1801 -11932 5 sky130_fd_sc_hd__fill_4_34/VPWR
flabel metal1 -2244 -11989 -2191 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_551/VPWR
flabel metal1 -2241 -11456 -2190 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_551/VGND
rlabel comment -2169 -11436 -2169 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_551/tapvpwrvgnd_1
rlabel metal1 -2261 -11484 -2169 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_551/VGND
rlabel metal1 -2261 -12028 -2169 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_551/VPWR
flabel locali 437 -11691 471 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A
flabel locali 1083 -11895 1117 -11861 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/X
flabel locali 1083 -11827 1117 -11793 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/X
flabel locali 1083 -11759 1117 -11725 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/X
flabel locali 1083 -11691 1117 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/X
flabel locali 1083 -11623 1117 -11589 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/X
flabel locali 1083 -11555 1117 -11521 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/X
flabel pwell 437 -11453 471 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/VNB
flabel nwell 437 -11997 471 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/VPB
flabel metal1 437 -11453 471 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/VGND
flabel metal1 437 -11997 471 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_132/VPWR
rlabel comment 407 -11436 407 -11436 2 sky130_fd_sc_hd__clkdlybuf4s50_1_132/clkdlybuf4s50_1
rlabel metal1 407 -11484 1143 -11388 5 sky130_fd_sc_hd__clkdlybuf4s50_1_132/VGND
rlabel metal1 407 -12028 1143 -11932 5 sky130_fd_sc_hd__clkdlybuf4s50_1_132/VPWR
flabel metal1 252 -11453 286 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_168/VGND
flabel metal1 252 -11997 286 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_168/VPWR
flabel nwell 252 -11997 286 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_168/VPB
flabel pwell 252 -11453 286 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_168/VNB
rlabel comment 315 -11436 315 -11436 8 sky130_fd_sc_hd__decap_4_168/decap_4
rlabel metal1 -53 -11484 315 -11388 5 sky130_fd_sc_hd__decap_4_168/VGND
rlabel metal1 -53 -12028 315 -11932 5 sky130_fd_sc_hd__decap_4_168/VPWR
flabel metal1 -852 -11997 -818 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_29/VPWR
flabel metal1 -852 -11453 -818 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_29/VGND
flabel nwell -852 -11997 -818 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_29/VPB
flabel pwell -852 -11453 -818 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_29/VNB
rlabel comment -881 -11436 -881 -11436 2 sky130_fd_sc_hd__decap_8_29/decap_8
rlabel metal1 -881 -11484 -145 -11388 5 sky130_fd_sc_hd__decap_8_29/VGND
rlabel metal1 -881 -12028 -145 -11932 5 sky130_fd_sc_hd__decap_8_29/VPWR
flabel metal1 332 -11989 385 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_338/VPWR
flabel metal1 335 -11456 386 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_338/VGND
rlabel comment 407 -11436 407 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_338/tapvpwrvgnd_1
rlabel metal1 315 -11484 407 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_338/VGND
rlabel metal1 315 -12028 407 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_338/VPWR
flabel metal1 -128 -11989 -75 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_339/VPWR
flabel metal1 -125 -11456 -74 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_339/VGND
rlabel comment -53 -11436 -53 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_339/tapvpwrvgnd_1
rlabel metal1 -145 -11484 -53 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_339/VGND
rlabel metal1 -145 -12028 -53 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_339/VPWR
flabel metal1 1540 -11453 1574 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_169/VGND
flabel metal1 1540 -11997 1574 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_169/VPWR
flabel nwell 1540 -11997 1574 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_169/VPB
flabel pwell 1540 -11453 1574 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_169/VNB
rlabel comment 1603 -11436 1603 -11436 8 sky130_fd_sc_hd__decap_4_169/decap_4
rlabel metal1 1235 -11484 1603 -11388 5 sky130_fd_sc_hd__decap_4_169/VGND
rlabel metal1 1235 -12028 1603 -11932 5 sky130_fd_sc_hd__decap_4_169/VPWR
flabel metal1 2828 -11453 2862 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_170/VGND
flabel metal1 2828 -11997 2862 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_170/VPWR
flabel nwell 2828 -11997 2862 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_170/VPB
flabel pwell 2828 -11453 2862 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_170/VNB
rlabel comment 2891 -11436 2891 -11436 8 sky130_fd_sc_hd__decap_4_170/decap_4
rlabel metal1 2523 -11484 2891 -11388 5 sky130_fd_sc_hd__decap_4_170/VGND
rlabel metal1 2523 -12028 2891 -11932 5 sky130_fd_sc_hd__decap_4_170/VPWR
flabel metal1 2368 -11997 2402 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_137/VPWR
flabel metal1 2368 -11453 2402 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_137/VGND
flabel nwell 2368 -11997 2402 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_137/VPB
flabel pwell 2368 -11453 2402 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_137/VNB
rlabel comment 2431 -11436 2431 -11436 8 sky130_fd_sc_hd__decap_8_137/decap_8
rlabel metal1 1695 -11484 2431 -11388 5 sky130_fd_sc_hd__decap_8_137/VGND
rlabel metal1 1695 -12028 2431 -11932 5 sky130_fd_sc_hd__decap_8_137/VPWR
flabel metal1 1160 -11989 1213 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_340/VPWR
flabel metal1 1163 -11456 1214 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_340/VGND
rlabel comment 1235 -11436 1235 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_340/tapvpwrvgnd_1
rlabel metal1 1143 -11484 1235 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_340/VGND
rlabel metal1 1143 -12028 1235 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_340/VPWR
flabel metal1 1620 -11989 1673 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_341/VPWR
flabel metal1 1623 -11456 1674 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_341/VGND
rlabel comment 1695 -11436 1695 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_341/tapvpwrvgnd_1
rlabel metal1 1603 -11484 1695 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_341/VGND
rlabel metal1 1603 -12028 1695 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_341/VPWR
flabel metal1 2448 -11989 2501 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_342/VPWR
flabel metal1 2451 -11456 2502 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_342/VGND
rlabel comment 2523 -11436 2523 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_342/tapvpwrvgnd_1
rlabel metal1 2431 -11484 2523 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_342/VGND
rlabel metal1 2431 -12028 2523 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_342/VPWR
flabel locali 3013 -11691 3047 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A
flabel locali 3659 -11895 3693 -11861 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/X
flabel locali 3659 -11827 3693 -11793 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/X
flabel locali 3659 -11759 3693 -11725 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/X
flabel locali 3659 -11691 3693 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/X
flabel locali 3659 -11623 3693 -11589 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/X
flabel locali 3659 -11555 3693 -11521 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/X
flabel pwell 3013 -11453 3047 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/VNB
flabel nwell 3013 -11997 3047 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/VPB
flabel metal1 3013 -11453 3047 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/VGND
flabel metal1 3013 -11997 3047 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_134/VPWR
rlabel comment 2983 -11436 2983 -11436 2 sky130_fd_sc_hd__clkdlybuf4s50_1_134/clkdlybuf4s50_1
rlabel metal1 2983 -11484 3719 -11388 5 sky130_fd_sc_hd__clkdlybuf4s50_1_134/VGND
rlabel metal1 2983 -12028 3719 -11932 5 sky130_fd_sc_hd__clkdlybuf4s50_1_134/VPWR
flabel metal1 4116 -11453 4150 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_171/VGND
flabel metal1 4116 -11997 4150 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_171/VPWR
flabel nwell 4116 -11997 4150 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_171/VPB
flabel pwell 4116 -11453 4150 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_171/VNB
rlabel comment 4179 -11436 4179 -11436 8 sky130_fd_sc_hd__decap_4_171/decap_4
rlabel metal1 3811 -11484 4179 -11388 5 sky130_fd_sc_hd__decap_4_171/VGND
rlabel metal1 3811 -12028 4179 -11932 5 sky130_fd_sc_hd__decap_4_171/VPWR
flabel metal1 4944 -11997 4978 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_143/VPWR
flabel metal1 4944 -11453 4978 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_143/VGND
flabel nwell 4944 -11997 4978 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_143/VPB
flabel pwell 4944 -11453 4978 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_143/VNB
rlabel comment 5007 -11436 5007 -11436 8 sky130_fd_sc_hd__decap_8_143/decap_8
rlabel metal1 4271 -11484 5007 -11388 5 sky130_fd_sc_hd__decap_8_143/VGND
rlabel metal1 4271 -12028 5007 -11932 5 sky130_fd_sc_hd__decap_8_143/VPWR
flabel metal1 2908 -11989 2961 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_343/VPWR
flabel metal1 2911 -11456 2962 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_343/VGND
rlabel comment 2983 -11436 2983 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_343/tapvpwrvgnd_1
rlabel metal1 2891 -11484 2983 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_343/VGND
rlabel metal1 2891 -12028 2983 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_343/VPWR
flabel metal1 3736 -11989 3789 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_344/VPWR
flabel metal1 3739 -11456 3790 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_344/VGND
rlabel comment 3811 -11436 3811 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_344/tapvpwrvgnd_1
rlabel metal1 3719 -11484 3811 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_344/VGND
rlabel metal1 3719 -12028 3811 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_344/VPWR
flabel metal1 4196 -11989 4249 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_345/VPWR
flabel metal1 4199 -11456 4250 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_345/VGND
rlabel comment 4271 -11436 4271 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_345/tapvpwrvgnd_1
rlabel metal1 4179 -11484 4271 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_345/VGND
rlabel metal1 4179 -12028 4271 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_345/VPWR
flabel locali 5589 -11691 5623 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A
flabel locali 6235 -11895 6269 -11861 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/X
flabel locali 6235 -11827 6269 -11793 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/X
flabel locali 6235 -11759 6269 -11725 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/X
flabel locali 6235 -11691 6269 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/X
flabel locali 6235 -11623 6269 -11589 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/X
flabel locali 6235 -11555 6269 -11521 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/X
flabel pwell 5589 -11453 5623 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/VNB
flabel nwell 5589 -11997 5623 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/VPB
flabel metal1 5589 -11453 5623 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/VGND
flabel metal1 5589 -11997 5623 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_136/VPWR
rlabel comment 5559 -11436 5559 -11436 2 sky130_fd_sc_hd__clkdlybuf4s50_1_136/clkdlybuf4s50_1
rlabel metal1 5559 -11484 6295 -11388 5 sky130_fd_sc_hd__clkdlybuf4s50_1_136/VGND
rlabel metal1 5559 -12028 6295 -11932 5 sky130_fd_sc_hd__clkdlybuf4s50_1_136/VPWR
flabel metal1 5404 -11453 5438 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_172/VGND
flabel metal1 5404 -11997 5438 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_172/VPWR
flabel nwell 5404 -11997 5438 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_172/VPB
flabel pwell 5404 -11453 5438 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_172/VNB
rlabel comment 5467 -11436 5467 -11436 8 sky130_fd_sc_hd__decap_4_172/decap_4
rlabel metal1 5099 -11484 5467 -11388 5 sky130_fd_sc_hd__decap_4_172/VGND
rlabel metal1 5099 -12028 5467 -11932 5 sky130_fd_sc_hd__decap_4_172/VPWR
flabel metal1 6692 -11453 6726 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_173/VGND
flabel metal1 6692 -11997 6726 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_173/VPWR
flabel nwell 6692 -11997 6726 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_173/VPB
flabel pwell 6692 -11453 6726 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_173/VNB
rlabel comment 6755 -11436 6755 -11436 8 sky130_fd_sc_hd__decap_4_173/decap_4
rlabel metal1 6387 -11484 6755 -11388 5 sky130_fd_sc_hd__decap_4_173/VGND
rlabel metal1 6387 -12028 6755 -11932 5 sky130_fd_sc_hd__decap_4_173/VPWR
flabel metal1 5024 -11989 5077 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_346/VPWR
flabel metal1 5027 -11456 5078 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_346/VGND
rlabel comment 5099 -11436 5099 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_346/tapvpwrvgnd_1
rlabel metal1 5007 -11484 5099 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_346/VGND
rlabel metal1 5007 -12028 5099 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_346/VPWR
flabel metal1 5484 -11989 5537 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_347/VPWR
flabel metal1 5487 -11456 5538 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_347/VGND
rlabel comment 5559 -11436 5559 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_347/tapvpwrvgnd_1
rlabel metal1 5467 -11484 5559 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_347/VGND
rlabel metal1 5467 -12028 5559 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_347/VPWR
flabel metal1 6312 -11989 6365 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_348/VPWR
flabel metal1 6315 -11456 6366 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_348/VGND
rlabel comment 6387 -11436 6387 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_348/tapvpwrvgnd_1
rlabel metal1 6295 -11484 6387 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_348/VGND
rlabel metal1 6295 -12028 6387 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_348/VPWR
flabel locali 8165 -11691 8199 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A
flabel locali 8811 -11895 8845 -11861 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/X
flabel locali 8811 -11827 8845 -11793 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/X
flabel locali 8811 -11759 8845 -11725 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/X
flabel locali 8811 -11691 8845 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/X
flabel locali 8811 -11623 8845 -11589 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/X
flabel locali 8811 -11555 8845 -11521 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/X
flabel pwell 8165 -11453 8199 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/VNB
flabel nwell 8165 -11997 8199 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/VPB
flabel metal1 8165 -11453 8199 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/VGND
flabel metal1 8165 -11997 8199 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_138/VPWR
rlabel comment 8135 -11436 8135 -11436 2 sky130_fd_sc_hd__clkdlybuf4s50_1_138/clkdlybuf4s50_1
rlabel metal1 8135 -11484 8871 -11388 5 sky130_fd_sc_hd__clkdlybuf4s50_1_138/VGND
rlabel metal1 8135 -12028 8871 -11932 5 sky130_fd_sc_hd__clkdlybuf4s50_1_138/VPWR
flabel metal1 7980 -11453 8014 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_174/VGND
flabel metal1 7980 -11997 8014 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_174/VPWR
flabel nwell 7980 -11997 8014 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_174/VPB
flabel pwell 7980 -11453 8014 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_174/VNB
rlabel comment 8043 -11436 8043 -11436 8 sky130_fd_sc_hd__decap_4_174/decap_4
rlabel metal1 7675 -11484 8043 -11388 5 sky130_fd_sc_hd__decap_4_174/VGND
rlabel metal1 7675 -12028 8043 -11932 5 sky130_fd_sc_hd__decap_4_174/VPWR
flabel metal1 7520 -11997 7554 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_153/VPWR
flabel metal1 7520 -11453 7554 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_153/VGND
flabel nwell 7520 -11997 7554 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_153/VPB
flabel pwell 7520 -11453 7554 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_153/VNB
rlabel comment 7583 -11436 7583 -11436 8 sky130_fd_sc_hd__decap_8_153/decap_8
rlabel metal1 6847 -11484 7583 -11388 5 sky130_fd_sc_hd__decap_8_153/VGND
rlabel metal1 6847 -12028 7583 -11932 5 sky130_fd_sc_hd__decap_8_153/VPWR
flabel metal1 6772 -11989 6825 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_349/VPWR
flabel metal1 6775 -11456 6826 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_349/VGND
rlabel comment 6847 -11436 6847 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_349/tapvpwrvgnd_1
rlabel metal1 6755 -11484 6847 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_349/VGND
rlabel metal1 6755 -12028 6847 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_349/VPWR
flabel metal1 7600 -11989 7653 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_350/VPWR
flabel metal1 7603 -11456 7654 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_350/VGND
rlabel comment 7675 -11436 7675 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_350/tapvpwrvgnd_1
rlabel metal1 7583 -11484 7675 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_350/VGND
rlabel metal1 7583 -12028 7675 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_350/VPWR
flabel metal1 8060 -11989 8113 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_351/VPWR
flabel metal1 8063 -11456 8114 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_351/VGND
rlabel comment 8135 -11436 8135 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_351/tapvpwrvgnd_1
rlabel metal1 8043 -11484 8135 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_351/VGND
rlabel metal1 8043 -12028 8135 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_351/VPWR
flabel metal1 9268 -11453 9302 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_175/VGND
flabel metal1 9268 -11997 9302 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_175/VPWR
flabel nwell 9268 -11997 9302 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_175/VPB
flabel pwell 9268 -11453 9302 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_175/VNB
rlabel comment 9331 -11436 9331 -11436 8 sky130_fd_sc_hd__decap_4_175/decap_4
rlabel metal1 8963 -11484 9331 -11388 5 sky130_fd_sc_hd__decap_4_175/VGND
rlabel metal1 8963 -12028 9331 -11932 5 sky130_fd_sc_hd__decap_4_175/VPWR
flabel metal1 10648 -11453 10682 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_176/VGND
flabel metal1 10648 -11997 10682 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_176/VPWR
flabel nwell 10648 -11997 10682 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_176/VPB
flabel pwell 10648 -11453 10682 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_176/VNB
rlabel comment 10711 -11436 10711 -11436 8 sky130_fd_sc_hd__decap_4_176/decap_4
rlabel metal1 10343 -11484 10711 -11388 5 sky130_fd_sc_hd__decap_4_176/VGND
rlabel metal1 10343 -12028 10711 -11932 5 sky130_fd_sc_hd__decap_4_176/VPWR
flabel metal1 10096 -11997 10130 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_164/VPWR
flabel metal1 10096 -11453 10130 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_164/VGND
flabel nwell 10096 -11997 10130 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_164/VPB
flabel pwell 10096 -11453 10130 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_164/VNB
rlabel comment 10159 -11436 10159 -11436 8 sky130_fd_sc_hd__decap_8_164/decap_8
rlabel metal1 9423 -11484 10159 -11388 5 sky130_fd_sc_hd__decap_8_164/VGND
rlabel metal1 9423 -12028 10159 -11932 5 sky130_fd_sc_hd__decap_8_164/VPWR
flabel metal1 10285 -11993 10321 -11963 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_48/VPWR
flabel metal1 10285 -11452 10321 -11423 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_48/VGND
flabel nwell 10292 -11987 10312 -11970 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_48/VPB
flabel pwell 10291 -11447 10315 -11425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_48/VNB
rlabel comment 10343 -11436 10343 -11436 8 sky130_fd_sc_hd__fill_1_48/fill_1
rlabel metal1 10251 -11484 10343 -11388 5 sky130_fd_sc_hd__fill_1_48/VGND
rlabel metal1 10251 -12028 10343 -11932 5 sky130_fd_sc_hd__fill_1_48/VPWR
flabel metal1 8888 -11989 8941 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_352/VPWR
flabel metal1 8891 -11456 8942 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_352/VGND
rlabel comment 8963 -11436 8963 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_352/tapvpwrvgnd_1
rlabel metal1 8871 -11484 8963 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_352/VGND
rlabel metal1 8871 -12028 8963 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_352/VPWR
flabel metal1 9348 -11989 9401 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_353/VPWR
flabel metal1 9351 -11456 9402 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_353/VGND
rlabel comment 9423 -11436 9423 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_353/tapvpwrvgnd_1
rlabel metal1 9331 -11484 9423 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_353/VGND
rlabel metal1 9331 -12028 9423 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_353/VPWR
flabel metal1 10176 -11989 10229 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_354/VPWR
flabel metal1 10179 -11456 10230 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_354/VGND
rlabel comment 10251 -11436 10251 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_354/tapvpwrvgnd_1
rlabel metal1 10159 -11484 10251 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_354/VGND
rlabel metal1 10159 -12028 10251 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_354/VPWR
flabel locali 10741 -11691 10775 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A
flabel locali 11387 -11895 11421 -11861 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/X
flabel locali 11387 -11827 11421 -11793 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/X
flabel locali 11387 -11759 11421 -11725 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/X
flabel locali 11387 -11691 11421 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/X
flabel locali 11387 -11623 11421 -11589 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/X
flabel locali 11387 -11555 11421 -11521 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/X
flabel pwell 10741 -11453 10775 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/VNB
flabel nwell 10741 -11997 10775 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/VPB
flabel metal1 10741 -11453 10775 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/VGND
flabel metal1 10741 -11997 10775 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_140/VPWR
rlabel comment 10711 -11436 10711 -11436 2 sky130_fd_sc_hd__clkdlybuf4s50_1_140/clkdlybuf4s50_1
rlabel metal1 10711 -11484 11447 -11388 5 sky130_fd_sc_hd__clkdlybuf4s50_1_140/VGND
rlabel metal1 10711 -12028 11447 -11932 5 sky130_fd_sc_hd__clkdlybuf4s50_1_140/VPWR
flabel metal1 11936 -11453 11970 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_177/VGND
flabel metal1 11936 -11997 11970 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_177/VPWR
flabel nwell 11936 -11997 11970 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_177/VPB
flabel pwell 11936 -11453 11970 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_177/VNB
rlabel comment 11999 -11436 11999 -11436 8 sky130_fd_sc_hd__decap_4_177/decap_4
rlabel metal1 11631 -11484 11999 -11388 5 sky130_fd_sc_hd__decap_4_177/VGND
rlabel metal1 11631 -12028 11999 -11932 5 sky130_fd_sc_hd__decap_4_177/VPWR
flabel metal1 10653 -11993 10689 -11963 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_49/VPWR
flabel metal1 10653 -11452 10689 -11423 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_49/VGND
flabel nwell 10660 -11987 10680 -11970 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_49/VPB
flabel pwell 10659 -11447 10683 -11425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_49/VNB
rlabel comment 10711 -11436 10711 -11436 8 sky130_fd_sc_hd__fill_1_49/fill_1
rlabel metal1 10619 -11484 10711 -11388 5 sky130_fd_sc_hd__fill_1_49/VGND
rlabel metal1 10619 -12028 10711 -11932 5 sky130_fd_sc_hd__fill_1_49/VPWR
flabel metal1 11573 -11993 11609 -11963 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_50/VPWR
flabel metal1 11573 -11452 11609 -11423 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_50/VGND
flabel nwell 11580 -11987 11600 -11970 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_50/VPB
flabel pwell 11579 -11447 11603 -11425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_50/VNB
rlabel comment 11631 -11436 11631 -11436 8 sky130_fd_sc_hd__fill_1_50/fill_1
rlabel metal1 11539 -11484 11631 -11388 5 sky130_fd_sc_hd__fill_1_50/VGND
rlabel metal1 11539 -12028 11631 -11932 5 sky130_fd_sc_hd__fill_1_50/VPWR
flabel metal1 12033 -11445 12056 -11426 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_11/VGND
flabel metal1 12033 -11988 12053 -11971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_11/VPWR
flabel nwell 12034 -11992 12059 -11966 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_11/VPB
flabel pwell 12034 -11448 12056 -11424 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_11/VNB
rlabel comment 11999 -11436 11999 -11436 2 sky130_fd_sc_hd__fill_4_11/fill_4
rlabel metal1 11999 -11484 12367 -11388 5 sky130_fd_sc_hd__fill_4_11/VGND
rlabel metal1 11999 -12028 12367 -11932 5 sky130_fd_sc_hd__fill_4_11/VPWR
flabel metal1 11464 -11989 11517 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_355/VPWR
flabel metal1 11467 -11456 11518 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_355/VGND
rlabel comment 11539 -11436 11539 -11436 8 sky130_fd_sc_hd__tapvpwrvgnd_1_355/tapvpwrvgnd_1
rlabel metal1 11447 -11484 11539 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_355/VGND
rlabel metal1 11447 -12028 11539 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_355/VPWR
flabel locali 15248 -11759 15282 -11725 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/X
flabel locali 15340 -11759 15374 -11725 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/X
flabel locali 15340 -11691 15374 -11657 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/X
flabel locali 15248 -11691 15282 -11657 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/X
flabel locali 15248 -11623 15282 -11589 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/X
flabel locali 15340 -11623 15374 -11589 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/X
flabel locali 13684 -11623 13718 -11589 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/A
flabel locali 13684 -11691 13718 -11657 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/A
flabel pwell 13684 -11453 13718 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/VNB
flabel pwell 13701 -11436 13701 -11436 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/VNB
flabel nwell 13684 -11997 13718 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/VPB
flabel nwell 13701 -11980 13701 -11980 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/VPB
flabel metal1 13684 -11453 13718 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/VGND
flabel metal1 13684 -11997 13718 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_11/VPWR
rlabel comment 13655 -11436 13655 -11436 2 sky130_fd_sc_hd__clkbuf_16_11/clkbuf_16
rlabel metal1 13655 -11484 15495 -11388 5 sky130_fd_sc_hd__clkbuf_16_11/VGND
rlabel metal1 13655 -12028 15495 -11932 5 sky130_fd_sc_hd__clkbuf_16_11/VPWR
flabel locali 12672 -11691 12706 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/A
flabel locali 12764 -11691 12798 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/A
flabel locali 13040 -11623 13074 -11589 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/Y
flabel locali 12580 -11691 12614 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/A
flabel locali 13040 -11759 13074 -11725 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/Y
flabel locali 12948 -11691 12982 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/A
flabel locali 12856 -11691 12890 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/A
flabel locali 13040 -11691 13074 -11657 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_8/Y
flabel pwell 12488 -11453 12522 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_8/VNB
flabel nwell 12488 -11997 12522 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_8/VPB
flabel metal1 12488 -11997 12522 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_8/VPWR
flabel metal1 12488 -11453 12522 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_8/VGND
rlabel comment 12459 -11436 12459 -11436 2 sky130_fd_sc_hd__clkinv_4_8/clkinv_4
rlabel metal1 12459 -11484 13103 -11388 5 sky130_fd_sc_hd__clkinv_4_8/VGND
rlabel metal1 12459 -12028 13103 -11932 5 sky130_fd_sc_hd__clkinv_4_8/VPWR
flabel metal1 13224 -11453 13258 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_178/VGND
flabel metal1 13224 -11997 13258 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_178/VPWR
flabel nwell 13224 -11997 13258 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_178/VPB
flabel pwell 13224 -11453 13258 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_178/VNB
rlabel comment 13195 -11436 13195 -11436 2 sky130_fd_sc_hd__decap_4_178/decap_4
rlabel metal1 13195 -11484 13563 -11388 5 sky130_fd_sc_hd__decap_4_178/VGND
rlabel metal1 13195 -12028 13563 -11932 5 sky130_fd_sc_hd__decap_4_178/VPWR
flabel metal1 12389 -11989 12442 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_356/VPWR
flabel metal1 12388 -11456 12439 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_356/VGND
rlabel comment 12367 -11436 12367 -11436 2 sky130_fd_sc_hd__tapvpwrvgnd_1_356/tapvpwrvgnd_1
rlabel metal1 12367 -11484 12459 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_356/VGND
rlabel metal1 12367 -12028 12459 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_356/VPWR
flabel metal1 13585 -11989 13638 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_357/VPWR
flabel metal1 13584 -11456 13635 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_357/VGND
rlabel comment 13563 -11436 13563 -11436 2 sky130_fd_sc_hd__tapvpwrvgnd_1_357/tapvpwrvgnd_1
rlabel metal1 13563 -11484 13655 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_357/VGND
rlabel metal1 13563 -12028 13655 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_357/VPWR
flabel metal1 13125 -11989 13178 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_358/VPWR
flabel metal1 13124 -11456 13175 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_358/VGND
rlabel comment 13103 -11436 13103 -11436 2 sky130_fd_sc_hd__tapvpwrvgnd_1_358/tapvpwrvgnd_1
rlabel metal1 13103 -11484 13195 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_358/VGND
rlabel metal1 13103 -12028 13195 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_358/VPWR
flabel metal1 15616 -11453 15650 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_24/VGND
flabel metal1 15616 -11997 15650 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_24/VPWR
flabel nwell 15616 -11997 15650 -11963 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_24/VPB
flabel pwell 15616 -11453 15650 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_24/VNB
rlabel comment 15587 -11436 15587 -11436 2 sky130_fd_sc_hd__decap_12_24/decap_12
rlabel metal1 15587 -11484 16691 -11388 5 sky130_fd_sc_hd__decap_12_24/VGND
rlabel metal1 15587 -12028 16691 -11932 5 sky130_fd_sc_hd__decap_12_24/VPWR
flabel metal1 15517 -11989 15570 -11960 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_359/VPWR
flabel metal1 15516 -11456 15567 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_359/VGND
rlabel comment 15495 -11436 15495 -11436 2 sky130_fd_sc_hd__tapvpwrvgnd_1_359/tapvpwrvgnd_1
rlabel metal1 15495 -11484 15587 -11388 5 sky130_fd_sc_hd__tapvpwrvgnd_1_359/VGND
rlabel metal1 15495 -12028 15587 -11932 5 sky130_fd_sc_hd__tapvpwrvgnd_1_359/VPWR
flabel metal1 -944 -10909 -910 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_31/VPWR
flabel metal1 -944 -11453 -910 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_31/VGND
flabel nwell -944 -10909 -910 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_31/VPB
flabel pwell -944 -11453 -910 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_31/VNB
rlabel comment -881 -11436 -881 -11436 6 sky130_fd_sc_hd__decap_8_31/decap_8
rlabel metal1 -1617 -11484 -881 -11388 1 sky130_fd_sc_hd__decap_8_31/VGND
rlabel metal1 -1617 -10940 -881 -10844 1 sky130_fd_sc_hd__decap_8_31/VPWR
flabel metal1 -2968 -10909 -2934 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_85/VPWR
flabel metal1 -2968 -11453 -2934 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_85/VGND
flabel nwell -2968 -10909 -2934 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_85/VPB
flabel pwell -2968 -11453 -2934 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_85/VNB
rlabel comment -2997 -11436 -2997 -11436 4 sky130_fd_sc_hd__decap_8_85/decap_8
rlabel metal1 -2997 -11484 -2261 -11388 1 sky130_fd_sc_hd__decap_8_85/VGND
rlabel metal1 -2997 -10940 -2261 -10844 1 sky130_fd_sc_hd__decap_8_85/VPWR
flabel metal1 -1781 -11450 -1728 -11418 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_24/VGND
flabel metal1 -1780 -10906 -1728 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_24/VPWR
flabel nwell -1773 -10901 -1739 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_24/VPB
flabel pwell -1770 -11446 -1738 -11424 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_24/VNB
rlabel comment -1801 -11436 -1801 -11436 4 sky130_fd_sc_hd__fill_2_24/fill_2
rlabel metal1 -1801 -11484 -1617 -11388 1 sky130_fd_sc_hd__fill_2_24/VGND
rlabel metal1 -1801 -10940 -1617 -10844 1 sky130_fd_sc_hd__fill_2_24/VPWR
flabel metal1 -2135 -11446 -2112 -11427 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_33/VGND
flabel metal1 -2135 -10901 -2115 -10884 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_33/VPWR
flabel nwell -2134 -10906 -2109 -10880 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_33/VPB
flabel pwell -2134 -11448 -2112 -11424 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_33/VNB
rlabel comment -2169 -11436 -2169 -11436 4 sky130_fd_sc_hd__fill_4_33/fill_4
rlabel metal1 -2169 -11484 -1801 -11388 1 sky130_fd_sc_hd__fill_4_33/VGND
rlabel metal1 -2169 -10940 -1801 -10844 1 sky130_fd_sc_hd__fill_4_33/VPWR
flabel metal1 -2239 -10912 -2186 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_550/VPWR
flabel metal1 -2240 -11454 -2189 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_550/VGND
rlabel comment -2261 -11436 -2261 -11436 4 sky130_fd_sc_hd__tapvpwrvgnd_1_550/tapvpwrvgnd_1
rlabel metal1 -2261 -11484 -2169 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_550/VGND
rlabel metal1 -2261 -10940 -2169 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_550/VPWR
flabel locali 1079 -11215 1113 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/A
flabel locali 433 -11011 467 -10977 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X
flabel locali 433 -11079 467 -11045 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X
flabel locali 433 -11147 467 -11113 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X
flabel locali 433 -11215 467 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X
flabel locali 433 -11283 467 -11249 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X
flabel locali 433 -11351 467 -11317 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X
flabel pwell 1079 -11453 1113 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/VNB
flabel nwell 1079 -10909 1113 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/VPB
flabel metal1 1079 -11453 1113 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/VGND
flabel metal1 1079 -10909 1113 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_142/VPWR
rlabel comment 1143 -11436 1143 -11436 6 sky130_fd_sc_hd__clkdlybuf4s50_1_142/clkdlybuf4s50_1
rlabel metal1 407 -11484 1143 -11388 1 sky130_fd_sc_hd__clkdlybuf4s50_1_142/VGND
rlabel metal1 407 -10940 1143 -10844 1 sky130_fd_sc_hd__clkdlybuf4s50_1_142/VPWR
flabel metal1 252 -11453 286 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_180/VGND
flabel metal1 252 -10909 286 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_180/VPWR
flabel nwell 252 -10909 286 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_180/VPB
flabel pwell 252 -11453 286 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_180/VNB
rlabel comment 315 -11436 315 -11436 6 sky130_fd_sc_hd__decap_4_180/decap_4
rlabel metal1 -53 -11484 315 -11388 1 sky130_fd_sc_hd__decap_4_180/VGND
rlabel metal1 -53 -10940 315 -10844 1 sky130_fd_sc_hd__decap_4_180/VPWR
flabel metal1 -208 -10909 -174 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_33/VPWR
flabel metal1 -208 -11453 -174 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_33/VGND
flabel nwell -208 -10909 -174 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_33/VPB
flabel pwell -208 -11453 -174 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_33/VNB
rlabel comment -145 -11436 -145 -11436 6 sky130_fd_sc_hd__decap_8_33/decap_8
rlabel metal1 -881 -11484 -145 -11388 1 sky130_fd_sc_hd__decap_8_33/VGND
rlabel metal1 -881 -10940 -145 -10844 1 sky130_fd_sc_hd__decap_8_33/VPWR
flabel metal1 332 -10912 385 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_362/VPWR
flabel metal1 335 -11454 386 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_362/VGND
rlabel comment 407 -11436 407 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_362/tapvpwrvgnd_1
rlabel metal1 315 -11484 407 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_362/VGND
rlabel metal1 315 -10940 407 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_362/VPWR
flabel metal1 -128 -10912 -75 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_363/VPWR
flabel metal1 -125 -11454 -74 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_363/VGND
rlabel comment -53 -11436 -53 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_363/tapvpwrvgnd_1
rlabel metal1 -145 -11484 -53 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_363/VGND
rlabel metal1 -145 -10940 -53 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_363/VPWR
flabel metal1 1540 -11453 1574 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_183/VGND
flabel metal1 1540 -10909 1574 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_183/VPWR
flabel nwell 1540 -10909 1574 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_183/VPB
flabel pwell 1540 -11453 1574 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_183/VNB
rlabel comment 1603 -11436 1603 -11436 6 sky130_fd_sc_hd__decap_4_183/decap_4
rlabel metal1 1235 -11484 1603 -11388 1 sky130_fd_sc_hd__decap_4_183/VGND
rlabel metal1 1235 -10940 1603 -10844 1 sky130_fd_sc_hd__decap_4_183/VPWR
flabel metal1 2828 -11453 2862 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_184/VGND
flabel metal1 2828 -10909 2862 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_184/VPWR
flabel nwell 2828 -10909 2862 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_184/VPB
flabel pwell 2828 -11453 2862 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_184/VNB
rlabel comment 2891 -11436 2891 -11436 6 sky130_fd_sc_hd__decap_4_184/decap_4
rlabel metal1 2523 -11484 2891 -11388 1 sky130_fd_sc_hd__decap_4_184/VGND
rlabel metal1 2523 -10940 2891 -10844 1 sky130_fd_sc_hd__decap_4_184/VPWR
flabel metal1 1724 -10909 1758 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_136/VPWR
flabel metal1 1724 -11453 1758 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_136/VGND
flabel nwell 1724 -10909 1758 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_136/VPB
flabel pwell 1724 -11453 1758 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_136/VNB
rlabel comment 1695 -11436 1695 -11436 4 sky130_fd_sc_hd__decap_8_136/decap_8
rlabel metal1 1695 -11484 2431 -11388 1 sky130_fd_sc_hd__decap_8_136/VGND
rlabel metal1 1695 -10940 2431 -10844 1 sky130_fd_sc_hd__decap_8_136/VPWR
flabel metal1 1160 -10912 1213 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_367/VPWR
flabel metal1 1163 -11454 1214 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_367/VGND
rlabel comment 1235 -11436 1235 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_367/tapvpwrvgnd_1
rlabel metal1 1143 -11484 1235 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_367/VGND
rlabel metal1 1143 -10940 1235 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_367/VPWR
flabel metal1 1620 -10912 1673 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_368/VPWR
flabel metal1 1623 -11454 1674 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_368/VGND
rlabel comment 1695 -11436 1695 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_368/tapvpwrvgnd_1
rlabel metal1 1603 -11484 1695 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_368/VGND
rlabel metal1 1603 -10940 1695 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_368/VPWR
flabel metal1 2448 -10912 2501 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_369/VPWR
flabel metal1 2451 -11454 2502 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_369/VGND
rlabel comment 2523 -11436 2523 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_369/tapvpwrvgnd_1
rlabel metal1 2431 -11484 2523 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_369/VGND
rlabel metal1 2431 -10940 2523 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_369/VPWR
flabel locali 3655 -11215 3689 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/A
flabel locali 3009 -11011 3043 -10977 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
flabel locali 3009 -11079 3043 -11045 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
flabel locali 3009 -11147 3043 -11113 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
flabel locali 3009 -11215 3043 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
flabel locali 3009 -11283 3043 -11249 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
flabel locali 3009 -11351 3043 -11317 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
flabel pwell 3655 -11453 3689 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/VNB
flabel nwell 3655 -10909 3689 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/VPB
flabel metal1 3655 -11453 3689 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/VGND
flabel metal1 3655 -10909 3689 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_147/VPWR
rlabel comment 3719 -11436 3719 -11436 6 sky130_fd_sc_hd__clkdlybuf4s50_1_147/clkdlybuf4s50_1
rlabel metal1 2983 -11484 3719 -11388 1 sky130_fd_sc_hd__clkdlybuf4s50_1_147/VGND
rlabel metal1 2983 -10940 3719 -10844 1 sky130_fd_sc_hd__clkdlybuf4s50_1_147/VPWR
flabel metal1 4116 -11453 4150 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_186/VGND
flabel metal1 4116 -10909 4150 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_186/VPWR
flabel nwell 4116 -10909 4150 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_186/VPB
flabel pwell 4116 -11453 4150 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_186/VNB
rlabel comment 4179 -11436 4179 -11436 6 sky130_fd_sc_hd__decap_4_186/decap_4
rlabel metal1 3811 -11484 4179 -11388 1 sky130_fd_sc_hd__decap_4_186/VGND
rlabel metal1 3811 -10940 4179 -10844 1 sky130_fd_sc_hd__decap_4_186/VPWR
flabel metal1 4300 -10909 4334 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_146/VPWR
flabel metal1 4300 -11453 4334 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_146/VGND
flabel nwell 4300 -10909 4334 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_146/VPB
flabel pwell 4300 -11453 4334 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_146/VNB
rlabel comment 4271 -11436 4271 -11436 4 sky130_fd_sc_hd__decap_8_146/decap_8
rlabel metal1 4271 -11484 5007 -11388 1 sky130_fd_sc_hd__decap_8_146/VGND
rlabel metal1 4271 -10940 5007 -10844 1 sky130_fd_sc_hd__decap_8_146/VPWR
flabel metal1 2908 -10912 2961 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_373/VPWR
flabel metal1 2911 -11454 2962 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_373/VGND
rlabel comment 2983 -11436 2983 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_373/tapvpwrvgnd_1
rlabel metal1 2891 -11484 2983 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_373/VGND
rlabel metal1 2891 -10940 2983 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_373/VPWR
flabel metal1 3736 -10912 3789 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_374/VPWR
flabel metal1 3739 -11454 3790 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_374/VGND
rlabel comment 3811 -11436 3811 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_374/tapvpwrvgnd_1
rlabel metal1 3719 -11484 3811 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_374/VGND
rlabel metal1 3719 -10940 3811 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_374/VPWR
flabel metal1 4196 -10912 4249 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_375/VPWR
flabel metal1 4199 -11454 4250 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_375/VGND
rlabel comment 4271 -11436 4271 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_375/tapvpwrvgnd_1
rlabel metal1 4179 -11484 4271 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_375/VGND
rlabel metal1 4179 -10940 4271 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_375/VPWR
flabel locali 6231 -11215 6265 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/A
flabel locali 5585 -11011 5619 -10977 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
flabel locali 5585 -11079 5619 -11045 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
flabel locali 5585 -11147 5619 -11113 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
flabel locali 5585 -11215 5619 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
flabel locali 5585 -11283 5619 -11249 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
flabel locali 5585 -11351 5619 -11317 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
flabel pwell 6231 -11453 6265 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/VNB
flabel nwell 6231 -10909 6265 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/VPB
flabel metal1 6231 -11453 6265 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/VGND
flabel metal1 6231 -10909 6265 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_150/VPWR
rlabel comment 6295 -11436 6295 -11436 6 sky130_fd_sc_hd__clkdlybuf4s50_1_150/clkdlybuf4s50_1
rlabel metal1 5559 -11484 6295 -11388 1 sky130_fd_sc_hd__clkdlybuf4s50_1_150/VGND
rlabel metal1 5559 -10940 6295 -10844 1 sky130_fd_sc_hd__clkdlybuf4s50_1_150/VPWR
flabel metal1 5404 -11453 5438 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_189/VGND
flabel metal1 5404 -10909 5438 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_189/VPWR
flabel nwell 5404 -10909 5438 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_189/VPB
flabel pwell 5404 -11453 5438 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_189/VNB
rlabel comment 5467 -11436 5467 -11436 6 sky130_fd_sc_hd__decap_4_189/decap_4
rlabel metal1 5099 -11484 5467 -11388 1 sky130_fd_sc_hd__decap_4_189/VGND
rlabel metal1 5099 -10940 5467 -10844 1 sky130_fd_sc_hd__decap_4_189/VPWR
flabel metal1 6692 -11453 6726 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_190/VGND
flabel metal1 6692 -10909 6726 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_190/VPWR
flabel nwell 6692 -10909 6726 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_190/VPB
flabel pwell 6692 -11453 6726 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_190/VNB
rlabel comment 6755 -11436 6755 -11436 6 sky130_fd_sc_hd__decap_4_190/decap_4
rlabel metal1 6387 -11484 6755 -11388 1 sky130_fd_sc_hd__decap_4_190/VGND
rlabel metal1 6387 -10940 6755 -10844 1 sky130_fd_sc_hd__decap_4_190/VPWR
flabel metal1 5024 -10912 5077 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_379/VPWR
flabel metal1 5027 -11454 5078 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_379/VGND
rlabel comment 5099 -11436 5099 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_379/tapvpwrvgnd_1
rlabel metal1 5007 -11484 5099 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_379/VGND
rlabel metal1 5007 -10940 5099 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_379/VPWR
flabel metal1 5484 -10912 5537 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_380/VPWR
flabel metal1 5487 -11454 5538 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_380/VGND
rlabel comment 5559 -11436 5559 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_380/tapvpwrvgnd_1
rlabel metal1 5467 -11484 5559 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_380/VGND
rlabel metal1 5467 -10940 5559 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_380/VPWR
flabel metal1 6312 -10912 6365 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_381/VPWR
flabel metal1 6315 -11454 6366 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_381/VGND
rlabel comment 6387 -11436 6387 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_381/tapvpwrvgnd_1
rlabel metal1 6295 -11484 6387 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_381/VGND
rlabel metal1 6295 -10940 6387 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_381/VPWR
flabel locali 8807 -11215 8841 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/A
flabel locali 8161 -11011 8195 -10977 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X
flabel locali 8161 -11079 8195 -11045 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X
flabel locali 8161 -11147 8195 -11113 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X
flabel locali 8161 -11215 8195 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X
flabel locali 8161 -11283 8195 -11249 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X
flabel locali 8161 -11351 8195 -11317 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X
flabel pwell 8807 -11453 8841 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/VNB
flabel nwell 8807 -10909 8841 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/VPB
flabel metal1 8807 -11453 8841 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/VGND
flabel metal1 8807 -10909 8841 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_154/VPWR
rlabel comment 8871 -11436 8871 -11436 6 sky130_fd_sc_hd__clkdlybuf4s50_1_154/clkdlybuf4s50_1
rlabel metal1 8135 -11484 8871 -11388 1 sky130_fd_sc_hd__clkdlybuf4s50_1_154/VGND
rlabel metal1 8135 -10940 8871 -10844 1 sky130_fd_sc_hd__clkdlybuf4s50_1_154/VPWR
flabel metal1 7980 -11453 8014 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_192/VGND
flabel metal1 7980 -10909 8014 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_192/VPWR
flabel nwell 7980 -10909 8014 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_192/VPB
flabel pwell 7980 -11453 8014 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_192/VNB
rlabel comment 8043 -11436 8043 -11436 6 sky130_fd_sc_hd__decap_4_192/decap_4
rlabel metal1 7675 -11484 8043 -11388 1 sky130_fd_sc_hd__decap_4_192/VGND
rlabel metal1 7675 -10940 8043 -10844 1 sky130_fd_sc_hd__decap_4_192/VPWR
flabel metal1 6876 -10909 6910 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_156/VPWR
flabel metal1 6876 -11453 6910 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_156/VGND
flabel nwell 6876 -10909 6910 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_156/VPB
flabel pwell 6876 -11453 6910 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_156/VNB
rlabel comment 6847 -11436 6847 -11436 4 sky130_fd_sc_hd__decap_8_156/decap_8
rlabel metal1 6847 -11484 7583 -11388 1 sky130_fd_sc_hd__decap_8_156/VGND
rlabel metal1 6847 -10940 7583 -10844 1 sky130_fd_sc_hd__decap_8_156/VPWR
flabel metal1 6772 -10912 6825 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_385/VPWR
flabel metal1 6775 -11454 6826 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_385/VGND
rlabel comment 6847 -11436 6847 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_385/tapvpwrvgnd_1
rlabel metal1 6755 -11484 6847 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_385/VGND
rlabel metal1 6755 -10940 6847 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_385/VPWR
flabel metal1 7600 -10912 7653 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_386/VPWR
flabel metal1 7603 -11454 7654 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_386/VGND
rlabel comment 7675 -11436 7675 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_386/tapvpwrvgnd_1
rlabel metal1 7583 -11484 7675 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_386/VGND
rlabel metal1 7583 -10940 7675 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_386/VPWR
flabel metal1 8060 -10912 8113 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_387/VPWR
flabel metal1 8063 -11454 8114 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_387/VGND
rlabel comment 8135 -11436 8135 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_387/tapvpwrvgnd_1
rlabel metal1 8043 -11484 8135 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_387/VGND
rlabel metal1 8043 -10940 8135 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_387/VPWR
flabel metal1 9268 -11453 9302 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_194/VGND
flabel metal1 9268 -10909 9302 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_194/VPWR
flabel nwell 9268 -10909 9302 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_194/VPB
flabel pwell 9268 -11453 9302 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_194/VNB
rlabel comment 9331 -11436 9331 -11436 6 sky130_fd_sc_hd__decap_4_194/decap_4
rlabel metal1 8963 -11484 9331 -11388 1 sky130_fd_sc_hd__decap_4_194/VGND
rlabel metal1 8963 -10940 9331 -10844 1 sky130_fd_sc_hd__decap_4_194/VPWR
flabel metal1 10648 -11453 10682 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_197/VGND
flabel metal1 10648 -10909 10682 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_197/VPWR
flabel nwell 10648 -10909 10682 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_197/VPB
flabel pwell 10648 -11453 10682 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_197/VNB
rlabel comment 10711 -11436 10711 -11436 6 sky130_fd_sc_hd__decap_4_197/decap_4
rlabel metal1 10343 -11484 10711 -11388 1 sky130_fd_sc_hd__decap_4_197/VGND
rlabel metal1 10343 -10940 10711 -10844 1 sky130_fd_sc_hd__decap_4_197/VPWR
flabel metal1 9452 -10909 9486 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_165/VPWR
flabel metal1 9452 -11453 9486 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_165/VGND
flabel nwell 9452 -10909 9486 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_165/VPB
flabel pwell 9452 -11453 9486 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_165/VNB
rlabel comment 9423 -11436 9423 -11436 4 sky130_fd_sc_hd__decap_8_165/decap_8
rlabel metal1 9423 -11484 10159 -11388 1 sky130_fd_sc_hd__decap_8_165/VGND
rlabel metal1 9423 -10940 10159 -10844 1 sky130_fd_sc_hd__decap_8_165/VPWR
flabel metal1 10285 -10909 10321 -10879 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_52/VPWR
flabel metal1 10285 -11449 10321 -11420 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_52/VGND
flabel nwell 10292 -10902 10312 -10885 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_52/VPB
flabel pwell 10291 -11447 10315 -11425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_52/VNB
rlabel comment 10343 -11436 10343 -11436 6 sky130_fd_sc_hd__fill_1_52/fill_1
rlabel metal1 10251 -11484 10343 -11388 1 sky130_fd_sc_hd__fill_1_52/VGND
rlabel metal1 10251 -10940 10343 -10844 1 sky130_fd_sc_hd__fill_1_52/VPWR
flabel metal1 8888 -10912 8941 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_391/VPWR
flabel metal1 8891 -11454 8942 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_391/VGND
rlabel comment 8963 -11436 8963 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_391/tapvpwrvgnd_1
rlabel metal1 8871 -11484 8963 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_391/VGND
rlabel metal1 8871 -10940 8963 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_391/VPWR
flabel metal1 9348 -10912 9401 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_392/VPWR
flabel metal1 9351 -11454 9402 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_392/VGND
rlabel comment 9423 -11436 9423 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_392/tapvpwrvgnd_1
rlabel metal1 9331 -11484 9423 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_392/VGND
rlabel metal1 9331 -10940 9423 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_392/VPWR
flabel metal1 10176 -10912 10229 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_393/VPWR
flabel metal1 10179 -11454 10230 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_393/VGND
rlabel comment 10251 -11436 10251 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_393/tapvpwrvgnd_1
rlabel metal1 10159 -11484 10251 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_393/VGND
rlabel metal1 10159 -10940 10251 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_393/VPWR
flabel locali 11383 -11215 11417 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A
flabel locali 10737 -11011 10771 -10977 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X
flabel locali 10737 -11079 10771 -11045 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X
flabel locali 10737 -11147 10771 -11113 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X
flabel locali 10737 -11215 10771 -11181 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X
flabel locali 10737 -11283 10771 -11249 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X
flabel locali 10737 -11351 10771 -11317 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X
flabel pwell 11383 -11453 11417 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/VNB
flabel nwell 11383 -10909 11417 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/VPB
flabel metal1 11383 -11453 11417 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/VGND
flabel metal1 11383 -10909 11417 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_158/VPWR
rlabel comment 11447 -11436 11447 -11436 6 sky130_fd_sc_hd__clkdlybuf4s50_1_158/clkdlybuf4s50_1
rlabel metal1 10711 -11484 11447 -11388 1 sky130_fd_sc_hd__clkdlybuf4s50_1_158/VGND
rlabel metal1 10711 -10940 11447 -10844 1 sky130_fd_sc_hd__clkdlybuf4s50_1_158/VPWR
flabel metal1 11936 -11453 11970 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_198/VGND
flabel metal1 11936 -10909 11970 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_198/VPWR
flabel nwell 11936 -10909 11970 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_198/VPB
flabel pwell 11936 -11453 11970 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_198/VNB
rlabel comment 11999 -11436 11999 -11436 6 sky130_fd_sc_hd__decap_4_198/decap_4
rlabel metal1 11631 -11484 11999 -11388 1 sky130_fd_sc_hd__decap_4_198/VGND
rlabel metal1 11631 -10940 11999 -10844 1 sky130_fd_sc_hd__decap_4_198/VPWR
flabel metal1 10653 -10909 10689 -10879 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_55/VPWR
flabel metal1 10653 -11449 10689 -11420 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_55/VGND
flabel nwell 10660 -10902 10680 -10885 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_55/VPB
flabel pwell 10659 -11447 10683 -11425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_55/VNB
rlabel comment 10711 -11436 10711 -11436 6 sky130_fd_sc_hd__fill_1_55/fill_1
rlabel metal1 10619 -11484 10711 -11388 1 sky130_fd_sc_hd__fill_1_55/VGND
rlabel metal1 10619 -10940 10711 -10844 1 sky130_fd_sc_hd__fill_1_55/VPWR
flabel metal1 11573 -10909 11609 -10879 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_56/VPWR
flabel metal1 11573 -11449 11609 -11420 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_56/VGND
flabel nwell 11580 -10902 11600 -10885 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_56/VPB
flabel pwell 11579 -11447 11603 -11425 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_56/VNB
rlabel comment 11631 -11436 11631 -11436 6 sky130_fd_sc_hd__fill_1_56/fill_1
rlabel metal1 11539 -11484 11631 -11388 1 sky130_fd_sc_hd__fill_1_56/VGND
rlabel metal1 11539 -10940 11631 -10844 1 sky130_fd_sc_hd__fill_1_56/VPWR
flabel metal1 12668 -11456 12700 -11426 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_26/VGND
flabel metal1 12668 -10913 12706 -10881 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_26/VPWR
flabel nwell 12658 -10914 12715 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_26/VPB
flabel pwell 12665 -11460 12709 -11426 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_26/VNB
rlabel comment 12735 -11436 12735 -11436 6 sky130_fd_sc_hd__fill_8_26/fill_8
rlabel metal1 11999 -11484 12735 -11388 1 sky130_fd_sc_hd__fill_8_26/VGND
rlabel metal1 11999 -10940 12735 -10844 1 sky130_fd_sc_hd__fill_8_26/VPWR
flabel metal1 11464 -10912 11517 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_395/VPWR
flabel metal1 11467 -11454 11518 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_395/VGND
rlabel comment 11539 -11436 11539 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_395/tapvpwrvgnd_1
rlabel metal1 11447 -11484 11539 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_395/VGND
rlabel metal1 11447 -10940 11539 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_395/VPWR
flabel metal1 14604 -11453 14638 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_26/VGND
flabel metal1 14604 -10909 14638 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_26/VPWR
flabel nwell 14604 -10909 14638 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_26/VPB
flabel pwell 14604 -11453 14638 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_26/VNB
rlabel comment 14667 -11436 14667 -11436 6 sky130_fd_sc_hd__decap_12_26/decap_12
rlabel metal1 13563 -11484 14667 -11388 1 sky130_fd_sc_hd__decap_12_26/VGND
rlabel metal1 13563 -10940 14667 -10844 1 sky130_fd_sc_hd__decap_12_26/VPWR
flabel metal1 13404 -11456 13436 -11426 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_28/VGND
flabel metal1 13404 -10913 13442 -10881 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_28/VPWR
flabel nwell 13394 -10914 13451 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_28/VPB
flabel pwell 13401 -11460 13445 -11426 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_28/VNB
rlabel comment 13471 -11436 13471 -11436 6 sky130_fd_sc_hd__fill_8_28/fill_8
rlabel metal1 12735 -11484 13471 -11388 1 sky130_fd_sc_hd__fill_8_28/VGND
rlabel metal1 12735 -10940 13471 -10844 1 sky130_fd_sc_hd__fill_8_28/VPWR
flabel metal1 13488 -10912 13541 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_397/VPWR
flabel metal1 13491 -11454 13542 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_397/VGND
rlabel comment 13563 -11436 13563 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_397/tapvpwrvgnd_1
rlabel metal1 13471 -11484 13563 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_397/VGND
rlabel metal1 13471 -10940 13563 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_397/VPWR
flabel metal1 16628 -10909 16662 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_35/VPWR
flabel metal1 16628 -11453 16662 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_35/VGND
flabel nwell 16628 -10909 16662 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_35/VPB
flabel pwell 16628 -11453 16662 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_35/VNB
rlabel comment 16691 -11436 16691 -11436 6 sky130_fd_sc_hd__decap_8_35/decap_8
rlabel metal1 15955 -11484 16691 -11388 1 sky130_fd_sc_hd__decap_8_35/VGND
rlabel metal1 15955 -10940 16691 -10844 1 sky130_fd_sc_hd__decap_8_35/VPWR
flabel metal1 15800 -11453 15834 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_28/VGND
flabel metal1 15800 -10909 15834 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_28/VPWR
flabel nwell 15800 -10909 15834 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_28/VPB
flabel pwell 15800 -11453 15834 -11419 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_28/VNB
rlabel comment 15863 -11436 15863 -11436 6 sky130_fd_sc_hd__decap_12_28/decap_12
rlabel metal1 14759 -11484 15863 -11388 1 sky130_fd_sc_hd__decap_12_28/VGND
rlabel metal1 14759 -10940 15863 -10844 1 sky130_fd_sc_hd__decap_12_28/VPWR
flabel metal1 14684 -10912 14737 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_400/VPWR
flabel metal1 14687 -11454 14738 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_400/VGND
rlabel comment 14759 -11436 14759 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_400/tapvpwrvgnd_1
rlabel metal1 14667 -11484 14759 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_400/VGND
rlabel metal1 14667 -10940 14759 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_400/VPWR
flabel metal1 15880 -10912 15933 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_401/VPWR
flabel metal1 15883 -11454 15934 -11416 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_401/VGND
rlabel comment 15955 -11436 15955 -11436 6 sky130_fd_sc_hd__tapvpwrvgnd_1_401/tapvpwrvgnd_1
rlabel metal1 15863 -11484 15955 -11388 1 sky130_fd_sc_hd__tapvpwrvgnd_1_401/VGND
rlabel metal1 15863 -10940 15955 -10844 1 sky130_fd_sc_hd__tapvpwrvgnd_1_401/VPWR
flabel metal1 -2244 -10901 -2191 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_549/VPWR
flabel metal1 -2241 -10368 -2190 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_549/VGND
rlabel comment -2169 -10348 -2169 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_549/tapvpwrvgnd_1
rlabel metal1 -2261 -10396 -2169 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_549/VGND
rlabel metal1 -2261 -10940 -2169 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_549/VPWR
flabel metal1 -2239 -9824 -2186 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_548/VPWR
flabel metal1 -2240 -10366 -2189 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_548/VGND
rlabel comment -2261 -10348 -2261 -10348 4 sky130_fd_sc_hd__tapvpwrvgnd_1_548/tapvpwrvgnd_1
rlabel metal1 -2261 -10396 -2169 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_548/VGND
rlabel metal1 -2261 -9852 -2169 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_548/VPWR
flabel metal1 -2324 -10909 -2290 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_84/VPWR
flabel metal1 -2324 -10365 -2290 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_84/VGND
flabel nwell -2324 -10909 -2290 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_84/VPB
flabel pwell -2324 -10365 -2290 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_84/VNB
rlabel comment -2261 -10348 -2261 -10348 8 sky130_fd_sc_hd__decap_8_84/decap_8
rlabel metal1 -2997 -10396 -2261 -10300 5 sky130_fd_sc_hd__decap_8_84/VGND
rlabel metal1 -2997 -10940 -2261 -10844 5 sky130_fd_sc_hd__decap_8_84/VPWR
flabel metal1 -2968 -9821 -2934 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_83/VPWR
flabel metal1 -2968 -10365 -2934 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_83/VGND
flabel nwell -2968 -9821 -2934 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_83/VPB
flabel pwell -2968 -10365 -2934 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_83/VNB
rlabel comment -2997 -10348 -2997 -10348 4 sky130_fd_sc_hd__decap_8_83/decap_8
rlabel metal1 -2997 -10396 -2261 -10300 1 sky130_fd_sc_hd__decap_8_83/VGND
rlabel metal1 -2997 -9852 -2261 -9756 1 sky130_fd_sc_hd__decap_8_83/VPWR
flabel metal1 -1692 -10901 -1639 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_525/VPWR
flabel metal1 -1689 -10368 -1638 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_525/VGND
rlabel comment -1617 -10348 -1617 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_525/tapvpwrvgnd_1
rlabel metal1 -1709 -10396 -1617 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_525/VGND
rlabel metal1 -1709 -10940 -1617 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_525/VPWR
flabel metal1 -2135 -10358 -2112 -10339 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_32/VGND
flabel metal1 -2135 -9813 -2115 -9796 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_32/VPWR
flabel nwell -2134 -9818 -2109 -9792 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_32/VPB
flabel pwell -2134 -10360 -2112 -10336 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_32/VNB
rlabel comment -2169 -10348 -2169 -10348 4 sky130_fd_sc_hd__fill_4_32/fill_4
rlabel metal1 -2169 -10396 -1801 -10300 1 sky130_fd_sc_hd__fill_4_32/VGND
rlabel metal1 -2169 -9852 -1801 -9756 1 sky130_fd_sc_hd__fill_4_32/VPWR
flabel metal1 -2058 -10366 -2005 -10334 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_23/VGND
flabel metal1 -2058 -10909 -2006 -10878 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_23/VPWR
flabel nwell -2047 -10901 -2013 -10883 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_23/VPB
flabel pwell -2048 -10360 -2016 -10338 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_23/VNB
rlabel comment -1985 -10348 -1985 -10348 8 sky130_fd_sc_hd__fill_2_23/fill_2
rlabel metal1 -2169 -10396 -1985 -10300 5 sky130_fd_sc_hd__fill_2_23/VGND
rlabel metal1 -2169 -10940 -1985 -10844 5 sky130_fd_sc_hd__fill_2_23/VPWR
flabel metal1 -1781 -10362 -1728 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_22/VGND
flabel metal1 -1780 -9818 -1728 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_22/VPWR
flabel nwell -1773 -9813 -1739 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_22/VPB
flabel pwell -1770 -10358 -1738 -10336 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_22/VNB
rlabel comment -1801 -10348 -1801 -10348 4 sky130_fd_sc_hd__fill_2_22/fill_2
rlabel metal1 -1801 -10396 -1617 -10300 1 sky130_fd_sc_hd__fill_2_22/VGND
rlabel metal1 -1801 -9852 -1617 -9756 1 sky130_fd_sc_hd__fill_2_22/VPWR
flabel metal1 -1588 -9821 -1554 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_36/VPWR
flabel metal1 -1588 -10365 -1554 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_36/VGND
flabel nwell -1588 -9821 -1554 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_36/VPB
flabel pwell -1588 -10365 -1554 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_36/VNB
rlabel comment -1617 -10348 -1617 -10348 4 sky130_fd_sc_hd__decap_8_36/decap_8
rlabel metal1 -1617 -10396 -881 -10300 1 sky130_fd_sc_hd__decap_8_36/VGND
rlabel metal1 -1617 -9852 -881 -9756 1 sky130_fd_sc_hd__decap_8_36/VPWR
flabel metal1 -944 -10909 -910 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_30/VPWR
flabel metal1 -944 -10365 -910 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_30/VGND
flabel nwell -944 -10909 -910 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_30/VPB
flabel pwell -944 -10365 -910 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_30/VNB
rlabel comment -881 -10348 -881 -10348 8 sky130_fd_sc_hd__decap_8_30/decap_8
rlabel metal1 -1617 -10396 -881 -10300 5 sky130_fd_sc_hd__decap_8_30/VGND
rlabel metal1 -1617 -10940 -881 -10844 5 sky130_fd_sc_hd__decap_8_30/VPWR
flabel locali -1772 -10535 -1738 -10501 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/Y
flabel locali -1772 -10603 -1738 -10569 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/Y
flabel locali -1864 -10671 -1830 -10637 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/Y
flabel locali -1864 -10603 -1830 -10569 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/Y
flabel locali -1864 -10535 -1830 -10501 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/Y
flabel locali -1956 -10467 -1922 -10433 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/A
flabel locali -1956 -10535 -1922 -10501 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/A
flabel locali -1956 -10603 -1922 -10569 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_6/A
flabel nwell -1956 -10909 -1922 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_6/VPB
flabel pwell -1956 -10365 -1922 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_6/VNB
flabel metal1 -1956 -10365 -1922 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_6/VGND
flabel metal1 -1956 -10909 -1922 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_6/VPWR
rlabel comment -1985 -10348 -1985 -10348 2 sky130_fd_sc_hd__clkinv_1_6/clkinv_1
rlabel metal1 -1985 -10396 -1709 -10300 5 sky130_fd_sc_hd__clkinv_1_6/VGND
rlabel metal1 -1985 -10940 -1709 -10844 5 sky130_fd_sc_hd__clkinv_1_6/VPWR
flabel metal1 -852 -9821 -818 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_37/VPWR
flabel metal1 -852 -10365 -818 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_37/VGND
flabel nwell -852 -9821 -818 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_37/VPB
flabel pwell -852 -10365 -818 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_37/VNB
rlabel comment -881 -10348 -881 -10348 4 sky130_fd_sc_hd__decap_8_37/decap_8
rlabel metal1 -881 -10396 -145 -10300 1 sky130_fd_sc_hd__decap_8_37/VGND
rlabel metal1 -881 -9852 -145 -9756 1 sky130_fd_sc_hd__decap_8_37/VPWR
flabel metal1 -208 -10909 -174 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_32/VPWR
flabel metal1 -208 -10365 -174 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_32/VGND
flabel nwell -208 -10909 -174 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_32/VPB
flabel pwell -208 -10365 -174 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_32/VNB
rlabel comment -145 -10348 -145 -10348 8 sky130_fd_sc_hd__decap_8_32/decap_8
rlabel metal1 -881 -10396 -145 -10300 5 sky130_fd_sc_hd__decap_8_32/VGND
rlabel metal1 -881 -10940 -145 -10844 5 sky130_fd_sc_hd__decap_8_32/VPWR
flabel metal1 332 -9824 385 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_403/VPWR
flabel metal1 335 -10366 386 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_403/VGND
rlabel comment 407 -10348 407 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_403/tapvpwrvgnd_1
rlabel metal1 315 -10396 407 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_403/VGND
rlabel metal1 315 -9852 407 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_403/VPWR
flabel metal1 -128 -9824 -75 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_402/VPWR
flabel metal1 -125 -10366 -74 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_402/VGND
rlabel comment -53 -10348 -53 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_402/tapvpwrvgnd_1
rlabel metal1 -145 -10396 -53 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_402/VGND
rlabel metal1 -145 -9852 -53 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_402/VPWR
flabel metal1 -128 -10901 -75 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_361/VPWR
flabel metal1 -125 -10368 -74 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_361/VGND
rlabel comment -53 -10348 -53 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_361/tapvpwrvgnd_1
rlabel metal1 -145 -10396 -53 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_361/VGND
rlabel metal1 -145 -10940 -53 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_361/VPWR
flabel metal1 332 -10901 385 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_360/VPWR
flabel metal1 335 -10368 386 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_360/VGND
rlabel comment 407 -10348 407 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_360/tapvpwrvgnd_1
rlabel metal1 315 -10396 407 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_360/VGND
rlabel metal1 315 -10940 407 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_360/VPWR
flabel metal1 252 -10365 286 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_199/VGND
flabel metal1 252 -9821 286 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_199/VPWR
flabel nwell 252 -9821 286 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_199/VPB
flabel pwell 252 -10365 286 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_199/VNB
rlabel comment 315 -10348 315 -10348 6 sky130_fd_sc_hd__decap_4_199/decap_4
rlabel metal1 -53 -10396 315 -10300 1 sky130_fd_sc_hd__decap_4_199/VGND
rlabel metal1 -53 -9852 315 -9756 1 sky130_fd_sc_hd__decap_4_199/VPWR
flabel metal1 252 -10365 286 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_179/VGND
flabel metal1 252 -10909 286 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_179/VPWR
flabel nwell 252 -10909 286 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_179/VPB
flabel pwell 252 -10365 286 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_179/VNB
rlabel comment 315 -10348 315 -10348 8 sky130_fd_sc_hd__decap_4_179/decap_4
rlabel metal1 -53 -10396 315 -10300 5 sky130_fd_sc_hd__decap_4_179/VGND
rlabel metal1 -53 -10940 315 -10844 5 sky130_fd_sc_hd__decap_4_179/VPWR
flabel locali 437 -10127 471 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/A
flabel locali 1083 -9923 1117 -9889 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/X
flabel locali 1083 -9991 1117 -9957 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/X
flabel locali 1083 -10059 1117 -10025 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/X
flabel locali 1083 -10127 1117 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/X
flabel locali 1083 -10195 1117 -10161 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/X
flabel locali 1083 -10263 1117 -10229 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/X
flabel pwell 437 -10365 471 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/VNB
flabel nwell 437 -9821 471 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/VPB
flabel metal1 437 -10365 471 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/VGND
flabel metal1 437 -9821 471 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_159/VPWR
rlabel comment 407 -10348 407 -10348 4 sky130_fd_sc_hd__clkdlybuf4s50_1_159/clkdlybuf4s50_1
rlabel metal1 407 -10396 1143 -10300 1 sky130_fd_sc_hd__clkdlybuf4s50_1_159/VGND
rlabel metal1 407 -9852 1143 -9756 1 sky130_fd_sc_hd__clkdlybuf4s50_1_159/VPWR
flabel locali 1079 -10603 1113 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/A
flabel locali 433 -10807 467 -10773 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/X
flabel locali 433 -10739 467 -10705 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/X
flabel locali 433 -10671 467 -10637 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/X
flabel locali 433 -10603 467 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/X
flabel locali 433 -10535 467 -10501 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/X
flabel locali 433 -10467 467 -10433 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/X
flabel pwell 1079 -10365 1113 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/VNB
flabel nwell 1079 -10909 1113 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/VPB
flabel metal1 1079 -10365 1113 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/VGND
flabel metal1 1079 -10909 1113 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_141/VPWR
rlabel comment 1143 -10348 1143 -10348 8 sky130_fd_sc_hd__clkdlybuf4s50_1_141/clkdlybuf4s50_1
rlabel metal1 407 -10396 1143 -10300 5 sky130_fd_sc_hd__clkdlybuf4s50_1_141/VGND
rlabel metal1 407 -10940 1143 -10844 5 sky130_fd_sc_hd__clkdlybuf4s50_1_141/VPWR
flabel metal1 1160 -9824 1213 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_406/VPWR
flabel metal1 1163 -10366 1214 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_406/VGND
rlabel comment 1235 -10348 1235 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_406/tapvpwrvgnd_1
rlabel metal1 1143 -10396 1235 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_406/VGND
rlabel metal1 1143 -9852 1235 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_406/VPWR
flabel metal1 1620 -9824 1673 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_405/VPWR
flabel metal1 1623 -10366 1674 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_405/VGND
rlabel comment 1695 -10348 1695 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_405/tapvpwrvgnd_1
rlabel metal1 1603 -10396 1695 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_405/VGND
rlabel metal1 1603 -9852 1695 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_405/VPWR
flabel metal1 1160 -10901 1213 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_365/VPWR
flabel metal1 1163 -10368 1214 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_365/VGND
rlabel comment 1235 -10348 1235 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_365/tapvpwrvgnd_1
rlabel metal1 1143 -10396 1235 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_365/VGND
rlabel metal1 1143 -10940 1235 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_365/VPWR
flabel metal1 1620 -10901 1673 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_364/VPWR
flabel metal1 1623 -10368 1674 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_364/VGND
rlabel comment 1695 -10348 1695 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_364/tapvpwrvgnd_1
rlabel metal1 1603 -10396 1695 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_364/VGND
rlabel metal1 1603 -10940 1695 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_364/VPWR
flabel metal1 1540 -10365 1574 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_201/VGND
flabel metal1 1540 -9821 1574 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_201/VPWR
flabel nwell 1540 -9821 1574 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_201/VPB
flabel pwell 1540 -10365 1574 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_201/VNB
rlabel comment 1603 -10348 1603 -10348 6 sky130_fd_sc_hd__decap_4_201/decap_4
rlabel metal1 1235 -10396 1603 -10300 1 sky130_fd_sc_hd__decap_4_201/VGND
rlabel metal1 1235 -9852 1603 -9756 1 sky130_fd_sc_hd__decap_4_201/VPWR
flabel metal1 1540 -10365 1574 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_181/VGND
flabel metal1 1540 -10909 1574 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_181/VPWR
flabel nwell 1540 -10909 1574 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_181/VPB
flabel pwell 1540 -10365 1574 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_181/VNB
rlabel comment 1603 -10348 1603 -10348 8 sky130_fd_sc_hd__decap_4_181/decap_4
rlabel metal1 1235 -10396 1603 -10300 5 sky130_fd_sc_hd__decap_4_181/VGND
rlabel metal1 1235 -10940 1603 -10844 5 sky130_fd_sc_hd__decap_4_181/VPWR
flabel metal1 2448 -9824 2501 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_404/VPWR
flabel metal1 2451 -10366 2502 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_404/VGND
rlabel comment 2523 -10348 2523 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_404/tapvpwrvgnd_1
rlabel metal1 2431 -10396 2523 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_404/VGND
rlabel metal1 2431 -9852 2523 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_404/VPWR
flabel metal1 2448 -10901 2501 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_366/VPWR
flabel metal1 2451 -10368 2502 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_366/VGND
rlabel comment 2523 -10348 2523 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_366/tapvpwrvgnd_1
rlabel metal1 2431 -10396 2523 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_366/VGND
rlabel metal1 2431 -10940 2523 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_366/VPWR
flabel metal1 2368 -10909 2402 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_135/VPWR
flabel metal1 2368 -10365 2402 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_135/VGND
flabel nwell 2368 -10909 2402 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_135/VPB
flabel pwell 2368 -10365 2402 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_135/VNB
rlabel comment 2431 -10348 2431 -10348 8 sky130_fd_sc_hd__decap_8_135/decap_8
rlabel metal1 1695 -10396 2431 -10300 5 sky130_fd_sc_hd__decap_8_135/VGND
rlabel metal1 1695 -10940 2431 -10844 5 sky130_fd_sc_hd__decap_8_135/VPWR
flabel metal1 1724 -9821 1758 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_134/VPWR
flabel metal1 1724 -10365 1758 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_134/VGND
flabel nwell 1724 -9821 1758 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_134/VPB
flabel pwell 1724 -10365 1758 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_134/VNB
rlabel comment 1695 -10348 1695 -10348 4 sky130_fd_sc_hd__decap_8_134/decap_8
rlabel metal1 1695 -10396 2431 -10300 1 sky130_fd_sc_hd__decap_8_134/VGND
rlabel metal1 1695 -9852 2431 -9756 1 sky130_fd_sc_hd__decap_8_134/VPWR
flabel metal1 2828 -10365 2862 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_200/VGND
flabel metal1 2828 -9821 2862 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_200/VPWR
flabel nwell 2828 -9821 2862 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_200/VPB
flabel pwell 2828 -10365 2862 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_200/VNB
rlabel comment 2891 -10348 2891 -10348 6 sky130_fd_sc_hd__decap_4_200/decap_4
rlabel metal1 2523 -10396 2891 -10300 1 sky130_fd_sc_hd__decap_4_200/VGND
rlabel metal1 2523 -9852 2891 -9756 1 sky130_fd_sc_hd__decap_4_200/VPWR
flabel metal1 2828 -10365 2862 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_182/VGND
flabel metal1 2828 -10909 2862 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_182/VPWR
flabel nwell 2828 -10909 2862 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_182/VPB
flabel pwell 2828 -10365 2862 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_182/VNB
rlabel comment 2891 -10348 2891 -10348 8 sky130_fd_sc_hd__decap_4_182/decap_4
rlabel metal1 2523 -10396 2891 -10300 5 sky130_fd_sc_hd__decap_4_182/VGND
rlabel metal1 2523 -10940 2891 -10844 5 sky130_fd_sc_hd__decap_4_182/VPWR
flabel metal1 2908 -9824 2961 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_409/VPWR
flabel metal1 2911 -10366 2962 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_409/VGND
rlabel comment 2983 -10348 2983 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_409/tapvpwrvgnd_1
rlabel metal1 2891 -10396 2983 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_409/VGND
rlabel metal1 2891 -9852 2983 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_409/VPWR
flabel metal1 2908 -10901 2961 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_372/VPWR
flabel metal1 2911 -10368 2962 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_372/VGND
rlabel comment 2983 -10348 2983 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_372/tapvpwrvgnd_1
rlabel metal1 2891 -10396 2983 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_372/VGND
rlabel metal1 2891 -10940 2983 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_372/VPWR
flabel locali 3013 -10127 3047 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A
flabel locali 3659 -9923 3693 -9889 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X
flabel locali 3659 -9991 3693 -9957 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X
flabel locali 3659 -10059 3693 -10025 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X
flabel locali 3659 -10127 3693 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X
flabel locali 3659 -10195 3693 -10161 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X
flabel locali 3659 -10263 3693 -10229 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X
flabel pwell 3013 -10365 3047 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/VNB
flabel nwell 3013 -9821 3047 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/VPB
flabel metal1 3013 -10365 3047 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/VGND
flabel metal1 3013 -9821 3047 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_162/VPWR
rlabel comment 2983 -10348 2983 -10348 4 sky130_fd_sc_hd__clkdlybuf4s50_1_162/clkdlybuf4s50_1
rlabel metal1 2983 -10396 3719 -10300 1 sky130_fd_sc_hd__clkdlybuf4s50_1_162/VGND
rlabel metal1 2983 -9852 3719 -9756 1 sky130_fd_sc_hd__clkdlybuf4s50_1_162/VPWR
flabel locali 3655 -10603 3689 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A
flabel locali 3009 -10807 3043 -10773 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
flabel locali 3009 -10739 3043 -10705 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
flabel locali 3009 -10671 3043 -10637 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
flabel locali 3009 -10603 3043 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
flabel locali 3009 -10535 3043 -10501 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
flabel locali 3009 -10467 3043 -10433 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
flabel pwell 3655 -10365 3689 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/VNB
flabel nwell 3655 -10909 3689 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/VPB
flabel metal1 3655 -10365 3689 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/VGND
flabel metal1 3655 -10909 3689 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_146/VPWR
rlabel comment 3719 -10348 3719 -10348 8 sky130_fd_sc_hd__clkdlybuf4s50_1_146/clkdlybuf4s50_1
rlabel metal1 2983 -10396 3719 -10300 5 sky130_fd_sc_hd__clkdlybuf4s50_1_146/VGND
rlabel metal1 2983 -10940 3719 -10844 5 sky130_fd_sc_hd__clkdlybuf4s50_1_146/VPWR
flabel metal1 4196 -9824 4249 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_408/VPWR
flabel metal1 4199 -10366 4250 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_408/VGND
rlabel comment 4271 -10348 4271 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_408/tapvpwrvgnd_1
rlabel metal1 4179 -10396 4271 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_408/VGND
rlabel metal1 4179 -9852 4271 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_408/VPWR
flabel metal1 3736 -9824 3789 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_407/VPWR
flabel metal1 3739 -10366 3790 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_407/VGND
rlabel comment 3811 -10348 3811 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_407/tapvpwrvgnd_1
rlabel metal1 3719 -10396 3811 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_407/VGND
rlabel metal1 3719 -9852 3811 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_407/VPWR
flabel metal1 3736 -10901 3789 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_371/VPWR
flabel metal1 3739 -10368 3790 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_371/VGND
rlabel comment 3811 -10348 3811 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_371/tapvpwrvgnd_1
rlabel metal1 3719 -10396 3811 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_371/VGND
rlabel metal1 3719 -10940 3811 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_371/VPWR
flabel metal1 4196 -10901 4249 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_370/VPWR
flabel metal1 4199 -10368 4250 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_370/VGND
rlabel comment 4271 -10348 4271 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_370/tapvpwrvgnd_1
rlabel metal1 4179 -10396 4271 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_370/VGND
rlabel metal1 4179 -10940 4271 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_370/VPWR
flabel metal1 4300 -9821 4334 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_148/VPWR
flabel metal1 4300 -10365 4334 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_148/VGND
flabel nwell 4300 -9821 4334 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_148/VPB
flabel pwell 4300 -10365 4334 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_148/VNB
rlabel comment 4271 -10348 4271 -10348 4 sky130_fd_sc_hd__decap_8_148/decap_8
rlabel metal1 4271 -10396 5007 -10300 1 sky130_fd_sc_hd__decap_8_148/VGND
rlabel metal1 4271 -9852 5007 -9756 1 sky130_fd_sc_hd__decap_8_148/VPWR
flabel metal1 4944 -10909 4978 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_145/VPWR
flabel metal1 4944 -10365 4978 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_145/VGND
flabel nwell 4944 -10909 4978 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_145/VPB
flabel pwell 4944 -10365 4978 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_145/VNB
rlabel comment 5007 -10348 5007 -10348 8 sky130_fd_sc_hd__decap_8_145/decap_8
rlabel metal1 4271 -10396 5007 -10300 5 sky130_fd_sc_hd__decap_8_145/VGND
rlabel metal1 4271 -10940 5007 -10844 5 sky130_fd_sc_hd__decap_8_145/VPWR
flabel metal1 4116 -10365 4150 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_202/VGND
flabel metal1 4116 -9821 4150 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_202/VPWR
flabel nwell 4116 -9821 4150 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_202/VPB
flabel pwell 4116 -10365 4150 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_202/VNB
rlabel comment 4179 -10348 4179 -10348 6 sky130_fd_sc_hd__decap_4_202/decap_4
rlabel metal1 3811 -10396 4179 -10300 1 sky130_fd_sc_hd__decap_4_202/VGND
rlabel metal1 3811 -9852 4179 -9756 1 sky130_fd_sc_hd__decap_4_202/VPWR
flabel metal1 4116 -10365 4150 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_185/VGND
flabel metal1 4116 -10909 4150 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_185/VPWR
flabel nwell 4116 -10909 4150 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_185/VPB
flabel pwell 4116 -10365 4150 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_185/VNB
rlabel comment 4179 -10348 4179 -10348 8 sky130_fd_sc_hd__decap_4_185/decap_4
rlabel metal1 3811 -10396 4179 -10300 5 sky130_fd_sc_hd__decap_4_185/VGND
rlabel metal1 3811 -10940 4179 -10844 5 sky130_fd_sc_hd__decap_4_185/VPWR
flabel metal1 5024 -9824 5077 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_412/VPWR
flabel metal1 5027 -10366 5078 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_412/VGND
rlabel comment 5099 -10348 5099 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_412/tapvpwrvgnd_1
rlabel metal1 5007 -10396 5099 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_412/VGND
rlabel metal1 5007 -9852 5099 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_412/VPWR
flabel metal1 5484 -9824 5537 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_411/VPWR
flabel metal1 5487 -10366 5538 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_411/VGND
rlabel comment 5559 -10348 5559 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_411/tapvpwrvgnd_1
rlabel metal1 5467 -10396 5559 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_411/VGND
rlabel metal1 5467 -9852 5559 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_411/VPWR
flabel metal1 5024 -10901 5077 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_378/VPWR
flabel metal1 5027 -10368 5078 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_378/VGND
rlabel comment 5099 -10348 5099 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_378/tapvpwrvgnd_1
rlabel metal1 5007 -10396 5099 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_378/VGND
rlabel metal1 5007 -10940 5099 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_378/VPWR
flabel metal1 5484 -10901 5537 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_377/VPWR
flabel metal1 5487 -10368 5538 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_377/VGND
rlabel comment 5559 -10348 5559 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_377/tapvpwrvgnd_1
rlabel metal1 5467 -10396 5559 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_377/VGND
rlabel metal1 5467 -10940 5559 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_377/VPWR
flabel metal1 5404 -10365 5438 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_204/VGND
flabel metal1 5404 -9821 5438 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_204/VPWR
flabel nwell 5404 -9821 5438 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_204/VPB
flabel pwell 5404 -10365 5438 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_204/VNB
rlabel comment 5467 -10348 5467 -10348 6 sky130_fd_sc_hd__decap_4_204/decap_4
rlabel metal1 5099 -10396 5467 -10300 1 sky130_fd_sc_hd__decap_4_204/VGND
rlabel metal1 5099 -9852 5467 -9756 1 sky130_fd_sc_hd__decap_4_204/VPWR
flabel metal1 5404 -10365 5438 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_188/VGND
flabel metal1 5404 -10909 5438 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_188/VPWR
flabel nwell 5404 -10909 5438 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_188/VPB
flabel pwell 5404 -10365 5438 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_188/VNB
rlabel comment 5467 -10348 5467 -10348 8 sky130_fd_sc_hd__decap_4_188/decap_4
rlabel metal1 5099 -10396 5467 -10300 5 sky130_fd_sc_hd__decap_4_188/VGND
rlabel metal1 5099 -10940 5467 -10844 5 sky130_fd_sc_hd__decap_4_188/VPWR
flabel metal1 6312 -9824 6365 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_410/VPWR
flabel metal1 6315 -10366 6366 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_410/VGND
rlabel comment 6387 -10348 6387 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_410/tapvpwrvgnd_1
rlabel metal1 6295 -10396 6387 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_410/VGND
rlabel metal1 6295 -9852 6387 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_410/VPWR
flabel metal1 6312 -10901 6365 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_376/VPWR
flabel metal1 6315 -10368 6366 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_376/VGND
rlabel comment 6387 -10348 6387 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_376/tapvpwrvgnd_1
rlabel metal1 6295 -10396 6387 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_376/VGND
rlabel metal1 6295 -10940 6387 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_376/VPWR
flabel locali 5589 -10127 5623 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A
flabel locali 6235 -9923 6269 -9889 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/X
flabel locali 6235 -9991 6269 -9957 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/X
flabel locali 6235 -10059 6269 -10025 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/X
flabel locali 6235 -10127 6269 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/X
flabel locali 6235 -10195 6269 -10161 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/X
flabel locali 6235 -10263 6269 -10229 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/X
flabel pwell 5589 -10365 5623 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/VNB
flabel nwell 5589 -9821 5623 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/VPB
flabel metal1 5589 -10365 5623 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/VGND
flabel metal1 5589 -9821 5623 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_163/VPWR
rlabel comment 5559 -10348 5559 -10348 4 sky130_fd_sc_hd__clkdlybuf4s50_1_163/clkdlybuf4s50_1
rlabel metal1 5559 -10396 6295 -10300 1 sky130_fd_sc_hd__clkdlybuf4s50_1_163/VGND
rlabel metal1 5559 -9852 6295 -9756 1 sky130_fd_sc_hd__clkdlybuf4s50_1_163/VPWR
flabel locali 6231 -10603 6265 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/A
flabel locali 5585 -10807 5619 -10773 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X
flabel locali 5585 -10739 5619 -10705 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X
flabel locali 5585 -10671 5619 -10637 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X
flabel locali 5585 -10603 5619 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X
flabel locali 5585 -10535 5619 -10501 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X
flabel locali 5585 -10467 5619 -10433 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X
flabel pwell 6231 -10365 6265 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/VNB
flabel nwell 6231 -10909 6265 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/VPB
flabel metal1 6231 -10365 6265 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/VGND
flabel metal1 6231 -10909 6265 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_149/VPWR
rlabel comment 6295 -10348 6295 -10348 8 sky130_fd_sc_hd__clkdlybuf4s50_1_149/clkdlybuf4s50_1
rlabel metal1 5559 -10396 6295 -10300 5 sky130_fd_sc_hd__clkdlybuf4s50_1_149/VGND
rlabel metal1 5559 -10940 6295 -10844 5 sky130_fd_sc_hd__clkdlybuf4s50_1_149/VPWR
flabel metal1 6692 -10365 6726 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_203/VGND
flabel metal1 6692 -9821 6726 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_203/VPWR
flabel nwell 6692 -9821 6726 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_203/VPB
flabel pwell 6692 -10365 6726 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_203/VNB
rlabel comment 6755 -10348 6755 -10348 6 sky130_fd_sc_hd__decap_4_203/decap_4
rlabel metal1 6387 -10396 6755 -10300 1 sky130_fd_sc_hd__decap_4_203/VGND
rlabel metal1 6387 -9852 6755 -9756 1 sky130_fd_sc_hd__decap_4_203/VPWR
flabel metal1 6692 -10365 6726 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_187/VGND
flabel metal1 6692 -10909 6726 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_187/VPWR
flabel nwell 6692 -10909 6726 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_187/VPB
flabel pwell 6692 -10365 6726 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_187/VNB
rlabel comment 6755 -10348 6755 -10348 8 sky130_fd_sc_hd__decap_4_187/decap_4
rlabel metal1 6387 -10396 6755 -10300 5 sky130_fd_sc_hd__decap_4_187/VGND
rlabel metal1 6387 -10940 6755 -10844 5 sky130_fd_sc_hd__decap_4_187/VPWR
flabel metal1 6772 -9824 6825 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_415/VPWR
flabel metal1 6775 -10366 6826 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_415/VGND
rlabel comment 6847 -10348 6847 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_415/tapvpwrvgnd_1
rlabel metal1 6755 -10396 6847 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_415/VGND
rlabel metal1 6755 -9852 6847 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_415/VPWR
flabel metal1 6772 -10901 6825 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_382/VPWR
flabel metal1 6775 -10368 6826 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_382/VGND
rlabel comment 6847 -10348 6847 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_382/tapvpwrvgnd_1
rlabel metal1 6755 -10396 6847 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_382/VGND
rlabel metal1 6755 -10940 6847 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_382/VPWR
flabel metal1 6876 -9821 6910 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_158/VPWR
flabel metal1 6876 -10365 6910 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_158/VGND
flabel nwell 6876 -9821 6910 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_158/VPB
flabel pwell 6876 -10365 6910 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_158/VNB
rlabel comment 6847 -10348 6847 -10348 4 sky130_fd_sc_hd__decap_8_158/decap_8
rlabel metal1 6847 -10396 7583 -10300 1 sky130_fd_sc_hd__decap_8_158/VGND
rlabel metal1 6847 -9852 7583 -9756 1 sky130_fd_sc_hd__decap_8_158/VPWR
flabel metal1 7520 -10909 7554 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_155/VPWR
flabel metal1 7520 -10365 7554 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_155/VGND
flabel nwell 7520 -10909 7554 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_155/VPB
flabel pwell 7520 -10365 7554 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_155/VNB
rlabel comment 7583 -10348 7583 -10348 8 sky130_fd_sc_hd__decap_8_155/decap_8
rlabel metal1 6847 -10396 7583 -10300 5 sky130_fd_sc_hd__decap_8_155/VGND
rlabel metal1 6847 -10940 7583 -10844 5 sky130_fd_sc_hd__decap_8_155/VPWR
flabel metal1 8060 -9824 8113 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_414/VPWR
flabel metal1 8063 -10366 8114 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_414/VGND
rlabel comment 8135 -10348 8135 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_414/tapvpwrvgnd_1
rlabel metal1 8043 -10396 8135 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_414/VGND
rlabel metal1 8043 -9852 8135 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_414/VPWR
flabel metal1 7600 -9824 7653 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_413/VPWR
flabel metal1 7603 -10366 7654 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_413/VGND
rlabel comment 7675 -10348 7675 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_413/tapvpwrvgnd_1
rlabel metal1 7583 -10396 7675 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_413/VGND
rlabel metal1 7583 -9852 7675 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_413/VPWR
flabel metal1 7600 -10901 7653 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_384/VPWR
flabel metal1 7603 -10368 7654 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_384/VGND
rlabel comment 7675 -10348 7675 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_384/tapvpwrvgnd_1
rlabel metal1 7583 -10396 7675 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_384/VGND
rlabel metal1 7583 -10940 7675 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_384/VPWR
flabel metal1 8060 -10901 8113 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_383/VPWR
flabel metal1 8063 -10368 8114 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_383/VGND
rlabel comment 8135 -10348 8135 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_383/tapvpwrvgnd_1
rlabel metal1 8043 -10396 8135 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_383/VGND
rlabel metal1 8043 -10940 8135 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_383/VPWR
flabel metal1 7980 -10365 8014 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_205/VGND
flabel metal1 7980 -9821 8014 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_205/VPWR
flabel nwell 7980 -9821 8014 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_205/VPB
flabel pwell 7980 -10365 8014 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_205/VNB
rlabel comment 8043 -10348 8043 -10348 6 sky130_fd_sc_hd__decap_4_205/decap_4
rlabel metal1 7675 -10396 8043 -10300 1 sky130_fd_sc_hd__decap_4_205/VGND
rlabel metal1 7675 -9852 8043 -9756 1 sky130_fd_sc_hd__decap_4_205/VPWR
flabel metal1 7980 -10365 8014 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_191/VGND
flabel metal1 7980 -10909 8014 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_191/VPWR
flabel nwell 7980 -10909 8014 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_191/VPB
flabel pwell 7980 -10365 8014 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_191/VNB
rlabel comment 8043 -10348 8043 -10348 8 sky130_fd_sc_hd__decap_4_191/decap_4
rlabel metal1 7675 -10396 8043 -10300 5 sky130_fd_sc_hd__decap_4_191/VGND
rlabel metal1 7675 -10940 8043 -10844 5 sky130_fd_sc_hd__decap_4_191/VPWR
flabel locali 8165 -10127 8199 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A
flabel locali 8811 -9923 8845 -9889 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/X
flabel locali 8811 -9991 8845 -9957 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/X
flabel locali 8811 -10059 8845 -10025 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/X
flabel locali 8811 -10127 8845 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/X
flabel locali 8811 -10195 8845 -10161 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/X
flabel locali 8811 -10263 8845 -10229 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/X
flabel pwell 8165 -10365 8199 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/VNB
flabel nwell 8165 -9821 8199 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/VPB
flabel metal1 8165 -10365 8199 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/VGND
flabel metal1 8165 -9821 8199 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_164/VPWR
rlabel comment 8135 -10348 8135 -10348 4 sky130_fd_sc_hd__clkdlybuf4s50_1_164/clkdlybuf4s50_1
rlabel metal1 8135 -10396 8871 -10300 1 sky130_fd_sc_hd__clkdlybuf4s50_1_164/VGND
rlabel metal1 8135 -9852 8871 -9756 1 sky130_fd_sc_hd__clkdlybuf4s50_1_164/VPWR
flabel locali 8807 -10603 8841 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/A
flabel locali 8161 -10807 8195 -10773 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X
flabel locali 8161 -10739 8195 -10705 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X
flabel locali 8161 -10671 8195 -10637 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X
flabel locali 8161 -10603 8195 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X
flabel locali 8161 -10535 8195 -10501 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X
flabel locali 8161 -10467 8195 -10433 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X
flabel pwell 8807 -10365 8841 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/VNB
flabel nwell 8807 -10909 8841 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/VPB
flabel metal1 8807 -10365 8841 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/VGND
flabel metal1 8807 -10909 8841 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_152/VPWR
rlabel comment 8871 -10348 8871 -10348 8 sky130_fd_sc_hd__clkdlybuf4s50_1_152/clkdlybuf4s50_1
rlabel metal1 8135 -10396 8871 -10300 5 sky130_fd_sc_hd__clkdlybuf4s50_1_152/VGND
rlabel metal1 8135 -10940 8871 -10844 5 sky130_fd_sc_hd__clkdlybuf4s50_1_152/VPWR
flabel metal1 8888 -9824 8941 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_418/VPWR
flabel metal1 8891 -10366 8942 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_418/VGND
rlabel comment 8963 -10348 8963 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_418/tapvpwrvgnd_1
rlabel metal1 8871 -10396 8963 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_418/VGND
rlabel metal1 8871 -9852 8963 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_418/VPWR
flabel metal1 8888 -10901 8941 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_388/VPWR
flabel metal1 8891 -10368 8942 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_388/VGND
rlabel comment 8963 -10348 8963 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_388/tapvpwrvgnd_1
rlabel metal1 8871 -10396 8963 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_388/VGND
rlabel metal1 8871 -10940 8963 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_388/VPWR
flabel metal1 9268 -10365 9302 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_206/VGND
flabel metal1 9268 -9821 9302 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_206/VPWR
flabel nwell 9268 -9821 9302 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_206/VPB
flabel pwell 9268 -10365 9302 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_206/VNB
rlabel comment 9331 -10348 9331 -10348 6 sky130_fd_sc_hd__decap_4_206/decap_4
rlabel metal1 8963 -10396 9331 -10300 1 sky130_fd_sc_hd__decap_4_206/VGND
rlabel metal1 8963 -9852 9331 -9756 1 sky130_fd_sc_hd__decap_4_206/VPWR
flabel metal1 9268 -10365 9302 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_193/VGND
flabel metal1 9268 -10909 9302 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_193/VPWR
flabel nwell 9268 -10909 9302 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_193/VPB
flabel pwell 9268 -10365 9302 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_193/VNB
rlabel comment 9331 -10348 9331 -10348 8 sky130_fd_sc_hd__decap_4_193/decap_4
rlabel metal1 8963 -10396 9331 -10300 5 sky130_fd_sc_hd__decap_4_193/VGND
rlabel metal1 8963 -10940 9331 -10844 5 sky130_fd_sc_hd__decap_4_193/VPWR
flabel metal1 9348 -9824 9401 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_417/VPWR
flabel metal1 9351 -10366 9402 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_417/VGND
rlabel comment 9423 -10348 9423 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_417/tapvpwrvgnd_1
rlabel metal1 9331 -10396 9423 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_417/VGND
rlabel metal1 9331 -9852 9423 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_417/VPWR
flabel metal1 9348 -10901 9401 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_389/VPWR
flabel metal1 9351 -10368 9402 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_389/VGND
rlabel comment 9423 -10348 9423 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_389/tapvpwrvgnd_1
rlabel metal1 9331 -10396 9423 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_389/VGND
rlabel metal1 9331 -10940 9423 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_389/VPWR
flabel metal1 9452 -9821 9486 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_167/VPWR
flabel metal1 9452 -10365 9486 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_167/VGND
flabel nwell 9452 -9821 9486 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_167/VPB
flabel pwell 9452 -10365 9486 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_167/VNB
rlabel comment 9423 -10348 9423 -10348 4 sky130_fd_sc_hd__decap_8_167/decap_8
rlabel metal1 9423 -10396 10159 -10300 1 sky130_fd_sc_hd__decap_8_167/VGND
rlabel metal1 9423 -9852 10159 -9756 1 sky130_fd_sc_hd__decap_8_167/VPWR
flabel metal1 10096 -10909 10130 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_166/VPWR
flabel metal1 10096 -10365 10130 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_166/VGND
flabel nwell 10096 -10909 10130 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_166/VPB
flabel pwell 10096 -10365 10130 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_166/VNB
rlabel comment 10159 -10348 10159 -10348 8 sky130_fd_sc_hd__decap_8_166/decap_8
rlabel metal1 9423 -10396 10159 -10300 5 sky130_fd_sc_hd__decap_8_166/VGND
rlabel metal1 9423 -10940 10159 -10844 5 sky130_fd_sc_hd__decap_8_166/VPWR
flabel metal1 10176 -9824 10229 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_416/VPWR
flabel metal1 10179 -10366 10230 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_416/VGND
rlabel comment 10251 -10348 10251 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_416/tapvpwrvgnd_1
rlabel metal1 10159 -10396 10251 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_416/VGND
rlabel metal1 10159 -9852 10251 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_416/VPWR
flabel metal1 10176 -10901 10229 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_390/VPWR
flabel metal1 10179 -10368 10230 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_390/VGND
rlabel comment 10251 -10348 10251 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_390/tapvpwrvgnd_1
rlabel metal1 10159 -10396 10251 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_390/VGND
rlabel metal1 10159 -10940 10251 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_390/VPWR
flabel metal1 10285 -9821 10321 -9791 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_57/VPWR
flabel metal1 10285 -10361 10321 -10332 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_57/VGND
flabel nwell 10292 -9814 10312 -9797 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_57/VPB
flabel pwell 10291 -10359 10315 -10337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_57/VNB
rlabel comment 10343 -10348 10343 -10348 6 sky130_fd_sc_hd__fill_1_57/fill_1
rlabel metal1 10251 -10396 10343 -10300 1 sky130_fd_sc_hd__fill_1_57/VGND
rlabel metal1 10251 -9852 10343 -9756 1 sky130_fd_sc_hd__fill_1_57/VPWR
flabel metal1 10285 -10905 10321 -10875 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_51/VPWR
flabel metal1 10285 -10364 10321 -10335 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_51/VGND
flabel nwell 10292 -10899 10312 -10882 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_51/VPB
flabel pwell 10291 -10359 10315 -10337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_51/VNB
rlabel comment 10343 -10348 10343 -10348 8 sky130_fd_sc_hd__fill_1_51/fill_1
rlabel metal1 10251 -10396 10343 -10300 5 sky130_fd_sc_hd__fill_1_51/VGND
rlabel metal1 10251 -10940 10343 -10844 5 sky130_fd_sc_hd__fill_1_51/VPWR
flabel metal1 10648 -10365 10682 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_208/VGND
flabel metal1 10648 -9821 10682 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_208/VPWR
flabel nwell 10648 -9821 10682 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_208/VPB
flabel pwell 10648 -10365 10682 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_208/VNB
rlabel comment 10711 -10348 10711 -10348 6 sky130_fd_sc_hd__decap_4_208/decap_4
rlabel metal1 10343 -10396 10711 -10300 1 sky130_fd_sc_hd__decap_4_208/VGND
rlabel metal1 10343 -9852 10711 -9756 1 sky130_fd_sc_hd__decap_4_208/VPWR
flabel metal1 10648 -10365 10682 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_196/VGND
flabel metal1 10648 -10909 10682 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_196/VPWR
flabel nwell 10648 -10909 10682 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_196/VPB
flabel pwell 10648 -10365 10682 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_196/VNB
rlabel comment 10711 -10348 10711 -10348 8 sky130_fd_sc_hd__decap_4_196/decap_4
rlabel metal1 10343 -10396 10711 -10300 5 sky130_fd_sc_hd__decap_4_196/VGND
rlabel metal1 10343 -10940 10711 -10844 5 sky130_fd_sc_hd__decap_4_196/VPWR
flabel metal1 10653 -9821 10689 -9791 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_59/VPWR
flabel metal1 10653 -10361 10689 -10332 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_59/VGND
flabel nwell 10660 -9814 10680 -9797 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_59/VPB
flabel pwell 10659 -10359 10683 -10337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_59/VNB
rlabel comment 10711 -10348 10711 -10348 6 sky130_fd_sc_hd__fill_1_59/fill_1
rlabel metal1 10619 -10396 10711 -10300 1 sky130_fd_sc_hd__fill_1_59/VGND
rlabel metal1 10619 -9852 10711 -9756 1 sky130_fd_sc_hd__fill_1_59/VPWR
flabel metal1 10653 -10905 10689 -10875 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_54/VPWR
flabel metal1 10653 -10364 10689 -10335 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_54/VGND
flabel nwell 10660 -10899 10680 -10882 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_54/VPB
flabel pwell 10659 -10359 10683 -10337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_54/VNB
rlabel comment 10711 -10348 10711 -10348 8 sky130_fd_sc_hd__fill_1_54/fill_1
rlabel metal1 10619 -10396 10711 -10300 5 sky130_fd_sc_hd__fill_1_54/VGND
rlabel metal1 10619 -10940 10711 -10844 5 sky130_fd_sc_hd__fill_1_54/VPWR
flabel locali 10741 -10127 10775 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A
flabel locali 11387 -9923 11421 -9889 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
flabel locali 11387 -9991 11421 -9957 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
flabel locali 11387 -10059 11421 -10025 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
flabel locali 11387 -10127 11421 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
flabel locali 11387 -10195 11421 -10161 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
flabel locali 11387 -10263 11421 -10229 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
flabel pwell 10741 -10365 10775 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/VNB
flabel nwell 10741 -9821 10775 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/VPB
flabel metal1 10741 -10365 10775 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/VGND
flabel metal1 10741 -9821 10775 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_167/VPWR
rlabel comment 10711 -10348 10711 -10348 4 sky130_fd_sc_hd__clkdlybuf4s50_1_167/clkdlybuf4s50_1
rlabel metal1 10711 -10396 11447 -10300 1 sky130_fd_sc_hd__clkdlybuf4s50_1_167/VGND
rlabel metal1 10711 -9852 11447 -9756 1 sky130_fd_sc_hd__clkdlybuf4s50_1_167/VPWR
flabel locali 11383 -10603 11417 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/A
flabel locali 10737 -10807 10771 -10773 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X
flabel locali 10737 -10739 10771 -10705 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X
flabel locali 10737 -10671 10771 -10637 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X
flabel locali 10737 -10603 10771 -10569 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X
flabel locali 10737 -10535 10771 -10501 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X
flabel locali 10737 -10467 10771 -10433 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X
flabel pwell 11383 -10365 11417 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/VNB
flabel nwell 11383 -10909 11417 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/VPB
flabel metal1 11383 -10365 11417 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/VGND
flabel metal1 11383 -10909 11417 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_157/VPWR
rlabel comment 11447 -10348 11447 -10348 8 sky130_fd_sc_hd__clkdlybuf4s50_1_157/clkdlybuf4s50_1
rlabel metal1 10711 -10396 11447 -10300 5 sky130_fd_sc_hd__clkdlybuf4s50_1_157/VGND
rlabel metal1 10711 -10940 11447 -10844 5 sky130_fd_sc_hd__clkdlybuf4s50_1_157/VPWR
flabel metal1 11464 -9824 11517 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_419/VPWR
flabel metal1 11467 -10366 11518 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_419/VGND
rlabel comment 11539 -10348 11539 -10348 6 sky130_fd_sc_hd__tapvpwrvgnd_1_419/tapvpwrvgnd_1
rlabel metal1 11447 -10396 11539 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_419/VGND
rlabel metal1 11447 -9852 11539 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_419/VPWR
flabel metal1 11464 -10901 11517 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_394/VPWR
flabel metal1 11467 -10368 11518 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_394/VGND
rlabel comment 11539 -10348 11539 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_394/tapvpwrvgnd_1
rlabel metal1 11447 -10396 11539 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_394/VGND
rlabel metal1 11447 -10940 11539 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_394/VPWR
flabel metal1 12668 -10358 12700 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_25/VGND
flabel metal1 12668 -10903 12706 -10871 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_25/VPWR
flabel nwell 12658 -10901 12715 -10870 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_25/VPB
flabel pwell 12665 -10358 12709 -10324 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_25/VNB
rlabel comment 12735 -10348 12735 -10348 8 sky130_fd_sc_hd__fill_8_25/fill_8
rlabel metal1 11999 -10396 12735 -10300 5 sky130_fd_sc_hd__fill_8_25/VGND
rlabel metal1 11999 -10940 12735 -10844 5 sky130_fd_sc_hd__fill_8_25/VPWR
flabel metal1 12033 -10358 12056 -10339 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_12/VGND
flabel metal1 12033 -9813 12053 -9796 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_12/VPWR
flabel nwell 12034 -9818 12059 -9792 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_12/VPB
flabel pwell 12034 -10360 12056 -10336 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_12/VNB
rlabel comment 11999 -10348 11999 -10348 4 sky130_fd_sc_hd__fill_4_12/fill_4
rlabel metal1 11999 -10396 12367 -10300 1 sky130_fd_sc_hd__fill_4_12/VGND
rlabel metal1 11999 -9852 12367 -9756 1 sky130_fd_sc_hd__fill_4_12/VPWR
flabel metal1 11573 -9821 11609 -9791 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_58/VPWR
flabel metal1 11573 -10361 11609 -10332 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_58/VGND
flabel nwell 11580 -9814 11600 -9797 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_58/VPB
flabel pwell 11579 -10359 11603 -10337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_58/VNB
rlabel comment 11631 -10348 11631 -10348 6 sky130_fd_sc_hd__fill_1_58/fill_1
rlabel metal1 11539 -10396 11631 -10300 1 sky130_fd_sc_hd__fill_1_58/VGND
rlabel metal1 11539 -9852 11631 -9756 1 sky130_fd_sc_hd__fill_1_58/VPWR
flabel metal1 11573 -10905 11609 -10875 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_53/VPWR
flabel metal1 11573 -10364 11609 -10335 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_53/VGND
flabel nwell 11580 -10899 11600 -10882 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_53/VPB
flabel pwell 11579 -10359 11603 -10337 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_53/VNB
rlabel comment 11631 -10348 11631 -10348 8 sky130_fd_sc_hd__fill_1_53/fill_1
rlabel metal1 11539 -10396 11631 -10300 5 sky130_fd_sc_hd__fill_1_53/VGND
rlabel metal1 11539 -10940 11631 -10844 5 sky130_fd_sc_hd__fill_1_53/VPWR
flabel metal1 11936 -10365 11970 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_207/VGND
flabel metal1 11936 -9821 11970 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_207/VPWR
flabel nwell 11936 -9821 11970 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_207/VPB
flabel pwell 11936 -10365 11970 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_207/VNB
rlabel comment 11999 -10348 11999 -10348 6 sky130_fd_sc_hd__decap_4_207/decap_4
rlabel metal1 11631 -10396 11999 -10300 1 sky130_fd_sc_hd__decap_4_207/VGND
rlabel metal1 11631 -9852 11999 -9756 1 sky130_fd_sc_hd__decap_4_207/VPWR
flabel metal1 11936 -10365 11970 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_195/VGND
flabel metal1 11936 -10909 11970 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_195/VPWR
flabel nwell 11936 -10909 11970 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_195/VPB
flabel pwell 11936 -10365 11970 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_195/VNB
rlabel comment 11999 -10348 11999 -10348 8 sky130_fd_sc_hd__decap_4_195/decap_4
rlabel metal1 11631 -10396 11999 -10300 5 sky130_fd_sc_hd__decap_4_195/VGND
rlabel metal1 11631 -10940 11999 -10844 5 sky130_fd_sc_hd__decap_4_195/VPWR
flabel locali 15248 -10059 15282 -10025 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/X
flabel locali 15340 -10059 15374 -10025 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/X
flabel locali 15340 -10127 15374 -10093 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/X
flabel locali 15248 -10127 15282 -10093 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/X
flabel locali 15248 -10195 15282 -10161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/X
flabel locali 15340 -10195 15374 -10161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/X
flabel locali 13684 -10195 13718 -10161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/A
flabel locali 13684 -10127 13718 -10093 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/A
flabel pwell 13684 -10365 13718 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/VNB
flabel pwell 13701 -10348 13701 -10348 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/VNB
flabel nwell 13684 -9821 13718 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/VPB
flabel nwell 13701 -9804 13701 -9804 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/VPB
flabel metal1 13684 -10365 13718 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/VGND
flabel metal1 13684 -9821 13718 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_12/VPWR
rlabel comment 13655 -10348 13655 -10348 4 sky130_fd_sc_hd__clkbuf_16_12/clkbuf_16
rlabel metal1 13655 -10396 15495 -10300 1 sky130_fd_sc_hd__clkbuf_16_12/VGND
rlabel metal1 13655 -9852 15495 -9756 1 sky130_fd_sc_hd__clkbuf_16_12/VPWR
flabel locali 12672 -10127 12706 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/A
flabel locali 12764 -10127 12798 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/A
flabel locali 13040 -10195 13074 -10161 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/Y
flabel locali 12580 -10127 12614 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/A
flabel locali 13040 -10059 13074 -10025 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/Y
flabel locali 12948 -10127 12982 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/A
flabel locali 12856 -10127 12890 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/A
flabel locali 13040 -10127 13074 -10093 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_9/Y
flabel pwell 12488 -10365 12522 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_9/VNB
flabel nwell 12488 -9821 12522 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_9/VPB
flabel metal1 12488 -9821 12522 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_9/VPWR
flabel metal1 12488 -10365 12522 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_9/VGND
rlabel comment 12459 -10348 12459 -10348 4 sky130_fd_sc_hd__clkinv_4_9/clkinv_4
rlabel metal1 12459 -10396 13103 -10300 1 sky130_fd_sc_hd__clkinv_4_9/VGND
rlabel metal1 12459 -9852 13103 -9756 1 sky130_fd_sc_hd__clkinv_4_9/VPWR
flabel metal1 13224 -10365 13258 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_209/VGND
flabel metal1 13224 -9821 13258 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_209/VPWR
flabel nwell 13224 -9821 13258 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_209/VPB
flabel pwell 13224 -10365 13258 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_209/VNB
rlabel comment 13195 -10348 13195 -10348 4 sky130_fd_sc_hd__decap_4_209/decap_4
rlabel metal1 13195 -10396 13563 -10300 1 sky130_fd_sc_hd__decap_4_209/VGND
rlabel metal1 13195 -9852 13563 -9756 1 sky130_fd_sc_hd__decap_4_209/VPWR
flabel metal1 14604 -10365 14638 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_25/VGND
flabel metal1 14604 -10909 14638 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_25/VPWR
flabel nwell 14604 -10909 14638 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_25/VPB
flabel pwell 14604 -10365 14638 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_25/VNB
rlabel comment 14667 -10348 14667 -10348 8 sky130_fd_sc_hd__decap_12_25/decap_12
rlabel metal1 13563 -10396 14667 -10300 5 sky130_fd_sc_hd__decap_12_25/VGND
rlabel metal1 13563 -10940 14667 -10844 5 sky130_fd_sc_hd__decap_12_25/VPWR
flabel metal1 13404 -10358 13436 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_27/VGND
flabel metal1 13404 -10903 13442 -10871 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_27/VPWR
flabel nwell 13394 -10901 13451 -10870 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_27/VPB
flabel pwell 13401 -10358 13445 -10324 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_27/VNB
rlabel comment 13471 -10348 13471 -10348 8 sky130_fd_sc_hd__fill_8_27/fill_8
rlabel metal1 12735 -10396 13471 -10300 5 sky130_fd_sc_hd__fill_8_27/VGND
rlabel metal1 12735 -10940 13471 -10844 5 sky130_fd_sc_hd__fill_8_27/VPWR
flabel metal1 13488 -10901 13541 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_396/VPWR
flabel metal1 13491 -10368 13542 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_396/VGND
rlabel comment 13563 -10348 13563 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_396/tapvpwrvgnd_1
rlabel metal1 13471 -10396 13563 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_396/VGND
rlabel metal1 13471 -10940 13563 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_396/VPWR
flabel metal1 13585 -9824 13638 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_420/VPWR
flabel metal1 13584 -10366 13635 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_420/VGND
rlabel comment 13563 -10348 13563 -10348 4 sky130_fd_sc_hd__tapvpwrvgnd_1_420/tapvpwrvgnd_1
rlabel metal1 13563 -10396 13655 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_420/VGND
rlabel metal1 13563 -9852 13655 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_420/VPWR
flabel metal1 13125 -9824 13178 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_421/VPWR
flabel metal1 13124 -10366 13175 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_421/VGND
rlabel comment 13103 -10348 13103 -10348 4 sky130_fd_sc_hd__tapvpwrvgnd_1_421/tapvpwrvgnd_1
rlabel metal1 13103 -10396 13195 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_421/VGND
rlabel metal1 13103 -9852 13195 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_421/VPWR
flabel metal1 12389 -9824 12442 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_422/VPWR
flabel metal1 12388 -10366 12439 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_422/VGND
rlabel comment 12367 -10348 12367 -10348 4 sky130_fd_sc_hd__tapvpwrvgnd_1_422/tapvpwrvgnd_1
rlabel metal1 12367 -10396 12459 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_422/VGND
rlabel metal1 12367 -9852 12459 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_422/VPWR
flabel metal1 16628 -10909 16662 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_34/VPWR
flabel metal1 16628 -10365 16662 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_34/VGND
flabel nwell 16628 -10909 16662 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_34/VPB
flabel pwell 16628 -10365 16662 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_34/VNB
rlabel comment 16691 -10348 16691 -10348 8 sky130_fd_sc_hd__decap_8_34/decap_8
rlabel metal1 15955 -10396 16691 -10300 5 sky130_fd_sc_hd__decap_8_34/VGND
rlabel metal1 15955 -10940 16691 -10844 5 sky130_fd_sc_hd__decap_8_34/VPWR
flabel metal1 15800 -10365 15834 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_27/VGND
flabel metal1 15800 -10909 15834 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_27/VPWR
flabel nwell 15800 -10909 15834 -10875 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_27/VPB
flabel pwell 15800 -10365 15834 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_27/VNB
rlabel comment 15863 -10348 15863 -10348 8 sky130_fd_sc_hd__decap_12_27/decap_12
rlabel metal1 14759 -10396 15863 -10300 5 sky130_fd_sc_hd__decap_12_27/VGND
rlabel metal1 14759 -10940 15863 -10844 5 sky130_fd_sc_hd__decap_12_27/VPWR
flabel metal1 15616 -10365 15650 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_29/VGND
flabel metal1 15616 -9821 15650 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_29/VPWR
flabel nwell 15616 -9821 15650 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_29/VPB
flabel pwell 15616 -10365 15650 -10331 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_29/VNB
rlabel comment 15587 -10348 15587 -10348 4 sky130_fd_sc_hd__decap_12_29/decap_12
rlabel metal1 15587 -10396 16691 -10300 1 sky130_fd_sc_hd__decap_12_29/VGND
rlabel metal1 15587 -9852 16691 -9756 1 sky130_fd_sc_hd__decap_12_29/VPWR
flabel metal1 14684 -10901 14737 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_398/VPWR
flabel metal1 14687 -10368 14738 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_398/VGND
rlabel comment 14759 -10348 14759 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_398/tapvpwrvgnd_1
rlabel metal1 14667 -10396 14759 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_398/VGND
rlabel metal1 14667 -10940 14759 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_398/VPWR
flabel metal1 15880 -10901 15933 -10872 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_399/VPWR
flabel metal1 15883 -10368 15934 -10330 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_399/VGND
rlabel comment 15955 -10348 15955 -10348 8 sky130_fd_sc_hd__tapvpwrvgnd_1_399/tapvpwrvgnd_1
rlabel metal1 15863 -10396 15955 -10300 5 sky130_fd_sc_hd__tapvpwrvgnd_1_399/VGND
rlabel metal1 15863 -10940 15955 -10844 5 sky130_fd_sc_hd__tapvpwrvgnd_1_399/VPWR
flabel metal1 15517 -9824 15570 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_423/VPWR
flabel metal1 15516 -10366 15567 -10328 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_423/VGND
rlabel comment 15495 -10348 15495 -10348 4 sky130_fd_sc_hd__tapvpwrvgnd_1_423/tapvpwrvgnd_1
rlabel metal1 15495 -10396 15587 -10300 1 sky130_fd_sc_hd__tapvpwrvgnd_1_423/VGND
rlabel metal1 15495 -9852 15587 -9756 1 sky130_fd_sc_hd__tapvpwrvgnd_1_423/VPWR
flabel metal1 -944 -9821 -910 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_38/VPWR
flabel metal1 -944 -9277 -910 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_38/VGND
flabel nwell -944 -9821 -910 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_38/VPB
flabel pwell -944 -9277 -910 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_38/VNB
rlabel comment -881 -9260 -881 -9260 8 sky130_fd_sc_hd__decap_8_38/decap_8
rlabel metal1 -1617 -9308 -881 -9212 5 sky130_fd_sc_hd__decap_8_38/VGND
rlabel metal1 -1617 -9852 -881 -9756 5 sky130_fd_sc_hd__decap_8_38/VPWR
flabel metal1 -2324 -9821 -2290 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_82/VPWR
flabel metal1 -2324 -9277 -2290 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_82/VGND
flabel nwell -2324 -9821 -2290 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_82/VPB
flabel pwell -2324 -9277 -2290 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_82/VNB
rlabel comment -2261 -9260 -2261 -9260 8 sky130_fd_sc_hd__decap_8_82/decap_8
rlabel metal1 -2997 -9308 -2261 -9212 5 sky130_fd_sc_hd__decap_8_82/VGND
rlabel metal1 -2997 -9852 -2261 -9756 5 sky130_fd_sc_hd__decap_8_82/VPWR
flabel metal1 -1690 -9278 -1637 -9246 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_21/VGND
flabel metal1 -1690 -9821 -1638 -9790 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_21/VPWR
flabel nwell -1679 -9813 -1645 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_21/VPB
flabel pwell -1680 -9272 -1648 -9250 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_21/VNB
rlabel comment -1617 -9260 -1617 -9260 8 sky130_fd_sc_hd__fill_2_21/fill_2
rlabel metal1 -1801 -9308 -1617 -9212 5 sky130_fd_sc_hd__fill_2_21/VGND
rlabel metal1 -1801 -9852 -1617 -9756 5 sky130_fd_sc_hd__fill_2_21/VPWR
flabel metal1 -1858 -9269 -1835 -9250 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_31/VGND
flabel metal1 -1855 -9812 -1835 -9795 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_31/VPWR
flabel nwell -1861 -9816 -1836 -9790 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_31/VPB
flabel pwell -1858 -9272 -1836 -9248 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_31/VNB
rlabel comment -1801 -9260 -1801 -9260 8 sky130_fd_sc_hd__fill_4_31/fill_4
rlabel metal1 -2169 -9308 -1801 -9212 5 sky130_fd_sc_hd__fill_4_31/VGND
rlabel metal1 -2169 -9852 -1801 -9756 5 sky130_fd_sc_hd__fill_4_31/VPWR
flabel metal1 -2244 -9813 -2191 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_547/VPWR
flabel metal1 -2241 -9280 -2190 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_547/VGND
rlabel comment -2169 -9260 -2169 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_547/tapvpwrvgnd_1
rlabel metal1 -2261 -9308 -2169 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_547/VGND
rlabel metal1 -2261 -9852 -2169 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_547/VPWR
flabel locali 1079 -9515 1113 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/A
flabel locali 433 -9719 467 -9685 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X
flabel locali 433 -9651 467 -9617 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X
flabel locali 433 -9583 467 -9549 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X
flabel locali 433 -9515 467 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X
flabel locali 433 -9447 467 -9413 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X
flabel locali 433 -9379 467 -9345 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X
flabel pwell 1079 -9277 1113 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/VNB
flabel nwell 1079 -9821 1113 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/VPB
flabel metal1 1079 -9277 1113 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/VGND
flabel metal1 1079 -9821 1113 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_168/VPWR
rlabel comment 1143 -9260 1143 -9260 8 sky130_fd_sc_hd__clkdlybuf4s50_1_168/clkdlybuf4s50_1
rlabel metal1 407 -9308 1143 -9212 5 sky130_fd_sc_hd__clkdlybuf4s50_1_168/VGND
rlabel metal1 407 -9852 1143 -9756 5 sky130_fd_sc_hd__clkdlybuf4s50_1_168/VPWR
flabel locali -209 -9515 -175 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A
flabel locali -855 -9719 -821 -9685 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X
flabel locali -855 -9651 -821 -9617 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X
flabel locali -855 -9583 -821 -9549 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X
flabel locali -855 -9515 -821 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X
flabel locali -855 -9447 -821 -9413 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X
flabel locali -855 -9379 -821 -9345 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/X
flabel pwell -209 -9277 -175 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/VNB
flabel nwell -209 -9821 -175 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/VPB
flabel metal1 -209 -9277 -175 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/VGND
flabel metal1 -209 -9821 -175 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_169/VPWR
rlabel comment -145 -9260 -145 -9260 8 sky130_fd_sc_hd__clkdlybuf4s50_1_169/clkdlybuf4s50_1
rlabel metal1 -881 -9308 -145 -9212 5 sky130_fd_sc_hd__clkdlybuf4s50_1_169/VGND
rlabel metal1 -881 -9852 -145 -9756 5 sky130_fd_sc_hd__clkdlybuf4s50_1_169/VPWR
flabel metal1 252 -9277 286 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_210/VGND
flabel metal1 252 -9821 286 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_210/VPWR
flabel nwell 252 -9821 286 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_210/VPB
flabel pwell 252 -9277 286 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_210/VNB
rlabel comment 315 -9260 315 -9260 8 sky130_fd_sc_hd__decap_4_210/decap_4
rlabel metal1 -53 -9308 315 -9212 5 sky130_fd_sc_hd__decap_4_210/VGND
rlabel metal1 -53 -9852 315 -9756 5 sky130_fd_sc_hd__decap_4_210/VPWR
flabel metal1 -128 -9813 -75 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_424/VPWR
flabel metal1 -125 -9280 -74 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_424/VGND
rlabel comment -53 -9260 -53 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_424/tapvpwrvgnd_1
rlabel metal1 -145 -9308 -53 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_424/VGND
rlabel metal1 -145 -9852 -53 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_424/VPWR
flabel metal1 332 -9813 385 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_425/VPWR
flabel metal1 335 -9280 386 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_425/VGND
rlabel comment 407 -9260 407 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_425/tapvpwrvgnd_1
rlabel metal1 315 -9308 407 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_425/VGND
rlabel metal1 315 -9852 407 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_425/VPWR
flabel metal1 2828 -9277 2862 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_211/VGND
flabel metal1 2828 -9821 2862 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_211/VPWR
flabel nwell 2828 -9821 2862 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_211/VPB
flabel pwell 2828 -9277 2862 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_211/VNB
rlabel comment 2891 -9260 2891 -9260 8 sky130_fd_sc_hd__decap_4_211/decap_4
rlabel metal1 2523 -9308 2891 -9212 5 sky130_fd_sc_hd__decap_4_211/VGND
rlabel metal1 2523 -9852 2891 -9756 5 sky130_fd_sc_hd__decap_4_211/VPWR
flabel metal1 1540 -9277 1574 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_212/VGND
flabel metal1 1540 -9821 1574 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_212/VPWR
flabel nwell 1540 -9821 1574 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_212/VPB
flabel pwell 1540 -9277 1574 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_212/VNB
rlabel comment 1603 -9260 1603 -9260 8 sky130_fd_sc_hd__decap_4_212/decap_4
rlabel metal1 1235 -9308 1603 -9212 5 sky130_fd_sc_hd__decap_4_212/VGND
rlabel metal1 1235 -9852 1603 -9756 5 sky130_fd_sc_hd__decap_4_212/VPWR
flabel metal1 2368 -9821 2402 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_133/VPWR
flabel metal1 2368 -9277 2402 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_133/VGND
flabel nwell 2368 -9821 2402 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_133/VPB
flabel pwell 2368 -9277 2402 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_133/VNB
rlabel comment 2431 -9260 2431 -9260 8 sky130_fd_sc_hd__decap_8_133/decap_8
rlabel metal1 1695 -9308 2431 -9212 5 sky130_fd_sc_hd__decap_8_133/VGND
rlabel metal1 1695 -9852 2431 -9756 5 sky130_fd_sc_hd__decap_8_133/VPWR
flabel metal1 2448 -9813 2501 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_426/VPWR
flabel metal1 2451 -9280 2502 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_426/VGND
rlabel comment 2523 -9260 2523 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_426/tapvpwrvgnd_1
rlabel metal1 2431 -9308 2523 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_426/VGND
rlabel metal1 2431 -9852 2523 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_426/VPWR
flabel metal1 1620 -9813 1673 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_427/VPWR
flabel metal1 1623 -9280 1674 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_427/VGND
rlabel comment 1695 -9260 1695 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_427/tapvpwrvgnd_1
rlabel metal1 1603 -9308 1695 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_427/VGND
rlabel metal1 1603 -9852 1695 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_427/VPWR
flabel metal1 1160 -9813 1213 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_428/VPWR
flabel metal1 1163 -9280 1214 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_428/VGND
rlabel comment 1235 -9260 1235 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_428/tapvpwrvgnd_1
rlabel metal1 1143 -9308 1235 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_428/VGND
rlabel metal1 1143 -9852 1235 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_428/VPWR
flabel locali 3655 -9515 3689 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A
flabel locali 3009 -9719 3043 -9685 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
flabel locali 3009 -9651 3043 -9617 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
flabel locali 3009 -9583 3043 -9549 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
flabel locali 3009 -9515 3043 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
flabel locali 3009 -9447 3043 -9413 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
flabel locali 3009 -9379 3043 -9345 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
flabel pwell 3655 -9277 3689 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/VNB
flabel nwell 3655 -9821 3689 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/VPB
flabel metal1 3655 -9277 3689 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/VGND
flabel metal1 3655 -9821 3689 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_172/VPWR
rlabel comment 3719 -9260 3719 -9260 8 sky130_fd_sc_hd__clkdlybuf4s50_1_172/clkdlybuf4s50_1
rlabel metal1 2983 -9308 3719 -9212 5 sky130_fd_sc_hd__clkdlybuf4s50_1_172/VGND
rlabel metal1 2983 -9852 3719 -9756 5 sky130_fd_sc_hd__clkdlybuf4s50_1_172/VPWR
flabel metal1 4116 -9277 4150 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_213/VGND
flabel metal1 4116 -9821 4150 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_213/VPWR
flabel nwell 4116 -9821 4150 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_213/VPB
flabel pwell 4116 -9277 4150 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_213/VNB
rlabel comment 4179 -9260 4179 -9260 8 sky130_fd_sc_hd__decap_4_213/decap_4
rlabel metal1 3811 -9308 4179 -9212 5 sky130_fd_sc_hd__decap_4_213/VGND
rlabel metal1 3811 -9852 4179 -9756 5 sky130_fd_sc_hd__decap_4_213/VPWR
flabel metal1 4944 -9821 4978 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_147/VPWR
flabel metal1 4944 -9277 4978 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_147/VGND
flabel nwell 4944 -9821 4978 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_147/VPB
flabel pwell 4944 -9277 4978 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_147/VNB
rlabel comment 5007 -9260 5007 -9260 8 sky130_fd_sc_hd__decap_8_147/decap_8
rlabel metal1 4271 -9308 5007 -9212 5 sky130_fd_sc_hd__decap_8_147/VGND
rlabel metal1 4271 -9852 5007 -9756 5 sky130_fd_sc_hd__decap_8_147/VPWR
flabel metal1 3736 -9813 3789 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_429/VPWR
flabel metal1 3739 -9280 3790 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_429/VGND
rlabel comment 3811 -9260 3811 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_429/tapvpwrvgnd_1
rlabel metal1 3719 -9308 3811 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_429/VGND
rlabel metal1 3719 -9852 3811 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_429/VPWR
flabel metal1 4196 -9813 4249 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_430/VPWR
flabel metal1 4199 -9280 4250 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_430/VGND
rlabel comment 4271 -9260 4271 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_430/tapvpwrvgnd_1
rlabel metal1 4179 -9308 4271 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_430/VGND
rlabel metal1 4179 -9852 4271 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_430/VPWR
flabel metal1 2908 -9813 2961 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_431/VPWR
flabel metal1 2911 -9280 2962 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_431/VGND
rlabel comment 2983 -9260 2983 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_431/tapvpwrvgnd_1
rlabel metal1 2891 -9308 2983 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_431/VGND
rlabel metal1 2891 -9852 2983 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_431/VPWR
flabel locali 6231 -9515 6265 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/A
flabel locali 5585 -9719 5619 -9685 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X
flabel locali 5585 -9651 5619 -9617 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X
flabel locali 5585 -9583 5619 -9549 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X
flabel locali 5585 -9515 5619 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X
flabel locali 5585 -9447 5619 -9413 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X
flabel locali 5585 -9379 5619 -9345 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X
flabel pwell 6231 -9277 6265 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/VNB
flabel nwell 6231 -9821 6265 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/VPB
flabel metal1 6231 -9277 6265 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/VGND
flabel metal1 6231 -9821 6265 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_173/VPWR
rlabel comment 6295 -9260 6295 -9260 8 sky130_fd_sc_hd__clkdlybuf4s50_1_173/clkdlybuf4s50_1
rlabel metal1 5559 -9308 6295 -9212 5 sky130_fd_sc_hd__clkdlybuf4s50_1_173/VGND
rlabel metal1 5559 -9852 6295 -9756 5 sky130_fd_sc_hd__clkdlybuf4s50_1_173/VPWR
flabel metal1 6692 -9277 6726 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_214/VGND
flabel metal1 6692 -9821 6726 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_214/VPWR
flabel nwell 6692 -9821 6726 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_214/VPB
flabel pwell 6692 -9277 6726 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_214/VNB
rlabel comment 6755 -9260 6755 -9260 8 sky130_fd_sc_hd__decap_4_214/decap_4
rlabel metal1 6387 -9308 6755 -9212 5 sky130_fd_sc_hd__decap_4_214/VGND
rlabel metal1 6387 -9852 6755 -9756 5 sky130_fd_sc_hd__decap_4_214/VPWR
flabel metal1 5404 -9277 5438 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_215/VGND
flabel metal1 5404 -9821 5438 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_215/VPWR
flabel nwell 5404 -9821 5438 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_215/VPB
flabel pwell 5404 -9277 5438 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_215/VNB
rlabel comment 5467 -9260 5467 -9260 8 sky130_fd_sc_hd__decap_4_215/decap_4
rlabel metal1 5099 -9308 5467 -9212 5 sky130_fd_sc_hd__decap_4_215/VGND
rlabel metal1 5099 -9852 5467 -9756 5 sky130_fd_sc_hd__decap_4_215/VPWR
flabel metal1 6312 -9813 6365 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_432/VPWR
flabel metal1 6315 -9280 6366 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_432/VGND
rlabel comment 6387 -9260 6387 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_432/tapvpwrvgnd_1
rlabel metal1 6295 -9308 6387 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_432/VGND
rlabel metal1 6295 -9852 6387 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_432/VPWR
flabel metal1 5484 -9813 5537 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_433/VPWR
flabel metal1 5487 -9280 5538 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_433/VGND
rlabel comment 5559 -9260 5559 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_433/tapvpwrvgnd_1
rlabel metal1 5467 -9308 5559 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_433/VGND
rlabel metal1 5467 -9852 5559 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_433/VPWR
flabel metal1 5024 -9813 5077 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_434/VPWR
flabel metal1 5027 -9280 5078 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_434/VGND
rlabel comment 5099 -9260 5099 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_434/tapvpwrvgnd_1
rlabel metal1 5007 -9308 5099 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_434/VGND
rlabel metal1 5007 -9852 5099 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_434/VPWR
flabel locali 8807 -9515 8841 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/A
flabel locali 8161 -9719 8195 -9685 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X
flabel locali 8161 -9651 8195 -9617 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X
flabel locali 8161 -9583 8195 -9549 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X
flabel locali 8161 -9515 8195 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X
flabel locali 8161 -9447 8195 -9413 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X
flabel locali 8161 -9379 8195 -9345 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X
flabel pwell 8807 -9277 8841 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/VNB
flabel nwell 8807 -9821 8841 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/VPB
flabel metal1 8807 -9277 8841 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/VGND
flabel metal1 8807 -9821 8841 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_174/VPWR
rlabel comment 8871 -9260 8871 -9260 8 sky130_fd_sc_hd__clkdlybuf4s50_1_174/clkdlybuf4s50_1
rlabel metal1 8135 -9308 8871 -9212 5 sky130_fd_sc_hd__clkdlybuf4s50_1_174/VGND
rlabel metal1 8135 -9852 8871 -9756 5 sky130_fd_sc_hd__clkdlybuf4s50_1_174/VPWR
flabel metal1 7980 -9277 8014 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_216/VGND
flabel metal1 7980 -9821 8014 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_216/VPWR
flabel nwell 7980 -9821 8014 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_216/VPB
flabel pwell 7980 -9277 8014 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_216/VNB
rlabel comment 8043 -9260 8043 -9260 8 sky130_fd_sc_hd__decap_4_216/decap_4
rlabel metal1 7675 -9308 8043 -9212 5 sky130_fd_sc_hd__decap_4_216/VGND
rlabel metal1 7675 -9852 8043 -9756 5 sky130_fd_sc_hd__decap_4_216/VPWR
flabel metal1 7520 -9821 7554 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_157/VPWR
flabel metal1 7520 -9277 7554 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_157/VGND
flabel nwell 7520 -9821 7554 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_157/VPB
flabel pwell 7520 -9277 7554 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_157/VNB
rlabel comment 7583 -9260 7583 -9260 8 sky130_fd_sc_hd__decap_8_157/decap_8
rlabel metal1 6847 -9308 7583 -9212 5 sky130_fd_sc_hd__decap_8_157/VGND
rlabel metal1 6847 -9852 7583 -9756 5 sky130_fd_sc_hd__decap_8_157/VPWR
flabel metal1 7600 -9813 7653 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_435/VPWR
flabel metal1 7603 -9280 7654 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_435/VGND
rlabel comment 7675 -9260 7675 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_435/tapvpwrvgnd_1
rlabel metal1 7583 -9308 7675 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_435/VGND
rlabel metal1 7583 -9852 7675 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_435/VPWR
flabel metal1 8060 -9813 8113 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_436/VPWR
flabel metal1 8063 -9280 8114 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_436/VGND
rlabel comment 8135 -9260 8135 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_436/tapvpwrvgnd_1
rlabel metal1 8043 -9308 8135 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_436/VGND
rlabel metal1 8043 -9852 8135 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_436/VPWR
flabel metal1 6772 -9813 6825 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_437/VPWR
flabel metal1 6775 -9280 6826 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_437/VGND
rlabel comment 6847 -9260 6847 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_437/tapvpwrvgnd_1
rlabel metal1 6755 -9308 6847 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_437/VGND
rlabel metal1 6755 -9852 6847 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_437/VPWR
flabel metal1 9268 -9277 9302 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_217/VGND
flabel metal1 9268 -9821 9302 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_217/VPWR
flabel nwell 9268 -9821 9302 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_217/VPB
flabel pwell 9268 -9277 9302 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_217/VNB
rlabel comment 9331 -9260 9331 -9260 8 sky130_fd_sc_hd__decap_4_217/decap_4
rlabel metal1 8963 -9308 9331 -9212 5 sky130_fd_sc_hd__decap_4_217/VGND
rlabel metal1 8963 -9852 9331 -9756 5 sky130_fd_sc_hd__decap_4_217/VPWR
flabel metal1 10648 -9277 10682 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_219/VGND
flabel metal1 10648 -9821 10682 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_219/VPWR
flabel nwell 10648 -9821 10682 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_219/VPB
flabel pwell 10648 -9277 10682 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_219/VNB
rlabel comment 10711 -9260 10711 -9260 8 sky130_fd_sc_hd__decap_4_219/decap_4
rlabel metal1 10343 -9308 10711 -9212 5 sky130_fd_sc_hd__decap_4_219/VGND
rlabel metal1 10343 -9852 10711 -9756 5 sky130_fd_sc_hd__decap_4_219/VPWR
flabel metal1 10096 -9821 10130 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_168/VPWR
flabel metal1 10096 -9277 10130 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_168/VGND
flabel nwell 10096 -9821 10130 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_168/VPB
flabel pwell 10096 -9277 10130 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_168/VNB
rlabel comment 10159 -9260 10159 -9260 8 sky130_fd_sc_hd__decap_8_168/decap_8
rlabel metal1 9423 -9308 10159 -9212 5 sky130_fd_sc_hd__decap_8_168/VGND
rlabel metal1 9423 -9852 10159 -9756 5 sky130_fd_sc_hd__decap_8_168/VPWR
flabel metal1 10285 -9817 10321 -9787 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_60/VPWR
flabel metal1 10285 -9276 10321 -9247 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_60/VGND
flabel nwell 10292 -9811 10312 -9794 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_60/VPB
flabel pwell 10291 -9271 10315 -9249 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_60/VNB
rlabel comment 10343 -9260 10343 -9260 8 sky130_fd_sc_hd__fill_1_60/fill_1
rlabel metal1 10251 -9308 10343 -9212 5 sky130_fd_sc_hd__fill_1_60/VGND
rlabel metal1 10251 -9852 10343 -9756 5 sky130_fd_sc_hd__fill_1_60/VPWR
flabel metal1 10176 -9813 10229 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_438/VPWR
flabel metal1 10179 -9280 10230 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_438/VGND
rlabel comment 10251 -9260 10251 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_438/tapvpwrvgnd_1
rlabel metal1 10159 -9308 10251 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_438/VGND
rlabel metal1 10159 -9852 10251 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_438/VPWR
flabel metal1 9348 -9813 9401 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_439/VPWR
flabel metal1 9351 -9280 9402 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_439/VGND
rlabel comment 9423 -9260 9423 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_439/tapvpwrvgnd_1
rlabel metal1 9331 -9308 9423 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_439/VGND
rlabel metal1 9331 -9852 9423 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_439/VPWR
flabel metal1 8888 -9813 8941 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_440/VPWR
flabel metal1 8891 -9280 8942 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_440/VGND
rlabel comment 8963 -9260 8963 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_440/tapvpwrvgnd_1
rlabel metal1 8871 -9308 8963 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_440/VGND
rlabel metal1 8871 -9852 8963 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_440/VPWR
flabel locali 11383 -9515 11417 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/A
flabel locali 10737 -9719 10771 -9685 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X
flabel locali 10737 -9651 10771 -9617 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X
flabel locali 10737 -9583 10771 -9549 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X
flabel locali 10737 -9515 10771 -9481 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X
flabel locali 10737 -9447 10771 -9413 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X
flabel locali 10737 -9379 10771 -9345 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X
flabel pwell 11383 -9277 11417 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/VNB
flabel nwell 11383 -9821 11417 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/VPB
flabel metal1 11383 -9277 11417 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/VGND
flabel metal1 11383 -9821 11417 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_177/VPWR
rlabel comment 11447 -9260 11447 -9260 8 sky130_fd_sc_hd__clkdlybuf4s50_1_177/clkdlybuf4s50_1
rlabel metal1 10711 -9308 11447 -9212 5 sky130_fd_sc_hd__clkdlybuf4s50_1_177/VGND
rlabel metal1 10711 -9852 11447 -9756 5 sky130_fd_sc_hd__clkdlybuf4s50_1_177/VPWR
flabel metal1 11936 -9277 11970 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_218/VGND
flabel metal1 11936 -9821 11970 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_218/VPWR
flabel nwell 11936 -9821 11970 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_218/VPB
flabel pwell 11936 -9277 11970 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_218/VNB
rlabel comment 11999 -9260 11999 -9260 8 sky130_fd_sc_hd__decap_4_218/decap_4
rlabel metal1 11631 -9308 11999 -9212 5 sky130_fd_sc_hd__decap_4_218/VGND
rlabel metal1 11631 -9852 11999 -9756 5 sky130_fd_sc_hd__decap_4_218/VPWR
flabel metal1 11573 -9817 11609 -9787 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_61/VPWR
flabel metal1 11573 -9276 11609 -9247 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_61/VGND
flabel nwell 11580 -9811 11600 -9794 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_61/VPB
flabel pwell 11579 -9271 11603 -9249 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_61/VNB
rlabel comment 11631 -9260 11631 -9260 8 sky130_fd_sc_hd__fill_1_61/fill_1
rlabel metal1 11539 -9308 11631 -9212 5 sky130_fd_sc_hd__fill_1_61/VGND
rlabel metal1 11539 -9852 11631 -9756 5 sky130_fd_sc_hd__fill_1_61/VPWR
flabel metal1 10653 -9817 10689 -9787 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_62/VPWR
flabel metal1 10653 -9276 10689 -9247 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_62/VGND
flabel nwell 10660 -9811 10680 -9794 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_62/VPB
flabel pwell 10659 -9271 10683 -9249 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_62/VNB
rlabel comment 10711 -9260 10711 -9260 8 sky130_fd_sc_hd__fill_1_62/fill_1
rlabel metal1 10619 -9308 10711 -9212 5 sky130_fd_sc_hd__fill_1_62/VGND
rlabel metal1 10619 -9852 10711 -9756 5 sky130_fd_sc_hd__fill_1_62/VPWR
flabel metal1 12668 -9270 12700 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_29/VGND
flabel metal1 12668 -9815 12706 -9783 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_29/VPWR
flabel nwell 12658 -9813 12715 -9782 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_29/VPB
flabel pwell 12665 -9270 12709 -9236 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_29/VNB
rlabel comment 12735 -9260 12735 -9260 8 sky130_fd_sc_hd__fill_8_29/fill_8
rlabel metal1 11999 -9308 12735 -9212 5 sky130_fd_sc_hd__fill_8_29/VGND
rlabel metal1 11999 -9852 12735 -9756 5 sky130_fd_sc_hd__fill_8_29/VPWR
flabel metal1 11464 -9813 11517 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_441/VPWR
flabel metal1 11467 -9280 11518 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_441/VGND
rlabel comment 11539 -9260 11539 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_441/tapvpwrvgnd_1
rlabel metal1 11447 -9308 11539 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_441/VGND
rlabel metal1 11447 -9852 11539 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_441/VPWR
flabel locali 15248 -9583 15282 -9549 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/X
flabel locali 15340 -9583 15374 -9549 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/X
flabel locali 15340 -9515 15374 -9481 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/X
flabel locali 15248 -9515 15282 -9481 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/X
flabel locali 15248 -9447 15282 -9413 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/X
flabel locali 15340 -9447 15374 -9413 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/X
flabel locali 13684 -9447 13718 -9413 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/A
flabel locali 13684 -9515 13718 -9481 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/A
flabel pwell 13684 -9277 13718 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/VNB
flabel pwell 13701 -9260 13701 -9260 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/VNB
flabel nwell 13684 -9821 13718 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/VPB
flabel nwell 13701 -9804 13701 -9804 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/VPB
flabel metal1 13684 -9277 13718 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/VGND
flabel metal1 13684 -9821 13718 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_13/VPWR
rlabel comment 13655 -9260 13655 -9260 2 sky130_fd_sc_hd__clkbuf_16_13/clkbuf_16
rlabel metal1 13655 -9308 15495 -9212 5 sky130_fd_sc_hd__clkbuf_16_13/VGND
rlabel metal1 13655 -9852 15495 -9756 5 sky130_fd_sc_hd__clkbuf_16_13/VPWR
flabel metal1 13505 -9817 13541 -9787 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_63/VPWR
flabel metal1 13505 -9276 13541 -9247 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_63/VGND
flabel nwell 13512 -9811 13532 -9794 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_63/VPB
flabel pwell 13511 -9271 13535 -9249 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_63/VNB
rlabel comment 13563 -9260 13563 -9260 8 sky130_fd_sc_hd__fill_1_63/fill_1
rlabel metal1 13471 -9308 13563 -9212 5 sky130_fd_sc_hd__fill_1_63/VGND
rlabel metal1 13471 -9852 13563 -9756 5 sky130_fd_sc_hd__fill_1_63/VPWR
flabel metal1 13404 -9270 13436 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_30/VGND
flabel metal1 13404 -9815 13442 -9783 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_30/VPWR
flabel nwell 13394 -9813 13451 -9782 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_30/VPB
flabel pwell 13401 -9270 13445 -9236 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_30/VNB
rlabel comment 13471 -9260 13471 -9260 8 sky130_fd_sc_hd__fill_8_30/fill_8
rlabel metal1 12735 -9308 13471 -9212 5 sky130_fd_sc_hd__fill_8_30/VGND
rlabel metal1 12735 -9852 13471 -9756 5 sky130_fd_sc_hd__fill_8_30/VPWR
flabel metal1 13580 -9813 13633 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_442/VPWR
flabel metal1 13583 -9280 13634 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_442/VGND
rlabel comment 13655 -9260 13655 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_442/tapvpwrvgnd_1
rlabel metal1 13563 -9308 13655 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_442/VGND
rlabel metal1 13563 -9852 13655 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_442/VPWR
flabel metal1 16628 -9277 16662 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_30/VGND
flabel metal1 16628 -9821 16662 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_30/VPWR
flabel nwell 16628 -9821 16662 -9787 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_30/VPB
flabel pwell 16628 -9277 16662 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_30/VNB
rlabel comment 16691 -9260 16691 -9260 8 sky130_fd_sc_hd__decap_12_30/decap_12
rlabel metal1 15587 -9308 16691 -9212 5 sky130_fd_sc_hd__decap_12_30/VGND
rlabel metal1 15587 -9852 16691 -9756 5 sky130_fd_sc_hd__decap_12_30/VPWR
flabel metal1 15512 -9813 15565 -9784 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_443/VPWR
flabel metal1 15515 -9280 15566 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_443/VGND
rlabel comment 15587 -9260 15587 -9260 8 sky130_fd_sc_hd__tapvpwrvgnd_1_443/tapvpwrvgnd_1
rlabel metal1 15495 -9308 15587 -9212 5 sky130_fd_sc_hd__tapvpwrvgnd_1_443/VGND
rlabel metal1 15495 -9852 15587 -9756 5 sky130_fd_sc_hd__tapvpwrvgnd_1_443/VPWR
flabel metal1 -1588 -8733 -1554 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_39/VPWR
flabel metal1 -1588 -9277 -1554 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_39/VGND
flabel nwell -1588 -8733 -1554 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_39/VPB
flabel pwell -1588 -9277 -1554 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_39/VNB
rlabel comment -1617 -9260 -1617 -9260 4 sky130_fd_sc_hd__decap_8_39/decap_8
rlabel metal1 -1617 -9308 -881 -9212 1 sky130_fd_sc_hd__decap_8_39/VGND
rlabel metal1 -1617 -8764 -881 -8668 1 sky130_fd_sc_hd__decap_8_39/VPWR
flabel metal1 -2968 -8733 -2934 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_81/VPWR
flabel metal1 -2968 -9277 -2934 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_81/VGND
flabel nwell -2968 -8733 -2934 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_81/VPB
flabel pwell -2968 -9277 -2934 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_81/VNB
rlabel comment -2997 -9260 -2997 -9260 4 sky130_fd_sc_hd__decap_8_81/decap_8
rlabel metal1 -2997 -9308 -2261 -9212 1 sky130_fd_sc_hd__decap_8_81/VGND
rlabel metal1 -2997 -8764 -2261 -8668 1 sky130_fd_sc_hd__decap_8_81/VPWR
flabel metal1 -1781 -9274 -1728 -9242 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_20/VGND
flabel metal1 -1780 -8730 -1728 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_20/VPWR
flabel nwell -1773 -8725 -1739 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_20/VPB
flabel pwell -1770 -9270 -1738 -9248 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_20/VNB
rlabel comment -1801 -9260 -1801 -9260 4 sky130_fd_sc_hd__fill_2_20/fill_2
rlabel metal1 -1801 -9308 -1617 -9212 1 sky130_fd_sc_hd__fill_2_20/VGND
rlabel metal1 -1801 -8764 -1617 -8668 1 sky130_fd_sc_hd__fill_2_20/VPWR
flabel metal1 -2135 -9270 -2112 -9251 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_30/VGND
flabel metal1 -2135 -8725 -2115 -8708 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_30/VPWR
flabel nwell -2134 -8730 -2109 -8704 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_30/VPB
flabel pwell -2134 -9272 -2112 -9248 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_30/VNB
rlabel comment -2169 -9260 -2169 -9260 4 sky130_fd_sc_hd__fill_4_30/fill_4
rlabel metal1 -2169 -9308 -1801 -9212 1 sky130_fd_sc_hd__fill_4_30/VGND
rlabel metal1 -2169 -8764 -1801 -8668 1 sky130_fd_sc_hd__fill_4_30/VPWR
flabel metal1 -2239 -8736 -2186 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_546/VPWR
flabel metal1 -2240 -9278 -2189 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_546/VGND
rlabel comment -2261 -9260 -2261 -9260 4 sky130_fd_sc_hd__tapvpwrvgnd_1_546/tapvpwrvgnd_1
rlabel metal1 -2261 -9308 -2169 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_546/VGND
rlabel metal1 -2261 -8764 -2169 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_546/VPWR
flabel locali 437 -9039 471 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/A
flabel locali 1083 -8835 1117 -8801 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/X
flabel locali 1083 -8903 1117 -8869 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/X
flabel locali 1083 -8971 1117 -8937 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/X
flabel locali 1083 -9039 1117 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/X
flabel locali 1083 -9107 1117 -9073 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/X
flabel locali 1083 -9175 1117 -9141 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/X
flabel pwell 437 -9277 471 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/VNB
flabel nwell 437 -8733 471 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/VPB
flabel metal1 437 -9277 471 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/VGND
flabel metal1 437 -8733 471 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_178/VPWR
rlabel comment 407 -9260 407 -9260 4 sky130_fd_sc_hd__clkdlybuf4s50_1_178/clkdlybuf4s50_1
rlabel metal1 407 -9308 1143 -9212 1 sky130_fd_sc_hd__clkdlybuf4s50_1_178/VGND
rlabel metal1 407 -8764 1143 -8668 1 sky130_fd_sc_hd__clkdlybuf4s50_1_178/VPWR
flabel metal1 252 -9277 286 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_220/VGND
flabel metal1 252 -8733 286 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_220/VPWR
flabel nwell 252 -8733 286 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_220/VPB
flabel pwell 252 -9277 286 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_220/VNB
rlabel comment 315 -9260 315 -9260 6 sky130_fd_sc_hd__decap_4_220/decap_4
rlabel metal1 -53 -9308 315 -9212 1 sky130_fd_sc_hd__decap_4_220/VGND
rlabel metal1 -53 -8764 315 -8668 1 sky130_fd_sc_hd__decap_4_220/VPWR
flabel metal1 -852 -8733 -818 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_40/VPWR
flabel metal1 -852 -9277 -818 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_40/VGND
flabel nwell -852 -8733 -818 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_40/VPB
flabel pwell -852 -9277 -818 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_40/VNB
rlabel comment -881 -9260 -881 -9260 4 sky130_fd_sc_hd__decap_8_40/decap_8
rlabel metal1 -881 -9308 -145 -9212 1 sky130_fd_sc_hd__decap_8_40/VGND
rlabel metal1 -881 -8764 -145 -8668 1 sky130_fd_sc_hd__decap_8_40/VPWR
flabel metal1 332 -8736 385 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_444/VPWR
flabel metal1 335 -9278 386 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_444/VGND
rlabel comment 407 -9260 407 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_444/tapvpwrvgnd_1
rlabel metal1 315 -9308 407 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_444/VGND
rlabel metal1 315 -8764 407 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_444/VPWR
flabel metal1 -128 -8736 -75 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_445/VPWR
flabel metal1 -125 -9278 -74 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_445/VGND
rlabel comment -53 -9260 -53 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_445/tapvpwrvgnd_1
rlabel metal1 -145 -9308 -53 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_445/VGND
rlabel metal1 -145 -8764 -53 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_445/VPWR
flabel metal1 1540 -9277 1574 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_221/VGND
flabel metal1 1540 -8733 1574 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_221/VPWR
flabel nwell 1540 -8733 1574 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_221/VPB
flabel pwell 1540 -9277 1574 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_221/VNB
rlabel comment 1603 -9260 1603 -9260 6 sky130_fd_sc_hd__decap_4_221/decap_4
rlabel metal1 1235 -9308 1603 -9212 1 sky130_fd_sc_hd__decap_4_221/VGND
rlabel metal1 1235 -8764 1603 -8668 1 sky130_fd_sc_hd__decap_4_221/VPWR
flabel metal1 2828 -9277 2862 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_222/VGND
flabel metal1 2828 -8733 2862 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_222/VPWR
flabel nwell 2828 -8733 2862 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_222/VPB
flabel pwell 2828 -9277 2862 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_222/VNB
rlabel comment 2891 -9260 2891 -9260 6 sky130_fd_sc_hd__decap_4_222/decap_4
rlabel metal1 2523 -9308 2891 -9212 1 sky130_fd_sc_hd__decap_4_222/VGND
rlabel metal1 2523 -8764 2891 -8668 1 sky130_fd_sc_hd__decap_4_222/VPWR
flabel metal1 1724 -8733 1758 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_132/VPWR
flabel metal1 1724 -9277 1758 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_132/VGND
flabel nwell 1724 -8733 1758 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_132/VPB
flabel pwell 1724 -9277 1758 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_132/VNB
rlabel comment 1695 -9260 1695 -9260 4 sky130_fd_sc_hd__decap_8_132/decap_8
rlabel metal1 1695 -9308 2431 -9212 1 sky130_fd_sc_hd__decap_8_132/VGND
rlabel metal1 1695 -8764 2431 -8668 1 sky130_fd_sc_hd__decap_8_132/VPWR
flabel metal1 1160 -8736 1213 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_446/VPWR
flabel metal1 1163 -9278 1214 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_446/VGND
rlabel comment 1235 -9260 1235 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_446/tapvpwrvgnd_1
rlabel metal1 1143 -9308 1235 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_446/VGND
rlabel metal1 1143 -8764 1235 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_446/VPWR
flabel metal1 1620 -8736 1673 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_447/VPWR
flabel metal1 1623 -9278 1674 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_447/VGND
rlabel comment 1695 -9260 1695 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_447/tapvpwrvgnd_1
rlabel metal1 1603 -9308 1695 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_447/VGND
rlabel metal1 1603 -8764 1695 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_447/VPWR
flabel metal1 2448 -8736 2501 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_448/VPWR
flabel metal1 2451 -9278 2502 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_448/VGND
rlabel comment 2523 -9260 2523 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_448/tapvpwrvgnd_1
rlabel metal1 2431 -9308 2523 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_448/VGND
rlabel metal1 2431 -8764 2523 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_448/VPWR
flabel locali 3013 -9039 3047 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A
flabel locali 3659 -8835 3693 -8801 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/X
flabel locali 3659 -8903 3693 -8869 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/X
flabel locali 3659 -8971 3693 -8937 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/X
flabel locali 3659 -9039 3693 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/X
flabel locali 3659 -9107 3693 -9073 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/X
flabel locali 3659 -9175 3693 -9141 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/X
flabel pwell 3013 -9277 3047 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/VNB
flabel nwell 3013 -8733 3047 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/VPB
flabel metal1 3013 -9277 3047 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/VGND
flabel metal1 3013 -8733 3047 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_180/VPWR
rlabel comment 2983 -9260 2983 -9260 4 sky130_fd_sc_hd__clkdlybuf4s50_1_180/clkdlybuf4s50_1
rlabel metal1 2983 -9308 3719 -9212 1 sky130_fd_sc_hd__clkdlybuf4s50_1_180/VGND
rlabel metal1 2983 -8764 3719 -8668 1 sky130_fd_sc_hd__clkdlybuf4s50_1_180/VPWR
flabel metal1 4116 -9277 4150 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_223/VGND
flabel metal1 4116 -8733 4150 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_223/VPWR
flabel nwell 4116 -8733 4150 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_223/VPB
flabel pwell 4116 -9277 4150 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_223/VNB
rlabel comment 4179 -9260 4179 -9260 6 sky130_fd_sc_hd__decap_4_223/decap_4
rlabel metal1 3811 -9308 4179 -9212 1 sky130_fd_sc_hd__decap_4_223/VGND
rlabel metal1 3811 -8764 4179 -8668 1 sky130_fd_sc_hd__decap_4_223/VPWR
flabel metal1 4300 -8733 4334 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_150/VPWR
flabel metal1 4300 -9277 4334 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_150/VGND
flabel nwell 4300 -8733 4334 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_150/VPB
flabel pwell 4300 -9277 4334 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_150/VNB
rlabel comment 4271 -9260 4271 -9260 4 sky130_fd_sc_hd__decap_8_150/decap_8
rlabel metal1 4271 -9308 5007 -9212 1 sky130_fd_sc_hd__decap_8_150/VGND
rlabel metal1 4271 -8764 5007 -8668 1 sky130_fd_sc_hd__decap_8_150/VPWR
flabel metal1 2908 -8736 2961 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_449/VPWR
flabel metal1 2911 -9278 2962 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_449/VGND
rlabel comment 2983 -9260 2983 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_449/tapvpwrvgnd_1
rlabel metal1 2891 -9308 2983 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_449/VGND
rlabel metal1 2891 -8764 2983 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_449/VPWR
flabel metal1 4196 -8736 4249 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_450/VPWR
flabel metal1 4199 -9278 4250 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_450/VGND
rlabel comment 4271 -9260 4271 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_450/tapvpwrvgnd_1
rlabel metal1 4179 -9308 4271 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_450/VGND
rlabel metal1 4179 -8764 4271 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_450/VPWR
flabel metal1 3736 -8736 3789 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_451/VPWR
flabel metal1 3739 -9278 3790 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_451/VGND
rlabel comment 3811 -9260 3811 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_451/tapvpwrvgnd_1
rlabel metal1 3719 -9308 3811 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_451/VGND
rlabel metal1 3719 -8764 3811 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_451/VPWR
flabel locali 5589 -9039 5623 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A
flabel locali 6235 -8835 6269 -8801 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/X
flabel locali 6235 -8903 6269 -8869 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/X
flabel locali 6235 -8971 6269 -8937 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/X
flabel locali 6235 -9039 6269 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/X
flabel locali 6235 -9107 6269 -9073 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/X
flabel locali 6235 -9175 6269 -9141 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/X
flabel pwell 5589 -9277 5623 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/VNB
flabel nwell 5589 -8733 5623 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/VPB
flabel metal1 5589 -9277 5623 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/VGND
flabel metal1 5589 -8733 5623 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_182/VPWR
rlabel comment 5559 -9260 5559 -9260 4 sky130_fd_sc_hd__clkdlybuf4s50_1_182/clkdlybuf4s50_1
rlabel metal1 5559 -9308 6295 -9212 1 sky130_fd_sc_hd__clkdlybuf4s50_1_182/VGND
rlabel metal1 5559 -8764 6295 -8668 1 sky130_fd_sc_hd__clkdlybuf4s50_1_182/VPWR
flabel metal1 5404 -9277 5438 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_224/VGND
flabel metal1 5404 -8733 5438 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_224/VPWR
flabel nwell 5404 -8733 5438 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_224/VPB
flabel pwell 5404 -9277 5438 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_224/VNB
rlabel comment 5467 -9260 5467 -9260 6 sky130_fd_sc_hd__decap_4_224/decap_4
rlabel metal1 5099 -9308 5467 -9212 1 sky130_fd_sc_hd__decap_4_224/VGND
rlabel metal1 5099 -8764 5467 -8668 1 sky130_fd_sc_hd__decap_4_224/VPWR
flabel metal1 6692 -9277 6726 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_225/VGND
flabel metal1 6692 -8733 6726 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_225/VPWR
flabel nwell 6692 -8733 6726 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_225/VPB
flabel pwell 6692 -9277 6726 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_225/VNB
rlabel comment 6755 -9260 6755 -9260 6 sky130_fd_sc_hd__decap_4_225/decap_4
rlabel metal1 6387 -9308 6755 -9212 1 sky130_fd_sc_hd__decap_4_225/VGND
rlabel metal1 6387 -8764 6755 -8668 1 sky130_fd_sc_hd__decap_4_225/VPWR
flabel metal1 5024 -8736 5077 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_452/VPWR
flabel metal1 5027 -9278 5078 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_452/VGND
rlabel comment 5099 -9260 5099 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_452/tapvpwrvgnd_1
rlabel metal1 5007 -9308 5099 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_452/VGND
rlabel metal1 5007 -8764 5099 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_452/VPWR
flabel metal1 5484 -8736 5537 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_453/VPWR
flabel metal1 5487 -9278 5538 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_453/VGND
rlabel comment 5559 -9260 5559 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_453/tapvpwrvgnd_1
rlabel metal1 5467 -9308 5559 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_453/VGND
rlabel metal1 5467 -8764 5559 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_453/VPWR
flabel metal1 6312 -8736 6365 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_454/VPWR
flabel metal1 6315 -9278 6366 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_454/VGND
rlabel comment 6387 -9260 6387 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_454/tapvpwrvgnd_1
rlabel metal1 6295 -9308 6387 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_454/VGND
rlabel metal1 6295 -8764 6387 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_454/VPWR
flabel locali 8165 -9039 8199 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A
flabel locali 8811 -8835 8845 -8801 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/X
flabel locali 8811 -8903 8845 -8869 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/X
flabel locali 8811 -8971 8845 -8937 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/X
flabel locali 8811 -9039 8845 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/X
flabel locali 8811 -9107 8845 -9073 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/X
flabel locali 8811 -9175 8845 -9141 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/X
flabel pwell 8165 -9277 8199 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/VNB
flabel nwell 8165 -8733 8199 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/VPB
flabel metal1 8165 -9277 8199 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/VGND
flabel metal1 8165 -8733 8199 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_184/VPWR
rlabel comment 8135 -9260 8135 -9260 4 sky130_fd_sc_hd__clkdlybuf4s50_1_184/clkdlybuf4s50_1
rlabel metal1 8135 -9308 8871 -9212 1 sky130_fd_sc_hd__clkdlybuf4s50_1_184/VGND
rlabel metal1 8135 -8764 8871 -8668 1 sky130_fd_sc_hd__clkdlybuf4s50_1_184/VPWR
flabel metal1 7980 -9277 8014 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_226/VGND
flabel metal1 7980 -8733 8014 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_226/VPWR
flabel nwell 7980 -8733 8014 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_226/VPB
flabel pwell 7980 -9277 8014 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_226/VNB
rlabel comment 8043 -9260 8043 -9260 6 sky130_fd_sc_hd__decap_4_226/decap_4
rlabel metal1 7675 -9308 8043 -9212 1 sky130_fd_sc_hd__decap_4_226/VGND
rlabel metal1 7675 -8764 8043 -8668 1 sky130_fd_sc_hd__decap_4_226/VPWR
flabel metal1 6876 -8733 6910 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_159/VPWR
flabel metal1 6876 -9277 6910 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_159/VGND
flabel nwell 6876 -8733 6910 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_159/VPB
flabel pwell 6876 -9277 6910 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_159/VNB
rlabel comment 6847 -9260 6847 -9260 4 sky130_fd_sc_hd__decap_8_159/decap_8
rlabel metal1 6847 -9308 7583 -9212 1 sky130_fd_sc_hd__decap_8_159/VGND
rlabel metal1 6847 -8764 7583 -8668 1 sky130_fd_sc_hd__decap_8_159/VPWR
flabel metal1 6772 -8736 6825 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_455/VPWR
flabel metal1 6775 -9278 6826 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_455/VGND
rlabel comment 6847 -9260 6847 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_455/tapvpwrvgnd_1
rlabel metal1 6755 -9308 6847 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_455/VGND
rlabel metal1 6755 -8764 6847 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_455/VPWR
flabel metal1 8060 -8736 8113 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_456/VPWR
flabel metal1 8063 -9278 8114 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_456/VGND
rlabel comment 8135 -9260 8135 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_456/tapvpwrvgnd_1
rlabel metal1 8043 -9308 8135 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_456/VGND
rlabel metal1 8043 -8764 8135 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_456/VPWR
flabel metal1 7600 -8736 7653 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_457/VPWR
flabel metal1 7603 -9278 7654 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_457/VGND
rlabel comment 7675 -9260 7675 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_457/tapvpwrvgnd_1
rlabel metal1 7583 -9308 7675 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_457/VGND
rlabel metal1 7583 -8764 7675 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_457/VPWR
flabel metal1 9268 -9277 9302 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_227/VGND
flabel metal1 9268 -8733 9302 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_227/VPWR
flabel nwell 9268 -8733 9302 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_227/VPB
flabel pwell 9268 -9277 9302 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_227/VNB
rlabel comment 9331 -9260 9331 -9260 6 sky130_fd_sc_hd__decap_4_227/decap_4
rlabel metal1 8963 -9308 9331 -9212 1 sky130_fd_sc_hd__decap_4_227/VGND
rlabel metal1 8963 -8764 9331 -8668 1 sky130_fd_sc_hd__decap_4_227/VPWR
flabel metal1 10648 -9277 10682 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_228/VGND
flabel metal1 10648 -8733 10682 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_228/VPWR
flabel nwell 10648 -8733 10682 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_228/VPB
flabel pwell 10648 -9277 10682 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_228/VNB
rlabel comment 10711 -9260 10711 -9260 6 sky130_fd_sc_hd__decap_4_228/decap_4
rlabel metal1 10343 -9308 10711 -9212 1 sky130_fd_sc_hd__decap_4_228/VGND
rlabel metal1 10343 -8764 10711 -8668 1 sky130_fd_sc_hd__decap_4_228/VPWR
flabel metal1 9452 -8733 9486 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_169/VPWR
flabel metal1 9452 -9277 9486 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_169/VGND
flabel nwell 9452 -8733 9486 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_169/VPB
flabel pwell 9452 -9277 9486 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_169/VNB
rlabel comment 9423 -9260 9423 -9260 4 sky130_fd_sc_hd__decap_8_169/decap_8
rlabel metal1 9423 -9308 10159 -9212 1 sky130_fd_sc_hd__decap_8_169/VGND
rlabel metal1 9423 -8764 10159 -8668 1 sky130_fd_sc_hd__decap_8_169/VPWR
flabel metal1 10285 -8733 10321 -8703 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_64/VPWR
flabel metal1 10285 -9273 10321 -9244 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_64/VGND
flabel nwell 10292 -8726 10312 -8709 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_64/VPB
flabel pwell 10291 -9271 10315 -9249 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_64/VNB
rlabel comment 10343 -9260 10343 -9260 6 sky130_fd_sc_hd__fill_1_64/fill_1
rlabel metal1 10251 -9308 10343 -9212 1 sky130_fd_sc_hd__fill_1_64/VGND
rlabel metal1 10251 -8764 10343 -8668 1 sky130_fd_sc_hd__fill_1_64/VPWR
flabel metal1 8888 -8736 8941 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_458/VPWR
flabel metal1 8891 -9278 8942 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_458/VGND
rlabel comment 8963 -9260 8963 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_458/tapvpwrvgnd_1
rlabel metal1 8871 -9308 8963 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_458/VGND
rlabel metal1 8871 -8764 8963 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_458/VPWR
flabel metal1 9348 -8736 9401 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_459/VPWR
flabel metal1 9351 -9278 9402 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_459/VGND
rlabel comment 9423 -9260 9423 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_459/tapvpwrvgnd_1
rlabel metal1 9331 -9308 9423 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_459/VGND
rlabel metal1 9331 -8764 9423 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_459/VPWR
flabel metal1 10176 -8736 10229 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_460/VPWR
flabel metal1 10179 -9278 10230 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_460/VGND
rlabel comment 10251 -9260 10251 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_460/tapvpwrvgnd_1
rlabel metal1 10159 -9308 10251 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_460/VGND
rlabel metal1 10159 -8764 10251 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_460/VPWR
flabel locali 10741 -9039 10775 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A
flabel locali 11387 -8835 11421 -8801 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X
flabel locali 11387 -8903 11421 -8869 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X
flabel locali 11387 -8971 11421 -8937 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X
flabel locali 11387 -9039 11421 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X
flabel locali 11387 -9107 11421 -9073 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X
flabel locali 11387 -9175 11421 -9141 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X
flabel pwell 10741 -9277 10775 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/VNB
flabel nwell 10741 -8733 10775 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/VPB
flabel metal1 10741 -9277 10775 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/VGND
flabel metal1 10741 -8733 10775 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_186/VPWR
rlabel comment 10711 -9260 10711 -9260 4 sky130_fd_sc_hd__clkdlybuf4s50_1_186/clkdlybuf4s50_1
rlabel metal1 10711 -9308 11447 -9212 1 sky130_fd_sc_hd__clkdlybuf4s50_1_186/VGND
rlabel metal1 10711 -8764 11447 -8668 1 sky130_fd_sc_hd__clkdlybuf4s50_1_186/VPWR
flabel metal1 11936 -9277 11970 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_229/VGND
flabel metal1 11936 -8733 11970 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_229/VPWR
flabel nwell 11936 -8733 11970 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_229/VPB
flabel pwell 11936 -9277 11970 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_229/VNB
rlabel comment 11999 -9260 11999 -9260 6 sky130_fd_sc_hd__decap_4_229/decap_4
rlabel metal1 11631 -9308 11999 -9212 1 sky130_fd_sc_hd__decap_4_229/VGND
rlabel metal1 11631 -8764 11999 -8668 1 sky130_fd_sc_hd__decap_4_229/VPWR
flabel metal1 10653 -8733 10689 -8703 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_65/VPWR
flabel metal1 10653 -9273 10689 -9244 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_65/VGND
flabel nwell 10660 -8726 10680 -8709 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_65/VPB
flabel pwell 10659 -9271 10683 -9249 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_65/VNB
rlabel comment 10711 -9260 10711 -9260 6 sky130_fd_sc_hd__fill_1_65/fill_1
rlabel metal1 10619 -9308 10711 -9212 1 sky130_fd_sc_hd__fill_1_65/VGND
rlabel metal1 10619 -8764 10711 -8668 1 sky130_fd_sc_hd__fill_1_65/VPWR
flabel metal1 11573 -8733 11609 -8703 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_66/VPWR
flabel metal1 11573 -9273 11609 -9244 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_66/VGND
flabel nwell 11580 -8726 11600 -8709 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_66/VPB
flabel pwell 11579 -9271 11603 -9249 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_66/VNB
rlabel comment 11631 -9260 11631 -9260 6 sky130_fd_sc_hd__fill_1_66/fill_1
rlabel metal1 11539 -9308 11631 -9212 1 sky130_fd_sc_hd__fill_1_66/VGND
rlabel metal1 11539 -8764 11631 -8668 1 sky130_fd_sc_hd__fill_1_66/VPWR
flabel metal1 12033 -9270 12056 -9251 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_13/VGND
flabel metal1 12033 -8725 12053 -8708 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_13/VPWR
flabel nwell 12034 -8730 12059 -8704 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_13/VPB
flabel pwell 12034 -9272 12056 -9248 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_13/VNB
rlabel comment 11999 -9260 11999 -9260 4 sky130_fd_sc_hd__fill_4_13/fill_4
rlabel metal1 11999 -9308 12367 -9212 1 sky130_fd_sc_hd__fill_4_13/VGND
rlabel metal1 11999 -8764 12367 -8668 1 sky130_fd_sc_hd__fill_4_13/VPWR
flabel metal1 11464 -8736 11517 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_461/VPWR
flabel metal1 11467 -9278 11518 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_461/VGND
rlabel comment 11539 -9260 11539 -9260 6 sky130_fd_sc_hd__tapvpwrvgnd_1_461/tapvpwrvgnd_1
rlabel metal1 11447 -9308 11539 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_461/VGND
rlabel metal1 11447 -8764 11539 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_461/VPWR
flabel locali 15248 -8971 15282 -8937 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/X
flabel locali 15340 -8971 15374 -8937 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/X
flabel locali 15340 -9039 15374 -9005 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/X
flabel locali 15248 -9039 15282 -9005 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/X
flabel locali 15248 -9107 15282 -9073 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/X
flabel locali 15340 -9107 15374 -9073 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/X
flabel locali 13684 -9107 13718 -9073 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/A
flabel locali 13684 -9039 13718 -9005 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/A
flabel pwell 13684 -9277 13718 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/VNB
flabel pwell 13701 -9260 13701 -9260 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/VNB
flabel nwell 13684 -8733 13718 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/VPB
flabel nwell 13701 -8716 13701 -8716 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/VPB
flabel metal1 13684 -9277 13718 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/VGND
flabel metal1 13684 -8733 13718 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_14/VPWR
rlabel comment 13655 -9260 13655 -9260 4 sky130_fd_sc_hd__clkbuf_16_14/clkbuf_16
rlabel metal1 13655 -9308 15495 -9212 1 sky130_fd_sc_hd__clkbuf_16_14/VGND
rlabel metal1 13655 -8764 15495 -8668 1 sky130_fd_sc_hd__clkbuf_16_14/VPWR
flabel locali 12672 -9039 12706 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/A
flabel locali 12764 -9039 12798 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/A
flabel locali 13040 -9107 13074 -9073 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/Y
flabel locali 12580 -9039 12614 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/A
flabel locali 13040 -8971 13074 -8937 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/Y
flabel locali 12948 -9039 12982 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/A
flabel locali 12856 -9039 12890 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/A
flabel locali 13040 -9039 13074 -9005 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_10/Y
flabel pwell 12488 -9277 12522 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_10/VNB
flabel nwell 12488 -8733 12522 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_10/VPB
flabel metal1 12488 -8733 12522 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_10/VPWR
flabel metal1 12488 -9277 12522 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_10/VGND
rlabel comment 12459 -9260 12459 -9260 4 sky130_fd_sc_hd__clkinv_4_10/clkinv_4
rlabel metal1 12459 -9308 13103 -9212 1 sky130_fd_sc_hd__clkinv_4_10/VGND
rlabel metal1 12459 -8764 13103 -8668 1 sky130_fd_sc_hd__clkinv_4_10/VPWR
flabel metal1 13224 -9277 13258 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_230/VGND
flabel metal1 13224 -8733 13258 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_230/VPWR
flabel nwell 13224 -8733 13258 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_230/VPB
flabel pwell 13224 -9277 13258 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_230/VNB
rlabel comment 13195 -9260 13195 -9260 4 sky130_fd_sc_hd__decap_4_230/decap_4
rlabel metal1 13195 -9308 13563 -9212 1 sky130_fd_sc_hd__decap_4_230/VGND
rlabel metal1 13195 -8764 13563 -8668 1 sky130_fd_sc_hd__decap_4_230/VPWR
flabel metal1 12389 -8736 12442 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_462/VPWR
flabel metal1 12388 -9278 12439 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_462/VGND
rlabel comment 12367 -9260 12367 -9260 4 sky130_fd_sc_hd__tapvpwrvgnd_1_462/tapvpwrvgnd_1
rlabel metal1 12367 -9308 12459 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_462/VGND
rlabel metal1 12367 -8764 12459 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_462/VPWR
flabel metal1 13125 -8736 13178 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_463/VPWR
flabel metal1 13124 -9278 13175 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_463/VGND
rlabel comment 13103 -9260 13103 -9260 4 sky130_fd_sc_hd__tapvpwrvgnd_1_463/tapvpwrvgnd_1
rlabel metal1 13103 -9308 13195 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_463/VGND
rlabel metal1 13103 -8764 13195 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_463/VPWR
flabel metal1 13585 -8736 13638 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_464/VPWR
flabel metal1 13584 -9278 13635 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_464/VGND
rlabel comment 13563 -9260 13563 -9260 4 sky130_fd_sc_hd__tapvpwrvgnd_1_464/tapvpwrvgnd_1
rlabel metal1 13563 -9308 13655 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_464/VGND
rlabel metal1 13563 -8764 13655 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_464/VPWR
flabel metal1 15616 -9277 15650 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_31/VGND
flabel metal1 15616 -8733 15650 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_31/VPWR
flabel nwell 15616 -8733 15650 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_31/VPB
flabel pwell 15616 -9277 15650 -9243 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_31/VNB
rlabel comment 15587 -9260 15587 -9260 4 sky130_fd_sc_hd__decap_12_31/decap_12
rlabel metal1 15587 -9308 16691 -9212 1 sky130_fd_sc_hd__decap_12_31/VGND
rlabel metal1 15587 -8764 16691 -8668 1 sky130_fd_sc_hd__decap_12_31/VPWR
flabel metal1 15517 -8736 15570 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_465/VPWR
flabel metal1 15516 -9278 15567 -9240 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_465/VGND
rlabel comment 15495 -9260 15495 -9260 4 sky130_fd_sc_hd__tapvpwrvgnd_1_465/tapvpwrvgnd_1
rlabel metal1 15495 -9308 15587 -9212 1 sky130_fd_sc_hd__tapvpwrvgnd_1_465/VGND
rlabel metal1 15495 -8764 15587 -8668 1 sky130_fd_sc_hd__tapvpwrvgnd_1_465/VPWR
flabel metal1 -944 -8733 -910 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_41/VPWR
flabel metal1 -944 -8189 -910 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_41/VGND
flabel nwell -944 -8733 -910 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_41/VPB
flabel pwell -944 -8189 -910 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_41/VNB
rlabel comment -881 -8172 -881 -8172 8 sky130_fd_sc_hd__decap_8_41/decap_8
rlabel metal1 -1617 -8220 -881 -8124 5 sky130_fd_sc_hd__decap_8_41/VGND
rlabel metal1 -1617 -8764 -881 -8668 5 sky130_fd_sc_hd__decap_8_41/VPWR
flabel metal1 -2324 -8733 -2290 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_80/VPWR
flabel metal1 -2324 -8189 -2290 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_80/VGND
flabel nwell -2324 -8733 -2290 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_80/VPB
flabel pwell -2324 -8189 -2290 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_80/VNB
rlabel comment -2261 -8172 -2261 -8172 8 sky130_fd_sc_hd__decap_8_80/decap_8
rlabel metal1 -2997 -8220 -2261 -8124 5 sky130_fd_sc_hd__decap_8_80/VGND
rlabel metal1 -2997 -8764 -2261 -8668 5 sky130_fd_sc_hd__decap_8_80/VPWR
flabel metal1 -1690 -8190 -1637 -8158 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_19/VGND
flabel metal1 -1690 -8733 -1638 -8702 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_19/VPWR
flabel nwell -1679 -8725 -1645 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_19/VPB
flabel pwell -1680 -8184 -1648 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_19/VNB
rlabel comment -1617 -8172 -1617 -8172 8 sky130_fd_sc_hd__fill_2_19/fill_2
rlabel metal1 -1801 -8220 -1617 -8124 5 sky130_fd_sc_hd__fill_2_19/VGND
rlabel metal1 -1801 -8764 -1617 -8668 5 sky130_fd_sc_hd__fill_2_19/VPWR
flabel metal1 -1858 -8181 -1835 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_29/VGND
flabel metal1 -1855 -8724 -1835 -8707 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_29/VPWR
flabel nwell -1861 -8728 -1836 -8702 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_29/VPB
flabel pwell -1858 -8184 -1836 -8160 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_29/VNB
rlabel comment -1801 -8172 -1801 -8172 8 sky130_fd_sc_hd__fill_4_29/fill_4
rlabel metal1 -2169 -8220 -1801 -8124 5 sky130_fd_sc_hd__fill_4_29/VGND
rlabel metal1 -2169 -8764 -1801 -8668 5 sky130_fd_sc_hd__fill_4_29/VPWR
flabel metal1 -2244 -8725 -2191 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_545/VPWR
flabel metal1 -2241 -8192 -2190 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_545/VGND
rlabel comment -2169 -8172 -2169 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_545/tapvpwrvgnd_1
rlabel metal1 -2261 -8220 -2169 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_545/VGND
rlabel metal1 -2261 -8764 -2169 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_545/VPWR
flabel locali 1079 -8427 1113 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/A
flabel locali 433 -8631 467 -8597 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
flabel locali 433 -8563 467 -8529 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
flabel locali 433 -8495 467 -8461 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
flabel locali 433 -8427 467 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
flabel locali 433 -8359 467 -8325 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
flabel locali 433 -8291 467 -8257 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
flabel pwell 1079 -8189 1113 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/VNB
flabel nwell 1079 -8733 1113 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/VPB
flabel metal1 1079 -8189 1113 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/VGND
flabel metal1 1079 -8733 1113 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_187/VPWR
rlabel comment 1143 -8172 1143 -8172 8 sky130_fd_sc_hd__clkdlybuf4s50_1_187/clkdlybuf4s50_1
rlabel metal1 407 -8220 1143 -8124 5 sky130_fd_sc_hd__clkdlybuf4s50_1_187/VGND
rlabel metal1 407 -8764 1143 -8668 5 sky130_fd_sc_hd__clkdlybuf4s50_1_187/VPWR
flabel metal1 252 -8189 286 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_231/VGND
flabel metal1 252 -8733 286 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_231/VPWR
flabel nwell 252 -8733 286 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_231/VPB
flabel pwell 252 -8189 286 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_231/VNB
rlabel comment 315 -8172 315 -8172 8 sky130_fd_sc_hd__decap_4_231/decap_4
rlabel metal1 -53 -8220 315 -8124 5 sky130_fd_sc_hd__decap_4_231/VGND
rlabel metal1 -53 -8764 315 -8668 5 sky130_fd_sc_hd__decap_4_231/VPWR
flabel metal1 -208 -8733 -174 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_42/VPWR
flabel metal1 -208 -8189 -174 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_42/VGND
flabel nwell -208 -8733 -174 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_42/VPB
flabel pwell -208 -8189 -174 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_42/VNB
rlabel comment -145 -8172 -145 -8172 8 sky130_fd_sc_hd__decap_8_42/decap_8
rlabel metal1 -881 -8220 -145 -8124 5 sky130_fd_sc_hd__decap_8_42/VGND
rlabel metal1 -881 -8764 -145 -8668 5 sky130_fd_sc_hd__decap_8_42/VPWR
flabel metal1 332 -8725 385 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_466/VPWR
flabel metal1 335 -8192 386 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_466/VGND
rlabel comment 407 -8172 407 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_466/tapvpwrvgnd_1
rlabel metal1 315 -8220 407 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_466/VGND
rlabel metal1 315 -8764 407 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_466/VPWR
flabel metal1 -128 -8725 -75 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_467/VPWR
flabel metal1 -125 -8192 -74 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_467/VGND
rlabel comment -53 -8172 -53 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_467/tapvpwrvgnd_1
rlabel metal1 -145 -8220 -53 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_467/VGND
rlabel metal1 -145 -8764 -53 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_467/VPWR
flabel metal1 1540 -8189 1574 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_232/VGND
flabel metal1 1540 -8733 1574 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_232/VPWR
flabel nwell 1540 -8733 1574 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_232/VPB
flabel pwell 1540 -8189 1574 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_232/VNB
rlabel comment 1603 -8172 1603 -8172 8 sky130_fd_sc_hd__decap_4_232/decap_4
rlabel metal1 1235 -8220 1603 -8124 5 sky130_fd_sc_hd__decap_4_232/VGND
rlabel metal1 1235 -8764 1603 -8668 5 sky130_fd_sc_hd__decap_4_232/VPWR
flabel metal1 2828 -8189 2862 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_233/VGND
flabel metal1 2828 -8733 2862 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_233/VPWR
flabel nwell 2828 -8733 2862 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_233/VPB
flabel pwell 2828 -8189 2862 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_233/VNB
rlabel comment 2891 -8172 2891 -8172 8 sky130_fd_sc_hd__decap_4_233/decap_4
rlabel metal1 2523 -8220 2891 -8124 5 sky130_fd_sc_hd__decap_4_233/VGND
rlabel metal1 2523 -8764 2891 -8668 5 sky130_fd_sc_hd__decap_4_233/VPWR
flabel metal1 2368 -8733 2402 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_131/VPWR
flabel metal1 2368 -8189 2402 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_131/VGND
flabel nwell 2368 -8733 2402 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_131/VPB
flabel pwell 2368 -8189 2402 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_131/VNB
rlabel comment 2431 -8172 2431 -8172 8 sky130_fd_sc_hd__decap_8_131/decap_8
rlabel metal1 1695 -8220 2431 -8124 5 sky130_fd_sc_hd__decap_8_131/VGND
rlabel metal1 1695 -8764 2431 -8668 5 sky130_fd_sc_hd__decap_8_131/VPWR
flabel metal1 1620 -8725 1673 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_468/VPWR
flabel metal1 1623 -8192 1674 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_468/VGND
rlabel comment 1695 -8172 1695 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_468/tapvpwrvgnd_1
rlabel metal1 1603 -8220 1695 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_468/VGND
rlabel metal1 1603 -8764 1695 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_468/VPWR
flabel metal1 1160 -8725 1213 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_469/VPWR
flabel metal1 1163 -8192 1214 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_469/VGND
rlabel comment 1235 -8172 1235 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_469/tapvpwrvgnd_1
rlabel metal1 1143 -8220 1235 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_469/VGND
rlabel metal1 1143 -8764 1235 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_469/VPWR
flabel metal1 2448 -8725 2501 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_470/VPWR
flabel metal1 2451 -8192 2502 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_470/VGND
rlabel comment 2523 -8172 2523 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_470/tapvpwrvgnd_1
rlabel metal1 2431 -8220 2523 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_470/VGND
rlabel metal1 2431 -8764 2523 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_470/VPWR
flabel locali 3655 -8427 3689 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A
flabel locali 3009 -8631 3043 -8597 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X
flabel locali 3009 -8563 3043 -8529 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X
flabel locali 3009 -8495 3043 -8461 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X
flabel locali 3009 -8427 3043 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X
flabel locali 3009 -8359 3043 -8325 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X
flabel locali 3009 -8291 3043 -8257 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X
flabel pwell 3655 -8189 3689 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/VNB
flabel nwell 3655 -8733 3689 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/VPB
flabel metal1 3655 -8189 3689 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/VGND
flabel metal1 3655 -8733 3689 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_190/VPWR
rlabel comment 3719 -8172 3719 -8172 8 sky130_fd_sc_hd__clkdlybuf4s50_1_190/clkdlybuf4s50_1
rlabel metal1 2983 -8220 3719 -8124 5 sky130_fd_sc_hd__clkdlybuf4s50_1_190/VGND
rlabel metal1 2983 -8764 3719 -8668 5 sky130_fd_sc_hd__clkdlybuf4s50_1_190/VPWR
flabel metal1 4116 -8189 4150 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_234/VGND
flabel metal1 4116 -8733 4150 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_234/VPWR
flabel nwell 4116 -8733 4150 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_234/VPB
flabel pwell 4116 -8189 4150 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_234/VNB
rlabel comment 4179 -8172 4179 -8172 8 sky130_fd_sc_hd__decap_4_234/decap_4
rlabel metal1 3811 -8220 4179 -8124 5 sky130_fd_sc_hd__decap_4_234/VGND
rlabel metal1 3811 -8764 4179 -8668 5 sky130_fd_sc_hd__decap_4_234/VPWR
flabel metal1 4944 -8733 4978 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_149/VPWR
flabel metal1 4944 -8189 4978 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_149/VGND
flabel nwell 4944 -8733 4978 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_149/VPB
flabel pwell 4944 -8189 4978 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_149/VNB
rlabel comment 5007 -8172 5007 -8172 8 sky130_fd_sc_hd__decap_8_149/decap_8
rlabel metal1 4271 -8220 5007 -8124 5 sky130_fd_sc_hd__decap_8_149/VGND
rlabel metal1 4271 -8764 5007 -8668 5 sky130_fd_sc_hd__decap_8_149/VPWR
flabel metal1 4196 -8725 4249 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_471/VPWR
flabel metal1 4199 -8192 4250 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_471/VGND
rlabel comment 4271 -8172 4271 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_471/tapvpwrvgnd_1
rlabel metal1 4179 -8220 4271 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_471/VGND
rlabel metal1 4179 -8764 4271 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_471/VPWR
flabel metal1 2908 -8725 2961 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_472/VPWR
flabel metal1 2911 -8192 2962 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_472/VGND
rlabel comment 2983 -8172 2983 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_472/tapvpwrvgnd_1
rlabel metal1 2891 -8220 2983 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_472/VGND
rlabel metal1 2891 -8764 2983 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_472/VPWR
flabel metal1 3736 -8725 3789 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_473/VPWR
flabel metal1 3739 -8192 3790 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_473/VGND
rlabel comment 3811 -8172 3811 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_473/tapvpwrvgnd_1
rlabel metal1 3719 -8220 3811 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_473/VGND
rlabel metal1 3719 -8764 3811 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_473/VPWR
flabel locali 6231 -8427 6265 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/A
flabel locali 5585 -8631 5619 -8597 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
flabel locali 5585 -8563 5619 -8529 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
flabel locali 5585 -8495 5619 -8461 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
flabel locali 5585 -8427 5619 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
flabel locali 5585 -8359 5619 -8325 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
flabel locali 5585 -8291 5619 -8257 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X
flabel pwell 6231 -8189 6265 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/VNB
flabel nwell 6231 -8733 6265 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/VPB
flabel metal1 6231 -8189 6265 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/VGND
flabel metal1 6231 -8733 6265 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_191/VPWR
rlabel comment 6295 -8172 6295 -8172 8 sky130_fd_sc_hd__clkdlybuf4s50_1_191/clkdlybuf4s50_1
rlabel metal1 5559 -8220 6295 -8124 5 sky130_fd_sc_hd__clkdlybuf4s50_1_191/VGND
rlabel metal1 5559 -8764 6295 -8668 5 sky130_fd_sc_hd__clkdlybuf4s50_1_191/VPWR
flabel metal1 6692 -8189 6726 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_235/VGND
flabel metal1 6692 -8733 6726 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_235/VPWR
flabel nwell 6692 -8733 6726 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_235/VPB
flabel pwell 6692 -8189 6726 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_235/VNB
rlabel comment 6755 -8172 6755 -8172 8 sky130_fd_sc_hd__decap_4_235/decap_4
rlabel metal1 6387 -8220 6755 -8124 5 sky130_fd_sc_hd__decap_4_235/VGND
rlabel metal1 6387 -8764 6755 -8668 5 sky130_fd_sc_hd__decap_4_235/VPWR
flabel metal1 5404 -8189 5438 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_236/VGND
flabel metal1 5404 -8733 5438 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_236/VPWR
flabel nwell 5404 -8733 5438 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_236/VPB
flabel pwell 5404 -8189 5438 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_236/VNB
rlabel comment 5467 -8172 5467 -8172 8 sky130_fd_sc_hd__decap_4_236/decap_4
rlabel metal1 5099 -8220 5467 -8124 5 sky130_fd_sc_hd__decap_4_236/VGND
rlabel metal1 5099 -8764 5467 -8668 5 sky130_fd_sc_hd__decap_4_236/VPWR
flabel metal1 6312 -8725 6365 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_474/VPWR
flabel metal1 6315 -8192 6366 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_474/VGND
rlabel comment 6387 -8172 6387 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_474/tapvpwrvgnd_1
rlabel metal1 6295 -8220 6387 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_474/VGND
rlabel metal1 6295 -8764 6387 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_474/VPWR
flabel metal1 5484 -8725 5537 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_475/VPWR
flabel metal1 5487 -8192 5538 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_475/VGND
rlabel comment 5559 -8172 5559 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_475/tapvpwrvgnd_1
rlabel metal1 5467 -8220 5559 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_475/VGND
rlabel metal1 5467 -8764 5559 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_475/VPWR
flabel metal1 5024 -8725 5077 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_476/VPWR
flabel metal1 5027 -8192 5078 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_476/VGND
rlabel comment 5099 -8172 5099 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_476/tapvpwrvgnd_1
rlabel metal1 5007 -8220 5099 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_476/VGND
rlabel metal1 5007 -8764 5099 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_476/VPWR
flabel locali 8807 -8427 8841 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/A
flabel locali 8161 -8631 8195 -8597 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X
flabel locali 8161 -8563 8195 -8529 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X
flabel locali 8161 -8495 8195 -8461 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X
flabel locali 8161 -8427 8195 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X
flabel locali 8161 -8359 8195 -8325 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X
flabel locali 8161 -8291 8195 -8257 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X
flabel pwell 8807 -8189 8841 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/VNB
flabel nwell 8807 -8733 8841 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/VPB
flabel metal1 8807 -8189 8841 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/VGND
flabel metal1 8807 -8733 8841 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_193/VPWR
rlabel comment 8871 -8172 8871 -8172 8 sky130_fd_sc_hd__clkdlybuf4s50_1_193/clkdlybuf4s50_1
rlabel metal1 8135 -8220 8871 -8124 5 sky130_fd_sc_hd__clkdlybuf4s50_1_193/VGND
rlabel metal1 8135 -8764 8871 -8668 5 sky130_fd_sc_hd__clkdlybuf4s50_1_193/VPWR
flabel metal1 7980 -8189 8014 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_237/VGND
flabel metal1 7980 -8733 8014 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_237/VPWR
flabel nwell 7980 -8733 8014 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_237/VPB
flabel pwell 7980 -8189 8014 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_237/VNB
rlabel comment 8043 -8172 8043 -8172 8 sky130_fd_sc_hd__decap_4_237/decap_4
rlabel metal1 7675 -8220 8043 -8124 5 sky130_fd_sc_hd__decap_4_237/VGND
rlabel metal1 7675 -8764 8043 -8668 5 sky130_fd_sc_hd__decap_4_237/VPWR
flabel metal1 7520 -8733 7554 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_160/VPWR
flabel metal1 7520 -8189 7554 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_160/VGND
flabel nwell 7520 -8733 7554 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_160/VPB
flabel pwell 7520 -8189 7554 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_160/VNB
rlabel comment 7583 -8172 7583 -8172 8 sky130_fd_sc_hd__decap_8_160/decap_8
rlabel metal1 6847 -8220 7583 -8124 5 sky130_fd_sc_hd__decap_8_160/VGND
rlabel metal1 6847 -8764 7583 -8668 5 sky130_fd_sc_hd__decap_8_160/VPWR
flabel metal1 6772 -8725 6825 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_477/VPWR
flabel metal1 6775 -8192 6826 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_477/VGND
rlabel comment 6847 -8172 6847 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_477/tapvpwrvgnd_1
rlabel metal1 6755 -8220 6847 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_477/VGND
rlabel metal1 6755 -8764 6847 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_477/VPWR
flabel metal1 8060 -8725 8113 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_478/VPWR
flabel metal1 8063 -8192 8114 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_478/VGND
rlabel comment 8135 -8172 8135 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_478/tapvpwrvgnd_1
rlabel metal1 8043 -8220 8135 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_478/VGND
rlabel metal1 8043 -8764 8135 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_478/VPWR
flabel metal1 7600 -8725 7653 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_479/VPWR
flabel metal1 7603 -8192 7654 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_479/VGND
rlabel comment 7675 -8172 7675 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_479/tapvpwrvgnd_1
rlabel metal1 7583 -8220 7675 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_479/VGND
rlabel metal1 7583 -8764 7675 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_479/VPWR
flabel metal1 9268 -8189 9302 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_238/VGND
flabel metal1 9268 -8733 9302 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_238/VPWR
flabel nwell 9268 -8733 9302 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_238/VPB
flabel pwell 9268 -8189 9302 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_238/VNB
rlabel comment 9331 -8172 9331 -8172 8 sky130_fd_sc_hd__decap_4_238/decap_4
rlabel metal1 8963 -8220 9331 -8124 5 sky130_fd_sc_hd__decap_4_238/VGND
rlabel metal1 8963 -8764 9331 -8668 5 sky130_fd_sc_hd__decap_4_238/VPWR
flabel metal1 10648 -8189 10682 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_240/VGND
flabel metal1 10648 -8733 10682 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_240/VPWR
flabel nwell 10648 -8733 10682 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_240/VPB
flabel pwell 10648 -8189 10682 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_240/VNB
rlabel comment 10711 -8172 10711 -8172 8 sky130_fd_sc_hd__decap_4_240/decap_4
rlabel metal1 10343 -8220 10711 -8124 5 sky130_fd_sc_hd__decap_4_240/VGND
rlabel metal1 10343 -8764 10711 -8668 5 sky130_fd_sc_hd__decap_4_240/VPWR
flabel metal1 10096 -8733 10130 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_170/VPWR
flabel metal1 10096 -8189 10130 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_170/VGND
flabel nwell 10096 -8733 10130 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_170/VPB
flabel pwell 10096 -8189 10130 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_170/VNB
rlabel comment 10159 -8172 10159 -8172 8 sky130_fd_sc_hd__decap_8_170/decap_8
rlabel metal1 9423 -8220 10159 -8124 5 sky130_fd_sc_hd__decap_8_170/VGND
rlabel metal1 9423 -8764 10159 -8668 5 sky130_fd_sc_hd__decap_8_170/VPWR
flabel metal1 10285 -8729 10321 -8699 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_67/VPWR
flabel metal1 10285 -8188 10321 -8159 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_67/VGND
flabel nwell 10292 -8723 10312 -8706 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_67/VPB
flabel pwell 10291 -8183 10315 -8161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_67/VNB
rlabel comment 10343 -8172 10343 -8172 8 sky130_fd_sc_hd__fill_1_67/fill_1
rlabel metal1 10251 -8220 10343 -8124 5 sky130_fd_sc_hd__fill_1_67/VGND
rlabel metal1 10251 -8764 10343 -8668 5 sky130_fd_sc_hd__fill_1_67/VPWR
flabel metal1 8888 -8725 8941 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_480/VPWR
flabel metal1 8891 -8192 8942 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_480/VGND
rlabel comment 8963 -8172 8963 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_480/tapvpwrvgnd_1
rlabel metal1 8871 -8220 8963 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_480/VGND
rlabel metal1 8871 -8764 8963 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_480/VPWR
flabel metal1 9348 -8725 9401 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_481/VPWR
flabel metal1 9351 -8192 9402 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_481/VGND
rlabel comment 9423 -8172 9423 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_481/tapvpwrvgnd_1
rlabel metal1 9331 -8220 9423 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_481/VGND
rlabel metal1 9331 -8764 9423 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_481/VPWR
flabel metal1 10176 -8725 10229 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_482/VPWR
flabel metal1 10179 -8192 10230 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_482/VGND
rlabel comment 10251 -8172 10251 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_482/tapvpwrvgnd_1
rlabel metal1 10159 -8220 10251 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_482/VGND
rlabel metal1 10159 -8764 10251 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_482/VPWR
flabel locali 11383 -8427 11417 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A
flabel locali 10737 -8631 10771 -8597 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
flabel locali 10737 -8563 10771 -8529 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
flabel locali 10737 -8495 10771 -8461 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
flabel locali 10737 -8427 10771 -8393 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
flabel locali 10737 -8359 10771 -8325 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
flabel locali 10737 -8291 10771 -8257 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
flabel pwell 11383 -8189 11417 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/VNB
flabel nwell 11383 -8733 11417 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/VPB
flabel metal1 11383 -8189 11417 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/VGND
flabel metal1 11383 -8733 11417 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_195/VPWR
rlabel comment 11447 -8172 11447 -8172 8 sky130_fd_sc_hd__clkdlybuf4s50_1_195/clkdlybuf4s50_1
rlabel metal1 10711 -8220 11447 -8124 5 sky130_fd_sc_hd__clkdlybuf4s50_1_195/VGND
rlabel metal1 10711 -8764 11447 -8668 5 sky130_fd_sc_hd__clkdlybuf4s50_1_195/VPWR
flabel metal1 11936 -8189 11970 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_239/VGND
flabel metal1 11936 -8733 11970 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_239/VPWR
flabel nwell 11936 -8733 11970 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_239/VPB
flabel pwell 11936 -8189 11970 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_239/VNB
rlabel comment 11999 -8172 11999 -8172 8 sky130_fd_sc_hd__decap_4_239/decap_4
rlabel metal1 11631 -8220 11999 -8124 5 sky130_fd_sc_hd__decap_4_239/VGND
rlabel metal1 11631 -8764 11999 -8668 5 sky130_fd_sc_hd__decap_4_239/VPWR
flabel metal1 11573 -8729 11609 -8699 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_68/VPWR
flabel metal1 11573 -8188 11609 -8159 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_68/VGND
flabel nwell 11580 -8723 11600 -8706 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_68/VPB
flabel pwell 11579 -8183 11603 -8161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_68/VNB
rlabel comment 11631 -8172 11631 -8172 8 sky130_fd_sc_hd__fill_1_68/fill_1
rlabel metal1 11539 -8220 11631 -8124 5 sky130_fd_sc_hd__fill_1_68/VGND
rlabel metal1 11539 -8764 11631 -8668 5 sky130_fd_sc_hd__fill_1_68/VPWR
flabel metal1 10653 -8729 10689 -8699 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_69/VPWR
flabel metal1 10653 -8188 10689 -8159 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_69/VGND
flabel nwell 10660 -8723 10680 -8706 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_69/VPB
flabel pwell 10659 -8183 10683 -8161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_69/VNB
rlabel comment 10711 -8172 10711 -8172 8 sky130_fd_sc_hd__fill_1_69/fill_1
rlabel metal1 10619 -8220 10711 -8124 5 sky130_fd_sc_hd__fill_1_69/VGND
rlabel metal1 10619 -8764 10711 -8668 5 sky130_fd_sc_hd__fill_1_69/VPWR
flabel metal1 12668 -8182 12700 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_31/VGND
flabel metal1 12668 -8727 12706 -8695 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_31/VPWR
flabel nwell 12658 -8725 12715 -8694 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_31/VPB
flabel pwell 12665 -8182 12709 -8148 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_31/VNB
rlabel comment 12735 -8172 12735 -8172 8 sky130_fd_sc_hd__fill_8_31/fill_8
rlabel metal1 11999 -8220 12735 -8124 5 sky130_fd_sc_hd__fill_8_31/VGND
rlabel metal1 11999 -8764 12735 -8668 5 sky130_fd_sc_hd__fill_8_31/VPWR
flabel metal1 11464 -8725 11517 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_483/VPWR
flabel metal1 11467 -8192 11518 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_483/VGND
rlabel comment 11539 -8172 11539 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_483/tapvpwrvgnd_1
rlabel metal1 11447 -8220 11539 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_483/VGND
rlabel metal1 11447 -8764 11539 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_483/VPWR
flabel locali 15248 -8495 15282 -8461 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/X
flabel locali 15340 -8495 15374 -8461 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/X
flabel locali 15340 -8427 15374 -8393 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/X
flabel locali 15248 -8427 15282 -8393 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/X
flabel locali 15248 -8359 15282 -8325 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/X
flabel locali 15340 -8359 15374 -8325 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/X
flabel locali 13684 -8359 13718 -8325 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/A
flabel locali 13684 -8427 13718 -8393 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/A
flabel pwell 13684 -8189 13718 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/VNB
flabel pwell 13701 -8172 13701 -8172 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/VNB
flabel nwell 13684 -8733 13718 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/VPB
flabel nwell 13701 -8716 13701 -8716 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/VPB
flabel metal1 13684 -8189 13718 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/VGND
flabel metal1 13684 -8733 13718 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_15/VPWR
rlabel comment 13655 -8172 13655 -8172 2 sky130_fd_sc_hd__clkbuf_16_15/clkbuf_16
rlabel metal1 13655 -8220 15495 -8124 5 sky130_fd_sc_hd__clkbuf_16_15/VGND
rlabel metal1 13655 -8764 15495 -8668 5 sky130_fd_sc_hd__clkbuf_16_15/VPWR
flabel metal1 13505 -8729 13541 -8699 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_70/VPWR
flabel metal1 13505 -8188 13541 -8159 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_70/VGND
flabel nwell 13512 -8723 13532 -8706 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_70/VPB
flabel pwell 13511 -8183 13535 -8161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_70/VNB
rlabel comment 13563 -8172 13563 -8172 8 sky130_fd_sc_hd__fill_1_70/fill_1
rlabel metal1 13471 -8220 13563 -8124 5 sky130_fd_sc_hd__fill_1_70/VGND
rlabel metal1 13471 -8764 13563 -8668 5 sky130_fd_sc_hd__fill_1_70/VPWR
flabel metal1 13404 -8182 13436 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_32/VGND
flabel metal1 13404 -8727 13442 -8695 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_32/VPWR
flabel nwell 13394 -8725 13451 -8694 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_32/VPB
flabel pwell 13401 -8182 13445 -8148 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_32/VNB
rlabel comment 13471 -8172 13471 -8172 8 sky130_fd_sc_hd__fill_8_32/fill_8
rlabel metal1 12735 -8220 13471 -8124 5 sky130_fd_sc_hd__fill_8_32/VGND
rlabel metal1 12735 -8764 13471 -8668 5 sky130_fd_sc_hd__fill_8_32/VPWR
flabel metal1 13580 -8725 13633 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_484/VPWR
flabel metal1 13583 -8192 13634 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_484/VGND
rlabel comment 13655 -8172 13655 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_484/tapvpwrvgnd_1
rlabel metal1 13563 -8220 13655 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_484/VGND
rlabel metal1 13563 -8764 13655 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_484/VPWR
flabel metal1 16628 -8189 16662 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_32/VGND
flabel metal1 16628 -8733 16662 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_32/VPWR
flabel nwell 16628 -8733 16662 -8699 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_32/VPB
flabel pwell 16628 -8189 16662 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_32/VNB
rlabel comment 16691 -8172 16691 -8172 8 sky130_fd_sc_hd__decap_12_32/decap_12
rlabel metal1 15587 -8220 16691 -8124 5 sky130_fd_sc_hd__decap_12_32/VGND
rlabel metal1 15587 -8764 16691 -8668 5 sky130_fd_sc_hd__decap_12_32/VPWR
flabel metal1 15512 -8725 15565 -8696 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_485/VPWR
flabel metal1 15515 -8192 15566 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_485/VGND
rlabel comment 15587 -8172 15587 -8172 8 sky130_fd_sc_hd__tapvpwrvgnd_1_485/tapvpwrvgnd_1
rlabel metal1 15495 -8220 15587 -8124 5 sky130_fd_sc_hd__tapvpwrvgnd_1_485/VGND
rlabel metal1 15495 -8764 15587 -8668 5 sky130_fd_sc_hd__tapvpwrvgnd_1_485/VPWR
flabel metal1 -1404 -8189 -1370 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_241/VGND
flabel metal1 -1404 -7645 -1370 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_241/VPWR
flabel nwell -1404 -7645 -1370 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_241/VPB
flabel pwell -1404 -8189 -1370 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_241/VNB
rlabel comment -1433 -8172 -1433 -8172 4 sky130_fd_sc_hd__decap_4_241/decap_4
rlabel metal1 -1433 -8220 -1065 -8124 1 sky130_fd_sc_hd__decap_4_241/VGND
rlabel metal1 -1433 -7676 -1065 -7580 1 sky130_fd_sc_hd__decap_4_241/VPWR
flabel metal1 -2968 -7645 -2934 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_79/VPWR
flabel metal1 -2968 -8189 -2934 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_79/VGND
flabel nwell -2968 -7645 -2934 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_79/VPB
flabel pwell -2968 -8189 -2934 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_79/VNB
rlabel comment -2997 -8172 -2997 -8172 4 sky130_fd_sc_hd__decap_8_79/decap_8
rlabel metal1 -2997 -8220 -2261 -8124 1 sky130_fd_sc_hd__decap_8_79/VGND
rlabel metal1 -2997 -7676 -2261 -7580 1 sky130_fd_sc_hd__decap_8_79/VPWR
flabel metal1 -1597 -8186 -1544 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_3/VGND
flabel metal1 -1596 -7642 -1544 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_3/VPWR
flabel nwell -1589 -7637 -1555 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_3/VPB
flabel pwell -1586 -8182 -1554 -8160 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_3/VNB
rlabel comment -1617 -8172 -1617 -8172 4 sky130_fd_sc_hd__fill_2_3/fill_2
rlabel metal1 -1617 -8220 -1433 -8124 1 sky130_fd_sc_hd__fill_2_3/VGND
rlabel metal1 -1617 -7676 -1433 -7580 1 sky130_fd_sc_hd__fill_2_3/VPWR
flabel metal1 -1781 -8186 -1728 -8154 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_18/VGND
flabel metal1 -1780 -7642 -1728 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_18/VPWR
flabel nwell -1773 -7637 -1739 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_18/VPB
flabel pwell -1770 -8182 -1738 -8160 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_18/VNB
rlabel comment -1801 -8172 -1801 -8172 4 sky130_fd_sc_hd__fill_2_18/fill_2
rlabel metal1 -1801 -8220 -1617 -8124 1 sky130_fd_sc_hd__fill_2_18/VGND
rlabel metal1 -1801 -7676 -1617 -7580 1 sky130_fd_sc_hd__fill_2_18/VPWR
flabel metal1 -2135 -8182 -2112 -8163 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_28/VGND
flabel metal1 -2135 -7637 -2115 -7620 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_28/VPWR
flabel nwell -2134 -7642 -2109 -7616 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_28/VPB
flabel pwell -2134 -8184 -2112 -8160 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_28/VNB
rlabel comment -2169 -8172 -2169 -8172 4 sky130_fd_sc_hd__fill_4_28/fill_4
rlabel metal1 -2169 -8220 -1801 -8124 1 sky130_fd_sc_hd__fill_4_28/VGND
rlabel metal1 -2169 -7676 -1801 -7580 1 sky130_fd_sc_hd__fill_4_28/VPWR
flabel metal1 -2239 -7648 -2186 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_544/VPWR
flabel metal1 -2240 -8190 -2189 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_544/VGND
rlabel comment -2261 -8172 -2261 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_544/tapvpwrvgnd_1
rlabel metal1 -2261 -8220 -2169 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_544/VGND
rlabel metal1 -2261 -7676 -2169 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_544/VPWR
flabel locali 68 -7951 102 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/A
flabel locali 160 -7951 194 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/A
flabel locali 436 -8019 470 -7985 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/Y
flabel locali -24 -7951 10 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/A
flabel locali 436 -7883 470 -7849 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/Y
flabel locali 344 -7951 378 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/A
flabel locali 252 -7951 286 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/A
flabel locali 436 -7951 470 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_11/Y
flabel pwell -116 -8189 -82 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_11/VNB
flabel nwell -116 -7645 -82 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_11/VPB
flabel metal1 -116 -7645 -82 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_11/VPWR
flabel metal1 -116 -8189 -82 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_11/VGND
rlabel comment -145 -8172 -145 -8172 4 sky130_fd_sc_hd__clkinv_4_11/clkinv_4
rlabel metal1 -145 -8220 499 -8124 1 sky130_fd_sc_hd__clkinv_4_11/VGND
rlabel metal1 -145 -7676 499 -7580 1 sky130_fd_sc_hd__clkinv_4_11/VPWR
flabel metal1 620 -8189 654 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_242/VGND
flabel metal1 620 -7645 654 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_242/VPWR
flabel nwell 620 -7645 654 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_242/VPB
flabel pwell 620 -8189 654 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_242/VNB
rlabel comment 591 -8172 591 -8172 4 sky130_fd_sc_hd__decap_4_242/decap_4
rlabel metal1 591 -8220 959 -8124 1 sky130_fd_sc_hd__decap_4_242/VGND
rlabel metal1 591 -7676 959 -7580 1 sky130_fd_sc_hd__decap_4_242/VPWR
flabel metal1 -576 -8189 -542 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_243/VGND
flabel metal1 -576 -7645 -542 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_243/VPWR
flabel nwell -576 -7645 -542 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_243/VPB
flabel pwell -576 -8189 -542 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_243/VNB
rlabel comment -605 -8172 -605 -8172 4 sky130_fd_sc_hd__decap_4_243/decap_4
rlabel metal1 -605 -8220 -237 -8124 1 sky130_fd_sc_hd__decap_4_243/VGND
rlabel metal1 -605 -7676 -237 -7580 1 sky130_fd_sc_hd__decap_4_243/VPWR
flabel locali -853 -8087 -819 -8053 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/Y
flabel locali -853 -8019 -819 -7985 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/Y
flabel locali -853 -7951 -819 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/Y
flabel locali -945 -7951 -911 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/B
flabel locali -761 -7951 -727 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/A
flabel nwell -945 -7645 -911 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VPB
flabel pwell -945 -8189 -911 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VNB
flabel metal1 -945 -8189 -911 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VGND
flabel metal1 -945 -7645 -911 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VPWR
rlabel comment -973 -8172 -973 -8172 4 sky130_fd_sc_hd__nand2_1_3/nand2_1
rlabel metal1 -973 -8220 -697 -8124 1 sky130_fd_sc_hd__nand2_1_3/VGND
rlabel metal1 -973 -7676 -697 -7580 1 sky130_fd_sc_hd__nand2_1_3/VPWR
flabel metal1 521 -7648 574 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_486/VPWR
flabel metal1 520 -8190 571 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_486/VGND
rlabel comment 499 -8172 499 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_486/tapvpwrvgnd_1
rlabel metal1 499 -8220 591 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_486/VGND
rlabel metal1 499 -7676 591 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_486/VPWR
flabel metal1 -215 -7648 -162 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_487/VPWR
flabel metal1 -216 -8190 -165 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_487/VGND
rlabel comment -237 -8172 -237 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_487/tapvpwrvgnd_1
rlabel metal1 -237 -8220 -145 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_487/VGND
rlabel metal1 -237 -7676 -145 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_487/VPWR
flabel metal1 -675 -7648 -622 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_488/VPWR
flabel metal1 -676 -8190 -625 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_488/VGND
rlabel comment -697 -8172 -697 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_488/tapvpwrvgnd_1
rlabel metal1 -697 -8220 -605 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_488/VGND
rlabel metal1 -697 -7676 -605 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_488/VPWR
flabel metal1 -1043 -7648 -990 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_489/VPWR
flabel metal1 -1044 -8190 -993 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_489/VGND
rlabel comment -1065 -8172 -1065 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_489/tapvpwrvgnd_1
rlabel metal1 -1065 -8220 -973 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_489/VGND
rlabel metal1 -1065 -7676 -973 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_489/VPWR
flabel locali 2369 -7951 2403 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/A
flabel locali 3015 -7747 3049 -7713 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/X
flabel locali 3015 -7815 3049 -7781 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/X
flabel locali 3015 -7883 3049 -7849 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/X
flabel locali 3015 -7951 3049 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/X
flabel locali 3015 -8019 3049 -7985 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/X
flabel locali 3015 -8087 3049 -8053 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/X
flabel pwell 2369 -8189 2403 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/VNB
flabel nwell 2369 -7645 2403 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/VPB
flabel metal1 2369 -8189 2403 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/VGND
flabel metal1 2369 -7645 2403 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_196/VPWR
rlabel comment 2339 -8172 2339 -8172 4 sky130_fd_sc_hd__clkdlybuf4s50_1_196/clkdlybuf4s50_1
rlabel metal1 2339 -8220 3075 -8124 1 sky130_fd_sc_hd__clkdlybuf4s50_1_196/VGND
rlabel metal1 2339 -7676 3075 -7580 1 sky130_fd_sc_hd__clkdlybuf4s50_1_196/VPWR
flabel locali 1264 -8019 1298 -7985 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/Y
flabel locali 1264 -7951 1298 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/Y
flabel locali 1172 -7883 1206 -7849 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/Y
flabel locali 1172 -7951 1206 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/Y
flabel locali 1172 -8019 1206 -7985 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/Y
flabel locali 1080 -8087 1114 -8053 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/A
flabel locali 1080 -8019 1114 -7985 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/A
flabel locali 1080 -7951 1114 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_3/A
flabel nwell 1080 -7645 1114 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_3/VPB
flabel pwell 1080 -8189 1114 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_3/VNB
flabel metal1 1080 -8189 1114 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_3/VGND
flabel metal1 1080 -7645 1114 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_3/VPWR
rlabel comment 1051 -8172 1051 -8172 4 sky130_fd_sc_hd__clkinv_1_3/clkinv_1
rlabel metal1 1051 -8220 1327 -8124 1 sky130_fd_sc_hd__clkinv_1_3/VGND
rlabel metal1 1051 -7676 1327 -7580 1 sky130_fd_sc_hd__clkinv_1_3/VPWR
flabel metal1 1448 -8189 1482 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_244/VGND
flabel metal1 1448 -7645 1482 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_244/VPWR
flabel nwell 1448 -7645 1482 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_244/VPB
flabel pwell 1448 -8189 1482 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_244/VNB
rlabel comment 1419 -8172 1419 -8172 4 sky130_fd_sc_hd__decap_4_244/decap_4
rlabel metal1 1419 -8220 1787 -8124 1 sky130_fd_sc_hd__decap_4_244/VGND
rlabel metal1 1419 -7676 1787 -7580 1 sky130_fd_sc_hd__decap_4_244/VPWR
flabel metal1 1908 -8189 1942 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_245/VGND
flabel metal1 1908 -7645 1942 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_245/VPWR
flabel nwell 1908 -7645 1942 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_245/VPB
flabel pwell 1908 -8189 1942 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_245/VNB
rlabel comment 1879 -8172 1879 -8172 4 sky130_fd_sc_hd__decap_4_245/decap_4
rlabel metal1 1879 -8220 2247 -8124 1 sky130_fd_sc_hd__decap_4_245/VGND
rlabel metal1 1879 -7676 2247 -7580 1 sky130_fd_sc_hd__decap_4_245/VPWR
flabel metal1 1349 -7648 1402 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_490/VPWR
flabel metal1 1348 -8190 1399 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_490/VGND
rlabel comment 1327 -8172 1327 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_490/tapvpwrvgnd_1
rlabel metal1 1327 -8220 1419 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_490/VGND
rlabel metal1 1327 -7676 1419 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_490/VPWR
flabel metal1 981 -7648 1034 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_491/VPWR
flabel metal1 980 -8190 1031 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_491/VGND
rlabel comment 959 -8172 959 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_491/tapvpwrvgnd_1
rlabel metal1 959 -8220 1051 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_491/VGND
rlabel metal1 959 -7676 1051 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_491/VPWR
flabel metal1 2269 -7648 2322 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_492/VPWR
flabel metal1 2268 -8190 2319 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_492/VGND
rlabel comment 2247 -8172 2247 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_492/tapvpwrvgnd_1
rlabel metal1 2247 -8220 2339 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_492/VGND
rlabel metal1 2247 -7676 2339 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_492/VPWR
flabel metal1 1809 -7648 1862 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_493/VPWR
flabel metal1 1808 -8190 1859 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_493/VGND
rlabel comment 1787 -8172 1787 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_493/tapvpwrvgnd_1
rlabel metal1 1787 -8220 1879 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_493/VGND
rlabel metal1 1787 -7676 1879 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_493/VPWR
flabel metal1 3196 -8189 3230 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_246/VGND
flabel metal1 3196 -7645 3230 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_246/VPWR
flabel nwell 3196 -7645 3230 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_246/VPB
flabel pwell 3196 -8189 3230 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_246/VNB
rlabel comment 3167 -8172 3167 -8172 4 sky130_fd_sc_hd__decap_4_246/decap_4
rlabel metal1 3167 -8220 3535 -8124 1 sky130_fd_sc_hd__decap_4_246/VGND
rlabel metal1 3167 -7676 3535 -7580 1 sky130_fd_sc_hd__decap_4_246/VPWR
flabel metal1 4392 -8189 4426 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_33/VGND
flabel metal1 4392 -7645 4426 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_33/VPWR
flabel nwell 4392 -7645 4426 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_33/VPB
flabel pwell 4392 -8189 4426 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_33/VNB
rlabel comment 4363 -8172 4363 -8172 4 sky130_fd_sc_hd__decap_12_33/decap_12
rlabel metal1 4363 -8220 5467 -8124 1 sky130_fd_sc_hd__decap_12_33/VGND
rlabel metal1 4363 -7676 5467 -7580 1 sky130_fd_sc_hd__decap_12_33/VPWR
flabel metal1 3662 -8192 3694 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_33/VGND
flabel metal1 3656 -7649 3694 -7617 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_33/VPWR
flabel nwell 3647 -7650 3704 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_33/VPB
flabel pwell 3653 -8196 3697 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_33/VNB
rlabel comment 3627 -8172 3627 -8172 4 sky130_fd_sc_hd__fill_8_33/fill_8
rlabel metal1 3627 -8220 4363 -8124 1 sky130_fd_sc_hd__fill_8_33/VGND
rlabel metal1 3627 -7676 4363 -7580 1 sky130_fd_sc_hd__fill_8_33/VPWR
flabel metal1 3097 -7648 3150 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_494/VPWR
flabel metal1 3096 -8190 3147 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_494/VGND
rlabel comment 3075 -8172 3075 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_494/tapvpwrvgnd_1
rlabel metal1 3075 -8220 3167 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_494/VGND
rlabel metal1 3075 -7676 3167 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_494/VPWR
flabel metal1 3557 -7648 3610 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_495/VPWR
flabel metal1 3556 -8190 3607 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_495/VGND
rlabel comment 3535 -8172 3535 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_495/tapvpwrvgnd_1
rlabel metal1 3535 -8220 3627 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_495/VGND
rlabel metal1 3535 -7676 3627 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_495/VPWR
flabel metal1 6416 -8189 6450 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_247/VGND
flabel metal1 6416 -7645 6450 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_247/VPWR
flabel nwell 6416 -7645 6450 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_247/VPB
flabel pwell 6416 -8189 6450 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_247/VNB
rlabel comment 6387 -8172 6387 -8172 4 sky130_fd_sc_hd__decap_4_247/decap_4
rlabel metal1 6387 -8220 6755 -8124 1 sky130_fd_sc_hd__decap_4_247/VGND
rlabel metal1 6387 -7676 6755 -7580 1 sky130_fd_sc_hd__decap_4_247/VPWR
flabel metal1 5857 -7645 5893 -7615 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_71/VPWR
flabel metal1 5857 -8185 5893 -8156 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_71/VGND
flabel nwell 5866 -7638 5886 -7621 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_71/VPB
flabel pwell 5863 -8183 5887 -8161 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_71/VNB
rlabel comment 5835 -8172 5835 -8172 4 sky130_fd_sc_hd__fill_1_71/fill_1
rlabel metal1 5835 -8220 5927 -8124 1 sky130_fd_sc_hd__fill_1_71/VGND
rlabel metal1 5835 -7676 5927 -7580 1 sky130_fd_sc_hd__fill_1_71/VPWR
flabel metal1 5961 -8182 5984 -8163 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_14/VGND
flabel metal1 5961 -7637 5981 -7620 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_14/VPWR
flabel nwell 5962 -7642 5987 -7616 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_14/VPB
flabel pwell 5962 -8184 5984 -8160 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_14/VNB
rlabel comment 5927 -8172 5927 -8172 4 sky130_fd_sc_hd__fill_4_14/fill_4
rlabel metal1 5927 -8220 6295 -8124 1 sky130_fd_sc_hd__fill_4_14/VGND
rlabel metal1 5927 -7676 6295 -7580 1 sky130_fd_sc_hd__fill_4_14/VPWR
flabel metal1 5501 -8182 5524 -8163 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_15/VGND
flabel metal1 5501 -7637 5521 -7620 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_15/VPWR
flabel nwell 5502 -7642 5527 -7616 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_15/VPB
flabel pwell 5502 -8184 5524 -8160 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_15/VNB
rlabel comment 5467 -8172 5467 -8172 4 sky130_fd_sc_hd__fill_4_15/fill_4
rlabel metal1 5467 -8220 5835 -8124 1 sky130_fd_sc_hd__fill_4_15/VGND
rlabel metal1 5467 -7676 5835 -7580 1 sky130_fd_sc_hd__fill_4_15/VPWR
flabel metal1 6317 -7648 6370 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_496/VPWR
flabel metal1 6316 -8190 6367 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_496/VGND
rlabel comment 6295 -8172 6295 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_496/tapvpwrvgnd_1
rlabel metal1 6295 -8220 6387 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_496/VGND
rlabel metal1 6295 -7676 6387 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_496/VPWR
flabel locali 6877 -7951 6911 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
flabel locali 7523 -7747 7557 -7713 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/X
flabel locali 7523 -7815 7557 -7781 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/X
flabel locali 7523 -7883 7557 -7849 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/X
flabel locali 7523 -7951 7557 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/X
flabel locali 7523 -8019 7557 -7985 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/X
flabel locali 7523 -8087 7557 -8053 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/X
flabel pwell 6877 -8189 6911 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/VNB
flabel nwell 6877 -7645 6911 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/VPB
flabel metal1 6877 -8189 6911 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/VGND
flabel metal1 6877 -7645 6911 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_197/VPWR
rlabel comment 6847 -8172 6847 -8172 4 sky130_fd_sc_hd__clkdlybuf4s50_1_197/clkdlybuf4s50_1
rlabel metal1 6847 -8220 7583 -8124 1 sky130_fd_sc_hd__clkdlybuf4s50_1_197/VGND
rlabel metal1 6847 -7676 7583 -7580 1 sky130_fd_sc_hd__clkdlybuf4s50_1_197/VPWR
flabel locali 8165 -7951 8199 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A
flabel locali 8811 -7747 8845 -7713 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/X
flabel locali 8811 -7815 8845 -7781 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/X
flabel locali 8811 -7883 8845 -7849 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/X
flabel locali 8811 -7951 8845 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/X
flabel locali 8811 -8019 8845 -7985 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/X
flabel locali 8811 -8087 8845 -8053 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/X
flabel pwell 8165 -8189 8199 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/VNB
flabel nwell 8165 -7645 8199 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/VPB
flabel metal1 8165 -8189 8199 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/VGND
flabel metal1 8165 -7645 8199 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_198/VPWR
rlabel comment 8135 -8172 8135 -8172 4 sky130_fd_sc_hd__clkdlybuf4s50_1_198/clkdlybuf4s50_1
rlabel metal1 8135 -8220 8871 -8124 1 sky130_fd_sc_hd__clkdlybuf4s50_1_198/VGND
rlabel metal1 8135 -7676 8871 -7580 1 sky130_fd_sc_hd__clkdlybuf4s50_1_198/VPWR
flabel metal1 7704 -8189 7738 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_248/VGND
flabel metal1 7704 -7645 7738 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_248/VPWR
flabel nwell 7704 -7645 7738 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_248/VPB
flabel pwell 7704 -8189 7738 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_248/VNB
rlabel comment 7675 -8172 7675 -8172 4 sky130_fd_sc_hd__decap_4_248/decap_4
rlabel metal1 7675 -8220 8043 -8124 1 sky130_fd_sc_hd__decap_4_248/VGND
rlabel metal1 7675 -7676 8043 -7580 1 sky130_fd_sc_hd__decap_4_248/VPWR
flabel metal1 6777 -7648 6830 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_497/VPWR
flabel metal1 6776 -8190 6827 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_497/VGND
rlabel comment 6755 -8172 6755 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_497/tapvpwrvgnd_1
rlabel metal1 6755 -8220 6847 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_497/VGND
rlabel metal1 6755 -7676 6847 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_497/VPWR
flabel metal1 8065 -7648 8118 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_498/VPWR
flabel metal1 8064 -8190 8115 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_498/VGND
rlabel comment 8043 -8172 8043 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_498/tapvpwrvgnd_1
rlabel metal1 8043 -8220 8135 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_498/VGND
rlabel metal1 8043 -7676 8135 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_498/VPWR
flabel metal1 7605 -7648 7658 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_499/VPWR
flabel metal1 7604 -8190 7655 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_499/VGND
rlabel comment 7583 -8172 7583 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_499/tapvpwrvgnd_1
rlabel metal1 7583 -8220 7675 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_499/VGND
rlabel metal1 7583 -7676 7675 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_499/VPWR
flabel locali 9453 -7951 9487 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A
flabel locali 10099 -7747 10133 -7713 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/X
flabel locali 10099 -7815 10133 -7781 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/X
flabel locali 10099 -7883 10133 -7849 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/X
flabel locali 10099 -7951 10133 -7917 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/X
flabel locali 10099 -8019 10133 -7985 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/X
flabel locali 10099 -8087 10133 -8053 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/X
flabel pwell 9453 -8189 9487 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/VNB
flabel nwell 9453 -7645 9487 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/VPB
flabel metal1 9453 -8189 9487 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/VGND
flabel metal1 9453 -7645 9487 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_199/VPWR
rlabel comment 9423 -8172 9423 -8172 4 sky130_fd_sc_hd__clkdlybuf4s50_1_199/clkdlybuf4s50_1
rlabel metal1 9423 -8220 10159 -8124 1 sky130_fd_sc_hd__clkdlybuf4s50_1_199/VGND
rlabel metal1 9423 -7676 10159 -7580 1 sky130_fd_sc_hd__clkdlybuf4s50_1_199/VPWR
flabel metal1 8992 -8189 9026 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_249/VGND
flabel metal1 8992 -7645 9026 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_249/VPWR
flabel nwell 8992 -7645 9026 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_249/VPB
flabel pwell 8992 -8189 9026 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_249/VNB
rlabel comment 8963 -8172 8963 -8172 4 sky130_fd_sc_hd__decap_4_249/decap_4
rlabel metal1 8963 -8220 9331 -8124 1 sky130_fd_sc_hd__decap_4_249/VGND
rlabel metal1 8963 -7676 9331 -7580 1 sky130_fd_sc_hd__decap_4_249/VPWR
flabel metal1 10280 -8189 10314 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_250/VGND
flabel metal1 10280 -7645 10314 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_250/VPWR
flabel nwell 10280 -7645 10314 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_250/VPB
flabel pwell 10280 -8189 10314 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_250/VNB
rlabel comment 10251 -8172 10251 -8172 4 sky130_fd_sc_hd__decap_4_250/decap_4
rlabel metal1 10251 -8220 10619 -8124 1 sky130_fd_sc_hd__decap_4_250/VGND
rlabel metal1 10251 -7676 10619 -7580 1 sky130_fd_sc_hd__decap_4_250/VPWR
flabel metal1 8893 -7648 8946 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_500/VPWR
flabel metal1 8892 -8190 8943 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_500/VGND
rlabel comment 8871 -8172 8871 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_500/tapvpwrvgnd_1
rlabel metal1 8871 -8220 8963 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_500/VGND
rlabel metal1 8871 -7676 8963 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_500/VPWR
flabel metal1 9353 -7648 9406 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_501/VPWR
flabel metal1 9352 -8190 9403 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_501/VGND
rlabel comment 9331 -8172 9331 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_501/tapvpwrvgnd_1
rlabel metal1 9331 -8220 9423 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_501/VGND
rlabel metal1 9331 -7676 9423 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_501/VPWR
flabel metal1 10181 -7648 10234 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_502/VPWR
flabel metal1 10180 -8190 10231 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_502/VGND
rlabel comment 10159 -8172 10159 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_502/tapvpwrvgnd_1
rlabel metal1 10159 -8220 10251 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_502/VGND
rlabel metal1 10159 -7676 10251 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_502/VPWR
flabel metal1 11660 -8189 11694 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_251/VGND
flabel metal1 11660 -7645 11694 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_251/VPWR
flabel nwell 11660 -7645 11694 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_251/VPB
flabel pwell 11660 -8189 11694 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_251/VNB
rlabel comment 11631 -8172 11631 -8172 4 sky130_fd_sc_hd__decap_4_251/decap_4
rlabel metal1 11631 -8220 11999 -8124 1 sky130_fd_sc_hd__decap_4_251/VGND
rlabel metal1 11631 -7676 11999 -7580 1 sky130_fd_sc_hd__decap_4_251/VPWR
flabel metal1 12034 -8192 12066 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_34/VGND
flabel metal1 12028 -7649 12066 -7617 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_34/VPWR
flabel nwell 12019 -7650 12076 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_34/VPB
flabel pwell 12025 -8196 12069 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_34/VNB
rlabel comment 11999 -8172 11999 -8172 4 sky130_fd_sc_hd__fill_8_34/fill_8
rlabel metal1 11999 -8220 12735 -8124 1 sky130_fd_sc_hd__fill_8_34/VGND
rlabel metal1 11999 -7676 12735 -7580 1 sky130_fd_sc_hd__fill_8_34/VPWR
flabel locali 11109 -7951 11143 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/Y
flabel locali 11109 -7883 11143 -7849 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/Y
flabel locali 11385 -7951 11419 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/A
flabel locali 11293 -7951 11327 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/A
flabel locali 11017 -7951 11051 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/B
flabel locali 10925 -7951 10959 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/B
flabel locali 10741 -7951 10775 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/B
flabel locali 10833 -7951 10867 -7917 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_3/B
flabel nwell 10741 -7645 10775 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_3/VPB
flabel pwell 10741 -8189 10775 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_3/VNB
flabel metal1 10741 -8189 10775 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_3/VGND
flabel metal1 10741 -7645 10775 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_3/VPWR
rlabel comment 10711 -8172 10711 -8172 4 sky130_fd_sc_hd__nand2_4_3/nand2_4
rlabel metal1 10711 -8220 11539 -8124 1 sky130_fd_sc_hd__nand2_4_3/VGND
rlabel metal1 10711 -7676 11539 -7580 1 sky130_fd_sc_hd__nand2_4_3/VPWR
flabel metal1 11561 -7648 11614 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_503/VPWR
flabel metal1 11560 -8190 11611 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_503/VGND
rlabel comment 11539 -8172 11539 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_503/tapvpwrvgnd_1
rlabel metal1 11539 -8220 11631 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_503/VGND
rlabel metal1 11539 -7676 11631 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_503/VPWR
flabel metal1 10641 -7648 10694 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_504/VPWR
flabel metal1 10640 -8190 10691 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_504/VGND
rlabel comment 10619 -8172 10619 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_504/tapvpwrvgnd_1
rlabel metal1 10619 -8220 10711 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_504/VGND
rlabel metal1 10619 -7676 10711 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_504/VPWR
flabel metal1 13592 -8189 13626 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_34/VGND
flabel metal1 13592 -7645 13626 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_34/VPWR
flabel nwell 13592 -7645 13626 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_34/VPB
flabel pwell 13592 -8189 13626 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_34/VNB
rlabel comment 13563 -8172 13563 -8172 4 sky130_fd_sc_hd__decap_12_34/decap_12
rlabel metal1 13563 -8220 14667 -8124 1 sky130_fd_sc_hd__decap_12_34/VGND
rlabel metal1 13563 -7676 14667 -7580 1 sky130_fd_sc_hd__decap_12_34/VPWR
flabel metal1 12770 -8192 12802 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_35/VGND
flabel metal1 12764 -7649 12802 -7617 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_35/VPWR
flabel nwell 12755 -7650 12812 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_35/VPB
flabel pwell 12761 -8196 12805 -8162 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_35/VNB
rlabel comment 12735 -8172 12735 -8172 4 sky130_fd_sc_hd__fill_8_35/fill_8
rlabel metal1 12735 -8220 13471 -8124 1 sky130_fd_sc_hd__fill_8_35/VGND
rlabel metal1 12735 -7676 13471 -7580 1 sky130_fd_sc_hd__fill_8_35/VPWR
flabel metal1 13493 -7648 13546 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_505/VPWR
flabel metal1 13492 -8190 13543 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_505/VGND
rlabel comment 13471 -8172 13471 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_505/tapvpwrvgnd_1
rlabel metal1 13471 -8220 13563 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_505/VGND
rlabel metal1 13471 -7676 13563 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_505/VPWR
flabel metal1 15984 -7645 16018 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_43/VPWR
flabel metal1 15984 -8189 16018 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_43/VGND
flabel nwell 15984 -7645 16018 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_43/VPB
flabel pwell 15984 -8189 16018 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_43/VNB
rlabel comment 15955 -8172 15955 -8172 4 sky130_fd_sc_hd__decap_8_43/decap_8
rlabel metal1 15955 -8220 16691 -8124 1 sky130_fd_sc_hd__decap_8_43/VGND
rlabel metal1 15955 -7676 16691 -7580 1 sky130_fd_sc_hd__decap_8_43/VPWR
flabel metal1 14788 -8189 14822 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_35/VGND
flabel metal1 14788 -7645 14822 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_35/VPWR
flabel nwell 14788 -7645 14822 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_35/VPB
flabel pwell 14788 -8189 14822 -8155 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_35/VNB
rlabel comment 14759 -8172 14759 -8172 4 sky130_fd_sc_hd__decap_12_35/decap_12
rlabel metal1 14759 -8220 15863 -8124 1 sky130_fd_sc_hd__decap_12_35/VGND
rlabel metal1 14759 -7676 15863 -7580 1 sky130_fd_sc_hd__decap_12_35/VPWR
flabel metal1 14689 -7648 14742 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_506/VPWR
flabel metal1 14688 -8190 14739 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_506/VGND
rlabel comment 14667 -8172 14667 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_506/tapvpwrvgnd_1
rlabel metal1 14667 -8220 14759 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_506/VGND
rlabel metal1 14667 -7676 14759 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_506/VPWR
flabel metal1 15885 -7648 15938 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_507/VPWR
flabel metal1 15884 -8190 15935 -8152 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_507/VGND
rlabel comment 15863 -8172 15863 -8172 4 sky130_fd_sc_hd__tapvpwrvgnd_1_507/tapvpwrvgnd_1
rlabel metal1 15863 -8220 15955 -8124 1 sky130_fd_sc_hd__tapvpwrvgnd_1_507/VGND
rlabel metal1 15863 -7676 15955 -7580 1 sky130_fd_sc_hd__tapvpwrvgnd_1_507/VPWR
flabel metal1 -1588 -7645 -1554 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_44/VPWR
flabel metal1 -1588 -7101 -1554 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_44/VGND
flabel nwell -1588 -7645 -1554 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_44/VPB
flabel pwell -1588 -7101 -1554 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_44/VNB
rlabel comment -1617 -7084 -1617 -7084 2 sky130_fd_sc_hd__decap_8_44/decap_8
rlabel metal1 -1617 -7132 -881 -7036 5 sky130_fd_sc_hd__decap_8_44/VGND
rlabel metal1 -1617 -7676 -881 -7580 5 sky130_fd_sc_hd__decap_8_44/VPWR
flabel metal1 -2324 -7645 -2290 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_78/VPWR
flabel metal1 -2324 -7101 -2290 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_78/VGND
flabel nwell -2324 -7645 -2290 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_78/VPB
flabel pwell -2324 -7101 -2290 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_78/VNB
rlabel comment -2261 -7084 -2261 -7084 8 sky130_fd_sc_hd__decap_8_78/decap_8
rlabel metal1 -2997 -7132 -2261 -7036 5 sky130_fd_sc_hd__decap_8_78/VGND
rlabel metal1 -2997 -7676 -2261 -7580 5 sky130_fd_sc_hd__decap_8_78/VPWR
flabel metal1 -1690 -7102 -1637 -7070 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_17/VGND
flabel metal1 -1690 -7645 -1638 -7614 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_17/VPWR
flabel nwell -1679 -7637 -1645 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_17/VPB
flabel pwell -1680 -7096 -1648 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_17/VNB
rlabel comment -1617 -7084 -1617 -7084 8 sky130_fd_sc_hd__fill_2_17/fill_2
rlabel metal1 -1801 -7132 -1617 -7036 5 sky130_fd_sc_hd__fill_2_17/VGND
rlabel metal1 -1801 -7676 -1617 -7580 5 sky130_fd_sc_hd__fill_2_17/VPWR
flabel metal1 -1858 -7093 -1835 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_17/VGND
flabel metal1 -1855 -7636 -1835 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_17/VPWR
flabel nwell -1861 -7640 -1836 -7614 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_17/VPB
flabel pwell -1858 -7096 -1836 -7072 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_17/VNB
rlabel comment -1801 -7084 -1801 -7084 8 sky130_fd_sc_hd__fill_4_17/fill_4
rlabel metal1 -2169 -7132 -1801 -7036 5 sky130_fd_sc_hd__fill_4_17/VGND
rlabel metal1 -2169 -7676 -1801 -7580 5 sky130_fd_sc_hd__fill_4_17/VPWR
flabel metal1 -2244 -7637 -2191 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_543/VPWR
flabel metal1 -2241 -7104 -2190 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_543/VGND
rlabel comment -2169 -7084 -2169 -7084 8 sky130_fd_sc_hd__tapvpwrvgnd_1_543/tapvpwrvgnd_1
rlabel metal1 -2261 -7132 -2169 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_543/VGND
rlabel metal1 -2261 -7676 -2169 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_543/VPWR
flabel metal1 -852 -7645 -818 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_45/VPWR
flabel metal1 -852 -7101 -818 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_45/VGND
flabel nwell -852 -7645 -818 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_45/VPB
flabel pwell -852 -7101 -818 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_45/VNB
rlabel comment -881 -7084 -881 -7084 2 sky130_fd_sc_hd__decap_8_45/decap_8
rlabel metal1 -881 -7132 -145 -7036 5 sky130_fd_sc_hd__decap_8_45/VGND
rlabel metal1 -881 -7676 -145 -7580 5 sky130_fd_sc_hd__decap_8_45/VPWR
flabel metal1 -24 -7645 10 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_48/VPWR
flabel metal1 -24 -7101 10 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_48/VGND
flabel nwell -24 -7645 10 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_48/VPB
flabel pwell -24 -7101 10 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_48/VNB
rlabel comment -53 -7084 -53 -7084 2 sky130_fd_sc_hd__decap_8_48/decap_8
rlabel metal1 -53 -7132 683 -7036 5 sky130_fd_sc_hd__decap_8_48/VGND
rlabel metal1 -53 -7676 683 -7580 5 sky130_fd_sc_hd__decap_8_48/VPWR
flabel metal1 712 -7645 746 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_49/VPWR
flabel metal1 712 -7101 746 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_49/VGND
flabel nwell 712 -7645 746 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_49/VPB
flabel pwell 712 -7101 746 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_49/VNB
rlabel comment 683 -7084 683 -7084 2 sky130_fd_sc_hd__decap_8_49/decap_8
rlabel metal1 683 -7132 1419 -7036 5 sky130_fd_sc_hd__decap_8_49/VGND
rlabel metal1 683 -7676 1419 -7580 5 sky130_fd_sc_hd__decap_8_49/VPWR
flabel metal1 -123 -7637 -70 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_514/VPWR
flabel metal1 -124 -7104 -73 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_514/VGND
rlabel comment -145 -7084 -145 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_514/tapvpwrvgnd_1
rlabel metal1 -145 -7132 -53 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_514/VGND
rlabel metal1 -145 -7676 -53 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_514/VPWR
flabel metal1 2552 -7101 2586 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_255/VGND
flabel metal1 2552 -7645 2586 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_255/VPWR
flabel nwell 2552 -7645 2586 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_255/VPB
flabel pwell 2552 -7101 2586 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_255/VNB
rlabel comment 2615 -7084 2615 -7084 8 sky130_fd_sc_hd__decap_4_255/decap_4
rlabel metal1 2247 -7132 2615 -7036 5 sky130_fd_sc_hd__decap_4_255/VGND
rlabel metal1 2247 -7676 2615 -7580 5 sky130_fd_sc_hd__decap_4_255/VPWR
flabel metal1 1540 -7645 1574 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_53/VPWR
flabel metal1 1540 -7101 1574 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_53/VGND
flabel nwell 1540 -7645 1574 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_53/VPB
flabel pwell 1540 -7101 1574 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_53/VNB
rlabel comment 1511 -7084 1511 -7084 2 sky130_fd_sc_hd__decap_8_53/decap_8
rlabel metal1 1511 -7132 2247 -7036 5 sky130_fd_sc_hd__decap_8_53/VGND
rlabel metal1 1511 -7676 2247 -7580 5 sky130_fd_sc_hd__decap_8_53/VPWR
flabel metal1 2726 -7102 2779 -7070 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_4/VGND
flabel metal1 2726 -7645 2778 -7614 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_4/VPWR
flabel nwell 2737 -7637 2771 -7619 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_4/VPB
flabel pwell 2736 -7096 2768 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_4/VNB
rlabel comment 2799 -7084 2799 -7084 8 sky130_fd_sc_hd__fill_2_4/fill_2
rlabel metal1 2615 -7132 2799 -7036 5 sky130_fd_sc_hd__fill_2_4/VGND
rlabel metal1 2615 -7676 2799 -7580 5 sky130_fd_sc_hd__fill_2_4/VPWR
flabel metal1 1441 -7637 1494 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_516/VPWR
flabel metal1 1440 -7104 1491 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_516/VGND
rlabel comment 1419 -7084 1419 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_516/tapvpwrvgnd_1
rlabel metal1 1419 -7132 1511 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_516/VGND
rlabel metal1 1419 -7676 1511 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_516/VPWR
flabel metal1 2816 -7637 2869 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_519/VPWR
flabel metal1 2819 -7104 2870 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_519/VGND
rlabel comment 2891 -7084 2891 -7084 8 sky130_fd_sc_hd__tapvpwrvgnd_1_519/tapvpwrvgnd_1
rlabel metal1 2799 -7132 2891 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_519/VGND
rlabel metal1 2799 -7676 2891 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_519/VPWR
flabel metal1 3649 -7637 3702 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_509/VPWR
flabel metal1 3648 -7104 3699 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_509/VGND
rlabel comment 3627 -7084 3627 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_509/tapvpwrvgnd_1
rlabel metal1 3627 -7132 3719 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_509/VGND
rlabel metal1 3627 -7676 3719 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_509/VPWR
flabel metal1 3189 -7637 3242 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_508/VPWR
flabel metal1 3188 -7104 3239 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_508/VGND
rlabel comment 3167 -7084 3167 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_508/tapvpwrvgnd_1
rlabel metal1 3167 -7132 3259 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_508/VGND
rlabel metal1 3167 -7676 3259 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_508/VPWR
flabel metal1 3564 -7101 3598 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_252/VGND
flabel metal1 3564 -7645 3598 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_252/VPWR
flabel nwell 3564 -7645 3598 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_252/VPB
flabel pwell 3564 -7101 3598 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_252/VNB
rlabel comment 3627 -7084 3627 -7084 8 sky130_fd_sc_hd__decap_4_252/decap_4
rlabel metal1 3259 -7132 3627 -7036 5 sky130_fd_sc_hd__decap_4_252/VGND
rlabel metal1 3259 -7676 3627 -7580 5 sky130_fd_sc_hd__decap_4_252/VPWR
flabel locali 2920 -7271 2954 -7237 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/Y
flabel locali 2920 -7339 2954 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/Y
flabel locali 3012 -7407 3046 -7373 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/Y
flabel locali 3012 -7339 3046 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/Y
flabel locali 3012 -7271 3046 -7237 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/Y
flabel locali 3104 -7203 3138 -7169 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/A
flabel locali 3104 -7271 3138 -7237 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/A
flabel locali 3104 -7339 3138 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_4/A
flabel nwell 3104 -7645 3138 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_4/VPB
flabel pwell 3104 -7101 3138 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_4/VNB
flabel metal1 3104 -7101 3138 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_4/VGND
flabel metal1 3104 -7645 3138 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_4/VPWR
rlabel comment 3167 -7084 3167 -7084 8 sky130_fd_sc_hd__clkinv_1_4/clkinv_1
rlabel metal1 2891 -7132 3167 -7036 5 sky130_fd_sc_hd__clkinv_1_4/VGND
rlabel metal1 2891 -7676 3167 -7580 5 sky130_fd_sc_hd__clkinv_1_4/VPWR
flabel metal1 4477 -7637 4530 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_511/VPWR
flabel metal1 4476 -7104 4527 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_511/VGND
rlabel comment 4455 -7084 4455 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_511/tapvpwrvgnd_1
rlabel metal1 4455 -7132 4547 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_511/VGND
rlabel metal1 4455 -7676 4547 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_511/VPWR
flabel metal1 4017 -7637 4070 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_510/VPWR
flabel metal1 4016 -7104 4067 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_510/VGND
rlabel comment 3995 -7084 3995 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_510/tapvpwrvgnd_1
rlabel metal1 3995 -7132 4087 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_510/VGND
rlabel metal1 3995 -7676 4087 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_510/VPWR
flabel locali 3839 -7203 3873 -7169 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_4/Y
flabel locali 3839 -7271 3873 -7237 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_4/Y
flabel locali 3839 -7339 3873 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_4/Y
flabel locali 3747 -7339 3781 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_4/B
flabel locali 3931 -7339 3965 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_4/A
flabel nwell 3747 -7645 3781 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_4/VPB
flabel pwell 3747 -7101 3781 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_4/VNB
flabel metal1 3747 -7101 3781 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_4/VGND
flabel metal1 3747 -7645 3781 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_4/VPWR
rlabel comment 3719 -7084 3719 -7084 2 sky130_fd_sc_hd__nand2_1_4/nand2_1
rlabel metal1 3719 -7132 3995 -7036 5 sky130_fd_sc_hd__nand2_1_4/VGND
rlabel metal1 3719 -7676 3995 -7580 5 sky130_fd_sc_hd__nand2_1_4/VPWR
flabel metal1 4577 -7101 4611 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__mux2_1_0/VGND
flabel metal1 4577 -7645 4611 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__mux2_1_0/VPWR
flabel locali 5221 -7407 5255 -7373 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/S
flabel locali 5129 -7407 5163 -7373 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/S
flabel locali 5037 -7271 5071 -7237 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/A1
flabel locali 5037 -7339 5071 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/A1
flabel locali 4945 -7339 4979 -7305 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/A0
flabel locali 4577 -7203 4611 -7169 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/X
flabel locali 4577 -7475 4611 -7441 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/X
flabel locali 4577 -7543 4611 -7509 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/X
flabel nwell 4621 -7645 4655 -7611 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/VPB
flabel pwell 4631 -7101 4665 -7067 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__mux2_1_0/VNB
rlabel comment 4547 -7084 4547 -7084 2 sky130_fd_sc_hd__mux2_1_0/mux2_1
rlabel metal1 4547 -7132 5375 -7036 5 sky130_fd_sc_hd__mux2_1_0/VGND
rlabel metal1 4547 -7676 5375 -7580 5 sky130_fd_sc_hd__mux2_1_0/VPWR
flabel metal1 4392 -7101 4426 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_253/VGND
flabel metal1 4392 -7645 4426 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_253/VPWR
flabel nwell 4392 -7645 4426 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_253/VPB
flabel pwell 4392 -7101 4426 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_253/VNB
rlabel comment 4455 -7084 4455 -7084 8 sky130_fd_sc_hd__decap_4_253/decap_4
rlabel metal1 4087 -7132 4455 -7036 5 sky130_fd_sc_hd__decap_4_253/VGND
rlabel metal1 4087 -7676 4455 -7580 5 sky130_fd_sc_hd__decap_4_253/VPWR
flabel metal1 5772 -7101 5806 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_254/VGND
flabel metal1 5772 -7645 5806 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_254/VPWR
flabel nwell 5772 -7645 5806 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_254/VPB
flabel pwell 5772 -7101 5806 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_254/VNB
rlabel comment 5835 -7084 5835 -7084 8 sky130_fd_sc_hd__decap_4_254/decap_4
rlabel metal1 5467 -7132 5835 -7036 5 sky130_fd_sc_hd__decap_4_254/VGND
rlabel metal1 5467 -7676 5835 -7580 5 sky130_fd_sc_hd__decap_4_254/VPWR
flabel metal1 7612 -7101 7646 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VGND
flabel metal1 7612 -7645 7646 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPWR
flabel locali 5956 -7422 5990 -7388 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q_N
flabel locali 7352 -7339 7386 -7305 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/D
flabel locali 7612 -7339 7646 -7305 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/CLK
flabel locali 6251 -7203 6285 -7169 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q
flabel pwell 7612 -7101 7646 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel pwell 7629 -7084 7629 -7084 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel nwell 7612 -7645 7646 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
flabel nwell 7629 -7628 7629 -7628 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
rlabel comment 7675 -7084 7675 -7084 8 sky130_fd_sc_hd__dfxbp_1_0/dfxbp_1
rlabel metal1 5927 -7132 7675 -7036 5 sky130_fd_sc_hd__dfxbp_1_0/VGND
rlabel metal1 5927 -7676 7675 -7580 5 sky130_fd_sc_hd__dfxbp_1_0/VPWR
flabel metal1 5397 -7637 5450 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_512/VPWR
flabel metal1 5396 -7104 5447 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_512/VGND
rlabel comment 5375 -7084 5375 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_512/tapvpwrvgnd_1
rlabel metal1 5375 -7132 5467 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_512/VGND
rlabel metal1 5375 -7676 5467 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_512/VPWR
flabel metal1 5857 -7637 5910 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_513/VPWR
flabel metal1 5856 -7104 5907 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_513/VGND
rlabel comment 5835 -7084 5835 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_513/tapvpwrvgnd_1
rlabel metal1 5835 -7132 5927 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_513/VGND
rlabel metal1 5835 -7676 5927 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_513/VPWR
flabel metal1 7796 -7645 7830 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_52/VPWR
flabel metal1 7796 -7101 7830 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_52/VGND
flabel nwell 7796 -7645 7830 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_52/VPB
flabel pwell 7796 -7101 7830 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_52/VNB
rlabel comment 7767 -7084 7767 -7084 2 sky130_fd_sc_hd__decap_8_52/decap_8
rlabel metal1 7767 -7132 8503 -7036 5 sky130_fd_sc_hd__decap_8_52/VGND
rlabel metal1 7767 -7676 8503 -7580 5 sky130_fd_sc_hd__decap_8_52/VPWR
flabel metal1 8532 -7645 8566 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_54/VPWR
flabel metal1 8532 -7101 8566 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_54/VGND
flabel nwell 8532 -7645 8566 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_54/VPB
flabel pwell 8532 -7101 8566 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_54/VNB
rlabel comment 8503 -7084 8503 -7084 2 sky130_fd_sc_hd__decap_8_54/decap_8
rlabel metal1 8503 -7132 9239 -7036 5 sky130_fd_sc_hd__decap_8_54/VGND
rlabel metal1 8503 -7676 9239 -7580 5 sky130_fd_sc_hd__decap_8_54/VPWR
flabel metal1 7697 -7637 7750 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_518/VPWR
flabel metal1 7696 -7104 7747 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_518/VGND
rlabel comment 7675 -7084 7675 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_518/tapvpwrvgnd_1
rlabel metal1 7675 -7132 7767 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_518/VGND
rlabel metal1 7675 -7676 7767 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_518/VPWR
flabel metal1 10000 -7094 10032 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_37/VGND
flabel metal1 10000 -7639 10038 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_37/VPWR
flabel nwell 9990 -7637 10047 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_37/VPB
flabel pwell 9997 -7094 10041 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_37/VNB
rlabel comment 10067 -7084 10067 -7084 8 sky130_fd_sc_hd__fill_8_37/fill_8
rlabel metal1 9331 -7132 10067 -7036 5 sky130_fd_sc_hd__fill_8_37/VGND
rlabel metal1 9331 -7676 10067 -7580 5 sky130_fd_sc_hd__fill_8_37/VPWR
flabel metal1 10736 -7094 10768 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_38/VGND
flabel metal1 10736 -7639 10774 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_38/VPWR
flabel nwell 10726 -7637 10783 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_38/VPB
flabel pwell 10733 -7094 10777 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_38/VNB
rlabel comment 10803 -7084 10803 -7084 8 sky130_fd_sc_hd__fill_8_38/fill_8
rlabel metal1 10067 -7132 10803 -7036 5 sky130_fd_sc_hd__fill_8_38/VGND
rlabel metal1 10067 -7676 10803 -7580 5 sky130_fd_sc_hd__fill_8_38/VPWR
flabel metal1 9261 -7637 9314 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_520/VPWR
flabel metal1 9260 -7104 9311 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_520/VGND
rlabel comment 9239 -7084 9239 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_520/tapvpwrvgnd_1
rlabel metal1 9239 -7132 9331 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_520/VGND
rlabel metal1 9239 -7676 9331 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_520/VPWR
flabel metal1 11472 -7094 11504 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_40/VGND
flabel metal1 11472 -7639 11510 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_40/VPWR
flabel nwell 11462 -7637 11519 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_40/VPB
flabel pwell 11469 -7094 11513 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_40/VNB
rlabel comment 11539 -7084 11539 -7084 8 sky130_fd_sc_hd__fill_8_40/fill_8
rlabel metal1 10803 -7132 11539 -7036 5 sky130_fd_sc_hd__fill_8_40/VGND
rlabel metal1 10803 -7676 11539 -7580 5 sky130_fd_sc_hd__fill_8_40/VPWR
flabel metal1 12208 -7094 12240 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_41/VGND
flabel metal1 12208 -7639 12246 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_41/VPWR
flabel nwell 12198 -7637 12255 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_41/VPB
flabel pwell 12205 -7094 12249 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_41/VNB
rlabel comment 12275 -7084 12275 -7084 8 sky130_fd_sc_hd__fill_8_41/fill_8
rlabel metal1 11539 -7132 12275 -7036 5 sky130_fd_sc_hd__fill_8_41/VGND
rlabel metal1 11539 -7676 12275 -7580 5 sky130_fd_sc_hd__fill_8_41/VPWR
flabel metal1 12944 -7094 12976 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_44/VGND
flabel metal1 12944 -7639 12982 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_44/VPWR
flabel nwell 12934 -7637 12991 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_44/VPB
flabel pwell 12941 -7094 12985 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_44/VNB
rlabel comment 13011 -7084 13011 -7084 8 sky130_fd_sc_hd__fill_8_44/fill_8
rlabel metal1 12275 -7132 13011 -7036 5 sky130_fd_sc_hd__fill_8_44/VGND
rlabel metal1 12275 -7676 13011 -7580 5 sky130_fd_sc_hd__fill_8_44/VPWR
flabel metal1 13680 -7094 13712 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_45/VGND
flabel metal1 13680 -7639 13718 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_45/VPWR
flabel nwell 13670 -7637 13727 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_45/VPB
flabel pwell 13677 -7094 13721 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_45/VNB
rlabel comment 13747 -7084 13747 -7084 8 sky130_fd_sc_hd__fill_8_45/fill_8
rlabel metal1 13011 -7132 13747 -7036 5 sky130_fd_sc_hd__fill_8_45/VGND
rlabel metal1 13011 -7676 13747 -7580 5 sky130_fd_sc_hd__fill_8_45/VPWR
flabel metal1 14416 -7094 14448 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_48/VGND
flabel metal1 14416 -7639 14454 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_48/VPWR
flabel nwell 14406 -7637 14463 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_48/VPB
flabel pwell 14413 -7094 14457 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_48/VNB
rlabel comment 14483 -7084 14483 -7084 8 sky130_fd_sc_hd__fill_8_48/fill_8
rlabel metal1 13747 -7132 14483 -7036 5 sky130_fd_sc_hd__fill_8_48/VGND
rlabel metal1 13747 -7676 14483 -7580 5 sky130_fd_sc_hd__fill_8_48/VPWR
flabel metal1 15984 -7645 16018 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_64/VPWR
flabel metal1 15984 -7101 16018 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_64/VGND
flabel nwell 15984 -7645 16018 -7611 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_64/VPB
flabel pwell 15984 -7101 16018 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_64/VNB
rlabel comment 15955 -7084 15955 -7084 2 sky130_fd_sc_hd__decap_8_64/decap_8
rlabel metal1 15955 -7132 16691 -7036 5 sky130_fd_sc_hd__decap_8_64/VGND
rlabel metal1 15955 -7676 16691 -7580 5 sky130_fd_sc_hd__decap_8_64/VPWR
flabel metal1 15152 -7094 15184 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_49/VGND
flabel metal1 15152 -7639 15190 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_49/VPWR
flabel nwell 15142 -7637 15199 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_49/VPB
flabel pwell 15149 -7094 15193 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_49/VNB
rlabel comment 15219 -7084 15219 -7084 8 sky130_fd_sc_hd__fill_8_49/fill_8
rlabel metal1 14483 -7132 15219 -7036 5 sky130_fd_sc_hd__fill_8_49/VGND
rlabel metal1 14483 -7676 15219 -7580 5 sky130_fd_sc_hd__fill_8_49/VPWR
flabel metal1 15888 -7094 15920 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_53/VGND
flabel metal1 15888 -7639 15926 -7607 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_53/VPWR
flabel nwell 15878 -7637 15935 -7606 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_53/VPB
flabel pwell 15885 -7094 15929 -7060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_53/VNB
rlabel comment 15955 -7084 15955 -7084 8 sky130_fd_sc_hd__fill_8_53/fill_8
rlabel metal1 15219 -7132 15955 -7036 5 sky130_fd_sc_hd__fill_8_53/VGND
rlabel metal1 15219 -7676 15955 -7580 5 sky130_fd_sc_hd__fill_8_53/VPWR
flabel metal1 15885 -7637 15938 -7608 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_524/VPWR
flabel metal1 15884 -7104 15935 -7066 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_524/VGND
rlabel comment 15863 -7084 15863 -7084 2 sky130_fd_sc_hd__tapvpwrvgnd_1_524/tapvpwrvgnd_1
rlabel metal1 15863 -7132 15955 -7036 5 sky130_fd_sc_hd__tapvpwrvgnd_1_524/VGND
rlabel metal1 15863 -7676 15955 -7580 5 sky130_fd_sc_hd__tapvpwrvgnd_1_524/VPWR
flabel metal1 -2968 -6557 -2934 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_3_0/VPWR
flabel metal1 -2968 -7101 -2934 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_3_0/VGND
flabel nwell -2968 -6557 -2934 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_3_0/VPB
flabel pwell -2968 -7101 -2934 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_3_0/VNB
rlabel comment -2997 -7084 -2997 -7084 4 sky130_fd_sc_hd__decap_3_0/decap_3
rlabel metal1 -2997 -7132 -2721 -7036 1 sky130_fd_sc_hd__decap_3_0/VGND
rlabel metal1 -2997 -6588 -2721 -6492 1 sky130_fd_sc_hd__decap_3_0/VPWR
flabel metal1 -1404 -6013 -1370 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_105/VGND
flabel metal1 -1404 -6557 -1370 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_105/VPWR
flabel nwell -1404 -6557 -1370 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_105/VPB
flabel pwell -1404 -6013 -1370 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_105/VNB
rlabel comment -1433 -5996 -1433 -5996 2 sky130_fd_sc_hd__decap_4_105/decap_4
rlabel metal1 -1433 -6044 -1065 -5948 5 sky130_fd_sc_hd__decap_4_105/VGND
rlabel metal1 -1433 -6588 -1065 -6492 5 sky130_fd_sc_hd__decap_4_105/VPWR
flabel metal1 -2324 -6557 -2290 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_76/VPWR
flabel metal1 -2324 -6013 -2290 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_76/VGND
flabel nwell -2324 -6557 -2290 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_76/VPB
flabel pwell -2324 -6013 -2290 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_76/VNB
rlabel comment -2261 -5996 -2261 -5996 8 sky130_fd_sc_hd__decap_8_76/decap_8
rlabel metal1 -2997 -6044 -2261 -5948 5 sky130_fd_sc_hd__decap_8_76/VGND
rlabel metal1 -2997 -6588 -2261 -6492 5 sky130_fd_sc_hd__decap_8_76/VPWR
flabel metal1 -2600 -7101 -2566 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VGND
flabel metal1 -2600 -6557 -2566 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPWR
flabel locali -944 -6780 -910 -6746 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/Q_N
flabel locali -2340 -6863 -2306 -6829 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/D
flabel locali -2600 -6863 -2566 -6829 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/CLK
flabel locali -1239 -6999 -1205 -6965 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/Q
flabel pwell -2600 -7101 -2566 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel pwell -2583 -7084 -2583 -7084 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel nwell -2600 -6557 -2566 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPB
flabel nwell -2583 -6540 -2583 -6540 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPB
rlabel comment -2629 -7084 -2629 -7084 4 sky130_fd_sc_hd__dfxbp_1_1/dfxbp_1
rlabel metal1 -2629 -7132 -881 -7036 1 sky130_fd_sc_hd__dfxbp_1_1/VGND
rlabel metal1 -2629 -6588 -881 -6492 1 sky130_fd_sc_hd__dfxbp_1_1/VPWR
flabel metal1 -1597 -6014 -1544 -5982 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VGND
flabel metal1 -1596 -6557 -1544 -6526 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VPWR
flabel nwell -1589 -6549 -1555 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VPB
flabel pwell -1586 -6008 -1554 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VNB
rlabel comment -1617 -5996 -1617 -5996 2 sky130_fd_sc_hd__fill_2_1/fill_2
rlabel metal1 -1617 -6044 -1433 -5948 5 sky130_fd_sc_hd__fill_2_1/VGND
rlabel metal1 -1617 -6588 -1433 -6492 5 sky130_fd_sc_hd__fill_2_1/VPWR
flabel metal1 -1690 -6014 -1637 -5982 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_13/VGND
flabel metal1 -1690 -6557 -1638 -6526 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_13/VPWR
flabel nwell -1679 -6549 -1645 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_13/VPB
flabel pwell -1680 -6008 -1648 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_13/VNB
rlabel comment -1617 -5996 -1617 -5996 8 sky130_fd_sc_hd__fill_2_13/fill_2
rlabel metal1 -1801 -6044 -1617 -5948 5 sky130_fd_sc_hd__fill_2_13/VGND
rlabel metal1 -1801 -6588 -1617 -6492 5 sky130_fd_sc_hd__fill_2_13/VPWR
flabel metal1 -1858 -6005 -1835 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_26/VGND
flabel metal1 -1855 -6548 -1835 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_26/VPWR
flabel nwell -1861 -6552 -1836 -6526 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_26/VPB
flabel pwell -1858 -6008 -1836 -5984 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_26/VNB
rlabel comment -1801 -5996 -1801 -5996 8 sky130_fd_sc_hd__fill_4_26/fill_4
rlabel metal1 -2169 -6044 -1801 -5948 5 sky130_fd_sc_hd__fill_4_26/VGND
rlabel metal1 -2169 -6588 -1801 -6492 5 sky130_fd_sc_hd__fill_4_26/VPWR
flabel metal1 -2704 -6560 -2651 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_523/VPWR
flabel metal1 -2701 -7102 -2650 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_523/VGND
rlabel comment -2629 -7084 -2629 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_523/tapvpwrvgnd_1
rlabel metal1 -2721 -7132 -2629 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_523/VGND
rlabel metal1 -2721 -6588 -2629 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_523/VPWR
flabel metal1 -2244 -6549 -2191 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_541/VPWR
flabel metal1 -2241 -6016 -2190 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_541/VGND
rlabel comment -2169 -5996 -2169 -5996 8 sky130_fd_sc_hd__tapvpwrvgnd_1_541/tapvpwrvgnd_1
rlabel metal1 -2261 -6044 -2169 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_541/VGND
rlabel metal1 -2261 -6588 -2169 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_541/VPWR
flabel metal1 -675 -6549 -622 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_213/VPWR
flabel metal1 -676 -6016 -625 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_213/VGND
rlabel comment -697 -5996 -697 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_213/tapvpwrvgnd_1
rlabel metal1 -697 -6044 -605 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_213/VGND
rlabel metal1 -697 -6588 -605 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_213/VPWR
flabel metal1 -1043 -6549 -990 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_212/VPWR
flabel metal1 -1044 -6016 -993 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_212/VGND
rlabel comment -1065 -5996 -1065 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_212/tapvpwrvgnd_1
rlabel metal1 -1065 -6044 -973 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_212/VGND
rlabel metal1 -1065 -6588 -973 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_212/VPWR
flabel locali -853 -6115 -819 -6081 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali -853 -6183 -819 -6149 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali -853 -6251 -819 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali -945 -6251 -911 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/B
flabel locali -761 -6251 -727 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/A
flabel nwell -945 -6557 -911 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VPB
flabel pwell -945 -6013 -911 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VNB
flabel metal1 -945 -6013 -911 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VGND
flabel metal1 -945 -6557 -911 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VPWR
rlabel comment -973 -5996 -973 -5996 2 sky130_fd_sc_hd__nand2_1_1/nand2_1
rlabel metal1 -973 -6044 -697 -5948 5 sky130_fd_sc_hd__nand2_1_1/VGND
rlabel metal1 -973 -6588 -697 -6492 5 sky130_fd_sc_hd__nand2_1_1/VPWR
flabel metal1 -208 -6557 -174 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_47/VPWR
flabel metal1 -208 -7101 -174 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_47/VGND
flabel nwell -208 -6557 -174 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_47/VPB
flabel pwell -208 -7101 -174 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_47/VNB
rlabel comment -145 -7084 -145 -7084 6 sky130_fd_sc_hd__decap_8_47/decap_8
rlabel metal1 -881 -7132 -145 -7036 1 sky130_fd_sc_hd__decap_8_47/VGND
rlabel metal1 -881 -6588 -145 -6492 1 sky130_fd_sc_hd__decap_8_47/VPWR
flabel metal1 -576 -6013 -542 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_106/VGND
flabel metal1 -576 -6557 -542 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_106/VPWR
flabel nwell -576 -6557 -542 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_106/VPB
flabel pwell -576 -6013 -542 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_106/VNB
rlabel comment -605 -5996 -605 -5996 2 sky130_fd_sc_hd__decap_4_106/decap_4
rlabel metal1 -605 -6044 -237 -5948 5 sky130_fd_sc_hd__decap_4_106/VGND
rlabel metal1 -605 -6588 -237 -6492 5 sky130_fd_sc_hd__decap_4_106/VPWR
flabel metal1 -128 -6560 -75 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_515/VPWR
flabel metal1 -125 -7102 -74 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_515/VGND
rlabel comment -53 -7084 -53 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_515/tapvpwrvgnd_1
rlabel metal1 -145 -7132 -53 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_515/VGND
rlabel metal1 -145 -6588 -53 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_515/VPWR
flabel metal1 521 -6549 574 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_217/VPWR
flabel metal1 520 -6016 571 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_217/VGND
rlabel comment 499 -5996 499 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_217/tapvpwrvgnd_1
rlabel metal1 499 -6044 591 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_217/VGND
rlabel metal1 499 -6588 591 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_217/VPWR
flabel metal1 -215 -6549 -162 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_216/VPWR
flabel metal1 -216 -6016 -165 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_216/VGND
rlabel comment -237 -5996 -237 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_216/tapvpwrvgnd_1
rlabel metal1 -237 -6044 -145 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_216/VGND
rlabel metal1 -237 -6588 -145 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_216/VPWR
flabel metal1 620 -6557 654 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_50/VPWR
flabel metal1 620 -7101 654 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_50/VGND
flabel nwell 620 -6557 654 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_50/VPB
flabel pwell 620 -7101 654 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_50/VNB
rlabel comment 683 -7084 683 -7084 6 sky130_fd_sc_hd__decap_8_50/decap_8
rlabel metal1 -53 -7132 683 -7036 1 sky130_fd_sc_hd__decap_8_50/VGND
rlabel metal1 -53 -6588 683 -6492 1 sky130_fd_sc_hd__decap_8_50/VPWR
flabel locali 68 -6251 102 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/A
flabel locali 160 -6251 194 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/A
flabel locali 436 -6183 470 -6149 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/Y
flabel locali -24 -6251 10 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/A
flabel locali 436 -6319 470 -6285 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/Y
flabel locali 344 -6251 378 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/A
flabel locali 252 -6251 286 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/A
flabel locali 436 -6251 470 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_5/Y
flabel pwell -116 -6013 -82 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_5/VNB
flabel nwell -116 -6557 -82 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_5/VPB
flabel metal1 -116 -6557 -82 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_5/VPWR
flabel metal1 -116 -6013 -82 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_5/VGND
rlabel comment -145 -5996 -145 -5996 2 sky130_fd_sc_hd__clkinv_4_5/clkinv_4
rlabel metal1 -145 -6044 499 -5948 5 sky130_fd_sc_hd__clkinv_4_5/VGND
rlabel metal1 -145 -6588 499 -6492 5 sky130_fd_sc_hd__clkinv_4_5/VPWR
flabel metal1 1356 -6557 1390 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_51/VPWR
flabel metal1 1356 -7101 1390 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_51/VGND
flabel nwell 1356 -6557 1390 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_51/VPB
flabel pwell 1356 -7101 1390 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_51/VNB
rlabel comment 1419 -7084 1419 -7084 6 sky130_fd_sc_hd__decap_8_51/decap_8
rlabel metal1 683 -7132 1419 -7036 1 sky130_fd_sc_hd__decap_8_51/VGND
rlabel metal1 683 -6588 1419 -6492 1 sky130_fd_sc_hd__decap_8_51/VPWR
flabel metal1 620 -6013 654 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_108/VGND
flabel metal1 620 -6557 654 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_108/VPWR
flabel nwell 620 -6557 654 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_108/VPB
flabel pwell 620 -6013 654 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_108/VNB
rlabel comment 591 -5996 591 -5996 2 sky130_fd_sc_hd__decap_4_108/decap_4
rlabel metal1 591 -6044 959 -5948 5 sky130_fd_sc_hd__decap_4_108/VGND
rlabel metal1 591 -6588 959 -6492 5 sky130_fd_sc_hd__decap_4_108/VPWR
flabel metal1 1436 -6560 1489 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_517/VPWR
flabel metal1 1439 -7102 1490 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_517/VGND
rlabel comment 1511 -7084 1511 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_517/tapvpwrvgnd_1
rlabel metal1 1419 -7132 1511 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_517/VGND
rlabel metal1 1419 -6588 1511 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_517/VPWR
flabel metal1 981 -6549 1034 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_219/VPWR
flabel metal1 980 -6016 1031 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_219/VGND
rlabel comment 959 -5996 959 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_219/tapvpwrvgnd_1
rlabel metal1 959 -6044 1051 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_219/VGND
rlabel metal1 959 -6588 1051 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_219/VPWR
flabel metal1 1349 -6549 1402 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_218/VPWR
flabel metal1 1348 -6016 1399 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_218/VGND
rlabel comment 1327 -5996 1327 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_218/tapvpwrvgnd_1
rlabel metal1 1327 -6044 1419 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_218/VGND
rlabel metal1 1327 -6588 1419 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_218/VPWR
flabel metal1 2184 -6557 2218 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_55/VPWR
flabel metal1 2184 -7101 2218 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_55/VGND
flabel nwell 2184 -6557 2218 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_55/VPB
flabel pwell 2184 -7101 2218 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_55/VNB
rlabel comment 2247 -7084 2247 -7084 6 sky130_fd_sc_hd__decap_8_55/decap_8
rlabel metal1 1511 -7132 2247 -7036 1 sky130_fd_sc_hd__decap_8_55/VGND
rlabel metal1 1511 -6588 2247 -6492 1 sky130_fd_sc_hd__decap_8_55/VPWR
flabel metal1 1448 -6013 1482 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_109/VGND
flabel metal1 1448 -6557 1482 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_109/VPWR
flabel nwell 1448 -6557 1482 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_109/VPB
flabel pwell 1448 -6013 1482 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_109/VNB
rlabel comment 1419 -5996 1419 -5996 2 sky130_fd_sc_hd__decap_4_109/decap_4
rlabel metal1 1419 -6044 1787 -5948 5 sky130_fd_sc_hd__decap_4_109/VGND
rlabel metal1 1419 -6588 1787 -6492 5 sky130_fd_sc_hd__decap_4_109/VPWR
flabel locali 1264 -6183 1298 -6149 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/Y
flabel locali 1264 -6251 1298 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/Y
flabel locali 1172 -6319 1206 -6285 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/Y
flabel locali 1172 -6251 1206 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/Y
flabel locali 1172 -6183 1206 -6149 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/Y
flabel locali 1080 -6115 1114 -6081 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/A
flabel locali 1080 -6183 1114 -6149 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/A
flabel locali 1080 -6251 1114 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_1/A
flabel nwell 1080 -6557 1114 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_1/VPB
flabel pwell 1080 -6013 1114 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_1/VNB
flabel metal1 1080 -6013 1114 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_1/VGND
flabel metal1 1080 -6557 1114 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_1/VPWR
rlabel comment 1051 -5996 1051 -5996 2 sky130_fd_sc_hd__clkinv_1_1/clkinv_1
rlabel metal1 1051 -6044 1327 -5948 5 sky130_fd_sc_hd__clkinv_1_1/VGND
rlabel metal1 1051 -6588 1327 -6492 5 sky130_fd_sc_hd__clkinv_1_1/VPWR
flabel metal1 1809 -6549 1862 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_222/VPWR
flabel metal1 1808 -6016 1859 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_222/VGND
rlabel comment 1787 -5996 1787 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_222/tapvpwrvgnd_1
rlabel metal1 1787 -6044 1879 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_222/VGND
rlabel metal1 1787 -6588 1879 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_222/VPWR
flabel metal1 2269 -6549 2322 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_221/VPWR
flabel metal1 2268 -6016 2319 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_221/VGND
rlabel comment 2247 -5996 2247 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_221/tapvpwrvgnd_1
rlabel metal1 2247 -6044 2339 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_221/VGND
rlabel metal1 2247 -6588 2339 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_221/VPWR
flabel metal1 2920 -6557 2954 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_56/VPWR
flabel metal1 2920 -7101 2954 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_56/VGND
flabel nwell 2920 -6557 2954 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_56/VPB
flabel pwell 2920 -7101 2954 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_56/VNB
rlabel comment 2983 -7084 2983 -7084 6 sky130_fd_sc_hd__decap_8_56/decap_8
rlabel metal1 2247 -7132 2983 -7036 1 sky130_fd_sc_hd__decap_8_56/VGND
rlabel metal1 2247 -6588 2983 -6492 1 sky130_fd_sc_hd__decap_8_56/VPWR
flabel metal1 1908 -6013 1942 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_111/VGND
flabel metal1 1908 -6557 1942 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_111/VPWR
flabel nwell 1908 -6557 1942 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_111/VPB
flabel pwell 1908 -6013 1942 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_111/VNB
rlabel comment 1879 -5996 1879 -5996 2 sky130_fd_sc_hd__decap_4_111/decap_4
rlabel metal1 1879 -6044 2247 -5948 5 sky130_fd_sc_hd__decap_4_111/VGND
rlabel metal1 1879 -6588 2247 -6492 5 sky130_fd_sc_hd__decap_4_111/VPWR
flabel locali 2369 -6251 2403 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A
flabel locali 3015 -6455 3049 -6421 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/X
flabel locali 3015 -6387 3049 -6353 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/X
flabel locali 3015 -6319 3049 -6285 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/X
flabel locali 3015 -6251 3049 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/X
flabel locali 3015 -6183 3049 -6149 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/X
flabel locali 3015 -6115 3049 -6081 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/X
flabel pwell 2369 -6013 2403 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/VNB
flabel nwell 2369 -6557 2403 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/VPB
flabel metal1 2369 -6013 2403 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/VGND
flabel metal1 2369 -6557 2403 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_89/VPWR
rlabel comment 2339 -5996 2339 -5996 2 sky130_fd_sc_hd__clkdlybuf4s50_1_89/clkdlybuf4s50_1
rlabel metal1 2339 -6044 3075 -5948 5 sky130_fd_sc_hd__clkdlybuf4s50_1_89/VGND
rlabel metal1 2339 -6588 3075 -6492 5 sky130_fd_sc_hd__clkdlybuf4s50_1_89/VPWR
flabel metal1 3000 -6560 3053 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_526/VPWR
flabel metal1 3003 -7102 3054 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_526/VGND
rlabel comment 3075 -7084 3075 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_526/tapvpwrvgnd_1
rlabel metal1 2983 -7132 3075 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_526/VGND
rlabel metal1 2983 -6588 3075 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_526/VPWR
flabel metal1 3557 -6549 3610 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_226/VPWR
flabel metal1 3556 -6016 3607 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_226/VGND
rlabel comment 3535 -5996 3535 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_226/tapvpwrvgnd_1
rlabel metal1 3535 -6044 3627 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_226/VGND
rlabel metal1 3535 -6588 3627 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_226/VPWR
flabel metal1 3097 -6549 3150 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_225/VPWR
flabel metal1 3096 -6016 3147 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_225/VGND
rlabel comment 3075 -5996 3075 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_225/tapvpwrvgnd_1
rlabel metal1 3075 -6044 3167 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_225/VGND
rlabel metal1 3075 -6588 3167 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_225/VPWR
flabel metal1 3662 -6006 3694 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_13/VGND
flabel metal1 3656 -6551 3694 -6519 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_13/VPWR
flabel nwell 3647 -6549 3704 -6518 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_13/VPB
flabel pwell 3653 -6006 3697 -5972 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_13/VNB
rlabel comment 3627 -5996 3627 -5996 2 sky130_fd_sc_hd__fill_8_13/fill_8
rlabel metal1 3627 -6044 4363 -5948 5 sky130_fd_sc_hd__fill_8_13/VGND
rlabel metal1 3627 -6588 4363 -6492 5 sky130_fd_sc_hd__fill_8_13/VPWR
flabel metal1 3748 -6557 3782 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_58/VPWR
flabel metal1 3748 -7101 3782 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_58/VGND
flabel nwell 3748 -6557 3782 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_58/VPB
flabel pwell 3748 -7101 3782 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_58/VNB
rlabel comment 3811 -7084 3811 -7084 6 sky130_fd_sc_hd__decap_8_58/decap_8
rlabel metal1 3075 -7132 3811 -7036 1 sky130_fd_sc_hd__decap_8_58/VGND
rlabel metal1 3075 -6588 3811 -6492 1 sky130_fd_sc_hd__decap_8_58/VPWR
flabel metal1 3196 -6013 3230 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_113/VGND
flabel metal1 3196 -6557 3230 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_113/VPWR
flabel nwell 3196 -6557 3230 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_113/VPB
flabel pwell 3196 -6013 3230 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_113/VNB
rlabel comment 3167 -5996 3167 -5996 2 sky130_fd_sc_hd__decap_4_113/decap_4
rlabel metal1 3167 -6044 3535 -5948 5 sky130_fd_sc_hd__decap_4_113/VGND
rlabel metal1 3167 -6588 3535 -6492 5 sky130_fd_sc_hd__decap_4_113/VPWR
flabel metal1 4564 -6560 4617 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_527/VPWR
flabel metal1 4567 -7102 4618 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_527/VGND
rlabel comment 4639 -7084 4639 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_527/tapvpwrvgnd_1
rlabel metal1 4547 -7132 4639 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_527/VGND
rlabel metal1 4547 -6588 4639 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_527/VPWR
flabel metal1 5312 -6557 5346 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_60/VPWR
flabel metal1 5312 -7101 5346 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_60/VGND
flabel nwell 5312 -6557 5346 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_60/VPB
flabel pwell 5312 -7101 5346 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_60/VNB
rlabel comment 5375 -7084 5375 -7084 6 sky130_fd_sc_hd__decap_8_60/decap_8
rlabel metal1 4639 -7132 5375 -7036 1 sky130_fd_sc_hd__decap_8_60/VGND
rlabel metal1 4639 -6588 5375 -6492 1 sky130_fd_sc_hd__decap_8_60/VPWR
flabel metal1 4484 -6557 4518 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_57/VPWR
flabel metal1 4484 -7101 4518 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_57/VGND
flabel nwell 4484 -6557 4518 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_57/VPB
flabel pwell 4484 -7101 4518 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_57/VNB
rlabel comment 4547 -7084 4547 -7084 6 sky130_fd_sc_hd__decap_8_57/decap_8
rlabel metal1 3811 -7132 4547 -7036 1 sky130_fd_sc_hd__decap_8_57/VGND
rlabel metal1 3811 -6588 4547 -6492 1 sky130_fd_sc_hd__decap_8_57/VPWR
flabel metal1 4392 -6013 4426 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_14/VGND
flabel metal1 4392 -6557 4426 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_14/VPWR
flabel nwell 4392 -6557 4426 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_14/VPB
flabel pwell 4392 -6013 4426 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_14/VNB
rlabel comment 4363 -5996 4363 -5996 2 sky130_fd_sc_hd__decap_12_14/decap_12
rlabel metal1 4363 -6044 5467 -5948 5 sky130_fd_sc_hd__decap_12_14/VGND
rlabel metal1 4363 -6588 5467 -6492 5 sky130_fd_sc_hd__decap_12_14/VPWR
flabel metal1 6416 -6013 6450 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_116/VGND
flabel metal1 6416 -6557 6450 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_116/VPWR
flabel nwell 6416 -6557 6450 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_116/VPB
flabel pwell 6416 -6013 6450 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_116/VNB
rlabel comment 6387 -5996 6387 -5996 2 sky130_fd_sc_hd__decap_4_116/decap_4
rlabel metal1 6387 -6044 6755 -5948 5 sky130_fd_sc_hd__decap_4_116/VGND
rlabel metal1 6387 -6588 6755 -6492 5 sky130_fd_sc_hd__decap_4_116/VPWR
flabel metal1 6048 -6557 6082 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_59/VPWR
flabel metal1 6048 -7101 6082 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_59/VGND
flabel nwell 6048 -6557 6082 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_59/VPB
flabel pwell 6048 -7101 6082 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_59/VNB
rlabel comment 6111 -7084 6111 -7084 6 sky130_fd_sc_hd__decap_8_59/decap_8
rlabel metal1 5375 -7132 6111 -7036 1 sky130_fd_sc_hd__decap_8_59/VGND
rlabel metal1 5375 -6588 6111 -6492 1 sky130_fd_sc_hd__decap_8_59/VPWR
flabel metal1 6876 -6557 6910 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_61/VPWR
flabel metal1 6876 -7101 6910 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_61/VGND
flabel nwell 6876 -6557 6910 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_61/VPB
flabel pwell 6876 -7101 6910 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_61/VNB
rlabel comment 6939 -7084 6939 -7084 6 sky130_fd_sc_hd__decap_8_61/decap_8
rlabel metal1 6203 -7132 6939 -7036 1 sky130_fd_sc_hd__decap_8_61/VGND
rlabel metal1 6203 -6588 6939 -6492 1 sky130_fd_sc_hd__decap_8_61/VPWR
flabel metal1 5857 -6553 5893 -6523 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_31/VPWR
flabel metal1 5857 -6012 5893 -5983 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_31/VGND
flabel nwell 5866 -6547 5886 -6530 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_31/VPB
flabel pwell 5863 -6007 5887 -5985 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_31/VNB
rlabel comment 5835 -5996 5835 -5996 2 sky130_fd_sc_hd__fill_1_31/fill_1
rlabel metal1 5835 -6044 5927 -5948 5 sky130_fd_sc_hd__fill_1_31/VGND
rlabel metal1 5835 -6588 5927 -6492 5 sky130_fd_sc_hd__fill_1_31/VPWR
flabel metal1 5961 -6005 5984 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_6/VGND
flabel metal1 5961 -6548 5981 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_6/VPWR
flabel nwell 5962 -6552 5987 -6526 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_6/VPB
flabel pwell 5962 -6008 5984 -5984 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_6/VNB
rlabel comment 5927 -5996 5927 -5996 2 sky130_fd_sc_hd__fill_4_6/fill_4
rlabel metal1 5927 -6044 6295 -5948 5 sky130_fd_sc_hd__fill_4_6/VGND
rlabel metal1 5927 -6588 6295 -6492 5 sky130_fd_sc_hd__fill_4_6/VPWR
flabel metal1 5501 -6005 5524 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_7/VGND
flabel metal1 5501 -6548 5521 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_7/VPWR
flabel nwell 5502 -6552 5527 -6526 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_7/VPB
flabel pwell 5502 -6008 5524 -5984 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_7/VNB
rlabel comment 5467 -5996 5467 -5996 2 sky130_fd_sc_hd__fill_4_7/fill_4
rlabel metal1 5467 -6044 5835 -5948 5 sky130_fd_sc_hd__fill_4_7/VGND
rlabel metal1 5467 -6588 5835 -6492 5 sky130_fd_sc_hd__fill_4_7/VPWR
flabel metal1 6317 -6549 6370 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_232/VPWR
flabel metal1 6316 -6016 6367 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_232/VGND
rlabel comment 6295 -5996 6295 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_232/tapvpwrvgnd_1
rlabel metal1 6295 -6044 6387 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_232/VGND
rlabel metal1 6295 -6588 6387 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_232/VPWR
flabel metal1 6128 -6560 6181 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_528/VPWR
flabel metal1 6131 -7102 6182 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_528/VGND
rlabel comment 6203 -7084 6203 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_528/tapvpwrvgnd_1
rlabel metal1 6111 -7132 6203 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_528/VGND
rlabel metal1 6111 -6588 6203 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_528/VPWR
flabel metal1 6777 -6549 6830 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_234/VPWR
flabel metal1 6776 -6016 6827 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_234/VGND
rlabel comment 6755 -5996 6755 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_234/tapvpwrvgnd_1
rlabel metal1 6755 -6044 6847 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_234/VGND
rlabel metal1 6755 -6588 6847 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_234/VPWR
flabel metal1 7612 -6557 7646 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_62/VPWR
flabel metal1 7612 -7101 7646 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_62/VGND
flabel nwell 7612 -6557 7646 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_62/VPB
flabel pwell 7612 -7101 7646 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_62/VNB
rlabel comment 7675 -7084 7675 -7084 6 sky130_fd_sc_hd__decap_8_62/decap_8
rlabel metal1 6939 -7132 7675 -7036 1 sky130_fd_sc_hd__decap_8_62/VGND
rlabel metal1 6939 -6588 7675 -6492 1 sky130_fd_sc_hd__decap_8_62/VPWR
flabel locali 6877 -6251 6911 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A
flabel locali 7523 -6455 7557 -6421 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/X
flabel locali 7523 -6387 7557 -6353 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/X
flabel locali 7523 -6319 7557 -6285 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/X
flabel locali 7523 -6251 7557 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/X
flabel locali 7523 -6183 7557 -6149 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/X
flabel locali 7523 -6115 7557 -6081 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/X
flabel pwell 6877 -6013 6911 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/VNB
flabel nwell 6877 -6557 6911 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/VPB
flabel metal1 6877 -6013 6911 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/VGND
flabel metal1 6877 -6557 6911 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_93/VPWR
rlabel comment 6847 -5996 6847 -5996 2 sky130_fd_sc_hd__clkdlybuf4s50_1_93/clkdlybuf4s50_1
rlabel metal1 6847 -6044 7583 -5948 5 sky130_fd_sc_hd__clkdlybuf4s50_1_93/VGND
rlabel metal1 6847 -6588 7583 -6492 5 sky130_fd_sc_hd__clkdlybuf4s50_1_93/VPWR
flabel metal1 7692 -6560 7745 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_529/VPWR
flabel metal1 7695 -7102 7746 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_529/VGND
rlabel comment 7767 -7084 7767 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_529/tapvpwrvgnd_1
rlabel metal1 7675 -7132 7767 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_529/VGND
rlabel metal1 7675 -6588 7767 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_529/VPWR
flabel metal1 7605 -6549 7658 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_237/VPWR
flabel metal1 7604 -6016 7655 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_237/VGND
rlabel comment 7583 -5996 7583 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_237/tapvpwrvgnd_1
rlabel metal1 7583 -6044 7675 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_237/VGND
rlabel metal1 7583 -6588 7675 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_237/VPWR
flabel metal1 8065 -6549 8118 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_236/VPWR
flabel metal1 8064 -6016 8115 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_236/VGND
rlabel comment 8043 -5996 8043 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_236/tapvpwrvgnd_1
rlabel metal1 8043 -6044 8135 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_236/VGND
rlabel metal1 8043 -6588 8135 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_236/VPWR
flabel metal1 8440 -6557 8474 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_63/VPWR
flabel metal1 8440 -7101 8474 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_63/VGND
flabel nwell 8440 -6557 8474 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_63/VPB
flabel pwell 8440 -7101 8474 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_63/VNB
rlabel comment 8503 -7084 8503 -7084 6 sky130_fd_sc_hd__decap_8_63/decap_8
rlabel metal1 7767 -7132 8503 -7036 1 sky130_fd_sc_hd__decap_8_63/VGND
rlabel metal1 7767 -6588 8503 -6492 1 sky130_fd_sc_hd__decap_8_63/VPWR
flabel metal1 7704 -6013 7738 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_118/VGND
flabel metal1 7704 -6557 7738 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_118/VPWR
flabel nwell 7704 -6557 7738 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_118/VPB
flabel pwell 7704 -6013 7738 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_118/VNB
rlabel comment 7675 -5996 7675 -5996 2 sky130_fd_sc_hd__decap_4_118/decap_4
rlabel metal1 7675 -6044 8043 -5948 5 sky130_fd_sc_hd__decap_4_118/VGND
rlabel metal1 7675 -6588 8043 -6492 5 sky130_fd_sc_hd__decap_4_118/VPWR
flabel locali 8165 -6251 8199 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A
flabel locali 8811 -6455 8845 -6421 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/X
flabel locali 8811 -6387 8845 -6353 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/X
flabel locali 8811 -6319 8845 -6285 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/X
flabel locali 8811 -6251 8845 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/X
flabel locali 8811 -6183 8845 -6149 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/X
flabel locali 8811 -6115 8845 -6081 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/X
flabel pwell 8165 -6013 8199 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/VNB
flabel nwell 8165 -6557 8199 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/VPB
flabel metal1 8165 -6013 8199 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/VGND
flabel metal1 8165 -6557 8199 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_95/VPWR
rlabel comment 8135 -5996 8135 -5996 2 sky130_fd_sc_hd__clkdlybuf4s50_1_95/clkdlybuf4s50_1
rlabel metal1 8135 -6044 8871 -5948 5 sky130_fd_sc_hd__clkdlybuf4s50_1_95/VGND
rlabel metal1 8135 -6588 8871 -6492 5 sky130_fd_sc_hd__clkdlybuf4s50_1_95/VPWR
flabel metal1 9176 -6557 9210 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_65/VPWR
flabel metal1 9176 -7101 9210 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_65/VGND
flabel nwell 9176 -6557 9210 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_65/VPB
flabel pwell 9176 -7101 9210 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_65/VNB
rlabel comment 9239 -7084 9239 -7084 6 sky130_fd_sc_hd__decap_8_65/decap_8
rlabel metal1 8503 -7132 9239 -7036 1 sky130_fd_sc_hd__decap_8_65/VGND
rlabel metal1 8503 -6588 9239 -6492 1 sky130_fd_sc_hd__decap_8_65/VPWR
flabel locali 9453 -6251 9487 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A
flabel locali 10099 -6455 10133 -6421 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/X
flabel locali 10099 -6387 10133 -6353 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/X
flabel locali 10099 -6319 10133 -6285 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/X
flabel locali 10099 -6251 10133 -6217 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/X
flabel locali 10099 -6183 10133 -6149 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/X
flabel locali 10099 -6115 10133 -6081 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/X
flabel pwell 9453 -6013 9487 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/VNB
flabel nwell 9453 -6557 9487 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/VPB
flabel metal1 9453 -6013 9487 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/VGND
flabel metal1 9453 -6557 9487 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_97/VPWR
rlabel comment 9423 -5996 9423 -5996 2 sky130_fd_sc_hd__clkdlybuf4s50_1_97/clkdlybuf4s50_1
rlabel metal1 9423 -6044 10159 -5948 5 sky130_fd_sc_hd__clkdlybuf4s50_1_97/VGND
rlabel metal1 9423 -6588 10159 -6492 5 sky130_fd_sc_hd__clkdlybuf4s50_1_97/VPWR
flabel metal1 8992 -6013 9026 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_120/VGND
flabel metal1 8992 -6557 9026 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_120/VPWR
flabel nwell 8992 -6557 9026 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_120/VPB
flabel pwell 8992 -6013 9026 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_120/VNB
rlabel comment 8963 -5996 8963 -5996 2 sky130_fd_sc_hd__decap_4_120/decap_4
rlabel metal1 8963 -6044 9331 -5948 5 sky130_fd_sc_hd__decap_4_120/VGND
rlabel metal1 8963 -6588 9331 -6492 5 sky130_fd_sc_hd__decap_4_120/VPWR
flabel metal1 10280 -6013 10314 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_122/VGND
flabel metal1 10280 -6557 10314 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_122/VPWR
flabel nwell 10280 -6557 10314 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_122/VPB
flabel pwell 10280 -6013 10314 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_122/VNB
rlabel comment 10251 -5996 10251 -5996 2 sky130_fd_sc_hd__decap_4_122/decap_4
rlabel metal1 10251 -6044 10619 -5948 5 sky130_fd_sc_hd__decap_4_122/VGND
rlabel metal1 10251 -6588 10619 -6492 5 sky130_fd_sc_hd__decap_4_122/VPWR
flabel metal1 9366 -7104 9398 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_36/VGND
flabel metal1 9360 -6561 9398 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_36/VPWR
flabel nwell 9351 -6562 9408 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_36/VPB
flabel pwell 9357 -7108 9401 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_36/VNB
rlabel comment 9331 -7084 9331 -7084 4 sky130_fd_sc_hd__fill_8_36/fill_8
rlabel metal1 9331 -7132 10067 -7036 1 sky130_fd_sc_hd__fill_8_36/VGND
rlabel metal1 9331 -6588 10067 -6492 1 sky130_fd_sc_hd__fill_8_36/VPWR
flabel metal1 10102 -7104 10134 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_39/VGND
flabel metal1 10096 -6561 10134 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_39/VPWR
flabel nwell 10087 -6562 10144 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_39/VPB
flabel pwell 10093 -7108 10137 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_39/VNB
rlabel comment 10067 -7084 10067 -7084 4 sky130_fd_sc_hd__fill_8_39/fill_8
rlabel metal1 10067 -7132 10803 -7036 1 sky130_fd_sc_hd__fill_8_39/VGND
rlabel metal1 10067 -6588 10803 -6492 1 sky130_fd_sc_hd__fill_8_39/VPWR
flabel metal1 8893 -6549 8946 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_240/VPWR
flabel metal1 8892 -6016 8943 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_240/VGND
rlabel comment 8871 -5996 8871 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_240/tapvpwrvgnd_1
rlabel metal1 8871 -6044 8963 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_240/VGND
rlabel metal1 8871 -6588 8963 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_240/VPWR
flabel metal1 9353 -6549 9406 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_242/VPWR
flabel metal1 9352 -6016 9403 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_242/VGND
rlabel comment 9331 -5996 9331 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_242/tapvpwrvgnd_1
rlabel metal1 9331 -6044 9423 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_242/VGND
rlabel metal1 9331 -6588 9423 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_242/VPWR
flabel metal1 10181 -6549 10234 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_244/VPWR
flabel metal1 10180 -6016 10231 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_244/VGND
rlabel comment 10159 -5996 10159 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_244/tapvpwrvgnd_1
rlabel metal1 10159 -6044 10251 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_244/VGND
rlabel metal1 10159 -6588 10251 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_244/VPWR
flabel metal1 9256 -6560 9309 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_530/VPWR
flabel metal1 9259 -7102 9310 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_530/VGND
rlabel comment 9331 -7084 9331 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_530/tapvpwrvgnd_1
rlabel metal1 9239 -7132 9331 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_530/VGND
rlabel metal1 9239 -6588 9331 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_530/VPWR
flabel metal1 11660 -6013 11694 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_124/VGND
flabel metal1 11660 -6557 11694 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_124/VPWR
flabel nwell 11660 -6557 11694 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_124/VPB
flabel pwell 11660 -6013 11694 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_124/VNB
rlabel comment 11631 -5996 11631 -5996 2 sky130_fd_sc_hd__decap_4_124/decap_4
rlabel metal1 11631 -6044 11999 -5948 5 sky130_fd_sc_hd__decap_4_124/VGND
rlabel metal1 11631 -6588 11999 -6492 5 sky130_fd_sc_hd__decap_4_124/VPWR
flabel metal1 12034 -6006 12066 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_14/VGND
flabel metal1 12028 -6551 12066 -6519 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_14/VPWR
flabel nwell 12019 -6549 12076 -6518 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_14/VPB
flabel pwell 12025 -6006 12069 -5972 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_14/VNB
rlabel comment 11999 -5996 11999 -5996 2 sky130_fd_sc_hd__fill_8_14/fill_8
rlabel metal1 11999 -6044 12735 -5948 5 sky130_fd_sc_hd__fill_8_14/VGND
rlabel metal1 11999 -6588 12735 -6492 5 sky130_fd_sc_hd__fill_8_14/VPWR
flabel metal1 10838 -7104 10870 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_42/VGND
flabel metal1 10832 -6561 10870 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_42/VPWR
flabel nwell 10823 -6562 10880 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_42/VPB
flabel pwell 10829 -7108 10873 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_42/VNB
rlabel comment 10803 -7084 10803 -7084 4 sky130_fd_sc_hd__fill_8_42/fill_8
rlabel metal1 10803 -7132 11539 -7036 1 sky130_fd_sc_hd__fill_8_42/VGND
rlabel metal1 10803 -6588 11539 -6492 1 sky130_fd_sc_hd__fill_8_42/VPWR
flabel metal1 11574 -7104 11606 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_43/VGND
flabel metal1 11568 -6561 11606 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_43/VPWR
flabel nwell 11559 -6562 11616 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_43/VPB
flabel pwell 11565 -7108 11609 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_43/VNB
rlabel comment 11539 -7084 11539 -7084 4 sky130_fd_sc_hd__fill_8_43/fill_8
rlabel metal1 11539 -7132 12275 -7036 1 sky130_fd_sc_hd__fill_8_43/VGND
rlabel metal1 11539 -6588 12275 -6492 1 sky130_fd_sc_hd__fill_8_43/VPWR
flabel metal1 12310 -7104 12342 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_46/VGND
flabel metal1 12304 -6561 12342 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_46/VPWR
flabel nwell 12295 -6562 12352 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_46/VPB
flabel pwell 12301 -7108 12345 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_46/VNB
rlabel comment 12275 -7084 12275 -7084 4 sky130_fd_sc_hd__fill_8_46/fill_8
rlabel metal1 12275 -7132 13011 -7036 1 sky130_fd_sc_hd__fill_8_46/VGND
rlabel metal1 12275 -6588 13011 -6492 1 sky130_fd_sc_hd__fill_8_46/VPWR
flabel locali 11109 -6251 11143 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/Y
flabel locali 11109 -6319 11143 -6285 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/Y
flabel locali 11385 -6251 11419 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/A
flabel locali 11293 -6251 11327 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/A
flabel locali 11017 -6251 11051 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 10925 -6251 10959 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 10741 -6251 10775 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 10833 -6251 10867 -6217 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel nwell 10741 -6557 10775 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VPB
flabel pwell 10741 -6013 10775 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VNB
flabel metal1 10741 -6013 10775 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VGND
flabel metal1 10741 -6557 10775 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VPWR
rlabel comment 10711 -5996 10711 -5996 2 sky130_fd_sc_hd__nand2_4_1/nand2_4
rlabel metal1 10711 -6044 11539 -5948 5 sky130_fd_sc_hd__nand2_4_1/VGND
rlabel metal1 10711 -6588 11539 -6492 5 sky130_fd_sc_hd__nand2_4_1/VPWR
flabel metal1 10641 -6549 10694 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_246/VPWR
flabel metal1 10640 -6016 10691 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_246/VGND
rlabel comment 10619 -5996 10619 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_246/tapvpwrvgnd_1
rlabel metal1 10619 -6044 10711 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_246/VGND
rlabel metal1 10619 -6588 10711 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_246/VPWR
flabel metal1 11561 -6549 11614 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_247/VPWR
flabel metal1 11560 -6016 11611 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_247/VGND
rlabel comment 11539 -5996 11539 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_247/tapvpwrvgnd_1
rlabel metal1 11539 -6044 11631 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_247/VGND
rlabel metal1 11539 -6588 11631 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_247/VPWR
flabel metal1 13592 -6013 13626 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_15/VGND
flabel metal1 13592 -6557 13626 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_15/VPWR
flabel nwell 13592 -6557 13626 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_15/VPB
flabel pwell 13592 -6013 13626 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_15/VNB
rlabel comment 13563 -5996 13563 -5996 2 sky130_fd_sc_hd__decap_12_15/decap_12
rlabel metal1 13563 -6044 14667 -5948 5 sky130_fd_sc_hd__decap_12_15/VGND
rlabel metal1 13563 -6588 14667 -6492 5 sky130_fd_sc_hd__decap_12_15/VPWR
flabel metal1 12770 -6006 12802 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_17/VGND
flabel metal1 12764 -6551 12802 -6519 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_17/VPWR
flabel nwell 12755 -6549 12812 -6518 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_17/VPB
flabel pwell 12761 -6006 12805 -5972 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_17/VNB
rlabel comment 12735 -5996 12735 -5996 2 sky130_fd_sc_hd__fill_8_17/fill_8
rlabel metal1 12735 -6044 13471 -5948 5 sky130_fd_sc_hd__fill_8_17/VGND
rlabel metal1 12735 -6588 13471 -6492 5 sky130_fd_sc_hd__fill_8_17/VPWR
flabel metal1 13046 -7104 13078 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_47/VGND
flabel metal1 13040 -6561 13078 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_47/VPWR
flabel nwell 13031 -6562 13088 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_47/VPB
flabel pwell 13037 -7108 13081 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_47/VNB
rlabel comment 13011 -7084 13011 -7084 4 sky130_fd_sc_hd__fill_8_47/fill_8
rlabel metal1 13011 -7132 13747 -7036 1 sky130_fd_sc_hd__fill_8_47/VGND
rlabel metal1 13011 -6588 13747 -6492 1 sky130_fd_sc_hd__fill_8_47/VPWR
flabel metal1 13782 -7104 13814 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_50/VGND
flabel metal1 13776 -6561 13814 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_50/VPWR
flabel nwell 13767 -6562 13824 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_50/VPB
flabel pwell 13773 -7108 13817 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_50/VNB
rlabel comment 13747 -7084 13747 -7084 4 sky130_fd_sc_hd__fill_8_50/fill_8
rlabel metal1 13747 -7132 14483 -7036 1 sky130_fd_sc_hd__fill_8_50/VGND
rlabel metal1 13747 -6588 14483 -6492 1 sky130_fd_sc_hd__fill_8_50/VPWR
flabel metal1 13493 -6549 13546 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_250/VPWR
flabel metal1 13492 -6016 13543 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_250/VGND
rlabel comment 13471 -5996 13471 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_250/tapvpwrvgnd_1
rlabel metal1 13471 -6044 13563 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_250/VGND
rlabel metal1 13471 -6588 13563 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_250/VPWR
flabel metal1 15984 -6557 16018 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_21/VPWR
flabel metal1 15984 -6013 16018 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_21/VGND
flabel nwell 15984 -6557 16018 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_21/VPB
flabel pwell 15984 -6013 16018 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_21/VNB
rlabel comment 15955 -5996 15955 -5996 2 sky130_fd_sc_hd__decap_8_21/decap_8
rlabel metal1 15955 -6044 16691 -5948 5 sky130_fd_sc_hd__decap_8_21/VGND
rlabel metal1 15955 -6588 16691 -6492 5 sky130_fd_sc_hd__decap_8_21/VPWR
flabel metal1 16628 -6557 16662 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_66/VPWR
flabel metal1 16628 -7101 16662 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_66/VGND
flabel nwell 16628 -6557 16662 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_66/VPB
flabel pwell 16628 -7101 16662 -7067 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_66/VNB
rlabel comment 16691 -7084 16691 -7084 6 sky130_fd_sc_hd__decap_8_66/decap_8
rlabel metal1 15955 -7132 16691 -7036 1 sky130_fd_sc_hd__decap_8_66/VGND
rlabel metal1 15955 -6588 16691 -6492 1 sky130_fd_sc_hd__decap_8_66/VPWR
flabel metal1 14788 -6013 14822 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_16/VGND
flabel metal1 14788 -6557 14822 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_16/VPWR
flabel nwell 14788 -6557 14822 -6523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_16/VPB
flabel pwell 14788 -6013 14822 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_16/VNB
rlabel comment 14759 -5996 14759 -5996 2 sky130_fd_sc_hd__decap_12_16/decap_12
rlabel metal1 14759 -6044 15863 -5948 5 sky130_fd_sc_hd__decap_12_16/VGND
rlabel metal1 14759 -6588 15863 -6492 5 sky130_fd_sc_hd__decap_12_16/VPWR
flabel metal1 14518 -7104 14550 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_51/VGND
flabel metal1 14512 -6561 14550 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_51/VPWR
flabel nwell 14503 -6562 14560 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_51/VPB
flabel pwell 14509 -7108 14553 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_51/VNB
rlabel comment 14483 -7084 14483 -7084 4 sky130_fd_sc_hd__fill_8_51/fill_8
rlabel metal1 14483 -7132 15219 -7036 1 sky130_fd_sc_hd__fill_8_51/VGND
rlabel metal1 14483 -6588 15219 -6492 1 sky130_fd_sc_hd__fill_8_51/VPWR
flabel metal1 15254 -7104 15286 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_52/VGND
flabel metal1 15248 -6561 15286 -6529 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_52/VPWR
flabel nwell 15239 -6562 15296 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_52/VPB
flabel pwell 15245 -7108 15289 -7074 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_52/VNB
rlabel comment 15219 -7084 15219 -7084 4 sky130_fd_sc_hd__fill_8_52/fill_8
rlabel metal1 15219 -7132 15955 -7036 1 sky130_fd_sc_hd__fill_8_52/VGND
rlabel metal1 15219 -6588 15955 -6492 1 sky130_fd_sc_hd__fill_8_52/VPWR
flabel metal1 14689 -6549 14742 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_251/VPWR
flabel metal1 14688 -6016 14739 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_251/VGND
rlabel comment 14667 -5996 14667 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_251/tapvpwrvgnd_1
rlabel metal1 14667 -6044 14759 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_251/VGND
rlabel metal1 14667 -6588 14759 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_251/VPWR
flabel metal1 15885 -6549 15938 -6520 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_253/VPWR
flabel metal1 15884 -6016 15935 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_253/VGND
rlabel comment 15863 -5996 15863 -5996 2 sky130_fd_sc_hd__tapvpwrvgnd_1_253/tapvpwrvgnd_1
rlabel metal1 15863 -6044 15955 -5948 5 sky130_fd_sc_hd__tapvpwrvgnd_1_253/VGND
rlabel metal1 15863 -6588 15955 -6492 5 sky130_fd_sc_hd__tapvpwrvgnd_1_253/VPWR
flabel metal1 15880 -6560 15933 -6531 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_521/VPWR
flabel metal1 15883 -7102 15934 -7064 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_521/VGND
rlabel comment 15955 -7084 15955 -7084 6 sky130_fd_sc_hd__tapvpwrvgnd_1_521/tapvpwrvgnd_1
rlabel metal1 15863 -7132 15955 -7036 1 sky130_fd_sc_hd__tapvpwrvgnd_1_521/VGND
rlabel metal1 15863 -6588 15955 -6492 1 sky130_fd_sc_hd__tapvpwrvgnd_1_521/VPWR
flabel metal1 -944 -5469 -910 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_19/VPWR
flabel metal1 -944 -6013 -910 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_19/VGND
flabel nwell -944 -5469 -910 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_19/VPB
flabel pwell -944 -6013 -910 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_19/VNB
rlabel comment -881 -5996 -881 -5996 6 sky130_fd_sc_hd__decap_8_19/decap_8
rlabel metal1 -1617 -6044 -881 -5948 1 sky130_fd_sc_hd__decap_8_19/VGND
rlabel metal1 -1617 -5500 -881 -5404 1 sky130_fd_sc_hd__decap_8_19/VPWR
flabel metal1 -2968 -5469 -2934 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_77/VPWR
flabel metal1 -2968 -6013 -2934 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_77/VGND
flabel nwell -2968 -5469 -2934 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_77/VPB
flabel pwell -2968 -6013 -2934 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_77/VNB
rlabel comment -2997 -5996 -2997 -5996 4 sky130_fd_sc_hd__decap_8_77/decap_8
rlabel metal1 -2997 -6044 -2261 -5948 1 sky130_fd_sc_hd__decap_8_77/VGND
rlabel metal1 -2997 -5500 -2261 -5404 1 sky130_fd_sc_hd__decap_8_77/VPWR
flabel metal1 -1781 -6010 -1728 -5978 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_14/VGND
flabel metal1 -1780 -5466 -1728 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_14/VPWR
flabel nwell -1773 -5461 -1739 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_14/VPB
flabel pwell -1770 -6006 -1738 -5984 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_14/VNB
rlabel comment -1801 -5996 -1801 -5996 4 sky130_fd_sc_hd__fill_2_14/fill_2
rlabel metal1 -1801 -6044 -1617 -5948 1 sky130_fd_sc_hd__fill_2_14/VGND
rlabel metal1 -1801 -5500 -1617 -5404 1 sky130_fd_sc_hd__fill_2_14/VPWR
flabel metal1 -2135 -6006 -2112 -5987 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_27/VGND
flabel metal1 -2135 -5461 -2115 -5444 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_27/VPWR
flabel nwell -2134 -5466 -2109 -5440 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_27/VPB
flabel pwell -2134 -6008 -2112 -5984 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_27/VNB
rlabel comment -2169 -5996 -2169 -5996 4 sky130_fd_sc_hd__fill_4_27/fill_4
rlabel metal1 -2169 -6044 -1801 -5948 1 sky130_fd_sc_hd__fill_4_27/VGND
rlabel metal1 -2169 -5500 -1801 -5404 1 sky130_fd_sc_hd__fill_4_27/VPWR
flabel metal1 -2239 -5472 -2186 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_542/VPWR
flabel metal1 -2240 -6014 -2189 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_542/VGND
rlabel comment -2261 -5996 -2261 -5996 4 sky130_fd_sc_hd__tapvpwrvgnd_1_542/tapvpwrvgnd_1
rlabel metal1 -2261 -6044 -2169 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_542/VGND
rlabel metal1 -2261 -5500 -2169 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_542/VPWR
flabel locali 1079 -5775 1113 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/A
flabel locali 433 -5571 467 -5537 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X
flabel locali 433 -5639 467 -5605 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X
flabel locali 433 -5707 467 -5673 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X
flabel locali 433 -5775 467 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X
flabel locali 433 -5843 467 -5809 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X
flabel locali 433 -5911 467 -5877 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X
flabel pwell 1079 -6013 1113 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/VNB
flabel nwell 1079 -5469 1113 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/VPB
flabel metal1 1079 -6013 1113 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/VGND
flabel metal1 1079 -5469 1113 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_87/VPWR
rlabel comment 1143 -5996 1143 -5996 6 sky130_fd_sc_hd__clkdlybuf4s50_1_87/clkdlybuf4s50_1
rlabel metal1 407 -6044 1143 -5948 1 sky130_fd_sc_hd__clkdlybuf4s50_1_87/VGND
rlabel metal1 407 -5500 1143 -5404 1 sky130_fd_sc_hd__clkdlybuf4s50_1_87/VPWR
flabel metal1 252 -6013 286 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_107/VGND
flabel metal1 252 -5469 286 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_107/VPWR
flabel nwell 252 -5469 286 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_107/VPB
flabel pwell 252 -6013 286 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_107/VNB
rlabel comment 315 -5996 315 -5996 6 sky130_fd_sc_hd__decap_4_107/decap_4
rlabel metal1 -53 -6044 315 -5948 1 sky130_fd_sc_hd__decap_4_107/VGND
rlabel metal1 -53 -5500 315 -5404 1 sky130_fd_sc_hd__decap_4_107/VPWR
flabel metal1 -208 -5469 -174 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_20/VPWR
flabel metal1 -208 -6013 -174 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_20/VGND
flabel nwell -208 -5469 -174 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_20/VPB
flabel pwell -208 -6013 -174 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_20/VNB
rlabel comment -145 -5996 -145 -5996 6 sky130_fd_sc_hd__decap_8_20/decap_8
rlabel metal1 -881 -6044 -145 -5948 1 sky130_fd_sc_hd__decap_8_20/VGND
rlabel metal1 -881 -5500 -145 -5404 1 sky130_fd_sc_hd__decap_8_20/VPWR
flabel metal1 -128 -5472 -75 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_214/VPWR
flabel metal1 -125 -6014 -74 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_214/VGND
rlabel comment -53 -5996 -53 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_214/tapvpwrvgnd_1
rlabel metal1 -145 -6044 -53 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_214/VGND
rlabel metal1 -145 -5500 -53 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_214/VPWR
flabel metal1 332 -5472 385 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_215/VPWR
flabel metal1 335 -6014 386 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_215/VGND
rlabel comment 407 -5996 407 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_215/tapvpwrvgnd_1
rlabel metal1 315 -6044 407 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_215/VGND
rlabel metal1 315 -5500 407 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_215/VPWR
flabel metal1 1540 -6013 1574 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_110/VGND
flabel metal1 1540 -5469 1574 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_110/VPWR
flabel nwell 1540 -5469 1574 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_110/VPB
flabel pwell 1540 -6013 1574 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_110/VNB
rlabel comment 1603 -5996 1603 -5996 6 sky130_fd_sc_hd__decap_4_110/decap_4
rlabel metal1 1235 -6044 1603 -5948 1 sky130_fd_sc_hd__decap_4_110/VGND
rlabel metal1 1235 -5500 1603 -5404 1 sky130_fd_sc_hd__decap_4_110/VPWR
flabel metal1 2828 -6013 2862 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_112/VGND
flabel metal1 2828 -5469 2862 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_112/VPWR
flabel nwell 2828 -5469 2862 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_112/VPB
flabel pwell 2828 -6013 2862 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_112/VNB
rlabel comment 2891 -5996 2891 -5996 6 sky130_fd_sc_hd__decap_4_112/decap_4
rlabel metal1 2523 -6044 2891 -5948 1 sky130_fd_sc_hd__decap_4_112/VGND
rlabel metal1 2523 -5500 2891 -5404 1 sky130_fd_sc_hd__decap_4_112/VPWR
flabel metal1 1724 -5469 1758 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_100/VPWR
flabel metal1 1724 -6013 1758 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_100/VGND
flabel nwell 1724 -5469 1758 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_100/VPB
flabel pwell 1724 -6013 1758 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_100/VNB
rlabel comment 1695 -5996 1695 -5996 4 sky130_fd_sc_hd__decap_8_100/decap_8
rlabel metal1 1695 -6044 2431 -5948 1 sky130_fd_sc_hd__decap_8_100/VGND
rlabel metal1 1695 -5500 2431 -5404 1 sky130_fd_sc_hd__decap_8_100/VPWR
flabel metal1 1160 -5472 1213 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_220/VPWR
flabel metal1 1163 -6014 1214 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_220/VGND
rlabel comment 1235 -5996 1235 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_220/tapvpwrvgnd_1
rlabel metal1 1143 -6044 1235 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_220/VGND
rlabel metal1 1143 -5500 1235 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_220/VPWR
flabel metal1 1620 -5472 1673 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_223/VPWR
flabel metal1 1623 -6014 1674 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_223/VGND
rlabel comment 1695 -5996 1695 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_223/tapvpwrvgnd_1
rlabel metal1 1603 -6044 1695 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_223/VGND
rlabel metal1 1603 -5500 1695 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_223/VPWR
flabel metal1 2448 -5472 2501 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_224/VPWR
flabel metal1 2451 -6014 2502 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_224/VGND
rlabel comment 2523 -5996 2523 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_224/tapvpwrvgnd_1
rlabel metal1 2431 -6044 2523 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_224/VGND
rlabel metal1 2431 -5500 2523 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_224/VPWR
flabel locali 3655 -5775 3689 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/A
flabel locali 3009 -5571 3043 -5537 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X
flabel locali 3009 -5639 3043 -5605 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X
flabel locali 3009 -5707 3043 -5673 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X
flabel locali 3009 -5775 3043 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X
flabel locali 3009 -5843 3043 -5809 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X
flabel locali 3009 -5911 3043 -5877 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X
flabel pwell 3655 -6013 3689 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/VNB
flabel nwell 3655 -5469 3689 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/VPB
flabel metal1 3655 -6013 3689 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/VGND
flabel metal1 3655 -5469 3689 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_90/VPWR
rlabel comment 3719 -5996 3719 -5996 6 sky130_fd_sc_hd__clkdlybuf4s50_1_90/clkdlybuf4s50_1
rlabel metal1 2983 -6044 3719 -5948 1 sky130_fd_sc_hd__clkdlybuf4s50_1_90/VGND
rlabel metal1 2983 -5500 3719 -5404 1 sky130_fd_sc_hd__clkdlybuf4s50_1_90/VPWR
flabel metal1 4116 -6013 4150 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_114/VGND
flabel metal1 4116 -5469 4150 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_114/VPWR
flabel nwell 4116 -5469 4150 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_114/VPB
flabel pwell 4116 -6013 4150 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_114/VNB
rlabel comment 4179 -5996 4179 -5996 6 sky130_fd_sc_hd__decap_4_114/decap_4
rlabel metal1 3811 -6044 4179 -5948 1 sky130_fd_sc_hd__decap_4_114/VGND
rlabel metal1 3811 -5500 4179 -5404 1 sky130_fd_sc_hd__decap_4_114/VPWR
flabel metal1 4300 -5469 4334 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_101/VPWR
flabel metal1 4300 -6013 4334 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_101/VGND
flabel nwell 4300 -5469 4334 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_101/VPB
flabel pwell 4300 -6013 4334 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_101/VNB
rlabel comment 4271 -5996 4271 -5996 4 sky130_fd_sc_hd__decap_8_101/decap_8
rlabel metal1 4271 -6044 5007 -5948 1 sky130_fd_sc_hd__decap_8_101/VGND
rlabel metal1 4271 -5500 5007 -5404 1 sky130_fd_sc_hd__decap_8_101/VPWR
flabel metal1 2908 -5472 2961 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_227/VPWR
flabel metal1 2911 -6014 2962 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_227/VGND
rlabel comment 2983 -5996 2983 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_227/tapvpwrvgnd_1
rlabel metal1 2891 -6044 2983 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_227/VGND
rlabel metal1 2891 -5500 2983 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_227/VPWR
flabel metal1 4196 -5472 4249 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_228/VPWR
flabel metal1 4199 -6014 4250 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_228/VGND
rlabel comment 4271 -5996 4271 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_228/tapvpwrvgnd_1
rlabel metal1 4179 -6044 4271 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_228/VGND
rlabel metal1 4179 -5500 4271 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_228/VPWR
flabel metal1 3736 -5472 3789 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_229/VPWR
flabel metal1 3739 -6014 3790 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_229/VGND
rlabel comment 3811 -5996 3811 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_229/tapvpwrvgnd_1
rlabel metal1 3719 -6044 3811 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_229/VGND
rlabel metal1 3719 -5500 3811 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_229/VPWR
flabel locali 6231 -5775 6265 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/A
flabel locali 5585 -5571 5619 -5537 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
flabel locali 5585 -5639 5619 -5605 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
flabel locali 5585 -5707 5619 -5673 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
flabel locali 5585 -5775 5619 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
flabel locali 5585 -5843 5619 -5809 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
flabel locali 5585 -5911 5619 -5877 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
flabel pwell 6231 -6013 6265 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/VNB
flabel nwell 6231 -5469 6265 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/VPB
flabel metal1 6231 -6013 6265 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/VGND
flabel metal1 6231 -5469 6265 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_92/VPWR
rlabel comment 6295 -5996 6295 -5996 6 sky130_fd_sc_hd__clkdlybuf4s50_1_92/clkdlybuf4s50_1
rlabel metal1 5559 -6044 6295 -5948 1 sky130_fd_sc_hd__clkdlybuf4s50_1_92/VGND
rlabel metal1 5559 -5500 6295 -5404 1 sky130_fd_sc_hd__clkdlybuf4s50_1_92/VPWR
flabel metal1 5404 -6013 5438 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_115/VGND
flabel metal1 5404 -5469 5438 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_115/VPWR
flabel nwell 5404 -5469 5438 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_115/VPB
flabel pwell 5404 -6013 5438 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_115/VNB
rlabel comment 5467 -5996 5467 -5996 6 sky130_fd_sc_hd__decap_4_115/decap_4
rlabel metal1 5099 -6044 5467 -5948 1 sky130_fd_sc_hd__decap_4_115/VGND
rlabel metal1 5099 -5500 5467 -5404 1 sky130_fd_sc_hd__decap_4_115/VPWR
flabel metal1 6692 -6013 6726 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_117/VGND
flabel metal1 6692 -5469 6726 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_117/VPWR
flabel nwell 6692 -5469 6726 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_117/VPB
flabel pwell 6692 -6013 6726 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_117/VNB
rlabel comment 6755 -5996 6755 -5996 6 sky130_fd_sc_hd__decap_4_117/decap_4
rlabel metal1 6387 -6044 6755 -5948 1 sky130_fd_sc_hd__decap_4_117/VGND
rlabel metal1 6387 -5500 6755 -5404 1 sky130_fd_sc_hd__decap_4_117/VPWR
flabel metal1 5024 -5472 5077 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_230/VPWR
flabel metal1 5027 -6014 5078 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_230/VGND
rlabel comment 5099 -5996 5099 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_230/tapvpwrvgnd_1
rlabel metal1 5007 -6044 5099 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_230/VGND
rlabel metal1 5007 -5500 5099 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_230/VPWR
flabel metal1 5484 -5472 5537 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_231/VPWR
flabel metal1 5487 -6014 5538 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_231/VGND
rlabel comment 5559 -5996 5559 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_231/tapvpwrvgnd_1
rlabel metal1 5467 -6044 5559 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_231/VGND
rlabel metal1 5467 -5500 5559 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_231/VPWR
flabel metal1 6312 -5472 6365 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_233/VPWR
flabel metal1 6315 -6014 6366 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_233/VGND
rlabel comment 6387 -5996 6387 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_233/tapvpwrvgnd_1
rlabel metal1 6295 -6044 6387 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_233/VGND
rlabel metal1 6295 -5500 6387 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_233/VPWR
flabel locali 8807 -5775 8841 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/A
flabel locali 8161 -5571 8195 -5537 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X
flabel locali 8161 -5639 8195 -5605 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X
flabel locali 8161 -5707 8195 -5673 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X
flabel locali 8161 -5775 8195 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X
flabel locali 8161 -5843 8195 -5809 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X
flabel locali 8161 -5911 8195 -5877 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X
flabel pwell 8807 -6013 8841 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/VNB
flabel nwell 8807 -5469 8841 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/VPB
flabel metal1 8807 -6013 8841 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/VGND
flabel metal1 8807 -5469 8841 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_96/VPWR
rlabel comment 8871 -5996 8871 -5996 6 sky130_fd_sc_hd__clkdlybuf4s50_1_96/clkdlybuf4s50_1
rlabel metal1 8135 -6044 8871 -5948 1 sky130_fd_sc_hd__clkdlybuf4s50_1_96/VGND
rlabel metal1 8135 -5500 8871 -5404 1 sky130_fd_sc_hd__clkdlybuf4s50_1_96/VPWR
flabel metal1 7980 -6013 8014 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_119/VGND
flabel metal1 7980 -5469 8014 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_119/VPWR
flabel nwell 7980 -5469 8014 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_119/VPB
flabel pwell 7980 -6013 8014 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_119/VNB
rlabel comment 8043 -5996 8043 -5996 6 sky130_fd_sc_hd__decap_4_119/decap_4
rlabel metal1 7675 -6044 8043 -5948 1 sky130_fd_sc_hd__decap_4_119/VGND
rlabel metal1 7675 -5500 8043 -5404 1 sky130_fd_sc_hd__decap_4_119/VPWR
flabel metal1 6876 -5469 6910 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_112/VPWR
flabel metal1 6876 -6013 6910 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_112/VGND
flabel nwell 6876 -5469 6910 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_112/VPB
flabel pwell 6876 -6013 6910 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_112/VNB
rlabel comment 6847 -5996 6847 -5996 4 sky130_fd_sc_hd__decap_8_112/decap_8
rlabel metal1 6847 -6044 7583 -5948 1 sky130_fd_sc_hd__decap_8_112/VGND
rlabel metal1 6847 -5500 7583 -5404 1 sky130_fd_sc_hd__decap_8_112/VPWR
flabel metal1 6772 -5472 6825 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_235/VPWR
flabel metal1 6775 -6014 6826 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_235/VGND
rlabel comment 6847 -5996 6847 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_235/tapvpwrvgnd_1
rlabel metal1 6755 -6044 6847 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_235/VGND
rlabel metal1 6755 -5500 6847 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_235/VPWR
flabel metal1 8060 -5472 8113 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_238/VPWR
flabel metal1 8063 -6014 8114 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_238/VGND
rlabel comment 8135 -5996 8135 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_238/tapvpwrvgnd_1
rlabel metal1 8043 -6044 8135 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_238/VGND
rlabel metal1 8043 -5500 8135 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_238/VPWR
flabel metal1 7600 -5472 7653 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_239/VPWR
flabel metal1 7603 -6014 7654 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_239/VGND
rlabel comment 7675 -5996 7675 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_239/tapvpwrvgnd_1
rlabel metal1 7583 -6044 7675 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_239/VGND
rlabel metal1 7583 -5500 7675 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_239/VPWR
flabel metal1 9268 -6013 9302 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_121/VGND
flabel metal1 9268 -5469 9302 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_121/VPWR
flabel nwell 9268 -5469 9302 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_121/VPB
flabel pwell 9268 -6013 9302 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_121/VNB
rlabel comment 9331 -5996 9331 -5996 6 sky130_fd_sc_hd__decap_4_121/decap_4
rlabel metal1 8963 -6044 9331 -5948 1 sky130_fd_sc_hd__decap_4_121/VGND
rlabel metal1 8963 -5500 9331 -5404 1 sky130_fd_sc_hd__decap_4_121/VPWR
flabel metal1 10648 -6013 10682 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_123/VGND
flabel metal1 10648 -5469 10682 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_123/VPWR
flabel nwell 10648 -5469 10682 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_123/VPB
flabel pwell 10648 -6013 10682 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_123/VNB
rlabel comment 10711 -5996 10711 -5996 6 sky130_fd_sc_hd__decap_4_123/decap_4
rlabel metal1 10343 -6044 10711 -5948 1 sky130_fd_sc_hd__decap_4_123/VGND
rlabel metal1 10343 -5500 10711 -5404 1 sky130_fd_sc_hd__decap_4_123/VPWR
flabel metal1 9452 -5469 9486 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_122/VPWR
flabel metal1 9452 -6013 9486 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_122/VGND
flabel nwell 9452 -5469 9486 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_122/VPB
flabel pwell 9452 -6013 9486 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_122/VNB
rlabel comment 9423 -5996 9423 -5996 4 sky130_fd_sc_hd__decap_8_122/decap_8
rlabel metal1 9423 -6044 10159 -5948 1 sky130_fd_sc_hd__decap_8_122/VGND
rlabel metal1 9423 -5500 10159 -5404 1 sky130_fd_sc_hd__decap_8_122/VPWR
flabel metal1 10285 -5469 10321 -5439 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_32/VPWR
flabel metal1 10285 -6009 10321 -5980 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_32/VGND
flabel nwell 10292 -5462 10312 -5445 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_32/VPB
flabel pwell 10291 -6007 10315 -5985 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_32/VNB
rlabel comment 10343 -5996 10343 -5996 6 sky130_fd_sc_hd__fill_1_32/fill_1
rlabel metal1 10251 -6044 10343 -5948 1 sky130_fd_sc_hd__fill_1_32/VGND
rlabel metal1 10251 -5500 10343 -5404 1 sky130_fd_sc_hd__fill_1_32/VPWR
flabel metal1 8888 -5472 8941 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_241/VPWR
flabel metal1 8891 -6014 8942 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_241/VGND
rlabel comment 8963 -5996 8963 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_241/tapvpwrvgnd_1
rlabel metal1 8871 -6044 8963 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_241/VGND
rlabel metal1 8871 -5500 8963 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_241/VPWR
flabel metal1 9348 -5472 9401 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_243/VPWR
flabel metal1 9351 -6014 9402 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_243/VGND
rlabel comment 9423 -5996 9423 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_243/tapvpwrvgnd_1
rlabel metal1 9331 -6044 9423 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_243/VGND
rlabel metal1 9331 -5500 9423 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_243/VPWR
flabel metal1 10176 -5472 10229 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_245/VPWR
flabel metal1 10179 -6014 10230 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_245/VGND
rlabel comment 10251 -5996 10251 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_245/tapvpwrvgnd_1
rlabel metal1 10159 -6044 10251 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_245/VGND
rlabel metal1 10159 -5500 10251 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_245/VPWR
flabel locali 11383 -5775 11417 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/A
flabel locali 10737 -5571 10771 -5537 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
flabel locali 10737 -5639 10771 -5605 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
flabel locali 10737 -5707 10771 -5673 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
flabel locali 10737 -5775 10771 -5741 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
flabel locali 10737 -5843 10771 -5809 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
flabel locali 10737 -5911 10771 -5877 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
flabel pwell 11383 -6013 11417 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/VNB
flabel nwell 11383 -5469 11417 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/VPB
flabel metal1 11383 -6013 11417 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/VGND
flabel metal1 11383 -5469 11417 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_99/VPWR
rlabel comment 11447 -5996 11447 -5996 6 sky130_fd_sc_hd__clkdlybuf4s50_1_99/clkdlybuf4s50_1
rlabel metal1 10711 -6044 11447 -5948 1 sky130_fd_sc_hd__clkdlybuf4s50_1_99/VGND
rlabel metal1 10711 -5500 11447 -5404 1 sky130_fd_sc_hd__clkdlybuf4s50_1_99/VPWR
flabel metal1 11936 -6013 11970 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_125/VGND
flabel metal1 11936 -5469 11970 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_125/VPWR
flabel nwell 11936 -5469 11970 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_125/VPB
flabel pwell 11936 -6013 11970 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_125/VNB
rlabel comment 11999 -5996 11999 -5996 6 sky130_fd_sc_hd__decap_4_125/decap_4
rlabel metal1 11631 -6044 11999 -5948 1 sky130_fd_sc_hd__decap_4_125/VGND
rlabel metal1 11631 -5500 11999 -5404 1 sky130_fd_sc_hd__decap_4_125/VPWR
flabel metal1 10653 -5469 10689 -5439 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_33/VPWR
flabel metal1 10653 -6009 10689 -5980 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_33/VGND
flabel nwell 10660 -5462 10680 -5445 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_33/VPB
flabel pwell 10659 -6007 10683 -5985 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_33/VNB
rlabel comment 10711 -5996 10711 -5996 6 sky130_fd_sc_hd__fill_1_33/fill_1
rlabel metal1 10619 -6044 10711 -5948 1 sky130_fd_sc_hd__fill_1_33/VGND
rlabel metal1 10619 -5500 10711 -5404 1 sky130_fd_sc_hd__fill_1_33/VPWR
flabel metal1 11573 -5469 11609 -5439 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_34/VPWR
flabel metal1 11573 -6009 11609 -5980 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_34/VGND
flabel nwell 11580 -5462 11600 -5445 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_34/VPB
flabel pwell 11579 -6007 11603 -5985 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_34/VNB
rlabel comment 11631 -5996 11631 -5996 6 sky130_fd_sc_hd__fill_1_34/fill_1
rlabel metal1 11539 -6044 11631 -5948 1 sky130_fd_sc_hd__fill_1_34/VGND
rlabel metal1 11539 -5500 11631 -5404 1 sky130_fd_sc_hd__fill_1_34/VPWR
flabel metal1 12668 -6016 12700 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_15/VGND
flabel metal1 12668 -5473 12706 -5441 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_15/VPWR
flabel nwell 12658 -5474 12715 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_15/VPB
flabel pwell 12665 -6020 12709 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_15/VNB
rlabel comment 12735 -5996 12735 -5996 6 sky130_fd_sc_hd__fill_8_15/fill_8
rlabel metal1 11999 -6044 12735 -5948 1 sky130_fd_sc_hd__fill_8_15/VGND
rlabel metal1 11999 -5500 12735 -5404 1 sky130_fd_sc_hd__fill_8_15/VPWR
flabel metal1 11464 -5472 11517 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_248/VPWR
flabel metal1 11467 -6014 11518 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_248/VGND
rlabel comment 11539 -5996 11539 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_248/tapvpwrvgnd_1
rlabel metal1 11447 -6044 11539 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_248/VGND
rlabel metal1 11447 -5500 11539 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_248/VPWR
flabel locali 15248 -5707 15282 -5673 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/X
flabel locali 15340 -5707 15374 -5673 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/X
flabel locali 15340 -5775 15374 -5741 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/X
flabel locali 15248 -5775 15282 -5741 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/X
flabel locali 15248 -5843 15282 -5809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/X
flabel locali 15340 -5843 15374 -5809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/X
flabel locali 13684 -5843 13718 -5809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/A
flabel locali 13684 -5775 13718 -5741 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/A
flabel pwell 13684 -6013 13718 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/VNB
flabel pwell 13701 -5996 13701 -5996 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/VNB
flabel nwell 13684 -5469 13718 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/VPB
flabel nwell 13701 -5452 13701 -5452 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/VPB
flabel metal1 13684 -6013 13718 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/VGND
flabel metal1 13684 -5469 13718 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_7/VPWR
rlabel comment 13655 -5996 13655 -5996 4 sky130_fd_sc_hd__clkbuf_16_7/clkbuf_16
rlabel metal1 13655 -6044 15495 -5948 1 sky130_fd_sc_hd__clkbuf_16_7/VGND
rlabel metal1 13655 -5500 15495 -5404 1 sky130_fd_sc_hd__clkbuf_16_7/VPWR
flabel metal1 13505 -5469 13541 -5439 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_35/VPWR
flabel metal1 13505 -6009 13541 -5980 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_35/VGND
flabel nwell 13512 -5462 13532 -5445 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_35/VPB
flabel pwell 13511 -6007 13535 -5985 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_35/VNB
rlabel comment 13563 -5996 13563 -5996 6 sky130_fd_sc_hd__fill_1_35/fill_1
rlabel metal1 13471 -6044 13563 -5948 1 sky130_fd_sc_hd__fill_1_35/VGND
rlabel metal1 13471 -5500 13563 -5404 1 sky130_fd_sc_hd__fill_1_35/VPWR
flabel metal1 13404 -6016 13436 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_16/VGND
flabel metal1 13404 -5473 13442 -5441 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_16/VPWR
flabel nwell 13394 -5474 13451 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_16/VPB
flabel pwell 13401 -6020 13445 -5986 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_16/VNB
rlabel comment 13471 -5996 13471 -5996 6 sky130_fd_sc_hd__fill_8_16/fill_8
rlabel metal1 12735 -6044 13471 -5948 1 sky130_fd_sc_hd__fill_8_16/VGND
rlabel metal1 12735 -5500 13471 -5404 1 sky130_fd_sc_hd__fill_8_16/VPWR
flabel metal1 13580 -5472 13633 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_249/VPWR
flabel metal1 13583 -6014 13634 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_249/VGND
rlabel comment 13655 -5996 13655 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_249/tapvpwrvgnd_1
rlabel metal1 13563 -6044 13655 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_249/VGND
rlabel metal1 13563 -5500 13655 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_249/VPWR
flabel metal1 16628 -6013 16662 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_17/VGND
flabel metal1 16628 -5469 16662 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_17/VPWR
flabel nwell 16628 -5469 16662 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_17/VPB
flabel pwell 16628 -6013 16662 -5979 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_17/VNB
rlabel comment 16691 -5996 16691 -5996 6 sky130_fd_sc_hd__decap_12_17/decap_12
rlabel metal1 15587 -6044 16691 -5948 1 sky130_fd_sc_hd__decap_12_17/VGND
rlabel metal1 15587 -5500 16691 -5404 1 sky130_fd_sc_hd__decap_12_17/VPWR
flabel metal1 15512 -5472 15565 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_252/VPWR
flabel metal1 15515 -6014 15566 -5976 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_252/VGND
rlabel comment 15587 -5996 15587 -5996 6 sky130_fd_sc_hd__tapvpwrvgnd_1_252/tapvpwrvgnd_1
rlabel metal1 15495 -6044 15587 -5948 1 sky130_fd_sc_hd__tapvpwrvgnd_1_252/VGND
rlabel metal1 15495 -5500 15587 -5404 1 sky130_fd_sc_hd__tapvpwrvgnd_1_252/VPWR
flabel metal1 -1588 -5469 -1554 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_17/VPWR
flabel metal1 -1588 -4925 -1554 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_17/VGND
flabel nwell -1588 -5469 -1554 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_17/VPB
flabel pwell -1588 -4925 -1554 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_17/VNB
rlabel comment -1617 -4908 -1617 -4908 2 sky130_fd_sc_hd__decap_8_17/decap_8
rlabel metal1 -1617 -4956 -881 -4860 5 sky130_fd_sc_hd__decap_8_17/VGND
rlabel metal1 -1617 -5500 -881 -5404 5 sky130_fd_sc_hd__decap_8_17/VPWR
flabel metal1 -2324 -5469 -2290 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_74/VPWR
flabel metal1 -2324 -4925 -2290 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_74/VGND
flabel nwell -2324 -5469 -2290 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_74/VPB
flabel pwell -2324 -4925 -2290 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_74/VNB
rlabel comment -2261 -4908 -2261 -4908 8 sky130_fd_sc_hd__decap_8_74/decap_8
rlabel metal1 -2997 -4956 -2261 -4860 5 sky130_fd_sc_hd__decap_8_74/VGND
rlabel metal1 -2997 -5500 -2261 -5404 5 sky130_fd_sc_hd__decap_8_74/VPWR
flabel metal1 -1690 -4926 -1637 -4894 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_11/VGND
flabel metal1 -1690 -5469 -1638 -5438 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_11/VPWR
flabel nwell -1679 -5461 -1645 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_11/VPB
flabel pwell -1680 -4920 -1648 -4898 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_11/VNB
rlabel comment -1617 -4908 -1617 -4908 8 sky130_fd_sc_hd__fill_2_11/fill_2
rlabel metal1 -1801 -4956 -1617 -4860 5 sky130_fd_sc_hd__fill_2_11/VGND
rlabel metal1 -1801 -5500 -1617 -5404 5 sky130_fd_sc_hd__fill_2_11/VPWR
flabel metal1 -1858 -4917 -1835 -4898 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_24/VGND
flabel metal1 -1855 -5460 -1835 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_24/VPWR
flabel nwell -1861 -5464 -1836 -5438 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_24/VPB
flabel pwell -1858 -4920 -1836 -4896 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_24/VNB
rlabel comment -1801 -4908 -1801 -4908 8 sky130_fd_sc_hd__fill_4_24/fill_4
rlabel metal1 -2169 -4956 -1801 -4860 5 sky130_fd_sc_hd__fill_4_24/VGND
rlabel metal1 -2169 -5500 -1801 -5404 5 sky130_fd_sc_hd__fill_4_24/VPWR
flabel metal1 -2244 -5461 -2191 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_539/VPWR
flabel metal1 -2241 -4928 -2190 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_539/VGND
rlabel comment -2169 -4908 -2169 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_539/tapvpwrvgnd_1
rlabel metal1 -2261 -4956 -2169 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_539/VGND
rlabel metal1 -2261 -5500 -2169 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_539/VPWR
flabel locali 437 -5163 471 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/A
flabel locali 1083 -5367 1117 -5333 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/X
flabel locali 1083 -5299 1117 -5265 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/X
flabel locali 1083 -5231 1117 -5197 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/X
flabel locali 1083 -5163 1117 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/X
flabel locali 1083 -5095 1117 -5061 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/X
flabel locali 1083 -5027 1117 -4993 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/X
flabel pwell 437 -4925 471 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/VNB
flabel nwell 437 -5469 471 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/VPB
flabel metal1 437 -4925 471 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/VGND
flabel metal1 437 -5469 471 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_78/VPWR
rlabel comment 407 -4908 407 -4908 2 sky130_fd_sc_hd__clkdlybuf4s50_1_78/clkdlybuf4s50_1
rlabel metal1 407 -4956 1143 -4860 5 sky130_fd_sc_hd__clkdlybuf4s50_1_78/VGND
rlabel metal1 407 -5500 1143 -5404 5 sky130_fd_sc_hd__clkdlybuf4s50_1_78/VPWR
flabel metal1 252 -4925 286 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_94/VGND
flabel metal1 252 -5469 286 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_94/VPWR
flabel nwell 252 -5469 286 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_94/VPB
flabel pwell 252 -4925 286 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_94/VNB
rlabel comment 315 -4908 315 -4908 8 sky130_fd_sc_hd__decap_4_94/decap_4
rlabel metal1 -53 -4956 315 -4860 5 sky130_fd_sc_hd__decap_4_94/VGND
rlabel metal1 -53 -5500 315 -5404 5 sky130_fd_sc_hd__decap_4_94/VPWR
flabel metal1 -852 -5469 -818 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_18/VPWR
flabel metal1 -852 -4925 -818 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_18/VGND
flabel nwell -852 -5469 -818 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_18/VPB
flabel pwell -852 -4925 -818 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_18/VNB
rlabel comment -881 -4908 -881 -4908 2 sky130_fd_sc_hd__decap_8_18/decap_8
rlabel metal1 -881 -4956 -145 -4860 5 sky130_fd_sc_hd__decap_8_18/VGND
rlabel metal1 -881 -5500 -145 -5404 5 sky130_fd_sc_hd__decap_8_18/VPWR
flabel metal1 -128 -5461 -75 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_190/VPWR
flabel metal1 -125 -4928 -74 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_190/VGND
rlabel comment -53 -4908 -53 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_190/tapvpwrvgnd_1
rlabel metal1 -145 -4956 -53 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_190/VGND
rlabel metal1 -145 -5500 -53 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_190/VPWR
flabel metal1 332 -5461 385 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_191/VPWR
flabel metal1 335 -4928 386 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_191/VGND
rlabel comment 407 -4908 407 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_191/tapvpwrvgnd_1
rlabel metal1 315 -4956 407 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_191/VGND
rlabel metal1 315 -5500 407 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_191/VPWR
flabel metal1 1540 -4925 1574 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_95/VGND
flabel metal1 1540 -5469 1574 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_95/VPWR
flabel nwell 1540 -5469 1574 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_95/VPB
flabel pwell 1540 -4925 1574 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_95/VNB
rlabel comment 1603 -4908 1603 -4908 8 sky130_fd_sc_hd__decap_4_95/decap_4
rlabel metal1 1235 -4956 1603 -4860 5 sky130_fd_sc_hd__decap_4_95/VGND
rlabel metal1 1235 -5500 1603 -5404 5 sky130_fd_sc_hd__decap_4_95/VPWR
flabel metal1 2828 -4925 2862 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_96/VGND
flabel metal1 2828 -5469 2862 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_96/VPWR
flabel nwell 2828 -5469 2862 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_96/VPB
flabel pwell 2828 -4925 2862 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_96/VNB
rlabel comment 2891 -4908 2891 -4908 8 sky130_fd_sc_hd__decap_4_96/decap_4
rlabel metal1 2523 -4956 2891 -4860 5 sky130_fd_sc_hd__decap_4_96/VGND
rlabel metal1 2523 -5500 2891 -5404 5 sky130_fd_sc_hd__decap_4_96/VPWR
flabel metal1 2368 -5469 2402 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_99/VPWR
flabel metal1 2368 -4925 2402 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_99/VGND
flabel nwell 2368 -5469 2402 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_99/VPB
flabel pwell 2368 -4925 2402 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_99/VNB
rlabel comment 2431 -4908 2431 -4908 8 sky130_fd_sc_hd__decap_8_99/decap_8
rlabel metal1 1695 -4956 2431 -4860 5 sky130_fd_sc_hd__decap_8_99/VGND
rlabel metal1 1695 -5500 2431 -5404 5 sky130_fd_sc_hd__decap_8_99/VPWR
flabel metal1 1160 -5461 1213 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_192/VPWR
flabel metal1 1163 -4928 1214 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_192/VGND
rlabel comment 1235 -4908 1235 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_192/tapvpwrvgnd_1
rlabel metal1 1143 -4956 1235 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_192/VGND
rlabel metal1 1143 -5500 1235 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_192/VPWR
flabel metal1 1620 -5461 1673 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_193/VPWR
flabel metal1 1623 -4928 1674 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_193/VGND
rlabel comment 1695 -4908 1695 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_193/tapvpwrvgnd_1
rlabel metal1 1603 -4956 1695 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_193/VGND
rlabel metal1 1603 -5500 1695 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_193/VPWR
flabel metal1 2448 -5461 2501 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_194/VPWR
flabel metal1 2451 -4928 2502 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_194/VGND
rlabel comment 2523 -4908 2523 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_194/tapvpwrvgnd_1
rlabel metal1 2431 -4956 2523 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_194/VGND
rlabel metal1 2431 -5500 2523 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_194/VPWR
flabel locali 3013 -5163 3047 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A
flabel locali 3659 -5367 3693 -5333 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/X
flabel locali 3659 -5299 3693 -5265 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/X
flabel locali 3659 -5231 3693 -5197 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/X
flabel locali 3659 -5163 3693 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/X
flabel locali 3659 -5095 3693 -5061 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/X
flabel locali 3659 -5027 3693 -4993 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/X
flabel pwell 3013 -4925 3047 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/VNB
flabel nwell 3013 -5469 3047 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/VPB
flabel metal1 3013 -4925 3047 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/VGND
flabel metal1 3013 -5469 3047 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_80/VPWR
rlabel comment 2983 -4908 2983 -4908 2 sky130_fd_sc_hd__clkdlybuf4s50_1_80/clkdlybuf4s50_1
rlabel metal1 2983 -4956 3719 -4860 5 sky130_fd_sc_hd__clkdlybuf4s50_1_80/VGND
rlabel metal1 2983 -5500 3719 -5404 5 sky130_fd_sc_hd__clkdlybuf4s50_1_80/VPWR
flabel metal1 4116 -4925 4150 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_97/VGND
flabel metal1 4116 -5469 4150 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_97/VPWR
flabel nwell 4116 -5469 4150 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_97/VPB
flabel pwell 4116 -4925 4150 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_97/VNB
rlabel comment 4179 -4908 4179 -4908 8 sky130_fd_sc_hd__decap_4_97/decap_4
rlabel metal1 3811 -4956 4179 -4860 5 sky130_fd_sc_hd__decap_4_97/VGND
rlabel metal1 3811 -5500 4179 -5404 5 sky130_fd_sc_hd__decap_4_97/VPWR
flabel metal1 4944 -5469 4978 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_103/VPWR
flabel metal1 4944 -4925 4978 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_103/VGND
flabel nwell 4944 -5469 4978 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_103/VPB
flabel pwell 4944 -4925 4978 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_103/VNB
rlabel comment 5007 -4908 5007 -4908 8 sky130_fd_sc_hd__decap_8_103/decap_8
rlabel metal1 4271 -4956 5007 -4860 5 sky130_fd_sc_hd__decap_8_103/VGND
rlabel metal1 4271 -5500 5007 -5404 5 sky130_fd_sc_hd__decap_8_103/VPWR
flabel metal1 3736 -5461 3789 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_195/VPWR
flabel metal1 3739 -4928 3790 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_195/VGND
rlabel comment 3811 -4908 3811 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_195/tapvpwrvgnd_1
rlabel metal1 3719 -4956 3811 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_195/VGND
rlabel metal1 3719 -5500 3811 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_195/VPWR
flabel metal1 2908 -5461 2961 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_196/VPWR
flabel metal1 2911 -4928 2962 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_196/VGND
rlabel comment 2983 -4908 2983 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_196/tapvpwrvgnd_1
rlabel metal1 2891 -4956 2983 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_196/VGND
rlabel metal1 2891 -5500 2983 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_196/VPWR
flabel metal1 4196 -5461 4249 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_197/VPWR
flabel metal1 4199 -4928 4250 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_197/VGND
rlabel comment 4271 -4908 4271 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_197/tapvpwrvgnd_1
rlabel metal1 4179 -4956 4271 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_197/VGND
rlabel metal1 4179 -5500 4271 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_197/VPWR
flabel locali 5589 -5163 5623 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A
flabel locali 6235 -5367 6269 -5333 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/X
flabel locali 6235 -5299 6269 -5265 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/X
flabel locali 6235 -5231 6269 -5197 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/X
flabel locali 6235 -5163 6269 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/X
flabel locali 6235 -5095 6269 -5061 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/X
flabel locali 6235 -5027 6269 -4993 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/X
flabel pwell 5589 -4925 5623 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/VNB
flabel nwell 5589 -5469 5623 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/VPB
flabel metal1 5589 -4925 5623 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/VGND
flabel metal1 5589 -5469 5623 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_82/VPWR
rlabel comment 5559 -4908 5559 -4908 2 sky130_fd_sc_hd__clkdlybuf4s50_1_82/clkdlybuf4s50_1
rlabel metal1 5559 -4956 6295 -4860 5 sky130_fd_sc_hd__clkdlybuf4s50_1_82/VGND
rlabel metal1 5559 -5500 6295 -5404 5 sky130_fd_sc_hd__clkdlybuf4s50_1_82/VPWR
flabel metal1 5404 -4925 5438 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_98/VGND
flabel metal1 5404 -5469 5438 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_98/VPWR
flabel nwell 5404 -5469 5438 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_98/VPB
flabel pwell 5404 -4925 5438 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_98/VNB
rlabel comment 5467 -4908 5467 -4908 8 sky130_fd_sc_hd__decap_4_98/decap_4
rlabel metal1 5099 -4956 5467 -4860 5 sky130_fd_sc_hd__decap_4_98/VGND
rlabel metal1 5099 -5500 5467 -5404 5 sky130_fd_sc_hd__decap_4_98/VPWR
flabel metal1 6692 -4925 6726 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_99/VGND
flabel metal1 6692 -5469 6726 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_99/VPWR
flabel nwell 6692 -5469 6726 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_99/VPB
flabel pwell 6692 -4925 6726 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_99/VNB
rlabel comment 6755 -4908 6755 -4908 8 sky130_fd_sc_hd__decap_4_99/decap_4
rlabel metal1 6387 -4956 6755 -4860 5 sky130_fd_sc_hd__decap_4_99/VGND
rlabel metal1 6387 -5500 6755 -5404 5 sky130_fd_sc_hd__decap_4_99/VPWR
flabel metal1 5024 -5461 5077 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_198/VPWR
flabel metal1 5027 -4928 5078 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_198/VGND
rlabel comment 5099 -4908 5099 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_198/tapvpwrvgnd_1
rlabel metal1 5007 -4956 5099 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_198/VGND
rlabel metal1 5007 -5500 5099 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_198/VPWR
flabel metal1 5484 -5461 5537 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_199/VPWR
flabel metal1 5487 -4928 5538 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_199/VGND
rlabel comment 5559 -4908 5559 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_199/tapvpwrvgnd_1
rlabel metal1 5467 -4956 5559 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_199/VGND
rlabel metal1 5467 -5500 5559 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_199/VPWR
flabel metal1 6312 -5461 6365 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_200/VPWR
flabel metal1 6315 -4928 6366 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_200/VGND
rlabel comment 6387 -4908 6387 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_200/tapvpwrvgnd_1
rlabel metal1 6295 -4956 6387 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_200/VGND
rlabel metal1 6295 -5500 6387 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_200/VPWR
flabel locali 8165 -5163 8199 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A
flabel locali 8811 -5367 8845 -5333 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/X
flabel locali 8811 -5299 8845 -5265 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/X
flabel locali 8811 -5231 8845 -5197 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/X
flabel locali 8811 -5163 8845 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/X
flabel locali 8811 -5095 8845 -5061 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/X
flabel locali 8811 -5027 8845 -4993 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/X
flabel pwell 8165 -4925 8199 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/VNB
flabel nwell 8165 -5469 8199 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/VPB
flabel metal1 8165 -4925 8199 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/VGND
flabel metal1 8165 -5469 8199 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_84/VPWR
rlabel comment 8135 -4908 8135 -4908 2 sky130_fd_sc_hd__clkdlybuf4s50_1_84/clkdlybuf4s50_1
rlabel metal1 8135 -4956 8871 -4860 5 sky130_fd_sc_hd__clkdlybuf4s50_1_84/VGND
rlabel metal1 8135 -5500 8871 -5404 5 sky130_fd_sc_hd__clkdlybuf4s50_1_84/VPWR
flabel metal1 7980 -4925 8014 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_100/VGND
flabel metal1 7980 -5469 8014 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_100/VPWR
flabel nwell 7980 -5469 8014 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_100/VPB
flabel pwell 7980 -4925 8014 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_100/VNB
rlabel comment 8043 -4908 8043 -4908 8 sky130_fd_sc_hd__decap_4_100/decap_4
rlabel metal1 7675 -4956 8043 -4860 5 sky130_fd_sc_hd__decap_4_100/VGND
rlabel metal1 7675 -5500 8043 -5404 5 sky130_fd_sc_hd__decap_4_100/VPWR
flabel metal1 7520 -5469 7554 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_111/VPWR
flabel metal1 7520 -4925 7554 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_111/VGND
flabel nwell 7520 -5469 7554 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_111/VPB
flabel pwell 7520 -4925 7554 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_111/VNB
rlabel comment 7583 -4908 7583 -4908 8 sky130_fd_sc_hd__decap_8_111/decap_8
rlabel metal1 6847 -4956 7583 -4860 5 sky130_fd_sc_hd__decap_8_111/VGND
rlabel metal1 6847 -5500 7583 -5404 5 sky130_fd_sc_hd__decap_8_111/VPWR
flabel metal1 6772 -5461 6825 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_201/VPWR
flabel metal1 6775 -4928 6826 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_201/VGND
rlabel comment 6847 -4908 6847 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_201/tapvpwrvgnd_1
rlabel metal1 6755 -4956 6847 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_201/VGND
rlabel metal1 6755 -5500 6847 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_201/VPWR
flabel metal1 7600 -5461 7653 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_202/VPWR
flabel metal1 7603 -4928 7654 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_202/VGND
rlabel comment 7675 -4908 7675 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_202/tapvpwrvgnd_1
rlabel metal1 7583 -4956 7675 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_202/VGND
rlabel metal1 7583 -5500 7675 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_202/VPWR
flabel metal1 8060 -5461 8113 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_203/VPWR
flabel metal1 8063 -4928 8114 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_203/VGND
rlabel comment 8135 -4908 8135 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_203/tapvpwrvgnd_1
rlabel metal1 8043 -4956 8135 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_203/VGND
rlabel metal1 8043 -5500 8135 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_203/VPWR
flabel metal1 9268 -4925 9302 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_101/VGND
flabel metal1 9268 -5469 9302 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_101/VPWR
flabel nwell 9268 -5469 9302 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_101/VPB
flabel pwell 9268 -4925 9302 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_101/VNB
rlabel comment 9331 -4908 9331 -4908 8 sky130_fd_sc_hd__decap_4_101/decap_4
rlabel metal1 8963 -4956 9331 -4860 5 sky130_fd_sc_hd__decap_4_101/VGND
rlabel metal1 8963 -5500 9331 -5404 5 sky130_fd_sc_hd__decap_4_101/VPWR
flabel metal1 10648 -4925 10682 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_102/VGND
flabel metal1 10648 -5469 10682 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_102/VPWR
flabel nwell 10648 -5469 10682 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_102/VPB
flabel pwell 10648 -4925 10682 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_102/VNB
rlabel comment 10711 -4908 10711 -4908 8 sky130_fd_sc_hd__decap_4_102/decap_4
rlabel metal1 10343 -4956 10711 -4860 5 sky130_fd_sc_hd__decap_4_102/VGND
rlabel metal1 10343 -5500 10711 -5404 5 sky130_fd_sc_hd__decap_4_102/VPWR
flabel metal1 10096 -5469 10130 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_121/VPWR
flabel metal1 10096 -4925 10130 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_121/VGND
flabel nwell 10096 -5469 10130 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_121/VPB
flabel pwell 10096 -4925 10130 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_121/VNB
rlabel comment 10159 -4908 10159 -4908 8 sky130_fd_sc_hd__decap_8_121/decap_8
rlabel metal1 9423 -4956 10159 -4860 5 sky130_fd_sc_hd__decap_8_121/VGND
rlabel metal1 9423 -5500 10159 -5404 5 sky130_fd_sc_hd__decap_8_121/VPWR
flabel metal1 10285 -5465 10321 -5435 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_28/VPWR
flabel metal1 10285 -4924 10321 -4895 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_28/VGND
flabel nwell 10292 -5459 10312 -5442 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_28/VPB
flabel pwell 10291 -4919 10315 -4897 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_28/VNB
rlabel comment 10343 -4908 10343 -4908 8 sky130_fd_sc_hd__fill_1_28/fill_1
rlabel metal1 10251 -4956 10343 -4860 5 sky130_fd_sc_hd__fill_1_28/VGND
rlabel metal1 10251 -5500 10343 -5404 5 sky130_fd_sc_hd__fill_1_28/VPWR
flabel metal1 9348 -5461 9401 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_204/VPWR
flabel metal1 9351 -4928 9402 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_204/VGND
rlabel comment 9423 -4908 9423 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_204/tapvpwrvgnd_1
rlabel metal1 9331 -4956 9423 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_204/VGND
rlabel metal1 9331 -5500 9423 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_204/VPWR
flabel metal1 8888 -5461 8941 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_205/VPWR
flabel metal1 8891 -4928 8942 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_205/VGND
rlabel comment 8963 -4908 8963 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_205/tapvpwrvgnd_1
rlabel metal1 8871 -4956 8963 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_205/VGND
rlabel metal1 8871 -5500 8963 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_205/VPWR
flabel metal1 10176 -5461 10229 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_206/VPWR
flabel metal1 10179 -4928 10230 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_206/VGND
rlabel comment 10251 -4908 10251 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_206/tapvpwrvgnd_1
rlabel metal1 10159 -4956 10251 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_206/VGND
rlabel metal1 10159 -5500 10251 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_206/VPWR
flabel locali 10741 -5163 10775 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A
flabel locali 11387 -5367 11421 -5333 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
flabel locali 11387 -5299 11421 -5265 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
flabel locali 11387 -5231 11421 -5197 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
flabel locali 11387 -5163 11421 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
flabel locali 11387 -5095 11421 -5061 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
flabel locali 11387 -5027 11421 -4993 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
flabel pwell 10741 -4925 10775 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/VNB
flabel nwell 10741 -5469 10775 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/VPB
flabel metal1 10741 -4925 10775 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/VGND
flabel metal1 10741 -5469 10775 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_86/VPWR
rlabel comment 10711 -4908 10711 -4908 2 sky130_fd_sc_hd__clkdlybuf4s50_1_86/clkdlybuf4s50_1
rlabel metal1 10711 -4956 11447 -4860 5 sky130_fd_sc_hd__clkdlybuf4s50_1_86/VGND
rlabel metal1 10711 -5500 11447 -5404 5 sky130_fd_sc_hd__clkdlybuf4s50_1_86/VPWR
flabel metal1 11936 -4925 11970 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_103/VGND
flabel metal1 11936 -5469 11970 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_103/VPWR
flabel nwell 11936 -5469 11970 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_103/VPB
flabel pwell 11936 -4925 11970 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_103/VNB
rlabel comment 11999 -4908 11999 -4908 8 sky130_fd_sc_hd__decap_4_103/decap_4
rlabel metal1 11631 -4956 11999 -4860 5 sky130_fd_sc_hd__decap_4_103/VGND
rlabel metal1 11631 -5500 11999 -5404 5 sky130_fd_sc_hd__decap_4_103/VPWR
flabel metal1 10653 -5465 10689 -5435 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_29/VPWR
flabel metal1 10653 -4924 10689 -4895 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_29/VGND
flabel nwell 10660 -5459 10680 -5442 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_29/VPB
flabel pwell 10659 -4919 10683 -4897 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_29/VNB
rlabel comment 10711 -4908 10711 -4908 8 sky130_fd_sc_hd__fill_1_29/fill_1
rlabel metal1 10619 -4956 10711 -4860 5 sky130_fd_sc_hd__fill_1_29/VGND
rlabel metal1 10619 -5500 10711 -5404 5 sky130_fd_sc_hd__fill_1_29/VPWR
flabel metal1 11573 -5465 11609 -5435 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_30/VPWR
flabel metal1 11573 -4924 11609 -4895 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_30/VGND
flabel nwell 11580 -5459 11600 -5442 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_30/VPB
flabel pwell 11579 -4919 11603 -4897 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_30/VNB
rlabel comment 11631 -4908 11631 -4908 8 sky130_fd_sc_hd__fill_1_30/fill_1
rlabel metal1 11539 -4956 11631 -4860 5 sky130_fd_sc_hd__fill_1_30/VGND
rlabel metal1 11539 -5500 11631 -5404 5 sky130_fd_sc_hd__fill_1_30/VPWR
flabel metal1 12033 -4917 12056 -4898 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_5/VGND
flabel metal1 12033 -5460 12053 -5443 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_5/VPWR
flabel nwell 12034 -5464 12059 -5438 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_5/VPB
flabel pwell 12034 -4920 12056 -4896 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_5/VNB
rlabel comment 11999 -4908 11999 -4908 2 sky130_fd_sc_hd__fill_4_5/fill_4
rlabel metal1 11999 -4956 12367 -4860 5 sky130_fd_sc_hd__fill_4_5/VGND
rlabel metal1 11999 -5500 12367 -5404 5 sky130_fd_sc_hd__fill_4_5/VPWR
flabel metal1 11464 -5461 11517 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_207/VPWR
flabel metal1 11467 -4928 11518 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_207/VGND
rlabel comment 11539 -4908 11539 -4908 8 sky130_fd_sc_hd__tapvpwrvgnd_1_207/tapvpwrvgnd_1
rlabel metal1 11447 -4956 11539 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_207/VGND
rlabel metal1 11447 -5500 11539 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_207/VPWR
flabel locali 15248 -5231 15282 -5197 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/X
flabel locali 15340 -5231 15374 -5197 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/X
flabel locali 15340 -5163 15374 -5129 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/X
flabel locali 15248 -5163 15282 -5129 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/X
flabel locali 15248 -5095 15282 -5061 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/X
flabel locali 15340 -5095 15374 -5061 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/X
flabel locali 13684 -5095 13718 -5061 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/A
flabel locali 13684 -5163 13718 -5129 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/A
flabel pwell 13684 -4925 13718 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/VNB
flabel pwell 13701 -4908 13701 -4908 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/VNB
flabel nwell 13684 -5469 13718 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/VPB
flabel nwell 13701 -5452 13701 -5452 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/VPB
flabel metal1 13684 -4925 13718 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/VGND
flabel metal1 13684 -5469 13718 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_6/VPWR
rlabel comment 13655 -4908 13655 -4908 2 sky130_fd_sc_hd__clkbuf_16_6/clkbuf_16
rlabel metal1 13655 -4956 15495 -4860 5 sky130_fd_sc_hd__clkbuf_16_6/VGND
rlabel metal1 13655 -5500 15495 -5404 5 sky130_fd_sc_hd__clkbuf_16_6/VPWR
flabel locali 12672 -5163 12706 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/A
flabel locali 12764 -5163 12798 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/A
flabel locali 13040 -5095 13074 -5061 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/Y
flabel locali 12580 -5163 12614 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/A
flabel locali 13040 -5231 13074 -5197 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/Y
flabel locali 12948 -5163 12982 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/A
flabel locali 12856 -5163 12890 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/A
flabel locali 13040 -5163 13074 -5129 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_4/Y
flabel pwell 12488 -4925 12522 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_4/VNB
flabel nwell 12488 -5469 12522 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_4/VPB
flabel metal1 12488 -5469 12522 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_4/VPWR
flabel metal1 12488 -4925 12522 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_4/VGND
rlabel comment 12459 -4908 12459 -4908 2 sky130_fd_sc_hd__clkinv_4_4/clkinv_4
rlabel metal1 12459 -4956 13103 -4860 5 sky130_fd_sc_hd__clkinv_4_4/VGND
rlabel metal1 12459 -5500 13103 -5404 5 sky130_fd_sc_hd__clkinv_4_4/VPWR
flabel metal1 13224 -4925 13258 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_104/VGND
flabel metal1 13224 -5469 13258 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_104/VPWR
flabel nwell 13224 -5469 13258 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_104/VPB
flabel pwell 13224 -4925 13258 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_104/VNB
rlabel comment 13195 -4908 13195 -4908 2 sky130_fd_sc_hd__decap_4_104/decap_4
rlabel metal1 13195 -4956 13563 -4860 5 sky130_fd_sc_hd__decap_4_104/VGND
rlabel metal1 13195 -5500 13563 -5404 5 sky130_fd_sc_hd__decap_4_104/VPWR
flabel metal1 12389 -5461 12442 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_208/VPWR
flabel metal1 12388 -4928 12439 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_208/VGND
rlabel comment 12367 -4908 12367 -4908 2 sky130_fd_sc_hd__tapvpwrvgnd_1_208/tapvpwrvgnd_1
rlabel metal1 12367 -4956 12459 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_208/VGND
rlabel metal1 12367 -5500 12459 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_208/VPWR
flabel metal1 13585 -5461 13638 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_209/VPWR
flabel metal1 13584 -4928 13635 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_209/VGND
rlabel comment 13563 -4908 13563 -4908 2 sky130_fd_sc_hd__tapvpwrvgnd_1_209/tapvpwrvgnd_1
rlabel metal1 13563 -4956 13655 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_209/VGND
rlabel metal1 13563 -5500 13655 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_209/VPWR
flabel metal1 13125 -5461 13178 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_210/VPWR
flabel metal1 13124 -4928 13175 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_210/VGND
rlabel comment 13103 -4908 13103 -4908 2 sky130_fd_sc_hd__tapvpwrvgnd_1_210/tapvpwrvgnd_1
rlabel metal1 13103 -4956 13195 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_210/VGND
rlabel metal1 13103 -5500 13195 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_210/VPWR
flabel metal1 15616 -4925 15650 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_13/VGND
flabel metal1 15616 -5469 15650 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_13/VPWR
flabel nwell 15616 -5469 15650 -5435 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_13/VPB
flabel pwell 15616 -4925 15650 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_13/VNB
rlabel comment 15587 -4908 15587 -4908 2 sky130_fd_sc_hd__decap_12_13/decap_12
rlabel metal1 15587 -4956 16691 -4860 5 sky130_fd_sc_hd__decap_12_13/VGND
rlabel metal1 15587 -5500 16691 -5404 5 sky130_fd_sc_hd__decap_12_13/VPWR
flabel metal1 15517 -5461 15570 -5432 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_211/VPWR
flabel metal1 15516 -4928 15567 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_211/VGND
rlabel comment 15495 -4908 15495 -4908 2 sky130_fd_sc_hd__tapvpwrvgnd_1_211/tapvpwrvgnd_1
rlabel metal1 15495 -4956 15587 -4860 5 sky130_fd_sc_hd__tapvpwrvgnd_1_211/VGND
rlabel metal1 15495 -5500 15587 -5404 5 sky130_fd_sc_hd__tapvpwrvgnd_1_211/VPWR
flabel metal1 -944 -4381 -910 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_16/VPWR
flabel metal1 -944 -4925 -910 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_16/VGND
flabel nwell -944 -4381 -910 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_16/VPB
flabel pwell -944 -4925 -910 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_16/VNB
rlabel comment -881 -4908 -881 -4908 6 sky130_fd_sc_hd__decap_8_16/decap_8
rlabel metal1 -1617 -4956 -881 -4860 1 sky130_fd_sc_hd__decap_8_16/VGND
rlabel metal1 -1617 -4412 -881 -4316 1 sky130_fd_sc_hd__decap_8_16/VPWR
flabel metal1 -2968 -4381 -2934 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_75/VPWR
flabel metal1 -2968 -4925 -2934 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_75/VGND
flabel nwell -2968 -4381 -2934 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_75/VPB
flabel pwell -2968 -4925 -2934 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_75/VNB
rlabel comment -2997 -4908 -2997 -4908 4 sky130_fd_sc_hd__decap_8_75/decap_8
rlabel metal1 -2997 -4956 -2261 -4860 1 sky130_fd_sc_hd__decap_8_75/VGND
rlabel metal1 -2997 -4412 -2261 -4316 1 sky130_fd_sc_hd__decap_8_75/VPWR
flabel metal1 -1781 -4922 -1728 -4890 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_12/VGND
flabel metal1 -1780 -4378 -1728 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_12/VPWR
flabel nwell -1773 -4373 -1739 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_12/VPB
flabel pwell -1770 -4918 -1738 -4896 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_12/VNB
rlabel comment -1801 -4908 -1801 -4908 4 sky130_fd_sc_hd__fill_2_12/fill_2
rlabel metal1 -1801 -4956 -1617 -4860 1 sky130_fd_sc_hd__fill_2_12/VGND
rlabel metal1 -1801 -4412 -1617 -4316 1 sky130_fd_sc_hd__fill_2_12/VPWR
flabel metal1 -2135 -4918 -2112 -4899 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_25/VGND
flabel metal1 -2135 -4373 -2115 -4356 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_25/VPWR
flabel nwell -2134 -4378 -2109 -4352 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_25/VPB
flabel pwell -2134 -4920 -2112 -4896 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_25/VNB
rlabel comment -2169 -4908 -2169 -4908 4 sky130_fd_sc_hd__fill_4_25/fill_4
rlabel metal1 -2169 -4956 -1801 -4860 1 sky130_fd_sc_hd__fill_4_25/VGND
rlabel metal1 -2169 -4412 -1801 -4316 1 sky130_fd_sc_hd__fill_4_25/VPWR
flabel metal1 -2239 -4384 -2186 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_540/VPWR
flabel metal1 -2240 -4926 -2189 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_540/VGND
rlabel comment -2261 -4908 -2261 -4908 4 sky130_fd_sc_hd__tapvpwrvgnd_1_540/tapvpwrvgnd_1
rlabel metal1 -2261 -4956 -2169 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_540/VGND
rlabel metal1 -2261 -4412 -2169 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_540/VPWR
flabel locali -209 -4687 -175 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A
flabel locali -855 -4483 -821 -4449 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/X
flabel locali -855 -4551 -821 -4517 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/X
flabel locali -855 -4619 -821 -4585 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/X
flabel locali -855 -4687 -821 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/X
flabel locali -855 -4755 -821 -4721 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/X
flabel locali -855 -4823 -821 -4789 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/X
flabel pwell -209 -4925 -175 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/VNB
flabel nwell -209 -4381 -175 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/VPB
flabel metal1 -209 -4925 -175 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/VGND
flabel metal1 -209 -4381 -175 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_68/VPWR
rlabel comment -145 -4908 -145 -4908 6 sky130_fd_sc_hd__clkdlybuf4s50_1_68/clkdlybuf4s50_1
rlabel metal1 -881 -4956 -145 -4860 1 sky130_fd_sc_hd__clkdlybuf4s50_1_68/VGND
rlabel metal1 -881 -4412 -145 -4316 1 sky130_fd_sc_hd__clkdlybuf4s50_1_68/VPWR
flabel locali 1079 -4687 1113 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/A
flabel locali 433 -4483 467 -4449 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X
flabel locali 433 -4551 467 -4517 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X
flabel locali 433 -4619 467 -4585 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X
flabel locali 433 -4687 467 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X
flabel locali 433 -4755 467 -4721 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X
flabel locali 433 -4823 467 -4789 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X
flabel pwell 1079 -4925 1113 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/VNB
flabel nwell 1079 -4381 1113 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/VPB
flabel metal1 1079 -4925 1113 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/VGND
flabel metal1 1079 -4381 1113 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_69/VPWR
rlabel comment 1143 -4908 1143 -4908 6 sky130_fd_sc_hd__clkdlybuf4s50_1_69/clkdlybuf4s50_1
rlabel metal1 407 -4956 1143 -4860 1 sky130_fd_sc_hd__clkdlybuf4s50_1_69/VGND
rlabel metal1 407 -4412 1143 -4316 1 sky130_fd_sc_hd__clkdlybuf4s50_1_69/VPWR
flabel metal1 252 -4925 286 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_84/VGND
flabel metal1 252 -4381 286 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_84/VPWR
flabel nwell 252 -4381 286 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_84/VPB
flabel pwell 252 -4925 286 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_84/VNB
rlabel comment 315 -4908 315 -4908 6 sky130_fd_sc_hd__decap_4_84/decap_4
rlabel metal1 -53 -4956 315 -4860 1 sky130_fd_sc_hd__decap_4_84/VGND
rlabel metal1 -53 -4412 315 -4316 1 sky130_fd_sc_hd__decap_4_84/VPWR
flabel metal1 -128 -4384 -75 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_170/VPWR
flabel metal1 -125 -4926 -74 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_170/VGND
rlabel comment -53 -4908 -53 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_170/tapvpwrvgnd_1
rlabel metal1 -145 -4956 -53 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_170/VGND
rlabel metal1 -145 -4412 -53 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_170/VPWR
flabel metal1 332 -4384 385 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_171/VPWR
flabel metal1 335 -4926 386 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_171/VGND
rlabel comment 407 -4908 407 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_171/tapvpwrvgnd_1
rlabel metal1 315 -4956 407 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_171/VGND
rlabel metal1 315 -4412 407 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_171/VPWR
flabel metal1 1540 -4925 1574 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_85/VGND
flabel metal1 1540 -4381 1574 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_85/VPWR
flabel nwell 1540 -4381 1574 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_85/VPB
flabel pwell 1540 -4925 1574 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_85/VNB
rlabel comment 1603 -4908 1603 -4908 6 sky130_fd_sc_hd__decap_4_85/decap_4
rlabel metal1 1235 -4956 1603 -4860 1 sky130_fd_sc_hd__decap_4_85/VGND
rlabel metal1 1235 -4412 1603 -4316 1 sky130_fd_sc_hd__decap_4_85/VPWR
flabel metal1 2828 -4925 2862 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_86/VGND
flabel metal1 2828 -4381 2862 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_86/VPWR
flabel nwell 2828 -4381 2862 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_86/VPB
flabel pwell 2828 -4925 2862 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_86/VNB
rlabel comment 2891 -4908 2891 -4908 6 sky130_fd_sc_hd__decap_4_86/decap_4
rlabel metal1 2523 -4956 2891 -4860 1 sky130_fd_sc_hd__decap_4_86/VGND
rlabel metal1 2523 -4412 2891 -4316 1 sky130_fd_sc_hd__decap_4_86/VPWR
flabel metal1 1724 -4381 1758 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_98/VPWR
flabel metal1 1724 -4925 1758 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_98/VGND
flabel nwell 1724 -4381 1758 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_98/VPB
flabel pwell 1724 -4925 1758 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_98/VNB
rlabel comment 1695 -4908 1695 -4908 4 sky130_fd_sc_hd__decap_8_98/decap_8
rlabel metal1 1695 -4956 2431 -4860 1 sky130_fd_sc_hd__decap_8_98/VGND
rlabel metal1 1695 -4412 2431 -4316 1 sky130_fd_sc_hd__decap_8_98/VPWR
flabel metal1 1160 -4384 1213 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_172/VPWR
flabel metal1 1163 -4926 1214 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_172/VGND
rlabel comment 1235 -4908 1235 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_172/tapvpwrvgnd_1
rlabel metal1 1143 -4956 1235 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_172/VGND
rlabel metal1 1143 -4412 1235 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_172/VPWR
flabel metal1 1620 -4384 1673 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_173/VPWR
flabel metal1 1623 -4926 1674 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_173/VGND
rlabel comment 1695 -4908 1695 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_173/tapvpwrvgnd_1
rlabel metal1 1603 -4956 1695 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_173/VGND
rlabel metal1 1603 -4412 1695 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_173/VPWR
flabel metal1 2448 -4384 2501 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_174/VPWR
flabel metal1 2451 -4926 2502 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_174/VGND
rlabel comment 2523 -4908 2523 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_174/tapvpwrvgnd_1
rlabel metal1 2431 -4956 2523 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_174/VGND
rlabel metal1 2431 -4412 2523 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_174/VPWR
flabel locali 3655 -4687 3689 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/A
flabel locali 3009 -4483 3043 -4449 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X
flabel locali 3009 -4551 3043 -4517 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X
flabel locali 3009 -4619 3043 -4585 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X
flabel locali 3009 -4687 3043 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X
flabel locali 3009 -4755 3043 -4721 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X
flabel locali 3009 -4823 3043 -4789 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X
flabel pwell 3655 -4925 3689 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/VNB
flabel nwell 3655 -4381 3689 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/VPB
flabel metal1 3655 -4925 3689 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/VGND
flabel metal1 3655 -4381 3689 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_71/VPWR
rlabel comment 3719 -4908 3719 -4908 6 sky130_fd_sc_hd__clkdlybuf4s50_1_71/clkdlybuf4s50_1
rlabel metal1 2983 -4956 3719 -4860 1 sky130_fd_sc_hd__clkdlybuf4s50_1_71/VGND
rlabel metal1 2983 -4412 3719 -4316 1 sky130_fd_sc_hd__clkdlybuf4s50_1_71/VPWR
flabel metal1 4116 -4925 4150 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_87/VGND
flabel metal1 4116 -4381 4150 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_87/VPWR
flabel nwell 4116 -4381 4150 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_87/VPB
flabel pwell 4116 -4925 4150 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_87/VNB
rlabel comment 4179 -4908 4179 -4908 6 sky130_fd_sc_hd__decap_4_87/decap_4
rlabel metal1 3811 -4956 4179 -4860 1 sky130_fd_sc_hd__decap_4_87/VGND
rlabel metal1 3811 -4412 4179 -4316 1 sky130_fd_sc_hd__decap_4_87/VPWR
flabel metal1 4300 -4381 4334 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_102/VPWR
flabel metal1 4300 -4925 4334 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_102/VGND
flabel nwell 4300 -4381 4334 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_102/VPB
flabel pwell 4300 -4925 4334 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_102/VNB
rlabel comment 4271 -4908 4271 -4908 4 sky130_fd_sc_hd__decap_8_102/decap_8
rlabel metal1 4271 -4956 5007 -4860 1 sky130_fd_sc_hd__decap_8_102/VGND
rlabel metal1 4271 -4412 5007 -4316 1 sky130_fd_sc_hd__decap_8_102/VPWR
flabel metal1 2908 -4384 2961 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_175/VPWR
flabel metal1 2911 -4926 2962 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_175/VGND
rlabel comment 2983 -4908 2983 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_175/tapvpwrvgnd_1
rlabel metal1 2891 -4956 2983 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_175/VGND
rlabel metal1 2891 -4412 2983 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_175/VPWR
flabel metal1 3736 -4384 3789 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_176/VPWR
flabel metal1 3739 -4926 3790 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_176/VGND
rlabel comment 3811 -4908 3811 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_176/tapvpwrvgnd_1
rlabel metal1 3719 -4956 3811 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_176/VGND
rlabel metal1 3719 -4412 3811 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_176/VPWR
flabel metal1 4196 -4384 4249 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_177/VPWR
flabel metal1 4199 -4926 4250 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_177/VGND
rlabel comment 4271 -4908 4271 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_177/tapvpwrvgnd_1
rlabel metal1 4179 -4956 4271 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_177/VGND
rlabel metal1 4179 -4412 4271 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_177/VPWR
flabel locali 6231 -4687 6265 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/A
flabel locali 5585 -4483 5619 -4449 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
flabel locali 5585 -4551 5619 -4517 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
flabel locali 5585 -4619 5619 -4585 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
flabel locali 5585 -4687 5619 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
flabel locali 5585 -4755 5619 -4721 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
flabel locali 5585 -4823 5619 -4789 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
flabel pwell 6231 -4925 6265 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/VNB
flabel nwell 6231 -4381 6265 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/VPB
flabel metal1 6231 -4925 6265 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/VGND
flabel metal1 6231 -4381 6265 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_73/VPWR
rlabel comment 6295 -4908 6295 -4908 6 sky130_fd_sc_hd__clkdlybuf4s50_1_73/clkdlybuf4s50_1
rlabel metal1 5559 -4956 6295 -4860 1 sky130_fd_sc_hd__clkdlybuf4s50_1_73/VGND
rlabel metal1 5559 -4412 6295 -4316 1 sky130_fd_sc_hd__clkdlybuf4s50_1_73/VPWR
flabel metal1 5404 -4925 5438 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_88/VGND
flabel metal1 5404 -4381 5438 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_88/VPWR
flabel nwell 5404 -4381 5438 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_88/VPB
flabel pwell 5404 -4925 5438 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_88/VNB
rlabel comment 5467 -4908 5467 -4908 6 sky130_fd_sc_hd__decap_4_88/decap_4
rlabel metal1 5099 -4956 5467 -4860 1 sky130_fd_sc_hd__decap_4_88/VGND
rlabel metal1 5099 -4412 5467 -4316 1 sky130_fd_sc_hd__decap_4_88/VPWR
flabel metal1 6692 -4925 6726 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_89/VGND
flabel metal1 6692 -4381 6726 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_89/VPWR
flabel nwell 6692 -4381 6726 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_89/VPB
flabel pwell 6692 -4925 6726 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_89/VNB
rlabel comment 6755 -4908 6755 -4908 6 sky130_fd_sc_hd__decap_4_89/decap_4
rlabel metal1 6387 -4956 6755 -4860 1 sky130_fd_sc_hd__decap_4_89/VGND
rlabel metal1 6387 -4412 6755 -4316 1 sky130_fd_sc_hd__decap_4_89/VPWR
flabel metal1 5024 -4384 5077 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_178/VPWR
flabel metal1 5027 -4926 5078 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_178/VGND
rlabel comment 5099 -4908 5099 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_178/tapvpwrvgnd_1
rlabel metal1 5007 -4956 5099 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_178/VGND
rlabel metal1 5007 -4412 5099 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_178/VPWR
flabel metal1 5484 -4384 5537 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_179/VPWR
flabel metal1 5487 -4926 5538 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_179/VGND
rlabel comment 5559 -4908 5559 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_179/tapvpwrvgnd_1
rlabel metal1 5467 -4956 5559 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_179/VGND
rlabel metal1 5467 -4412 5559 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_179/VPWR
flabel metal1 6312 -4384 6365 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_180/VPWR
flabel metal1 6315 -4926 6366 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_180/VGND
rlabel comment 6387 -4908 6387 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_180/tapvpwrvgnd_1
rlabel metal1 6295 -4956 6387 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_180/VGND
rlabel metal1 6295 -4412 6387 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_180/VPWR
flabel locali 8807 -4687 8841 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/A
flabel locali 8161 -4483 8195 -4449 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
flabel locali 8161 -4551 8195 -4517 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
flabel locali 8161 -4619 8195 -4585 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
flabel locali 8161 -4687 8195 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
flabel locali 8161 -4755 8195 -4721 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
flabel locali 8161 -4823 8195 -4789 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
flabel pwell 8807 -4925 8841 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/VNB
flabel nwell 8807 -4381 8841 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/VPB
flabel metal1 8807 -4925 8841 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/VGND
flabel metal1 8807 -4381 8841 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_75/VPWR
rlabel comment 8871 -4908 8871 -4908 6 sky130_fd_sc_hd__clkdlybuf4s50_1_75/clkdlybuf4s50_1
rlabel metal1 8135 -4956 8871 -4860 1 sky130_fd_sc_hd__clkdlybuf4s50_1_75/VGND
rlabel metal1 8135 -4412 8871 -4316 1 sky130_fd_sc_hd__clkdlybuf4s50_1_75/VPWR
flabel metal1 7980 -4925 8014 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_90/VGND
flabel metal1 7980 -4381 8014 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_90/VPWR
flabel nwell 7980 -4381 8014 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_90/VPB
flabel pwell 7980 -4925 8014 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_90/VNB
rlabel comment 8043 -4908 8043 -4908 6 sky130_fd_sc_hd__decap_4_90/decap_4
rlabel metal1 7675 -4956 8043 -4860 1 sky130_fd_sc_hd__decap_4_90/VGND
rlabel metal1 7675 -4412 8043 -4316 1 sky130_fd_sc_hd__decap_4_90/VPWR
flabel metal1 6876 -4381 6910 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_114/VPWR
flabel metal1 6876 -4925 6910 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_114/VGND
flabel nwell 6876 -4381 6910 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_114/VPB
flabel pwell 6876 -4925 6910 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_114/VNB
rlabel comment 6847 -4908 6847 -4908 4 sky130_fd_sc_hd__decap_8_114/decap_8
rlabel metal1 6847 -4956 7583 -4860 1 sky130_fd_sc_hd__decap_8_114/VGND
rlabel metal1 6847 -4412 7583 -4316 1 sky130_fd_sc_hd__decap_8_114/VPWR
flabel metal1 6772 -4384 6825 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_181/VPWR
flabel metal1 6775 -4926 6826 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_181/VGND
rlabel comment 6847 -4908 6847 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_181/tapvpwrvgnd_1
rlabel metal1 6755 -4956 6847 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_181/VGND
rlabel metal1 6755 -4412 6847 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_181/VPWR
flabel metal1 7600 -4384 7653 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_182/VPWR
flabel metal1 7603 -4926 7654 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_182/VGND
rlabel comment 7675 -4908 7675 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_182/tapvpwrvgnd_1
rlabel metal1 7583 -4956 7675 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_182/VGND
rlabel metal1 7583 -4412 7675 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_182/VPWR
flabel metal1 8060 -4384 8113 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_183/VPWR
flabel metal1 8063 -4926 8114 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_183/VGND
rlabel comment 8135 -4908 8135 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_183/tapvpwrvgnd_1
rlabel metal1 8043 -4956 8135 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_183/VGND
rlabel metal1 8043 -4412 8135 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_183/VPWR
flabel metal1 9268 -4925 9302 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_91/VGND
flabel metal1 9268 -4381 9302 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_91/VPWR
flabel nwell 9268 -4381 9302 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_91/VPB
flabel pwell 9268 -4925 9302 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_91/VNB
rlabel comment 9331 -4908 9331 -4908 6 sky130_fd_sc_hd__decap_4_91/decap_4
rlabel metal1 8963 -4956 9331 -4860 1 sky130_fd_sc_hd__decap_4_91/VGND
rlabel metal1 8963 -4412 9331 -4316 1 sky130_fd_sc_hd__decap_4_91/VPWR
flabel metal1 10648 -4925 10682 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_92/VGND
flabel metal1 10648 -4381 10682 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_92/VPWR
flabel nwell 10648 -4381 10682 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_92/VPB
flabel pwell 10648 -4925 10682 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_92/VNB
rlabel comment 10711 -4908 10711 -4908 6 sky130_fd_sc_hd__decap_4_92/decap_4
rlabel metal1 10343 -4956 10711 -4860 1 sky130_fd_sc_hd__decap_4_92/VGND
rlabel metal1 10343 -4412 10711 -4316 1 sky130_fd_sc_hd__decap_4_92/VPWR
flabel metal1 9452 -4381 9486 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_124/VPWR
flabel metal1 9452 -4925 9486 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_124/VGND
flabel nwell 9452 -4381 9486 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_124/VPB
flabel pwell 9452 -4925 9486 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_124/VNB
rlabel comment 9423 -4908 9423 -4908 4 sky130_fd_sc_hd__decap_8_124/decap_8
rlabel metal1 9423 -4956 10159 -4860 1 sky130_fd_sc_hd__decap_8_124/VGND
rlabel metal1 9423 -4412 10159 -4316 1 sky130_fd_sc_hd__decap_8_124/VPWR
flabel metal1 10285 -4381 10321 -4351 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_24/VPWR
flabel metal1 10285 -4921 10321 -4892 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_24/VGND
flabel nwell 10292 -4374 10312 -4357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_24/VPB
flabel pwell 10291 -4919 10315 -4897 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_24/VNB
rlabel comment 10343 -4908 10343 -4908 6 sky130_fd_sc_hd__fill_1_24/fill_1
rlabel metal1 10251 -4956 10343 -4860 1 sky130_fd_sc_hd__fill_1_24/VGND
rlabel metal1 10251 -4412 10343 -4316 1 sky130_fd_sc_hd__fill_1_24/VPWR
flabel metal1 9348 -4384 9401 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_184/VPWR
flabel metal1 9351 -4926 9402 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_184/VGND
rlabel comment 9423 -4908 9423 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_184/tapvpwrvgnd_1
rlabel metal1 9331 -4956 9423 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_184/VGND
rlabel metal1 9331 -4412 9423 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_184/VPWR
flabel metal1 8888 -4384 8941 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_185/VPWR
flabel metal1 8891 -4926 8942 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_185/VGND
rlabel comment 8963 -4908 8963 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_185/tapvpwrvgnd_1
rlabel metal1 8871 -4956 8963 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_185/VGND
rlabel metal1 8871 -4412 8963 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_185/VPWR
flabel metal1 10176 -4384 10229 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_186/VPWR
flabel metal1 10179 -4926 10230 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_186/VGND
rlabel comment 10251 -4908 10251 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_186/tapvpwrvgnd_1
rlabel metal1 10159 -4956 10251 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_186/VGND
rlabel metal1 10159 -4412 10251 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_186/VPWR
flabel locali 11383 -4687 11417 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/A
flabel locali 10737 -4483 10771 -4449 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
flabel locali 10737 -4551 10771 -4517 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
flabel locali 10737 -4619 10771 -4585 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
flabel locali 10737 -4687 10771 -4653 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
flabel locali 10737 -4755 10771 -4721 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
flabel locali 10737 -4823 10771 -4789 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
flabel pwell 11383 -4925 11417 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/VNB
flabel nwell 11383 -4381 11417 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/VPB
flabel metal1 11383 -4925 11417 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/VGND
flabel metal1 11383 -4381 11417 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_77/VPWR
rlabel comment 11447 -4908 11447 -4908 6 sky130_fd_sc_hd__clkdlybuf4s50_1_77/clkdlybuf4s50_1
rlabel metal1 10711 -4956 11447 -4860 1 sky130_fd_sc_hd__clkdlybuf4s50_1_77/VGND
rlabel metal1 10711 -4412 11447 -4316 1 sky130_fd_sc_hd__clkdlybuf4s50_1_77/VPWR
flabel metal1 11936 -4925 11970 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_93/VGND
flabel metal1 11936 -4381 11970 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_93/VPWR
flabel nwell 11936 -4381 11970 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_93/VPB
flabel pwell 11936 -4925 11970 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_93/VNB
rlabel comment 11999 -4908 11999 -4908 6 sky130_fd_sc_hd__decap_4_93/decap_4
rlabel metal1 11631 -4956 11999 -4860 1 sky130_fd_sc_hd__decap_4_93/VGND
rlabel metal1 11631 -4412 11999 -4316 1 sky130_fd_sc_hd__decap_4_93/VPWR
flabel metal1 10653 -4381 10689 -4351 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_25/VPWR
flabel metal1 10653 -4921 10689 -4892 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_25/VGND
flabel nwell 10660 -4374 10680 -4357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_25/VPB
flabel pwell 10659 -4919 10683 -4897 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_25/VNB
rlabel comment 10711 -4908 10711 -4908 6 sky130_fd_sc_hd__fill_1_25/fill_1
rlabel metal1 10619 -4956 10711 -4860 1 sky130_fd_sc_hd__fill_1_25/VGND
rlabel metal1 10619 -4412 10711 -4316 1 sky130_fd_sc_hd__fill_1_25/VPWR
flabel metal1 11573 -4381 11609 -4351 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_26/VPWR
flabel metal1 11573 -4921 11609 -4892 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_26/VGND
flabel nwell 11580 -4374 11600 -4357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_26/VPB
flabel pwell 11579 -4919 11603 -4897 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_26/VNB
rlabel comment 11631 -4908 11631 -4908 6 sky130_fd_sc_hd__fill_1_26/fill_1
rlabel metal1 11539 -4956 11631 -4860 1 sky130_fd_sc_hd__fill_1_26/VGND
rlabel metal1 11539 -4412 11631 -4316 1 sky130_fd_sc_hd__fill_1_26/VPWR
flabel metal1 12668 -4928 12700 -4898 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_11/VGND
flabel metal1 12668 -4385 12706 -4353 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_11/VPWR
flabel nwell 12658 -4386 12715 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_11/VPB
flabel pwell 12665 -4932 12709 -4898 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_11/VNB
rlabel comment 12735 -4908 12735 -4908 6 sky130_fd_sc_hd__fill_8_11/fill_8
rlabel metal1 11999 -4956 12735 -4860 1 sky130_fd_sc_hd__fill_8_11/VGND
rlabel metal1 11999 -4412 12735 -4316 1 sky130_fd_sc_hd__fill_8_11/VPWR
flabel metal1 11464 -4384 11517 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_187/VPWR
flabel metal1 11467 -4926 11518 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_187/VGND
rlabel comment 11539 -4908 11539 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_187/tapvpwrvgnd_1
rlabel metal1 11447 -4956 11539 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_187/VGND
rlabel metal1 11447 -4412 11539 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_187/VPWR
flabel locali 15248 -4619 15282 -4585 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/X
flabel locali 15340 -4619 15374 -4585 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/X
flabel locali 15340 -4687 15374 -4653 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/X
flabel locali 15248 -4687 15282 -4653 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/X
flabel locali 15248 -4755 15282 -4721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/X
flabel locali 15340 -4755 15374 -4721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/X
flabel locali 13684 -4755 13718 -4721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/A
flabel locali 13684 -4687 13718 -4653 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/A
flabel pwell 13684 -4925 13718 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/VNB
flabel pwell 13701 -4908 13701 -4908 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/VNB
flabel nwell 13684 -4381 13718 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/VPB
flabel nwell 13701 -4364 13701 -4364 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/VPB
flabel metal1 13684 -4925 13718 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/VGND
flabel metal1 13684 -4381 13718 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_5/VPWR
rlabel comment 13655 -4908 13655 -4908 4 sky130_fd_sc_hd__clkbuf_16_5/clkbuf_16
rlabel metal1 13655 -4956 15495 -4860 1 sky130_fd_sc_hd__clkbuf_16_5/VGND
rlabel metal1 13655 -4412 15495 -4316 1 sky130_fd_sc_hd__clkbuf_16_5/VPWR
flabel metal1 13505 -4381 13541 -4351 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_27/VPWR
flabel metal1 13505 -4921 13541 -4892 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_27/VGND
flabel nwell 13512 -4374 13532 -4357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_27/VPB
flabel pwell 13511 -4919 13535 -4897 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_27/VNB
rlabel comment 13563 -4908 13563 -4908 6 sky130_fd_sc_hd__fill_1_27/fill_1
rlabel metal1 13471 -4956 13563 -4860 1 sky130_fd_sc_hd__fill_1_27/VGND
rlabel metal1 13471 -4412 13563 -4316 1 sky130_fd_sc_hd__fill_1_27/VPWR
flabel metal1 13404 -4928 13436 -4898 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_12/VGND
flabel metal1 13404 -4385 13442 -4353 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_12/VPWR
flabel nwell 13394 -4386 13451 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_12/VPB
flabel pwell 13401 -4932 13445 -4898 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_12/VNB
rlabel comment 13471 -4908 13471 -4908 6 sky130_fd_sc_hd__fill_8_12/fill_8
rlabel metal1 12735 -4956 13471 -4860 1 sky130_fd_sc_hd__fill_8_12/VGND
rlabel metal1 12735 -4412 13471 -4316 1 sky130_fd_sc_hd__fill_8_12/VPWR
flabel metal1 13580 -4384 13633 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_188/VPWR
flabel metal1 13583 -4926 13634 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_188/VGND
rlabel comment 13655 -4908 13655 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_188/tapvpwrvgnd_1
rlabel metal1 13563 -4956 13655 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_188/VGND
rlabel metal1 13563 -4412 13655 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_188/VPWR
flabel metal1 16628 -4925 16662 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_12/VGND
flabel metal1 16628 -4381 16662 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_12/VPWR
flabel nwell 16628 -4381 16662 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_12/VPB
flabel pwell 16628 -4925 16662 -4891 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_12/VNB
rlabel comment 16691 -4908 16691 -4908 6 sky130_fd_sc_hd__decap_12_12/decap_12
rlabel metal1 15587 -4956 16691 -4860 1 sky130_fd_sc_hd__decap_12_12/VGND
rlabel metal1 15587 -4412 16691 -4316 1 sky130_fd_sc_hd__decap_12_12/VPWR
flabel metal1 15512 -4384 15565 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_189/VPWR
flabel metal1 15515 -4926 15566 -4888 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_189/VGND
rlabel comment 15587 -4908 15587 -4908 6 sky130_fd_sc_hd__tapvpwrvgnd_1_189/tapvpwrvgnd_1
rlabel metal1 15495 -4956 15587 -4860 1 sky130_fd_sc_hd__tapvpwrvgnd_1_189/VGND
rlabel metal1 15495 -4412 15587 -4316 1 sky130_fd_sc_hd__tapvpwrvgnd_1_189/VPWR
flabel metal1 -1588 -4381 -1554 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_14/VPWR
flabel metal1 -1588 -3837 -1554 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_14/VGND
flabel nwell -1588 -4381 -1554 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_14/VPB
flabel pwell -1588 -3837 -1554 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_14/VNB
rlabel comment -1617 -3820 -1617 -3820 2 sky130_fd_sc_hd__decap_8_14/decap_8
rlabel metal1 -1617 -3868 -881 -3772 5 sky130_fd_sc_hd__decap_8_14/VGND
rlabel metal1 -1617 -4412 -881 -4316 5 sky130_fd_sc_hd__decap_8_14/VPWR
flabel metal1 -2324 -4381 -2290 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_73/VPWR
flabel metal1 -2324 -3837 -2290 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_73/VGND
flabel nwell -2324 -4381 -2290 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_73/VPB
flabel pwell -2324 -3837 -2290 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_73/VNB
rlabel comment -2261 -3820 -2261 -3820 8 sky130_fd_sc_hd__decap_8_73/decap_8
rlabel metal1 -2997 -3868 -2261 -3772 5 sky130_fd_sc_hd__decap_8_73/VGND
rlabel metal1 -2997 -4412 -2261 -4316 5 sky130_fd_sc_hd__decap_8_73/VPWR
flabel metal1 -1690 -3838 -1637 -3806 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_10/VGND
flabel metal1 -1690 -4381 -1638 -4350 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_10/VPWR
flabel nwell -1679 -4373 -1645 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_10/VPB
flabel pwell -1680 -3832 -1648 -3810 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_10/VNB
rlabel comment -1617 -3820 -1617 -3820 8 sky130_fd_sc_hd__fill_2_10/fill_2
rlabel metal1 -1801 -3868 -1617 -3772 5 sky130_fd_sc_hd__fill_2_10/VGND
rlabel metal1 -1801 -4412 -1617 -4316 5 sky130_fd_sc_hd__fill_2_10/VPWR
flabel metal1 -1858 -3829 -1835 -3810 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_23/VGND
flabel metal1 -1855 -4372 -1835 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_23/VPWR
flabel nwell -1861 -4376 -1836 -4350 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_23/VPB
flabel pwell -1858 -3832 -1836 -3808 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_23/VNB
rlabel comment -1801 -3820 -1801 -3820 8 sky130_fd_sc_hd__fill_4_23/fill_4
rlabel metal1 -2169 -3868 -1801 -3772 5 sky130_fd_sc_hd__fill_4_23/VGND
rlabel metal1 -2169 -4412 -1801 -4316 5 sky130_fd_sc_hd__fill_4_23/VPWR
flabel metal1 -2244 -4373 -2191 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_538/VPWR
flabel metal1 -2241 -3840 -2190 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_538/VGND
rlabel comment -2169 -3820 -2169 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_538/tapvpwrvgnd_1
rlabel metal1 -2261 -3868 -2169 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_538/VGND
rlabel metal1 -2261 -4412 -2169 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_538/VPWR
flabel locali 437 -4075 471 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/A
flabel locali 1083 -4279 1117 -4245 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/X
flabel locali 1083 -4211 1117 -4177 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/X
flabel locali 1083 -4143 1117 -4109 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/X
flabel locali 1083 -4075 1117 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/X
flabel locali 1083 -4007 1117 -3973 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/X
flabel locali 1083 -3939 1117 -3905 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/X
flabel pwell 437 -3837 471 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/VNB
flabel nwell 437 -4381 471 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/VPB
flabel metal1 437 -3837 471 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/VGND
flabel metal1 437 -4381 471 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_59/VPWR
rlabel comment 407 -3820 407 -3820 2 sky130_fd_sc_hd__clkdlybuf4s50_1_59/clkdlybuf4s50_1
rlabel metal1 407 -3868 1143 -3772 5 sky130_fd_sc_hd__clkdlybuf4s50_1_59/VGND
rlabel metal1 407 -4412 1143 -4316 5 sky130_fd_sc_hd__clkdlybuf4s50_1_59/VPWR
flabel metal1 252 -3837 286 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_73/VGND
flabel metal1 252 -4381 286 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_73/VPWR
flabel nwell 252 -4381 286 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_73/VPB
flabel pwell 252 -3837 286 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_73/VNB
rlabel comment 315 -3820 315 -3820 8 sky130_fd_sc_hd__decap_4_73/decap_4
rlabel metal1 -53 -3868 315 -3772 5 sky130_fd_sc_hd__decap_4_73/VGND
rlabel metal1 -53 -4412 315 -4316 5 sky130_fd_sc_hd__decap_4_73/VPWR
flabel metal1 -852 -4381 -818 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_15/VPWR
flabel metal1 -852 -3837 -818 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_15/VGND
flabel nwell -852 -4381 -818 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_15/VPB
flabel pwell -852 -3837 -818 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_15/VNB
rlabel comment -881 -3820 -881 -3820 2 sky130_fd_sc_hd__decap_8_15/decap_8
rlabel metal1 -881 -3868 -145 -3772 5 sky130_fd_sc_hd__decap_8_15/VGND
rlabel metal1 -881 -4412 -145 -4316 5 sky130_fd_sc_hd__decap_8_15/VPWR
flabel metal1 -128 -4373 -75 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_148/VPWR
flabel metal1 -125 -3840 -74 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_148/VGND
rlabel comment -53 -3820 -53 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_148/tapvpwrvgnd_1
rlabel metal1 -145 -3868 -53 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_148/VGND
rlabel metal1 -145 -4412 -53 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_148/VPWR
flabel metal1 332 -4373 385 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_149/VPWR
flabel metal1 335 -3840 386 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_149/VGND
rlabel comment 407 -3820 407 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_149/tapvpwrvgnd_1
rlabel metal1 315 -3868 407 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_149/VGND
rlabel metal1 315 -4412 407 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_149/VPWR
flabel metal1 1540 -3837 1574 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_74/VGND
flabel metal1 1540 -4381 1574 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_74/VPWR
flabel nwell 1540 -4381 1574 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_74/VPB
flabel pwell 1540 -3837 1574 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_74/VNB
rlabel comment 1603 -3820 1603 -3820 8 sky130_fd_sc_hd__decap_4_74/decap_4
rlabel metal1 1235 -3868 1603 -3772 5 sky130_fd_sc_hd__decap_4_74/VGND
rlabel metal1 1235 -4412 1603 -4316 5 sky130_fd_sc_hd__decap_4_74/VPWR
flabel metal1 2828 -3837 2862 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_75/VGND
flabel metal1 2828 -4381 2862 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_75/VPWR
flabel nwell 2828 -4381 2862 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_75/VPB
flabel pwell 2828 -3837 2862 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_75/VNB
rlabel comment 2891 -3820 2891 -3820 8 sky130_fd_sc_hd__decap_4_75/decap_4
rlabel metal1 2523 -3868 2891 -3772 5 sky130_fd_sc_hd__decap_4_75/VGND
rlabel metal1 2523 -4412 2891 -4316 5 sky130_fd_sc_hd__decap_4_75/VPWR
flabel metal1 2368 -4381 2402 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_97/VPWR
flabel metal1 2368 -3837 2402 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_97/VGND
flabel nwell 2368 -4381 2402 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_97/VPB
flabel pwell 2368 -3837 2402 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_97/VNB
rlabel comment 2431 -3820 2431 -3820 8 sky130_fd_sc_hd__decap_8_97/decap_8
rlabel metal1 1695 -3868 2431 -3772 5 sky130_fd_sc_hd__decap_8_97/VGND
rlabel metal1 1695 -4412 2431 -4316 5 sky130_fd_sc_hd__decap_8_97/VPWR
flabel metal1 1160 -4373 1213 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_150/VPWR
flabel metal1 1163 -3840 1214 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_150/VGND
rlabel comment 1235 -3820 1235 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_150/tapvpwrvgnd_1
rlabel metal1 1143 -3868 1235 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_150/VGND
rlabel metal1 1143 -4412 1235 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_150/VPWR
flabel metal1 1620 -4373 1673 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_151/VPWR
flabel metal1 1623 -3840 1674 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_151/VGND
rlabel comment 1695 -3820 1695 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_151/tapvpwrvgnd_1
rlabel metal1 1603 -3868 1695 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_151/VGND
rlabel metal1 1603 -4412 1695 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_151/VPWR
flabel metal1 2448 -4373 2501 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_152/VPWR
flabel metal1 2451 -3840 2502 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_152/VGND
rlabel comment 2523 -3820 2523 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_152/tapvpwrvgnd_1
rlabel metal1 2431 -3868 2523 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_152/VGND
rlabel metal1 2431 -4412 2523 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_152/VPWR
flabel locali 3013 -4075 3047 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A
flabel locali 3659 -4279 3693 -4245 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/X
flabel locali 3659 -4211 3693 -4177 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/X
flabel locali 3659 -4143 3693 -4109 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/X
flabel locali 3659 -4075 3693 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/X
flabel locali 3659 -4007 3693 -3973 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/X
flabel locali 3659 -3939 3693 -3905 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/X
flabel pwell 3013 -3837 3047 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/VNB
flabel nwell 3013 -4381 3047 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/VPB
flabel metal1 3013 -3837 3047 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/VGND
flabel metal1 3013 -4381 3047 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_61/VPWR
rlabel comment 2983 -3820 2983 -3820 2 sky130_fd_sc_hd__clkdlybuf4s50_1_61/clkdlybuf4s50_1
rlabel metal1 2983 -3868 3719 -3772 5 sky130_fd_sc_hd__clkdlybuf4s50_1_61/VGND
rlabel metal1 2983 -4412 3719 -4316 5 sky130_fd_sc_hd__clkdlybuf4s50_1_61/VPWR
flabel metal1 4116 -3837 4150 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_76/VGND
flabel metal1 4116 -4381 4150 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_76/VPWR
flabel nwell 4116 -4381 4150 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_76/VPB
flabel pwell 4116 -3837 4150 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_76/VNB
rlabel comment 4179 -3820 4179 -3820 8 sky130_fd_sc_hd__decap_4_76/decap_4
rlabel metal1 3811 -3868 4179 -3772 5 sky130_fd_sc_hd__decap_4_76/VGND
rlabel metal1 3811 -4412 4179 -4316 5 sky130_fd_sc_hd__decap_4_76/VPWR
flabel metal1 4944 -4381 4978 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_105/VPWR
flabel metal1 4944 -3837 4978 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_105/VGND
flabel nwell 4944 -4381 4978 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_105/VPB
flabel pwell 4944 -3837 4978 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_105/VNB
rlabel comment 5007 -3820 5007 -3820 8 sky130_fd_sc_hd__decap_8_105/decap_8
rlabel metal1 4271 -3868 5007 -3772 5 sky130_fd_sc_hd__decap_8_105/VGND
rlabel metal1 4271 -4412 5007 -4316 5 sky130_fd_sc_hd__decap_8_105/VPWR
flabel metal1 2908 -4373 2961 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_153/VPWR
flabel metal1 2911 -3840 2962 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_153/VGND
rlabel comment 2983 -3820 2983 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_153/tapvpwrvgnd_1
rlabel metal1 2891 -3868 2983 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_153/VGND
rlabel metal1 2891 -4412 2983 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_153/VPWR
flabel metal1 3736 -4373 3789 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_154/VPWR
flabel metal1 3739 -3840 3790 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_154/VGND
rlabel comment 3811 -3820 3811 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_154/tapvpwrvgnd_1
rlabel metal1 3719 -3868 3811 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_154/VGND
rlabel metal1 3719 -4412 3811 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_154/VPWR
flabel metal1 4196 -4373 4249 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_155/VPWR
flabel metal1 4199 -3840 4250 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_155/VGND
rlabel comment 4271 -3820 4271 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_155/tapvpwrvgnd_1
rlabel metal1 4179 -3868 4271 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_155/VGND
rlabel metal1 4179 -4412 4271 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_155/VPWR
flabel locali 5589 -4075 5623 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A
flabel locali 6235 -4279 6269 -4245 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/X
flabel locali 6235 -4211 6269 -4177 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/X
flabel locali 6235 -4143 6269 -4109 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/X
flabel locali 6235 -4075 6269 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/X
flabel locali 6235 -4007 6269 -3973 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/X
flabel locali 6235 -3939 6269 -3905 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/X
flabel pwell 5589 -3837 5623 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/VNB
flabel nwell 5589 -4381 5623 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/VPB
flabel metal1 5589 -3837 5623 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/VGND
flabel metal1 5589 -4381 5623 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_63/VPWR
rlabel comment 5559 -3820 5559 -3820 2 sky130_fd_sc_hd__clkdlybuf4s50_1_63/clkdlybuf4s50_1
rlabel metal1 5559 -3868 6295 -3772 5 sky130_fd_sc_hd__clkdlybuf4s50_1_63/VGND
rlabel metal1 5559 -4412 6295 -4316 5 sky130_fd_sc_hd__clkdlybuf4s50_1_63/VPWR
flabel metal1 5404 -3837 5438 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_77/VGND
flabel metal1 5404 -4381 5438 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_77/VPWR
flabel nwell 5404 -4381 5438 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_77/VPB
flabel pwell 5404 -3837 5438 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_77/VNB
rlabel comment 5467 -3820 5467 -3820 8 sky130_fd_sc_hd__decap_4_77/decap_4
rlabel metal1 5099 -3868 5467 -3772 5 sky130_fd_sc_hd__decap_4_77/VGND
rlabel metal1 5099 -4412 5467 -4316 5 sky130_fd_sc_hd__decap_4_77/VPWR
flabel metal1 6692 -3837 6726 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_78/VGND
flabel metal1 6692 -4381 6726 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_78/VPWR
flabel nwell 6692 -4381 6726 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_78/VPB
flabel pwell 6692 -3837 6726 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_78/VNB
rlabel comment 6755 -3820 6755 -3820 8 sky130_fd_sc_hd__decap_4_78/decap_4
rlabel metal1 6387 -3868 6755 -3772 5 sky130_fd_sc_hd__decap_4_78/VGND
rlabel metal1 6387 -4412 6755 -4316 5 sky130_fd_sc_hd__decap_4_78/VPWR
flabel metal1 5024 -4373 5077 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_156/VPWR
flabel metal1 5027 -3840 5078 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_156/VGND
rlabel comment 5099 -3820 5099 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_156/tapvpwrvgnd_1
rlabel metal1 5007 -3868 5099 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_156/VGND
rlabel metal1 5007 -4412 5099 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_156/VPWR
flabel metal1 5484 -4373 5537 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_157/VPWR
flabel metal1 5487 -3840 5538 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_157/VGND
rlabel comment 5559 -3820 5559 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_157/tapvpwrvgnd_1
rlabel metal1 5467 -3868 5559 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_157/VGND
rlabel metal1 5467 -4412 5559 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_157/VPWR
flabel metal1 6312 -4373 6365 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_158/VPWR
flabel metal1 6315 -3840 6366 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_158/VGND
rlabel comment 6387 -3820 6387 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_158/tapvpwrvgnd_1
rlabel metal1 6295 -3868 6387 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_158/VGND
rlabel metal1 6295 -4412 6387 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_158/VPWR
flabel locali 8165 -4075 8199 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A
flabel locali 8811 -4279 8845 -4245 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/X
flabel locali 8811 -4211 8845 -4177 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/X
flabel locali 8811 -4143 8845 -4109 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/X
flabel locali 8811 -4075 8845 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/X
flabel locali 8811 -4007 8845 -3973 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/X
flabel locali 8811 -3939 8845 -3905 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/X
flabel pwell 8165 -3837 8199 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/VNB
flabel nwell 8165 -4381 8199 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/VPB
flabel metal1 8165 -3837 8199 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/VGND
flabel metal1 8165 -4381 8199 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_65/VPWR
rlabel comment 8135 -3820 8135 -3820 2 sky130_fd_sc_hd__clkdlybuf4s50_1_65/clkdlybuf4s50_1
rlabel metal1 8135 -3868 8871 -3772 5 sky130_fd_sc_hd__clkdlybuf4s50_1_65/VGND
rlabel metal1 8135 -4412 8871 -4316 5 sky130_fd_sc_hd__clkdlybuf4s50_1_65/VPWR
flabel metal1 7980 -3837 8014 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_79/VGND
flabel metal1 7980 -4381 8014 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_79/VPWR
flabel nwell 7980 -4381 8014 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_79/VPB
flabel pwell 7980 -3837 8014 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_79/VNB
rlabel comment 8043 -3820 8043 -3820 8 sky130_fd_sc_hd__decap_4_79/decap_4
rlabel metal1 7675 -3868 8043 -3772 5 sky130_fd_sc_hd__decap_4_79/VGND
rlabel metal1 7675 -4412 8043 -4316 5 sky130_fd_sc_hd__decap_4_79/VPWR
flabel metal1 7520 -4381 7554 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_113/VPWR
flabel metal1 7520 -3837 7554 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_113/VGND
flabel nwell 7520 -4381 7554 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_113/VPB
flabel pwell 7520 -3837 7554 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_113/VNB
rlabel comment 7583 -3820 7583 -3820 8 sky130_fd_sc_hd__decap_8_113/decap_8
rlabel metal1 6847 -3868 7583 -3772 5 sky130_fd_sc_hd__decap_8_113/VGND
rlabel metal1 6847 -4412 7583 -4316 5 sky130_fd_sc_hd__decap_8_113/VPWR
flabel metal1 6772 -4373 6825 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_159/VPWR
flabel metal1 6775 -3840 6826 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_159/VGND
rlabel comment 6847 -3820 6847 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_159/tapvpwrvgnd_1
rlabel metal1 6755 -3868 6847 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_159/VGND
rlabel metal1 6755 -4412 6847 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_159/VPWR
flabel metal1 7600 -4373 7653 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_160/VPWR
flabel metal1 7603 -3840 7654 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_160/VGND
rlabel comment 7675 -3820 7675 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_160/tapvpwrvgnd_1
rlabel metal1 7583 -3868 7675 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_160/VGND
rlabel metal1 7583 -4412 7675 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_160/VPWR
flabel metal1 8060 -4373 8113 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_161/VPWR
flabel metal1 8063 -3840 8114 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_161/VGND
rlabel comment 8135 -3820 8135 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_161/tapvpwrvgnd_1
rlabel metal1 8043 -3868 8135 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_161/VGND
rlabel metal1 8043 -4412 8135 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_161/VPWR
flabel metal1 9268 -3837 9302 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_80/VGND
flabel metal1 9268 -4381 9302 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_80/VPWR
flabel nwell 9268 -4381 9302 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_80/VPB
flabel pwell 9268 -3837 9302 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_80/VNB
rlabel comment 9331 -3820 9331 -3820 8 sky130_fd_sc_hd__decap_4_80/decap_4
rlabel metal1 8963 -3868 9331 -3772 5 sky130_fd_sc_hd__decap_4_80/VGND
rlabel metal1 8963 -4412 9331 -4316 5 sky130_fd_sc_hd__decap_4_80/VPWR
flabel metal1 10648 -3837 10682 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_81/VGND
flabel metal1 10648 -4381 10682 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_81/VPWR
flabel nwell 10648 -4381 10682 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_81/VPB
flabel pwell 10648 -3837 10682 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_81/VNB
rlabel comment 10711 -3820 10711 -3820 8 sky130_fd_sc_hd__decap_4_81/decap_4
rlabel metal1 10343 -3868 10711 -3772 5 sky130_fd_sc_hd__decap_4_81/VGND
rlabel metal1 10343 -4412 10711 -4316 5 sky130_fd_sc_hd__decap_4_81/VPWR
flabel metal1 10096 -4381 10130 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_123/VPWR
flabel metal1 10096 -3837 10130 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_123/VGND
flabel nwell 10096 -4381 10130 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_123/VPB
flabel pwell 10096 -3837 10130 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_123/VNB
rlabel comment 10159 -3820 10159 -3820 8 sky130_fd_sc_hd__decap_8_123/decap_8
rlabel metal1 9423 -3868 10159 -3772 5 sky130_fd_sc_hd__decap_8_123/VGND
rlabel metal1 9423 -4412 10159 -4316 5 sky130_fd_sc_hd__decap_8_123/VPWR
flabel metal1 10285 -4377 10321 -4347 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_21/VPWR
flabel metal1 10285 -3836 10321 -3807 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_21/VGND
flabel nwell 10292 -4371 10312 -4354 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_21/VPB
flabel pwell 10291 -3831 10315 -3809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_21/VNB
rlabel comment 10343 -3820 10343 -3820 8 sky130_fd_sc_hd__fill_1_21/fill_1
rlabel metal1 10251 -3868 10343 -3772 5 sky130_fd_sc_hd__fill_1_21/VGND
rlabel metal1 10251 -4412 10343 -4316 5 sky130_fd_sc_hd__fill_1_21/VPWR
flabel metal1 9348 -4373 9401 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_162/VPWR
flabel metal1 9351 -3840 9402 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_162/VGND
rlabel comment 9423 -3820 9423 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_162/tapvpwrvgnd_1
rlabel metal1 9331 -3868 9423 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_162/VGND
rlabel metal1 9331 -4412 9423 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_162/VPWR
flabel metal1 8888 -4373 8941 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_163/VPWR
flabel metal1 8891 -3840 8942 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_163/VGND
rlabel comment 8963 -3820 8963 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_163/tapvpwrvgnd_1
rlabel metal1 8871 -3868 8963 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_163/VGND
rlabel metal1 8871 -4412 8963 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_163/VPWR
flabel metal1 10176 -4373 10229 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_164/VPWR
flabel metal1 10179 -3840 10230 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_164/VGND
rlabel comment 10251 -3820 10251 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_164/tapvpwrvgnd_1
rlabel metal1 10159 -3868 10251 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_164/VGND
rlabel metal1 10159 -4412 10251 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_164/VPWR
flabel locali 10741 -4075 10775 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A
flabel locali 11387 -4279 11421 -4245 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X
flabel locali 11387 -4211 11421 -4177 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X
flabel locali 11387 -4143 11421 -4109 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X
flabel locali 11387 -4075 11421 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X
flabel locali 11387 -4007 11421 -3973 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X
flabel locali 11387 -3939 11421 -3905 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X
flabel pwell 10741 -3837 10775 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/VNB
flabel nwell 10741 -4381 10775 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/VPB
flabel metal1 10741 -3837 10775 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/VGND
flabel metal1 10741 -4381 10775 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_67/VPWR
rlabel comment 10711 -3820 10711 -3820 2 sky130_fd_sc_hd__clkdlybuf4s50_1_67/clkdlybuf4s50_1
rlabel metal1 10711 -3868 11447 -3772 5 sky130_fd_sc_hd__clkdlybuf4s50_1_67/VGND
rlabel metal1 10711 -4412 11447 -4316 5 sky130_fd_sc_hd__clkdlybuf4s50_1_67/VPWR
flabel metal1 11936 -3837 11970 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_82/VGND
flabel metal1 11936 -4381 11970 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_82/VPWR
flabel nwell 11936 -4381 11970 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_82/VPB
flabel pwell 11936 -3837 11970 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_82/VNB
rlabel comment 11999 -3820 11999 -3820 8 sky130_fd_sc_hd__decap_4_82/decap_4
rlabel metal1 11631 -3868 11999 -3772 5 sky130_fd_sc_hd__decap_4_82/VGND
rlabel metal1 11631 -4412 11999 -4316 5 sky130_fd_sc_hd__decap_4_82/VPWR
flabel metal1 10653 -4377 10689 -4347 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_22/VPWR
flabel metal1 10653 -3836 10689 -3807 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_22/VGND
flabel nwell 10660 -4371 10680 -4354 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_22/VPB
flabel pwell 10659 -3831 10683 -3809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_22/VNB
rlabel comment 10711 -3820 10711 -3820 8 sky130_fd_sc_hd__fill_1_22/fill_1
rlabel metal1 10619 -3868 10711 -3772 5 sky130_fd_sc_hd__fill_1_22/VGND
rlabel metal1 10619 -4412 10711 -4316 5 sky130_fd_sc_hd__fill_1_22/VPWR
flabel metal1 11573 -4377 11609 -4347 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_23/VPWR
flabel metal1 11573 -3836 11609 -3807 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_23/VGND
flabel nwell 11580 -4371 11600 -4354 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_23/VPB
flabel pwell 11579 -3831 11603 -3809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_23/VNB
rlabel comment 11631 -3820 11631 -3820 8 sky130_fd_sc_hd__fill_1_23/fill_1
rlabel metal1 11539 -3868 11631 -3772 5 sky130_fd_sc_hd__fill_1_23/VGND
rlabel metal1 11539 -4412 11631 -4316 5 sky130_fd_sc_hd__fill_1_23/VPWR
flabel metal1 12033 -3829 12056 -3810 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_4/VGND
flabel metal1 12033 -4372 12053 -4355 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_4/VPWR
flabel nwell 12034 -4376 12059 -4350 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_4/VPB
flabel pwell 12034 -3832 12056 -3808 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_4/VNB
rlabel comment 11999 -3820 11999 -3820 2 sky130_fd_sc_hd__fill_4_4/fill_4
rlabel metal1 11999 -3868 12367 -3772 5 sky130_fd_sc_hd__fill_4_4/VGND
rlabel metal1 11999 -4412 12367 -4316 5 sky130_fd_sc_hd__fill_4_4/VPWR
flabel metal1 11464 -4373 11517 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_165/VPWR
flabel metal1 11467 -3840 11518 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_165/VGND
rlabel comment 11539 -3820 11539 -3820 8 sky130_fd_sc_hd__tapvpwrvgnd_1_165/tapvpwrvgnd_1
rlabel metal1 11447 -3868 11539 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_165/VGND
rlabel metal1 11447 -4412 11539 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_165/VPWR
flabel locali 15248 -4143 15282 -4109 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/X
flabel locali 15340 -4143 15374 -4109 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/X
flabel locali 15340 -4075 15374 -4041 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/X
flabel locali 15248 -4075 15282 -4041 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/X
flabel locali 15248 -4007 15282 -3973 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/X
flabel locali 15340 -4007 15374 -3973 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/X
flabel locali 13684 -4007 13718 -3973 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/A
flabel locali 13684 -4075 13718 -4041 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/A
flabel pwell 13684 -3837 13718 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/VNB
flabel pwell 13701 -3820 13701 -3820 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/VNB
flabel nwell 13684 -4381 13718 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/VPB
flabel nwell 13701 -4364 13701 -4364 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/VPB
flabel metal1 13684 -3837 13718 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/VGND
flabel metal1 13684 -4381 13718 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_4/VPWR
rlabel comment 13655 -3820 13655 -3820 2 sky130_fd_sc_hd__clkbuf_16_4/clkbuf_16
rlabel metal1 13655 -3868 15495 -3772 5 sky130_fd_sc_hd__clkbuf_16_4/VGND
rlabel metal1 13655 -4412 15495 -4316 5 sky130_fd_sc_hd__clkbuf_16_4/VPWR
flabel locali 12672 -4075 12706 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/A
flabel locali 12764 -4075 12798 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/A
flabel locali 13040 -4007 13074 -3973 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/Y
flabel locali 12580 -4075 12614 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/A
flabel locali 13040 -4143 13074 -4109 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/Y
flabel locali 12948 -4075 12982 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/A
flabel locali 12856 -4075 12890 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/A
flabel locali 13040 -4075 13074 -4041 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_3/Y
flabel pwell 12488 -3837 12522 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_3/VNB
flabel nwell 12488 -4381 12522 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_3/VPB
flabel metal1 12488 -4381 12522 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_3/VPWR
flabel metal1 12488 -3837 12522 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_3/VGND
rlabel comment 12459 -3820 12459 -3820 2 sky130_fd_sc_hd__clkinv_4_3/clkinv_4
rlabel metal1 12459 -3868 13103 -3772 5 sky130_fd_sc_hd__clkinv_4_3/VGND
rlabel metal1 12459 -4412 13103 -4316 5 sky130_fd_sc_hd__clkinv_4_3/VPWR
flabel metal1 13224 -3837 13258 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_83/VGND
flabel metal1 13224 -4381 13258 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_83/VPWR
flabel nwell 13224 -4381 13258 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_83/VPB
flabel pwell 13224 -3837 13258 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_83/VNB
rlabel comment 13195 -3820 13195 -3820 2 sky130_fd_sc_hd__decap_4_83/decap_4
rlabel metal1 13195 -3868 13563 -3772 5 sky130_fd_sc_hd__decap_4_83/VGND
rlabel metal1 13195 -4412 13563 -4316 5 sky130_fd_sc_hd__decap_4_83/VPWR
flabel metal1 12389 -4373 12442 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_166/VPWR
flabel metal1 12388 -3840 12439 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_166/VGND
rlabel comment 12367 -3820 12367 -3820 2 sky130_fd_sc_hd__tapvpwrvgnd_1_166/tapvpwrvgnd_1
rlabel metal1 12367 -3868 12459 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_166/VGND
rlabel metal1 12367 -4412 12459 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_166/VPWR
flabel metal1 13585 -4373 13638 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_167/VPWR
flabel metal1 13584 -3840 13635 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_167/VGND
rlabel comment 13563 -3820 13563 -3820 2 sky130_fd_sc_hd__tapvpwrvgnd_1_167/tapvpwrvgnd_1
rlabel metal1 13563 -3868 13655 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_167/VGND
rlabel metal1 13563 -4412 13655 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_167/VPWR
flabel metal1 13125 -4373 13178 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_168/VPWR
flabel metal1 13124 -3840 13175 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_168/VGND
rlabel comment 13103 -3820 13103 -3820 2 sky130_fd_sc_hd__tapvpwrvgnd_1_168/tapvpwrvgnd_1
rlabel metal1 13103 -3868 13195 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_168/VGND
rlabel metal1 13103 -4412 13195 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_168/VPWR
flabel metal1 15616 -3837 15650 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_11/VGND
flabel metal1 15616 -4381 15650 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_11/VPWR
flabel nwell 15616 -4381 15650 -4347 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_11/VPB
flabel pwell 15616 -3837 15650 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_11/VNB
rlabel comment 15587 -3820 15587 -3820 2 sky130_fd_sc_hd__decap_12_11/decap_12
rlabel metal1 15587 -3868 16691 -3772 5 sky130_fd_sc_hd__decap_12_11/VGND
rlabel metal1 15587 -4412 16691 -4316 5 sky130_fd_sc_hd__decap_12_11/VPWR
flabel metal1 15517 -4373 15570 -4344 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_169/VPWR
flabel metal1 15516 -3840 15567 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_169/VGND
rlabel comment 15495 -3820 15495 -3820 2 sky130_fd_sc_hd__tapvpwrvgnd_1_169/tapvpwrvgnd_1
rlabel metal1 15495 -3868 15587 -3772 5 sky130_fd_sc_hd__tapvpwrvgnd_1_169/VGND
rlabel metal1 15495 -4412 15587 -4316 5 sky130_fd_sc_hd__tapvpwrvgnd_1_169/VPWR
flabel metal1 -2239 -3296 -2186 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_537/VPWR
flabel metal1 -2240 -3838 -2189 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_537/VGND
rlabel comment -2261 -3820 -2261 -3820 4 sky130_fd_sc_hd__tapvpwrvgnd_1_537/tapvpwrvgnd_1
rlabel metal1 -2261 -3868 -2169 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_537/VGND
rlabel metal1 -2261 -3324 -2169 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_537/VPWR
flabel metal1 -2244 -3285 -2191 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_536/VPWR
flabel metal1 -2241 -2752 -2190 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_536/VGND
rlabel comment -2169 -2732 -2169 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_536/tapvpwrvgnd_1
rlabel metal1 -2261 -2780 -2169 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_536/VGND
rlabel metal1 -2261 -3324 -2169 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_536/VPWR
flabel metal1 -2968 -3293 -2934 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_72/VPWR
flabel metal1 -2968 -3837 -2934 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_72/VGND
flabel nwell -2968 -3293 -2934 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_72/VPB
flabel pwell -2968 -3837 -2934 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_72/VNB
rlabel comment -2997 -3820 -2997 -3820 4 sky130_fd_sc_hd__decap_8_72/decap_8
rlabel metal1 -2997 -3868 -2261 -3772 1 sky130_fd_sc_hd__decap_8_72/VGND
rlabel metal1 -2997 -3324 -2261 -3228 1 sky130_fd_sc_hd__decap_8_72/VPWR
flabel metal1 -2324 -3293 -2290 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_71/VPWR
flabel metal1 -2324 -2749 -2290 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_71/VGND
flabel nwell -2324 -3293 -2290 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_71/VPB
flabel pwell -2324 -2749 -2290 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_71/VNB
rlabel comment -2261 -2732 -2261 -2732 8 sky130_fd_sc_hd__decap_8_71/decap_8
rlabel metal1 -2997 -2780 -2261 -2684 5 sky130_fd_sc_hd__decap_8_71/VGND
rlabel metal1 -2997 -3324 -2261 -3228 5 sky130_fd_sc_hd__decap_8_71/VPWR
flabel metal1 -1692 -3285 -1639 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_522/VPWR
flabel metal1 -1689 -2752 -1638 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_522/VGND
rlabel comment -1617 -2732 -1617 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_522/tapvpwrvgnd_1
rlabel metal1 -1709 -2780 -1617 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_522/VGND
rlabel metal1 -1709 -3324 -1617 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_522/VPWR
flabel metal1 -2135 -3830 -2112 -3811 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_22/VGND
flabel metal1 -2135 -3285 -2115 -3268 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_22/VPWR
flabel nwell -2134 -3290 -2109 -3264 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_22/VPB
flabel pwell -2134 -3832 -2112 -3808 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_22/VNB
rlabel comment -2169 -3820 -2169 -3820 4 sky130_fd_sc_hd__fill_4_22/fill_4
rlabel metal1 -2169 -3868 -1801 -3772 1 sky130_fd_sc_hd__fill_4_22/VGND
rlabel metal1 -2169 -3324 -1801 -3228 1 sky130_fd_sc_hd__fill_4_22/VPWR
flabel metal1 -1781 -3834 -1728 -3802 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_9/VGND
flabel metal1 -1780 -3290 -1728 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_9/VPWR
flabel nwell -1773 -3285 -1739 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_9/VPB
flabel pwell -1770 -3830 -1738 -3808 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_9/VNB
rlabel comment -1801 -3820 -1801 -3820 4 sky130_fd_sc_hd__fill_2_9/fill_2
rlabel metal1 -1801 -3868 -1617 -3772 1 sky130_fd_sc_hd__fill_2_9/VGND
rlabel metal1 -1801 -3324 -1617 -3228 1 sky130_fd_sc_hd__fill_2_9/VPWR
flabel metal1 -2058 -2750 -2005 -2718 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_8/VGND
flabel metal1 -2058 -3293 -2006 -3262 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_8/VPWR
flabel nwell -2047 -3285 -2013 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_8/VPB
flabel pwell -2048 -2744 -2016 -2722 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_8/VNB
rlabel comment -1985 -2732 -1985 -2732 8 sky130_fd_sc_hd__fill_2_8/fill_2
rlabel metal1 -2169 -2780 -1985 -2684 5 sky130_fd_sc_hd__fill_2_8/VGND
rlabel metal1 -2169 -3324 -1985 -3228 5 sky130_fd_sc_hd__fill_2_8/VPWR
flabel metal1 -944 -3293 -910 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_11/VPWR
flabel metal1 -944 -3837 -910 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_11/VGND
flabel nwell -944 -3293 -910 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_11/VPB
flabel pwell -944 -3837 -910 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_11/VNB
rlabel comment -881 -3820 -881 -3820 6 sky130_fd_sc_hd__decap_8_11/decap_8
rlabel metal1 -1617 -3868 -881 -3772 1 sky130_fd_sc_hd__decap_8_11/VGND
rlabel metal1 -1617 -3324 -881 -3228 1 sky130_fd_sc_hd__decap_8_11/VPWR
flabel metal1 -944 -3293 -910 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_7/VPWR
flabel metal1 -944 -2749 -910 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_7/VGND
flabel nwell -944 -3293 -910 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_7/VPB
flabel pwell -944 -2749 -910 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_7/VNB
rlabel comment -881 -2732 -881 -2732 8 sky130_fd_sc_hd__decap_8_7/decap_8
rlabel metal1 -1617 -2780 -881 -2684 5 sky130_fd_sc_hd__decap_8_7/VGND
rlabel metal1 -1617 -3324 -881 -3228 5 sky130_fd_sc_hd__decap_8_7/VPWR
flabel locali -1772 -2919 -1738 -2885 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/Y
flabel locali -1772 -2987 -1738 -2953 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/Y
flabel locali -1864 -3055 -1830 -3021 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/Y
flabel locali -1864 -2987 -1830 -2953 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/Y
flabel locali -1864 -2919 -1830 -2885 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/Y
flabel locali -1956 -2851 -1922 -2817 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/A
flabel locali -1956 -2919 -1922 -2885 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/A
flabel locali -1956 -2987 -1922 -2953 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_5/A
flabel nwell -1956 -3293 -1922 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_5/VPB
flabel pwell -1956 -2749 -1922 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_5/VNB
flabel metal1 -1956 -2749 -1922 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_5/VGND
flabel metal1 -1956 -3293 -1922 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_5/VPWR
rlabel comment -1985 -2732 -1985 -2732 2 sky130_fd_sc_hd__clkinv_1_5/clkinv_1
rlabel metal1 -1985 -2780 -1709 -2684 5 sky130_fd_sc_hd__clkinv_1_5/VGND
rlabel metal1 -1985 -3324 -1709 -3228 5 sky130_fd_sc_hd__clkinv_1_5/VPWR
flabel metal1 -208 -3293 -174 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_12/VPWR
flabel metal1 -208 -3837 -174 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_12/VGND
flabel nwell -208 -3293 -174 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_12/VPB
flabel pwell -208 -3837 -174 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_12/VNB
rlabel comment -145 -3820 -145 -3820 6 sky130_fd_sc_hd__decap_8_12/decap_8
rlabel metal1 -881 -3868 -145 -3772 1 sky130_fd_sc_hd__decap_8_12/VGND
rlabel metal1 -881 -3324 -145 -3228 1 sky130_fd_sc_hd__decap_8_12/VPWR
flabel metal1 -208 -3293 -174 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_8/VPWR
flabel metal1 -208 -2749 -174 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_8/VGND
flabel nwell -208 -3293 -174 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_8/VPB
flabel pwell -208 -2749 -174 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_8/VNB
rlabel comment -145 -2732 -145 -2732 8 sky130_fd_sc_hd__decap_8_8/decap_8
rlabel metal1 -881 -2780 -145 -2684 5 sky130_fd_sc_hd__decap_8_8/VGND
rlabel metal1 -881 -3324 -145 -3228 5 sky130_fd_sc_hd__decap_8_8/VPWR
flabel metal1 332 -3296 385 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_110/VPWR
flabel metal1 335 -3838 386 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_110/VGND
rlabel comment 407 -3820 407 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_110/tapvpwrvgnd_1
rlabel metal1 315 -3868 407 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_110/VGND
rlabel metal1 315 -3324 407 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_110/VPWR
flabel metal1 -128 -3296 -75 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_109/VPWR
flabel metal1 -125 -3838 -74 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_109/VGND
rlabel comment -53 -3820 -53 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_109/tapvpwrvgnd_1
rlabel metal1 -145 -3868 -53 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_109/VGND
rlabel metal1 -145 -3324 -53 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_109/VPWR
flabel metal1 -128 -3285 -75 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_90/VPWR
flabel metal1 -125 -2752 -74 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_90/VGND
rlabel comment -53 -2732 -53 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_90/tapvpwrvgnd_1
rlabel metal1 -145 -2780 -53 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_90/VGND
rlabel metal1 -145 -3324 -53 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_90/VPWR
flabel metal1 332 -3285 385 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_89/VPWR
flabel metal1 335 -2752 386 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_89/VGND
rlabel comment 407 -2732 407 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_89/tapvpwrvgnd_1
rlabel metal1 315 -2780 407 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_89/VGND
rlabel metal1 315 -3324 407 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_89/VPWR
flabel metal1 252 -3837 286 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_61/VGND
flabel metal1 252 -3293 286 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_61/VPWR
flabel nwell 252 -3293 286 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_61/VPB
flabel pwell 252 -3837 286 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_61/VNB
rlabel comment 315 -3820 315 -3820 6 sky130_fd_sc_hd__decap_4_61/decap_4
rlabel metal1 -53 -3868 315 -3772 1 sky130_fd_sc_hd__decap_4_61/VGND
rlabel metal1 -53 -3324 315 -3228 1 sky130_fd_sc_hd__decap_4_61/VPWR
flabel metal1 252 -2749 286 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_50/VGND
flabel metal1 252 -3293 286 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_50/VPWR
flabel nwell 252 -3293 286 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_50/VPB
flabel pwell 252 -2749 286 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_50/VNB
rlabel comment 315 -2732 315 -2732 8 sky130_fd_sc_hd__decap_4_50/decap_4
rlabel metal1 -53 -2780 315 -2684 5 sky130_fd_sc_hd__decap_4_50/VGND
rlabel metal1 -53 -3324 315 -3228 5 sky130_fd_sc_hd__decap_4_50/VPWR
flabel locali 1079 -3599 1113 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/A
flabel locali 433 -3395 467 -3361 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X
flabel locali 433 -3463 467 -3429 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X
flabel locali 433 -3531 467 -3497 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X
flabel locali 433 -3599 467 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X
flabel locali 433 -3667 467 -3633 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X
flabel locali 433 -3735 467 -3701 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/X
flabel pwell 1079 -3837 1113 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/VNB
flabel nwell 1079 -3293 1113 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/VPB
flabel metal1 1079 -3837 1113 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/VGND
flabel metal1 1079 -3293 1113 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_50/VPWR
rlabel comment 1143 -3820 1143 -3820 6 sky130_fd_sc_hd__clkdlybuf4s50_1_50/clkdlybuf4s50_1
rlabel metal1 407 -3868 1143 -3772 1 sky130_fd_sc_hd__clkdlybuf4s50_1_50/VGND
rlabel metal1 407 -3324 1143 -3228 1 sky130_fd_sc_hd__clkdlybuf4s50_1_50/VPWR
flabel locali 1079 -2987 1113 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A
flabel locali 433 -3191 467 -3157 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/X
flabel locali 433 -3123 467 -3089 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/X
flabel locali 433 -3055 467 -3021 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/X
flabel locali 433 -2987 467 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/X
flabel locali 433 -2919 467 -2885 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/X
flabel locali 433 -2851 467 -2817 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/X
flabel pwell 1079 -2749 1113 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/VNB
flabel nwell 1079 -3293 1113 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/VPB
flabel metal1 1079 -2749 1113 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/VGND
flabel metal1 1079 -3293 1113 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_39/VPWR
rlabel comment 1143 -2732 1143 -2732 8 sky130_fd_sc_hd__clkdlybuf4s50_1_39/clkdlybuf4s50_1
rlabel metal1 407 -2780 1143 -2684 5 sky130_fd_sc_hd__clkdlybuf4s50_1_39/VGND
rlabel metal1 407 -3324 1143 -3228 5 sky130_fd_sc_hd__clkdlybuf4s50_1_39/VPWR
flabel metal1 1620 -3296 1673 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_124/VPWR
flabel metal1 1623 -3838 1674 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_124/VGND
rlabel comment 1695 -3820 1695 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_124/tapvpwrvgnd_1
rlabel metal1 1603 -3868 1695 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_124/VGND
rlabel metal1 1603 -3324 1695 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_124/VPWR
flabel metal1 1160 -3296 1213 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_122/VPWR
flabel metal1 1163 -3838 1214 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_122/VGND
rlabel comment 1235 -3820 1235 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_122/tapvpwrvgnd_1
rlabel metal1 1143 -3868 1235 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_122/VGND
rlabel metal1 1143 -3324 1235 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_122/VPWR
flabel metal1 1620 -3285 1673 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_91/VPWR
flabel metal1 1623 -2752 1674 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_91/VGND
rlabel comment 1695 -2732 1695 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_91/tapvpwrvgnd_1
rlabel metal1 1603 -2780 1695 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_91/VGND
rlabel metal1 1603 -3324 1695 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_91/VPWR
flabel metal1 1160 -3285 1213 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_88/VPWR
flabel metal1 1163 -2752 1214 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_88/VGND
rlabel comment 1235 -2732 1235 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_88/tapvpwrvgnd_1
rlabel metal1 1143 -2780 1235 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_88/VGND
rlabel metal1 1143 -3324 1235 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_88/VPWR
flabel metal1 1540 -3837 1574 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_64/VGND
flabel metal1 1540 -3293 1574 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_64/VPWR
flabel nwell 1540 -3293 1574 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_64/VPB
flabel pwell 1540 -3837 1574 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_64/VNB
rlabel comment 1603 -3820 1603 -3820 6 sky130_fd_sc_hd__decap_4_64/decap_4
rlabel metal1 1235 -3868 1603 -3772 1 sky130_fd_sc_hd__decap_4_64/VGND
rlabel metal1 1235 -3324 1603 -3228 1 sky130_fd_sc_hd__decap_4_64/VPWR
flabel metal1 1540 -2749 1574 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_51/VGND
flabel metal1 1540 -3293 1574 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_51/VPWR
flabel nwell 1540 -3293 1574 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_51/VPB
flabel pwell 1540 -2749 1574 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_51/VNB
rlabel comment 1603 -2732 1603 -2732 8 sky130_fd_sc_hd__decap_4_51/decap_4
rlabel metal1 1235 -2780 1603 -2684 5 sky130_fd_sc_hd__decap_4_51/VGND
rlabel metal1 1235 -3324 1603 -3228 5 sky130_fd_sc_hd__decap_4_51/VPWR
flabel metal1 2448 -3296 2501 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_126/VPWR
flabel metal1 2451 -3838 2502 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_126/VGND
rlabel comment 2523 -3820 2523 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_126/tapvpwrvgnd_1
rlabel metal1 2431 -3868 2523 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_126/VGND
rlabel metal1 2431 -3324 2523 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_126/VPWR
flabel metal1 2448 -3285 2501 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_74/VPWR
flabel metal1 2451 -2752 2502 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_74/VGND
rlabel comment 2523 -2732 2523 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_74/tapvpwrvgnd_1
rlabel metal1 2431 -2780 2523 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_74/VGND
rlabel metal1 2431 -3324 2523 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_74/VPWR
flabel metal1 1724 -3293 1758 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_96/VPWR
flabel metal1 1724 -3837 1758 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_96/VGND
flabel nwell 1724 -3293 1758 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_96/VPB
flabel pwell 1724 -3837 1758 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_96/VNB
rlabel comment 1695 -3820 1695 -3820 4 sky130_fd_sc_hd__decap_8_96/decap_8
rlabel metal1 1695 -3868 2431 -3772 1 sky130_fd_sc_hd__decap_8_96/VGND
rlabel metal1 1695 -3324 2431 -3228 1 sky130_fd_sc_hd__decap_8_96/VPWR
flabel metal1 2368 -3293 2402 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_95/VPWR
flabel metal1 2368 -2749 2402 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_95/VGND
flabel nwell 2368 -3293 2402 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_95/VPB
flabel pwell 2368 -2749 2402 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_95/VNB
rlabel comment 2431 -2732 2431 -2732 8 sky130_fd_sc_hd__decap_8_95/decap_8
rlabel metal1 1695 -2780 2431 -2684 5 sky130_fd_sc_hd__decap_8_95/VGND
rlabel metal1 1695 -3324 2431 -3228 5 sky130_fd_sc_hd__decap_8_95/VPWR
flabel metal1 2828 -3837 2862 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_65/VGND
flabel metal1 2828 -3293 2862 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_65/VPWR
flabel nwell 2828 -3293 2862 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_65/VPB
flabel pwell 2828 -3837 2862 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_65/VNB
rlabel comment 2891 -3820 2891 -3820 6 sky130_fd_sc_hd__decap_4_65/decap_4
rlabel metal1 2523 -3868 2891 -3772 1 sky130_fd_sc_hd__decap_4_65/VGND
rlabel metal1 2523 -3324 2891 -3228 1 sky130_fd_sc_hd__decap_4_65/VPWR
flabel metal1 2828 -2749 2862 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_42/VGND
flabel metal1 2828 -3293 2862 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_42/VPWR
flabel nwell 2828 -3293 2862 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_42/VPB
flabel pwell 2828 -2749 2862 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_42/VNB
rlabel comment 2891 -2732 2891 -2732 8 sky130_fd_sc_hd__decap_4_42/decap_4
rlabel metal1 2523 -2780 2891 -2684 5 sky130_fd_sc_hd__decap_4_42/VGND
rlabel metal1 2523 -3324 2891 -3228 5 sky130_fd_sc_hd__decap_4_42/VPWR
flabel metal1 2908 -3296 2961 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_127/VPWR
flabel metal1 2911 -3838 2962 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_127/VGND
rlabel comment 2983 -3820 2983 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_127/tapvpwrvgnd_1
rlabel metal1 2891 -3868 2983 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_127/VGND
rlabel metal1 2891 -3324 2983 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_127/VPWR
flabel metal1 2908 -3285 2961 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_75/VPWR
flabel metal1 2911 -2752 2962 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_75/VGND
rlabel comment 2983 -2732 2983 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_75/tapvpwrvgnd_1
rlabel metal1 2891 -2780 2983 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_75/VGND
rlabel metal1 2891 -3324 2983 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_75/VPWR
flabel locali 3655 -3599 3689 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/A
flabel locali 3009 -3395 3043 -3361 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
flabel locali 3009 -3463 3043 -3429 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
flabel locali 3009 -3531 3043 -3497 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
flabel locali 3009 -3599 3043 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
flabel locali 3009 -3667 3043 -3633 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
flabel locali 3009 -3735 3043 -3701 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
flabel pwell 3655 -3837 3689 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/VNB
flabel nwell 3655 -3293 3689 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/VPB
flabel metal1 3655 -3837 3689 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/VGND
flabel metal1 3655 -3293 3689 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_52/VPWR
rlabel comment 3719 -3820 3719 -3820 6 sky130_fd_sc_hd__clkdlybuf4s50_1_52/clkdlybuf4s50_1
rlabel metal1 2983 -3868 3719 -3772 1 sky130_fd_sc_hd__clkdlybuf4s50_1_52/VGND
rlabel metal1 2983 -3324 3719 -3228 1 sky130_fd_sc_hd__clkdlybuf4s50_1_52/VPWR
flabel locali 3655 -2987 3689 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/A
flabel locali 3009 -3191 3043 -3157 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X
flabel locali 3009 -3123 3043 -3089 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X
flabel locali 3009 -3055 3043 -3021 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X
flabel locali 3009 -2987 3043 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X
flabel locali 3009 -2919 3043 -2885 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X
flabel locali 3009 -2851 3043 -2817 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/X
flabel pwell 3655 -2749 3689 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/VNB
flabel nwell 3655 -3293 3689 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/VPB
flabel metal1 3655 -2749 3689 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/VGND
flabel metal1 3655 -3293 3689 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_32/VPWR
rlabel comment 3719 -2732 3719 -2732 8 sky130_fd_sc_hd__clkdlybuf4s50_1_32/clkdlybuf4s50_1
rlabel metal1 2983 -2780 3719 -2684 5 sky130_fd_sc_hd__clkdlybuf4s50_1_32/VGND
rlabel metal1 2983 -3324 3719 -3228 5 sky130_fd_sc_hd__clkdlybuf4s50_1_32/VPWR
flabel metal1 4196 -3296 4249 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_134/VPWR
flabel metal1 4199 -3838 4250 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_134/VGND
rlabel comment 4271 -3820 4271 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_134/tapvpwrvgnd_1
rlabel metal1 4179 -3868 4271 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_134/VGND
rlabel metal1 4179 -3324 4271 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_134/VPWR
flabel metal1 3736 -3296 3789 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_129/VPWR
flabel metal1 3739 -3838 3790 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_129/VGND
rlabel comment 3811 -3820 3811 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_129/tapvpwrvgnd_1
rlabel metal1 3719 -3868 3811 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_129/VGND
rlabel metal1 3719 -3324 3811 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_129/VPWR
flabel metal1 4196 -3285 4249 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_77/VPWR
flabel metal1 4199 -2752 4250 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_77/VGND
rlabel comment 4271 -2732 4271 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_77/tapvpwrvgnd_1
rlabel metal1 4179 -2780 4271 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_77/VGND
rlabel metal1 4179 -3324 4271 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_77/VPWR
flabel metal1 3736 -3285 3789 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_76/VPWR
flabel metal1 3739 -2752 3790 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_76/VGND
rlabel comment 3811 -2732 3811 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_76/tapvpwrvgnd_1
rlabel metal1 3719 -2780 3811 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_76/VGND
rlabel metal1 3719 -3324 3811 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_76/VPWR
flabel metal1 4944 -3293 4978 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_106/VPWR
flabel metal1 4944 -2749 4978 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_106/VGND
flabel nwell 4944 -3293 4978 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_106/VPB
flabel pwell 4944 -2749 4978 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_106/VNB
rlabel comment 5007 -2732 5007 -2732 8 sky130_fd_sc_hd__decap_8_106/decap_8
rlabel metal1 4271 -2780 5007 -2684 5 sky130_fd_sc_hd__decap_8_106/VGND
rlabel metal1 4271 -3324 5007 -3228 5 sky130_fd_sc_hd__decap_8_106/VPWR
flabel metal1 4300 -3293 4334 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_104/VPWR
flabel metal1 4300 -3837 4334 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_104/VGND
flabel nwell 4300 -3293 4334 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_104/VPB
flabel pwell 4300 -3837 4334 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_104/VNB
rlabel comment 4271 -3820 4271 -3820 4 sky130_fd_sc_hd__decap_8_104/decap_8
rlabel metal1 4271 -3868 5007 -3772 1 sky130_fd_sc_hd__decap_8_104/VGND
rlabel metal1 4271 -3324 5007 -3228 1 sky130_fd_sc_hd__decap_8_104/VPWR
flabel metal1 4116 -3837 4150 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_66/VGND
flabel metal1 4116 -3293 4150 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_66/VPWR
flabel nwell 4116 -3293 4150 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_66/VPB
flabel pwell 4116 -3837 4150 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_66/VNB
rlabel comment 4179 -3820 4179 -3820 6 sky130_fd_sc_hd__decap_4_66/decap_4
rlabel metal1 3811 -3868 4179 -3772 1 sky130_fd_sc_hd__decap_4_66/VGND
rlabel metal1 3811 -3324 4179 -3228 1 sky130_fd_sc_hd__decap_4_66/VPWR
flabel metal1 4116 -2749 4150 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_43/VGND
flabel metal1 4116 -3293 4150 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_43/VPWR
flabel nwell 4116 -3293 4150 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_43/VPB
flabel pwell 4116 -2749 4150 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_43/VNB
rlabel comment 4179 -2732 4179 -2732 8 sky130_fd_sc_hd__decap_4_43/decap_4
rlabel metal1 3811 -2780 4179 -2684 5 sky130_fd_sc_hd__decap_4_43/VGND
rlabel metal1 3811 -3324 4179 -3228 5 sky130_fd_sc_hd__decap_4_43/VPWR
flabel metal1 5484 -3296 5537 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_136/VPWR
flabel metal1 5487 -3838 5538 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_136/VGND
rlabel comment 5559 -3820 5559 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_136/tapvpwrvgnd_1
rlabel metal1 5467 -3868 5559 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_136/VGND
rlabel metal1 5467 -3324 5559 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_136/VPWR
flabel metal1 5024 -3296 5077 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_135/VPWR
flabel metal1 5027 -3838 5078 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_135/VGND
rlabel comment 5099 -3820 5099 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_135/tapvpwrvgnd_1
rlabel metal1 5007 -3868 5099 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_135/VGND
rlabel metal1 5007 -3324 5099 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_135/VPWR
flabel metal1 5024 -3285 5077 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_79/VPWR
flabel metal1 5027 -2752 5078 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_79/VGND
rlabel comment 5099 -2732 5099 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_79/tapvpwrvgnd_1
rlabel metal1 5007 -2780 5099 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_79/VGND
rlabel metal1 5007 -3324 5099 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_79/VPWR
flabel metal1 5484 -3285 5537 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_78/VPWR
flabel metal1 5487 -2752 5538 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_78/VGND
rlabel comment 5559 -2732 5559 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_78/tapvpwrvgnd_1
rlabel metal1 5467 -2780 5559 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_78/VGND
rlabel metal1 5467 -3324 5559 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_78/VPWR
flabel metal1 5404 -3837 5438 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_67/VGND
flabel metal1 5404 -3293 5438 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_67/VPWR
flabel nwell 5404 -3293 5438 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_67/VPB
flabel pwell 5404 -3837 5438 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_67/VNB
rlabel comment 5467 -3820 5467 -3820 6 sky130_fd_sc_hd__decap_4_67/decap_4
rlabel metal1 5099 -3868 5467 -3772 1 sky130_fd_sc_hd__decap_4_67/VGND
rlabel metal1 5099 -3324 5467 -3228 1 sky130_fd_sc_hd__decap_4_67/VPWR
flabel metal1 5404 -2749 5438 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_44/VGND
flabel metal1 5404 -3293 5438 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_44/VPWR
flabel nwell 5404 -3293 5438 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_44/VPB
flabel pwell 5404 -2749 5438 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_44/VNB
rlabel comment 5467 -2732 5467 -2732 8 sky130_fd_sc_hd__decap_4_44/decap_4
rlabel metal1 5099 -2780 5467 -2684 5 sky130_fd_sc_hd__decap_4_44/VGND
rlabel metal1 5099 -3324 5467 -3228 5 sky130_fd_sc_hd__decap_4_44/VPWR
flabel metal1 6312 -3296 6365 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_137/VPWR
flabel metal1 6315 -3838 6366 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_137/VGND
rlabel comment 6387 -3820 6387 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_137/tapvpwrvgnd_1
rlabel metal1 6295 -3868 6387 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_137/VGND
rlabel metal1 6295 -3324 6387 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_137/VPWR
flabel metal1 6312 -3285 6365 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_80/VPWR
flabel metal1 6315 -2752 6366 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_80/VGND
rlabel comment 6387 -2732 6387 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_80/tapvpwrvgnd_1
rlabel metal1 6295 -2780 6387 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_80/VGND
rlabel metal1 6295 -3324 6387 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_80/VPWR
flabel locali 6231 -3599 6265 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/A
flabel locali 5585 -3395 5619 -3361 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X
flabel locali 5585 -3463 5619 -3429 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X
flabel locali 5585 -3531 5619 -3497 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X
flabel locali 5585 -3599 5619 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X
flabel locali 5585 -3667 5619 -3633 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X
flabel locali 5585 -3735 5619 -3701 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X
flabel pwell 6231 -3837 6265 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/VNB
flabel nwell 6231 -3293 6265 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/VPB
flabel metal1 6231 -3837 6265 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/VGND
flabel metal1 6231 -3293 6265 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_54/VPWR
rlabel comment 6295 -3820 6295 -3820 6 sky130_fd_sc_hd__clkdlybuf4s50_1_54/clkdlybuf4s50_1
rlabel metal1 5559 -3868 6295 -3772 1 sky130_fd_sc_hd__clkdlybuf4s50_1_54/VGND
rlabel metal1 5559 -3324 6295 -3228 1 sky130_fd_sc_hd__clkdlybuf4s50_1_54/VPWR
flabel locali 6231 -2987 6265 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/A
flabel locali 5585 -3191 5619 -3157 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X
flabel locali 5585 -3123 5619 -3089 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X
flabel locali 5585 -3055 5619 -3021 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X
flabel locali 5585 -2987 5619 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X
flabel locali 5585 -2919 5619 -2885 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X
flabel locali 5585 -2851 5619 -2817 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X
flabel pwell 6231 -2749 6265 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/VNB
flabel nwell 6231 -3293 6265 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/VPB
flabel metal1 6231 -2749 6265 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/VGND
flabel metal1 6231 -3293 6265 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_34/VPWR
rlabel comment 6295 -2732 6295 -2732 8 sky130_fd_sc_hd__clkdlybuf4s50_1_34/clkdlybuf4s50_1
rlabel metal1 5559 -2780 6295 -2684 5 sky130_fd_sc_hd__clkdlybuf4s50_1_34/VGND
rlabel metal1 5559 -3324 6295 -3228 5 sky130_fd_sc_hd__clkdlybuf4s50_1_34/VPWR
flabel metal1 6692 -3837 6726 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_68/VGND
flabel metal1 6692 -3293 6726 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_68/VPWR
flabel nwell 6692 -3293 6726 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_68/VPB
flabel pwell 6692 -3837 6726 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_68/VNB
rlabel comment 6755 -3820 6755 -3820 6 sky130_fd_sc_hd__decap_4_68/decap_4
rlabel metal1 6387 -3868 6755 -3772 1 sky130_fd_sc_hd__decap_4_68/VGND
rlabel metal1 6387 -3324 6755 -3228 1 sky130_fd_sc_hd__decap_4_68/VPWR
flabel metal1 6692 -2749 6726 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_45/VGND
flabel metal1 6692 -3293 6726 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_45/VPWR
flabel nwell 6692 -3293 6726 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_45/VPB
flabel pwell 6692 -2749 6726 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_45/VNB
rlabel comment 6755 -2732 6755 -2732 8 sky130_fd_sc_hd__decap_4_45/decap_4
rlabel metal1 6387 -2780 6755 -2684 5 sky130_fd_sc_hd__decap_4_45/VGND
rlabel metal1 6387 -3324 6755 -3228 5 sky130_fd_sc_hd__decap_4_45/VPWR
flabel metal1 6772 -3296 6825 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_138/VPWR
flabel metal1 6775 -3838 6826 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_138/VGND
rlabel comment 6847 -3820 6847 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_138/tapvpwrvgnd_1
rlabel metal1 6755 -3868 6847 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_138/VGND
rlabel metal1 6755 -3324 6847 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_138/VPWR
flabel metal1 6772 -3285 6825 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_81/VPWR
flabel metal1 6775 -2752 6826 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_81/VGND
rlabel comment 6847 -2732 6847 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_81/tapvpwrvgnd_1
rlabel metal1 6755 -2780 6847 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_81/VGND
rlabel metal1 6755 -3324 6847 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_81/VPWR
flabel metal1 6876 -3293 6910 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_116/VPWR
flabel metal1 6876 -3837 6910 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_116/VGND
flabel nwell 6876 -3293 6910 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_116/VPB
flabel pwell 6876 -3837 6910 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_116/VNB
rlabel comment 6847 -3820 6847 -3820 4 sky130_fd_sc_hd__decap_8_116/decap_8
rlabel metal1 6847 -3868 7583 -3772 1 sky130_fd_sc_hd__decap_8_116/VGND
rlabel metal1 6847 -3324 7583 -3228 1 sky130_fd_sc_hd__decap_8_116/VPWR
flabel metal1 7520 -3293 7554 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_115/VPWR
flabel metal1 7520 -2749 7554 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_115/VGND
flabel nwell 7520 -3293 7554 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_115/VPB
flabel pwell 7520 -2749 7554 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_115/VNB
rlabel comment 7583 -2732 7583 -2732 8 sky130_fd_sc_hd__decap_8_115/decap_8
rlabel metal1 6847 -2780 7583 -2684 5 sky130_fd_sc_hd__decap_8_115/VGND
rlabel metal1 6847 -3324 7583 -3228 5 sky130_fd_sc_hd__decap_8_115/VPWR
flabel metal1 8060 -3296 8113 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_140/VPWR
flabel metal1 8063 -3838 8114 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_140/VGND
rlabel comment 8135 -3820 8135 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_140/tapvpwrvgnd_1
rlabel metal1 8043 -3868 8135 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_140/VGND
rlabel metal1 8043 -3324 8135 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_140/VPWR
flabel metal1 7600 -3296 7653 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_139/VPWR
flabel metal1 7603 -3838 7654 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_139/VGND
rlabel comment 7675 -3820 7675 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_139/tapvpwrvgnd_1
rlabel metal1 7583 -3868 7675 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_139/VGND
rlabel metal1 7583 -3324 7675 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_139/VPWR
flabel metal1 8060 -3285 8113 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_83/VPWR
flabel metal1 8063 -2752 8114 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_83/VGND
rlabel comment 8135 -2732 8135 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_83/tapvpwrvgnd_1
rlabel metal1 8043 -2780 8135 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_83/VGND
rlabel metal1 8043 -3324 8135 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_83/VPWR
flabel metal1 7600 -3285 7653 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_82/VPWR
flabel metal1 7603 -2752 7654 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_82/VGND
rlabel comment 7675 -2732 7675 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_82/tapvpwrvgnd_1
rlabel metal1 7583 -2780 7675 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_82/VGND
rlabel metal1 7583 -3324 7675 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_82/VPWR
flabel metal1 7980 -3837 8014 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_69/VGND
flabel metal1 7980 -3293 8014 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_69/VPWR
flabel nwell 7980 -3293 8014 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_69/VPB
flabel pwell 7980 -3837 8014 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_69/VNB
rlabel comment 8043 -3820 8043 -3820 6 sky130_fd_sc_hd__decap_4_69/decap_4
rlabel metal1 7675 -3868 8043 -3772 1 sky130_fd_sc_hd__decap_4_69/VGND
rlabel metal1 7675 -3324 8043 -3228 1 sky130_fd_sc_hd__decap_4_69/VPWR
flabel metal1 7980 -2749 8014 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_46/VGND
flabel metal1 7980 -3293 8014 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_46/VPWR
flabel nwell 7980 -3293 8014 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_46/VPB
flabel pwell 7980 -2749 8014 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_46/VNB
rlabel comment 8043 -2732 8043 -2732 8 sky130_fd_sc_hd__decap_4_46/decap_4
rlabel metal1 7675 -2780 8043 -2684 5 sky130_fd_sc_hd__decap_4_46/VGND
rlabel metal1 7675 -3324 8043 -3228 5 sky130_fd_sc_hd__decap_4_46/VPWR
flabel locali 8807 -3599 8841 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/A
flabel locali 8161 -3395 8195 -3361 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X
flabel locali 8161 -3463 8195 -3429 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X
flabel locali 8161 -3531 8195 -3497 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X
flabel locali 8161 -3599 8195 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X
flabel locali 8161 -3667 8195 -3633 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X
flabel locali 8161 -3735 8195 -3701 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X
flabel pwell 8807 -3837 8841 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/VNB
flabel nwell 8807 -3293 8841 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/VPB
flabel metal1 8807 -3837 8841 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/VGND
flabel metal1 8807 -3293 8841 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_56/VPWR
rlabel comment 8871 -3820 8871 -3820 6 sky130_fd_sc_hd__clkdlybuf4s50_1_56/clkdlybuf4s50_1
rlabel metal1 8135 -3868 8871 -3772 1 sky130_fd_sc_hd__clkdlybuf4s50_1_56/VGND
rlabel metal1 8135 -3324 8871 -3228 1 sky130_fd_sc_hd__clkdlybuf4s50_1_56/VPWR
flabel locali 8807 -2987 8841 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/A
flabel locali 8161 -3191 8195 -3157 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
flabel locali 8161 -3123 8195 -3089 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
flabel locali 8161 -3055 8195 -3021 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
flabel locali 8161 -2987 8195 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
flabel locali 8161 -2919 8195 -2885 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
flabel locali 8161 -2851 8195 -2817 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
flabel pwell 8807 -2749 8841 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/VNB
flabel nwell 8807 -3293 8841 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/VPB
flabel metal1 8807 -2749 8841 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/VGND
flabel metal1 8807 -3293 8841 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_36/VPWR
rlabel comment 8871 -2732 8871 -2732 8 sky130_fd_sc_hd__clkdlybuf4s50_1_36/clkdlybuf4s50_1
rlabel metal1 8135 -2780 8871 -2684 5 sky130_fd_sc_hd__clkdlybuf4s50_1_36/VGND
rlabel metal1 8135 -3324 8871 -3228 5 sky130_fd_sc_hd__clkdlybuf4s50_1_36/VPWR
flabel metal1 8888 -3296 8941 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_142/VPWR
flabel metal1 8891 -3838 8942 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_142/VGND
rlabel comment 8963 -3820 8963 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_142/tapvpwrvgnd_1
rlabel metal1 8871 -3868 8963 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_142/VGND
rlabel metal1 8871 -3324 8963 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_142/VPWR
flabel metal1 8888 -3285 8941 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_84/VPWR
flabel metal1 8891 -2752 8942 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_84/VGND
rlabel comment 8963 -2732 8963 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_84/tapvpwrvgnd_1
rlabel metal1 8871 -2780 8963 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_84/VGND
rlabel metal1 8871 -3324 8963 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_84/VPWR
flabel metal1 9268 -3837 9302 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_70/VGND
flabel metal1 9268 -3293 9302 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_70/VPWR
flabel nwell 9268 -3293 9302 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_70/VPB
flabel pwell 9268 -3837 9302 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_70/VNB
rlabel comment 9331 -3820 9331 -3820 6 sky130_fd_sc_hd__decap_4_70/decap_4
rlabel metal1 8963 -3868 9331 -3772 1 sky130_fd_sc_hd__decap_4_70/VGND
rlabel metal1 8963 -3324 9331 -3228 1 sky130_fd_sc_hd__decap_4_70/VPWR
flabel metal1 9268 -2749 9302 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_47/VGND
flabel metal1 9268 -3293 9302 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_47/VPWR
flabel nwell 9268 -3293 9302 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_47/VPB
flabel pwell 9268 -2749 9302 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_47/VNB
rlabel comment 9331 -2732 9331 -2732 8 sky130_fd_sc_hd__decap_4_47/decap_4
rlabel metal1 8963 -2780 9331 -2684 5 sky130_fd_sc_hd__decap_4_47/VGND
rlabel metal1 8963 -3324 9331 -3228 5 sky130_fd_sc_hd__decap_4_47/VPWR
flabel metal1 9348 -3296 9401 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_141/VPWR
flabel metal1 9351 -3838 9402 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_141/VGND
rlabel comment 9423 -3820 9423 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_141/tapvpwrvgnd_1
rlabel metal1 9331 -3868 9423 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_141/VGND
rlabel metal1 9331 -3324 9423 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_141/VPWR
flabel metal1 9348 -3285 9401 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_85/VPWR
flabel metal1 9351 -2752 9402 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_85/VGND
rlabel comment 9423 -2732 9423 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_85/tapvpwrvgnd_1
rlabel metal1 9331 -2780 9423 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_85/VGND
rlabel metal1 9331 -3324 9423 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_85/VPWR
flabel metal1 9452 -3293 9486 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_126/VPWR
flabel metal1 9452 -3837 9486 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_126/VGND
flabel nwell 9452 -3293 9486 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_126/VPB
flabel pwell 9452 -3837 9486 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_126/VNB
rlabel comment 9423 -3820 9423 -3820 4 sky130_fd_sc_hd__decap_8_126/decap_8
rlabel metal1 9423 -3868 10159 -3772 1 sky130_fd_sc_hd__decap_8_126/VGND
rlabel metal1 9423 -3324 10159 -3228 1 sky130_fd_sc_hd__decap_8_126/VPWR
flabel metal1 10096 -3293 10130 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_125/VPWR
flabel metal1 10096 -2749 10130 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_125/VGND
flabel nwell 10096 -3293 10130 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_125/VPB
flabel pwell 10096 -2749 10130 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_125/VNB
rlabel comment 10159 -2732 10159 -2732 8 sky130_fd_sc_hd__decap_8_125/decap_8
rlabel metal1 9423 -2780 10159 -2684 5 sky130_fd_sc_hd__decap_8_125/VGND
rlabel metal1 9423 -3324 10159 -3228 5 sky130_fd_sc_hd__decap_8_125/VPWR
flabel metal1 10176 -3296 10229 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_143/VPWR
flabel metal1 10179 -3838 10230 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_143/VGND
rlabel comment 10251 -3820 10251 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_143/tapvpwrvgnd_1
rlabel metal1 10159 -3868 10251 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_143/VGND
rlabel metal1 10159 -3324 10251 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_143/VPWR
flabel metal1 10176 -3285 10229 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_86/VPWR
flabel metal1 10179 -2752 10230 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_86/VGND
rlabel comment 10251 -2732 10251 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_86/tapvpwrvgnd_1
rlabel metal1 10159 -2780 10251 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_86/VGND
rlabel metal1 10159 -3324 10251 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_86/VPWR
flabel metal1 10285 -3293 10321 -3263 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_18/VPWR
flabel metal1 10285 -3833 10321 -3804 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_18/VGND
flabel nwell 10292 -3286 10312 -3269 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_18/VPB
flabel pwell 10291 -3831 10315 -3809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_18/VNB
rlabel comment 10343 -3820 10343 -3820 6 sky130_fd_sc_hd__fill_1_18/fill_1
rlabel metal1 10251 -3868 10343 -3772 1 sky130_fd_sc_hd__fill_1_18/VGND
rlabel metal1 10251 -3324 10343 -3228 1 sky130_fd_sc_hd__fill_1_18/VPWR
flabel metal1 10285 -3289 10321 -3259 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_12/VPWR
flabel metal1 10285 -2748 10321 -2719 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_12/VGND
flabel nwell 10292 -3283 10312 -3266 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_12/VPB
flabel pwell 10291 -2743 10315 -2721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_12/VNB
rlabel comment 10343 -2732 10343 -2732 8 sky130_fd_sc_hd__fill_1_12/fill_1
rlabel metal1 10251 -2780 10343 -2684 5 sky130_fd_sc_hd__fill_1_12/VGND
rlabel metal1 10251 -3324 10343 -3228 5 sky130_fd_sc_hd__fill_1_12/VPWR
flabel metal1 10648 -3837 10682 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_71/VGND
flabel metal1 10648 -3293 10682 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_71/VPWR
flabel nwell 10648 -3293 10682 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_71/VPB
flabel pwell 10648 -3837 10682 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_71/VNB
rlabel comment 10711 -3820 10711 -3820 6 sky130_fd_sc_hd__decap_4_71/decap_4
rlabel metal1 10343 -3868 10711 -3772 1 sky130_fd_sc_hd__decap_4_71/VGND
rlabel metal1 10343 -3324 10711 -3228 1 sky130_fd_sc_hd__decap_4_71/VPWR
flabel metal1 10648 -2749 10682 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_48/VGND
flabel metal1 10648 -3293 10682 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_48/VPWR
flabel nwell 10648 -3293 10682 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_48/VPB
flabel pwell 10648 -2749 10682 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_48/VNB
rlabel comment 10711 -2732 10711 -2732 8 sky130_fd_sc_hd__decap_4_48/decap_4
rlabel metal1 10343 -2780 10711 -2684 5 sky130_fd_sc_hd__decap_4_48/VGND
rlabel metal1 10343 -3324 10711 -3228 5 sky130_fd_sc_hd__decap_4_48/VPWR
flabel metal1 10653 -3293 10689 -3263 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_19/VPWR
flabel metal1 10653 -3833 10689 -3804 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_19/VGND
flabel nwell 10660 -3286 10680 -3269 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_19/VPB
flabel pwell 10659 -3831 10683 -3809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_19/VNB
rlabel comment 10711 -3820 10711 -3820 6 sky130_fd_sc_hd__fill_1_19/fill_1
rlabel metal1 10619 -3868 10711 -3772 1 sky130_fd_sc_hd__fill_1_19/VGND
rlabel metal1 10619 -3324 10711 -3228 1 sky130_fd_sc_hd__fill_1_19/VPWR
flabel metal1 10653 -3289 10689 -3259 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_13/VPWR
flabel metal1 10653 -2748 10689 -2719 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_13/VGND
flabel nwell 10660 -3283 10680 -3266 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_13/VPB
flabel pwell 10659 -2743 10683 -2721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_13/VNB
rlabel comment 10711 -2732 10711 -2732 8 sky130_fd_sc_hd__fill_1_13/fill_1
rlabel metal1 10619 -2780 10711 -2684 5 sky130_fd_sc_hd__fill_1_13/VGND
rlabel metal1 10619 -3324 10711 -3228 5 sky130_fd_sc_hd__fill_1_13/VPWR
flabel locali 11383 -3599 11417 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A
flabel locali 10737 -3395 10771 -3361 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
flabel locali 10737 -3463 10771 -3429 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
flabel locali 10737 -3531 10771 -3497 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
flabel locali 10737 -3599 10771 -3565 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
flabel locali 10737 -3667 10771 -3633 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
flabel locali 10737 -3735 10771 -3701 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
flabel pwell 11383 -3837 11417 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/VNB
flabel nwell 11383 -3293 11417 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/VPB
flabel metal1 11383 -3837 11417 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/VGND
flabel metal1 11383 -3293 11417 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_58/VPWR
rlabel comment 11447 -3820 11447 -3820 6 sky130_fd_sc_hd__clkdlybuf4s50_1_58/clkdlybuf4s50_1
rlabel metal1 10711 -3868 11447 -3772 1 sky130_fd_sc_hd__clkdlybuf4s50_1_58/VGND
rlabel metal1 10711 -3324 11447 -3228 1 sky130_fd_sc_hd__clkdlybuf4s50_1_58/VPWR
flabel locali 11383 -2987 11417 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A
flabel locali 10737 -3191 10771 -3157 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X
flabel locali 10737 -3123 10771 -3089 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X
flabel locali 10737 -3055 10771 -3021 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X
flabel locali 10737 -2987 10771 -2953 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X
flabel locali 10737 -2919 10771 -2885 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X
flabel locali 10737 -2851 10771 -2817 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X
flabel pwell 11383 -2749 11417 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/VNB
flabel nwell 11383 -3293 11417 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/VPB
flabel metal1 11383 -2749 11417 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/VGND
flabel metal1 11383 -3293 11417 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_38/VPWR
rlabel comment 11447 -2732 11447 -2732 8 sky130_fd_sc_hd__clkdlybuf4s50_1_38/clkdlybuf4s50_1
rlabel metal1 10711 -2780 11447 -2684 5 sky130_fd_sc_hd__clkdlybuf4s50_1_38/VGND
rlabel metal1 10711 -3324 11447 -3228 5 sky130_fd_sc_hd__clkdlybuf4s50_1_38/VPWR
flabel metal1 11464 -3296 11517 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_144/VPWR
flabel metal1 11467 -3838 11518 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_144/VGND
rlabel comment 11539 -3820 11539 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_144/tapvpwrvgnd_1
rlabel metal1 11447 -3868 11539 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_144/VGND
rlabel metal1 11447 -3324 11539 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_144/VPWR
flabel metal1 11464 -3285 11517 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_87/VPWR
flabel metal1 11467 -2752 11518 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_87/VGND
rlabel comment 11539 -2732 11539 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_87/tapvpwrvgnd_1
rlabel metal1 11447 -2780 11539 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_87/VGND
rlabel metal1 11447 -3324 11539 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_87/VPWR
flabel metal1 12668 -3840 12700 -3810 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_9/VGND
flabel metal1 12668 -3297 12706 -3265 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_9/VPWR
flabel nwell 12658 -3298 12715 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_9/VPB
flabel pwell 12665 -3844 12709 -3810 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_9/VNB
rlabel comment 12735 -3820 12735 -3820 6 sky130_fd_sc_hd__fill_8_9/fill_8
rlabel metal1 11999 -3868 12735 -3772 1 sky130_fd_sc_hd__fill_8_9/VGND
rlabel metal1 11999 -3324 12735 -3228 1 sky130_fd_sc_hd__fill_8_9/VPWR
flabel metal1 12668 -2742 12700 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_8/VGND
flabel metal1 12668 -3287 12706 -3255 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_8/VPWR
flabel nwell 12658 -3285 12715 -3254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_8/VPB
flabel pwell 12665 -2742 12709 -2708 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_8/VNB
rlabel comment 12735 -2732 12735 -2732 8 sky130_fd_sc_hd__fill_8_8/fill_8
rlabel metal1 11999 -2780 12735 -2684 5 sky130_fd_sc_hd__fill_8_8/VGND
rlabel metal1 11999 -3324 12735 -3228 5 sky130_fd_sc_hd__fill_8_8/VPWR
flabel metal1 11573 -3293 11609 -3263 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_20/VPWR
flabel metal1 11573 -3833 11609 -3804 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_20/VGND
flabel nwell 11580 -3286 11600 -3269 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_20/VPB
flabel pwell 11579 -3831 11603 -3809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_20/VNB
rlabel comment 11631 -3820 11631 -3820 6 sky130_fd_sc_hd__fill_1_20/fill_1
rlabel metal1 11539 -3868 11631 -3772 1 sky130_fd_sc_hd__fill_1_20/VGND
rlabel metal1 11539 -3324 11631 -3228 1 sky130_fd_sc_hd__fill_1_20/VPWR
flabel metal1 11573 -3289 11609 -3259 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_14/VPWR
flabel metal1 11573 -2748 11609 -2719 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_14/VGND
flabel nwell 11580 -3283 11600 -3266 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_14/VPB
flabel pwell 11579 -2743 11603 -2721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_14/VNB
rlabel comment 11631 -2732 11631 -2732 8 sky130_fd_sc_hd__fill_1_14/fill_1
rlabel metal1 11539 -2780 11631 -2684 5 sky130_fd_sc_hd__fill_1_14/VGND
rlabel metal1 11539 -3324 11631 -3228 5 sky130_fd_sc_hd__fill_1_14/VPWR
flabel metal1 11936 -3837 11970 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_72/VGND
flabel metal1 11936 -3293 11970 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_72/VPWR
flabel nwell 11936 -3293 11970 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_72/VPB
flabel pwell 11936 -3837 11970 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_72/VNB
rlabel comment 11999 -3820 11999 -3820 6 sky130_fd_sc_hd__decap_4_72/decap_4
rlabel metal1 11631 -3868 11999 -3772 1 sky130_fd_sc_hd__decap_4_72/VGND
rlabel metal1 11631 -3324 11999 -3228 1 sky130_fd_sc_hd__decap_4_72/VPWR
flabel metal1 11936 -2749 11970 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_49/VGND
flabel metal1 11936 -3293 11970 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_49/VPWR
flabel nwell 11936 -3293 11970 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_49/VPB
flabel pwell 11936 -2749 11970 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_49/VNB
rlabel comment 11999 -2732 11999 -2732 8 sky130_fd_sc_hd__decap_4_49/decap_4
rlabel metal1 11631 -2780 11999 -2684 5 sky130_fd_sc_hd__decap_4_49/VGND
rlabel metal1 11631 -3324 11999 -3228 5 sky130_fd_sc_hd__decap_4_49/VPWR
flabel metal1 14604 -2749 14638 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_7/VGND
flabel metal1 14604 -3293 14638 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_7/VPWR
flabel nwell 14604 -3293 14638 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_7/VPB
flabel pwell 14604 -2749 14638 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_7/VNB
rlabel comment 14667 -2732 14667 -2732 8 sky130_fd_sc_hd__decap_12_7/decap_12
rlabel metal1 13563 -2780 14667 -2684 5 sky130_fd_sc_hd__decap_12_7/VGND
rlabel metal1 13563 -3324 14667 -3228 5 sky130_fd_sc_hd__decap_12_7/VPWR
flabel metal1 14604 -3837 14638 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_9/VGND
flabel metal1 14604 -3293 14638 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_9/VPWR
flabel nwell 14604 -3293 14638 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_9/VPB
flabel pwell 14604 -3837 14638 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_9/VNB
rlabel comment 14667 -3820 14667 -3820 6 sky130_fd_sc_hd__decap_12_9/decap_12
rlabel metal1 13563 -3868 14667 -3772 1 sky130_fd_sc_hd__decap_12_9/VGND
rlabel metal1 13563 -3324 14667 -3228 1 sky130_fd_sc_hd__decap_12_9/VPWR
flabel metal1 13404 -2742 13436 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_7/VGND
flabel metal1 13404 -3287 13442 -3255 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_7/VPWR
flabel nwell 13394 -3285 13451 -3254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_7/VPB
flabel pwell 13401 -2742 13445 -2708 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_7/VNB
rlabel comment 13471 -2732 13471 -2732 8 sky130_fd_sc_hd__fill_8_7/fill_8
rlabel metal1 12735 -2780 13471 -2684 5 sky130_fd_sc_hd__fill_8_7/VGND
rlabel metal1 12735 -3324 13471 -3228 5 sky130_fd_sc_hd__fill_8_7/VPWR
flabel metal1 13404 -3840 13436 -3810 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_10/VGND
flabel metal1 13404 -3297 13442 -3265 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_10/VPWR
flabel nwell 13394 -3298 13451 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_10/VPB
flabel pwell 13401 -3844 13445 -3810 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_10/VNB
rlabel comment 13471 -3820 13471 -3820 6 sky130_fd_sc_hd__fill_8_10/fill_8
rlabel metal1 12735 -3868 13471 -3772 1 sky130_fd_sc_hd__fill_8_10/VGND
rlabel metal1 12735 -3324 13471 -3228 1 sky130_fd_sc_hd__fill_8_10/VPWR
flabel metal1 13488 -3285 13541 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_131/VPWR
flabel metal1 13491 -2752 13542 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_131/VGND
rlabel comment 13563 -2732 13563 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_131/tapvpwrvgnd_1
rlabel metal1 13471 -2780 13563 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_131/VGND
rlabel metal1 13471 -3324 13563 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_131/VPWR
flabel metal1 13488 -3296 13541 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_145/VPWR
flabel metal1 13491 -3838 13542 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_145/VGND
rlabel comment 13563 -3820 13563 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_145/tapvpwrvgnd_1
rlabel metal1 13471 -3868 13563 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_145/VGND
rlabel metal1 13471 -3324 13563 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_145/VPWR
flabel metal1 16628 -3293 16662 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_10/VPWR
flabel metal1 16628 -2749 16662 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_10/VGND
flabel nwell 16628 -3293 16662 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_10/VPB
flabel pwell 16628 -2749 16662 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_10/VNB
rlabel comment 16691 -2732 16691 -2732 8 sky130_fd_sc_hd__decap_8_10/decap_8
rlabel metal1 15955 -2780 16691 -2684 5 sky130_fd_sc_hd__decap_8_10/VGND
rlabel metal1 15955 -3324 16691 -3228 5 sky130_fd_sc_hd__decap_8_10/VPWR
flabel metal1 16628 -3293 16662 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_13/VPWR
flabel metal1 16628 -3837 16662 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_13/VGND
flabel nwell 16628 -3293 16662 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_13/VPB
flabel pwell 16628 -3837 16662 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_13/VNB
rlabel comment 16691 -3820 16691 -3820 6 sky130_fd_sc_hd__decap_8_13/decap_8
rlabel metal1 15955 -3868 16691 -3772 1 sky130_fd_sc_hd__decap_8_13/VGND
rlabel metal1 15955 -3324 16691 -3228 1 sky130_fd_sc_hd__decap_8_13/VPWR
flabel metal1 15800 -2749 15834 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_8/VGND
flabel metal1 15800 -3293 15834 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_8/VPWR
flabel nwell 15800 -3293 15834 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_8/VPB
flabel pwell 15800 -2749 15834 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_8/VNB
rlabel comment 15863 -2732 15863 -2732 8 sky130_fd_sc_hd__decap_12_8/decap_12
rlabel metal1 14759 -2780 15863 -2684 5 sky130_fd_sc_hd__decap_12_8/VGND
rlabel metal1 14759 -3324 15863 -3228 5 sky130_fd_sc_hd__decap_12_8/VPWR
flabel metal1 15800 -3837 15834 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_10/VGND
flabel metal1 15800 -3293 15834 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_10/VPWR
flabel nwell 15800 -3293 15834 -3259 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_10/VPB
flabel pwell 15800 -3837 15834 -3803 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_10/VNB
rlabel comment 15863 -3820 15863 -3820 6 sky130_fd_sc_hd__decap_12_10/decap_12
rlabel metal1 14759 -3868 15863 -3772 1 sky130_fd_sc_hd__decap_12_10/VGND
rlabel metal1 14759 -3324 15863 -3228 1 sky130_fd_sc_hd__decap_12_10/VPWR
flabel metal1 14684 -3285 14737 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_132/VPWR
flabel metal1 14687 -2752 14738 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_132/VGND
rlabel comment 14759 -2732 14759 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_132/tapvpwrvgnd_1
rlabel metal1 14667 -2780 14759 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_132/VGND
rlabel metal1 14667 -3324 14759 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_132/VPWR
flabel metal1 15880 -3285 15933 -3256 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_133/VPWR
flabel metal1 15883 -2752 15934 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_133/VGND
rlabel comment 15955 -2732 15955 -2732 8 sky130_fd_sc_hd__tapvpwrvgnd_1_133/tapvpwrvgnd_1
rlabel metal1 15863 -2780 15955 -2684 5 sky130_fd_sc_hd__tapvpwrvgnd_1_133/VGND
rlabel metal1 15863 -3324 15955 -3228 5 sky130_fd_sc_hd__tapvpwrvgnd_1_133/VPWR
flabel metal1 14684 -3296 14737 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_146/VPWR
flabel metal1 14687 -3838 14738 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_146/VGND
rlabel comment 14759 -3820 14759 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_146/tapvpwrvgnd_1
rlabel metal1 14667 -3868 14759 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_146/VGND
rlabel metal1 14667 -3324 14759 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_146/VPWR
flabel metal1 15880 -3296 15933 -3267 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_147/VPWR
flabel metal1 15883 -3838 15934 -3800 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_147/VGND
rlabel comment 15955 -3820 15955 -3820 6 sky130_fd_sc_hd__tapvpwrvgnd_1_147/tapvpwrvgnd_1
rlabel metal1 15863 -3868 15955 -3772 1 sky130_fd_sc_hd__tapvpwrvgnd_1_147/VGND
rlabel metal1 15863 -3324 15955 -3228 1 sky130_fd_sc_hd__tapvpwrvgnd_1_147/VPWR
flabel metal1 -1588 -2205 -1554 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_5/VPWR
flabel metal1 -1588 -2749 -1554 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_5/VGND
flabel nwell -1588 -2205 -1554 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_5/VPB
flabel pwell -1588 -2749 -1554 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_5/VNB
rlabel comment -1617 -2732 -1617 -2732 4 sky130_fd_sc_hd__decap_8_5/decap_8
rlabel metal1 -1617 -2780 -881 -2684 1 sky130_fd_sc_hd__decap_8_5/VGND
rlabel metal1 -1617 -2236 -881 -2140 1 sky130_fd_sc_hd__decap_8_5/VPWR
flabel metal1 -2968 -2205 -2934 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_70/VPWR
flabel metal1 -2968 -2749 -2934 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_70/VGND
flabel nwell -2968 -2205 -2934 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_70/VPB
flabel pwell -2968 -2749 -2934 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_70/VNB
rlabel comment -2997 -2732 -2997 -2732 4 sky130_fd_sc_hd__decap_8_70/decap_8
rlabel metal1 -2997 -2780 -2261 -2684 1 sky130_fd_sc_hd__decap_8_70/VGND
rlabel metal1 -2997 -2236 -2261 -2140 1 sky130_fd_sc_hd__decap_8_70/VPWR
flabel metal1 -1781 -2746 -1728 -2714 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_6/VGND
flabel metal1 -1780 -2202 -1728 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_6/VPWR
flabel nwell -1773 -2197 -1739 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_6/VPB
flabel pwell -1770 -2742 -1738 -2720 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_6/VNB
rlabel comment -1801 -2732 -1801 -2732 4 sky130_fd_sc_hd__fill_2_6/fill_2
rlabel metal1 -1801 -2780 -1617 -2684 1 sky130_fd_sc_hd__fill_2_6/VGND
rlabel metal1 -1801 -2236 -1617 -2140 1 sky130_fd_sc_hd__fill_2_6/VPWR
flabel metal1 -2135 -2742 -2112 -2723 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_21/VGND
flabel metal1 -2135 -2197 -2115 -2180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_21/VPWR
flabel nwell -2134 -2202 -2109 -2176 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_21/VPB
flabel pwell -2134 -2744 -2112 -2720 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_21/VNB
rlabel comment -2169 -2732 -2169 -2732 4 sky130_fd_sc_hd__fill_4_21/fill_4
rlabel metal1 -2169 -2780 -1801 -2684 1 sky130_fd_sc_hd__fill_4_21/VGND
rlabel metal1 -2169 -2236 -1801 -2140 1 sky130_fd_sc_hd__fill_4_21/VPWR
flabel metal1 -2239 -2208 -2186 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_535/VPWR
flabel metal1 -2240 -2750 -2189 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_535/VGND
rlabel comment -2261 -2732 -2261 -2732 4 sky130_fd_sc_hd__tapvpwrvgnd_1_535/tapvpwrvgnd_1
rlabel metal1 -2261 -2780 -2169 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_535/VGND
rlabel metal1 -2261 -2236 -2169 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_535/VPWR
flabel locali 437 -2511 471 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/A
flabel locali 1083 -2307 1117 -2273 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X
flabel locali 1083 -2375 1117 -2341 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X
flabel locali 1083 -2443 1117 -2409 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X
flabel locali 1083 -2511 1117 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X
flabel locali 1083 -2579 1117 -2545 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X
flabel locali 1083 -2647 1117 -2613 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X
flabel pwell 437 -2749 471 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/VNB
flabel nwell 437 -2205 471 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/VPB
flabel metal1 437 -2749 471 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/VGND
flabel metal1 437 -2205 471 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_47/VPWR
rlabel comment 407 -2732 407 -2732 4 sky130_fd_sc_hd__clkdlybuf4s50_1_47/clkdlybuf4s50_1
rlabel metal1 407 -2780 1143 -2684 1 sky130_fd_sc_hd__clkdlybuf4s50_1_47/VGND
rlabel metal1 407 -2236 1143 -2140 1 sky130_fd_sc_hd__clkdlybuf4s50_1_47/VPWR
flabel metal1 252 -2749 286 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_58/VGND
flabel metal1 252 -2205 286 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_58/VPWR
flabel nwell 252 -2205 286 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_58/VPB
flabel pwell 252 -2749 286 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_58/VNB
rlabel comment 315 -2732 315 -2732 6 sky130_fd_sc_hd__decap_4_58/decap_4
rlabel metal1 -53 -2780 315 -2684 1 sky130_fd_sc_hd__decap_4_58/VGND
rlabel metal1 -53 -2236 315 -2140 1 sky130_fd_sc_hd__decap_4_58/VPWR
flabel metal1 -852 -2205 -818 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_6/VPWR
flabel metal1 -852 -2749 -818 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_6/VGND
flabel nwell -852 -2205 -818 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_6/VPB
flabel pwell -852 -2749 -818 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_6/VNB
rlabel comment -881 -2732 -881 -2732 4 sky130_fd_sc_hd__decap_8_6/decap_8
rlabel metal1 -881 -2780 -145 -2684 1 sky130_fd_sc_hd__decap_8_6/VGND
rlabel metal1 -881 -2236 -145 -2140 1 sky130_fd_sc_hd__decap_8_6/VPWR
flabel metal1 332 -2208 385 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_104/VPWR
flabel metal1 335 -2750 386 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_104/VGND
rlabel comment 407 -2732 407 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_104/tapvpwrvgnd_1
rlabel metal1 315 -2780 407 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_104/VGND
rlabel metal1 315 -2236 407 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_104/VPWR
flabel metal1 -128 -2208 -75 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_106/VPWR
flabel metal1 -125 -2750 -74 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_106/VGND
rlabel comment -53 -2732 -53 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_106/tapvpwrvgnd_1
rlabel metal1 -145 -2780 -53 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_106/VGND
rlabel metal1 -145 -2236 -53 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_106/VPWR
flabel metal1 2828 -2749 2862 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_34/VGND
flabel metal1 2828 -2205 2862 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_34/VPWR
flabel nwell 2828 -2205 2862 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_34/VPB
flabel pwell 2828 -2749 2862 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_34/VNB
rlabel comment 2891 -2732 2891 -2732 6 sky130_fd_sc_hd__decap_4_34/decap_4
rlabel metal1 2523 -2780 2891 -2684 1 sky130_fd_sc_hd__decap_4_34/VGND
rlabel metal1 2523 -2236 2891 -2140 1 sky130_fd_sc_hd__decap_4_34/VPWR
flabel metal1 1540 -2749 1574 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_56/VGND
flabel metal1 1540 -2205 1574 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_56/VPWR
flabel nwell 1540 -2205 1574 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_56/VPB
flabel pwell 1540 -2749 1574 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_56/VNB
rlabel comment 1603 -2732 1603 -2732 6 sky130_fd_sc_hd__decap_4_56/decap_4
rlabel metal1 1235 -2780 1603 -2684 1 sky130_fd_sc_hd__decap_4_56/VGND
rlabel metal1 1235 -2236 1603 -2140 1 sky130_fd_sc_hd__decap_4_56/VPWR
flabel metal1 1724 -2205 1758 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_94/VPWR
flabel metal1 1724 -2749 1758 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_94/VGND
flabel nwell 1724 -2205 1758 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_94/VPB
flabel pwell 1724 -2749 1758 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_94/VNB
rlabel comment 1695 -2732 1695 -2732 4 sky130_fd_sc_hd__decap_8_94/decap_8
rlabel metal1 1695 -2780 2431 -2684 1 sky130_fd_sc_hd__decap_8_94/VGND
rlabel metal1 1695 -2236 2431 -2140 1 sky130_fd_sc_hd__decap_8_94/VPWR
flabel metal1 2448 -2208 2501 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_60/VPWR
flabel metal1 2451 -2750 2502 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_60/VGND
rlabel comment 2523 -2732 2523 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_60/tapvpwrvgnd_1
rlabel metal1 2431 -2780 2523 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_60/VGND
rlabel metal1 2431 -2236 2523 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_60/VPWR
flabel metal1 1160 -2208 1213 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_100/VPWR
flabel metal1 1163 -2750 1214 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_100/VGND
rlabel comment 1235 -2732 1235 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_100/tapvpwrvgnd_1
rlabel metal1 1143 -2780 1235 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_100/VGND
rlabel metal1 1143 -2236 1235 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_100/VPWR
flabel metal1 1620 -2208 1673 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_101/VPWR
flabel metal1 1623 -2750 1674 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_101/VGND
rlabel comment 1695 -2732 1695 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_101/tapvpwrvgnd_1
rlabel metal1 1603 -2780 1695 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_101/VGND
rlabel metal1 1603 -2236 1695 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_101/VPWR
flabel locali 3013 -2511 3047 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A
flabel locali 3659 -2307 3693 -2273 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/X
flabel locali 3659 -2375 3693 -2341 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/X
flabel locali 3659 -2443 3693 -2409 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/X
flabel locali 3659 -2511 3693 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/X
flabel locali 3659 -2579 3693 -2545 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/X
flabel locali 3659 -2647 3693 -2613 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/X
flabel pwell 3013 -2749 3047 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/VNB
flabel nwell 3013 -2205 3047 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/VPB
flabel metal1 3013 -2749 3047 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/VGND
flabel metal1 3013 -2205 3047 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_25/VPWR
rlabel comment 2983 -2732 2983 -2732 4 sky130_fd_sc_hd__clkdlybuf4s50_1_25/clkdlybuf4s50_1
rlabel metal1 2983 -2780 3719 -2684 1 sky130_fd_sc_hd__clkdlybuf4s50_1_25/VGND
rlabel metal1 2983 -2236 3719 -2140 1 sky130_fd_sc_hd__clkdlybuf4s50_1_25/VPWR
flabel metal1 4116 -2749 4150 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_35/VGND
flabel metal1 4116 -2205 4150 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_35/VPWR
flabel nwell 4116 -2205 4150 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_35/VPB
flabel pwell 4116 -2749 4150 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_35/VNB
rlabel comment 4179 -2732 4179 -2732 6 sky130_fd_sc_hd__decap_4_35/decap_4
rlabel metal1 3811 -2780 4179 -2684 1 sky130_fd_sc_hd__decap_4_35/VGND
rlabel metal1 3811 -2236 4179 -2140 1 sky130_fd_sc_hd__decap_4_35/VPWR
flabel metal1 4300 -2205 4334 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_109/VPWR
flabel metal1 4300 -2749 4334 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_109/VGND
flabel nwell 4300 -2205 4334 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_109/VPB
flabel pwell 4300 -2749 4334 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_109/VNB
rlabel comment 4271 -2732 4271 -2732 4 sky130_fd_sc_hd__decap_8_109/decap_8
rlabel metal1 4271 -2780 5007 -2684 1 sky130_fd_sc_hd__decap_8_109/VGND
rlabel metal1 4271 -2236 5007 -2140 1 sky130_fd_sc_hd__decap_8_109/VPWR
flabel metal1 2908 -2208 2961 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_61/VPWR
flabel metal1 2911 -2750 2962 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_61/VGND
rlabel comment 2983 -2732 2983 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_61/tapvpwrvgnd_1
rlabel metal1 2891 -2780 2983 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_61/VGND
rlabel metal1 2891 -2236 2983 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_61/VPWR
flabel metal1 3736 -2208 3789 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_62/VPWR
flabel metal1 3739 -2750 3790 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_62/VGND
rlabel comment 3811 -2732 3811 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_62/tapvpwrvgnd_1
rlabel metal1 3719 -2780 3811 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_62/VGND
rlabel metal1 3719 -2236 3811 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_62/VPWR
flabel metal1 4196 -2208 4249 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_63/VPWR
flabel metal1 4199 -2750 4250 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_63/VGND
rlabel comment 4271 -2732 4271 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_63/tapvpwrvgnd_1
rlabel metal1 4179 -2780 4271 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_63/VGND
rlabel metal1 4179 -2236 4271 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_63/VPWR
flabel locali 5589 -2511 5623 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A
flabel locali 6235 -2307 6269 -2273 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/X
flabel locali 6235 -2375 6269 -2341 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/X
flabel locali 6235 -2443 6269 -2409 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/X
flabel locali 6235 -2511 6269 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/X
flabel locali 6235 -2579 6269 -2545 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/X
flabel locali 6235 -2647 6269 -2613 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/X
flabel pwell 5589 -2749 5623 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/VNB
flabel nwell 5589 -2205 5623 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/VPB
flabel metal1 5589 -2749 5623 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/VGND
flabel metal1 5589 -2205 5623 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_27/VPWR
rlabel comment 5559 -2732 5559 -2732 4 sky130_fd_sc_hd__clkdlybuf4s50_1_27/clkdlybuf4s50_1
rlabel metal1 5559 -2780 6295 -2684 1 sky130_fd_sc_hd__clkdlybuf4s50_1_27/VGND
rlabel metal1 5559 -2236 6295 -2140 1 sky130_fd_sc_hd__clkdlybuf4s50_1_27/VPWR
flabel metal1 5404 -2749 5438 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_36/VGND
flabel metal1 5404 -2205 5438 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_36/VPWR
flabel nwell 5404 -2205 5438 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_36/VPB
flabel pwell 5404 -2749 5438 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_36/VNB
rlabel comment 5467 -2732 5467 -2732 6 sky130_fd_sc_hd__decap_4_36/decap_4
rlabel metal1 5099 -2780 5467 -2684 1 sky130_fd_sc_hd__decap_4_36/VGND
rlabel metal1 5099 -2236 5467 -2140 1 sky130_fd_sc_hd__decap_4_36/VPWR
flabel metal1 6692 -2749 6726 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_37/VGND
flabel metal1 6692 -2205 6726 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_37/VPWR
flabel nwell 6692 -2205 6726 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_37/VPB
flabel pwell 6692 -2749 6726 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_37/VNB
rlabel comment 6755 -2732 6755 -2732 6 sky130_fd_sc_hd__decap_4_37/decap_4
rlabel metal1 6387 -2780 6755 -2684 1 sky130_fd_sc_hd__decap_4_37/VGND
rlabel metal1 6387 -2236 6755 -2140 1 sky130_fd_sc_hd__decap_4_37/VPWR
flabel metal1 5024 -2208 5077 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_64/VPWR
flabel metal1 5027 -2750 5078 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_64/VGND
rlabel comment 5099 -2732 5099 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_64/tapvpwrvgnd_1
rlabel metal1 5007 -2780 5099 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_64/VGND
rlabel metal1 5007 -2236 5099 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_64/VPWR
flabel metal1 5484 -2208 5537 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_65/VPWR
flabel metal1 5487 -2750 5538 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_65/VGND
rlabel comment 5559 -2732 5559 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_65/tapvpwrvgnd_1
rlabel metal1 5467 -2780 5559 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_65/VGND
rlabel metal1 5467 -2236 5559 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_65/VPWR
flabel metal1 6312 -2208 6365 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_66/VPWR
flabel metal1 6315 -2750 6366 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_66/VGND
rlabel comment 6387 -2732 6387 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_66/tapvpwrvgnd_1
rlabel metal1 6295 -2780 6387 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_66/VGND
rlabel metal1 6295 -2236 6387 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_66/VPWR
flabel locali 8165 -2511 8199 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A
flabel locali 8811 -2307 8845 -2273 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/X
flabel locali 8811 -2375 8845 -2341 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/X
flabel locali 8811 -2443 8845 -2409 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/X
flabel locali 8811 -2511 8845 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/X
flabel locali 8811 -2579 8845 -2545 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/X
flabel locali 8811 -2647 8845 -2613 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/X
flabel pwell 8165 -2749 8199 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/VNB
flabel nwell 8165 -2205 8199 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/VPB
flabel metal1 8165 -2749 8199 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/VGND
flabel metal1 8165 -2205 8199 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_29/VPWR
rlabel comment 8135 -2732 8135 -2732 4 sky130_fd_sc_hd__clkdlybuf4s50_1_29/clkdlybuf4s50_1
rlabel metal1 8135 -2780 8871 -2684 1 sky130_fd_sc_hd__clkdlybuf4s50_1_29/VGND
rlabel metal1 8135 -2236 8871 -2140 1 sky130_fd_sc_hd__clkdlybuf4s50_1_29/VPWR
flabel metal1 7980 -2749 8014 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_38/VGND
flabel metal1 7980 -2205 8014 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_38/VPWR
flabel nwell 7980 -2205 8014 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_38/VPB
flabel pwell 7980 -2749 8014 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_38/VNB
rlabel comment 8043 -2732 8043 -2732 6 sky130_fd_sc_hd__decap_4_38/decap_4
rlabel metal1 7675 -2780 8043 -2684 1 sky130_fd_sc_hd__decap_4_38/VGND
rlabel metal1 7675 -2236 8043 -2140 1 sky130_fd_sc_hd__decap_4_38/VPWR
flabel metal1 6876 -2205 6910 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_118/VPWR
flabel metal1 6876 -2749 6910 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_118/VGND
flabel nwell 6876 -2205 6910 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_118/VPB
flabel pwell 6876 -2749 6910 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_118/VNB
rlabel comment 6847 -2732 6847 -2732 4 sky130_fd_sc_hd__decap_8_118/decap_8
rlabel metal1 6847 -2780 7583 -2684 1 sky130_fd_sc_hd__decap_8_118/VGND
rlabel metal1 6847 -2236 7583 -2140 1 sky130_fd_sc_hd__decap_8_118/VPWR
flabel metal1 6772 -2208 6825 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_67/VPWR
flabel metal1 6775 -2750 6826 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_67/VGND
rlabel comment 6847 -2732 6847 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_67/tapvpwrvgnd_1
rlabel metal1 6755 -2780 6847 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_67/VGND
rlabel metal1 6755 -2236 6847 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_67/VPWR
flabel metal1 7600 -2208 7653 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_68/VPWR
flabel metal1 7603 -2750 7654 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_68/VGND
rlabel comment 7675 -2732 7675 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_68/tapvpwrvgnd_1
rlabel metal1 7583 -2780 7675 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_68/VGND
rlabel metal1 7583 -2236 7675 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_68/VPWR
flabel metal1 8060 -2208 8113 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_69/VPWR
flabel metal1 8063 -2750 8114 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_69/VGND
rlabel comment 8135 -2732 8135 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_69/tapvpwrvgnd_1
rlabel metal1 8043 -2780 8135 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_69/VGND
rlabel metal1 8043 -2236 8135 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_69/VPWR
flabel metal1 9268 -2749 9302 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_39/VGND
flabel metal1 9268 -2205 9302 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_39/VPWR
flabel nwell 9268 -2205 9302 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_39/VPB
flabel pwell 9268 -2749 9302 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_39/VNB
rlabel comment 9331 -2732 9331 -2732 6 sky130_fd_sc_hd__decap_4_39/decap_4
rlabel metal1 8963 -2780 9331 -2684 1 sky130_fd_sc_hd__decap_4_39/VGND
rlabel metal1 8963 -2236 9331 -2140 1 sky130_fd_sc_hd__decap_4_39/VPWR
flabel metal1 10648 -2749 10682 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_40/VGND
flabel metal1 10648 -2205 10682 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_40/VPWR
flabel nwell 10648 -2205 10682 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_40/VPB
flabel pwell 10648 -2749 10682 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_40/VNB
rlabel comment 10711 -2732 10711 -2732 6 sky130_fd_sc_hd__decap_4_40/decap_4
rlabel metal1 10343 -2780 10711 -2684 1 sky130_fd_sc_hd__decap_4_40/VGND
rlabel metal1 10343 -2236 10711 -2140 1 sky130_fd_sc_hd__decap_4_40/VPWR
flabel metal1 9452 -2205 9486 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_128/VPWR
flabel metal1 9452 -2749 9486 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_128/VGND
flabel nwell 9452 -2205 9486 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_128/VPB
flabel pwell 9452 -2749 9486 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_128/VNB
rlabel comment 9423 -2732 9423 -2732 4 sky130_fd_sc_hd__decap_8_128/decap_8
rlabel metal1 9423 -2780 10159 -2684 1 sky130_fd_sc_hd__decap_8_128/VGND
rlabel metal1 9423 -2236 10159 -2140 1 sky130_fd_sc_hd__decap_8_128/VPWR
flabel metal1 10285 -2205 10321 -2175 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_9/VPWR
flabel metal1 10285 -2745 10321 -2716 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_9/VGND
flabel nwell 10292 -2198 10312 -2181 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_9/VPB
flabel pwell 10291 -2743 10315 -2721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_9/VNB
rlabel comment 10343 -2732 10343 -2732 6 sky130_fd_sc_hd__fill_1_9/fill_1
rlabel metal1 10251 -2780 10343 -2684 1 sky130_fd_sc_hd__fill_1_9/VGND
rlabel metal1 10251 -2236 10343 -2140 1 sky130_fd_sc_hd__fill_1_9/VPWR
flabel metal1 8888 -2208 8941 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_70/VPWR
flabel metal1 8891 -2750 8942 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_70/VGND
rlabel comment 8963 -2732 8963 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_70/tapvpwrvgnd_1
rlabel metal1 8871 -2780 8963 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_70/VGND
rlabel metal1 8871 -2236 8963 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_70/VPWR
flabel metal1 9348 -2208 9401 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_71/VPWR
flabel metal1 9351 -2750 9402 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_71/VGND
rlabel comment 9423 -2732 9423 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_71/tapvpwrvgnd_1
rlabel metal1 9331 -2780 9423 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_71/VGND
rlabel metal1 9331 -2236 9423 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_71/VPWR
flabel metal1 10176 -2208 10229 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_72/VPWR
flabel metal1 10179 -2750 10230 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_72/VGND
rlabel comment 10251 -2732 10251 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_72/tapvpwrvgnd_1
rlabel metal1 10159 -2780 10251 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_72/VGND
rlabel metal1 10159 -2236 10251 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_72/VPWR
flabel locali 10741 -2511 10775 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A
flabel locali 11387 -2307 11421 -2273 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X
flabel locali 11387 -2375 11421 -2341 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X
flabel locali 11387 -2443 11421 -2409 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X
flabel locali 11387 -2511 11421 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X
flabel locali 11387 -2579 11421 -2545 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X
flabel locali 11387 -2647 11421 -2613 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X
flabel pwell 10741 -2749 10775 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/VNB
flabel nwell 10741 -2205 10775 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/VPB
flabel metal1 10741 -2749 10775 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/VGND
flabel metal1 10741 -2205 10775 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_31/VPWR
rlabel comment 10711 -2732 10711 -2732 4 sky130_fd_sc_hd__clkdlybuf4s50_1_31/clkdlybuf4s50_1
rlabel metal1 10711 -2780 11447 -2684 1 sky130_fd_sc_hd__clkdlybuf4s50_1_31/VGND
rlabel metal1 10711 -2236 11447 -2140 1 sky130_fd_sc_hd__clkdlybuf4s50_1_31/VPWR
flabel metal1 11936 -2749 11970 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_41/VGND
flabel metal1 11936 -2205 11970 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_41/VPWR
flabel nwell 11936 -2205 11970 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_41/VPB
flabel pwell 11936 -2749 11970 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_41/VNB
rlabel comment 11999 -2732 11999 -2732 6 sky130_fd_sc_hd__decap_4_41/decap_4
rlabel metal1 11631 -2780 11999 -2684 1 sky130_fd_sc_hd__decap_4_41/VGND
rlabel metal1 11631 -2236 11999 -2140 1 sky130_fd_sc_hd__decap_4_41/VPWR
flabel metal1 10653 -2205 10689 -2175 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_10/VPWR
flabel metal1 10653 -2745 10689 -2716 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_10/VGND
flabel nwell 10660 -2198 10680 -2181 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_10/VPB
flabel pwell 10659 -2743 10683 -2721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_10/VNB
rlabel comment 10711 -2732 10711 -2732 6 sky130_fd_sc_hd__fill_1_10/fill_1
rlabel metal1 10619 -2780 10711 -2684 1 sky130_fd_sc_hd__fill_1_10/VGND
rlabel metal1 10619 -2236 10711 -2140 1 sky130_fd_sc_hd__fill_1_10/VPWR
flabel metal1 11573 -2205 11609 -2175 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_11/VPWR
flabel metal1 11573 -2745 11609 -2716 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_11/VGND
flabel nwell 11580 -2198 11600 -2181 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_11/VPB
flabel pwell 11579 -2743 11603 -2721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_11/VNB
rlabel comment 11631 -2732 11631 -2732 6 sky130_fd_sc_hd__fill_1_11/fill_1
rlabel metal1 11539 -2780 11631 -2684 1 sky130_fd_sc_hd__fill_1_11/VGND
rlabel metal1 11539 -2236 11631 -2140 1 sky130_fd_sc_hd__fill_1_11/VPWR
flabel metal1 12033 -2742 12056 -2723 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_3/VGND
flabel metal1 12033 -2197 12053 -2180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_3/VPWR
flabel nwell 12034 -2202 12059 -2176 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_3/VPB
flabel pwell 12034 -2744 12056 -2720 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_3/VNB
rlabel comment 11999 -2732 11999 -2732 4 sky130_fd_sc_hd__fill_4_3/fill_4
rlabel metal1 11999 -2780 12367 -2684 1 sky130_fd_sc_hd__fill_4_3/VGND
rlabel metal1 11999 -2236 12367 -2140 1 sky130_fd_sc_hd__fill_4_3/VPWR
flabel metal1 11464 -2208 11517 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_73/VPWR
flabel metal1 11467 -2750 11518 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_73/VGND
rlabel comment 11539 -2732 11539 -2732 6 sky130_fd_sc_hd__tapvpwrvgnd_1_73/tapvpwrvgnd_1
rlabel metal1 11447 -2780 11539 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_73/VGND
rlabel metal1 11447 -2236 11539 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_73/VPWR
flabel locali 15248 -2443 15282 -2409 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/X
flabel locali 15340 -2443 15374 -2409 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/X
flabel locali 15340 -2511 15374 -2477 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/X
flabel locali 15248 -2511 15282 -2477 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/X
flabel locali 15248 -2579 15282 -2545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/X
flabel locali 15340 -2579 15374 -2545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/X
flabel locali 13684 -2579 13718 -2545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/A
flabel locali 13684 -2511 13718 -2477 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/A
flabel pwell 13684 -2749 13718 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/VNB
flabel pwell 13701 -2732 13701 -2732 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/VNB
flabel nwell 13684 -2205 13718 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/VPB
flabel nwell 13701 -2188 13701 -2188 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/VPB
flabel metal1 13684 -2749 13718 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/VGND
flabel metal1 13684 -2205 13718 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_3/VPWR
rlabel comment 13655 -2732 13655 -2732 4 sky130_fd_sc_hd__clkbuf_16_3/clkbuf_16
rlabel metal1 13655 -2780 15495 -2684 1 sky130_fd_sc_hd__clkbuf_16_3/VGND
rlabel metal1 13655 -2236 15495 -2140 1 sky130_fd_sc_hd__clkbuf_16_3/VPWR
flabel locali 12672 -2511 12706 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/A
flabel locali 12764 -2511 12798 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/A
flabel locali 13040 -2579 13074 -2545 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/Y
flabel locali 12580 -2511 12614 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/A
flabel locali 13040 -2443 13074 -2409 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/Y
flabel locali 12948 -2511 12982 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/A
flabel locali 12856 -2511 12890 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/A
flabel locali 13040 -2511 13074 -2477 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_2/Y
flabel pwell 12488 -2749 12522 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_2/VNB
flabel nwell 12488 -2205 12522 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_2/VPB
flabel metal1 12488 -2205 12522 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_2/VPWR
flabel metal1 12488 -2749 12522 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_2/VGND
rlabel comment 12459 -2732 12459 -2732 4 sky130_fd_sc_hd__clkinv_4_2/clkinv_4
rlabel metal1 12459 -2780 13103 -2684 1 sky130_fd_sc_hd__clkinv_4_2/VGND
rlabel metal1 12459 -2236 13103 -2140 1 sky130_fd_sc_hd__clkinv_4_2/VPWR
flabel metal1 13224 -2749 13258 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_63/VGND
flabel metal1 13224 -2205 13258 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_63/VPWR
flabel nwell 13224 -2205 13258 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_63/VPB
flabel pwell 13224 -2749 13258 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_63/VNB
rlabel comment 13195 -2732 13195 -2732 4 sky130_fd_sc_hd__decap_4_63/decap_4
rlabel metal1 13195 -2780 13563 -2684 1 sky130_fd_sc_hd__decap_4_63/VGND
rlabel metal1 13195 -2236 13563 -2140 1 sky130_fd_sc_hd__decap_4_63/VPWR
flabel metal1 12389 -2208 12442 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_114/VPWR
flabel metal1 12388 -2750 12439 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_114/VGND
rlabel comment 12367 -2732 12367 -2732 4 sky130_fd_sc_hd__tapvpwrvgnd_1_114/tapvpwrvgnd_1
rlabel metal1 12367 -2780 12459 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_114/VGND
rlabel metal1 12367 -2236 12459 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_114/VPWR
flabel metal1 13125 -2208 13178 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_115/VPWR
flabel metal1 13124 -2750 13175 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_115/VGND
rlabel comment 13103 -2732 13103 -2732 4 sky130_fd_sc_hd__tapvpwrvgnd_1_115/tapvpwrvgnd_1
rlabel metal1 13103 -2780 13195 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_115/VGND
rlabel metal1 13103 -2236 13195 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_115/VPWR
flabel metal1 13585 -2208 13638 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_116/VPWR
flabel metal1 13584 -2750 13635 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_116/VGND
rlabel comment 13563 -2732 13563 -2732 4 sky130_fd_sc_hd__tapvpwrvgnd_1_116/tapvpwrvgnd_1
rlabel metal1 13563 -2780 13655 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_116/VGND
rlabel metal1 13563 -2236 13655 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_116/VPWR
flabel metal1 15616 -2749 15650 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_6/VGND
flabel metal1 15616 -2205 15650 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_6/VPWR
flabel nwell 15616 -2205 15650 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_6/VPB
flabel pwell 15616 -2749 15650 -2715 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_6/VNB
rlabel comment 15587 -2732 15587 -2732 4 sky130_fd_sc_hd__decap_12_6/decap_12
rlabel metal1 15587 -2780 16691 -2684 1 sky130_fd_sc_hd__decap_12_6/VGND
rlabel metal1 15587 -2236 16691 -2140 1 sky130_fd_sc_hd__decap_12_6/VPWR
flabel metal1 15517 -2208 15570 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_130/VPWR
flabel metal1 15516 -2750 15567 -2712 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_130/VGND
rlabel comment 15495 -2732 15495 -2732 4 sky130_fd_sc_hd__tapvpwrvgnd_1_130/tapvpwrvgnd_1
rlabel metal1 15495 -2780 15587 -2684 1 sky130_fd_sc_hd__tapvpwrvgnd_1_130/VGND
rlabel metal1 15495 -2236 15587 -2140 1 sky130_fd_sc_hd__tapvpwrvgnd_1_130/VPWR
flabel metal1 -944 -2205 -910 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_4/VPWR
flabel metal1 -944 -1661 -910 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_4/VGND
flabel nwell -944 -2205 -910 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_4/VPB
flabel pwell -944 -1661 -910 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_4/VNB
rlabel comment -881 -1644 -881 -1644 8 sky130_fd_sc_hd__decap_8_4/decap_8
rlabel metal1 -1617 -1692 -881 -1596 5 sky130_fd_sc_hd__decap_8_4/VGND
rlabel metal1 -1617 -2236 -881 -2140 5 sky130_fd_sc_hd__decap_8_4/VPWR
flabel metal1 -2324 -2205 -2290 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_69/VPWR
flabel metal1 -2324 -1661 -2290 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_69/VGND
flabel nwell -2324 -2205 -2290 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_69/VPB
flabel pwell -2324 -1661 -2290 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_69/VNB
rlabel comment -2261 -1644 -2261 -1644 8 sky130_fd_sc_hd__decap_8_69/decap_8
rlabel metal1 -2997 -1692 -2261 -1596 5 sky130_fd_sc_hd__decap_8_69/VGND
rlabel metal1 -2997 -2236 -2261 -2140 5 sky130_fd_sc_hd__decap_8_69/VPWR
flabel metal1 -1690 -1662 -1637 -1630 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_7/VGND
flabel metal1 -1690 -2205 -1638 -2174 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_7/VPWR
flabel nwell -1679 -2197 -1645 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_7/VPB
flabel pwell -1680 -1656 -1648 -1634 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_7/VNB
rlabel comment -1617 -1644 -1617 -1644 8 sky130_fd_sc_hd__fill_2_7/fill_2
rlabel metal1 -1801 -1692 -1617 -1596 5 sky130_fd_sc_hd__fill_2_7/VGND
rlabel metal1 -1801 -2236 -1617 -2140 5 sky130_fd_sc_hd__fill_2_7/VPWR
flabel metal1 -1858 -1653 -1835 -1634 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_20/VGND
flabel metal1 -1855 -2196 -1835 -2179 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_20/VPWR
flabel nwell -1861 -2200 -1836 -2174 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_20/VPB
flabel pwell -1858 -1656 -1836 -1632 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_20/VNB
rlabel comment -1801 -1644 -1801 -1644 8 sky130_fd_sc_hd__fill_4_20/fill_4
rlabel metal1 -2169 -1692 -1801 -1596 5 sky130_fd_sc_hd__fill_4_20/VGND
rlabel metal1 -2169 -2236 -1801 -2140 5 sky130_fd_sc_hd__fill_4_20/VPWR
flabel metal1 -2244 -2197 -2191 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_534/VPWR
flabel metal1 -2241 -1664 -2190 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_534/VGND
rlabel comment -2169 -1644 -2169 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_534/tapvpwrvgnd_1
rlabel metal1 -2261 -1692 -2169 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_534/VGND
rlabel metal1 -2261 -2236 -2169 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_534/VPWR
flabel locali 1079 -1899 1113 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A
flabel locali 433 -2103 467 -2069 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X
flabel locali 433 -2035 467 -2001 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X
flabel locali 433 -1967 467 -1933 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X
flabel locali 433 -1899 467 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X
flabel locali 433 -1831 467 -1797 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X
flabel locali 433 -1763 467 -1729 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X
flabel pwell 1079 -1661 1113 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/VNB
flabel nwell 1079 -2205 1113 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/VPB
flabel metal1 1079 -1661 1113 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/VGND
flabel metal1 1079 -2205 1113 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_48/VPWR
rlabel comment 1143 -1644 1143 -1644 8 sky130_fd_sc_hd__clkdlybuf4s50_1_48/clkdlybuf4s50_1
rlabel metal1 407 -1692 1143 -1596 5 sky130_fd_sc_hd__clkdlybuf4s50_1_48/VGND
rlabel metal1 407 -2236 1143 -2140 5 sky130_fd_sc_hd__clkdlybuf4s50_1_48/VPWR
flabel locali -209 -1899 -175 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A
flabel locali -855 -2103 -821 -2069 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X
flabel locali -855 -2035 -821 -2001 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X
flabel locali -855 -1967 -821 -1933 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X
flabel locali -855 -1899 -821 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X
flabel locali -855 -1831 -821 -1797 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X
flabel locali -855 -1763 -821 -1729 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/X
flabel pwell -209 -1661 -175 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/VNB
flabel nwell -209 -2205 -175 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/VPB
flabel metal1 -209 -1661 -175 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/VGND
flabel metal1 -209 -2205 -175 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_49/VPWR
rlabel comment -145 -1644 -145 -1644 8 sky130_fd_sc_hd__clkdlybuf4s50_1_49/clkdlybuf4s50_1
rlabel metal1 -881 -1692 -145 -1596 5 sky130_fd_sc_hd__clkdlybuf4s50_1_49/VGND
rlabel metal1 -881 -2236 -145 -2140 5 sky130_fd_sc_hd__clkdlybuf4s50_1_49/VPWR
flabel metal1 252 -1661 286 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_59/VGND
flabel metal1 252 -2205 286 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_59/VPWR
flabel nwell 252 -2205 286 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_59/VPB
flabel pwell 252 -1661 286 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_59/VNB
rlabel comment 315 -1644 315 -1644 8 sky130_fd_sc_hd__decap_4_59/decap_4
rlabel metal1 -53 -1692 315 -1596 5 sky130_fd_sc_hd__decap_4_59/VGND
rlabel metal1 -53 -2236 315 -2140 5 sky130_fd_sc_hd__decap_4_59/VPWR
flabel metal1 332 -2197 385 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_105/VPWR
flabel metal1 335 -1664 386 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_105/VGND
rlabel comment 407 -1644 407 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_105/tapvpwrvgnd_1
rlabel metal1 315 -1692 407 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_105/VGND
rlabel metal1 315 -2236 407 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_105/VPWR
flabel metal1 -128 -2197 -75 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_107/VPWR
flabel metal1 -125 -1664 -74 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_107/VGND
rlabel comment -53 -1644 -53 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_107/tapvpwrvgnd_1
rlabel metal1 -145 -1692 -53 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_107/VGND
rlabel metal1 -145 -2236 -53 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_107/VPWR
flabel metal1 2828 -1661 2862 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_18/VGND
flabel metal1 2828 -2205 2862 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_18/VPWR
flabel nwell 2828 -2205 2862 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_18/VPB
flabel pwell 2828 -1661 2862 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_18/VNB
rlabel comment 2891 -1644 2891 -1644 8 sky130_fd_sc_hd__decap_4_18/decap_4
rlabel metal1 2523 -1692 2891 -1596 5 sky130_fd_sc_hd__decap_4_18/VGND
rlabel metal1 2523 -2236 2891 -2140 5 sky130_fd_sc_hd__decap_4_18/VPWR
flabel metal1 1540 -1661 1574 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_57/VGND
flabel metal1 1540 -2205 1574 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_57/VPWR
flabel nwell 1540 -2205 1574 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_57/VPB
flabel pwell 1540 -1661 1574 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_57/VNB
rlabel comment 1603 -1644 1603 -1644 8 sky130_fd_sc_hd__decap_4_57/decap_4
rlabel metal1 1235 -1692 1603 -1596 5 sky130_fd_sc_hd__decap_4_57/VGND
rlabel metal1 1235 -2236 1603 -2140 5 sky130_fd_sc_hd__decap_4_57/VPWR
flabel metal1 2368 -2205 2402 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_93/VPWR
flabel metal1 2368 -1661 2402 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_93/VGND
flabel nwell 2368 -2205 2402 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_93/VPB
flabel pwell 2368 -1661 2402 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_93/VNB
rlabel comment 2431 -1644 2431 -1644 8 sky130_fd_sc_hd__decap_8_93/decap_8
rlabel metal1 1695 -1692 2431 -1596 5 sky130_fd_sc_hd__decap_8_93/VGND
rlabel metal1 1695 -2236 2431 -2140 5 sky130_fd_sc_hd__decap_8_93/VPWR
flabel metal1 2448 -2197 2501 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_32/VPWR
flabel metal1 2451 -1664 2502 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_32/VGND
rlabel comment 2523 -1644 2523 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_32/tapvpwrvgnd_1
rlabel metal1 2431 -1692 2523 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_32/VGND
rlabel metal1 2431 -2236 2523 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_32/VPWR
flabel metal1 1160 -2197 1213 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_102/VPWR
flabel metal1 1163 -1664 1214 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_102/VGND
rlabel comment 1235 -1644 1235 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_102/tapvpwrvgnd_1
rlabel metal1 1143 -1692 1235 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_102/VGND
rlabel metal1 1143 -2236 1235 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_102/VPWR
flabel metal1 1620 -2197 1673 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_103/VPWR
flabel metal1 1623 -1664 1674 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_103/VGND
rlabel comment 1695 -1644 1695 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_103/tapvpwrvgnd_1
rlabel metal1 1603 -1692 1695 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_103/VGND
rlabel metal1 1603 -2236 1695 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_103/VPWR
flabel locali 3655 -1899 3689 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/A
flabel locali 3009 -2103 3043 -2069 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X
flabel locali 3009 -2035 3043 -2001 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X
flabel locali 3009 -1967 3043 -1933 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X
flabel locali 3009 -1899 3043 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X
flabel locali 3009 -1831 3043 -1797 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X
flabel locali 3009 -1763 3043 -1729 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/X
flabel pwell 3655 -1661 3689 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/VNB
flabel nwell 3655 -2205 3689 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/VPB
flabel metal1 3655 -1661 3689 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/VGND
flabel metal1 3655 -2205 3689 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_11/VPWR
rlabel comment 3719 -1644 3719 -1644 8 sky130_fd_sc_hd__clkdlybuf4s50_1_11/clkdlybuf4s50_1
rlabel metal1 2983 -1692 3719 -1596 5 sky130_fd_sc_hd__clkdlybuf4s50_1_11/VGND
rlabel metal1 2983 -2236 3719 -2140 5 sky130_fd_sc_hd__clkdlybuf4s50_1_11/VPWR
flabel metal1 4116 -1661 4150 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_19/VGND
flabel metal1 4116 -2205 4150 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_19/VPWR
flabel nwell 4116 -2205 4150 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_19/VPB
flabel pwell 4116 -1661 4150 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_19/VNB
rlabel comment 4179 -1644 4179 -1644 8 sky130_fd_sc_hd__decap_4_19/decap_4
rlabel metal1 3811 -1692 4179 -1596 5 sky130_fd_sc_hd__decap_4_19/VGND
rlabel metal1 3811 -2236 4179 -2140 5 sky130_fd_sc_hd__decap_4_19/VPWR
flabel metal1 4944 -2205 4978 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_110/VPWR
flabel metal1 4944 -1661 4978 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_110/VGND
flabel nwell 4944 -2205 4978 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_110/VPB
flabel pwell 4944 -1661 4978 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_110/VNB
rlabel comment 5007 -1644 5007 -1644 8 sky130_fd_sc_hd__decap_8_110/decap_8
rlabel metal1 4271 -1692 5007 -1596 5 sky130_fd_sc_hd__decap_8_110/VGND
rlabel metal1 4271 -2236 5007 -2140 5 sky130_fd_sc_hd__decap_8_110/VPWR
flabel metal1 2908 -2197 2961 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_33/VPWR
flabel metal1 2911 -1664 2962 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_33/VGND
rlabel comment 2983 -1644 2983 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_33/tapvpwrvgnd_1
rlabel metal1 2891 -1692 2983 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_33/VGND
rlabel metal1 2891 -2236 2983 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_33/VPWR
flabel metal1 3736 -2197 3789 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_34/VPWR
flabel metal1 3739 -1664 3790 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_34/VGND
rlabel comment 3811 -1644 3811 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_34/tapvpwrvgnd_1
rlabel metal1 3719 -1692 3811 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_34/VGND
rlabel metal1 3719 -2236 3811 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_34/VPWR
flabel metal1 4196 -2197 4249 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_35/VPWR
flabel metal1 4199 -1664 4250 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_35/VGND
rlabel comment 4271 -1644 4271 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_35/tapvpwrvgnd_1
rlabel metal1 4179 -1692 4271 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_35/VGND
rlabel metal1 4179 -2236 4271 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_35/VPWR
flabel locali 6231 -1899 6265 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/A
flabel locali 5585 -2103 5619 -2069 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
flabel locali 5585 -2035 5619 -2001 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
flabel locali 5585 -1967 5619 -1933 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
flabel locali 5585 -1899 5619 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
flabel locali 5585 -1831 5619 -1797 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
flabel locali 5585 -1763 5619 -1729 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
flabel pwell 6231 -1661 6265 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/VNB
flabel nwell 6231 -2205 6265 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/VPB
flabel metal1 6231 -1661 6265 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/VGND
flabel metal1 6231 -2205 6265 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_13/VPWR
rlabel comment 6295 -1644 6295 -1644 8 sky130_fd_sc_hd__clkdlybuf4s50_1_13/clkdlybuf4s50_1
rlabel metal1 5559 -1692 6295 -1596 5 sky130_fd_sc_hd__clkdlybuf4s50_1_13/VGND
rlabel metal1 5559 -2236 6295 -2140 5 sky130_fd_sc_hd__clkdlybuf4s50_1_13/VPWR
flabel metal1 5404 -1661 5438 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_20/VGND
flabel metal1 5404 -2205 5438 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_20/VPWR
flabel nwell 5404 -2205 5438 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_20/VPB
flabel pwell 5404 -1661 5438 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_20/VNB
rlabel comment 5467 -1644 5467 -1644 8 sky130_fd_sc_hd__decap_4_20/decap_4
rlabel metal1 5099 -1692 5467 -1596 5 sky130_fd_sc_hd__decap_4_20/VGND
rlabel metal1 5099 -2236 5467 -2140 5 sky130_fd_sc_hd__decap_4_20/VPWR
flabel metal1 6692 -1661 6726 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_21/VGND
flabel metal1 6692 -2205 6726 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_21/VPWR
flabel nwell 6692 -2205 6726 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_21/VPB
flabel pwell 6692 -1661 6726 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_21/VNB
rlabel comment 6755 -1644 6755 -1644 8 sky130_fd_sc_hd__decap_4_21/decap_4
rlabel metal1 6387 -1692 6755 -1596 5 sky130_fd_sc_hd__decap_4_21/VGND
rlabel metal1 6387 -2236 6755 -2140 5 sky130_fd_sc_hd__decap_4_21/VPWR
flabel metal1 5024 -2197 5077 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_36/VPWR
flabel metal1 5027 -1664 5078 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_36/VGND
rlabel comment 5099 -1644 5099 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_36/tapvpwrvgnd_1
rlabel metal1 5007 -1692 5099 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_36/VGND
rlabel metal1 5007 -2236 5099 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_36/VPWR
flabel metal1 5484 -2197 5537 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_37/VPWR
flabel metal1 5487 -1664 5538 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_37/VGND
rlabel comment 5559 -1644 5559 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_37/tapvpwrvgnd_1
rlabel metal1 5467 -1692 5559 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_37/VGND
rlabel metal1 5467 -2236 5559 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_37/VPWR
flabel metal1 6312 -2197 6365 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_38/VPWR
flabel metal1 6315 -1664 6366 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_38/VGND
rlabel comment 6387 -1644 6387 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_38/tapvpwrvgnd_1
rlabel metal1 6295 -1692 6387 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_38/VGND
rlabel metal1 6295 -2236 6387 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_38/VPWR
flabel locali 8807 -1899 8841 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/A
flabel locali 8161 -2103 8195 -2069 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X
flabel locali 8161 -2035 8195 -2001 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X
flabel locali 8161 -1967 8195 -1933 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X
flabel locali 8161 -1899 8195 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X
flabel locali 8161 -1831 8195 -1797 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X
flabel locali 8161 -1763 8195 -1729 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X
flabel pwell 8807 -1661 8841 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/VNB
flabel nwell 8807 -2205 8841 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/VPB
flabel metal1 8807 -1661 8841 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/VGND
flabel metal1 8807 -2205 8841 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_15/VPWR
rlabel comment 8871 -1644 8871 -1644 8 sky130_fd_sc_hd__clkdlybuf4s50_1_15/clkdlybuf4s50_1
rlabel metal1 8135 -1692 8871 -1596 5 sky130_fd_sc_hd__clkdlybuf4s50_1_15/VGND
rlabel metal1 8135 -2236 8871 -2140 5 sky130_fd_sc_hd__clkdlybuf4s50_1_15/VPWR
flabel metal1 7980 -1661 8014 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_22/VGND
flabel metal1 7980 -2205 8014 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_22/VPWR
flabel nwell 7980 -2205 8014 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_22/VPB
flabel pwell 7980 -1661 8014 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_22/VNB
rlabel comment 8043 -1644 8043 -1644 8 sky130_fd_sc_hd__decap_4_22/decap_4
rlabel metal1 7675 -1692 8043 -1596 5 sky130_fd_sc_hd__decap_4_22/VGND
rlabel metal1 7675 -2236 8043 -2140 5 sky130_fd_sc_hd__decap_4_22/VPWR
flabel metal1 7520 -2205 7554 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_117/VPWR
flabel metal1 7520 -1661 7554 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_117/VGND
flabel nwell 7520 -2205 7554 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_117/VPB
flabel pwell 7520 -1661 7554 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_117/VNB
rlabel comment 7583 -1644 7583 -1644 8 sky130_fd_sc_hd__decap_8_117/decap_8
rlabel metal1 6847 -1692 7583 -1596 5 sky130_fd_sc_hd__decap_8_117/VGND
rlabel metal1 6847 -2236 7583 -2140 5 sky130_fd_sc_hd__decap_8_117/VPWR
flabel metal1 6772 -2197 6825 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_39/VPWR
flabel metal1 6775 -1664 6826 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_39/VGND
rlabel comment 6847 -1644 6847 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_39/tapvpwrvgnd_1
rlabel metal1 6755 -1692 6847 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_39/VGND
rlabel metal1 6755 -2236 6847 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_39/VPWR
flabel metal1 7600 -2197 7653 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_40/VPWR
flabel metal1 7603 -1664 7654 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_40/VGND
rlabel comment 7675 -1644 7675 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_40/tapvpwrvgnd_1
rlabel metal1 7583 -1692 7675 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_40/VGND
rlabel metal1 7583 -2236 7675 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_40/VPWR
flabel metal1 8060 -2197 8113 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_41/VPWR
flabel metal1 8063 -1664 8114 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_41/VGND
rlabel comment 8135 -1644 8135 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_41/tapvpwrvgnd_1
rlabel metal1 8043 -1692 8135 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_41/VGND
rlabel metal1 8043 -2236 8135 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_41/VPWR
flabel metal1 9268 -1661 9302 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_23/VGND
flabel metal1 9268 -2205 9302 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_23/VPWR
flabel nwell 9268 -2205 9302 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_23/VPB
flabel pwell 9268 -1661 9302 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_23/VNB
rlabel comment 9331 -1644 9331 -1644 8 sky130_fd_sc_hd__decap_4_23/decap_4
rlabel metal1 8963 -1692 9331 -1596 5 sky130_fd_sc_hd__decap_4_23/VGND
rlabel metal1 8963 -2236 9331 -2140 5 sky130_fd_sc_hd__decap_4_23/VPWR
flabel metal1 10648 -1661 10682 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_24/VGND
flabel metal1 10648 -2205 10682 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_24/VPWR
flabel nwell 10648 -2205 10682 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_24/VPB
flabel pwell 10648 -1661 10682 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_24/VNB
rlabel comment 10711 -1644 10711 -1644 8 sky130_fd_sc_hd__decap_4_24/decap_4
rlabel metal1 10343 -1692 10711 -1596 5 sky130_fd_sc_hd__decap_4_24/VGND
rlabel metal1 10343 -2236 10711 -2140 5 sky130_fd_sc_hd__decap_4_24/VPWR
flabel metal1 10096 -2205 10130 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_127/VPWR
flabel metal1 10096 -1661 10130 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_127/VGND
flabel nwell 10096 -2205 10130 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_127/VPB
flabel pwell 10096 -1661 10130 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_127/VNB
rlabel comment 10159 -1644 10159 -1644 8 sky130_fd_sc_hd__decap_8_127/decap_8
rlabel metal1 9423 -1692 10159 -1596 5 sky130_fd_sc_hd__decap_8_127/VGND
rlabel metal1 9423 -2236 10159 -2140 5 sky130_fd_sc_hd__decap_8_127/VPWR
flabel metal1 10285 -2201 10321 -2171 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_2/VPWR
flabel metal1 10285 -1660 10321 -1631 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_2/VGND
flabel nwell 10292 -2195 10312 -2178 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_2/VPB
flabel pwell 10291 -1655 10315 -1633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_2/VNB
rlabel comment 10343 -1644 10343 -1644 8 sky130_fd_sc_hd__fill_1_2/fill_1
rlabel metal1 10251 -1692 10343 -1596 5 sky130_fd_sc_hd__fill_1_2/VGND
rlabel metal1 10251 -2236 10343 -2140 5 sky130_fd_sc_hd__fill_1_2/VPWR
flabel metal1 8888 -2197 8941 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_42/VPWR
flabel metal1 8891 -1664 8942 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_42/VGND
rlabel comment 8963 -1644 8963 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_42/tapvpwrvgnd_1
rlabel metal1 8871 -1692 8963 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_42/VGND
rlabel metal1 8871 -2236 8963 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_42/VPWR
flabel metal1 9348 -2197 9401 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_43/VPWR
flabel metal1 9351 -1664 9402 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_43/VGND
rlabel comment 9423 -1644 9423 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_43/tapvpwrvgnd_1
rlabel metal1 9331 -1692 9423 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_43/VGND
rlabel metal1 9331 -2236 9423 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_43/VPWR
flabel metal1 10176 -2197 10229 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_44/VPWR
flabel metal1 10179 -1664 10230 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_44/VGND
rlabel comment 10251 -1644 10251 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_44/tapvpwrvgnd_1
rlabel metal1 10159 -1692 10251 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_44/VGND
rlabel metal1 10159 -2236 10251 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_44/VPWR
flabel locali 11383 -1899 11417 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/A
flabel locali 10737 -2103 10771 -2069 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X
flabel locali 10737 -2035 10771 -2001 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X
flabel locali 10737 -1967 10771 -1933 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X
flabel locali 10737 -1899 10771 -1865 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X
flabel locali 10737 -1831 10771 -1797 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X
flabel locali 10737 -1763 10771 -1729 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X
flabel pwell 11383 -1661 11417 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/VNB
flabel nwell 11383 -2205 11417 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/VPB
flabel metal1 11383 -1661 11417 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/VGND
flabel metal1 11383 -2205 11417 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_17/VPWR
rlabel comment 11447 -1644 11447 -1644 8 sky130_fd_sc_hd__clkdlybuf4s50_1_17/clkdlybuf4s50_1
rlabel metal1 10711 -1692 11447 -1596 5 sky130_fd_sc_hd__clkdlybuf4s50_1_17/VGND
rlabel metal1 10711 -2236 11447 -2140 5 sky130_fd_sc_hd__clkdlybuf4s50_1_17/VPWR
flabel metal1 11936 -1661 11970 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_25/VGND
flabel metal1 11936 -2205 11970 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_25/VPWR
flabel nwell 11936 -2205 11970 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_25/VPB
flabel pwell 11936 -1661 11970 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_25/VNB
rlabel comment 11999 -1644 11999 -1644 8 sky130_fd_sc_hd__decap_4_25/decap_4
rlabel metal1 11631 -1692 11999 -1596 5 sky130_fd_sc_hd__decap_4_25/VGND
rlabel metal1 11631 -2236 11999 -2140 5 sky130_fd_sc_hd__decap_4_25/VPWR
flabel metal1 10653 -2201 10689 -2171 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_4/VPWR
flabel metal1 10653 -1660 10689 -1631 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_4/VGND
flabel nwell 10660 -2195 10680 -2178 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_4/VPB
flabel pwell 10659 -1655 10683 -1633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_4/VNB
rlabel comment 10711 -1644 10711 -1644 8 sky130_fd_sc_hd__fill_1_4/fill_1
rlabel metal1 10619 -1692 10711 -1596 5 sky130_fd_sc_hd__fill_1_4/VGND
rlabel metal1 10619 -2236 10711 -2140 5 sky130_fd_sc_hd__fill_1_4/VPWR
flabel metal1 11573 -2201 11609 -2171 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_5/VPWR
flabel metal1 11573 -1660 11609 -1631 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_5/VGND
flabel nwell 11580 -2195 11600 -2178 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_5/VPB
flabel pwell 11579 -1655 11603 -1633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_5/VNB
rlabel comment 11631 -1644 11631 -1644 8 sky130_fd_sc_hd__fill_1_5/fill_1
rlabel metal1 11539 -1692 11631 -1596 5 sky130_fd_sc_hd__fill_1_5/VGND
rlabel metal1 11539 -2236 11631 -2140 5 sky130_fd_sc_hd__fill_1_5/VPWR
flabel metal1 12668 -1654 12700 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_0/VGND
flabel metal1 12668 -2199 12706 -2167 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_0/VPWR
flabel nwell 12658 -2197 12715 -2166 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_0/VPB
flabel pwell 12665 -1654 12709 -1620 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_0/VNB
rlabel comment 12735 -1644 12735 -1644 8 sky130_fd_sc_hd__fill_8_0/fill_8
rlabel metal1 11999 -1692 12735 -1596 5 sky130_fd_sc_hd__fill_8_0/VGND
rlabel metal1 11999 -2236 12735 -2140 5 sky130_fd_sc_hd__fill_8_0/VPWR
flabel metal1 11464 -2197 11517 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_45/VPWR
flabel metal1 11467 -1664 11518 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_45/VGND
rlabel comment 11539 -1644 11539 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_45/tapvpwrvgnd_1
rlabel metal1 11447 -1692 11539 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_45/VGND
rlabel metal1 11447 -2236 11539 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_45/VPWR
flabel locali 15248 -1967 15282 -1933 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/X
flabel locali 15340 -1967 15374 -1933 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/X
flabel locali 15340 -1899 15374 -1865 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/X
flabel locali 15248 -1899 15282 -1865 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/X
flabel locali 15248 -1831 15282 -1797 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/X
flabel locali 15340 -1831 15374 -1797 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/X
flabel locali 13684 -1831 13718 -1797 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/A
flabel locali 13684 -1899 13718 -1865 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/A
flabel pwell 13684 -1661 13718 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/VNB
flabel pwell 13701 -1644 13701 -1644 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/VNB
flabel nwell 13684 -2205 13718 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/VPB
flabel nwell 13701 -2188 13701 -2188 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/VPB
flabel metal1 13684 -1661 13718 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/VGND
flabel metal1 13684 -2205 13718 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_1/VPWR
rlabel comment 13655 -1644 13655 -1644 2 sky130_fd_sc_hd__clkbuf_16_1/clkbuf_16
rlabel metal1 13655 -1692 15495 -1596 5 sky130_fd_sc_hd__clkbuf_16_1/VGND
rlabel metal1 13655 -2236 15495 -2140 5 sky130_fd_sc_hd__clkbuf_16_1/VPWR
flabel metal1 13505 -2201 13541 -2171 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_15/VPWR
flabel metal1 13505 -1660 13541 -1631 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_15/VGND
flabel nwell 13512 -2195 13532 -2178 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_15/VPB
flabel pwell 13511 -1655 13535 -1633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_15/VNB
rlabel comment 13563 -1644 13563 -1644 8 sky130_fd_sc_hd__fill_1_15/fill_1
rlabel metal1 13471 -1692 13563 -1596 5 sky130_fd_sc_hd__fill_1_15/VGND
rlabel metal1 13471 -2236 13563 -2140 5 sky130_fd_sc_hd__fill_1_15/VPWR
flabel metal1 13404 -1654 13436 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_1/VGND
flabel metal1 13404 -2199 13442 -2167 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_1/VPWR
flabel nwell 13394 -2197 13451 -2166 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_1/VPB
flabel pwell 13401 -1654 13445 -1620 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_1/VNB
rlabel comment 13471 -1644 13471 -1644 8 sky130_fd_sc_hd__fill_8_1/fill_8
rlabel metal1 12735 -1692 13471 -1596 5 sky130_fd_sc_hd__fill_8_1/VGND
rlabel metal1 12735 -2236 13471 -2140 5 sky130_fd_sc_hd__fill_8_1/VPWR
flabel metal1 13580 -2197 13633 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_117/VPWR
flabel metal1 13583 -1664 13634 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_117/VGND
rlabel comment 13655 -1644 13655 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_117/tapvpwrvgnd_1
rlabel metal1 13563 -1692 13655 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_117/VGND
rlabel metal1 13563 -2236 13655 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_117/VPWR
flabel metal1 16628 -1661 16662 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_5/VGND
flabel metal1 16628 -2205 16662 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_5/VPWR
flabel nwell 16628 -2205 16662 -2171 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_5/VPB
flabel pwell 16628 -1661 16662 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_5/VNB
rlabel comment 16691 -1644 16691 -1644 8 sky130_fd_sc_hd__decap_12_5/decap_12
rlabel metal1 15587 -1692 16691 -1596 5 sky130_fd_sc_hd__decap_12_5/VGND
rlabel metal1 15587 -2236 16691 -2140 5 sky130_fd_sc_hd__decap_12_5/VPWR
flabel metal1 15512 -2197 15565 -2168 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_128/VPWR
flabel metal1 15515 -1664 15566 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_128/VGND
rlabel comment 15587 -1644 15587 -1644 8 sky130_fd_sc_hd__tapvpwrvgnd_1_128/tapvpwrvgnd_1
rlabel metal1 15495 -1692 15587 -1596 5 sky130_fd_sc_hd__tapvpwrvgnd_1_128/VGND
rlabel metal1 15495 -2236 15587 -2140 5 sky130_fd_sc_hd__tapvpwrvgnd_1_128/VPWR
flabel metal1 -1588 -1117 -1554 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_2/VPWR
flabel metal1 -1588 -1661 -1554 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_2/VGND
flabel nwell -1588 -1117 -1554 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_2/VPB
flabel pwell -1588 -1661 -1554 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_2/VNB
rlabel comment -1617 -1644 -1617 -1644 4 sky130_fd_sc_hd__decap_8_2/decap_8
rlabel metal1 -1617 -1692 -881 -1596 1 sky130_fd_sc_hd__decap_8_2/VGND
rlabel metal1 -1617 -1148 -881 -1052 1 sky130_fd_sc_hd__decap_8_2/VPWR
flabel metal1 -2968 -1117 -2934 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_68/VPWR
flabel metal1 -2968 -1661 -2934 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_68/VGND
flabel nwell -2968 -1117 -2934 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_68/VPB
flabel pwell -2968 -1661 -2934 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_68/VNB
rlabel comment -2997 -1644 -2997 -1644 4 sky130_fd_sc_hd__decap_8_68/decap_8
rlabel metal1 -2997 -1692 -2261 -1596 1 sky130_fd_sc_hd__decap_8_68/VGND
rlabel metal1 -2997 -1148 -2261 -1052 1 sky130_fd_sc_hd__decap_8_68/VPWR
flabel metal1 -1781 -1658 -1728 -1626 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_5/VGND
flabel metal1 -1780 -1114 -1728 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_5/VPWR
flabel nwell -1773 -1109 -1739 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_5/VPB
flabel pwell -1770 -1654 -1738 -1632 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_5/VNB
rlabel comment -1801 -1644 -1801 -1644 4 sky130_fd_sc_hd__fill_2_5/fill_2
rlabel metal1 -1801 -1692 -1617 -1596 1 sky130_fd_sc_hd__fill_2_5/VGND
rlabel metal1 -1801 -1148 -1617 -1052 1 sky130_fd_sc_hd__fill_2_5/VPWR
flabel metal1 -2135 -1654 -2112 -1635 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_19/VGND
flabel metal1 -2135 -1109 -2115 -1092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_19/VPWR
flabel nwell -2134 -1114 -2109 -1088 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_19/VPB
flabel pwell -2134 -1656 -2112 -1632 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_19/VNB
rlabel comment -2169 -1644 -2169 -1644 4 sky130_fd_sc_hd__fill_4_19/fill_4
rlabel metal1 -2169 -1692 -1801 -1596 1 sky130_fd_sc_hd__fill_4_19/VGND
rlabel metal1 -2169 -1148 -1801 -1052 1 sky130_fd_sc_hd__fill_4_19/VPWR
flabel metal1 -2239 -1120 -2186 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_533/VPWR
flabel metal1 -2240 -1662 -2189 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_533/VGND
rlabel comment -2261 -1644 -2261 -1644 4 sky130_fd_sc_hd__tapvpwrvgnd_1_533/tapvpwrvgnd_1
rlabel metal1 -2261 -1692 -2169 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_533/VGND
rlabel metal1 -2261 -1148 -2169 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_533/VPWR
flabel locali 437 -1423 471 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A
flabel locali 1083 -1219 1117 -1185 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X
flabel locali 1083 -1287 1117 -1253 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X
flabel locali 1083 -1355 1117 -1321 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X
flabel locali 1083 -1423 1117 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X
flabel locali 1083 -1491 1117 -1457 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X
flabel locali 1083 -1559 1117 -1525 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X
flabel pwell 437 -1661 471 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/VNB
flabel nwell 437 -1117 471 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/VPB
flabel metal1 437 -1661 471 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/VGND
flabel metal1 437 -1117 471 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_44/VPWR
rlabel comment 407 -1644 407 -1644 4 sky130_fd_sc_hd__clkdlybuf4s50_1_44/clkdlybuf4s50_1
rlabel metal1 407 -1692 1143 -1596 1 sky130_fd_sc_hd__clkdlybuf4s50_1_44/VGND
rlabel metal1 407 -1148 1143 -1052 1 sky130_fd_sc_hd__clkdlybuf4s50_1_44/VPWR
flabel metal1 252 -1661 286 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_55/VGND
flabel metal1 252 -1117 286 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_55/VPWR
flabel nwell 252 -1117 286 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_55/VPB
flabel pwell 252 -1661 286 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_55/VNB
rlabel comment 315 -1644 315 -1644 6 sky130_fd_sc_hd__decap_4_55/decap_4
rlabel metal1 -53 -1692 315 -1596 1 sky130_fd_sc_hd__decap_4_55/VGND
rlabel metal1 -53 -1148 315 -1052 1 sky130_fd_sc_hd__decap_4_55/VPWR
flabel metal1 -852 -1117 -818 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_3/VPWR
flabel metal1 -852 -1661 -818 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_3/VGND
flabel nwell -852 -1117 -818 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_3/VPB
flabel pwell -852 -1661 -818 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_3/VNB
rlabel comment -881 -1644 -881 -1644 4 sky130_fd_sc_hd__decap_8_3/decap_8
rlabel metal1 -881 -1692 -145 -1596 1 sky130_fd_sc_hd__decap_8_3/VGND
rlabel metal1 -881 -1148 -145 -1052 1 sky130_fd_sc_hd__decap_8_3/VPWR
flabel metal1 332 -1120 385 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_98/VPWR
flabel metal1 335 -1662 386 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_98/VGND
rlabel comment 407 -1644 407 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_98/tapvpwrvgnd_1
rlabel metal1 315 -1692 407 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_98/VGND
rlabel metal1 315 -1148 407 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_98/VPWR
flabel metal1 -128 -1120 -75 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_99/VPWR
flabel metal1 -125 -1662 -74 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_99/VGND
rlabel comment -53 -1644 -53 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_99/tapvpwrvgnd_1
rlabel metal1 -145 -1692 -53 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_99/VGND
rlabel metal1 -145 -1148 -53 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_99/VPWR
flabel metal1 2828 -1661 2862 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_26/VGND
flabel metal1 2828 -1117 2862 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_26/VPWR
flabel nwell 2828 -1117 2862 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_26/VPB
flabel pwell 2828 -1661 2862 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_26/VNB
rlabel comment 2891 -1644 2891 -1644 6 sky130_fd_sc_hd__decap_4_26/decap_4
rlabel metal1 2523 -1692 2891 -1596 1 sky130_fd_sc_hd__decap_4_26/VGND
rlabel metal1 2523 -1148 2891 -1052 1 sky130_fd_sc_hd__decap_4_26/VPWR
flabel metal1 1540 -1661 1574 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_54/VGND
flabel metal1 1540 -1117 1574 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_54/VPWR
flabel nwell 1540 -1117 1574 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_54/VPB
flabel pwell 1540 -1661 1574 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_54/VNB
rlabel comment 1603 -1644 1603 -1644 6 sky130_fd_sc_hd__decap_4_54/decap_4
rlabel metal1 1235 -1692 1603 -1596 1 sky130_fd_sc_hd__decap_4_54/VGND
rlabel metal1 1235 -1148 1603 -1052 1 sky130_fd_sc_hd__decap_4_54/VPWR
flabel metal1 1724 -1117 1758 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_92/VPWR
flabel metal1 1724 -1661 1758 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_92/VGND
flabel nwell 1724 -1117 1758 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_92/VPB
flabel pwell 1724 -1661 1758 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_92/VNB
rlabel comment 1695 -1644 1695 -1644 4 sky130_fd_sc_hd__decap_8_92/decap_8
rlabel metal1 1695 -1692 2431 -1596 1 sky130_fd_sc_hd__decap_8_92/VGND
rlabel metal1 1695 -1148 2431 -1052 1 sky130_fd_sc_hd__decap_8_92/VPWR
flabel metal1 2448 -1120 2501 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_46/VPWR
flabel metal1 2451 -1662 2502 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_46/VGND
rlabel comment 2523 -1644 2523 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_46/tapvpwrvgnd_1
rlabel metal1 2431 -1692 2523 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_46/VGND
rlabel metal1 2431 -1148 2523 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_46/VPWR
flabel metal1 1160 -1120 1213 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_96/VPWR
flabel metal1 1163 -1662 1214 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_96/VGND
rlabel comment 1235 -1644 1235 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_96/tapvpwrvgnd_1
rlabel metal1 1143 -1692 1235 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_96/VGND
rlabel metal1 1143 -1148 1235 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_96/VPWR
flabel metal1 1620 -1120 1673 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_97/VPWR
flabel metal1 1623 -1662 1674 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_97/VGND
rlabel comment 1695 -1644 1695 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_97/tapvpwrvgnd_1
rlabel metal1 1603 -1692 1695 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_97/VGND
rlabel metal1 1603 -1148 1695 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_97/VPWR
flabel locali 3013 -1423 3047 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A
flabel locali 3659 -1219 3693 -1185 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/X
flabel locali 3659 -1287 3693 -1253 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/X
flabel locali 3659 -1355 3693 -1321 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/X
flabel locali 3659 -1423 3693 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/X
flabel locali 3659 -1491 3693 -1457 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/X
flabel locali 3659 -1559 3693 -1525 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/X
flabel pwell 3013 -1661 3047 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/VNB
flabel nwell 3013 -1117 3047 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/VPB
flabel metal1 3013 -1661 3047 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/VGND
flabel metal1 3013 -1117 3047 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_18/VPWR
rlabel comment 2983 -1644 2983 -1644 4 sky130_fd_sc_hd__clkdlybuf4s50_1_18/clkdlybuf4s50_1
rlabel metal1 2983 -1692 3719 -1596 1 sky130_fd_sc_hd__clkdlybuf4s50_1_18/VGND
rlabel metal1 2983 -1148 3719 -1052 1 sky130_fd_sc_hd__clkdlybuf4s50_1_18/VPWR
flabel metal1 4116 -1661 4150 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_27/VGND
flabel metal1 4116 -1117 4150 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_27/VPWR
flabel nwell 4116 -1117 4150 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_27/VPB
flabel pwell 4116 -1661 4150 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_27/VNB
rlabel comment 4179 -1644 4179 -1644 6 sky130_fd_sc_hd__decap_4_27/decap_4
rlabel metal1 3811 -1692 4179 -1596 1 sky130_fd_sc_hd__decap_4_27/VGND
rlabel metal1 3811 -1148 4179 -1052 1 sky130_fd_sc_hd__decap_4_27/VPWR
flabel metal1 4300 -1117 4334 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_107/VPWR
flabel metal1 4300 -1661 4334 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_107/VGND
flabel nwell 4300 -1117 4334 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_107/VPB
flabel pwell 4300 -1661 4334 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_107/VNB
rlabel comment 4271 -1644 4271 -1644 4 sky130_fd_sc_hd__decap_8_107/decap_8
rlabel metal1 4271 -1692 5007 -1596 1 sky130_fd_sc_hd__decap_8_107/VGND
rlabel metal1 4271 -1148 5007 -1052 1 sky130_fd_sc_hd__decap_8_107/VPWR
flabel metal1 2908 -1120 2961 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_47/VPWR
flabel metal1 2911 -1662 2962 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_47/VGND
rlabel comment 2983 -1644 2983 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_47/tapvpwrvgnd_1
rlabel metal1 2891 -1692 2983 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_47/VGND
rlabel metal1 2891 -1148 2983 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_47/VPWR
flabel metal1 3736 -1120 3789 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_48/VPWR
flabel metal1 3739 -1662 3790 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_48/VGND
rlabel comment 3811 -1644 3811 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_48/tapvpwrvgnd_1
rlabel metal1 3719 -1692 3811 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_48/VGND
rlabel metal1 3719 -1148 3811 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_48/VPWR
flabel metal1 4196 -1120 4249 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_49/VPWR
flabel metal1 4199 -1662 4250 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_49/VGND
rlabel comment 4271 -1644 4271 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_49/tapvpwrvgnd_1
rlabel metal1 4179 -1692 4271 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_49/VGND
rlabel metal1 4179 -1148 4271 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_49/VPWR
flabel locali 5589 -1423 5623 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A
flabel locali 6235 -1219 6269 -1185 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/X
flabel locali 6235 -1287 6269 -1253 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/X
flabel locali 6235 -1355 6269 -1321 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/X
flabel locali 6235 -1423 6269 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/X
flabel locali 6235 -1491 6269 -1457 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/X
flabel locali 6235 -1559 6269 -1525 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/X
flabel pwell 5589 -1661 5623 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/VNB
flabel nwell 5589 -1117 5623 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/VPB
flabel metal1 5589 -1661 5623 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/VGND
flabel metal1 5589 -1117 5623 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_20/VPWR
rlabel comment 5559 -1644 5559 -1644 4 sky130_fd_sc_hd__clkdlybuf4s50_1_20/clkdlybuf4s50_1
rlabel metal1 5559 -1692 6295 -1596 1 sky130_fd_sc_hd__clkdlybuf4s50_1_20/VGND
rlabel metal1 5559 -1148 6295 -1052 1 sky130_fd_sc_hd__clkdlybuf4s50_1_20/VPWR
flabel metal1 5404 -1661 5438 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_28/VGND
flabel metal1 5404 -1117 5438 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_28/VPWR
flabel nwell 5404 -1117 5438 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_28/VPB
flabel pwell 5404 -1661 5438 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_28/VNB
rlabel comment 5467 -1644 5467 -1644 6 sky130_fd_sc_hd__decap_4_28/decap_4
rlabel metal1 5099 -1692 5467 -1596 1 sky130_fd_sc_hd__decap_4_28/VGND
rlabel metal1 5099 -1148 5467 -1052 1 sky130_fd_sc_hd__decap_4_28/VPWR
flabel metal1 6692 -1661 6726 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_29/VGND
flabel metal1 6692 -1117 6726 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_29/VPWR
flabel nwell 6692 -1117 6726 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_29/VPB
flabel pwell 6692 -1661 6726 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_29/VNB
rlabel comment 6755 -1644 6755 -1644 6 sky130_fd_sc_hd__decap_4_29/decap_4
rlabel metal1 6387 -1692 6755 -1596 1 sky130_fd_sc_hd__decap_4_29/VGND
rlabel metal1 6387 -1148 6755 -1052 1 sky130_fd_sc_hd__decap_4_29/VPWR
flabel metal1 5484 -1120 5537 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_50/VPWR
flabel metal1 5487 -1662 5538 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_50/VGND
rlabel comment 5559 -1644 5559 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_50/tapvpwrvgnd_1
rlabel metal1 5467 -1692 5559 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_50/VGND
rlabel metal1 5467 -1148 5559 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_50/VPWR
flabel metal1 5024 -1120 5077 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_51/VPWR
flabel metal1 5027 -1662 5078 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_51/VGND
rlabel comment 5099 -1644 5099 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_51/tapvpwrvgnd_1
rlabel metal1 5007 -1692 5099 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_51/VGND
rlabel metal1 5007 -1148 5099 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_51/VPWR
flabel metal1 6312 -1120 6365 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_52/VPWR
flabel metal1 6315 -1662 6366 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_52/VGND
rlabel comment 6387 -1644 6387 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_52/tapvpwrvgnd_1
rlabel metal1 6295 -1692 6387 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_52/VGND
rlabel metal1 6295 -1148 6387 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_52/VPWR
flabel locali 8165 -1423 8199 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A
flabel locali 8811 -1219 8845 -1185 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/X
flabel locali 8811 -1287 8845 -1253 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/X
flabel locali 8811 -1355 8845 -1321 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/X
flabel locali 8811 -1423 8845 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/X
flabel locali 8811 -1491 8845 -1457 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/X
flabel locali 8811 -1559 8845 -1525 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/X
flabel pwell 8165 -1661 8199 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/VNB
flabel nwell 8165 -1117 8199 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/VPB
flabel metal1 8165 -1661 8199 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/VGND
flabel metal1 8165 -1117 8199 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_22/VPWR
rlabel comment 8135 -1644 8135 -1644 4 sky130_fd_sc_hd__clkdlybuf4s50_1_22/clkdlybuf4s50_1
rlabel metal1 8135 -1692 8871 -1596 1 sky130_fd_sc_hd__clkdlybuf4s50_1_22/VGND
rlabel metal1 8135 -1148 8871 -1052 1 sky130_fd_sc_hd__clkdlybuf4s50_1_22/VPWR
flabel metal1 7980 -1661 8014 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_30/VGND
flabel metal1 7980 -1117 8014 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_30/VPWR
flabel nwell 7980 -1117 8014 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_30/VPB
flabel pwell 7980 -1661 8014 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_30/VNB
rlabel comment 8043 -1644 8043 -1644 6 sky130_fd_sc_hd__decap_4_30/decap_4
rlabel metal1 7675 -1692 8043 -1596 1 sky130_fd_sc_hd__decap_4_30/VGND
rlabel metal1 7675 -1148 8043 -1052 1 sky130_fd_sc_hd__decap_4_30/VPWR
flabel metal1 6876 -1117 6910 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_120/VPWR
flabel metal1 6876 -1661 6910 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_120/VGND
flabel nwell 6876 -1117 6910 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_120/VPB
flabel pwell 6876 -1661 6910 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_120/VNB
rlabel comment 6847 -1644 6847 -1644 4 sky130_fd_sc_hd__decap_8_120/decap_8
rlabel metal1 6847 -1692 7583 -1596 1 sky130_fd_sc_hd__decap_8_120/VGND
rlabel metal1 6847 -1148 7583 -1052 1 sky130_fd_sc_hd__decap_8_120/VPWR
flabel metal1 6772 -1120 6825 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_53/VPWR
flabel metal1 6775 -1662 6826 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_53/VGND
rlabel comment 6847 -1644 6847 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_53/tapvpwrvgnd_1
rlabel metal1 6755 -1692 6847 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_53/VGND
rlabel metal1 6755 -1148 6847 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_53/VPWR
flabel metal1 7600 -1120 7653 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_54/VPWR
flabel metal1 7603 -1662 7654 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_54/VGND
rlabel comment 7675 -1644 7675 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_54/tapvpwrvgnd_1
rlabel metal1 7583 -1692 7675 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_54/VGND
rlabel metal1 7583 -1148 7675 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_54/VPWR
flabel metal1 8060 -1120 8113 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_55/VPWR
flabel metal1 8063 -1662 8114 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_55/VGND
rlabel comment 8135 -1644 8135 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_55/tapvpwrvgnd_1
rlabel metal1 8043 -1692 8135 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_55/VGND
rlabel metal1 8043 -1148 8135 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_55/VPWR
flabel metal1 9268 -1661 9302 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_31/VGND
flabel metal1 9268 -1117 9302 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_31/VPWR
flabel nwell 9268 -1117 9302 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_31/VPB
flabel pwell 9268 -1661 9302 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_31/VNB
rlabel comment 9331 -1644 9331 -1644 6 sky130_fd_sc_hd__decap_4_31/decap_4
rlabel metal1 8963 -1692 9331 -1596 1 sky130_fd_sc_hd__decap_4_31/VGND
rlabel metal1 8963 -1148 9331 -1052 1 sky130_fd_sc_hd__decap_4_31/VPWR
flabel metal1 10648 -1661 10682 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_32/VGND
flabel metal1 10648 -1117 10682 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_32/VPWR
flabel nwell 10648 -1117 10682 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_32/VPB
flabel pwell 10648 -1661 10682 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_32/VNB
rlabel comment 10711 -1644 10711 -1644 6 sky130_fd_sc_hd__decap_4_32/decap_4
rlabel metal1 10343 -1692 10711 -1596 1 sky130_fd_sc_hd__decap_4_32/VGND
rlabel metal1 10343 -1148 10711 -1052 1 sky130_fd_sc_hd__decap_4_32/VPWR
flabel metal1 9452 -1117 9486 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_130/VPWR
flabel metal1 9452 -1661 9486 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_130/VGND
flabel nwell 9452 -1117 9486 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_130/VPB
flabel pwell 9452 -1661 9486 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_130/VNB
rlabel comment 9423 -1644 9423 -1644 4 sky130_fd_sc_hd__decap_8_130/decap_8
rlabel metal1 9423 -1692 10159 -1596 1 sky130_fd_sc_hd__decap_8_130/VGND
rlabel metal1 9423 -1148 10159 -1052 1 sky130_fd_sc_hd__decap_8_130/VPWR
flabel metal1 10285 -1117 10321 -1087 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_6/VPWR
flabel metal1 10285 -1657 10321 -1628 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_6/VGND
flabel nwell 10292 -1110 10312 -1093 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_6/VPB
flabel pwell 10291 -1655 10315 -1633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_6/VNB
rlabel comment 10343 -1644 10343 -1644 6 sky130_fd_sc_hd__fill_1_6/fill_1
rlabel metal1 10251 -1692 10343 -1596 1 sky130_fd_sc_hd__fill_1_6/VGND
rlabel metal1 10251 -1148 10343 -1052 1 sky130_fd_sc_hd__fill_1_6/VPWR
flabel metal1 8888 -1120 8941 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_56/VPWR
flabel metal1 8891 -1662 8942 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_56/VGND
rlabel comment 8963 -1644 8963 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_56/tapvpwrvgnd_1
rlabel metal1 8871 -1692 8963 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_56/VGND
rlabel metal1 8871 -1148 8963 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_56/VPWR
flabel metal1 9348 -1120 9401 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_57/VPWR
flabel metal1 9351 -1662 9402 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_57/VGND
rlabel comment 9423 -1644 9423 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_57/tapvpwrvgnd_1
rlabel metal1 9331 -1692 9423 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_57/VGND
rlabel metal1 9331 -1148 9423 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_57/VPWR
flabel metal1 10176 -1120 10229 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_58/VPWR
flabel metal1 10179 -1662 10230 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_58/VGND
rlabel comment 10251 -1644 10251 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_58/tapvpwrvgnd_1
rlabel metal1 10159 -1692 10251 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_58/VGND
rlabel metal1 10159 -1148 10251 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_58/VPWR
flabel locali 10741 -1423 10775 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A
flabel locali 11387 -1219 11421 -1185 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
flabel locali 11387 -1287 11421 -1253 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
flabel locali 11387 -1355 11421 -1321 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
flabel locali 11387 -1423 11421 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
flabel locali 11387 -1491 11421 -1457 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
flabel locali 11387 -1559 11421 -1525 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
flabel pwell 10741 -1661 10775 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/VNB
flabel nwell 10741 -1117 10775 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/VPB
flabel metal1 10741 -1661 10775 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/VGND
flabel metal1 10741 -1117 10775 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_24/VPWR
rlabel comment 10711 -1644 10711 -1644 4 sky130_fd_sc_hd__clkdlybuf4s50_1_24/clkdlybuf4s50_1
rlabel metal1 10711 -1692 11447 -1596 1 sky130_fd_sc_hd__clkdlybuf4s50_1_24/VGND
rlabel metal1 10711 -1148 11447 -1052 1 sky130_fd_sc_hd__clkdlybuf4s50_1_24/VPWR
flabel metal1 11936 -1661 11970 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_33/VGND
flabel metal1 11936 -1117 11970 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_33/VPWR
flabel nwell 11936 -1117 11970 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_33/VPB
flabel pwell 11936 -1661 11970 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_33/VNB
rlabel comment 11999 -1644 11999 -1644 6 sky130_fd_sc_hd__decap_4_33/decap_4
rlabel metal1 11631 -1692 11999 -1596 1 sky130_fd_sc_hd__decap_4_33/VGND
rlabel metal1 11631 -1148 11999 -1052 1 sky130_fd_sc_hd__decap_4_33/VPWR
flabel metal1 10653 -1117 10689 -1087 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_7/VPWR
flabel metal1 10653 -1657 10689 -1628 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_7/VGND
flabel nwell 10660 -1110 10680 -1093 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_7/VPB
flabel pwell 10659 -1655 10683 -1633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_7/VNB
rlabel comment 10711 -1644 10711 -1644 6 sky130_fd_sc_hd__fill_1_7/fill_1
rlabel metal1 10619 -1692 10711 -1596 1 sky130_fd_sc_hd__fill_1_7/VGND
rlabel metal1 10619 -1148 10711 -1052 1 sky130_fd_sc_hd__fill_1_7/VPWR
flabel metal1 11573 -1117 11609 -1087 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_8/VPWR
flabel metal1 11573 -1657 11609 -1628 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_8/VGND
flabel nwell 11580 -1110 11600 -1093 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_8/VPB
flabel pwell 11579 -1655 11603 -1633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_8/VNB
rlabel comment 11631 -1644 11631 -1644 6 sky130_fd_sc_hd__fill_1_8/fill_1
rlabel metal1 11539 -1692 11631 -1596 1 sky130_fd_sc_hd__fill_1_8/VGND
rlabel metal1 11539 -1148 11631 -1052 1 sky130_fd_sc_hd__fill_1_8/VPWR
flabel metal1 12033 -1654 12056 -1635 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_2/VGND
flabel metal1 12033 -1109 12053 -1092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_2/VPWR
flabel nwell 12034 -1114 12059 -1088 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_2/VPB
flabel pwell 12034 -1656 12056 -1632 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_2/VNB
rlabel comment 11999 -1644 11999 -1644 4 sky130_fd_sc_hd__fill_4_2/fill_4
rlabel metal1 11999 -1692 12367 -1596 1 sky130_fd_sc_hd__fill_4_2/VGND
rlabel metal1 11999 -1148 12367 -1052 1 sky130_fd_sc_hd__fill_4_2/VPWR
flabel metal1 11464 -1120 11517 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_59/VPWR
flabel metal1 11467 -1662 11518 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_59/VGND
rlabel comment 11539 -1644 11539 -1644 6 sky130_fd_sc_hd__tapvpwrvgnd_1_59/tapvpwrvgnd_1
rlabel metal1 11447 -1692 11539 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_59/VGND
rlabel metal1 11447 -1148 11539 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_59/VPWR
flabel locali 15248 -1355 15282 -1321 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/X
flabel locali 15340 -1355 15374 -1321 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/X
flabel locali 15340 -1423 15374 -1389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/X
flabel locali 15248 -1423 15282 -1389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/X
flabel locali 15248 -1491 15282 -1457 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/X
flabel locali 15340 -1491 15374 -1457 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/X
flabel locali 13684 -1491 13718 -1457 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/A
flabel locali 13684 -1423 13718 -1389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/A
flabel pwell 13684 -1661 13718 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/VNB
flabel pwell 13701 -1644 13701 -1644 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/VNB
flabel nwell 13684 -1117 13718 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/VPB
flabel nwell 13701 -1100 13701 -1100 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/VPB
flabel metal1 13684 -1661 13718 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/VGND
flabel metal1 13684 -1117 13718 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_2/VPWR
rlabel comment 13655 -1644 13655 -1644 4 sky130_fd_sc_hd__clkbuf_16_2/clkbuf_16
rlabel metal1 13655 -1692 15495 -1596 1 sky130_fd_sc_hd__clkbuf_16_2/VGND
rlabel metal1 13655 -1148 15495 -1052 1 sky130_fd_sc_hd__clkbuf_16_2/VPWR
flabel locali 12672 -1423 12706 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/A
flabel locali 12764 -1423 12798 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/A
flabel locali 13040 -1491 13074 -1457 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/Y
flabel locali 12580 -1423 12614 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/A
flabel locali 13040 -1355 13074 -1321 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/Y
flabel locali 12948 -1423 12982 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/A
flabel locali 12856 -1423 12890 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/A
flabel locali 13040 -1423 13074 -1389 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_1/Y
flabel pwell 12488 -1661 12522 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_1/VNB
flabel nwell 12488 -1117 12522 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_1/VPB
flabel metal1 12488 -1117 12522 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_1/VPWR
flabel metal1 12488 -1661 12522 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_1/VGND
rlabel comment 12459 -1644 12459 -1644 4 sky130_fd_sc_hd__clkinv_4_1/clkinv_4
rlabel metal1 12459 -1692 13103 -1596 1 sky130_fd_sc_hd__clkinv_4_1/VGND
rlabel metal1 12459 -1148 13103 -1052 1 sky130_fd_sc_hd__clkinv_4_1/VPWR
flabel metal1 13224 -1661 13258 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_62/VGND
flabel metal1 13224 -1117 13258 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_62/VPWR
flabel nwell 13224 -1117 13258 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_62/VPB
flabel pwell 13224 -1661 13258 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_62/VNB
rlabel comment 13195 -1644 13195 -1644 4 sky130_fd_sc_hd__decap_4_62/decap_4
rlabel metal1 13195 -1692 13563 -1596 1 sky130_fd_sc_hd__decap_4_62/VGND
rlabel metal1 13195 -1148 13563 -1052 1 sky130_fd_sc_hd__decap_4_62/VPWR
flabel metal1 13125 -1120 13178 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_111/VPWR
flabel metal1 13124 -1662 13175 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_111/VGND
rlabel comment 13103 -1644 13103 -1644 4 sky130_fd_sc_hd__tapvpwrvgnd_1_111/tapvpwrvgnd_1
rlabel metal1 13103 -1692 13195 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_111/VGND
rlabel metal1 13103 -1148 13195 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_111/VPWR
flabel metal1 13585 -1120 13638 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_112/VPWR
flabel metal1 13584 -1662 13635 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_112/VGND
rlabel comment 13563 -1644 13563 -1644 4 sky130_fd_sc_hd__tapvpwrvgnd_1_112/tapvpwrvgnd_1
rlabel metal1 13563 -1692 13655 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_112/VGND
rlabel metal1 13563 -1148 13655 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_112/VPWR
flabel metal1 12389 -1120 12442 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_113/VPWR
flabel metal1 12388 -1662 12439 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_113/VGND
rlabel comment 12367 -1644 12367 -1644 4 sky130_fd_sc_hd__tapvpwrvgnd_1_113/tapvpwrvgnd_1
rlabel metal1 12367 -1692 12459 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_113/VGND
rlabel metal1 12367 -1148 12459 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_113/VPWR
flabel metal1 15616 -1661 15650 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_3/VGND
flabel metal1 15616 -1117 15650 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_3/VPWR
flabel nwell 15616 -1117 15650 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_3/VPB
flabel pwell 15616 -1661 15650 -1627 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_3/VNB
rlabel comment 15587 -1644 15587 -1644 4 sky130_fd_sc_hd__decap_12_3/decap_12
rlabel metal1 15587 -1692 16691 -1596 1 sky130_fd_sc_hd__decap_12_3/VGND
rlabel metal1 15587 -1148 16691 -1052 1 sky130_fd_sc_hd__decap_12_3/VPWR
flabel metal1 15517 -1120 15570 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_123/VPWR
flabel metal1 15516 -1662 15567 -1624 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_123/VGND
rlabel comment 15495 -1644 15495 -1644 4 sky130_fd_sc_hd__tapvpwrvgnd_1_123/tapvpwrvgnd_1
rlabel metal1 15495 -1692 15587 -1596 1 sky130_fd_sc_hd__tapvpwrvgnd_1_123/VGND
rlabel metal1 15495 -1148 15587 -1052 1 sky130_fd_sc_hd__tapvpwrvgnd_1_123/VPWR
flabel metal1 -944 -1117 -910 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_1/VPWR
flabel metal1 -944 -573 -910 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_1/VGND
flabel nwell -944 -1117 -910 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_1/VPB
flabel pwell -944 -573 -910 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_1/VNB
rlabel comment -881 -556 -881 -556 8 sky130_fd_sc_hd__decap_8_1/decap_8
rlabel metal1 -1617 -604 -881 -508 5 sky130_fd_sc_hd__decap_8_1/VGND
rlabel metal1 -1617 -1148 -881 -1052 5 sky130_fd_sc_hd__decap_8_1/VPWR
flabel metal1 -2324 -1117 -2290 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_67/VPWR
flabel metal1 -2324 -573 -2290 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_67/VGND
flabel nwell -2324 -1117 -2290 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_67/VPB
flabel pwell -2324 -573 -2290 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_67/VNB
rlabel comment -2261 -556 -2261 -556 8 sky130_fd_sc_hd__decap_8_67/decap_8
rlabel metal1 -2997 -604 -2261 -508 5 sky130_fd_sc_hd__decap_8_67/VGND
rlabel metal1 -2997 -1148 -2261 -1052 5 sky130_fd_sc_hd__decap_8_67/VPWR
flabel metal1 -1690 -574 -1637 -542 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VGND
flabel metal1 -1690 -1117 -1638 -1086 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VPWR
flabel nwell -1679 -1109 -1645 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VPB
flabel pwell -1680 -568 -1648 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VNB
rlabel comment -1617 -556 -1617 -556 8 sky130_fd_sc_hd__fill_2_0/fill_2
rlabel metal1 -1801 -604 -1617 -508 5 sky130_fd_sc_hd__fill_2_0/VGND
rlabel metal1 -1801 -1148 -1617 -1052 5 sky130_fd_sc_hd__fill_2_0/VPWR
flabel metal1 -1858 -565 -1835 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_18/VGND
flabel metal1 -1855 -1108 -1835 -1091 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_18/VPWR
flabel nwell -1861 -1112 -1836 -1086 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_18/VPB
flabel pwell -1858 -568 -1836 -544 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_18/VNB
rlabel comment -1801 -556 -1801 -556 8 sky130_fd_sc_hd__fill_4_18/fill_4
rlabel metal1 -2169 -604 -1801 -508 5 sky130_fd_sc_hd__fill_4_18/VGND
rlabel metal1 -2169 -1148 -1801 -1052 5 sky130_fd_sc_hd__fill_4_18/VPWR
flabel metal1 -2244 -1109 -2191 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_532/VPWR
flabel metal1 -2241 -576 -2190 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_532/VGND
rlabel comment -2169 -556 -2169 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_532/tapvpwrvgnd_1
rlabel metal1 -2261 -604 -2169 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_532/VGND
rlabel metal1 -2261 -1148 -2169 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_532/VPWR
flabel locali 1079 -811 1113 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A
flabel locali 433 -1015 467 -981 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X
flabel locali 433 -947 467 -913 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X
flabel locali 433 -879 467 -845 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X
flabel locali 433 -811 467 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X
flabel locali 433 -743 467 -709 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X
flabel locali 433 -675 467 -641 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/X
flabel pwell 1079 -573 1113 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/VNB
flabel nwell 1079 -1117 1113 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/VPB
flabel metal1 1079 -573 1113 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/VGND
flabel metal1 1079 -1117 1113 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_42/VPWR
rlabel comment 1143 -556 1143 -556 8 sky130_fd_sc_hd__clkdlybuf4s50_1_42/clkdlybuf4s50_1
rlabel metal1 407 -604 1143 -508 5 sky130_fd_sc_hd__clkdlybuf4s50_1_42/VGND
rlabel metal1 407 -1148 1143 -1052 5 sky130_fd_sc_hd__clkdlybuf4s50_1_42/VPWR
flabel metal1 252 -573 286 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_53/VGND
flabel metal1 252 -1117 286 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_53/VPWR
flabel nwell 252 -1117 286 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_53/VPB
flabel pwell 252 -573 286 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_53/VNB
rlabel comment 315 -556 315 -556 8 sky130_fd_sc_hd__decap_4_53/decap_4
rlabel metal1 -53 -604 315 -508 5 sky130_fd_sc_hd__decap_4_53/VGND
rlabel metal1 -53 -1148 315 -1052 5 sky130_fd_sc_hd__decap_4_53/VPWR
flabel metal1 -208 -1117 -174 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_0/VPWR
flabel metal1 -208 -573 -174 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_0/VGND
flabel nwell -208 -1117 -174 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_0/VPB
flabel pwell -208 -573 -174 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_0/VNB
rlabel comment -145 -556 -145 -556 8 sky130_fd_sc_hd__decap_8_0/decap_8
rlabel metal1 -881 -604 -145 -508 5 sky130_fd_sc_hd__decap_8_0/VGND
rlabel metal1 -881 -1148 -145 -1052 5 sky130_fd_sc_hd__decap_8_0/VPWR
flabel metal1 332 -1109 385 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_94/VPWR
flabel metal1 335 -576 386 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_94/VGND
rlabel comment 407 -556 407 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_94/tapvpwrvgnd_1
rlabel metal1 315 -604 407 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_94/VGND
rlabel metal1 315 -1148 407 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_94/VPWR
flabel metal1 -128 -1109 -75 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_95/VPWR
flabel metal1 -125 -576 -74 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_95/VGND
rlabel comment -53 -556 -53 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_95/tapvpwrvgnd_1
rlabel metal1 -145 -604 -53 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_95/VGND
rlabel metal1 -145 -1148 -53 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_95/VPWR
flabel metal1 2828 -573 2862 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_17/VGND
flabel metal1 2828 -1117 2862 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_17/VPWR
flabel nwell 2828 -1117 2862 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_17/VPB
flabel pwell 2828 -573 2862 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_17/VNB
rlabel comment 2891 -556 2891 -556 8 sky130_fd_sc_hd__decap_4_17/decap_4
rlabel metal1 2523 -604 2891 -508 5 sky130_fd_sc_hd__decap_4_17/VGND
rlabel metal1 2523 -1148 2891 -1052 5 sky130_fd_sc_hd__decap_4_17/VPWR
flabel metal1 1540 -573 1574 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_52/VGND
flabel metal1 1540 -1117 1574 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_52/VPWR
flabel nwell 1540 -1117 1574 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_52/VPB
flabel pwell 1540 -573 1574 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_52/VNB
rlabel comment 1603 -556 1603 -556 8 sky130_fd_sc_hd__decap_4_52/decap_4
rlabel metal1 1235 -604 1603 -508 5 sky130_fd_sc_hd__decap_4_52/VGND
rlabel metal1 1235 -1148 1603 -1052 5 sky130_fd_sc_hd__decap_4_52/VPWR
flabel metal1 2368 -1117 2402 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_91/VPWR
flabel metal1 2368 -573 2402 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_91/VGND
flabel nwell 2368 -1117 2402 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_91/VPB
flabel pwell 2368 -573 2402 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_91/VNB
rlabel comment 2431 -556 2431 -556 8 sky130_fd_sc_hd__decap_8_91/decap_8
rlabel metal1 1695 -604 2431 -508 5 sky130_fd_sc_hd__decap_8_91/VGND
rlabel metal1 1695 -1148 2431 -1052 5 sky130_fd_sc_hd__decap_8_91/VPWR
flabel metal1 2448 -1109 2501 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_31/VPWR
flabel metal1 2451 -576 2502 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_31/VGND
rlabel comment 2523 -556 2523 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_31/tapvpwrvgnd_1
rlabel metal1 2431 -604 2523 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_31/VGND
rlabel metal1 2431 -1148 2523 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_31/VPWR
flabel metal1 1160 -1109 1213 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_92/VPWR
flabel metal1 1163 -576 1214 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_92/VGND
rlabel comment 1235 -556 1235 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_92/tapvpwrvgnd_1
rlabel metal1 1143 -604 1235 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_92/VGND
rlabel metal1 1143 -1148 1235 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_92/VPWR
flabel metal1 1620 -1109 1673 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_93/VPWR
flabel metal1 1623 -576 1674 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_93/VGND
rlabel comment 1695 -556 1695 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_93/tapvpwrvgnd_1
rlabel metal1 1603 -604 1695 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_93/VGND
rlabel metal1 1603 -1148 1695 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_93/VPWR
flabel locali 3655 -811 3689 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/A
flabel locali 3009 -1015 3043 -981 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X
flabel locali 3009 -947 3043 -913 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X
flabel locali 3009 -879 3043 -845 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X
flabel locali 3009 -811 3043 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X
flabel locali 3009 -743 3043 -709 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X
flabel locali 3009 -675 3043 -641 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/X
flabel pwell 3655 -573 3689 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/VNB
flabel nwell 3655 -1117 3689 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/VPB
flabel metal1 3655 -573 3689 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/VGND
flabel metal1 3655 -1117 3689 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_10/VPWR
rlabel comment 3719 -556 3719 -556 8 sky130_fd_sc_hd__clkdlybuf4s50_1_10/clkdlybuf4s50_1
rlabel metal1 2983 -604 3719 -508 5 sky130_fd_sc_hd__clkdlybuf4s50_1_10/VGND
rlabel metal1 2983 -1148 3719 -1052 5 sky130_fd_sc_hd__clkdlybuf4s50_1_10/VPWR
flabel metal1 4116 -573 4150 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_16/VGND
flabel metal1 4116 -1117 4150 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_16/VPWR
flabel nwell 4116 -1117 4150 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_16/VPB
flabel pwell 4116 -573 4150 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_16/VNB
rlabel comment 4179 -556 4179 -556 8 sky130_fd_sc_hd__decap_4_16/decap_4
rlabel metal1 3811 -604 4179 -508 5 sky130_fd_sc_hd__decap_4_16/VGND
rlabel metal1 3811 -1148 4179 -1052 5 sky130_fd_sc_hd__decap_4_16/VPWR
flabel metal1 4944 -1117 4978 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_108/VPWR
flabel metal1 4944 -573 4978 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_108/VGND
flabel nwell 4944 -1117 4978 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_108/VPB
flabel pwell 4944 -573 4978 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_108/VNB
rlabel comment 5007 -556 5007 -556 8 sky130_fd_sc_hd__decap_8_108/decap_8
rlabel metal1 4271 -604 5007 -508 5 sky130_fd_sc_hd__decap_8_108/VGND
rlabel metal1 4271 -1148 5007 -1052 5 sky130_fd_sc_hd__decap_8_108/VPWR
flabel metal1 4196 -1109 4249 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_28/VPWR
flabel metal1 4199 -576 4250 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_28/VGND
rlabel comment 4271 -556 4271 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_28/tapvpwrvgnd_1
rlabel metal1 4179 -604 4271 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_28/VGND
rlabel metal1 4179 -1148 4271 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_28/VPWR
flabel metal1 3736 -1109 3789 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_29/VPWR
flabel metal1 3739 -576 3790 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_29/VGND
rlabel comment 3811 -556 3811 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_29/tapvpwrvgnd_1
rlabel metal1 3719 -604 3811 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_29/VGND
rlabel metal1 3719 -1148 3811 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_29/VPWR
flabel metal1 2908 -1109 2961 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_30/VPWR
flabel metal1 2911 -576 2962 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_30/VGND
rlabel comment 2983 -556 2983 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_30/tapvpwrvgnd_1
rlabel metal1 2891 -604 2983 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_30/VGND
rlabel metal1 2891 -1148 2983 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_30/VPWR
flabel locali 6231 -811 6265 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A
flabel locali 5585 -1015 5619 -981 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
flabel locali 5585 -947 5619 -913 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
flabel locali 5585 -879 5619 -845 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
flabel locali 5585 -811 5619 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
flabel locali 5585 -743 5619 -709 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
flabel locali 5585 -675 5619 -641 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
flabel pwell 6231 -573 6265 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/VNB
flabel nwell 6231 -1117 6265 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/VPB
flabel metal1 6231 -573 6265 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/VGND
flabel metal1 6231 -1117 6265 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_8/VPWR
rlabel comment 6295 -556 6295 -556 8 sky130_fd_sc_hd__clkdlybuf4s50_1_8/clkdlybuf4s50_1
rlabel metal1 5559 -604 6295 -508 5 sky130_fd_sc_hd__clkdlybuf4s50_1_8/VGND
rlabel metal1 5559 -1148 6295 -1052 5 sky130_fd_sc_hd__clkdlybuf4s50_1_8/VPWR
flabel metal1 6692 -573 6726 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_14/VGND
flabel metal1 6692 -1117 6726 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_14/VPWR
flabel nwell 6692 -1117 6726 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_14/VPB
flabel pwell 6692 -573 6726 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_14/VNB
rlabel comment 6755 -556 6755 -556 8 sky130_fd_sc_hd__decap_4_14/decap_4
rlabel metal1 6387 -604 6755 -508 5 sky130_fd_sc_hd__decap_4_14/VGND
rlabel metal1 6387 -1148 6755 -1052 5 sky130_fd_sc_hd__decap_4_14/VPWR
flabel metal1 5404 -573 5438 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_15/VGND
flabel metal1 5404 -1117 5438 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_15/VPWR
flabel nwell 5404 -1117 5438 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_15/VPB
flabel pwell 5404 -573 5438 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_15/VNB
rlabel comment 5467 -556 5467 -556 8 sky130_fd_sc_hd__decap_4_15/decap_4
rlabel metal1 5099 -604 5467 -508 5 sky130_fd_sc_hd__decap_4_15/VGND
rlabel metal1 5099 -1148 5467 -1052 5 sky130_fd_sc_hd__decap_4_15/VPWR
flabel metal1 6312 -1109 6365 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_25/VPWR
flabel metal1 6315 -576 6366 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_25/VGND
rlabel comment 6387 -556 6387 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_25/tapvpwrvgnd_1
rlabel metal1 6295 -604 6387 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_25/VGND
rlabel metal1 6295 -1148 6387 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_25/VPWR
flabel metal1 5484 -1109 5537 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_26/VPWR
flabel metal1 5487 -576 5538 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_26/VGND
rlabel comment 5559 -556 5559 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_26/tapvpwrvgnd_1
rlabel metal1 5467 -604 5559 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_26/VGND
rlabel metal1 5467 -1148 5559 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_26/VPWR
flabel metal1 5024 -1109 5077 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_27/VPWR
flabel metal1 5027 -576 5078 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_27/VGND
rlabel comment 5099 -556 5099 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_27/tapvpwrvgnd_1
rlabel metal1 5007 -604 5099 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_27/VGND
rlabel metal1 5007 -1148 5099 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_27/VPWR
flabel locali 8807 -811 8841 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A
flabel locali 8161 -1015 8195 -981 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/X
flabel locali 8161 -947 8195 -913 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/X
flabel locali 8161 -879 8195 -845 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/X
flabel locali 8161 -811 8195 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/X
flabel locali 8161 -743 8195 -709 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/X
flabel locali 8161 -675 8195 -641 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/X
flabel pwell 8807 -573 8841 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/VNB
flabel nwell 8807 -1117 8841 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/VPB
flabel metal1 8807 -573 8841 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/VGND
flabel metal1 8807 -1117 8841 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_6/VPWR
rlabel comment 8871 -556 8871 -556 8 sky130_fd_sc_hd__clkdlybuf4s50_1_6/clkdlybuf4s50_1
rlabel metal1 8135 -604 8871 -508 5 sky130_fd_sc_hd__clkdlybuf4s50_1_6/VGND
rlabel metal1 8135 -1148 8871 -1052 5 sky130_fd_sc_hd__clkdlybuf4s50_1_6/VPWR
flabel metal1 7980 -573 8014 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_13/VGND
flabel metal1 7980 -1117 8014 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_13/VPWR
flabel nwell 7980 -1117 8014 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_13/VPB
flabel pwell 7980 -573 8014 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_13/VNB
rlabel comment 8043 -556 8043 -556 8 sky130_fd_sc_hd__decap_4_13/decap_4
rlabel metal1 7675 -604 8043 -508 5 sky130_fd_sc_hd__decap_4_13/VGND
rlabel metal1 7675 -1148 8043 -1052 5 sky130_fd_sc_hd__decap_4_13/VPWR
flabel metal1 7520 -1117 7554 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_119/VPWR
flabel metal1 7520 -573 7554 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_119/VGND
flabel nwell 7520 -1117 7554 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_119/VPB
flabel pwell 7520 -573 7554 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_119/VNB
rlabel comment 7583 -556 7583 -556 8 sky130_fd_sc_hd__decap_8_119/decap_8
rlabel metal1 6847 -604 7583 -508 5 sky130_fd_sc_hd__decap_8_119/VGND
rlabel metal1 6847 -1148 7583 -1052 5 sky130_fd_sc_hd__decap_8_119/VPWR
flabel metal1 8060 -1109 8113 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_22/VPWR
flabel metal1 8063 -576 8114 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_22/VGND
rlabel comment 8135 -556 8135 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_22/tapvpwrvgnd_1
rlabel metal1 8043 -604 8135 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_22/VGND
rlabel metal1 8043 -1148 8135 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_22/VPWR
flabel metal1 7600 -1109 7653 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_23/VPWR
flabel metal1 7603 -576 7654 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_23/VGND
rlabel comment 7675 -556 7675 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_23/tapvpwrvgnd_1
rlabel metal1 7583 -604 7675 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_23/VGND
rlabel metal1 7583 -1148 7675 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_23/VPWR
flabel metal1 6772 -1109 6825 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_24/VPWR
flabel metal1 6775 -576 6826 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_24/VGND
rlabel comment 6847 -556 6847 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_24/tapvpwrvgnd_1
rlabel metal1 6755 -604 6847 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_24/VGND
rlabel metal1 6755 -1148 6847 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_24/VPWR
flabel metal1 10648 -573 10682 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_11/VGND
flabel metal1 10648 -1117 10682 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_11/VPWR
flabel nwell 10648 -1117 10682 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_11/VPB
flabel pwell 10648 -573 10682 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_11/VNB
rlabel comment 10711 -556 10711 -556 8 sky130_fd_sc_hd__decap_4_11/decap_4
rlabel metal1 10343 -604 10711 -508 5 sky130_fd_sc_hd__decap_4_11/VGND
rlabel metal1 10343 -1148 10711 -1052 5 sky130_fd_sc_hd__decap_4_11/VPWR
flabel metal1 9268 -573 9302 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_12/VGND
flabel metal1 9268 -1117 9302 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_12/VPWR
flabel nwell 9268 -1117 9302 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_12/VPB
flabel pwell 9268 -573 9302 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_12/VNB
rlabel comment 9331 -556 9331 -556 8 sky130_fd_sc_hd__decap_4_12/decap_4
rlabel metal1 8963 -604 9331 -508 5 sky130_fd_sc_hd__decap_4_12/VGND
rlabel metal1 8963 -1148 9331 -1052 5 sky130_fd_sc_hd__decap_4_12/VPWR
flabel metal1 10096 -1117 10130 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_129/VPWR
flabel metal1 10096 -573 10130 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_129/VGND
flabel nwell 10096 -1117 10130 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_129/VPB
flabel pwell 10096 -573 10130 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_129/VNB
rlabel comment 10159 -556 10159 -556 8 sky130_fd_sc_hd__decap_8_129/decap_8
rlabel metal1 9423 -604 10159 -508 5 sky130_fd_sc_hd__decap_8_129/VGND
rlabel metal1 9423 -1148 10159 -1052 5 sky130_fd_sc_hd__decap_8_129/VPWR
flabel metal1 10285 -1113 10321 -1083 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_3/VPWR
flabel metal1 10285 -572 10321 -543 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_3/VGND
flabel nwell 10292 -1107 10312 -1090 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_3/VPB
flabel pwell 10291 -567 10315 -545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_3/VNB
rlabel comment 10343 -556 10343 -556 8 sky130_fd_sc_hd__fill_1_3/fill_1
rlabel metal1 10251 -604 10343 -508 5 sky130_fd_sc_hd__fill_1_3/VGND
rlabel metal1 10251 -1148 10343 -1052 5 sky130_fd_sc_hd__fill_1_3/VPWR
flabel metal1 10176 -1109 10229 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_19/VPWR
flabel metal1 10179 -576 10230 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_19/VGND
rlabel comment 10251 -556 10251 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_19/tapvpwrvgnd_1
rlabel metal1 10159 -604 10251 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_19/VGND
rlabel metal1 10159 -1148 10251 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_19/VPWR
flabel metal1 9348 -1109 9401 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_20/VPWR
flabel metal1 9351 -576 9402 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_20/VGND
rlabel comment 9423 -556 9423 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_20/tapvpwrvgnd_1
rlabel metal1 9331 -604 9423 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_20/VGND
rlabel metal1 9331 -1148 9423 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_20/VPWR
flabel metal1 8888 -1109 8941 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_21/VPWR
flabel metal1 8891 -576 8942 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_21/VGND
rlabel comment 8963 -556 8963 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_21/tapvpwrvgnd_1
rlabel metal1 8871 -604 8963 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_21/VGND
rlabel metal1 8871 -1148 8963 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_21/VPWR
flabel locali 11383 -811 11417 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A
flabel locali 10737 -1015 10771 -981 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X
flabel locali 10737 -947 10771 -913 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X
flabel locali 10737 -879 10771 -845 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X
flabel locali 10737 -811 10771 -777 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X
flabel locali 10737 -743 10771 -709 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X
flabel locali 10737 -675 10771 -641 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X
flabel pwell 11383 -573 11417 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/VNB
flabel nwell 11383 -1117 11417 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/VPB
flabel metal1 11383 -573 11417 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/VGND
flabel metal1 11383 -1117 11417 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_5/VPWR
rlabel comment 11447 -556 11447 -556 8 sky130_fd_sc_hd__clkdlybuf4s50_1_5/clkdlybuf4s50_1
rlabel metal1 10711 -604 11447 -508 5 sky130_fd_sc_hd__clkdlybuf4s50_1_5/VGND
rlabel metal1 10711 -1148 11447 -1052 5 sky130_fd_sc_hd__clkdlybuf4s50_1_5/VPWR
flabel metal1 11936 -573 11970 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_10/VGND
flabel metal1 11936 -1117 11970 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_10/VPWR
flabel nwell 11936 -1117 11970 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_10/VPB
flabel pwell 11936 -573 11970 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_10/VNB
rlabel comment 11999 -556 11999 -556 8 sky130_fd_sc_hd__decap_4_10/decap_4
rlabel metal1 11631 -604 11999 -508 5 sky130_fd_sc_hd__decap_4_10/VGND
rlabel metal1 11631 -1148 11999 -1052 5 sky130_fd_sc_hd__decap_4_10/VPWR
flabel metal1 11573 -1113 11609 -1083 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_0/VPWR
flabel metal1 11573 -572 11609 -543 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_0/VGND
flabel nwell 11580 -1107 11600 -1090 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_0/VPB
flabel pwell 11579 -567 11603 -545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_0/VNB
rlabel comment 11631 -556 11631 -556 8 sky130_fd_sc_hd__fill_1_0/fill_1
rlabel metal1 11539 -604 11631 -508 5 sky130_fd_sc_hd__fill_1_0/VGND
rlabel metal1 11539 -1148 11631 -1052 5 sky130_fd_sc_hd__fill_1_0/VPWR
flabel metal1 10653 -1113 10689 -1083 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_1/VPWR
flabel metal1 10653 -572 10689 -543 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_1/VGND
flabel nwell 10660 -1107 10680 -1090 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_1/VPB
flabel pwell 10659 -567 10683 -545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_1/VNB
rlabel comment 10711 -556 10711 -556 8 sky130_fd_sc_hd__fill_1_1/fill_1
rlabel metal1 10619 -604 10711 -508 5 sky130_fd_sc_hd__fill_1_1/VGND
rlabel metal1 10619 -1148 10711 -1052 5 sky130_fd_sc_hd__fill_1_1/VPWR
flabel metal1 12668 -566 12700 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_3/VGND
flabel metal1 12668 -1111 12706 -1079 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_3/VPWR
flabel nwell 12658 -1109 12715 -1078 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_3/VPB
flabel pwell 12665 -566 12709 -532 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_3/VNB
rlabel comment 12735 -556 12735 -556 8 sky130_fd_sc_hd__fill_8_3/fill_8
rlabel metal1 11999 -604 12735 -508 5 sky130_fd_sc_hd__fill_8_3/VGND
rlabel metal1 11999 -1148 12735 -1052 5 sky130_fd_sc_hd__fill_8_3/VPWR
flabel metal1 11464 -1109 11517 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_18/VPWR
flabel metal1 11467 -576 11518 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_18/VGND
rlabel comment 11539 -556 11539 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_18/tapvpwrvgnd_1
rlabel metal1 11447 -604 11539 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_18/VGND
rlabel metal1 11447 -1148 11539 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_18/VPWR
flabel locali 15248 -879 15282 -845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/X
flabel locali 15340 -879 15374 -845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/X
flabel locali 15340 -811 15374 -777 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/X
flabel locali 15248 -811 15282 -777 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/X
flabel locali 15248 -743 15282 -709 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/X
flabel locali 15340 -743 15374 -709 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/X
flabel locali 13684 -743 13718 -709 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/A
flabel locali 13684 -811 13718 -777 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/A
flabel pwell 13684 -573 13718 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/VNB
flabel pwell 13701 -556 13701 -556 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/VNB
flabel nwell 13684 -1117 13718 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/VPB
flabel nwell 13701 -1100 13701 -1100 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/VPB
flabel metal1 13684 -573 13718 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/VGND
flabel metal1 13684 -1117 13718 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkbuf_16_0/VPWR
rlabel comment 13655 -556 13655 -556 2 sky130_fd_sc_hd__clkbuf_16_0/clkbuf_16
rlabel metal1 13655 -604 15495 -508 5 sky130_fd_sc_hd__clkbuf_16_0/VGND
rlabel metal1 13655 -1148 15495 -1052 5 sky130_fd_sc_hd__clkbuf_16_0/VPWR
flabel metal1 13505 -1113 13541 -1083 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_17/VPWR
flabel metal1 13505 -572 13541 -543 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_17/VGND
flabel nwell 13512 -1107 13532 -1090 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_17/VPB
flabel pwell 13511 -567 13535 -545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_17/VNB
rlabel comment 13563 -556 13563 -556 8 sky130_fd_sc_hd__fill_1_17/fill_1
rlabel metal1 13471 -604 13563 -508 5 sky130_fd_sc_hd__fill_1_17/VGND
rlabel metal1 13471 -1148 13563 -1052 5 sky130_fd_sc_hd__fill_1_17/VPWR
flabel metal1 13404 -566 13436 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_4/VGND
flabel metal1 13404 -1111 13442 -1079 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_4/VPWR
flabel nwell 13394 -1109 13451 -1078 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_4/VPB
flabel pwell 13401 -566 13445 -532 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_4/VNB
rlabel comment 13471 -556 13471 -556 8 sky130_fd_sc_hd__fill_8_4/fill_8
rlabel metal1 12735 -604 13471 -508 5 sky130_fd_sc_hd__fill_8_4/VGND
rlabel metal1 12735 -1148 13471 -1052 5 sky130_fd_sc_hd__fill_8_4/VPWR
flabel metal1 13580 -1109 13633 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_118/VPWR
flabel metal1 13583 -576 13634 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_118/VGND
rlabel comment 13655 -556 13655 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_118/tapvpwrvgnd_1
rlabel metal1 13563 -604 13655 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_118/VGND
rlabel metal1 13563 -1148 13655 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_118/VPWR
flabel metal1 16628 -573 16662 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_4/VGND
flabel metal1 16628 -1117 16662 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_4/VPWR
flabel nwell 16628 -1117 16662 -1083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_4/VPB
flabel pwell 16628 -573 16662 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_4/VNB
rlabel comment 16691 -556 16691 -556 8 sky130_fd_sc_hd__decap_12_4/decap_12
rlabel metal1 15587 -604 16691 -508 5 sky130_fd_sc_hd__decap_12_4/VGND
rlabel metal1 15587 -1148 16691 -1052 5 sky130_fd_sc_hd__decap_12_4/VPWR
flabel metal1 15512 -1109 15565 -1080 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_125/VPWR
flabel metal1 15515 -576 15566 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_125/VGND
rlabel comment 15587 -556 15587 -556 8 sky130_fd_sc_hd__tapvpwrvgnd_1_125/tapvpwrvgnd_1
rlabel metal1 15495 -604 15587 -508 5 sky130_fd_sc_hd__tapvpwrvgnd_1_125/VGND
rlabel metal1 15495 -1148 15587 -1052 5 sky130_fd_sc_hd__tapvpwrvgnd_1_125/VPWR
flabel metal1 -1404 -573 -1370 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VGND
flabel metal1 -1404 -29 -1370 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VPWR
flabel nwell -1404 -29 -1370 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VPB
flabel pwell -1404 -573 -1370 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_0/VNB
rlabel comment -1433 -556 -1433 -556 4 sky130_fd_sc_hd__decap_4_0/decap_4
rlabel metal1 -1433 -604 -1065 -508 1 sky130_fd_sc_hd__decap_4_0/VGND
rlabel metal1 -1433 -60 -1065 36 1 sky130_fd_sc_hd__decap_4_0/VPWR
flabel metal1 -2968 -29 -2934 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_46/VPWR
flabel metal1 -2968 -573 -2934 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_46/VGND
flabel nwell -2968 -29 -2934 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_46/VPB
flabel pwell -2968 -573 -2934 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_46/VNB
rlabel comment -2997 -556 -2997 -556 4 sky130_fd_sc_hd__decap_8_46/decap_8
rlabel metal1 -2997 -604 -2261 -508 1 sky130_fd_sc_hd__decap_8_46/VGND
rlabel metal1 -2997 -60 -2261 36 1 sky130_fd_sc_hd__decap_8_46/VPWR
flabel metal1 -1597 -570 -1544 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_15/VGND
flabel metal1 -1596 -26 -1544 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_15/VPWR
flabel nwell -1589 -21 -1555 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_15/VPB
flabel pwell -1586 -566 -1554 -544 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_15/VNB
rlabel comment -1617 -556 -1617 -556 4 sky130_fd_sc_hd__fill_2_15/fill_2
rlabel metal1 -1617 -604 -1433 -508 1 sky130_fd_sc_hd__fill_2_15/VGND
rlabel metal1 -1617 -60 -1433 36 1 sky130_fd_sc_hd__fill_2_15/VPWR
flabel metal1 -1690 -570 -1637 -538 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_16/VGND
flabel metal1 -1690 -26 -1638 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_16/VPWR
flabel nwell -1679 -21 -1645 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_16/VPB
flabel pwell -1680 -566 -1648 -544 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_16/VNB
rlabel comment -1617 -556 -1617 -556 6 sky130_fd_sc_hd__fill_2_16/fill_2
rlabel metal1 -1801 -604 -1617 -508 1 sky130_fd_sc_hd__fill_2_16/VGND
rlabel metal1 -1801 -60 -1617 36 1 sky130_fd_sc_hd__fill_2_16/VPWR
flabel metal1 -2135 -566 -2112 -547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_16/VGND
flabel metal1 -2135 -21 -2115 -4 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_16/VPWR
flabel nwell -2134 -26 -2109 0 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_16/VPB
flabel pwell -2134 -568 -2112 -544 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_16/VNB
rlabel comment -2169 -556 -2169 -556 4 sky130_fd_sc_hd__fill_4_16/fill_4
rlabel metal1 -2169 -604 -1801 -508 1 sky130_fd_sc_hd__fill_4_16/VGND
rlabel metal1 -2169 -60 -1801 36 1 sky130_fd_sc_hd__fill_4_16/VPWR
flabel metal1 -2239 -32 -2186 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_531/VPWR
flabel metal1 -2240 -574 -2189 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_531/VGND
rlabel comment -2261 -556 -2261 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_531/tapvpwrvgnd_1
rlabel metal1 -2261 -604 -2169 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_531/VGND
rlabel metal1 -2261 -60 -2169 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_531/VPWR
flabel locali 68 -335 102 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/A
flabel locali 160 -335 194 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/A
flabel locali 436 -403 470 -369 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/Y
flabel locali -24 -335 10 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/A
flabel locali 436 -267 470 -233 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/Y
flabel locali 344 -335 378 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/A
flabel locali 252 -335 286 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/A
flabel locali 436 -335 470 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkinv_4_0/Y
flabel pwell -116 -573 -82 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_0/VNB
flabel nwell -116 -29 -82 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_0/VPB
flabel metal1 -116 -29 -82 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_0/VPWR
flabel metal1 -116 -573 -82 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_4_0/VGND
rlabel comment -145 -556 -145 -556 4 sky130_fd_sc_hd__clkinv_4_0/clkinv_4
rlabel metal1 -145 -604 499 -508 1 sky130_fd_sc_hd__clkinv_4_0/VGND
rlabel metal1 -145 -60 499 36 1 sky130_fd_sc_hd__clkinv_4_0/VPWR
flabel metal1 620 -573 654 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VGND
flabel metal1 620 -29 654 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VPWR
flabel nwell 620 -29 654 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VPB
flabel pwell 620 -573 654 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_1/VNB
rlabel comment 591 -556 591 -556 4 sky130_fd_sc_hd__decap_4_1/decap_4
rlabel metal1 591 -604 959 -508 1 sky130_fd_sc_hd__decap_4_1/VGND
rlabel metal1 591 -60 959 36 1 sky130_fd_sc_hd__decap_4_1/VPWR
flabel metal1 -576 -573 -542 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_8/VGND
flabel metal1 -576 -29 -542 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_8/VPWR
flabel nwell -576 -29 -542 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_8/VPB
flabel pwell -576 -573 -542 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_8/VNB
rlabel comment -605 -556 -605 -556 4 sky130_fd_sc_hd__decap_4_8/decap_4
rlabel metal1 -605 -604 -237 -508 1 sky130_fd_sc_hd__decap_4_8/VGND
rlabel metal1 -605 -60 -237 36 1 sky130_fd_sc_hd__decap_4_8/VPWR
flabel locali -853 -471 -819 -437 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali -853 -403 -819 -369 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali -853 -335 -819 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali -945 -335 -911 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/B
flabel locali -761 -335 -727 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/A
flabel nwell -945 -29 -911 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPB
flabel pwell -945 -573 -911 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VNB
flabel metal1 -945 -573 -911 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VGND
flabel metal1 -945 -29 -911 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPWR
rlabel comment -973 -556 -973 -556 4 sky130_fd_sc_hd__nand2_1_0/nand2_1
rlabel metal1 -973 -604 -697 -508 1 sky130_fd_sc_hd__nand2_1_0/VGND
rlabel metal1 -973 -60 -697 36 1 sky130_fd_sc_hd__nand2_1_0/VPWR
flabel metal1 -1043 -32 -990 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 -1044 -574 -993 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment -1065 -556 -1065 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
rlabel metal1 -1065 -604 -973 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel metal1 -1065 -60 -973 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 -675 -32 -622 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 -676 -574 -625 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment -697 -556 -697 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
rlabel metal1 -697 -604 -605 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel metal1 -697 -60 -605 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 -215 -32 -162 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR
flabel metal1 -216 -574 -165 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
rlabel comment -237 -556 -237 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_2/tapvpwrvgnd_1
rlabel metal1 -237 -604 -145 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
rlabel metal1 -237 -60 -145 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR
flabel metal1 521 -32 574 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VPWR
flabel metal1 520 -574 571 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VGND
rlabel comment 499 -556 499 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_4/tapvpwrvgnd_1
rlabel metal1 499 -604 591 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VGND
rlabel metal1 499 -60 591 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VPWR
flabel locali 2369 -335 2403 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/A
flabel locali 3015 -131 3049 -97 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/X
flabel locali 3015 -199 3049 -165 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/X
flabel locali 3015 -267 3049 -233 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/X
flabel locali 3015 -335 3049 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/X
flabel locali 3015 -403 3049 -369 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/X
flabel locali 3015 -471 3049 -437 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/X
flabel pwell 2369 -573 2403 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/VNB
flabel nwell 2369 -29 2403 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/VPB
flabel metal1 2369 -573 2403 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/VGND
flabel metal1 2369 -29 2403 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_0/VPWR
rlabel comment 2339 -556 2339 -556 4 sky130_fd_sc_hd__clkdlybuf4s50_1_0/clkdlybuf4s50_1
rlabel metal1 2339 -604 3075 -508 1 sky130_fd_sc_hd__clkdlybuf4s50_1_0/VGND
rlabel metal1 2339 -60 3075 36 1 sky130_fd_sc_hd__clkdlybuf4s50_1_0/VPWR
flabel locali 1264 -403 1298 -369 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/Y
flabel locali 1264 -335 1298 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/Y
flabel locali 1172 -267 1206 -233 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/Y
flabel locali 1172 -335 1206 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/Y
flabel locali 1172 -403 1206 -369 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/Y
flabel locali 1080 -471 1114 -437 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/A
flabel locali 1080 -403 1114 -369 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/A
flabel locali 1080 -335 1114 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__clkinv_1_0/A
flabel nwell 1080 -29 1114 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_0/VPB
flabel pwell 1080 -573 1114 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_0/VNB
flabel metal1 1080 -573 1114 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_0/VGND
flabel metal1 1080 -29 1114 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkinv_1_0/VPWR
rlabel comment 1051 -556 1051 -556 4 sky130_fd_sc_hd__clkinv_1_0/clkinv_1
rlabel metal1 1051 -604 1327 -508 1 sky130_fd_sc_hd__clkinv_1_0/VGND
rlabel metal1 1051 -60 1327 36 1 sky130_fd_sc_hd__clkinv_1_0/VPWR
flabel metal1 1448 -573 1482 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_2/VGND
flabel metal1 1448 -29 1482 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_2/VPWR
flabel nwell 1448 -29 1482 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_2/VPB
flabel pwell 1448 -573 1482 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_2/VNB
rlabel comment 1419 -556 1419 -556 4 sky130_fd_sc_hd__decap_4_2/decap_4
rlabel metal1 1419 -604 1787 -508 1 sky130_fd_sc_hd__decap_4_2/VGND
rlabel metal1 1419 -60 1787 36 1 sky130_fd_sc_hd__decap_4_2/VPWR
flabel metal1 1908 -573 1942 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_3/VGND
flabel metal1 1908 -29 1942 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_3/VPWR
flabel nwell 1908 -29 1942 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_3/VPB
flabel pwell 1908 -573 1942 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_3/VNB
rlabel comment 1879 -556 1879 -556 4 sky130_fd_sc_hd__decap_4_3/decap_4
rlabel metal1 1879 -604 2247 -508 1 sky130_fd_sc_hd__decap_4_3/VGND
rlabel metal1 1879 -60 2247 36 1 sky130_fd_sc_hd__decap_4_3/VPWR
flabel metal1 981 -32 1034 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VPWR
flabel metal1 980 -574 1031 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VGND
rlabel comment 959 -556 959 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_5/tapvpwrvgnd_1
rlabel metal1 959 -604 1051 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VGND
rlabel metal1 959 -60 1051 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VPWR
flabel metal1 1349 -32 1402 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VPWR
flabel metal1 1348 -574 1399 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VGND
rlabel comment 1327 -556 1327 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_6/tapvpwrvgnd_1
rlabel metal1 1327 -604 1419 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VGND
rlabel metal1 1327 -60 1419 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VPWR
flabel metal1 1809 -32 1862 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VPWR
flabel metal1 1808 -574 1859 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VGND
rlabel comment 1787 -556 1787 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_7/tapvpwrvgnd_1
rlabel metal1 1787 -604 1879 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VGND
rlabel metal1 1787 -60 1879 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VPWR
flabel metal1 2269 -32 2322 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VPWR
flabel metal1 2268 -574 2319 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VGND
rlabel comment 2247 -556 2247 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_8/tapvpwrvgnd_1
rlabel metal1 2247 -604 2339 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VGND
rlabel metal1 2247 -60 2339 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VPWR
flabel metal1 3196 -573 3230 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_60/VGND
flabel metal1 3196 -29 3230 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_60/VPWR
flabel nwell 3196 -29 3230 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_60/VPB
flabel pwell 3196 -573 3230 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_60/VNB
rlabel comment 3167 -556 3167 -556 4 sky130_fd_sc_hd__decap_4_60/decap_4
rlabel metal1 3167 -604 3535 -508 1 sky130_fd_sc_hd__decap_4_60/VGND
rlabel metal1 3167 -60 3535 36 1 sky130_fd_sc_hd__decap_4_60/VPWR
flabel metal1 4392 -573 4426 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VGND
flabel metal1 4392 -29 4426 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VPWR
flabel nwell 4392 -29 4426 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VPB
flabel pwell 4392 -573 4426 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VNB
rlabel comment 4363 -556 4363 -556 4 sky130_fd_sc_hd__decap_12_0/decap_12
rlabel metal1 4363 -604 5467 -508 1 sky130_fd_sc_hd__decap_12_0/VGND
rlabel metal1 4363 -60 5467 36 1 sky130_fd_sc_hd__decap_12_0/VPWR
flabel metal1 3662 -576 3694 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_2/VGND
flabel metal1 3656 -33 3694 -1 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_2/VPWR
flabel nwell 3647 -34 3704 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_2/VPB
flabel pwell 3653 -580 3697 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_2/VNB
rlabel comment 3627 -556 3627 -556 4 sky130_fd_sc_hd__fill_8_2/fill_8
rlabel metal1 3627 -604 4363 -508 1 sky130_fd_sc_hd__fill_8_2/VGND
rlabel metal1 3627 -60 4363 36 1 sky130_fd_sc_hd__fill_8_2/VPWR
flabel metal1 3557 -32 3610 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VPWR
flabel metal1 3556 -574 3607 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VGND
rlabel comment 3535 -556 3535 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_3/tapvpwrvgnd_1
rlabel metal1 3535 -604 3627 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VGND
rlabel metal1 3535 -60 3627 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VPWR
flabel metal1 3097 -32 3150 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_108/VPWR
flabel metal1 3096 -574 3147 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_108/VGND
rlabel comment 3075 -556 3075 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_108/tapvpwrvgnd_1
rlabel metal1 3075 -604 3167 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_108/VGND
rlabel metal1 3075 -60 3167 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_108/VPWR
flabel metal1 6416 -573 6450 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_4/VGND
flabel metal1 6416 -29 6450 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_4/VPWR
flabel nwell 6416 -29 6450 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_4/VPB
flabel pwell 6416 -573 6450 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_4/VNB
rlabel comment 6387 -556 6387 -556 4 sky130_fd_sc_hd__decap_4_4/decap_4
rlabel metal1 6387 -604 6755 -508 1 sky130_fd_sc_hd__decap_4_4/VGND
rlabel metal1 6387 -60 6755 36 1 sky130_fd_sc_hd__decap_4_4/VPWR
flabel metal1 5857 -29 5893 1 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_16/VPWR
flabel metal1 5857 -569 5893 -540 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__fill_1_16/VGND
flabel nwell 5866 -22 5886 -5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_16/VPB
flabel pwell 5863 -567 5887 -545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_1_16/VNB
rlabel comment 5835 -556 5835 -556 4 sky130_fd_sc_hd__fill_1_16/fill_1
rlabel metal1 5835 -604 5927 -508 1 sky130_fd_sc_hd__fill_1_16/VGND
rlabel metal1 5835 -60 5927 36 1 sky130_fd_sc_hd__fill_1_16/VPWR
flabel metal1 5961 -566 5984 -547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_0/VGND
flabel metal1 5961 -21 5981 -4 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_0/VPWR
flabel nwell 5962 -26 5987 0 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_0/VPB
flabel pwell 5962 -568 5984 -544 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_0/VNB
rlabel comment 5927 -556 5927 -556 4 sky130_fd_sc_hd__fill_4_0/fill_4
rlabel metal1 5927 -604 6295 -508 1 sky130_fd_sc_hd__fill_4_0/VGND
rlabel metal1 5927 -60 6295 36 1 sky130_fd_sc_hd__fill_4_0/VPWR
flabel metal1 5501 -566 5524 -547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_1/VGND
flabel metal1 5501 -21 5521 -4 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_1/VPWR
flabel nwell 5502 -26 5527 0 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_1/VPB
flabel pwell 5502 -568 5524 -544 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_4_1/VNB
rlabel comment 5467 -556 5467 -556 4 sky130_fd_sc_hd__fill_4_1/fill_4
rlabel metal1 5467 -604 5835 -508 1 sky130_fd_sc_hd__fill_4_1/VGND
rlabel metal1 5467 -60 5835 36 1 sky130_fd_sc_hd__fill_4_1/VPWR
flabel metal1 6317 -32 6370 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VPWR
flabel metal1 6316 -574 6367 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VGND
rlabel comment 6295 -556 6295 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_9/tapvpwrvgnd_1
rlabel metal1 6295 -604 6387 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VGND
rlabel metal1 6295 -60 6387 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VPWR
flabel locali 6877 -335 6911 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A
flabel locali 7523 -131 7557 -97 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/X
flabel locali 7523 -199 7557 -165 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/X
flabel locali 7523 -267 7557 -233 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/X
flabel locali 7523 -335 7557 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/X
flabel locali 7523 -403 7557 -369 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/X
flabel locali 7523 -471 7557 -437 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/X
flabel pwell 6877 -573 6911 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/VNB
flabel nwell 6877 -29 6911 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/VPB
flabel metal1 6877 -573 6911 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/VGND
flabel metal1 6877 -29 6911 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_1/VPWR
rlabel comment 6847 -556 6847 -556 4 sky130_fd_sc_hd__clkdlybuf4s50_1_1/clkdlybuf4s50_1
rlabel metal1 6847 -604 7583 -508 1 sky130_fd_sc_hd__clkdlybuf4s50_1_1/VGND
rlabel metal1 6847 -60 7583 36 1 sky130_fd_sc_hd__clkdlybuf4s50_1_1/VPWR
flabel locali 8165 -335 8199 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A
flabel locali 8811 -131 8845 -97 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/X
flabel locali 8811 -199 8845 -165 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/X
flabel locali 8811 -267 8845 -233 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/X
flabel locali 8811 -335 8845 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/X
flabel locali 8811 -403 8845 -369 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/X
flabel locali 8811 -471 8845 -437 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/X
flabel pwell 8165 -573 8199 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/VNB
flabel nwell 8165 -29 8199 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/VPB
flabel metal1 8165 -573 8199 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/VGND
flabel metal1 8165 -29 8199 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_2/VPWR
rlabel comment 8135 -556 8135 -556 4 sky130_fd_sc_hd__clkdlybuf4s50_1_2/clkdlybuf4s50_1
rlabel metal1 8135 -604 8871 -508 1 sky130_fd_sc_hd__clkdlybuf4s50_1_2/VGND
rlabel metal1 8135 -60 8871 36 1 sky130_fd_sc_hd__clkdlybuf4s50_1_2/VPWR
flabel metal1 7704 -573 7738 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_5/VGND
flabel metal1 7704 -29 7738 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_5/VPWR
flabel nwell 7704 -29 7738 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_5/VPB
flabel pwell 7704 -573 7738 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_5/VNB
rlabel comment 7675 -556 7675 -556 4 sky130_fd_sc_hd__decap_4_5/decap_4
rlabel metal1 7675 -604 8043 -508 1 sky130_fd_sc_hd__decap_4_5/VGND
rlabel metal1 7675 -60 8043 36 1 sky130_fd_sc_hd__decap_4_5/VPWR
flabel metal1 6777 -32 6830 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_10/VPWR
flabel metal1 6776 -574 6827 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_10/VGND
rlabel comment 6755 -556 6755 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_10/tapvpwrvgnd_1
rlabel metal1 6755 -604 6847 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_10/VGND
rlabel metal1 6755 -60 6847 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_10/VPWR
flabel metal1 7605 -32 7658 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_11/VPWR
flabel metal1 7604 -574 7655 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_11/VGND
rlabel comment 7583 -556 7583 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_11/tapvpwrvgnd_1
rlabel metal1 7583 -604 7675 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_11/VGND
rlabel metal1 7583 -60 7675 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_11/VPWR
flabel metal1 8065 -32 8118 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_12/VPWR
flabel metal1 8064 -574 8115 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_12/VGND
rlabel comment 8043 -556 8043 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_12/tapvpwrvgnd_1
rlabel metal1 8043 -604 8135 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_12/VGND
rlabel metal1 8043 -60 8135 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_12/VPWR
flabel locali 9453 -335 9487 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A
flabel locali 10099 -131 10133 -97 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/X
flabel locali 10099 -199 10133 -165 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/X
flabel locali 10099 -267 10133 -233 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/X
flabel locali 10099 -335 10133 -301 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/X
flabel locali 10099 -403 10133 -369 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/X
flabel locali 10099 -471 10133 -437 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/X
flabel pwell 9453 -573 9487 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/VNB
flabel nwell 9453 -29 9487 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/VPB
flabel metal1 9453 -573 9487 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/VGND
flabel metal1 9453 -29 9487 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__clkdlybuf4s50_1_3/VPWR
rlabel comment 9423 -556 9423 -556 4 sky130_fd_sc_hd__clkdlybuf4s50_1_3/clkdlybuf4s50_1
rlabel metal1 9423 -604 10159 -508 1 sky130_fd_sc_hd__clkdlybuf4s50_1_3/VGND
rlabel metal1 9423 -60 10159 36 1 sky130_fd_sc_hd__clkdlybuf4s50_1_3/VPWR
flabel metal1 8992 -573 9026 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_6/VGND
flabel metal1 8992 -29 9026 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_6/VPWR
flabel nwell 8992 -29 9026 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_6/VPB
flabel pwell 8992 -573 9026 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_6/VNB
rlabel comment 8963 -556 8963 -556 4 sky130_fd_sc_hd__decap_4_6/decap_4
rlabel metal1 8963 -604 9331 -508 1 sky130_fd_sc_hd__decap_4_6/VGND
rlabel metal1 8963 -60 9331 36 1 sky130_fd_sc_hd__decap_4_6/VPWR
flabel metal1 10280 -573 10314 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_7/VGND
flabel metal1 10280 -29 10314 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_7/VPWR
flabel nwell 10280 -29 10314 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_7/VPB
flabel pwell 10280 -573 10314 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_7/VNB
rlabel comment 10251 -556 10251 -556 4 sky130_fd_sc_hd__decap_4_7/decap_4
rlabel metal1 10251 -604 10619 -508 1 sky130_fd_sc_hd__decap_4_7/VGND
rlabel metal1 10251 -60 10619 36 1 sky130_fd_sc_hd__decap_4_7/VPWR
flabel metal1 8893 -32 8946 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_13/VPWR
flabel metal1 8892 -574 8943 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_13/VGND
rlabel comment 8871 -556 8871 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_13/tapvpwrvgnd_1
rlabel metal1 8871 -604 8963 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_13/VGND
rlabel metal1 8871 -60 8963 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_13/VPWR
flabel metal1 9353 -32 9406 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_14/VPWR
flabel metal1 9352 -574 9403 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_14/VGND
rlabel comment 9331 -556 9331 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_14/tapvpwrvgnd_1
rlabel metal1 9331 -604 9423 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_14/VGND
rlabel metal1 9331 -60 9423 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_14/VPWR
flabel metal1 10181 -32 10234 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_15/VPWR
flabel metal1 10180 -574 10231 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_15/VGND
rlabel comment 10159 -556 10159 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_15/tapvpwrvgnd_1
rlabel metal1 10159 -604 10251 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_15/VGND
rlabel metal1 10159 -60 10251 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_15/VPWR
flabel metal1 11660 -573 11694 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_9/VGND
flabel metal1 11660 -29 11694 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_9/VPWR
flabel nwell 11660 -29 11694 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_9/VPB
flabel pwell 11660 -573 11694 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_4_9/VNB
rlabel comment 11631 -556 11631 -556 4 sky130_fd_sc_hd__decap_4_9/decap_4
rlabel metal1 11631 -604 11999 -508 1 sky130_fd_sc_hd__decap_4_9/VGND
rlabel metal1 11631 -60 11999 36 1 sky130_fd_sc_hd__decap_4_9/VPWR
flabel metal1 12034 -576 12066 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_5/VGND
flabel metal1 12028 -33 12066 -1 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_5/VPWR
flabel nwell 12019 -34 12076 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_5/VPB
flabel pwell 12025 -580 12069 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_5/VNB
rlabel comment 11999 -556 11999 -556 4 sky130_fd_sc_hd__fill_8_5/fill_8
rlabel metal1 11999 -604 12735 -508 1 sky130_fd_sc_hd__fill_8_5/VGND
rlabel metal1 11999 -60 12735 36 1 sky130_fd_sc_hd__fill_8_5/VPWR
flabel locali 11109 -335 11143 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/Y
flabel locali 11109 -267 11143 -233 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/Y
flabel locali 11385 -335 11419 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/A
flabel locali 11293 -335 11327 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/A
flabel locali 11017 -335 11051 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 10925 -335 10959 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 10741 -335 10775 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 10833 -335 10867 -301 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel nwell 10741 -29 10775 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VPB
flabel pwell 10741 -573 10775 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VNB
flabel metal1 10741 -573 10775 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VGND
flabel metal1 10741 -29 10775 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VPWR
rlabel comment 10711 -556 10711 -556 4 sky130_fd_sc_hd__nand2_4_0/nand2_4
rlabel metal1 10711 -604 11539 -508 1 sky130_fd_sc_hd__nand2_4_0/VGND
rlabel metal1 10711 -60 11539 36 1 sky130_fd_sc_hd__nand2_4_0/VPWR
flabel metal1 10641 -32 10694 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_16/VPWR
flabel metal1 10640 -574 10691 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_16/VGND
rlabel comment 10619 -556 10619 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_16/tapvpwrvgnd_1
rlabel metal1 10619 -604 10711 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_16/VGND
rlabel metal1 10619 -60 10711 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_16/VPWR
flabel metal1 11561 -32 11614 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_17/VPWR
flabel metal1 11560 -574 11611 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_17/VGND
rlabel comment 11539 -556 11539 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_17/tapvpwrvgnd_1
rlabel metal1 11539 -604 11631 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_17/VGND
rlabel metal1 11539 -60 11631 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_17/VPWR
flabel metal1 13592 -573 13626 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VGND
flabel metal1 13592 -29 13626 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VPWR
flabel nwell 13592 -29 13626 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VPB
flabel pwell 13592 -573 13626 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VNB
rlabel comment 13563 -556 13563 -556 4 sky130_fd_sc_hd__decap_12_1/decap_12
rlabel metal1 13563 -604 14667 -508 1 sky130_fd_sc_hd__decap_12_1/VGND
rlabel metal1 13563 -60 14667 36 1 sky130_fd_sc_hd__decap_12_1/VPWR
flabel metal1 12770 -576 12802 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_6/VGND
flabel metal1 12764 -33 12802 -1 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_6/VPWR
flabel nwell 12755 -34 12812 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_6/VPB
flabel pwell 12761 -580 12805 -546 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_8_6/VNB
rlabel comment 12735 -556 12735 -556 4 sky130_fd_sc_hd__fill_8_6/fill_8
rlabel metal1 12735 -604 13471 -508 1 sky130_fd_sc_hd__fill_8_6/VGND
rlabel metal1 12735 -60 13471 36 1 sky130_fd_sc_hd__fill_8_6/VPWR
flabel metal1 13493 -32 13546 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_119/VPWR
flabel metal1 13492 -574 13543 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_119/VGND
rlabel comment 13471 -556 13471 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_119/tapvpwrvgnd_1
rlabel metal1 13471 -604 13563 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_119/VGND
rlabel metal1 13471 -60 13563 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_119/VPWR
flabel metal1 15984 -29 16018 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_9/VPWR
flabel metal1 15984 -573 16018 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_9/VGND
flabel nwell 15984 -29 16018 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_9/VPB
flabel pwell 15984 -573 16018 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_8_9/VNB
rlabel comment 15955 -556 15955 -556 4 sky130_fd_sc_hd__decap_8_9/decap_8
rlabel metal1 15955 -604 16691 -508 1 sky130_fd_sc_hd__decap_8_9/VGND
rlabel metal1 15955 -60 16691 36 1 sky130_fd_sc_hd__decap_8_9/VPWR
flabel metal1 14788 -573 14822 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_2/VGND
flabel metal1 14788 -29 14822 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_2/VPWR
flabel nwell 14788 -29 14822 5 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_2/VPB
flabel pwell 14788 -573 14822 -539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_2/VNB
rlabel comment 14759 -556 14759 -556 4 sky130_fd_sc_hd__decap_12_2/decap_12
rlabel metal1 14759 -604 15863 -508 1 sky130_fd_sc_hd__decap_12_2/VGND
rlabel metal1 14759 -60 15863 36 1 sky130_fd_sc_hd__decap_12_2/VPWR
flabel metal1 14689 -32 14742 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_120/VPWR
flabel metal1 14688 -574 14739 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_120/VGND
rlabel comment 14667 -556 14667 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_120/tapvpwrvgnd_1
rlabel metal1 14667 -604 14759 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_120/VGND
rlabel metal1 14667 -60 14759 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_120/VPWR
flabel metal1 15885 -32 15938 -3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_121/VPWR
flabel metal1 15884 -574 15935 -536 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_121/VGND
rlabel comment 15863 -556 15863 -556 4 sky130_fd_sc_hd__tapvpwrvgnd_1_121/tapvpwrvgnd_1
rlabel metal1 15863 -604 15955 -508 1 sky130_fd_sc_hd__tapvpwrvgnd_1_121/VGND
rlabel metal1 15863 -60 15955 36 1 sky130_fd_sc_hd__tapvpwrvgnd_1_121/VPWR
<< end >>
