* NGSPICE file created from ota_v2.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_YVTR7C a_n207_n140# a_n1039_n205# a_29_n205# a_327_n140#
+ a_n683_n205# a_n1275_n140# a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_1097_n205#
+ a_n505_n205# a_n741_n140# a_563_n205# a_861_n140# w_n1311_n241# a_919_n205# a_n327_n205#
+ a_n563_n140# a_385_n205# a_683_n140# a_n919_n140# a_n149_n205# a_1039_n140# a_n385_n140#
+ a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_327_n140# a_207_n205# a_149_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_149_n140# a_29_n205# a_n29_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_861_n140# a_741_n205# a_683_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_n140# a_n327_n205# a_n385_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1097_n205# a_1097_n205# a_1039_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n741_n140# a_n861_n205# a_n919_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n1097_n140# a_n1275_n140# a_n1275_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_683_n140# a_563_n205# a_505_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1039_n140# a_919_n205# a_861_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n29_n140# a_n149_n205# a_n207_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n563_n140# a_n683_n205# a_n741_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_741_n205# a_n149_n205# 0.01fF
C1 a_327_n140# a_505_n140# 0.06fF
C2 a_149_n140# a_683_n140# 0.02fF
C3 a_327_n140# a_n29_n140# 0.03fF
C4 a_n683_n205# a_563_n205# 0.01fF
C5 a_1097_n205# a_861_n140# 0.03fF
C6 a_n563_n140# a_505_n140# 0.01fF
C7 a_n29_n140# a_n563_n140# 0.02fF
C8 a_n207_n140# a_n385_n140# 0.06fF
C9 a_n683_n205# w_n1311_n241# 0.20fF
C10 a_n741_n140# a_n385_n140# 0.03fF
C11 a_1039_n140# a_n207_n140# 0.01fF
C12 a_741_n205# a_919_n205# 0.10fF
C13 a_n505_n205# a_n149_n205# 0.03fF
C14 a_29_n205# a_563_n205# 0.02fF
C15 a_563_n205# a_n327_n205# 0.01fF
C16 a_29_n205# w_n1311_n241# 0.19fF
C17 a_n1039_n205# a_385_n205# 0.01fF
C18 w_n1311_n241# a_n327_n205# 0.20fF
C19 a_n505_n205# a_919_n205# 0.01fF
C20 w_n1311_n241# a_n385_n140# 0.02fF
C21 w_n1311_n241# a_1039_n140# 0.01fF
C22 a_149_n140# a_861_n140# 0.01fF
C23 a_207_n205# a_n1039_n205# 0.01fF
C24 a_n1275_n140# a_149_n140# 0.01fF
C25 a_29_n205# a_1097_n205# 0.01fF
C26 a_n1097_n140# a_327_n140# 0.01fF
C27 a_1097_n205# a_n327_n205# 0.00fF
C28 a_919_n205# a_n149_n205# 0.01fF
C29 a_327_n140# a_683_n140# 0.03fF
C30 a_n1097_n140# a_n563_n140# 0.02fF
C31 a_1097_n205# a_n385_n140# 0.01fF
C32 a_741_n205# a_n861_n205# 0.01fF
C33 a_1097_n205# a_1039_n140# 0.06fF
C34 a_n563_n140# a_683_n140# 0.01fF
C35 a_n505_n205# a_n861_n205# 0.03fF
C36 a_n1039_n205# a_563_n205# 0.01fF
C37 a_207_n205# a_385_n205# 0.10fF
C38 w_n1311_n241# a_n1039_n205# 0.20fF
C39 a_149_n140# a_n385_n140# 0.02fF
C40 a_327_n140# a_861_n140# 0.02fF
C41 a_149_n140# a_1039_n140# 0.01fF
C42 a_n1275_n140# a_327_n140# 0.01fF
C43 a_n861_n205# a_n149_n205# 0.01fF
C44 a_861_n140# a_n563_n140# 0.01fF
C45 a_n1275_n140# a_n563_n140# 0.01fF
C46 a_385_n205# a_563_n205# 0.10fF
C47 w_n1311_n241# a_385_n205# 0.17fF
C48 a_n919_n140# a_505_n140# 0.01fF
C49 a_n919_n140# a_n29_n140# 0.01fF
C50 a_n741_n140# a_n207_n140# 0.02fF
C51 a_207_n205# a_563_n205# 0.03fF
C52 a_327_n140# a_n385_n140# 0.01fF
C53 a_327_n140# a_1039_n140# 0.01fF
C54 a_207_n205# w_n1311_n241# 0.18fF
C55 a_n563_n140# a_n385_n140# 0.06fF
C56 a_1039_n140# a_n563_n140# 0.01fF
C57 a_1097_n205# a_385_n205# 0.01fF
C58 w_n1311_n241# a_n207_n140# 0.02fF
C59 a_n741_n140# w_n1311_n241# 0.02fF
C60 a_207_n205# a_1097_n205# 0.01fF
C61 a_n29_n140# a_505_n140# 0.02fF
C62 a_n505_n205# a_n1275_n140# 0.01fF
C63 a_n683_n205# a_741_n205# 0.01fF
C64 w_n1311_n241# a_563_n205# 0.16fF
C65 a_1097_n205# a_n207_n140# 0.01fF
C66 a_n919_n140# a_n1097_n140# 0.06fF
C67 a_n919_n140# a_683_n140# 0.01fF
C68 a_n683_n205# a_n505_n205# 0.10fF
C69 a_29_n205# a_741_n205# 0.01fF
C70 a_n1275_n140# a_n149_n205# 0.01fF
C71 a_741_n205# a_n327_n205# 0.01fF
C72 a_1097_n205# a_563_n205# 0.01fF
C73 w_n1311_n241# a_1097_n205# 0.28fF
C74 a_149_n140# a_n207_n140# 0.03fF
C75 a_n741_n140# a_149_n140# 0.01fF
C76 a_29_n205# a_n505_n205# 0.02fF
C77 a_n683_n205# a_n149_n205# 0.02fF
C78 a_n505_n205# a_n327_n205# 0.10fF
C79 a_n1097_n140# a_505_n140# 0.01fF
C80 a_n1097_n140# a_n29_n140# 0.01fF
C81 a_505_n140# a_683_n140# 0.06fF
C82 a_n29_n140# a_683_n140# 0.01fF
C83 a_n919_n140# a_n1275_n140# 0.03fF
C84 a_n683_n205# a_919_n205# 0.01fF
C85 a_29_n205# a_n149_n205# 0.10fF
C86 a_n327_n205# a_n149_n205# 0.10fF
C87 w_n1311_n241# a_149_n140# 0.02fF
C88 a_29_n205# a_919_n205# 0.01fF
C89 a_919_n205# a_n327_n205# 0.01fF
C90 a_n1275_n140# a_n861_n205# 0.02fF
C91 a_1097_n205# a_149_n140# 0.01fF
C92 a_861_n140# a_505_n140# 0.03fF
C93 a_861_n140# a_n29_n140# 0.01fF
C94 a_327_n140# a_n207_n140# 0.02fF
C95 a_n741_n140# a_327_n140# 0.01fF
C96 a_n1275_n140# a_n29_n140# 0.01fF
C97 a_n207_n140# a_n563_n140# 0.03fF
C98 a_n919_n140# a_n385_n140# 0.02fF
C99 a_n741_n140# a_n563_n140# 0.06fF
C100 a_n505_n205# a_n1039_n205# 0.02fF
C101 a_n683_n205# a_n861_n205# 0.10fF
C102 w_n1311_n241# a_327_n140# 0.02fF
C103 a_29_n205# a_n861_n205# 0.01fF
C104 a_n861_n205# a_n327_n205# 0.02fF
C105 a_n1039_n205# a_n149_n205# 0.01fF
C106 w_n1311_n241# a_n563_n140# 0.02fF
C107 a_741_n205# a_385_n205# 0.03fF
C108 a_n385_n140# a_505_n140# 0.01fF
C109 a_n29_n140# a_n385_n140# 0.03fF
C110 a_1097_n205# a_327_n140# 0.01fF
C111 a_1039_n140# a_n29_n140# 0.01fF
C112 a_1039_n140# a_505_n140# 0.02fF
C113 a_861_n140# a_683_n140# 0.06fF
C114 a_n1097_n140# a_n1275_n140# 0.06fF
C115 a_207_n205# a_741_n205# 0.02fF
C116 a_n505_n205# a_385_n205# 0.01fF
C117 a_207_n205# a_n505_n205# 0.01fF
C118 a_385_n205# a_n149_n205# 0.02fF
C119 a_149_n140# a_327_n140# 0.06fF
C120 a_149_n140# a_n563_n140# 0.01fF
C121 a_919_n205# a_385_n205# 0.02fF
C122 a_207_n205# a_n149_n205# 0.03fF
C123 a_741_n205# a_563_n205# 0.10fF
C124 a_n1039_n205# a_n861_n205# 0.10fF
C125 a_n1097_n140# a_n385_n140# 0.01fF
C126 a_741_n205# w_n1311_n241# 0.15fF
C127 a_n385_n140# a_683_n140# 0.01fF
C128 a_1039_n140# a_683_n140# 0.03fF
C129 a_207_n205# a_919_n205# 0.01fF
C130 a_n505_n205# a_563_n205# 0.01fF
C131 a_n505_n205# w_n1311_n241# 0.20fF
C132 a_741_n205# a_1097_n205# 0.02fF
C133 a_n683_n205# a_n1275_n140# 0.01fF
C134 a_563_n205# a_n149_n205# 0.01fF
C135 a_n861_n205# a_385_n205# 0.01fF
C136 w_n1311_n241# a_n149_n205# 0.19fF
C137 a_n505_n205# a_1097_n205# 0.00fF
C138 a_29_n205# a_n1275_n140# 0.00fF
C139 a_861_n140# a_n385_n140# 0.01fF
C140 a_n919_n140# a_n207_n140# 0.01fF
C141 a_n1275_n140# a_n327_n205# 0.01fF
C142 a_n919_n140# a_n741_n140# 0.06fF
C143 a_861_n140# a_1039_n140# 0.06fF
C144 a_327_n140# a_n563_n140# 0.01fF
C145 a_919_n205# a_563_n205# 0.03fF
C146 a_n1275_n140# a_n385_n140# 0.01fF
C147 a_207_n205# a_n861_n205# 0.01fF
C148 a_919_n205# w_n1311_n241# 0.14fF
C149 a_1097_n205# a_n149_n205# 0.00fF
C150 a_29_n205# a_n683_n205# 0.01fF
C151 a_n683_n205# a_n327_n205# 0.03fF
C152 a_n919_n140# w_n1311_n241# 0.02fF
C153 a_919_n205# a_1097_n205# 0.07fF
C154 a_29_n205# a_n327_n205# 0.03fF
C155 a_n207_n140# a_505_n140# 0.01fF
C156 a_n207_n140# a_n29_n140# 0.06fF
C157 a_n741_n140# a_505_n140# 0.01fF
C158 a_n741_n140# a_n29_n140# 0.01fF
C159 a_n861_n205# a_563_n205# 0.01fF
C160 a_1039_n140# a_n385_n140# 0.01fF
C161 w_n1311_n241# a_n861_n205# 0.20fF
C162 a_n1275_n140# a_n1039_n205# 0.07fF
C163 w_n1311_n241# a_n29_n140# 0.02fF
C164 w_n1311_n241# a_505_n140# 0.02fF
C165 a_n683_n205# a_n1039_n205# 0.03fF
C166 a_n919_n140# a_149_n140# 0.01fF
C167 a_1097_n205# a_505_n140# 0.01fF
C168 a_n1097_n140# a_n207_n140# 0.01fF
C169 a_1097_n205# a_n29_n140# 0.01fF
C170 a_n741_n140# a_n1097_n140# 0.03fF
C171 a_n207_n140# a_683_n140# 0.01fF
C172 a_n741_n140# a_683_n140# 0.01fF
C173 a_29_n205# a_n1039_n205# 0.01fF
C174 a_n1039_n205# a_n327_n205# 0.01fF
C175 a_n1275_n140# a_385_n205# 0.00fF
C176 w_n1311_n241# a_n1097_n140# 0.02fF
C177 a_207_n205# a_n1275_n140# 0.00fF
C178 w_n1311_n241# a_683_n140# 0.02fF
C179 a_149_n140# a_505_n140# 0.03fF
C180 a_149_n140# a_n29_n140# 0.06fF
C181 a_n683_n205# a_385_n205# 0.01fF
C182 a_861_n140# a_n207_n140# 0.01fF
C183 a_n741_n140# a_861_n140# 0.01fF
C184 a_n919_n140# a_327_n140# 0.01fF
C185 a_n1275_n140# a_n207_n140# 0.01fF
C186 a_207_n205# a_n683_n205# 0.01fF
C187 a_n741_n140# a_n1275_n140# 0.02fF
C188 a_1097_n205# a_683_n140# 0.02fF
C189 a_n919_n140# a_n563_n140# 0.03fF
C190 a_29_n205# a_385_n205# 0.03fF
C191 a_385_n205# a_n327_n205# 0.01fF
C192 a_n505_n205# a_741_n205# 0.01fF
C193 a_29_n205# a_207_n205# 0.10fF
C194 a_207_n205# a_n327_n205# 0.02fF
C195 w_n1311_n241# a_861_n140# 0.01fF
C196 w_n1311_n241# a_n1275_n140# 0.33fF
C197 a_n1097_n140# a_149_n140# 0.01fF
C198 w_n1311_n241# VSUBS 3.79fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AKSJZW a_n149_n195# a_n207_n140# a_207_n195# a_327_n140#
+ a_n1275_n140# a_n861_n195# a_n29_n140# a_149_n140# a_n1097_n140# a_n1039_n195# a_29_n195#
+ a_n683_n195# a_n741_n140# a_741_n195# a_861_n140# a_1097_n195# a_n563_n140# a_n505_n195#
+ a_563_n195# a_683_n140# a_n919_n140# a_919_n195# a_1039_n140# a_n385_n140# a_n327_n195#
+ a_385_n195# a_505_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n195# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n195# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n195# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n195# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_327_n140# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_861_n140# a_741_n195# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n207_n140# a_n327_n195# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_1097_n195# a_1097_n195# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n195# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1275_n140# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n195# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n195# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n861_n195# a_207_n195# 0.01fF
C1 a_n683_n195# a_n1275_n140# 0.01fF
C2 a_385_n195# a_741_n195# 0.03fF
C3 a_149_n140# a_n385_n140# 0.02fF
C4 a_1097_n195# a_n327_n195# 0.00fF
C5 a_1097_n195# a_683_n140# 0.02fF
C6 a_505_n140# a_683_n140# 0.06fF
C7 a_1097_n195# a_919_n195# 0.06fF
C8 a_n919_n140# a_n1097_n140# 0.06fF
C9 a_741_n195# a_207_n195# 0.02fF
C10 a_563_n195# a_29_n195# 0.02fF
C11 a_683_n140# a_n385_n140# 0.01fF
C12 a_385_n195# a_n327_n195# 0.01fF
C13 a_n505_n195# a_n149_n195# 0.03fF
C14 a_385_n195# a_919_n195# 0.02fF
C15 a_n919_n140# a_n1275_n140# 0.03fF
C16 a_n327_n195# a_207_n195# 0.02fF
C17 a_149_n140# a_861_n140# 0.01fF
C18 a_563_n195# a_n861_n195# 0.01fF
C19 a_919_n195# a_207_n195# 0.01fF
C20 a_385_n195# a_n1039_n195# 0.01fF
C21 a_1097_n195# a_327_n140# 0.01fF
C22 a_n149_n195# a_n1275_n140# 0.01fF
C23 a_149_n140# a_n741_n140# 0.01fF
C24 a_505_n140# a_327_n140# 0.06fF
C25 a_n29_n140# a_149_n140# 0.06fF
C26 a_1097_n195# a_n207_n140# 0.01fF
C27 a_n207_n140# a_505_n140# 0.01fF
C28 a_861_n140# a_683_n140# 0.06fF
C29 a_n1039_n195# a_207_n195# 0.01fF
C30 a_741_n195# a_563_n195# 0.10fF
C31 a_n741_n140# a_683_n140# 0.01fF
C32 a_327_n140# a_n385_n140# 0.01fF
C33 a_n29_n140# a_683_n140# 0.01fF
C34 a_n207_n140# a_n385_n140# 0.06fF
C35 a_n861_n195# a_29_n195# 0.01fF
C36 a_n327_n195# a_563_n195# 0.01fF
C37 a_149_n140# a_n563_n140# 0.01fF
C38 a_919_n195# a_563_n195# 0.03fF
C39 a_385_n195# a_n683_n195# 0.01fF
C40 a_741_n195# a_29_n195# 0.01fF
C41 a_n563_n140# a_683_n140# 0.01fF
C42 a_n505_n195# a_n1275_n140# 0.01fF
C43 a_327_n140# a_861_n140# 0.02fF
C44 a_n1039_n195# a_563_n195# 0.01fF
C45 a_n683_n195# a_207_n195# 0.01fF
C46 a_n919_n140# a_505_n140# 0.01fF
C47 a_n207_n140# a_861_n140# 0.01fF
C48 a_327_n140# a_n741_n140# 0.01fF
C49 a_n327_n195# a_29_n195# 0.03fF
C50 a_n29_n140# a_327_n140# 0.03fF
C51 a_n207_n140# a_n741_n140# 0.02fF
C52 a_n1275_n140# a_n1097_n140# 0.06fF
C53 a_n29_n140# a_n207_n140# 0.06fF
C54 a_n919_n140# a_n385_n140# 0.02fF
C55 a_741_n195# a_n861_n195# 0.01fF
C56 a_1097_n195# a_n149_n195# 0.00fF
C57 a_919_n195# a_29_n195# 0.01fF
C58 a_385_n195# a_n149_n195# 0.02fF
C59 a_n327_n195# a_n861_n195# 0.02fF
C60 a_n1039_n195# a_29_n195# 0.01fF
C61 a_327_n140# a_n563_n140# 0.01fF
C62 a_1097_n195# a_1039_n140# 0.06fF
C63 a_1039_n140# a_505_n140# 0.02fF
C64 a_n207_n140# a_n563_n140# 0.03fF
C65 a_563_n195# a_n683_n195# 0.01fF
C66 a_n149_n195# a_207_n195# 0.03fF
C67 a_741_n195# a_n327_n195# 0.01fF
C68 a_1039_n140# a_n385_n140# 0.01fF
C69 a_149_n140# a_683_n140# 0.02fF
C70 a_n1039_n195# a_n861_n195# 0.10fF
C71 a_n919_n140# a_n741_n140# 0.06fF
C72 a_741_n195# a_919_n195# 0.10fF
C73 a_n29_n140# a_n919_n140# 0.01fF
C74 a_1097_n195# a_n505_n195# 0.00fF
C75 a_29_n195# a_n683_n195# 0.01fF
C76 a_n327_n195# a_919_n195# 0.01fF
C77 a_505_n140# a_n1097_n140# 0.01fF
C78 a_385_n195# a_n505_n195# 0.01fF
C79 a_n149_n195# a_563_n195# 0.01fF
C80 a_1039_n140# a_861_n140# 0.06fF
C81 a_n327_n195# a_n1039_n195# 0.01fF
C82 a_n919_n140# a_n563_n140# 0.03fF
C83 a_n385_n140# a_n1097_n140# 0.01fF
C84 a_149_n140# a_327_n140# 0.06fF
C85 a_n505_n195# a_207_n195# 0.01fF
C86 a_n861_n195# a_n683_n195# 0.10fF
C87 a_n29_n140# a_1039_n140# 0.01fF
C88 a_149_n140# a_n207_n140# 0.03fF
C89 a_n385_n140# a_n1275_n140# 0.01fF
C90 a_385_n195# a_n1275_n140# 0.00fF
C91 a_327_n140# a_683_n140# 0.03fF
C92 a_n207_n140# a_683_n140# 0.01fF
C93 a_741_n195# a_n683_n195# 0.01fF
C94 a_n149_n195# a_29_n195# 0.10fF
C95 a_207_n195# a_n1275_n140# 0.00fF
C96 a_1039_n140# a_n563_n140# 0.01fF
C97 a_n327_n195# a_n683_n195# 0.03fF
C98 a_n741_n140# a_n1097_n140# 0.03fF
C99 a_n505_n195# a_563_n195# 0.01fF
C100 a_n29_n140# a_n1097_n140# 0.01fF
C101 a_919_n195# a_n683_n195# 0.01fF
C102 a_n149_n195# a_n861_n195# 0.01fF
C103 a_149_n140# a_n919_n140# 0.01fF
C104 a_n741_n140# a_n1275_n140# 0.02fF
C105 a_n29_n140# a_n1275_n140# 0.01fF
C106 a_n1039_n195# a_n683_n195# 0.03fF
C107 a_n207_n140# a_327_n140# 0.02fF
C108 a_n149_n195# a_741_n195# 0.01fF
C109 a_1097_n195# a_505_n140# 0.01fF
C110 a_n919_n140# a_683_n140# 0.01fF
C111 a_n563_n140# a_n1097_n140# 0.02fF
C112 a_n505_n195# a_29_n195# 0.02fF
C113 a_385_n195# a_1097_n195# 0.01fF
C114 a_1097_n195# a_n385_n140# 0.01fF
C115 a_505_n140# a_n385_n140# 0.01fF
C116 a_n149_n195# a_n327_n195# 0.10fF
C117 a_n563_n140# a_n1275_n140# 0.01fF
C118 a_149_n140# a_1039_n140# 0.01fF
C119 a_n149_n195# a_919_n195# 0.01fF
C120 a_1097_n195# a_207_n195# 0.01fF
C121 a_n505_n195# a_n861_n195# 0.03fF
C122 a_29_n195# a_n1275_n140# 0.00fF
C123 a_1039_n140# a_683_n140# 0.03fF
C124 a_n149_n195# a_n1039_n195# 0.01fF
C125 a_n919_n140# a_327_n140# 0.01fF
C126 a_385_n195# a_207_n195# 0.10fF
C127 a_n207_n140# a_n919_n140# 0.01fF
C128 a_n505_n195# a_741_n195# 0.01fF
C129 a_1097_n195# a_861_n140# 0.03fF
C130 a_505_n140# a_861_n140# 0.03fF
C131 a_n861_n195# a_n1275_n140# 0.02fF
C132 a_505_n140# a_n741_n140# 0.01fF
C133 a_n29_n140# a_1097_n195# 0.01fF
C134 a_n29_n140# a_505_n140# 0.02fF
C135 a_149_n140# a_n1097_n140# 0.01fF
C136 a_861_n140# a_n385_n140# 0.01fF
C137 a_n505_n195# a_n327_n195# 0.10fF
C138 a_n741_n140# a_n385_n140# 0.03fF
C139 a_1097_n195# a_563_n195# 0.01fF
C140 a_n505_n195# a_919_n195# 0.01fF
C141 a_n29_n140# a_n385_n140# 0.03fF
C142 a_149_n140# a_n1275_n140# 0.01fF
C143 a_1039_n140# a_327_n140# 0.01fF
C144 a_n149_n195# a_n683_n195# 0.02fF
C145 a_n207_n140# a_1039_n140# 0.01fF
C146 a_385_n195# a_563_n195# 0.10fF
C147 a_n505_n195# a_n1039_n195# 0.02fF
C148 a_505_n140# a_n563_n140# 0.01fF
C149 a_n327_n195# a_n1275_n140# 0.01fF
C150 a_563_n195# a_207_n195# 0.03fF
C151 a_n563_n140# a_n385_n140# 0.06fF
C152 a_1097_n195# a_29_n195# 0.01fF
C153 a_n741_n140# a_861_n140# 0.01fF
C154 a_n29_n140# a_861_n140# 0.01fF
C155 a_n1039_n195# a_n1275_n140# 0.06fF
C156 a_n29_n140# a_n741_n140# 0.01fF
C157 a_385_n195# a_29_n195# 0.03fF
C158 a_327_n140# a_n1097_n140# 0.01fF
C159 a_n207_n140# a_n1097_n140# 0.01fF
C160 a_n505_n195# a_n683_n195# 0.10fF
C161 a_29_n195# a_207_n195# 0.10fF
C162 a_327_n140# a_n1275_n140# 0.01fF
C163 a_861_n140# a_n563_n140# 0.01fF
C164 a_n207_n140# a_n1275_n140# 0.01fF
C165 a_385_n195# a_n861_n195# 0.01fF
C166 a_n741_n140# a_n563_n140# 0.06fF
C167 a_1097_n195# a_741_n195# 0.02fF
C168 a_149_n140# a_1097_n195# 0.01fF
C169 a_149_n140# a_505_n140# 0.03fF
C170 a_n29_n140# a_n563_n140# 0.02fF
C171 a_1039_n140# VSUBS 0.01fF
C172 a_861_n140# VSUBS 0.01fF
C173 a_683_n140# VSUBS 0.02fF
C174 a_505_n140# VSUBS 0.02fF
C175 a_327_n140# VSUBS 0.02fF
C176 a_149_n140# VSUBS 0.02fF
C177 a_n29_n140# VSUBS 0.02fF
C178 a_n207_n140# VSUBS 0.02fF
C179 a_n385_n140# VSUBS 0.02fF
C180 a_n563_n140# VSUBS 0.02fF
C181 a_n741_n140# VSUBS 0.02fF
C182 a_n919_n140# VSUBS 0.02fF
C183 a_n1097_n140# VSUBS 0.02fF
C184 a_1097_n195# VSUBS 0.31fF
C185 a_919_n195# VSUBS 0.19fF
C186 a_741_n195# VSUBS 0.20fF
C187 a_563_n195# VSUBS 0.21fF
C188 a_385_n195# VSUBS 0.22fF
C189 a_207_n195# VSUBS 0.23fF
C190 a_29_n195# VSUBS 0.23fF
C191 a_n149_n195# VSUBS 0.24fF
C192 a_n327_n195# VSUBS 0.24fF
C193 a_n505_n195# VSUBS 0.24fF
C194 a_n683_n195# VSUBS 0.24fF
C195 a_n861_n195# VSUBS 0.24fF
C196 a_n1039_n195# VSUBS 0.24fF
C197 a_n1275_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_K7HVMB a_664_n120# a_n608_n120# a_n86_n120# a_72_n208#
+ a_240_n120# a_n184_n120# a_n562_142# a_n510_n120# a_28_n120# a_n298_n120# a_126_n120#
+ a_452_n120# a_n396_n120# a_284_142# a_n138_142# a_550_n120# a_496_n208# a_338_n120#
+ a_n350_n208# a_n820_n120# VSUBS
X0 a_n820_n120# a_n820_n120# a_n820_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X1 a_n510_n120# a_n562_142# a_n608_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X2 a_664_n120# a_664_n120# a_664_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X3 a_n298_n120# a_n350_n208# a_n396_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X4 a_550_n120# a_496_n208# a_452_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X5 a_126_n120# a_72_n208# a_28_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X6 a_n86_n120# a_n138_142# a_n184_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X7 a_338_n120# a_284_142# a_240_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
C0 a_452_n120# a_n184_n120# 0.01fF
C1 a_n298_n120# a_n510_n120# 0.04fF
C2 a_n820_n120# a_n86_n120# 0.02fF
C3 a_72_n208# a_664_n120# 0.00fF
C4 a_n396_n120# a_n86_n120# 0.03fF
C5 a_n510_n120# a_n184_n120# 0.02fF
C6 a_n298_n120# a_126_n120# 0.02fF
C7 a_240_n120# a_28_n120# 0.04fF
C8 a_n298_n120# a_n608_n120# 0.03fF
C9 a_n820_n120# a_452_n120# 0.01fF
C10 a_28_n120# a_664_n120# 0.02fF
C11 a_126_n120# a_n184_n120# 0.03fF
C12 a_n396_n120# a_452_n120# 0.01fF
C13 a_n608_n120# a_n184_n120# 0.02fF
C14 a_n298_n120# a_550_n120# 0.01fF
C15 a_496_n208# a_n562_142# 0.00fF
C16 a_n820_n120# a_n510_n120# 0.06fF
C17 a_550_n120# a_n184_n120# 0.01fF
C18 a_n510_n120# a_n396_n120# 0.09fF
C19 a_n562_142# a_n138_142# 0.01fF
C20 a_n820_n120# a_126_n120# 0.02fF
C21 a_452_n120# a_n86_n120# 0.01fF
C22 a_n820_n120# a_n608_n120# 0.13fF
C23 a_126_n120# a_n396_n120# 0.01fF
C24 a_240_n120# a_664_n120# 0.03fF
C25 a_n608_n120# a_n396_n120# 0.04fF
C26 a_n298_n120# a_338_n120# 0.01fF
C27 a_n820_n120# a_550_n120# 0.01fF
C28 a_n510_n120# a_n86_n120# 0.02fF
C29 a_338_n120# a_n184_n120# 0.01fF
C30 a_550_n120# a_n396_n120# 0.01fF
C31 a_496_n208# a_72_n208# 0.01fF
C32 a_n562_142# a_284_142# 0.01fF
C33 a_126_n120# a_n86_n120# 0.04fF
C34 a_n820_n120# a_n562_142# 0.01fF
C35 a_72_n208# a_n138_142# 0.01fF
C36 a_n510_n120# a_452_n120# 0.01fF
C37 a_n608_n120# a_n86_n120# 0.01fF
C38 a_n298_n120# a_28_n120# 0.02fF
C39 a_126_n120# a_452_n120# 0.02fF
C40 a_n820_n120# a_338_n120# 0.01fF
C41 a_550_n120# a_n86_n120# 0.01fF
C42 a_n562_142# a_n350_n208# 0.01fF
C43 a_n608_n120# a_452_n120# 0.01fF
C44 a_n396_n120# a_338_n120# 0.01fF
C45 a_28_n120# a_n184_n120# 0.04fF
C46 a_n510_n120# a_126_n120# 0.01fF
C47 a_550_n120# a_452_n120# 0.11fF
C48 a_72_n208# a_284_142# 0.01fF
C49 a_n510_n120# a_n608_n120# 0.11fF
C50 a_n820_n120# a_72_n208# 0.00fF
C51 a_n510_n120# a_550_n120# 0.01fF
C52 a_n86_n120# a_338_n120# 0.02fF
C53 a_126_n120# a_n608_n120# 0.01fF
C54 a_n820_n120# a_28_n120# 0.02fF
C55 a_496_n208# a_664_n120# 0.01fF
C56 a_n298_n120# a_240_n120# 0.01fF
C57 a_28_n120# a_n396_n120# 0.02fF
C58 a_72_n208# a_n350_n208# 0.01fF
C59 a_126_n120# a_550_n120# 0.02fF
C60 a_n138_142# a_664_n120# 0.00fF
C61 a_n298_n120# a_664_n120# 0.01fF
C62 a_n510_n120# a_n562_142# 0.00fF
C63 a_240_n120# a_n184_n120# 0.02fF
C64 a_452_n120# a_338_n120# 0.09fF
C65 a_550_n120# a_n608_n120# 0.01fF
C66 a_n184_n120# a_664_n120# 0.02fF
C67 a_n510_n120# a_338_n120# 0.01fF
C68 a_28_n120# a_n86_n120# 0.09fF
C69 a_240_n120# a_284_142# 0.00fF
C70 a_n820_n120# a_240_n120# 0.01fF
C71 a_126_n120# a_338_n120# 0.04fF
C72 a_284_142# a_664_n120# 0.01fF
C73 a_240_n120# a_n396_n120# 0.01fF
C74 a_n820_n120# a_664_n120# 0.02fF
C75 a_n608_n120# a_338_n120# 0.01fF
C76 a_28_n120# a_452_n120# 0.02fF
C77 a_n396_n120# a_664_n120# 0.01fF
C78 a_550_n120# a_338_n120# 0.04fF
C79 a_28_n120# a_n510_n120# 0.01fF
C80 a_n350_n208# a_664_n120# 0.00fF
C81 a_240_n120# a_n86_n120# 0.02fF
C82 a_496_n208# a_n138_142# 0.00fF
C83 a_28_n120# a_126_n120# 0.11fF
C84 a_n86_n120# a_664_n120# 0.02fF
C85 a_28_n120# a_n608_n120# 0.01fF
C86 a_240_n120# a_452_n120# 0.04fF
C87 a_28_n120# a_550_n120# 0.01fF
C88 a_452_n120# a_664_n120# 0.06fF
C89 a_n298_n120# a_n184_n120# 0.09fF
C90 a_72_n208# a_n562_142# 0.00fF
C91 a_240_n120# a_n510_n120# 0.01fF
C92 a_496_n208# a_284_142# 0.01fF
C93 a_n820_n120# a_496_n208# 0.00fF
C94 a_n510_n120# a_664_n120# 0.01fF
C95 a_240_n120# a_126_n120# 0.09fF
C96 a_284_142# a_n138_142# 0.01fF
C97 a_240_n120# a_n608_n120# 0.01fF
C98 a_n820_n120# a_n138_142# 0.00fF
C99 a_n820_n120# a_n298_n120# 0.03fF
C100 a_126_n120# a_664_n120# 0.03fF
C101 a_28_n120# a_338_n120# 0.03fF
C102 a_n298_n120# a_n396_n120# 0.11fF
C103 a_n608_n120# a_664_n120# 0.01fF
C104 a_496_n208# a_n350_n208# 0.01fF
C105 a_240_n120# a_550_n120# 0.03fF
C106 a_n820_n120# a_n184_n120# 0.03fF
C107 a_n396_n120# a_n184_n120# 0.04fF
C108 a_550_n120# a_664_n120# 0.13fF
C109 a_n350_n208# a_n138_142# 0.01fF
C110 a_n298_n120# a_n350_n208# 0.00fF
C111 a_28_n120# a_72_n208# 0.00fF
C112 a_n820_n120# a_284_142# 0.00fF
C113 a_n86_n120# a_n138_142# 0.00fF
C114 a_n298_n120# a_n86_n120# 0.04fF
C115 a_n562_142# a_664_n120# 0.00fF
C116 a_496_n208# a_452_n120# 0.00fF
C117 a_240_n120# a_338_n120# 0.11fF
C118 a_n86_n120# a_n184_n120# 0.11fF
C119 a_n820_n120# a_n396_n120# 0.04fF
C120 a_n298_n120# a_452_n120# 0.01fF
C121 a_338_n120# a_664_n120# 0.04fF
C122 a_284_142# a_n350_n208# 0.00fF
C123 a_n820_n120# a_n350_n208# 0.01fF
C124 a_550_n120# VSUBS 0.01fF
C125 a_452_n120# VSUBS 0.01fF
C126 a_338_n120# VSUBS 0.01fF
C127 a_240_n120# VSUBS 0.01fF
C128 a_126_n120# VSUBS 0.02fF
C129 a_28_n120# VSUBS 0.01fF
C130 a_n86_n120# VSUBS 0.01fF
C131 a_n184_n120# VSUBS 0.02fF
C132 a_n298_n120# VSUBS 0.02fF
C133 a_n396_n120# VSUBS 0.02fF
C134 a_n510_n120# VSUBS 0.02fF
C135 a_n608_n120# VSUBS 0.02fF
C136 a_496_n208# VSUBS 0.11fF
C137 a_664_n120# VSUBS 0.17fF
C138 a_72_n208# VSUBS 0.10fF
C139 a_284_142# VSUBS 0.10fF
C140 a_n350_n208# VSUBS 0.12fF
C141 a_n138_142# VSUBS 0.11fF
C142 a_n820_n120# VSUBS 0.20fF
C143 a_n562_142# VSUBS 0.14fF
.ends

.subckt sky130_fd_pr__nfet_01v8_S6RQQZ a_n149_n194# a_n207_n140# a_207_n194# a_1453_n194#
+ a_n1217_n194# a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140#
+ a_n1097_n140# a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194#
+ a_861_n140# a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140#
+ a_n919_n140# a_919_n194# a_n1631_n140# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194#
+ a_n1395_n194# a_505_n140# a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n1453_n140# a_n1631_n140# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1453_n194# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1217_n194# a_n149_n194# 0.01fF
C1 a_n683_n194# a_n1631_n140# 0.01fF
C2 a_n1631_n140# a_n919_n140# 0.01fF
C3 a_1275_n194# a_n327_n194# 0.01fF
C4 a_207_n194# a_1453_n194# 0.00fF
C5 a_1395_n140# a_505_n140# 0.01fF
C6 a_29_n194# a_385_n194# 0.03fF
C7 a_741_n194# a_n683_n194# 0.01fF
C8 a_n385_n140# a_n1453_n140# 0.01fF
C9 a_683_n140# a_1039_n140# 0.03fF
C10 a_n563_n140# a_n919_n140# 0.03fF
C11 a_683_n140# a_149_n140# 0.02fF
C12 a_861_n140# a_505_n140# 0.03fF
C13 a_741_n194# a_563_n194# 0.10fF
C14 a_n207_n140# a_n29_n140# 0.06fF
C15 a_1097_n194# a_919_n194# 0.10fF
C16 a_385_n194# a_n149_n194# 0.02fF
C17 a_207_n194# a_n327_n194# 0.02fF
C18 a_29_n194# a_n683_n194# 0.01fF
C19 a_n919_n140# a_n1453_n140# 0.02fF
C20 a_n861_n194# a_n505_n194# 0.03fF
C21 a_n1395_n194# a_n1631_n140# 0.06fF
C22 a_505_n140# a_1217_n140# 0.01fF
C23 a_n385_n140# a_861_n140# 0.01fF
C24 a_29_n194# a_563_n194# 0.02fF
C25 a_n505_n194# a_919_n194# 0.01fF
C26 a_n683_n194# a_n149_n194# 0.02fF
C27 a_n385_n140# a_1217_n140# 0.01fF
C28 a_207_n194# a_n1217_n194# 0.01fF
C29 a_29_n194# a_n1395_n194# 0.01fF
C30 a_563_n194# a_n149_n194# 0.01fF
C31 a_327_n140# a_1039_n140# 0.01fF
C32 a_n1631_n140# a_n1097_n140# 0.02fF
C33 a_385_n194# a_1275_n194# 0.01fF
C34 a_149_n140# a_327_n140# 0.06fF
C35 a_n563_n140# a_n1097_n140# 0.02fF
C36 a_n741_n140# a_n1631_n140# 0.01fF
C37 a_n1275_n140# a_n385_n140# 0.01fF
C38 a_n741_n140# a_n563_n140# 0.06fF
C39 a_n1395_n194# a_n149_n194# 0.01fF
C40 a_385_n194# a_207_n194# 0.10fF
C41 a_n1097_n140# a_n1453_n140# 0.03fF
C42 a_505_n140# a_1453_n194# 0.01fF
C43 a_683_n140# a_n563_n140# 0.01fF
C44 a_n1275_n140# a_n919_n140# 0.03fF
C45 a_n741_n140# a_n1453_n140# 0.01fF
C46 a_n1631_n140# a_n1039_n194# 0.01fF
C47 a_563_n194# a_1275_n194# 0.01fF
C48 a_n1217_n194# a_n327_n194# 0.01fF
C49 a_n683_n194# a_207_n194# 0.01fF
C50 a_385_n194# a_1453_n194# 0.01fF
C51 a_n207_n140# a_1039_n140# 0.01fF
C52 a_n207_n140# a_149_n140# 0.03fF
C53 a_1039_n140# a_n29_n140# 0.01fF
C54 a_149_n140# a_n29_n140# 0.06fF
C55 a_563_n194# a_207_n194# 0.03fF
C56 a_29_n194# a_n1039_n194# 0.01fF
C57 a_n741_n140# a_861_n140# 0.01fF
C58 a_1395_n140# a_683_n140# 0.01fF
C59 a_385_n194# a_n327_n194# 0.01fF
C60 a_861_n140# a_683_n140# 0.06fF
C61 a_n1039_n194# a_n149_n194# 0.01fF
C62 a_n1395_n194# a_207_n194# 0.01fF
C63 a_741_n194# a_1097_n194# 0.03fF
C64 a_563_n194# a_1453_n194# 0.01fF
C65 a_n563_n140# a_327_n140# 0.01fF
C66 a_n683_n194# a_n327_n194# 0.03fF
C67 a_n1275_n140# a_n1097_n140# 0.06fF
C68 a_n505_n194# a_n1631_n140# 0.01fF
C69 a_n1275_n140# a_n741_n140# 0.02fF
C70 a_683_n140# a_1217_n140# 0.02fF
C71 a_741_n194# a_n505_n194# 0.01fF
C72 a_385_n194# a_n1217_n194# 0.01fF
C73 a_29_n194# a_1097_n194# 0.01fF
C74 a_563_n194# a_n327_n194# 0.01fF
C75 a_n385_n140# a_505_n140# 0.01fF
C76 a_1097_n194# a_n149_n194# 0.01fF
C77 a_29_n194# a_n505_n194# 0.02fF
C78 a_1395_n140# a_327_n140# 0.01fF
C79 a_n683_n194# a_n1217_n194# 0.02fF
C80 a_n1395_n194# a_n327_n194# 0.01fF
C81 a_n207_n140# a_n1631_n140# 0.01fF
C82 a_505_n140# a_n919_n140# 0.01fF
C83 a_n1631_n140# a_n29_n140# 0.01fF
C84 a_n207_n140# a_n563_n140# 0.03fF
C85 a_861_n140# a_327_n140# 0.02fF
C86 a_n563_n140# a_n29_n140# 0.02fF
C87 a_207_n194# a_n1039_n194# 0.01fF
C88 a_n505_n194# a_n149_n194# 0.03fF
C89 a_149_n140# a_1039_n140# 0.01fF
C90 a_385_n194# a_n683_n194# 0.01fF
C91 a_683_n140# a_1453_n194# 0.01fF
C92 a_n207_n140# a_n1453_n140# 0.01fF
C93 a_n385_n140# a_n919_n140# 0.02fF
C94 a_327_n140# a_1217_n140# 0.01fF
C95 a_n1453_n140# a_n29_n140# 0.01fF
C96 a_n1395_n194# a_n1217_n194# 0.10fF
C97 a_1097_n194# a_1275_n194# 0.10fF
C98 a_385_n194# a_563_n194# 0.10fF
C99 a_n861_n194# a_n1631_n140# 0.01fF
C100 a_n1275_n140# a_327_n140# 0.01fF
C101 a_1395_n140# a_n207_n140# 0.01fF
C102 a_741_n194# a_n861_n194# 0.01fF
C103 a_1395_n140# a_n29_n140# 0.01fF
C104 a_1097_n194# a_207_n194# 0.01fF
C105 a_861_n140# a_n207_n140# 0.01fF
C106 a_n327_n194# a_n1039_n194# 0.01fF
C107 a_n683_n194# a_563_n194# 0.01fF
C108 a_861_n140# a_n29_n140# 0.01fF
C109 a_741_n194# a_919_n194# 0.10fF
C110 a_505_n140# a_n1097_n140# 0.01fF
C111 a_29_n194# a_n861_n194# 0.01fF
C112 a_n741_n140# a_505_n140# 0.01fF
C113 a_n207_n140# a_1217_n140# 0.01fF
C114 a_n505_n194# a_207_n194# 0.01fF
C115 a_n683_n194# a_n1395_n194# 0.01fF
C116 a_1097_n194# a_1453_n194# 0.02fF
C117 a_1217_n140# a_n29_n140# 0.01fF
C118 a_327_n140# a_1453_n194# 0.01fF
C119 a_29_n194# a_919_n194# 0.01fF
C120 a_n385_n140# a_n1097_n140# 0.01fF
C121 a_683_n140# a_505_n140# 0.06fF
C122 a_n861_n194# a_n149_n194# 0.01fF
C123 a_n1217_n194# a_n1039_n194# 0.10fF
C124 a_n1275_n140# a_n207_n140# 0.01fF
C125 a_n385_n140# a_n741_n140# 0.03fF
C126 a_n1275_n140# a_n29_n140# 0.01fF
C127 a_1097_n194# a_n327_n194# 0.01fF
C128 a_n563_n140# a_1039_n140# 0.01fF
C129 a_n563_n140# a_149_n140# 0.01fF
C130 a_n149_n194# a_919_n194# 0.01fF
C131 a_n1097_n140# a_n919_n140# 0.06fF
C132 a_n385_n140# a_683_n140# 0.01fF
C133 a_n741_n140# a_n919_n140# 0.06fF
C134 a_385_n194# a_n1039_n194# 0.01fF
C135 a_n505_n194# a_n327_n194# 0.10fF
C136 a_149_n140# a_n1453_n140# 0.01fF
C137 a_683_n140# a_n919_n140# 0.01fF
C138 a_1453_n194# a_n29_n140# 0.01fF
C139 a_1395_n140# a_1039_n140# 0.03fF
C140 a_n683_n194# a_n1039_n194# 0.03fF
C141 a_505_n140# a_327_n140# 0.06fF
C142 a_1395_n140# a_149_n140# 0.01fF
C143 a_1275_n194# a_919_n194# 0.03fF
C144 a_n861_n194# a_207_n194# 0.01fF
C145 a_861_n140# a_1039_n140# 0.06fF
C146 a_563_n194# a_n1039_n194# 0.01fF
C147 a_861_n140# a_149_n140# 0.01fF
C148 a_n505_n194# a_n1217_n194# 0.01fF
C149 a_1097_n194# a_385_n194# 0.01fF
C150 a_n385_n140# a_327_n140# 0.01fF
C151 a_207_n194# a_919_n194# 0.01fF
C152 a_1217_n140# a_1039_n140# 0.06fF
C153 a_149_n140# a_1217_n140# 0.01fF
C154 a_n1395_n194# a_n1039_n194# 0.03fF
C155 a_n741_n140# a_n1097_n140# 0.03fF
C156 a_n563_n140# a_n1631_n140# 0.01fF
C157 a_n505_n194# a_385_n194# 0.01fF
C158 a_327_n140# a_n919_n140# 0.01fF
C159 a_n1275_n140# a_149_n140# 0.01fF
C160 a_1453_n194# a_919_n194# 0.01fF
C161 a_n207_n140# a_505_n140# 0.01fF
C162 a_n861_n194# a_n327_n194# 0.02fF
C163 a_1097_n194# a_563_n194# 0.02fF
C164 a_n741_n140# a_683_n140# 0.01fF
C165 a_505_n140# a_n29_n140# 0.02fF
C166 a_n1631_n140# a_n1453_n140# 0.06fF
C167 a_29_n194# a_n1631_n140# 0.00fF
C168 a_29_n194# a_741_n194# 0.01fF
C169 a_n563_n140# a_n1453_n140# 0.01fF
C170 a_n505_n194# a_n683_n194# 0.10fF
C171 a_n327_n194# a_919_n194# 0.01fF
C172 a_n385_n140# a_n207_n140# 0.06fF
C173 a_n505_n194# a_563_n194# 0.01fF
C174 a_n385_n140# a_n29_n140# 0.03fF
C175 a_n1631_n140# a_n149_n194# 0.00fF
C176 a_741_n194# a_n149_n194# 0.01fF
C177 a_1453_n194# a_1039_n140# 0.02fF
C178 a_n861_n194# a_n1217_n194# 0.03fF
C179 a_149_n140# a_1453_n194# 0.01fF
C180 a_n207_n140# a_n919_n140# 0.01fF
C181 a_861_n140# a_n563_n140# 0.01fF
C182 a_n505_n194# a_n1395_n194# 0.01fF
C183 a_n919_n140# a_n29_n140# 0.01fF
C184 a_29_n194# a_n149_n194# 0.10fF
C185 a_n1097_n140# a_327_n140# 0.01fF
C186 a_n741_n140# a_327_n140# 0.01fF
C187 a_n861_n194# a_385_n194# 0.01fF
C188 a_741_n194# a_1275_n194# 0.02fF
C189 a_n1275_n140# a_n1631_n140# 0.03fF
C190 a_683_n140# a_327_n140# 0.03fF
C191 a_n1275_n140# a_n563_n140# 0.01fF
C192 a_385_n194# a_919_n194# 0.02fF
C193 a_1395_n140# a_861_n140# 0.02fF
C194 a_n861_n194# a_n683_n194# 0.10fF
C195 a_741_n194# a_207_n194# 0.02fF
C196 a_29_n194# a_1275_n194# 0.01fF
C197 a_505_n140# a_1039_n140# 0.02fF
C198 a_n861_n194# a_563_n194# 0.01fF
C199 a_n1275_n140# a_n1453_n140# 0.06fF
C200 a_505_n140# a_149_n140# 0.03fF
C201 a_n683_n194# a_919_n194# 0.01fF
C202 a_1395_n140# a_1217_n140# 0.06fF
C203 a_n207_n140# a_n1097_n140# 0.01fF
C204 a_n505_n194# a_n1039_n194# 0.02fF
C205 a_n1097_n140# a_n29_n140# 0.01fF
C206 a_n741_n140# a_n207_n140# 0.02fF
C207 a_29_n194# a_207_n194# 0.10fF
C208 a_1275_n194# a_n149_n194# 0.01fF
C209 a_861_n140# a_1217_n140# 0.03fF
C210 a_563_n194# a_919_n194# 0.03fF
C211 a_n741_n140# a_n29_n140# 0.01fF
C212 a_741_n194# a_1453_n194# 0.01fF
C213 a_n385_n140# a_1039_n140# 0.01fF
C214 a_n861_n194# a_n1395_n194# 0.02fF
C215 a_n385_n140# a_149_n140# 0.02fF
C216 a_683_n140# a_n207_n140# 0.01fF
C217 a_683_n140# a_n29_n140# 0.01fF
C218 a_n1631_n140# a_n327_n194# 0.00fF
C219 a_207_n194# a_n149_n194# 0.03fF
C220 a_29_n194# a_1453_n194# 0.00fF
C221 a_741_n194# a_n327_n194# 0.01fF
C222 a_149_n140# a_n919_n140# 0.01fF
C223 a_n505_n194# a_1097_n194# 0.01fF
C224 a_1395_n140# a_1453_n194# 0.06fF
C225 a_1453_n194# a_n149_n194# 0.00fF
C226 a_29_n194# a_n327_n194# 0.03fF
C227 a_n1631_n140# a_n1217_n194# 0.02fF
C228 a_861_n140# a_1453_n194# 0.01fF
C229 a_207_n194# a_1275_n194# 0.01fF
C230 a_n861_n194# a_n1039_n194# 0.10fF
C231 a_n327_n194# a_n149_n194# 0.10fF
C232 a_n563_n140# a_505_n140# 0.01fF
C233 a_n207_n140# a_327_n140# 0.02fF
C234 a_327_n140# a_n29_n140# 0.03fF
C235 a_1217_n140# a_1453_n194# 0.03fF
C236 a_29_n194# a_n1217_n194# 0.01fF
C237 a_n385_n140# a_n1631_n140# 0.01fF
C238 a_1275_n194# a_1453_n194# 0.06fF
C239 a_741_n194# a_385_n194# 0.03fF
C240 a_149_n140# a_n1097_n140# 0.01fF
C241 a_n385_n140# a_n563_n140# 0.06fF
C242 a_n741_n140# a_149_n140# 0.01fF
C243 a_1395_n140# VSUBS 0.01fF
C244 a_1217_n140# VSUBS 0.01fF
C245 a_1039_n140# VSUBS 0.02fF
C246 a_861_n140# VSUBS 0.02fF
C247 a_683_n140# VSUBS 0.02fF
C248 a_505_n140# VSUBS 0.02fF
C249 a_327_n140# VSUBS 0.02fF
C250 a_149_n140# VSUBS 0.02fF
C251 a_n29_n140# VSUBS 0.02fF
C252 a_n207_n140# VSUBS 0.02fF
C253 a_n385_n140# VSUBS 0.02fF
C254 a_n563_n140# VSUBS 0.02fF
C255 a_n741_n140# VSUBS 0.02fF
C256 a_n919_n140# VSUBS 0.02fF
C257 a_n1097_n140# VSUBS 0.02fF
C258 a_n1275_n140# VSUBS 0.02fF
C259 a_n1453_n140# VSUBS 0.02fF
C260 a_1453_n194# VSUBS 0.31fF
C261 a_1275_n194# VSUBS 0.19fF
C262 a_1097_n194# VSUBS 0.20fF
C263 a_919_n194# VSUBS 0.21fF
C264 a_741_n194# VSUBS 0.22fF
C265 a_563_n194# VSUBS 0.23fF
C266 a_385_n194# VSUBS 0.23fF
C267 a_207_n194# VSUBS 0.24fF
C268 a_29_n194# VSUBS 0.24fF
C269 a_n149_n194# VSUBS 0.24fF
C270 a_n327_n194# VSUBS 0.24fF
C271 a_n505_n194# VSUBS 0.24fF
C272 a_n683_n194# VSUBS 0.24fF
C273 a_n861_n194# VSUBS 0.24fF
C274 a_n1039_n194# VSUBS 0.24fF
C275 a_n1217_n194# VSUBS 0.24fF
C276 a_n1395_n194# VSUBS 0.24fF
C277 a_n1631_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_6RUDQZ a_n594_n195# a_n1008_n140# a_n652_n140# a_652_n195#
+ a_772_n140# a_n60_n195# a_n474_n140# a_n416_n195# a_474_n195# a_594_n140# a_n296_n140#
+ a_n238_n195# a_60_n140# a_296_n195# a_416_n140# a_n118_n140# a_118_n195# a_238_n140#
+ a_n772_n195# a_n830_n140# a_830_n195# VSUBS
X0 a_772_n140# a_652_n195# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n195# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n195# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n195# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n195# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_830_n195# a_830_n195# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n1008_n140# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n195# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n195# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n195# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n195# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_772_n140# a_n474_n140# 0.01fF
C1 a_594_n140# a_n652_n140# 0.01fF
C2 a_474_n195# a_652_n195# 0.10fF
C3 a_n772_n195# a_n238_n195# 0.02fF
C4 a_n1008_n140# a_n594_n195# 0.02fF
C5 a_238_n140# a_416_n140# 0.06fF
C6 a_118_n195# a_n60_n195# 0.10fF
C7 a_n118_n140# a_60_n140# 0.06fF
C8 a_n1008_n140# a_594_n140# 0.01fF
C9 a_296_n195# a_n1008_n140# 0.00fF
C10 a_416_n140# a_n652_n140# 0.01fF
C11 a_n1008_n140# a_652_n195# 0.00fF
C12 a_594_n140# a_n296_n140# 0.01fF
C13 a_n238_n195# a_n416_n195# 0.10fF
C14 a_238_n140# a_830_n195# 0.01fF
C15 a_474_n195# a_830_n195# 0.02fF
C16 a_n1008_n140# a_416_n140# 0.01fF
C17 a_n830_n140# a_594_n140# 0.01fF
C18 a_594_n140# a_772_n140# 0.06fF
C19 a_830_n195# a_n652_n140# 0.01fF
C20 a_n772_n195# a_474_n195# 0.01fF
C21 a_416_n140# a_n296_n140# 0.01fF
C22 a_n830_n140# a_416_n140# 0.01fF
C23 a_594_n140# a_n474_n140# 0.01fF
C24 a_118_n195# a_n238_n195# 0.03fF
C25 a_n238_n195# a_n60_n195# 0.10fF
C26 a_416_n140# a_772_n140# 0.03fF
C27 a_n1008_n140# a_n772_n195# 0.06fF
C28 a_238_n140# a_n118_n140# 0.03fF
C29 a_416_n140# a_n474_n140# 0.01fF
C30 a_474_n195# a_n416_n195# 0.01fF
C31 a_830_n195# a_n296_n140# 0.01fF
C32 a_n118_n140# a_n652_n140# 0.02fF
C33 a_772_n140# a_830_n195# 0.06fF
C34 a_296_n195# a_n594_n195# 0.01fF
C35 a_830_n195# a_n474_n140# 0.01fF
C36 a_n594_n195# a_652_n195# 0.01fF
C37 a_n1008_n140# a_n118_n140# 0.01fF
C38 a_118_n195# a_474_n195# 0.03fF
C39 a_n1008_n140# a_n416_n195# 0.01fF
C40 a_474_n195# a_n60_n195# 0.02fF
C41 a_296_n195# a_652_n195# 0.03fF
C42 a_n118_n140# a_n296_n140# 0.06fF
C43 a_594_n140# a_416_n140# 0.06fF
C44 a_n830_n140# a_n118_n140# 0.01fF
C45 a_n118_n140# a_772_n140# 0.01fF
C46 a_n1008_n140# a_118_n195# 0.01fF
C47 a_n1008_n140# a_n60_n195# 0.01fF
C48 a_238_n140# a_60_n140# 0.06fF
C49 a_n594_n195# a_830_n195# 0.00fF
C50 a_n118_n140# a_n474_n140# 0.03fF
C51 a_n652_n140# a_60_n140# 0.01fF
C52 a_594_n140# a_830_n195# 0.03fF
C53 a_n772_n195# a_n594_n195# 0.10fF
C54 a_296_n195# a_830_n195# 0.01fF
C55 a_474_n195# a_n238_n195# 0.01fF
C56 a_830_n195# a_652_n195# 0.06fF
C57 a_296_n195# a_n772_n195# 0.01fF
C58 a_n1008_n140# a_60_n140# 0.01fF
C59 a_416_n140# a_830_n195# 0.02fF
C60 a_n772_n195# a_652_n195# 0.01fF
C61 a_n594_n195# a_n416_n195# 0.10fF
C62 a_n296_n140# a_60_n140# 0.03fF
C63 a_n830_n140# a_60_n140# 0.01fF
C64 a_n1008_n140# a_n238_n195# 0.01fF
C65 a_n118_n140# a_594_n140# 0.01fF
C66 a_296_n195# a_n416_n195# 0.01fF
C67 a_772_n140# a_60_n140# 0.01fF
C68 a_n416_n195# a_652_n195# 0.01fF
C69 a_n772_n195# a_830_n195# 0.00fF
C70 a_n474_n140# a_60_n140# 0.02fF
C71 a_118_n195# a_n594_n195# 0.01fF
C72 a_n118_n140# a_416_n140# 0.02fF
C73 a_n594_n195# a_n60_n195# 0.02fF
C74 a_238_n140# a_n652_n140# 0.01fF
C75 a_296_n195# a_118_n195# 0.10fF
C76 a_296_n195# a_n60_n195# 0.03fF
C77 a_238_n140# a_n1008_n140# 0.01fF
C78 a_118_n195# a_652_n195# 0.02fF
C79 a_n1008_n140# a_474_n195# 0.00fF
C80 a_652_n195# a_n60_n195# 0.01fF
C81 a_n118_n140# a_830_n195# 0.01fF
C82 a_830_n195# a_n416_n195# 0.00fF
C83 a_n1008_n140# a_n652_n140# 0.03fF
C84 a_238_n140# a_n296_n140# 0.02fF
C85 a_n772_n195# a_n416_n195# 0.03fF
C86 a_n830_n140# a_238_n140# 0.01fF
C87 a_594_n140# a_60_n140# 0.02fF
C88 a_n296_n140# a_n652_n140# 0.03fF
C89 a_238_n140# a_772_n140# 0.02fF
C90 a_n830_n140# a_n652_n140# 0.06fF
C91 a_n594_n195# a_n238_n195# 0.03fF
C92 a_118_n195# a_830_n195# 0.01fF
C93 a_830_n195# a_n60_n195# 0.01fF
C94 a_772_n140# a_n652_n140# 0.01fF
C95 a_416_n140# a_60_n140# 0.03fF
C96 a_238_n140# a_n474_n140# 0.01fF
C97 a_296_n195# a_n238_n195# 0.02fF
C98 a_n1008_n140# a_n296_n140# 0.01fF
C99 a_n772_n195# a_118_n195# 0.01fF
C100 a_n830_n140# a_n1008_n140# 0.06fF
C101 a_n772_n195# a_n60_n195# 0.01fF
C102 a_n474_n140# a_n652_n140# 0.06fF
C103 a_n238_n195# a_652_n195# 0.01fF
C104 a_n830_n140# a_n296_n140# 0.02fF
C105 a_830_n195# a_60_n140# 0.01fF
C106 a_n1008_n140# a_n474_n140# 0.02fF
C107 a_772_n140# a_n296_n140# 0.01fF
C108 a_n830_n140# a_772_n140# 0.01fF
C109 a_474_n195# a_n594_n195# 0.01fF
C110 a_118_n195# a_n416_n195# 0.02fF
C111 a_n416_n195# a_n60_n195# 0.03fF
C112 a_n296_n140# a_n474_n140# 0.06fF
C113 a_238_n140# a_594_n140# 0.03fF
C114 a_n238_n195# a_830_n195# 0.01fF
C115 a_296_n195# a_474_n195# 0.10fF
C116 a_n830_n140# a_n474_n140# 0.03fF
C117 a_772_n140# VSUBS 0.01fF
C118 a_594_n140# VSUBS 0.01fF
C119 a_416_n140# VSUBS 0.02fF
C120 a_238_n140# VSUBS 0.02fF
C121 a_60_n140# VSUBS 0.02fF
C122 a_n118_n140# VSUBS 0.02fF
C123 a_n296_n140# VSUBS 0.02fF
C124 a_n474_n140# VSUBS 0.02fF
C125 a_n652_n140# VSUBS 0.02fF
C126 a_n830_n140# VSUBS 0.02fF
C127 a_830_n195# VSUBS 0.31fF
C128 a_652_n195# VSUBS 0.19fF
C129 a_474_n195# VSUBS 0.20fF
C130 a_296_n195# VSUBS 0.21fF
C131 a_118_n195# VSUBS 0.22fF
C132 a_n60_n195# VSUBS 0.23fF
C133 a_n238_n195# VSUBS 0.23fF
C134 a_n416_n195# VSUBS 0.24fF
C135 a_n594_n195# VSUBS 0.24fF
C136 a_n772_n195# VSUBS 0.24fF
C137 a_n1008_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_SD55Q9 a_352_607# a_644_607# a_174_607# a_60_607#
+ a_232_553# a_n232_n389# a_466_607# a_n524_n389# a_524_553# a_n410_n887# a_n702_n887#
+ a_n994_n887# a_644_n389# a_352_n389# a_60_n389# a_524_55# a_n60_55# a_n352_55# a_n232_n887#
+ a_n524_n887# a_174_n389# a_n352_n445# a_466_n389# a_n60_n445# a_n644_n445# a_644_n887#
+ a_352_n887# a_n118_n389# a_60_n887# a_174_n887# a_n352_n943# a_466_n887# a_n118_n887#
+ a_n60_n943# a_n644_n943# a_232_n445# a_n118_109# a_n410_109# a_758_n887# a_524_n445#
+ a_n232_109# a_n702_109# a_n644_55# a_n524_109# a_352_109# a_232_55# a_n352_553#
+ a_644_109# a_174_109# a_60_109# a_n644_553# a_n60_553# a_466_109# a_n410_607# a_524_n943#
+ a_232_n943# a_n410_n389# a_n118_607# a_n702_n389# a_n232_607# a_n702_607# a_n524_607#
+ VSUBS
X0 a_60_n389# a_n60_n445# a_n118_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_644_n887# a_524_n943# a_466_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_644_607# a_524_553# a_466_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n524_607# a_n644_553# a_n702_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_352_n389# a_232_n445# a_174_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_644_n389# a_524_n445# a_466_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n232_n887# a_n352_n943# a_n410_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_644_109# a_524_55# a_466_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n524_n887# a_n644_n943# a_n702_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_352_607# a_232_553# a_174_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n524_109# a_n644_55# a_n702_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n232_607# a_n352_553# a_n410_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n232_n389# a_n352_n445# a_n410_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n524_n389# a_n644_n445# a_n702_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_60_607# a_n60_553# a_n118_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_352_109# a_232_55# a_174_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n232_109# a_n352_55# a_n410_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_60_n887# a_n60_n943# a_n118_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_60_109# a_n60_55# a_n118_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_352_n887# a_232_n943# a_174_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_644_109# a_758_n887# 0.33fF
C1 a_758_n887# a_n994_n887# 0.07fF
C2 a_466_n887# a_n232_n887# 0.03fF
C3 a_174_n887# a_n994_n887# 0.04fF
C4 a_644_109# a_174_109# 0.04fF
C5 a_174_109# a_n994_n887# 0.04fF
C6 a_524_n943# a_n994_n887# 0.01fF
C7 a_466_109# a_758_n887# 0.12fF
C8 a_174_n389# a_352_n389# 0.13fF
C9 a_352_109# a_n118_109# 0.04fF
C10 a_60_607# a_n524_607# 0.03fF
C11 a_466_109# a_174_109# 0.07fF
C12 a_466_n887# a_n524_n887# 0.02fF
C13 a_174_607# a_60_607# 0.25fF
C14 a_524_553# a_524_n445# 0.03fF
C15 a_466_n887# a_758_n887# 0.12fF
C16 a_n60_n943# a_n994_n887# 0.01fF
C17 a_n702_n389# a_n702_n887# 0.01fF
C18 a_n410_109# a_n232_109# 0.13fF
C19 a_n702_n887# a_n702_109# 0.00fF
C20 a_232_n943# a_n352_n943# 0.02fF
C21 a_644_n887# a_60_n887# 0.03fF
C22 a_466_607# a_352_607# 0.25fF
C23 a_n118_607# a_n994_n887# 0.05fF
C24 a_n118_n389# a_352_n389# 0.04fF
C25 a_644_109# a_n524_109# 0.02fF
C26 a_524_55# a_n352_55# 0.01fF
C27 a_466_n887# a_174_n887# 0.07fF
C28 a_n524_109# a_n994_n887# 0.12fF
C29 a_232_553# a_n352_553# 0.02fF
C30 a_758_n887# a_n60_n445# 0.01fF
C31 a_352_n887# a_n702_n887# 0.02fF
C32 a_n644_n943# a_n352_n943# 0.04fF
C33 a_n702_607# a_n524_607# 0.13fF
C34 a_644_607# a_758_n887# 0.33fF
C35 a_n524_109# a_466_109# 0.02fF
C36 a_n232_607# a_n232_n887# 0.00fF
C37 a_174_607# a_n702_607# 0.02fF
C38 a_n702_n389# a_466_n389# 0.02fF
C39 a_n702_n389# a_n702_607# 0.00fF
C40 a_n702_109# a_n702_607# 0.01fF
C41 a_n60_55# a_758_n887# 0.01fF
C42 a_174_n389# a_758_n887# 0.06fF
C43 a_466_607# a_n410_607# 0.02fF
C44 a_n994_n887# a_524_55# 0.01fF
C45 a_n60_553# a_n994_n887# 0.01fF
C46 a_n644_553# a_n644_55# 0.15fF
C47 a_n60_n943# a_n60_n445# 0.15fF
C48 a_174_n389# a_174_n887# 0.01fF
C49 a_644_n887# a_n232_n887# 0.02fF
C50 a_174_109# a_174_n389# 0.01fF
C51 a_n232_607# a_758_n887# 0.04fF
C52 a_60_607# a_n994_n887# 0.04fF
C53 a_n702_n887# a_n994_n887# 0.33fF
C54 a_n118_n389# a_758_n887# 0.04fF
C55 a_n118_109# a_60_109# 0.13fF
C56 a_n118_607# a_644_607# 0.03fF
C57 a_n60_55# a_n60_n943# 0.03fF
C58 a_n232_n887# a_60_n887# 0.07fF
C59 a_n410_n389# a_466_n389# 0.02fF
C60 a_644_n887# a_n524_n887# 0.02fF
C61 a_644_n887# a_758_n887# 0.33fF
C62 a_232_n943# a_n994_n887# 0.01fF
C63 a_n60_553# a_n60_n445# 0.03fF
C64 a_644_n887# a_174_n887# 0.04fF
C65 a_466_n389# a_n994_n887# 0.03fF
C66 a_n702_607# a_n994_n887# 0.33fF
C67 a_n352_553# a_n352_n445# 0.03fF
C68 a_758_n887# a_n644_55# 0.01fF
C69 a_60_n887# a_n524_n887# 0.03fF
C70 a_n644_n943# a_n994_n887# 0.05fF
C71 a_466_n887# a_n702_n887# 0.02fF
C72 a_n118_607# a_n232_607# 0.25fF
C73 a_232_55# a_n352_55# 0.02fF
C74 a_758_n887# a_60_n887# 0.05fF
C75 a_n118_607# a_n118_n389# 0.00fF
C76 a_352_109# a_n702_109# 0.02fF
C77 a_466_109# a_466_n389# 0.01fF
C78 a_n524_n389# a_n524_607# 0.00fF
C79 a_n60_55# a_n60_553# 0.15fF
C80 a_n60_55# a_524_55# 0.02fF
C81 a_n410_109# a_n410_n887# 0.00fF
C82 a_60_n887# a_174_n887# 0.25fF
C83 a_n702_n389# a_644_n389# 0.01fF
C84 a_n702_n389# a_n524_n389# 0.13fF
C85 a_n410_109# a_n410_607# 0.01fF
C86 a_352_109# a_352_n887# 0.00fF
C87 a_60_607# a_644_607# 0.03fF
C88 a_232_553# a_232_n445# 0.03fF
C89 a_352_n389# a_758_n887# 0.08fF
C90 a_466_n887# a_466_n389# 0.01fF
C91 a_758_n887# a_n644_553# 0.01fF
C92 a_232_55# a_n994_n887# 0.01fF
C93 a_n232_n887# a_n524_n887# 0.07fF
C94 a_n644_n445# a_n994_n887# 0.05fF
C95 a_n410_109# a_n118_109# 0.07fF
C96 a_758_n887# a_n232_n887# 0.04fF
C97 a_n118_109# a_n232_109# 0.25fF
C98 a_60_607# a_n232_607# 0.07fF
C99 a_n702_607# a_644_607# 0.01fF
C100 a_n410_n389# a_644_n389# 0.02fF
C101 a_n232_n887# a_174_n887# 0.05fF
C102 a_n410_n389# a_n524_n389# 0.25fF
C103 a_n232_n389# a_n702_n389# 0.04fF
C104 a_174_n389# a_466_n389# 0.07fF
C105 a_644_109# a_352_109# 0.07fF
C106 a_352_109# a_n994_n887# 0.03fF
C107 a_758_n887# a_n524_n887# 0.03fF
C108 a_n644_55# a_524_55# 0.01fF
C109 a_644_109# a_644_n389# 0.01fF
C110 a_644_n389# a_n994_n887# 0.02fF
C111 a_n702_n887# a_644_n887# 0.01fF
C112 a_174_n887# a_n524_n887# 0.03fF
C113 a_n524_n389# a_n994_n887# 0.12fF
C114 a_466_607# a_n524_607# 0.02fF
C115 a_466_109# a_352_109# 0.25fF
C116 a_n702_607# a_n232_607# 0.04fF
C117 a_524_553# a_n994_n887# 0.01fF
C118 a_758_n887# a_174_n887# 0.06fF
C119 a_174_607# a_466_607# 0.07fF
C120 a_174_109# a_758_n887# 0.06fF
C121 a_n644_n445# a_n60_n445# 0.02fF
C122 a_n118_n389# a_466_n389# 0.03fF
C123 a_524_n943# a_758_n887# 0.05fF
C124 a_n702_109# a_60_109# 0.03fF
C125 a_60_607# a_60_n887# 0.00fF
C126 a_174_109# a_174_n887# 0.00fF
C127 a_n410_n389# a_n232_n389# 0.13fF
C128 a_n702_n887# a_60_n887# 0.03fF
C129 a_n118_n887# a_n410_n887# 0.07fF
C130 a_n60_553# a_n644_553# 0.02fF
C131 a_n352_n943# a_n352_553# 0.01fF
C132 a_n352_n445# a_232_n445# 0.02fF
C133 a_n60_55# a_232_55# 0.04fF
C134 a_232_n445# a_524_n445# 0.04fF
C135 a_n410_607# a_352_607# 0.03fF
C136 a_n60_n943# a_758_n887# 0.01fF
C137 a_n524_109# a_n524_n887# 0.00fF
C138 a_n118_607# a_758_n887# 0.04fF
C139 a_n232_n389# a_n994_n887# 0.06fF
C140 a_n524_109# a_758_n887# 0.03fF
C141 a_n644_n943# a_n644_55# 0.03fF
C142 a_n60_n943# a_524_n943# 0.02fF
C143 a_n410_n887# a_n410_607# 0.00fF
C144 a_n524_109# a_174_109# 0.03fF
C145 a_644_607# a_644_n389# 0.00fF
C146 a_n118_109# a_n118_n887# 0.00fF
C147 a_n702_n887# a_n232_n887# 0.04fF
C148 a_174_n389# a_644_n389# 0.04fF
C149 a_352_n389# a_466_n389# 0.25fF
C150 a_466_607# a_n994_n887# 0.03fF
C151 a_n352_553# a_n352_55# 0.15fF
C152 a_n524_n389# a_174_n389# 0.03fF
C153 a_644_109# a_60_109# 0.03fF
C154 a_n60_553# a_758_n887# 0.01fF
C155 a_60_109# a_n994_n887# 0.04fF
C156 a_758_n887# a_524_55# 0.05fF
C157 a_n644_n943# a_n644_553# 0.01fF
C158 a_232_55# a_n644_55# 0.01fF
C159 a_466_109# a_466_607# 0.01fF
C160 a_524_n943# a_524_55# 0.03fF
C161 a_n702_n887# a_n524_n887# 0.13fF
C162 a_n410_109# a_n702_109# 0.07fF
C163 a_466_109# a_60_109# 0.05fF
C164 a_60_607# a_758_n887# 0.05fF
C165 a_n644_n445# a_n644_55# 0.15fF
C166 a_n118_n389# a_644_n389# 0.03fF
C167 a_n702_n887# a_758_n887# 0.02fF
C168 a_n702_109# a_n232_109# 0.04fF
C169 a_n524_n389# a_n118_n389# 0.05fF
C170 a_n702_n389# a_60_n389# 0.03fF
C171 a_n352_553# a_n994_n887# 0.02fF
C172 a_n702_n887# a_174_n887# 0.02fF
C173 a_n352_n445# a_524_n445# 0.01fF
C174 a_466_607# a_466_n887# 0.00fF
C175 a_n60_n943# a_n60_553# 0.01fF
C176 a_644_n887# a_644_n389# 0.01fF
C177 a_n232_n389# a_174_n389# 0.05fF
C178 a_232_n943# a_758_n887# 0.02fF
C179 a_466_n389# a_758_n887# 0.12fF
C180 a_n702_607# a_758_n887# 0.02fF
C181 a_n644_n445# a_n644_553# 0.03fF
C182 a_n644_n943# a_758_n887# 0.01fF
C183 a_n410_n389# a_n410_109# 0.01fF
C184 a_466_607# a_644_607# 0.13fF
C185 a_232_n943# a_524_n943# 0.04fF
C186 a_n232_n389# a_n232_607# 0.00fF
C187 a_n118_607# a_60_607# 0.13fF
C188 a_n232_n389# a_n118_n389# 0.25fF
C189 a_n410_n389# a_60_n389# 0.04fF
C190 a_352_109# a_352_n389# 0.01fF
C191 a_n644_n943# a_524_n943# 0.01fF
C192 a_644_109# a_n410_109# 0.02fF
C193 a_n410_109# a_n994_n887# 0.08fF
C194 a_n60_n943# a_232_n943# 0.04fF
C195 a_352_n389# a_644_n389# 0.07fF
C196 a_n524_n389# a_352_n389# 0.02fF
C197 a_644_109# a_n232_109# 0.02fF
C198 a_n994_n887# a_n232_109# 0.06fF
C199 a_60_n389# a_n994_n887# 0.04fF
C200 a_466_607# a_n232_607# 0.03fF
C201 a_n60_n943# a_n644_n943# 0.02fF
C202 a_466_109# a_n410_109# 0.02fF
C203 a_n118_607# a_n702_607# 0.03fF
C204 a_232_55# a_758_n887# 0.02fF
C205 a_n644_553# a_524_553# 0.01fF
C206 a_n524_607# a_352_607# 0.02fF
C207 a_466_109# a_n232_109# 0.03fF
C208 a_174_607# a_352_607# 0.13fF
C209 a_n644_n445# a_758_n887# 0.01fF
C210 a_352_n887# a_352_607# 0.00fF
C211 a_352_n887# a_n118_n887# 0.04fF
C212 a_n232_n389# a_352_n389# 0.03fF
C213 a_352_109# a_758_n887# 0.08fF
C214 a_n524_607# a_n410_607# 0.25fF
C215 a_n524_n389# a_n524_n887# 0.01fF
C216 a_644_n389# a_758_n887# 0.33fF
C217 a_174_607# a_n410_607# 0.03fF
C218 a_n524_n389# a_758_n887# 0.03fF
C219 a_232_553# a_n994_n887# 0.01fF
C220 a_352_109# a_174_109# 0.13fF
C221 a_60_109# a_60_n887# 0.00fF
C222 a_n994_n887# a_232_n445# 0.01fF
C223 a_n352_n943# a_n352_n445# 0.15fF
C224 a_758_n887# a_524_553# 0.05fF
C225 a_352_n887# a_n410_n887# 0.03fF
C226 a_n702_607# a_60_607# 0.03fF
C227 a_n232_n389# a_n232_n887# 0.01fF
C228 a_n702_n887# a_n702_607# 0.00fF
C229 a_524_n943# a_524_553# 0.01fF
C230 a_60_n389# a_174_n389# 0.25fF
C231 a_n702_109# a_n118_109# 0.03fF
C232 a_n994_n887# a_352_607# 0.03fF
C233 a_n118_n887# a_n994_n887# 0.05fF
C234 a_232_55# a_524_55# 0.04fF
C235 a_n524_109# a_352_109# 0.02fF
C236 a_n410_n389# a_n410_n887# 0.01fF
C237 a_232_n943# a_n644_n943# 0.01fF
C238 a_n232_607# a_n232_109# 0.01fF
C239 a_n232_n389# a_758_n887# 0.04fF
C240 a_n410_n389# a_n410_607# 0.00fF
C241 a_n524_109# a_n524_n389# 0.01fF
C242 a_n118_n389# a_60_n389# 0.13fF
C243 a_n60_n445# a_232_n445# 0.04fF
C244 a_n352_n445# a_n352_55# 0.15fF
C245 a_n352_553# a_n644_553# 0.04fF
C246 a_n994_n887# a_n410_n887# 0.08fF
C247 a_n994_n887# a_n410_607# 0.08fF
C248 a_466_n887# a_n118_n887# 0.03fF
C249 a_466_607# a_758_n887# 0.12fF
C250 a_232_n943# a_232_55# 0.03fF
C251 a_758_n887# a_60_109# 0.05fF
C252 a_n60_553# a_524_553# 0.02fF
C253 a_524_553# a_524_55# 0.15fF
C254 a_n352_n445# a_n994_n887# 0.02fF
C255 a_n994_n887# a_524_n445# 0.01fF
C256 a_644_109# a_n118_109# 0.03fF
C257 a_60_n389# a_60_n887# 0.01fF
C258 a_174_109# a_60_109# 0.25fF
C259 a_n118_109# a_n994_n887# 0.05fF
C260 a_644_607# a_352_607# 0.07fF
C261 a_466_n887# a_n410_n887# 0.02fF
C262 a_n644_n445# a_n644_n943# 0.15fF
C263 a_466_109# a_n118_109# 0.03fF
C264 a_n352_553# a_758_n887# 0.01fF
C265 a_60_n389# a_352_n389# 0.07fF
C266 a_466_607# a_n118_607# 0.03fF
C267 a_n524_109# a_60_109# 0.03fF
C268 a_644_607# a_n410_607# 0.02fF
C269 a_n232_607# a_352_607# 0.03fF
C270 a_466_n389# a_644_n389# 0.13fF
C271 a_n524_n389# a_466_n389# 0.02fF
C272 a_n232_n887# a_n232_109# 0.00fF
C273 a_n60_n445# a_n352_n445# 0.04fF
C274 a_n118_n389# a_n118_n887# 0.01fF
C275 a_n60_n445# a_524_n445# 0.02fF
C276 a_174_607# a_n524_607# 0.03fF
C277 a_644_n887# a_n118_n887# 0.03fF
C278 a_n702_n389# a_n702_109# 0.01fF
C279 a_n410_109# a_758_n887# 0.03fF
C280 a_n232_607# a_n410_607# 0.13fF
C281 a_758_n887# a_n232_109# 0.04fF
C282 a_n352_n943# a_n352_55# 0.03fF
C283 a_60_n389# a_758_n887# 0.05fF
C284 a_232_553# a_n644_553# 0.01fF
C285 a_n410_109# a_174_109# 0.03fF
C286 a_466_607# a_60_607# 0.05fF
C287 a_n232_n389# a_466_n389# 0.03fF
C288 a_n118_n887# a_60_n887# 0.13fF
C289 a_644_n887# a_n410_n887# 0.02fF
C290 a_174_109# a_n232_109# 0.05fF
C291 a_60_607# a_60_109# 0.01fF
C292 a_n352_553# a_n60_553# 0.04fF
C293 a_352_n389# a_352_607# 0.00fF
C294 a_n118_n389# a_n118_109# 0.01fF
C295 a_n410_n389# a_n702_n389# 0.07fF
C296 a_60_n887# a_n410_n887# 0.04fF
C297 a_n352_n943# a_n994_n887# 0.02fF
C298 a_n524_109# a_n410_109# 0.25fF
C299 a_466_607# a_466_n389# 0.00fF
C300 a_466_607# a_n702_607# 0.02fF
C301 a_n524_109# a_n232_109# 0.07fF
C302 a_n524_607# a_n994_n887# 0.12fF
C303 a_174_607# a_n994_n887# 0.04fF
C304 a_n524_n389# a_644_n389# 0.02fF
C305 a_n702_n389# a_n994_n887# 0.33fF
C306 a_644_109# a_n702_109# 0.01fF
C307 a_n232_n887# a_n118_n887# 0.25fF
C308 a_232_553# a_758_n887# 0.02fF
C309 a_n702_109# a_n994_n887# 0.33fF
C310 a_758_n887# a_232_n445# 0.02fF
C311 a_352_n887# a_n994_n887# 0.03fF
C312 a_466_109# a_n702_109# 0.02fF
C313 a_n232_n887# a_n410_n887# 0.13fF
C314 a_n118_n887# a_n524_n887# 0.05fF
C315 a_n994_n887# a_n352_55# 0.02fF
C316 a_758_n887# a_352_607# 0.08fF
C317 a_758_n887# a_n118_n887# 0.04fF
C318 a_n232_n389# a_644_n389# 0.02fF
C319 a_n118_n887# a_174_n887# 0.07fF
C320 a_n410_n389# a_n994_n887# 0.08fF
C321 a_n232_n389# a_n524_n389# 0.07fF
C322 a_60_n389# a_60_607# 0.00fF
C323 a_n524_n887# a_n410_n887# 0.25fF
C324 a_352_n887# a_466_n887# 0.25fF
C325 a_n524_607# a_644_607# 0.02fF
C326 a_758_n887# a_n410_n887# 0.03fF
C327 a_174_607# a_644_607# 0.04fF
C328 a_644_109# a_n994_n887# 0.02fF
C329 a_758_n887# a_n410_607# 0.03fF
C330 a_174_n887# a_n410_n887# 0.03fF
C331 a_352_109# a_60_109# 0.07fF
C332 a_174_607# a_174_n389# 0.00fF
C333 a_n702_n389# a_174_n389# 0.02fF
C334 a_n118_607# a_352_607# 0.04fF
C335 a_n118_607# a_n118_n887# 0.00fF
C336 a_644_109# a_466_109# 0.13fF
C337 a_60_n389# a_466_n389# 0.05fF
C338 a_232_553# a_n60_553# 0.04fF
C339 a_466_109# a_n994_n887# 0.03fF
C340 a_758_n887# a_n352_n445# 0.01fF
C341 a_n524_607# a_n232_607# 0.07fF
C342 a_758_n887# a_524_n445# 0.06fF
C343 a_n118_109# a_758_n887# 0.04fF
C344 a_174_607# a_n232_607# 0.05fF
C345 a_466_n887# a_n994_n887# 0.03fF
C346 a_n60_55# a_n352_55# 0.04fF
C347 a_n702_n389# a_n118_n389# 0.03fF
C348 a_174_109# a_n118_109# 0.07fF
C349 a_524_n943# a_524_n445# 0.15fF
C350 a_n118_607# a_n410_607# 0.07fF
C351 a_n60_n445# a_n994_n887# 0.01fF
C352 a_n352_553# a_524_553# 0.01fF
C353 a_466_109# a_466_n887# 0.00fF
C354 a_n410_n389# a_174_n389# 0.03fF
C355 a_232_n943# a_232_553# 0.01fF
C356 a_644_109# a_644_607# 0.01fF
C357 a_232_n943# a_232_n445# 0.15fF
C358 a_644_607# a_n994_n887# 0.02fF
C359 a_60_607# a_352_607# 0.07fF
C360 a_352_n887# a_644_n887# 0.07fF
C361 a_n702_n887# a_n118_n887# 0.03fF
C362 a_n118_607# a_n118_109# 0.01fF
C363 a_n60_55# a_n994_n887# 0.01fF
C364 a_n524_109# a_n118_109# 0.05fF
C365 a_174_n389# a_n994_n887# 0.04fF
C366 a_n410_n389# a_n118_n389# 0.07fF
C367 a_352_109# a_n410_109# 0.03fF
C368 a_352_109# a_n232_109# 0.03fF
C369 a_352_n887# a_60_n887# 0.07fF
C370 a_n702_n887# a_n410_n887# 0.07fF
C371 a_n232_607# a_n994_n887# 0.06fF
C372 a_n702_n389# a_352_n389# 0.02fF
C373 a_n702_607# a_352_607# 0.02fF
C374 a_60_607# a_n410_607# 0.04fF
C375 a_n644_55# a_n352_55# 0.04fF
C376 a_60_n389# a_644_n389# 0.03fF
C377 a_n118_n389# a_n994_n887# 0.05fF
C378 a_n524_n389# a_60_n389# 0.03fF
C379 a_524_55# a_524_n445# 0.15fF
C380 a_352_n887# a_352_n389# 0.01fF
C381 a_232_553# a_232_55# 0.15fF
C382 a_232_55# a_232_n445# 0.15fF
C383 a_644_109# a_644_n887# 0.00fF
C384 a_644_n887# a_n994_n887# 0.02fF
C385 a_n60_55# a_n60_n445# 0.15fF
C386 a_n644_n445# a_232_n445# 0.01fF
C387 a_n702_607# a_n410_607# 0.07fF
C388 a_n644_55# a_n994_n887# 0.05fF
C389 a_352_n887# a_n232_n887# 0.03fF
C390 a_n352_n943# a_758_n887# 0.01fF
C391 a_n524_607# a_n524_n887# 0.00fF
C392 a_n410_n389# a_352_n389# 0.03fF
C393 a_60_n887# a_n994_n887# 0.04fF
C394 a_n232_n389# a_n232_109# 0.01fF
C395 a_n232_n389# a_60_n389# 0.07fF
C396 a_n524_607# a_758_n887# 0.03fF
C397 a_n352_n943# a_524_n943# 0.01fF
C398 a_174_607# a_758_n887# 0.06fF
C399 a_n702_n389# a_758_n887# 0.02fF
C400 a_466_n887# a_644_n887# 0.13fF
C401 a_n702_109# a_758_n887# 0.02fF
C402 a_n232_607# a_644_607# 0.02fF
C403 a_352_n389# a_n994_n887# 0.03fF
C404 a_352_n887# a_n524_n887# 0.02fF
C405 a_174_607# a_174_n887# 0.00fF
C406 a_174_607# a_174_109# 0.01fF
C407 a_232_553# a_524_553# 0.04fF
C408 a_n644_553# a_n994_n887# 0.05fF
C409 a_n702_109# a_174_109# 0.02fF
C410 a_352_n887# a_758_n887# 0.08fF
C411 a_n410_109# a_60_109# 0.04fF
C412 a_n60_n943# a_n352_n943# 0.04fF
C413 a_352_109# a_352_607# 0.01fF
C414 a_n118_n389# a_174_n389# 0.07fF
C415 a_466_n887# a_60_n887# 0.05fF
C416 a_352_n887# a_174_n887# 0.13fF
C417 a_60_109# a_n232_109# 0.07fF
C418 a_644_n887# a_644_607# 0.00fF
C419 a_60_n389# a_60_109# 0.01fF
C420 a_758_n887# a_n352_55# 0.01fF
C421 a_n232_n887# a_n994_n887# 0.06fF
C422 a_n118_607# a_n524_607# 0.05fF
C423 a_n524_109# a_n524_607# 0.01fF
C424 a_174_607# a_n118_607# 0.07fF
C425 a_n410_n389# a_758_n887# 0.03fF
C426 a_n524_109# a_n702_109# 0.13fF
C427 a_n60_55# a_n644_55# 0.02fF
C428 a_n644_n445# a_n352_n445# 0.04fF
C429 a_n644_n445# a_524_n445# 0.01fF
C430 a_n994_n887# a_n524_n887# 0.12fF
C431 a_644_n887# VSUBS 0.01fF
C432 a_466_n887# VSUBS 0.01fF
C433 a_352_n887# VSUBS 0.01fF
C434 a_174_n887# VSUBS 0.01fF
C435 a_60_n887# VSUBS 0.01fF
C436 a_n118_n887# VSUBS 0.01fF
C437 a_n232_n887# VSUBS 0.01fF
C438 a_n410_n887# VSUBS 0.01fF
C439 a_n524_n887# VSUBS 0.01fF
C440 a_n702_n887# VSUBS 0.01fF
C441 a_524_n943# VSUBS 0.17fF
C442 a_232_n943# VSUBS 0.19fF
C443 a_n60_n943# VSUBS 0.20fF
C444 a_n352_n943# VSUBS 0.21fF
C445 a_n644_n943# VSUBS 0.22fF
C446 a_644_n389# VSUBS 0.01fF
C447 a_466_n389# VSUBS 0.01fF
C448 a_352_n389# VSUBS 0.01fF
C449 a_174_n389# VSUBS 0.01fF
C450 a_60_n389# VSUBS 0.01fF
C451 a_n118_n389# VSUBS 0.01fF
C452 a_n232_n389# VSUBS 0.01fF
C453 a_n410_n389# VSUBS 0.01fF
C454 a_n524_n389# VSUBS 0.01fF
C455 a_n702_n389# VSUBS 0.01fF
C456 a_524_n445# VSUBS 0.16fF
C457 a_232_n445# VSUBS 0.17fF
C458 a_n60_n445# VSUBS 0.18fF
C459 a_n352_n445# VSUBS 0.19fF
C460 a_n644_n445# VSUBS 0.20fF
C461 a_644_109# VSUBS 0.01fF
C462 a_466_109# VSUBS 0.01fF
C463 a_352_109# VSUBS 0.01fF
C464 a_174_109# VSUBS 0.01fF
C465 a_60_109# VSUBS 0.01fF
C466 a_n118_109# VSUBS 0.01fF
C467 a_n232_109# VSUBS 0.01fF
C468 a_n410_109# VSUBS 0.01fF
C469 a_n524_109# VSUBS 0.01fF
C470 a_n702_109# VSUBS 0.01fF
C471 a_524_55# VSUBS 0.17fF
C472 a_232_55# VSUBS 0.18fF
C473 a_n60_55# VSUBS 0.19fF
C474 a_n352_55# VSUBS 0.20fF
C475 a_n644_55# VSUBS 0.21fF
C476 a_644_607# VSUBS 0.02fF
C477 a_466_607# VSUBS 0.02fF
C478 a_352_607# VSUBS 0.02fF
C479 a_174_607# VSUBS 0.02fF
C480 a_60_607# VSUBS 0.02fF
C481 a_n118_607# VSUBS 0.02fF
C482 a_n232_607# VSUBS 0.02fF
C483 a_n410_607# VSUBS 0.02fF
C484 a_n524_607# VSUBS 0.02fF
C485 a_n702_607# VSUBS 0.02fF
C486 a_758_n887# VSUBS 1.37fF
C487 a_524_553# VSUBS 0.20fF
C488 a_232_553# VSUBS 0.22fF
C489 a_n60_553# VSUBS 0.23fF
C490 a_n352_553# VSUBS 0.24fF
C491 a_n644_553# VSUBS 0.25fF
C492 a_n994_n887# VSUBS 1.65fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EZNTQN a_n830_109# a_n652_n887# a_n652_109# a_n772_55#
+ a_118_553# a_594_n389# a_n772_n445# a_60_607# a_772_n887# a_n474_109# a_772_109#
+ a_n296_109# a_n772_553# a_n296_n389# a_594_109# a_n594_55# a_n594_553# a_n474_n887#
+ a_118_n943# a_60_n389# a_n594_n445# a_n60_55# a_n830_607# a_n772_n943# a_416_n389#
+ a_n652_607# a_594_n887# a_652_n445# a_n416_55# a_n474_607# a_772_607# a_n296_607#
+ a_n60_n445# a_594_607# a_n296_n887# a_n118_n389# a_652_553# a_60_n887# a_n238_55#
+ a_474_553# a_n594_n943# a_238_n389# a_n416_n445# a_416_n887# a_474_n445# a_296_553#
+ a_652_n943# a_n830_n389# a_652_55# a_n118_n887# a_n60_n943# a_n118_109# a_n238_n445#
+ a_416_109# a_n416_553# a_296_n445# a_238_109# a_474_55# a_n238_553# a_238_n887#
+ a_n416_n943# a_n1110_n1061# a_474_n943# a_n652_n389# a_n830_n887# a_60_109# a_772_n389#
+ a_n60_553# a_296_55# a_n118_607# a_n238_n943# a_416_607# a_296_n943# a_n474_n389#
+ a_118_n445# a_118_55# a_238_607#
X0 a_n652_109# a_n772_55# a_n830_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_60_n389# a_n60_n445# a_n118_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_594_n389# a_474_n445# a_416_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1110_n1061# a_n1110_n1061# a_772_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n830_n887# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n474_n887# a_n594_n943# a_n652_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_594_607# a_474_553# a_416_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_109# a_n416_55# a_n474_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_416_n887# a_296_n943# a_238_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n474_607# a_n594_553# a_n652_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n296_n887# a_n416_n943# a_n474_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1110_n1061# a_n1110_n1061# a_772_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1110_n1061# a_n1110_n1061# a_772_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_238_607# a_118_553# a_60_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_238_n887# a_118_n943# a_60_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n830_n389# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n474_n389# a_n594_n445# a_n652_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n830_607# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n118_607# a_n238_553# a_n296_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_594_109# a_474_55# a_416_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_416_n389# a_296_n445# a_238_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_772_n887# a_652_n943# a_594_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n474_109# a_n594_55# a_n652_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n296_n389# a_n416_n445# a_n474_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1110_n1061# a_n1110_n1061# a_772_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_238_109# a_118_55# a_60_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_238_n389# a_118_n445# a_60_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_607# a_296_553# a_238_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n830_109# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n118_109# a_n238_55# a_n296_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n118_n887# a_n238_n943# a_n296_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_60_607# a_n60_553# a_n118_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_772_n389# a_652_n445# a_594_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_772_607# a_652_553# a_594_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_n652_n887# a_n772_n943# a_n830_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_594_n887# a_474_n943# a_416_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_n652_607# a_n772_553# a_n830_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_60_n887# a_n60_n943# a_n118_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_416_109# a_296_55# a_238_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n118_n389# a_n238_n445# a_n296_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_60_109# a_n60_55# a_n118_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X41 a_n296_607# a_n416_553# a_n474_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X42 a_772_109# a_652_55# a_594_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_n652_n389# a_n772_n445# a_n830_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_652_553# a_n594_553# 0.01fF
C1 a_n594_n445# a_474_n445# 0.01fF
C2 a_n118_n389# a_n118_n887# 0.00fF
C3 a_n60_n943# a_n416_n943# 0.03fF
C4 a_296_n943# a_296_55# 0.03fF
C5 a_416_109# a_n830_109# 0.01fF
C6 a_60_607# a_594_607# 0.02fF
C7 a_416_607# a_416_n389# 0.00fF
C8 a_n238_55# a_652_55# 0.01fF
C9 a_n474_n389# a_n830_n389# 0.03fF
C10 a_n60_n445# a_n60_55# 0.15fF
C11 a_n60_55# a_118_55# 0.10fF
C12 a_n830_607# a_n830_109# 0.00fF
C13 a_772_607# a_n296_607# 0.01fF
C14 a_60_n887# a_60_109# 0.00fF
C15 a_n118_n887# a_n474_n887# 0.03fF
C16 a_60_n887# a_416_n887# 0.03fF
C17 a_60_109# a_772_109# 0.01fF
C18 a_n118_n389# a_772_n389# 0.01fF
C19 a_238_607# a_594_607# 0.03fF
C20 a_474_n943# a_n594_n943# 0.01fF
C21 a_n118_109# a_60_109# 0.06fF
C22 a_238_n887# a_n474_n887# 0.01fF
C23 a_n60_n943# a_652_n943# 0.01fF
C24 a_n594_n943# a_n594_553# 0.01fF
C25 a_n416_55# a_n594_55# 0.10fF
C26 a_n474_109# a_n296_109# 0.06fF
C27 a_652_553# a_n416_553# 0.01fF
C28 a_n118_n389# a_60_n389# 0.06fF
C29 a_118_55# a_652_55# 0.02fF
C30 a_652_n445# a_n60_n445# 0.01fF
C31 a_n238_n445# a_118_n445# 0.03fF
C32 a_n118_n389# a_n118_607# 0.00fF
C33 a_238_n887# a_238_109# 0.00fF
C34 a_416_n887# a_n652_n887# 0.01fF
C35 a_594_607# a_n118_607# 0.01fF
C36 a_238_607# a_238_109# 0.00fF
C37 a_652_553# a_n238_553# 0.01fF
C38 a_594_n887# a_594_109# 0.00fF
C39 a_n474_109# a_594_109# 0.01fF
C40 a_n60_n445# a_474_n445# 0.02fF
C41 a_n772_553# a_474_553# 0.01fF
C42 a_n772_553# a_n772_n445# 0.03fF
C43 a_296_553# a_n772_553# 0.01fF
C44 a_n60_553# a_652_553# 0.01fF
C45 a_60_607# a_60_109# 0.00fF
C46 a_n474_n389# a_594_n389# 0.01fF
C47 a_652_n445# a_n772_n445# 0.01fF
C48 a_n118_n887# a_416_n887# 0.02fF
C49 a_238_n389# a_n474_n389# 0.01fF
C50 a_238_109# a_n652_109# 0.01fF
C51 a_238_n887# a_416_n887# 0.06fF
C52 a_n416_553# a_n594_553# 0.10fF
C53 a_n60_55# a_296_55# 0.03fF
C54 a_118_553# a_652_553# 0.02fF
C55 a_n118_n389# a_n296_n389# 0.06fF
C56 a_n830_607# a_594_607# 0.01fF
C57 a_n594_n943# a_n594_n445# 0.15fF
C58 a_n830_n887# a_n296_n887# 0.02fF
C59 a_474_55# a_n238_55# 0.01fF
C60 a_n830_n389# a_772_n389# 0.01fF
C61 a_296_n943# a_n416_n943# 0.01fF
C62 a_n594_n943# a_n238_n943# 0.03fF
C63 a_n772_n943# a_n594_n943# 0.10fF
C64 a_n772_n445# a_474_n445# 0.01fF
C65 a_474_553# a_474_n445# 0.03fF
C66 a_n594_553# a_n238_553# 0.03fF
C67 a_238_109# a_416_109# 0.06fF
C68 a_60_n389# a_n830_n389# 0.01fF
C69 a_60_109# a_60_n389# 0.00fF
C70 a_296_55# a_652_55# 0.03fF
C71 a_n594_n445# a_n594_553# 0.03fF
C72 a_594_n887# a_n296_n887# 0.01fF
C73 a_n474_607# a_416_607# 0.01fF
C74 a_474_n943# a_n238_n943# 0.01fF
C75 a_474_55# a_118_55# 0.03fF
C76 a_474_n943# a_n772_n943# 0.01fF
C77 a_296_n943# a_652_n943# 0.03fF
C78 a_n60_553# a_n594_553# 0.02fF
C79 a_60_109# a_n652_109# 0.01fF
C80 a_n594_n445# a_296_n445# 0.01fF
C81 a_118_n943# a_n594_n943# 0.01fF
C82 a_238_109# a_n830_109# 0.01fF
C83 a_118_553# a_n594_553# 0.01fF
C84 a_n416_553# a_n238_553# 0.10fF
C85 a_n416_55# a_n772_55# 0.03fF
C86 a_n652_607# a_416_607# 0.01fF
C87 a_60_n887# a_n830_n887# 0.01fF
C88 a_n296_607# a_n296_109# 0.00fF
C89 a_n772_55# a_n594_55# 0.10fF
C90 a_474_n943# a_118_n943# 0.03fF
C91 a_60_109# a_416_109# 0.03fF
C92 a_238_n887# a_238_n389# 0.00fF
C93 a_652_n445# a_n416_n445# 0.01fF
C94 a_416_n887# a_416_109# 0.00fF
C95 a_n830_607# a_n830_n389# 0.00fF
C96 a_n60_553# a_n416_553# 0.03fF
C97 a_238_n389# a_238_607# 0.00fF
C98 a_474_55# a_474_553# 0.15fF
C99 a_594_n389# a_772_n389# 0.06fF
C100 a_652_553# a_474_553# 0.10fF
C101 a_772_n887# a_n296_n887# 0.01fF
C102 a_n830_n389# a_n296_n389# 0.02fF
C103 a_60_607# a_416_607# 0.03fF
C104 a_238_n389# a_772_n389# 0.02fF
C105 a_296_553# a_652_553# 0.03fF
C106 a_416_n389# a_n652_n389# 0.01fF
C107 a_n474_109# a_n474_n389# 0.00fF
C108 a_60_n887# a_594_n887# 0.02fF
C109 a_n652_n887# a_n830_n887# 0.06fF
C110 a_n238_n943# a_n238_553# 0.01fF
C111 a_594_n389# a_60_n389# 0.02fF
C112 a_118_553# a_n416_553# 0.02fF
C113 a_n474_109# a_772_109# 0.01fF
C114 a_772_109# a_772_607# 0.00fF
C115 a_238_607# a_416_607# 0.06fF
C116 a_238_n389# a_60_n389# 0.06fF
C117 a_n416_n445# a_474_n445# 0.01fF
C118 a_n60_553# a_n238_553# 0.10fF
C119 a_n118_109# a_n474_109# 0.03fF
C120 a_n830_n389# a_n830_109# 0.00fF
C121 a_60_109# a_n830_109# 0.01fF
C122 a_n474_607# a_n474_109# 0.00fF
C123 a_n474_607# a_772_607# 0.01fF
C124 a_n60_n445# a_296_n445# 0.03fF
C125 a_474_55# a_296_55# 0.10fF
C126 a_n772_n943# a_n238_n943# 0.02fF
C127 a_594_n887# a_n652_n887# 0.01fF
C128 a_118_553# a_n238_553# 0.03fF
C129 a_594_109# a_n296_109# 0.01fF
C130 a_416_607# a_n118_607# 0.02fF
C131 a_n238_55# a_n238_553# 0.15fF
C132 a_n118_n887# a_n830_n887# 0.01fF
C133 a_n60_n943# a_296_n943# 0.03fF
C134 a_474_n943# a_474_553# 0.01fF
C135 a_118_553# a_n60_553# 0.10fF
C136 a_474_553# a_n594_553# 0.01fF
C137 a_238_n887# a_n830_n887# 0.01fF
C138 a_n238_55# a_n238_n943# 0.03fF
C139 a_n652_607# a_772_607# 0.01fF
C140 a_60_n887# a_772_n887# 0.01fF
C141 a_296_553# a_n594_553# 0.01fF
C142 a_772_n887# a_772_109# 0.00fF
C143 a_118_n943# a_n238_n943# 0.03fF
C144 a_652_55# a_652_n943# 0.03fF
C145 a_594_n389# a_n296_n389# 0.01fF
C146 a_652_n445# a_652_n943# 0.15fF
C147 a_n118_n887# a_594_n887# 0.01fF
C148 a_118_n943# a_n772_n943# 0.01fF
C149 a_238_n389# a_n296_n389# 0.02fF
C150 a_n296_607# a_n296_n887# 0.00fF
C151 a_652_n445# a_118_n445# 0.02fF
C152 a_60_607# a_772_607# 0.01fF
C153 a_n60_n445# a_n594_n445# 0.02fF
C154 a_n772_n445# a_296_n445# 0.01fF
C155 a_238_n887# a_594_n887# 0.03fF
C156 a_296_553# a_296_n445# 0.03fF
C157 a_416_607# a_416_109# 0.00fF
C158 a_772_n887# a_n652_n887# 0.01fF
C159 a_416_607# a_n830_607# 0.01fF
C160 a_n60_553# a_n60_n445# 0.03fF
C161 a_118_553# a_118_n943# 0.01fF
C162 a_n416_55# a_n60_55# 0.03fF
C163 a_238_607# a_772_607# 0.02fF
C164 a_474_553# a_n416_553# 0.01fF
C165 a_n118_n389# a_n830_n389# 0.01fF
C166 a_n296_n887# a_n296_109# 0.00fF
C167 a_772_607# a_772_n389# 0.00fF
C168 a_n60_55# a_n594_55# 0.02fF
C169 a_296_553# a_n416_553# 0.01fF
C170 a_n474_n389# a_n652_n389# 0.06fF
C171 a_118_n445# a_474_n445# 0.03fF
C172 a_118_553# a_118_55# 0.15fF
C173 a_296_55# a_296_n445# 0.15fF
C174 a_416_n887# a_n474_n887# 0.01fF
C175 a_474_553# a_n238_553# 0.01fF
C176 a_n416_55# a_652_55# 0.01fF
C177 a_n238_55# a_118_55# 0.03fF
C178 a_772_607# a_n118_607# 0.01fF
C179 a_296_553# a_n238_553# 0.02fF
C180 a_652_55# a_n594_55# 0.01fF
C181 a_n772_n445# a_n594_n445# 0.10fF
C182 a_n118_n887# a_772_n887# 0.01fF
C183 a_118_n943# a_118_55# 0.03fF
C184 a_n474_109# a_n652_109# 0.06fF
C185 a_238_109# a_60_109# 0.06fF
C186 a_n652_n887# a_n652_n389# 0.00fF
C187 a_238_n887# a_772_n887# 0.02fF
C188 a_n60_553# a_474_553# 0.02fF
C189 a_n772_n943# a_n772_n445# 0.15fF
C190 a_n830_607# a_n830_n887# 0.00fF
C191 a_296_553# a_n60_553# 0.03fF
C192 a_n60_n943# a_n60_55# 0.03fF
C193 a_772_n887# a_772_n389# 0.00fF
C194 a_n474_607# a_n296_607# 0.06fF
C195 a_118_553# a_474_553# 0.03fF
C196 a_n652_607# a_n652_n389# 0.00fF
C197 a_n474_109# a_416_109# 0.01fF
C198 a_118_553# a_296_553# 0.10fF
C199 a_296_n445# a_n416_n445# 0.01fF
C200 a_772_109# a_n296_109# 0.01fF
C201 a_652_553# a_652_n943# 0.01fF
C202 a_n830_n887# a_n830_109# 0.00fF
C203 a_n830_607# a_772_607# 0.01fF
C204 a_n118_109# a_n296_109# 0.06fF
C205 a_n118_n389# a_594_n389# 0.01fF
C206 a_n594_n943# a_n416_n943# 0.10fF
C207 a_n118_n389# a_238_n389# 0.03fF
C208 a_652_n445# a_n238_n445# 0.01fF
C209 a_594_n389# a_594_607# 0.00fF
C210 a_n416_553# a_n416_n445# 0.03fF
C211 a_n652_607# a_n296_607# 0.03fF
C212 a_474_n943# a_n416_n943# 0.01fF
C213 a_n474_109# a_n830_109# 0.03fF
C214 a_n60_n445# a_n772_n445# 0.01fF
C215 a_772_109# a_594_109# 0.06fF
C216 a_772_n389# a_n652_n389# 0.01fF
C217 a_n118_109# a_594_109# 0.01fF
C218 a_n594_n943# a_652_n943# 0.01fF
C219 a_n238_55# a_296_55# 0.02fF
C220 a_n238_n445# a_474_n445# 0.01fF
C221 a_416_607# a_594_607# 0.06fF
C222 a_60_607# a_n296_607# 0.03fF
C223 a_n474_n389# a_416_n389# 0.01fF
C224 a_n594_n445# a_n416_n445# 0.10fF
C225 a_474_55# a_n416_55# 0.01fF
C226 a_238_n389# a_238_109# 0.00fF
C227 a_60_n389# a_n652_n389# 0.01fF
C228 a_474_55# a_n594_55# 0.01fF
C229 a_238_607# a_n296_607# 0.02fF
C230 a_474_n943# a_652_n943# 0.10fF
C231 a_n60_55# a_n772_55# 0.01fF
C232 a_n652_109# a_n652_n389# 0.00fF
C233 a_296_55# a_118_55# 0.10fF
C234 a_n416_553# a_n416_n943# 0.01fF
C235 a_n772_553# a_n772_55# 0.15fF
C236 a_296_553# a_474_553# 0.10fF
C237 a_n118_607# a_n296_607# 0.06fF
C238 a_118_n445# a_296_n445# 0.10fF
C239 a_n772_55# a_652_55# 0.01fF
C240 a_594_n389# a_n830_n389# 0.01fF
C241 a_60_n887# a_n296_n887# 0.03fF
C242 a_n594_n943# a_n594_55# 0.03fF
C243 a_238_n389# a_n830_n389# 0.01fF
C244 a_n830_n887# a_n474_n887# 0.03fF
C245 a_n296_n389# a_n652_n389# 0.03fF
C246 a_n238_n943# a_n416_n943# 0.10fF
C247 a_594_607# a_594_n887# 0.00fF
C248 a_n772_n943# a_n416_n943# 0.03fF
C249 a_n60_n445# a_n416_n445# 0.03fF
C250 a_n594_553# a_n594_55# 0.15fF
C251 a_416_607# a_416_n887# 0.00fF
C252 a_594_607# a_772_607# 0.06fF
C253 a_n652_n887# a_n296_n887# 0.03fF
C254 a_296_553# a_296_55# 0.15fF
C255 a_n652_109# a_n296_109# 0.03fF
C256 a_594_n887# a_n474_n887# 0.01fF
C257 a_n474_109# a_n474_n887# 0.00fF
C258 a_n830_607# a_n296_607# 0.02fF
C259 a_118_n445# a_n594_n445# 0.01fF
C260 a_416_n389# a_772_n389# 0.03fF
C261 a_n60_n943# a_n594_n943# 0.02fF
C262 a_n296_n389# a_n296_607# 0.00fF
C263 a_n238_n943# a_652_n943# 0.01fF
C264 a_n772_n943# a_652_n943# 0.01fF
C265 a_n474_109# a_238_109# 0.01fF
C266 a_n416_55# a_n416_553# 0.15fF
C267 a_416_109# a_n296_109# 0.01fF
C268 a_n652_109# a_594_109# 0.01fF
C269 a_60_n389# a_416_n389# 0.03fF
C270 a_118_n943# a_n416_n943# 0.02fF
C271 a_474_n943# a_n60_n943# 0.02fF
C272 a_n118_n887# a_n296_n887# 0.06fF
C273 a_n474_607# a_n474_n389# 0.00fF
C274 a_n772_n445# a_n416_n445# 0.03fF
C275 a_n296_n389# a_n296_109# 0.00fF
C276 a_n830_n389# a_n830_n887# 0.00fF
C277 a_n118_109# a_772_109# 0.01fF
C278 a_238_n887# a_n296_n887# 0.02fF
C279 a_416_n887# a_n830_n887# 0.01fF
C280 a_118_553# a_118_n445# 0.03fF
C281 a_238_n389# a_594_n389# 0.03fF
C282 a_772_n887# a_n474_n887# 0.01fF
C283 a_416_109# a_594_109# 0.06fF
C284 a_118_n943# a_652_n943# 0.02fF
C285 a_474_55# a_n772_55# 0.01fF
C286 a_60_n887# a_n652_n887# 0.01fF
C287 a_n594_n445# a_n594_55# 0.15fF
C288 a_n830_109# a_n296_109# 0.02fF
C289 a_118_n943# a_118_n445# 0.15fF
C290 a_n238_n445# a_296_n445# 0.02fF
C291 a_416_n887# a_594_n887# 0.06fF
C292 a_n474_109# a_60_109# 0.02fF
C293 a_416_109# a_416_n389# 0.00fF
C294 a_118_n445# a_n60_n445# 0.10fF
C295 a_n60_55# a_652_55# 0.01fF
C296 a_118_n445# a_118_55# 0.15fF
C297 a_n118_n389# a_n652_n389# 0.02fF
C298 a_416_n389# a_n296_n389# 0.01fF
C299 a_n830_109# a_594_109# 0.01fF
C300 a_n652_607# a_n474_607# 0.06fF
C301 a_n238_55# a_n416_55# 0.10fF
C302 a_60_607# a_60_n887# 0.00fF
C303 a_60_n887# a_n118_n887# 0.06fF
C304 a_n238_55# a_n594_55# 0.03fF
C305 a_n238_n445# a_n238_553# 0.03fF
C306 a_n118_109# a_n118_n887# 0.00fF
C307 a_60_n887# a_238_n887# 0.06fF
C308 a_652_n445# a_652_55# 0.15fF
C309 a_60_607# a_n474_607# 0.02fF
C310 a_n652_607# a_n652_n887# 0.00fF
C311 a_n238_n445# a_n594_n445# 0.03fF
C312 a_n474_n389# a_772_n389# 0.01fF
C313 a_n60_n943# a_n238_n943# 0.10fF
C314 a_296_n943# a_n594_n943# 0.01fF
C315 a_n60_n943# a_n60_553# 0.01fF
C316 a_n60_n943# a_n772_n943# 0.01fF
C317 a_n238_n445# a_n238_n943# 0.15fF
C318 a_772_109# a_772_n389# 0.00fF
C319 a_594_607# a_n296_607# 0.01fF
C320 a_772_n887# a_416_n887# 0.03fF
C321 a_n474_607# a_238_607# 0.01fF
C322 a_n416_55# a_118_55# 0.02fF
C323 a_n118_n887# a_n652_n887# 0.02fF
C324 a_118_n445# a_n772_n445# 0.01fF
C325 a_n474_n389# a_60_n389# 0.02fF
C326 a_118_55# a_n594_55# 0.01fF
C327 a_n296_n389# a_n296_n887# 0.00fF
C328 a_60_n887# a_60_n389# 0.00fF
C329 a_238_n887# a_n652_n887# 0.01fF
C330 a_474_n943# a_296_n943# 0.10fF
C331 a_652_n445# a_474_n445# 0.10fF
C332 a_594_n389# a_594_n887# 0.00fF
C333 a_60_607# a_n652_607# 0.01fF
C334 a_n118_109# a_n118_607# 0.00fF
C335 a_n474_607# a_n118_607# 0.03fF
C336 a_n238_55# a_n238_n445# 0.15fF
C337 a_118_n943# a_n60_n943# 0.10fF
C338 a_772_109# a_n652_109# 0.01fF
C339 a_n652_607# a_238_607# 0.01fF
C340 a_n118_109# a_n652_109# 0.02fF
C341 a_296_n943# a_296_n445# 0.15fF
C342 a_n830_n389# a_n652_n389# 0.06fF
C343 a_416_607# a_772_607# 0.03fF
C344 a_474_55# a_n60_55# 0.02fF
C345 a_238_n887# a_n118_n887# 0.03fF
C346 a_n60_n943# a_n60_n445# 0.15fF
C347 a_238_109# a_n296_109# 0.02fF
C348 a_594_607# a_594_109# 0.00fF
C349 a_60_607# a_238_607# 0.06fF
C350 a_n416_n445# a_n416_n943# 0.15fF
C351 a_n238_n445# a_n60_n445# 0.10fF
C352 a_n652_n887# a_n652_109# 0.00fF
C353 a_772_109# a_416_109# 0.03fF
C354 a_n772_553# a_652_553# 0.01fF
C355 a_n118_n389# a_416_n389# 0.02fF
C356 a_n474_n389# a_n296_n389# 0.06fF
C357 a_n652_607# a_n118_607# 0.02fF
C358 a_238_n887# a_238_607# 0.00fF
C359 a_n118_109# a_416_109# 0.02fF
C360 a_474_55# a_652_55# 0.10fF
C361 a_n474_607# a_n830_607# 0.03fF
C362 a_60_607# a_60_n389# 0.00fF
C363 a_652_553# a_652_55# 0.15fF
C364 a_n652_607# a_n652_109# 0.00fF
C365 a_652_n445# a_652_553# 0.03fF
C366 a_n772_n943# a_n772_55# 0.03fF
C367 a_238_109# a_594_109# 0.03fF
C368 a_60_607# a_n118_607# 0.06fF
C369 a_n118_n887# a_n118_607# 0.00fF
C370 a_n416_55# a_296_55# 0.01fF
C371 a_118_n445# a_n416_n445# 0.02fF
C372 a_594_n887# a_n830_n887# 0.01fF
C373 a_296_55# a_n594_55# 0.01fF
C374 a_296_n943# a_n238_n943# 0.02fF
C375 a_772_109# a_n830_109# 0.01fF
C376 a_60_n389# a_772_n389# 0.01fF
C377 a_60_109# a_n296_109# 0.03fF
C378 a_238_607# a_n118_607# 0.03fF
C379 a_n772_n943# a_296_n943# 0.01fF
C380 a_n118_109# a_n830_109# 0.01fF
C381 a_n238_n445# a_n772_n445# 0.02fF
C382 a_474_55# a_474_n445# 0.15fF
C383 a_n238_55# a_n772_55# 0.02fF
C384 a_n652_607# a_n830_607# 0.06fF
C385 a_594_n389# a_n652_n389# 0.01fF
C386 a_238_n389# a_n652_n389# 0.01fF
C387 a_n772_553# a_n594_553# 0.10fF
C388 a_n474_n887# a_n296_n887# 0.06fF
C389 a_60_109# a_594_109# 0.02fF
C390 a_60_607# a_n830_607# 0.01fF
C391 a_n416_55# a_n416_n445# 0.15fF
C392 a_n772_55# a_118_55# 0.01fF
C393 a_118_n943# a_296_n943# 0.10fF
C394 a_n416_n943# a_652_n943# 0.01fF
C395 a_772_n887# a_n830_n887# 0.01fF
C396 a_238_607# a_n830_607# 0.01fF
C397 a_n830_n389# a_416_n389# 0.01fF
C398 a_416_n887# a_416_n389# 0.00fF
C399 a_772_n389# a_n296_n389# 0.01fF
C400 a_652_n445# a_296_n445# 0.03fF
C401 a_474_n943# a_474_n445# 0.15fF
C402 a_n772_553# a_n416_553# 0.03fF
C403 a_n118_n389# a_n474_n389# 0.03fF
C404 a_772_n887# a_594_n887# 0.06fF
C405 a_416_607# a_n296_607# 0.01fF
C406 a_n830_607# a_n118_607# 0.01fF
C407 a_60_n389# a_n296_n389# 0.03fF
C408 a_772_n887# a_772_607# 0.00fF
C409 a_n118_109# a_n118_n389# 0.00fF
C410 a_416_109# a_n652_109# 0.01fF
C411 a_n772_n445# a_n772_55# 0.15fF
C412 a_n474_n389# a_n474_n887# 0.00fF
C413 a_n772_553# a_n238_553# 0.02fF
C414 a_n416_55# a_n416_n943# 0.03fF
C415 a_n238_n445# a_n416_n445# 0.10fF
C416 a_60_n887# a_n474_n887# 0.02fF
C417 a_296_n445# a_474_n445# 0.10fF
C418 a_n474_607# a_594_607# 0.01fF
C419 a_416_n887# a_n296_n887# 0.01fF
C420 a_n60_553# a_n60_55# 0.15fF
C421 a_n474_607# a_n474_n887# 0.00fF
C422 a_594_n389# a_594_109# 0.00fF
C423 a_n772_553# a_n60_553# 0.01fF
C424 a_n772_n943# a_n772_553# 0.01fF
C425 a_652_n445# a_n594_n445# 0.01fF
C426 a_296_553# a_296_n943# 0.01fF
C427 a_238_109# a_772_109# 0.02fF
C428 a_n652_109# a_n830_109# 0.06fF
C429 a_n118_109# a_238_109# 0.03fF
C430 a_n652_n887# a_n474_n887# 0.06fF
C431 a_n772_55# a_296_55# 0.01fF
C432 a_n238_55# a_n60_55# 0.10fF
C433 a_594_n389# a_416_n389# 0.06fF
C434 a_118_553# a_n772_553# 0.01fF
C435 a_238_n389# a_416_n389# 0.06fF
C436 a_474_55# a_474_n943# 0.03fF
C437 a_n652_607# a_594_607# 0.01fF
C438 a_772_n887# a_n1110_n1061# 0.10fF
C439 a_594_n887# a_n1110_n1061# 0.06fF
C440 a_416_n887# a_n1110_n1061# 0.05fF
C441 a_238_n887# a_n1110_n1061# 0.05fF
C442 a_60_n887# a_n1110_n1061# 0.04fF
C443 a_n118_n887# a_n1110_n1061# 0.04fF
C444 a_n296_n887# a_n1110_n1061# 0.05fF
C445 a_n474_n887# a_n1110_n1061# 0.05fF
C446 a_n652_n887# a_n1110_n1061# 0.06fF
C447 a_n830_n887# a_n1110_n1061# 0.10fF
C448 a_652_n943# a_n1110_n1061# 0.27fF
C449 a_474_n943# a_n1110_n1061# 0.24fF
C450 a_296_n943# a_n1110_n1061# 0.24fF
C451 a_118_n943# a_n1110_n1061# 0.24fF
C452 a_n60_n943# a_n1110_n1061# 0.25fF
C453 a_n238_n943# a_n1110_n1061# 0.26fF
C454 a_n416_n943# a_n1110_n1061# 0.26fF
C455 a_n594_n943# a_n1110_n1061# 0.27fF
C456 a_n772_n943# a_n1110_n1061# 0.32fF
C457 a_772_n389# a_n1110_n1061# 0.10fF
C458 a_594_n389# a_n1110_n1061# 0.06fF
C459 a_416_n389# a_n1110_n1061# 0.05fF
C460 a_238_n389# a_n1110_n1061# 0.04fF
C461 a_60_n389# a_n1110_n1061# 0.04fF
C462 a_n118_n389# a_n1110_n1061# 0.04fF
C463 a_n296_n389# a_n1110_n1061# 0.04fF
C464 a_n474_n389# a_n1110_n1061# 0.05fF
C465 a_n652_n389# a_n1110_n1061# 0.06fF
C466 a_n830_n389# a_n1110_n1061# 0.10fF
C467 a_652_n445# a_n1110_n1061# 0.22fF
C468 a_474_n445# a_n1110_n1061# 0.19fF
C469 a_296_n445# a_n1110_n1061# 0.19fF
C470 a_118_n445# a_n1110_n1061# 0.19fF
C471 a_n60_n445# a_n1110_n1061# 0.20fF
C472 a_n238_n445# a_n1110_n1061# 0.21fF
C473 a_n416_n445# a_n1110_n1061# 0.21fF
C474 a_n594_n445# a_n1110_n1061# 0.22fF
C475 a_n772_n445# a_n1110_n1061# 0.27fF
C476 a_772_109# a_n1110_n1061# 0.10fF
C477 a_594_109# a_n1110_n1061# 0.06fF
C478 a_416_109# a_n1110_n1061# 0.05fF
C479 a_238_109# a_n1110_n1061# 0.05fF
C480 a_60_109# a_n1110_n1061# 0.04fF
C481 a_n118_109# a_n1110_n1061# 0.04fF
C482 a_n296_109# a_n1110_n1061# 0.05fF
C483 a_n474_109# a_n1110_n1061# 0.05fF
C484 a_n652_109# a_n1110_n1061# 0.06fF
C485 a_n830_109# a_n1110_n1061# 0.10fF
C486 a_652_55# a_n1110_n1061# 0.23fF
C487 a_474_55# a_n1110_n1061# 0.20fF
C488 a_296_55# a_n1110_n1061# 0.20fF
C489 a_118_55# a_n1110_n1061# 0.21fF
C490 a_n60_55# a_n1110_n1061# 0.21fF
C491 a_n238_55# a_n1110_n1061# 0.22fF
C492 a_n416_55# a_n1110_n1061# 0.23fF
C493 a_n594_55# a_n1110_n1061# 0.24fF
C494 a_n772_55# a_n1110_n1061# 0.28fF
C495 a_772_607# a_n1110_n1061# 0.10fF
C496 a_594_607# a_n1110_n1061# 0.06fF
C497 a_416_607# a_n1110_n1061# 0.06fF
C498 a_238_607# a_n1110_n1061# 0.05fF
C499 a_60_607# a_n1110_n1061# 0.05fF
C500 a_n118_607# a_n1110_n1061# 0.05fF
C501 a_n296_607# a_n1110_n1061# 0.05fF
C502 a_n474_607# a_n1110_n1061# 0.06fF
C503 a_n652_607# a_n1110_n1061# 0.07fF
C504 a_n830_607# a_n1110_n1061# 0.10fF
C505 a_652_553# a_n1110_n1061# 0.30fF
C506 a_474_553# a_n1110_n1061# 0.27fF
C507 a_296_553# a_n1110_n1061# 0.27fF
C508 a_118_553# a_n1110_n1061# 0.27fF
C509 a_n60_553# a_n1110_n1061# 0.28fF
C510 a_n238_553# a_n1110_n1061# 0.29fF
C511 a_n416_553# a_n1110_n1061# 0.29fF
C512 a_n594_553# a_n1110_n1061# 0.30fF
C513 a_n772_553# a_n1110_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__pfet_01v8_JJWXCM a_n207_n140# a_29_n205# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n205# a_563_n205# a_n741_n140# a_n327_n205# a_n563_n140# a_385_n205#
+ w_n777_n241# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# VSUBS
X0 a_n385_n140# a_n505_n205# a_n563_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n205# a_149_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n205# a_n29_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n327_n205# a_n385_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_563_n205# a_563_n205# a_505_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n29_n140# a_n149_n205# a_n207_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_505_n140# a_385_n205# a_327_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n29_n140# a_n741_n140# 0.01fF
C1 a_n741_n140# a_n327_n205# 0.02fF
C2 a_n29_n140# a_n563_n140# 0.04fF
C3 a_563_n205# a_n149_n205# 0.01fF
C4 a_n29_n140# a_n207_n140# 0.13fF
C5 a_385_n205# a_n741_n140# 0.01fF
C6 a_327_n140# a_n385_n140# 0.03fF
C7 w_n777_n241# a_n385_n140# 0.02fF
C8 a_n29_n140# a_149_n140# 0.13fF
C9 a_563_n205# a_505_n140# 0.06fF
C10 a_207_n205# a_n149_n205# 0.03fF
C11 a_29_n205# a_n327_n205# 0.03fF
C12 a_n149_n205# a_n505_n205# 0.03fF
C13 a_n741_n140# a_n385_n140# 0.03fF
C14 a_29_n205# a_385_n205# 0.03fF
C15 a_n385_n140# a_n563_n140# 0.13fF
C16 a_n385_n140# a_n207_n140# 0.13fF
C17 w_n777_n241# a_n149_n205# 0.17fF
C18 a_563_n205# a_207_n205# 0.02fF
C19 a_563_n205# a_n505_n205# 0.01fF
C20 a_n385_n140# a_149_n140# 0.04fF
C21 a_385_n205# a_n327_n205# 0.01fF
C22 a_n741_n140# a_n149_n205# 0.01fF
C23 a_327_n140# a_505_n140# 0.13fF
C24 w_n777_n241# a_505_n140# 0.02fF
C25 a_563_n205# a_327_n140# 0.03fF
C26 w_n777_n241# a_563_n205# 0.28fF
C27 a_n29_n140# a_n385_n140# 0.06fF
C28 a_207_n205# a_n505_n205# 0.01fF
C29 a_n741_n140# a_505_n140# 0.01fF
C30 a_n563_n140# a_505_n140# 0.02fF
C31 a_563_n205# a_n741_n140# 0.01fF
C32 a_n207_n140# a_505_n140# 0.03fF
C33 a_563_n205# a_n563_n140# 0.01fF
C34 a_29_n205# a_n149_n205# 0.10fF
C35 a_563_n205# a_n207_n140# 0.01fF
C36 w_n777_n241# a_207_n205# 0.15fF
C37 w_n777_n241# a_n505_n205# 0.19fF
C38 a_149_n140# a_505_n140# 0.06fF
C39 a_563_n205# a_149_n140# 0.02fF
C40 a_207_n205# a_n741_n140# 0.01fF
C41 w_n777_n241# a_327_n140# 0.02fF
C42 a_n149_n205# a_n327_n205# 0.10fF
C43 a_29_n205# a_563_n205# 0.01fF
C44 a_n741_n140# a_n505_n205# 0.07fF
C45 a_385_n205# a_n149_n205# 0.02fF
C46 a_n29_n140# a_505_n140# 0.04fF
C47 a_327_n140# a_n741_n140# 0.01fF
C48 w_n777_n241# a_n741_n140# 0.33fF
C49 a_n29_n140# a_563_n205# 0.01fF
C50 a_327_n140# a_n563_n140# 0.02fF
C51 w_n777_n241# a_n563_n140# 0.02fF
C52 a_563_n205# a_n327_n205# 0.01fF
C53 a_327_n140# a_n207_n140# 0.04fF
C54 w_n777_n241# a_n207_n140# 0.02fF
C55 a_29_n205# a_207_n205# 0.10fF
C56 a_29_n205# a_n505_n205# 0.02fF
C57 a_385_n205# a_563_n205# 0.07fF
C58 a_n741_n140# a_n563_n140# 0.06fF
C59 a_327_n140# a_149_n140# 0.13fF
C60 w_n777_n241# a_149_n140# 0.02fF
C61 a_n741_n140# a_n207_n140# 0.02fF
C62 w_n777_n241# a_29_n205# 0.16fF
C63 a_n207_n140# a_n563_n140# 0.06fF
C64 a_207_n205# a_n327_n205# 0.02fF
C65 a_n385_n140# a_505_n140# 0.02fF
C66 a_n327_n205# a_n505_n205# 0.10fF
C67 a_385_n205# a_207_n205# 0.10fF
C68 a_n741_n140# a_149_n140# 0.01fF
C69 a_563_n205# a_n385_n140# 0.01fF
C70 a_385_n205# a_n505_n205# 0.01fF
C71 a_n563_n140# a_149_n140# 0.03fF
C72 a_29_n205# a_n741_n140# 0.01fF
C73 a_n29_n140# a_327_n140# 0.06fF
C74 w_n777_n241# a_n29_n140# 0.02fF
C75 a_n207_n140# a_149_n140# 0.06fF
C76 w_n777_n241# a_n327_n205# 0.18fF
C77 w_n777_n241# a_385_n205# 0.14fF
C78 w_n777_n241# VSUBS 2.25fF
.ends

.subckt sky130_fd_pr__nfet_01v8_LJREPQ a_n149_n195# a_n207_n140# a_207_n195# a_n29_n140#
+ a_149_n140# a_29_n195# a_n385_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_207_n195# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n385_n140# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n385_n140# a_n207_n140# 0.06fF
C1 a_n29_n140# a_207_n195# 0.03fF
C2 a_n385_n140# a_149_n140# 0.02fF
C3 a_n385_n140# a_207_n195# 0.03fF
C4 a_207_n195# a_n149_n195# 0.02fF
C5 a_n385_n140# a_n29_n140# 0.03fF
C6 a_207_n195# a_29_n195# 0.06fF
C7 a_n207_n140# a_149_n140# 0.03fF
C8 a_207_n195# a_n207_n140# 0.02fF
C9 a_n385_n140# a_n149_n195# 0.06fF
C10 a_n29_n140# a_n207_n140# 0.06fF
C11 a_207_n195# a_149_n140# 0.06fF
C12 a_n385_n140# a_29_n195# 0.02fF
C13 a_n29_n140# a_149_n140# 0.06fF
C14 a_29_n195# a_n149_n195# 0.10fF
C15 a_149_n140# VSUBS 0.01fF
C16 a_n29_n140# VSUBS 0.01fF
C17 a_n207_n140# VSUBS 0.02fF
C18 a_207_n195# VSUBS 0.31fF
C19 a_29_n195# VSUBS 0.19fF
C20 a_n149_n195# VSUBS 0.20fF
C21 a_n385_n140# VSUBS 0.33fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_SAWXCM a_n207_n140# a_29_n205# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n205# a_563_n205# a_n741_n140# a_n327_n205# a_n563_n140# a_385_n205#
+ w_n777_n241# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# VSUBS
X0 a_505_n140# a_385_n205# a_327_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n385_n140# a_n505_n205# a_n563_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_327_n140# a_207_n205# a_149_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_149_n140# a_29_n205# a_n29_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n205# a_n385_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_563_n205# a_563_n205# a_505_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n29_n140# a_n149_n205# a_n207_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n741_n140# a_327_n140# 0.01fF
C1 a_505_n140# a_327_n140# 0.13fF
C2 a_29_n205# a_n741_n140# 0.01fF
C3 a_207_n205# a_29_n205# 0.10fF
C4 a_563_n205# a_385_n205# 0.07fF
C5 a_327_n140# a_n207_n140# 0.04fF
C6 w_n777_n241# a_n741_n140# 0.33fF
C7 a_207_n205# w_n777_n241# 0.15fF
C8 a_505_n140# w_n777_n241# 0.02fF
C9 a_563_n205# a_n505_n205# 0.01fF
C10 w_n777_n241# a_n207_n140# 0.02fF
C11 a_n741_n140# a_149_n140# 0.01fF
C12 a_505_n140# a_149_n140# 0.06fF
C13 a_n149_n205# a_n327_n205# 0.10fF
C14 a_149_n140# a_n207_n140# 0.06fF
C15 a_n563_n140# a_327_n140# 0.02fF
C16 a_n29_n140# a_327_n140# 0.06fF
C17 w_n777_n241# a_n563_n140# 0.02fF
C18 a_29_n205# a_n327_n205# 0.03fF
C19 a_n29_n140# w_n777_n241# 0.02fF
C20 a_n385_n140# a_327_n140# 0.03fF
C21 a_563_n205# a_n741_n140# 0.01fF
C22 w_n777_n241# a_n327_n205# 0.18fF
C23 a_207_n205# a_563_n205# 0.02fF
C24 a_563_n205# a_505_n140# 0.06fF
C25 a_149_n140# a_n563_n140# 0.03fF
C26 a_n29_n140# a_149_n140# 0.13fF
C27 a_n505_n205# a_385_n205# 0.01fF
C28 a_563_n205# a_n207_n140# 0.01fF
C29 w_n777_n241# a_n385_n140# 0.02fF
C30 a_149_n140# a_n385_n140# 0.04fF
C31 a_563_n205# a_n563_n140# 0.01fF
C32 a_n149_n205# a_29_n205# 0.10fF
C33 a_n29_n140# a_563_n205# 0.01fF
C34 a_563_n205# a_n327_n205# 0.01fF
C35 a_n149_n205# w_n777_n241# 0.17fF
C36 a_n741_n140# a_385_n205# 0.01fF
C37 a_207_n205# a_385_n205# 0.10fF
C38 a_563_n205# a_n385_n140# 0.01fF
C39 w_n777_n241# a_327_n140# 0.02fF
C40 a_n741_n140# a_n505_n205# 0.07fF
C41 a_207_n205# a_n505_n205# 0.01fF
C42 w_n777_n241# a_29_n205# 0.16fF
C43 a_149_n140# a_327_n140# 0.13fF
C44 w_n777_n241# a_149_n140# 0.02fF
C45 a_563_n205# a_n149_n205# 0.01fF
C46 a_n327_n205# a_385_n205# 0.01fF
C47 a_207_n205# a_n741_n140# 0.01fF
C48 a_505_n140# a_n741_n140# 0.01fF
C49 a_563_n205# a_327_n140# 0.03fF
C50 a_n327_n205# a_n505_n205# 0.10fF
C51 a_563_n205# a_29_n205# 0.01fF
C52 a_n741_n140# a_n207_n140# 0.02fF
C53 a_505_n140# a_n207_n140# 0.03fF
C54 a_563_n205# w_n777_n241# 0.28fF
C55 a_563_n205# a_149_n140# 0.02fF
C56 a_n741_n140# a_n563_n140# 0.06fF
C57 a_n29_n140# a_n741_n140# 0.01fF
C58 a_505_n140# a_n563_n140# 0.02fF
C59 a_n29_n140# a_505_n140# 0.04fF
C60 a_n149_n205# a_385_n205# 0.02fF
C61 a_n741_n140# a_n327_n205# 0.02fF
C62 a_n563_n140# a_n207_n140# 0.06fF
C63 a_207_n205# a_n327_n205# 0.02fF
C64 a_n29_n140# a_n207_n140# 0.13fF
C65 a_n149_n205# a_n505_n205# 0.03fF
C66 a_n741_n140# a_n385_n140# 0.03fF
C67 a_29_n205# a_385_n205# 0.03fF
C68 a_505_n140# a_n385_n140# 0.02fF
C69 w_n777_n241# a_385_n205# 0.14fF
C70 a_29_n205# a_n505_n205# 0.02fF
C71 a_n385_n140# a_n207_n140# 0.13fF
C72 w_n777_n241# a_n505_n205# 0.19fF
C73 a_n29_n140# a_n563_n140# 0.04fF
C74 a_n149_n205# a_n741_n140# 0.01fF
C75 a_n563_n140# a_n385_n140# 0.13fF
C76 a_207_n205# a_n149_n205# 0.03fF
C77 a_n29_n140# a_n385_n140# 0.06fF
C78 w_n777_n241# VSUBS 2.25fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_28TRYY a_385_553# a_n1097_109# a_n149_55# a_919_n445#
+ a_29_55# a_n29_n389# a_n207_n887# a_1097_n943# a_n1555_n1061# a_n1097_n389# a_n327_n445#
+ a_149_n389# a_n207_109# a_385_n445# a_563_55# a_n505_n943# a_n1275_n887# a_327_n887#
+ a_505_109# a_563_n943# a_n505_553# a_n741_n389# a_327_109# a_n327_553# a_n1275_607#
+ a_n1217_55# a_861_n389# a_149_109# a_n149_553# a_n1097_607# a_385_55# a_n149_n445#
+ a_n29_109# a_919_n943# a_n29_n887# a_n327_n943# a_n1097_n887# a_149_n887# a_n207_607#
+ a_207_n445# a_385_n943# a_n563_n389# a_1097_553# a_n1039_55# a_1217_n389# a_207_55#
+ a_n1217_n445# a_505_607# a_n741_n887# a_327_607# a_n861_n445# a_683_n389# a_n861_55#
+ a_149_607# a_861_n887# a_n919_n389# a_207_553# a_n741_109# a_n919_109# a_n29_607#
+ a_n149_n943# a_1217_109# a_n563_109# a_919_55# a_n1217_553# a_n385_n389# a_1039_109#
+ a_1039_n389# a_861_109# a_n1039_n445# a_n385_109# a_207_n943# a_n861_553# a_n683_55#
+ a_n563_n887# a_n1039_553# a_29_n445# a_1217_n887# a_683_109# a_n683_n445# a_n1217_n943#
+ a_n683_553# a_29_553# a_505_n389# a_n861_n943# a_683_n887# a_741_n445# a_n505_55#
+ a_n919_n887# a_n741_607# a_n919_607# a_1217_607# a_n563_607# a_1097_55# a_1097_n445#
+ a_n207_n389# a_n385_n887# a_1039_607# a_1039_n887# a_861_607# a_n1039_n943# a_n385_607#
+ a_29_n943# a_n327_55# a_n1275_n389# a_683_607# a_n505_n445# a_327_n389# a_n683_n943#
+ a_919_553# a_741_553# a_563_n445# a_505_n887# a_563_553# a_741_n943# a_741_55# a_n1275_109#
X0 a_n919_607# a_n1039_553# a_n1097_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1039_607# a_919_553# a_861_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_109# a_29_55# a_n29_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1097_n887# a_n1217_n943# a_n1275_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_683_n887# a_563_n943# a_505_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n207_n389# a_n327_n445# a_n385_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_607# a_n327_553# a_n385_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n1275_109# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=3.248e+12p ps=2.704e+07u w=1.4e+06u l=600000u
X8 a_683_109# a_563_55# a_505_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_1217_n389# a_1097_n445# a_1039_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1275_n389# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n563_109# a_n683_55# a_n741_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1555_n1061# a_n1555_n1061# a_1217_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_n741_n389# a_n861_n445# a_n919_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n29_n887# a_n149_n943# a_n207_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n919_109# a_n1039_55# a_n1097_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_327_109# a_207_55# a_149_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1039_109# a_919_55# a_861_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1097_n389# a_n1217_n445# a_n1275_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_683_n389# a_563_n445# a_505_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_1039_n389# a_919_n445# a_861_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_505_607# a_385_553# a_327_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n207_109# a_n327_55# a_n385_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_n563_n887# a_n683_n943# a_n741_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_1217_607# a_1097_553# a_1039_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n919_n887# a_n1039_n943# a_n1097_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_505_n887# a_385_n943# a_327_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_861_607# a_741_553# a_683_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_n29_n389# a_n149_n445# a_n207_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n385_n887# a_n505_n943# a_n563_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n741_607# a_n861_553# a_n919_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_n1555_n1061# a_n1555_n1061# a_1217_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X32 a_n29_607# a_n149_553# a_n207_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_505_109# a_385_55# a_327_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_327_n887# a_207_n943# a_149_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X35 a_n563_n389# a_n683_n445# a_n741_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_149_n887# a_29_n943# a_n29_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_n1097_607# a_n1217_553# a_n1275_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X38 a_1217_109# a_1097_55# a_1039_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n919_n389# a_n1039_n445# a_n1097_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_505_n389# a_385_n445# a_327_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X41 a_n385_607# a_n505_553# a_n563_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X42 a_861_109# a_741_55# a_683_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_861_n887# a_741_n943# a_683_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X44 a_n385_n389# a_n505_n445# a_n563_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X45 a_n741_109# a_n861_55# a_n919_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X46 a_n1555_n1061# a_n1555_n1061# a_1217_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X47 a_n29_109# a_n149_55# a_n207_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X48 a_327_n389# a_207_n445# a_149_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X49 a_149_n389# a_29_n445# a_n29_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X50 a_149_607# a_29_553# a_n29_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X51 a_n1097_109# a_n1217_55# a_n1275_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X52 a_n207_n887# a_n327_n943# a_n385_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X53 a_n1275_607# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X54 a_683_607# a_563_553# a_505_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X55 a_n385_109# a_n505_55# a_n563_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X56 a_861_n389# a_741_n445# a_683_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X57 a_1217_n887# a_1097_n943# a_1039_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X58 a_n1275_n887# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X59 a_n563_607# a_n683_553# a_n741_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X60 a_n1555_n1061# a_n1555_n1061# a_1217_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X61 a_n741_n887# a_n861_n943# a_n919_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X62 a_327_607# a_207_553# a_149_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X63 a_1039_n887# a_919_n943# a_861_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1039_n445# a_563_n445# 0.01fF
C1 a_385_55# a_1097_55# 0.01fF
C2 a_n149_n943# a_207_n943# 0.03fF
C3 a_n1217_n943# a_n149_n943# 0.01fF
C4 a_n207_n389# a_n741_n389# 0.02fF
C5 a_207_n445# a_n505_n445# 0.01fF
C6 a_149_607# a_683_607# 0.02fF
C7 a_919_n943# a_1097_n943# 0.10fF
C8 a_1039_607# a_n385_607# 0.01fF
C9 a_29_553# a_n505_553# 0.02fF
C10 a_1217_109# a_n207_109# 0.01fF
C11 a_n1217_n943# a_207_n943# 0.01fF
C12 a_n385_109# a_n207_109# 0.06fF
C13 a_n149_553# a_n149_n445# 0.03fF
C14 a_327_n887# a_n1275_n887# 0.01fF
C15 a_n327_553# a_n861_553# 0.02fF
C16 a_n683_553# a_385_553# 0.01fF
C17 a_149_109# a_n1097_109# 0.01fF
C18 a_861_n389# a_n385_n389# 0.01fF
C19 a_1039_n887# a_n385_n887# 0.01fF
C20 a_207_55# a_n149_55# 0.03fF
C21 a_n1217_n445# a_n505_n445# 0.01fF
C22 a_n149_553# a_n505_553# 0.03fF
C23 a_n683_55# a_n683_n943# 0.03fF
C24 a_n207_607# a_683_607# 0.01fF
C25 a_207_n445# a_563_n445# 0.03fF
C26 a_1039_607# a_n563_607# 0.01fF
C27 a_n385_109# a_n563_109# 0.06fF
C28 a_1217_n389# a_327_n389# 0.01fF
C29 a_n1039_55# a_n327_55# 0.01fF
C30 a_29_n445# a_29_55# 0.15fF
C31 a_n919_607# a_n919_109# 0.00fF
C32 a_n741_n389# a_505_n389# 0.01fF
C33 a_n1217_553# a_n1039_553# 0.10fF
C34 a_n385_n389# a_n919_n389# 0.02fF
C35 a_n1097_n389# a_n385_n389# 0.01fF
C36 a_n149_553# a_n149_55# 0.15fF
C37 a_919_55# a_n327_55# 0.01fF
C38 a_919_55# a_919_n943# 0.03fF
C39 a_149_607# a_n207_607# 0.03fF
C40 a_861_109# a_1039_109# 0.06fF
C41 a_861_607# a_1039_607# 0.06fF
C42 a_n207_109# a_327_109# 0.02fF
C43 a_n1217_55# a_n149_55# 0.01fF
C44 a_n741_109# a_n207_109# 0.02fF
C45 a_n207_n389# a_n207_607# 0.00fF
C46 a_563_n943# a_741_n943# 0.10fF
C47 a_327_n887# a_n385_n887# 0.01fF
C48 a_n1097_607# a_505_607# 0.01fF
C49 a_n861_55# a_207_55# 0.01fF
C50 a_n683_55# a_741_55# 0.01fF
C51 a_n327_n445# a_n505_n445# 0.10fF
C52 a_n505_553# a_207_553# 0.01fF
C53 a_n207_n389# a_505_n389# 0.01fF
C54 a_n1039_n943# a_n1039_553# 0.01fF
C55 a_n563_109# a_327_109# 0.01fF
C56 a_741_n943# a_n149_n943# 0.01fF
C57 a_n741_109# a_n563_109# 0.06fF
C58 a_n1275_n887# a_n1275_n389# 0.00fF
C59 a_n385_n389# a_n385_n887# 0.00fF
C60 a_n1039_55# a_563_55# 0.01fF
C61 a_n1275_n389# a_n919_n389# 0.03fF
C62 a_505_109# a_505_n389# 0.00fF
C63 a_1039_n389# a_1217_n389# 0.06fF
C64 a_n1097_n389# a_n1275_n389# 0.06fF
C65 a_741_n943# a_207_n943# 0.02fF
C66 a_n1039_n943# a_29_n943# 0.01fF
C67 a_563_n943# a_385_n943# 0.10fF
C68 a_919_55# a_563_55# 0.03fF
C69 a_327_n887# a_327_n389# 0.00fF
C70 a_505_n887# a_1217_n887# 0.01fF
C71 a_n385_607# a_683_607# 0.01fF
C72 a_207_55# a_207_n445# 0.15fF
C73 a_1097_n943# a_29_n943# 0.01fF
C74 a_207_55# a_1097_55# 0.01fF
C75 a_n919_109# a_n207_109# 0.01fF
C76 a_741_55# a_29_55# 0.01fF
C77 a_n683_553# a_n683_n445# 0.03fF
C78 a_n861_55# a_n1217_55# 0.03fF
C79 a_861_109# a_861_n389# 0.00fF
C80 a_n1097_109# a_505_109# 0.01fF
C81 a_n29_607# a_n1275_607# 0.01fF
C82 a_1039_n887# a_1039_n389# 0.00fF
C83 a_149_607# a_n385_607# 0.02fF
C84 a_n505_553# a_1097_553# 0.01fF
C85 a_n1097_607# a_n29_607# 0.01fF
C86 a_n327_n445# a_563_n445# 0.01fF
C87 a_n149_n943# a_385_n943# 0.02fF
C88 a_n563_n389# a_149_n389# 0.01fF
C89 a_n385_n389# a_327_n389# 0.01fF
C90 a_n861_n445# a_n149_n445# 0.01fF
C91 a_n1039_55# a_n1039_553# 0.15fF
C92 a_385_n445# a_385_n943# 0.15fF
C93 a_207_n943# a_385_n943# 0.10fF
C94 a_n563_109# a_n919_109# 0.03fF
C95 a_n1217_553# a_385_553# 0.01fF
C96 a_505_607# a_1217_607# 0.01fF
C97 a_n1217_n943# a_385_n943# 0.01fF
C98 a_683_607# a_n563_607# 0.01fF
C99 a_385_553# a_n1039_553# 0.01fF
C100 a_n327_n445# a_n327_n943# 0.15fF
C101 a_n861_553# a_n683_553# 0.10fF
C102 a_n861_n943# a_n505_n943# 0.03fF
C103 a_n861_n445# a_741_n445# 0.01fF
C104 a_n149_n445# a_n149_n943# 0.15fF
C105 a_1217_109# a_n29_109# 0.01fF
C106 a_n385_607# a_n207_607# 0.06fF
C107 a_1217_109# a_1217_n389# 0.00fF
C108 a_149_607# a_n563_607# 0.01fF
C109 a_n207_n887# a_n741_n887# 0.02fF
C110 a_n29_n887# a_n919_n887# 0.01fF
C111 a_n385_109# a_n29_109# 0.03fF
C112 a_861_607# a_683_607# 0.06fF
C113 a_29_n445# a_n505_n445# 0.02fF
C114 a_919_553# a_n505_553# 0.01fF
C115 a_n861_n943# a_n683_n943# 0.10fF
C116 a_n1039_55# a_n1039_n943# 0.03fF
C117 a_385_n445# a_n149_n445# 0.02fF
C118 a_1217_109# a_1217_607# 0.00fF
C119 a_683_n389# a_n29_n389# 0.01fF
C120 a_n741_607# a_n741_n389# 0.00fF
C121 a_919_n445# a_919_553# 0.03fF
C122 a_n505_n445# a_n505_n943# 0.15fF
C123 a_n1217_n445# a_n1217_55# 0.15fF
C124 a_861_607# a_149_607# 0.01fF
C125 a_n1275_n389# a_327_n389# 0.01fF
C126 a_n741_607# a_683_607# 0.01fF
C127 a_149_n887# a_149_n389# 0.00fF
C128 a_n29_607# a_n29_109# 0.00fF
C129 a_207_n445# a_207_553# 0.03fF
C130 a_385_n445# a_741_n445# 0.03fF
C131 a_n1275_109# a_n1275_n887# 0.00fF
C132 a_1039_n389# a_n385_n389# 0.01fF
C133 a_n683_55# a_n683_553# 0.15fF
C134 a_919_n445# a_385_n445# 0.02fF
C135 a_n149_n943# a_n149_55# 0.03fF
C136 a_n29_607# a_1217_607# 0.01fF
C137 a_n741_607# a_149_607# 0.01fF
C138 a_n207_607# a_n563_607# 0.03fF
C139 a_861_n887# a_1217_n887# 0.03fF
C140 a_n1039_n445# a_n861_n445# 0.10fF
C141 a_29_n445# a_563_n445# 0.02fF
C142 a_n29_109# a_327_109# 0.03fF
C143 a_683_109# a_n207_109# 0.01fF
C144 a_n741_109# a_n29_109# 0.01fF
C145 a_563_553# a_n327_553# 0.01fF
C146 a_861_607# a_n207_607# 0.01fF
C147 a_n919_607# a_683_607# 0.01fF
C148 a_n505_55# a_n505_553# 0.15fF
C149 a_385_55# a_741_55# 0.03fF
C150 a_149_109# a_n207_109# 0.03fF
C151 a_n861_55# a_n861_n445# 0.15fF
C152 a_1097_55# a_1097_553# 0.15fF
C153 a_n683_55# a_n327_55# 0.03fF
C154 a_n919_607# a_149_607# 0.01fF
C155 a_741_n943# a_385_n943# 0.03fF
C156 a_n741_607# a_n207_607# 0.02fF
C157 a_n1039_n445# a_385_n445# 0.01fF
C158 a_n505_55# a_n149_55# 0.03fF
C159 a_683_109# a_n563_109# 0.01fF
C160 a_1217_n887# a_149_n887# 0.01fF
C161 a_683_n887# a_1217_n887# 0.02fF
C162 a_n207_n887# a_n1275_n887# 0.01fF
C163 a_n505_n943# a_n327_n943# 0.10fF
C164 a_149_109# a_n563_109# 0.01fF
C165 a_1217_n389# a_149_n389# 0.01fF
C166 a_n385_n389# a_n385_109# 0.00fF
C167 a_n683_n943# a_n327_n943# 0.03fF
C168 a_n327_55# a_29_55# 0.03fF
C169 a_n29_109# a_n919_109# 0.01fF
C170 a_207_n445# a_n861_n445# 0.01fF
C171 a_n919_607# a_n207_607# 0.01fF
C172 a_505_n887# a_505_109# 0.00fF
C173 a_n385_607# a_n563_607# 0.06fF
C174 a_n327_553# a_n327_n943# 0.01fF
C175 a_29_553# a_29_n445# 0.03fF
C176 a_n1217_553# a_n861_553# 0.03fF
C177 a_327_n887# a_327_109# 0.00fF
C178 a_n683_55# a_563_55# 0.01fF
C179 a_741_n943# a_741_n445# 0.15fF
C180 a_741_553# a_n327_553# 0.01fF
C181 a_861_607# a_n385_607# 0.01fF
C182 a_n861_553# a_n1039_553# 0.10fF
C183 a_505_n887# a_n29_n887# 0.02fF
C184 a_385_n445# a_207_n445# 0.10fF
C185 a_n1217_n445# a_n861_n445# 0.03fF
C186 a_n505_55# a_n861_55# 0.03fF
C187 a_207_n445# a_207_n943# 0.15fF
C188 a_683_n887# a_683_109# 0.00fF
C189 a_n29_n887# a_n563_n887# 0.02fF
C190 a_n207_n887# a_n385_n887# 0.06fF
C191 a_505_n887# a_505_n389# 0.00fF
C192 a_n563_n389# a_n741_n389# 0.06fF
C193 a_n207_n389# a_n207_109# 0.00fF
C194 a_n741_607# a_n385_607# 0.03fF
C195 a_861_n389# a_n29_n389# 0.01fF
C196 a_149_109# a_149_n887# 0.00fF
C197 a_741_553# a_741_55# 0.15fF
C198 a_563_55# a_29_55# 0.02fF
C199 a_683_n389# a_861_n389# 0.06fF
C200 a_29_553# a_n327_553# 0.03fF
C201 a_1217_n389# a_1217_n887# 0.00fF
C202 a_505_109# a_n207_109# 0.01fF
C203 a_1217_n887# a_1217_607# 0.00fF
C204 a_385_n445# a_n1217_n445# 0.01fF
C205 a_n1217_n445# a_n1217_n943# 0.15fF
C206 a_861_607# a_n563_607# 0.01fF
C207 a_n505_55# a_1097_55# 0.01fF
C208 a_n505_n445# a_1097_n445# 0.01fF
C209 a_n919_607# a_n919_n887# 0.00fF
C210 a_n29_n389# a_n919_n389# 0.01fF
C211 a_n1097_n389# a_n29_n389# 0.01fF
C212 a_n207_607# a_n207_109# 0.00fF
C213 a_1039_n887# a_1217_n887# 0.06fF
C214 a_1217_607# a_1039_607# 0.06fF
C215 a_n919_607# a_n385_607# 0.02fF
C216 a_n207_n389# a_n563_n389# 0.03fF
C217 a_683_n389# a_n919_n389# 0.01fF
C218 a_n149_553# a_n327_553# 0.10fF
C219 a_n327_n445# a_n861_n445# 0.02fF
C220 a_207_55# a_741_55# 0.02fF
C221 a_n741_607# a_n563_607# 0.06fF
C222 a_505_n887# a_n919_n887# 0.01fF
C223 a_n385_n389# a_149_n389# 0.02fF
C224 a_1217_109# a_861_109# 0.03fF
C225 a_n29_n887# a_n1097_n887# 0.01fF
C226 a_741_n445# a_n149_n445# 0.01fF
C227 a_n563_109# a_505_109# 0.01fF
C228 a_861_109# a_n385_109# 0.01fF
C229 a_n919_n887# a_n563_n887# 0.03fF
C230 a_1039_n887# a_1039_607# 0.00fF
C231 a_563_553# a_n683_553# 0.01fF
C232 a_919_n445# a_n149_n445# 0.01fF
C233 a_n29_109# a_683_109# 0.01fF
C234 a_861_607# a_n741_607# 0.01fF
C235 a_683_n887# a_683_607# 0.00fF
C236 a_n149_n445# a_n149_55# 0.15fF
C237 a_29_n943# a_29_55# 0.03fF
C238 a_919_n445# a_741_n445# 0.10fF
C239 a_563_n445# a_1097_n445# 0.02fF
C240 a_149_109# a_n29_109# 0.06fF
C241 a_n1097_109# a_n207_109# 0.01fF
C242 a_385_n445# a_n327_n445# 0.01fF
C243 a_385_55# a_n327_55# 0.01fF
C244 a_n919_607# a_n563_607# 0.03fF
C245 a_1217_n887# a_327_n887# 0.01fF
C246 a_149_n887# a_149_607# 0.00fF
C247 a_149_607# a_n1275_607# 0.01fF
C248 a_n1097_n887# a_n1097_109# 0.00fF
C249 a_n861_553# a_385_553# 0.01fF
C250 a_861_n887# a_n29_n887# 0.01fF
C251 a_n563_n389# a_505_n389# 0.01fF
C252 a_n1097_607# a_149_607# 0.01fF
C253 a_n327_553# a_207_553# 0.02fF
C254 a_n1275_n389# a_149_n389# 0.01fF
C255 a_n563_n887# a_n563_607# 0.00fF
C256 a_861_109# a_327_109# 0.02fF
C257 a_n741_109# a_861_109# 0.01fF
C258 a_n1039_n445# a_n149_n445# 0.01fF
C259 a_n563_109# a_n1097_109# 0.02fF
C260 a_n1039_55# a_n683_55# 0.03fF
C261 a_n1275_109# a_n385_109# 0.01fF
C262 a_n919_n887# a_n1097_n887# 0.06fF
C263 a_327_607# a_327_n389# 0.00fF
C264 a_n741_n887# a_n1275_n887# 0.02fF
C265 a_n919_607# a_n741_607# 0.06fF
C266 a_919_55# a_n683_55# 0.01fF
C267 a_n1275_607# a_n207_607# 0.01fF
C268 a_n29_n389# a_327_n389# 0.03fF
C269 a_741_553# a_n683_553# 0.01fF
C270 a_n1097_607# a_n207_607# 0.01fF
C271 a_683_n887# a_n29_n887# 0.01fF
C272 a_385_55# a_563_55# 0.10fF
C273 a_n29_n887# a_149_n887# 0.06fF
C274 a_683_n389# a_327_n389# 0.03fF
C275 a_563_n943# a_n505_n943# 0.01fF
C276 a_29_n445# a_n861_n445# 0.01fF
C277 a_n327_553# a_1097_553# 0.01fF
C278 a_n1039_55# a_29_55# 0.01fF
C279 a_n683_n943# a_563_n943# 0.01fF
C280 a_1217_607# a_683_607# 0.02fF
C281 a_563_553# a_563_55# 0.15fF
C282 a_919_55# a_29_55# 0.01fF
C283 a_n1275_109# a_327_109# 0.01fF
C284 a_n741_109# a_n1275_109# 0.02fF
C285 a_919_n943# a_n327_n943# 0.01fF
C286 a_29_553# a_n683_553# 0.01fF
C287 a_n327_n943# a_n327_55# 0.03fF
C288 a_207_n445# a_n149_n445# 0.03fF
C289 a_n505_n943# a_n149_n943# 0.03fF
C290 a_n741_n887# a_n385_n887# 0.03fF
C291 a_29_n445# a_385_n445# 0.03fF
C292 a_1217_n389# a_n207_n389# 0.01fF
C293 a_149_607# a_1217_607# 0.01fF
C294 a_n861_55# a_n149_55# 0.01fF
C295 a_n1097_607# a_n1097_109# 0.00fF
C296 a_n683_n943# a_n149_n943# 0.02fF
C297 a_n861_n943# a_29_n943# 0.01fF
C298 a_n505_n943# a_207_n943# 0.01fF
C299 a_n1217_n943# a_n505_n943# 0.01fF
C300 a_207_n445# a_741_n445# 0.02fF
C301 a_n29_109# a_505_109# 0.02fF
C302 a_n563_109# a_n563_607# 0.00fF
C303 a_1039_n389# a_n29_n389# 0.01fF
C304 a_563_55# a_563_n445# 0.15fF
C305 a_n327_553# a_919_553# 0.01fF
C306 a_n563_n389# a_n563_607# 0.00fF
C307 a_919_n445# a_207_n445# 0.01fF
C308 a_505_n887# a_n563_n887# 0.01fF
C309 a_1039_n389# a_683_n389# 0.03fF
C310 a_149_n887# a_n919_n887# 0.01fF
C311 a_n683_n943# a_207_n943# 0.01fF
C312 a_n149_553# a_n683_553# 0.02fF
C313 a_683_n887# a_n919_n887# 0.01fF
C314 a_n1217_n943# a_n683_n943# 0.02fF
C315 a_n1039_n943# a_n861_n943# 0.10fF
C316 a_n1217_n445# a_n149_n445# 0.01fF
C317 a_n1275_607# a_n385_607# 0.01fF
C318 a_563_553# a_n1039_553# 0.01fF
C319 a_1097_55# a_n149_55# 0.01fF
C320 a_n29_n887# a_n29_109# 0.00fF
C321 a_207_55# a_n327_55# 0.02fF
C322 a_1217_607# a_n207_607# 0.01fF
C323 a_n1097_607# a_n385_607# 0.01fF
C324 a_505_607# a_327_607# 0.06fF
C325 a_n1275_109# a_n919_109# 0.03fF
C326 a_861_n887# a_861_607# 0.00fF
C327 a_n505_55# a_n505_n943# 0.03fF
C328 a_n1097_n389# a_n919_n389# 0.06fF
C329 a_1217_n389# a_505_n389# 0.01fF
C330 a_n683_55# a_n683_n445# 0.15fF
C331 a_1039_n887# a_n29_n887# 0.01fF
C332 a_n385_n389# a_n741_n389# 0.03fF
C333 a_n1039_n445# a_207_n445# 0.01fF
C334 a_n29_109# a_n1097_109# 0.01fF
C335 a_n1275_607# a_n563_607# 0.01fF
C336 a_n1217_55# a_n327_55# 0.01fF
C337 a_n683_553# a_207_553# 0.01fF
C338 a_505_n887# a_n1097_n887# 0.01fF
C339 a_n1097_607# a_n563_607# 0.02fF
C340 a_n1275_n887# a_n385_n887# 0.01fF
C341 a_n1097_n887# a_n563_n887# 0.02fF
C342 a_n327_n445# a_n149_n445# 0.10fF
C343 a_207_55# a_563_55# 0.03fF
C344 a_861_109# a_683_109# 0.06fF
C345 a_385_55# a_n1039_55# 0.01fF
C346 a_n29_607# a_327_607# 0.03fF
C347 a_n385_n389# a_n207_n389# 0.06fF
C348 a_n1039_n445# a_n1217_n445# 0.10fF
C349 a_n327_n445# a_741_n445# 0.01fF
C350 a_1039_n389# a_1039_109# 0.00fF
C351 a_n505_55# a_741_55# 0.01fF
C352 a_n29_n887# a_327_n887# 0.03fF
C353 a_385_55# a_919_55# 0.02fF
C354 a_n327_n943# a_29_n943# 0.03fF
C355 a_861_n389# a_327_n389# 0.02fF
C356 a_n563_109# a_n563_n887# 0.00fF
C357 a_1097_553# a_1097_n445# 0.03fF
C358 a_n741_607# a_n1275_607# 0.02fF
C359 a_919_n445# a_n327_n445# 0.01fF
C360 a_385_55# a_385_553# 0.15fF
C361 a_149_109# a_861_109# 0.01fF
C362 a_741_n943# a_n505_n943# 0.01fF
C363 a_n563_n389# a_n563_n887# 0.00fF
C364 a_n29_607# a_n29_n389# 0.00fF
C365 a_1217_607# a_n385_607# 0.01fF
C366 a_n741_n389# a_n1275_n389# 0.02fF
C367 a_861_n887# a_505_n887# 0.03fF
C368 a_n1097_607# a_n741_607# 0.03fF
C369 a_861_n887# a_n563_n887# 0.01fF
C370 a_29_553# a_n1217_553# 0.01fF
C371 a_n1039_n943# a_n327_n943# 0.01fF
C372 a_n683_n943# a_741_n943# 0.01fF
C373 a_327_109# a_327_607# 0.00fF
C374 a_563_553# a_385_553# 0.10fF
C375 a_1097_n943# a_n327_n943# 0.01fF
C376 a_n919_n389# a_327_n389# 0.01fF
C377 a_29_553# a_n1039_553# 0.01fF
C378 a_n1097_n389# a_327_n389# 0.01fF
C379 a_n919_607# a_n1275_607# 0.03fF
C380 a_n207_n389# a_n1275_n389# 0.01fF
C381 a_29_553# a_29_n943# 0.01fF
C382 a_n385_n389# a_505_n389# 0.01fF
C383 a_n919_607# a_n1097_607# 0.06fF
C384 a_n149_553# a_n1217_553# 0.01fF
C385 a_n505_n943# a_385_n943# 0.01fF
C386 a_n1039_n445# a_n327_n445# 0.01fF
C387 a_207_n445# a_n1217_n445# 0.01fF
C388 a_n563_109# a_n207_109# 0.03fF
C389 a_505_n887# a_149_n887# 0.03fF
C390 a_1217_n887# a_n207_n887# 0.01fF
C391 a_505_n887# a_683_n887# 0.06fF
C392 a_149_109# a_n1275_109# 0.01fF
C393 a_149_n887# a_n563_n887# 0.01fF
C394 a_n1217_553# a_n1217_55# 0.15fF
C395 a_683_n887# a_n563_n887# 0.01fF
C396 a_327_n887# a_n919_n887# 0.01fF
C397 a_1039_n389# a_861_n389# 0.06fF
C398 a_919_553# a_n683_553# 0.01fF
C399 a_n149_553# a_n1039_553# 0.01fF
C400 a_n683_n943# a_385_n943# 0.01fF
C401 a_741_n943# a_741_55# 0.03fF
C402 a_29_n445# a_n149_n445# 0.10fF
C403 a_861_607# a_1217_607# 0.03fF
C404 a_1217_109# a_1039_109# 0.06fF
C405 a_n683_55# a_29_55# 0.01fF
C406 a_385_n445# a_1097_n445# 0.01fF
C407 a_n385_109# a_1039_109# 0.01fF
C408 a_n29_n389# a_149_n389# 0.06fF
C409 a_919_n943# a_563_n943# 0.03fF
C410 a_683_n389# a_149_n389# 0.02fF
C411 a_29_n445# a_741_n445# 0.01fF
C412 a_n563_n389# a_n563_109# 0.00fF
C413 a_29_n445# a_919_n445# 0.01fF
C414 a_741_553# a_385_553# 0.03fF
C415 a_n505_553# a_n505_n943# 0.01fF
C416 a_n385_n389# a_n385_607# 0.00fF
C417 a_919_n943# a_919_553# 0.01fF
C418 a_n1217_553# a_207_553# 0.01fF
C419 a_861_109# a_505_109# 0.03fF
C420 a_207_n445# a_n327_n445# 0.02fF
C421 a_919_n943# a_n149_n943# 0.01fF
C422 a_n505_n445# a_n683_n445# 0.10fF
C423 a_207_553# a_n1039_553# 0.01fF
C424 a_n1039_55# a_207_55# 0.01fF
C425 a_149_n887# a_n1097_n887# 0.01fF
C426 a_n741_109# a_n741_n887# 0.00fF
C427 a_327_109# a_1039_109# 0.01fF
C428 a_919_n943# a_207_n943# 0.01fF
C429 a_n1097_607# a_n1097_n887# 0.00fF
C430 a_919_55# a_207_55# 0.01fF
C431 a_n327_553# a_n505_553# 0.10fF
C432 a_29_553# a_385_553# 0.03fF
C433 a_563_55# a_563_n943# 0.03fF
C434 a_n861_553# a_n861_n943# 0.01fF
C435 a_n327_n445# a_n1217_n445# 0.01fF
C436 a_29_n445# a_n1039_n445# 0.01fF
C437 a_1039_607# a_327_607# 0.01fF
C438 a_861_n887# a_683_n887# 0.06fF
C439 a_1039_n887# a_505_n887# 0.02fF
C440 a_861_n887# a_149_n887# 0.01fF
C441 a_n1039_55# a_n1217_55# 0.10fF
C442 a_741_n445# a_741_55# 0.15fF
C443 a_563_n445# a_n683_n445# 0.01fF
C444 a_n505_55# a_n327_55# 0.10fF
C445 a_n149_553# a_385_553# 0.02fF
C446 a_1039_n887# a_n563_n887# 0.01fF
C447 a_563_553# a_n861_553# 0.01fF
C448 a_741_55# a_n149_55# 0.01fF
C449 a_1039_n389# a_327_n389# 0.01fF
C450 a_n29_109# a_n207_109# 0.06fF
C451 a_385_55# a_n683_55# 0.01fF
C452 a_563_n943# a_29_n943# 0.02fF
C453 a_505_n887# a_327_n887# 0.06fF
C454 a_683_n887# a_149_n887# 0.02fF
C455 a_29_n445# a_207_n445# 0.10fF
C456 a_1097_n943# a_1097_553# 0.01fF
C457 a_683_n389# a_683_109# 0.00fF
C458 a_327_n887# a_n563_n887# 0.01fF
C459 a_n1097_607# a_n1275_607# 0.06fF
C460 a_n207_n887# a_n207_n389# 0.00fF
C461 a_n385_109# a_n385_n887# 0.00fF
C462 a_207_553# a_385_553# 0.10fF
C463 a_n29_109# a_n563_109# 0.02fF
C464 a_n505_55# a_563_55# 0.01fF
C465 a_n1039_n943# a_563_n943# 0.01fF
C466 a_n1217_553# a_n1217_n943# 0.01fF
C467 a_n1275_109# a_n1097_109# 0.06fF
C468 a_1097_n943# a_563_n943# 0.02fF
C469 a_919_n943# a_741_n943# 0.10fF
C470 a_385_55# a_29_55# 0.03fF
C471 a_n149_n943# a_29_n943# 0.10fF
C472 a_861_n389# a_149_n389# 0.01fF
C473 a_29_n445# a_n1217_n445# 0.01fF
C474 a_n861_55# a_741_55# 0.01fF
C475 a_29_n943# a_207_n943# 0.10fF
C476 a_n207_n887# a_n207_607# 0.00fF
C477 a_n1039_n943# a_n149_n943# 0.01fF
C478 a_741_553# a_n861_553# 0.01fF
C479 a_n1217_n943# a_29_n943# 0.01fF
C480 a_n149_n445# a_1097_n445# 0.01fF
C481 a_n207_n887# a_n29_n887# 0.06fF
C482 a_1039_607# a_1039_109# 0.00fF
C483 a_1097_n943# a_n149_n943# 0.01fF
C484 a_861_n887# a_1039_n887# 0.06fF
C485 a_861_607# a_861_109# 0.00fF
C486 a_n1039_n943# a_207_n943# 0.01fF
C487 a_1097_553# a_385_553# 0.01fF
C488 a_683_607# a_327_607# 0.03fF
C489 a_n741_n389# a_n29_n389# 0.01fF
C490 a_149_n389# a_n919_n389# 0.01fF
C491 a_n1217_n943# a_n1039_n943# 0.10fF
C492 a_n1097_n389# a_149_n389# 0.01fF
C493 a_327_n887# a_n1097_n887# 0.01fF
C494 a_741_n445# a_1097_n445# 0.03fF
C495 a_919_n943# a_385_n943# 0.02fF
C496 a_1097_n943# a_207_n943# 0.01fF
C497 a_683_n389# a_n741_n389# 0.01fF
C498 a_1097_55# a_741_55# 0.03fF
C499 a_919_n445# a_1097_n445# 0.10fF
C500 a_n919_n389# a_n919_109# 0.00fF
C501 a_149_607# a_327_607# 0.06fF
C502 a_n505_553# a_n683_553# 0.10fF
C503 a_29_553# a_n861_553# 0.01fF
C504 a_683_n389# a_683_607# 0.00fF
C505 a_683_109# a_1039_109# 0.03fF
C506 a_29_n445# a_n327_n445# 0.03fF
C507 a_n207_n389# a_n29_n389# 0.06fF
C508 a_149_109# a_1039_109# 0.01fF
C509 a_1039_n887# a_149_n887# 0.01fF
C510 a_861_n887# a_327_n887# 0.02fF
C511 a_1039_n887# a_683_n887# 0.03fF
C512 a_919_55# a_919_553# 0.15fF
C513 a_919_553# a_385_553# 0.02fF
C514 a_683_n389# a_n207_n389# 0.01fF
C515 a_327_109# a_327_n389# 0.00fF
C516 a_n149_553# a_n861_553# 0.01fF
C517 a_n207_n887# a_n919_n887# 0.01fF
C518 a_n207_607# a_327_607# 0.02fF
C519 a_n683_55# a_207_55# 0.01fF
C520 a_n385_n389# a_n563_n389# 0.06fF
C521 a_919_n445# a_919_n943# 0.15fF
C522 a_385_n445# a_385_553# 0.03fF
C523 a_n327_553# a_n327_n445# 0.03fF
C524 a_n29_n887# a_n29_n389# 0.00fF
C525 a_n327_55# a_n149_55# 0.10fF
C526 a_741_n943# a_29_n943# 0.01fF
C527 a_149_n887# a_327_n887# 0.06fF
C528 a_683_n887# a_327_n887# 0.03fF
C529 a_n741_n887# a_n741_n389# 0.00fF
C530 a_n505_55# a_n1039_55# 0.02fF
C531 a_149_n389# a_327_n389# 0.06fF
C532 a_n29_n389# a_505_n389# 0.02fF
C533 a_29_553# a_29_55# 0.15fF
C534 a_207_55# a_29_55# 0.10fF
C535 a_n683_55# a_n1217_55# 0.02fF
C536 a_683_n389# a_505_n389# 0.06fF
C537 a_n505_55# a_919_55# 0.01fF
C538 a_n861_553# a_207_553# 0.01fF
C539 a_1217_n389# a_1217_607# 0.00fF
C540 a_1217_n887# a_n385_n887# 0.01fF
C541 a_1097_n943# a_741_n943# 0.03fF
C542 a_n563_n389# a_n1275_n389# 0.01fF
C543 a_207_n445# a_1097_n445# 0.01fF
C544 a_1097_55# a_1097_n445# 0.15fF
C545 a_n29_607# a_505_607# 0.02fF
C546 a_29_n943# a_385_n943# 0.03fF
C547 a_1217_109# a_n385_109# 0.01fF
C548 a_861_109# a_n207_109# 0.01fF
C549 a_n385_607# a_327_607# 0.01fF
C550 a_n1217_55# a_29_55# 0.01fF
C551 a_563_55# a_n149_55# 0.01fF
C552 a_n861_n445# a_n683_n445# 0.10fF
C553 a_n861_55# a_n327_55# 0.02fF
C554 a_n1039_n943# a_385_n943# 0.01fF
C555 a_505_109# a_1039_109# 0.02fF
C556 a_n505_n445# a_563_n445# 0.01fF
C557 a_n1217_553# a_n505_553# 0.01fF
C558 a_1039_n389# a_149_n389# 0.01fF
C559 a_n861_n943# a_n327_n943# 0.02fF
C560 a_1097_n943# a_385_n943# 0.01fF
C561 a_861_n389# a_n741_n389# 0.01fF
C562 a_n683_n943# a_n505_n943# 0.10fF
C563 a_861_109# a_n563_109# 0.01fF
C564 a_n29_n887# a_n741_n887# 0.01fF
C565 a_563_553# a_563_n445# 0.03fF
C566 a_n505_553# a_n1039_553# 0.02fF
C567 a_n1275_607# a_n1275_n389# 0.00fF
C568 a_385_n445# a_n683_n445# 0.01fF
C569 a_861_n887# a_861_109# 0.00fF
C570 a_n563_607# a_327_607# 0.01fF
C571 a_1097_55# a_n327_55# 0.01fF
C572 a_1217_109# a_327_109# 0.01fF
C573 a_n385_109# a_327_109# 0.01fF
C574 a_n861_553# a_n861_n445# 0.03fF
C575 a_n741_109# a_n385_109# 0.03fF
C576 a_n1275_109# a_n207_109# 0.01fF
C577 a_1039_n887# a_327_n887# 0.01fF
C578 a_n741_n389# a_n919_n389# 0.06fF
C579 a_n1097_n389# a_n741_n389# 0.03fF
C580 a_505_n887# a_n207_n887# 0.01fF
C581 a_861_607# a_327_607# 0.02fF
C582 a_861_n389# a_n207_n389# 0.01fF
C583 a_1217_n389# a_n385_n389# 0.01fF
C584 a_n861_55# a_563_55# 0.01fF
C585 a_n207_n887# a_n563_n887# 0.03fF
C586 a_741_553# a_563_553# 0.10fF
C587 a_n327_n445# a_1097_n445# 0.01fF
C588 a_n741_607# a_327_607# 0.01fF
C589 a_385_n943# a_385_553# 0.01fF
C590 a_385_55# a_207_55# 0.10fF
C591 a_n1275_109# a_n563_109# 0.01fF
C592 a_n1039_n445# a_n1039_553# 0.03fF
C593 a_n207_n389# a_n919_n389# 0.01fF
C594 a_n1097_n389# a_n207_n389# 0.01fF
C595 a_n919_n887# a_n741_n887# 0.06fF
C596 a_1097_55# a_563_55# 0.02fF
C597 a_n741_109# a_327_109# 0.01fF
C598 a_1039_n389# a_1039_607# 0.00fF
C599 a_29_553# a_563_553# 0.02fF
C600 a_n385_109# a_n919_109# 0.02fF
C601 a_n207_n887# a_n207_109# 0.00fF
C602 a_861_n389# a_505_n389# 0.03fF
C603 a_n1039_n445# a_n1039_n943# 0.15fF
C604 a_n919_607# a_327_607# 0.01fF
C605 a_n207_n887# a_n1097_n887# 0.01fF
C606 a_n29_n887# a_n1275_n887# 0.01fF
C607 a_385_55# a_n1217_55# 0.01fF
C608 a_n327_n445# a_n327_55# 0.15fF
C609 a_n505_553# a_385_553# 0.01fF
C610 a_563_553# a_n149_553# 0.01fF
C611 a_919_n445# a_919_55# 0.15fF
C612 a_n1039_55# a_n149_55# 0.01fF
C613 a_n1275_109# a_n1275_607# 0.00fF
C614 a_505_607# a_1039_607# 0.02fF
C615 a_n919_n389# a_505_n389# 0.01fF
C616 a_n741_n389# a_327_n389# 0.01fF
C617 a_n1097_n389# a_505_n389# 0.01fF
C618 a_919_55# a_n149_55# 0.01fF
C619 a_1217_109# a_1217_n887# 0.00fF
C620 a_n919_109# a_327_109# 0.01fF
C621 a_861_109# a_n29_109# 0.01fF
C622 a_861_n887# a_n207_n887# 0.01fF
C623 a_n505_55# a_n683_55# 0.10fF
C624 a_n741_109# a_n919_109# 0.06fF
C625 a_n1217_553# a_n1217_n445# 0.03fF
C626 a_n1097_n389# a_n1097_109# 0.00fF
C627 a_29_n445# a_1097_n445# 0.01fF
C628 a_n1039_55# a_n1039_n445# 0.15fF
C629 a_n29_n887# a_n385_n887# 0.03fF
C630 a_29_553# a_741_553# 0.01fF
C631 a_n741_n887# a_n741_607# 0.00fF
C632 a_n207_n389# a_327_n389# 0.02fF
C633 a_n919_n887# a_n1275_n887# 0.03fF
C634 a_1097_n943# a_1097_55# 0.03fF
C635 a_563_553# a_207_553# 0.03fF
C636 a_n919_n887# a_n919_n389# 0.00fF
C637 a_n505_55# a_29_55# 0.02fF
C638 a_n861_55# a_n1039_55# 0.10fF
C639 a_n29_607# a_1039_607# 0.01fF
C640 a_n207_n887# a_149_n887# 0.03fF
C641 a_683_n887# a_n207_n887# 0.01fF
C642 a_n683_n943# a_n683_553# 0.01fF
C643 a_741_553# a_n149_553# 0.01fF
C644 a_1217_109# a_683_109# 0.02fF
C645 a_n385_n389# a_n1275_n389# 0.01fF
C646 a_n149_n445# a_n683_n445# 0.02fF
C647 a_n1275_109# a_n29_109# 0.01fF
C648 a_n385_109# a_683_109# 0.01fF
C649 a_n327_553# a_n683_553# 0.03fF
C650 a_n861_n943# a_563_n943# 0.01fF
C651 a_149_109# a_1217_109# 0.01fF
C652 a_861_607# a_861_n389# 0.00fF
C653 a_149_109# a_n385_109# 0.02fF
C654 a_505_n887# a_n741_n887# 0.01fF
C655 a_563_553# a_1097_553# 0.02fF
C656 a_919_n943# a_n505_n943# 0.01fF
C657 a_n861_n943# a_n861_n445# 0.15fF
C658 a_741_n445# a_n683_n445# 0.01fF
C659 a_327_n389# a_505_n389# 0.06fF
C660 a_n919_n887# a_n385_n887# 0.02fF
C661 a_n563_n389# a_n29_n389# 0.02fF
C662 a_n741_n887# a_n563_n887# 0.06fF
C663 a_29_553# a_n149_553# 0.10fF
C664 a_919_n445# a_n683_n445# 0.01fF
C665 a_919_55# a_1097_55# 0.10fF
C666 a_1039_n389# a_n207_n389# 0.01fF
C667 a_n385_n887# a_n385_607# 0.00fF
C668 a_683_n389# a_n563_n389# 0.01fF
C669 a_919_n943# a_n683_n943# 0.01fF
C670 a_207_55# a_n1217_55# 0.01fF
C671 a_n861_n943# a_n149_n943# 0.01fF
C672 a_n505_n445# a_n861_n445# 0.03fF
C673 a_505_607# a_683_607# 0.06fF
C674 a_563_553# a_563_n943# 0.01fF
C675 a_741_553# a_207_553# 0.02fF
C676 a_683_109# a_327_109# 0.03fF
C677 a_n741_109# a_683_109# 0.01fF
C678 a_n327_553# a_n327_55# 0.15fF
C679 a_n861_n943# a_207_n943# 0.01fF
C680 a_n1217_n943# a_n861_n943# 0.03fF
C681 a_505_607# a_149_607# 0.03fF
C682 a_n1275_607# a_327_607# 0.01fF
C683 a_149_109# a_327_109# 0.06fF
C684 a_563_553# a_919_553# 0.03fF
C685 a_385_55# a_385_n445# 0.15fF
C686 a_149_109# a_n741_109# 0.01fF
C687 a_n505_553# a_n861_553# 0.03fF
C688 a_385_n445# a_n505_n445# 0.01fF
C689 a_n1097_607# a_327_607# 0.01fF
C690 a_n1039_n445# a_n683_n445# 0.03fF
C691 a_563_n445# a_563_n943# 0.15fF
C692 a_n207_109# a_1039_109# 0.01fF
C693 a_29_553# a_207_553# 0.10fF
C694 a_207_55# a_207_553# 0.15fF
C695 a_741_55# a_n327_55# 0.01fF
C696 a_1039_n389# a_505_n389# 0.02fF
C697 a_n741_n887# a_n1097_n887# 0.03fF
C698 a_505_607# a_505_109# 0.00fF
C699 a_683_n887# a_683_n389# 0.00fF
C700 a_563_n445# a_n861_n445# 0.01fF
C701 a_741_553# a_1097_553# 0.03fF
C702 a_1039_n887# a_n207_n887# 0.01fF
C703 a_n919_607# a_n919_n389# 0.00fF
C704 a_n29_607# a_683_607# 0.01fF
C705 a_505_607# a_n207_607# 0.01fF
C706 a_385_55# a_n505_55# 0.01fF
C707 a_563_n943# a_n327_n943# 0.01fF
C708 a_683_109# a_n919_109# 0.01fF
C709 a_n505_55# a_n505_n445# 0.15fF
C710 a_n563_109# a_1039_109# 0.01fF
C711 a_149_109# a_149_n389# 0.00fF
C712 a_n149_553# a_207_553# 0.03fF
C713 a_n1275_n887# a_n563_n887# 0.01fF
C714 a_1217_109# a_505_109# 0.01fF
C715 a_n741_109# a_n741_n389# 0.00fF
C716 a_n29_607# a_149_607# 0.06fF
C717 a_861_n887# a_n741_n887# 0.01fF
C718 a_385_n445# a_563_n445# 0.10fF
C719 a_n385_109# a_505_109# 0.01fF
C720 a_149_109# a_n919_109# 0.01fF
C721 a_505_607# a_505_n389# 0.00fF
C722 a_29_553# a_1097_553# 0.01fF
C723 a_n683_55# a_n149_55# 0.02fF
C724 a_29_n445# a_29_n943# 0.15fF
C725 a_207_n445# a_n683_n445# 0.01fF
C726 a_n207_n887# a_327_n887# 0.02fF
C727 a_563_55# a_741_55# 0.10fF
C728 a_n327_n943# a_n149_n943# 0.10fF
C729 a_n505_n943# a_29_n943# 0.02fF
C730 a_741_553# a_919_553# 0.10fF
C731 a_n327_553# a_n1217_553# 0.01fF
C732 a_n861_55# a_n861_553# 0.15fF
C733 a_1217_607# a_327_607# 0.01fF
C734 a_n327_n943# a_207_n943# 0.02fF
C735 a_n683_n943# a_29_n943# 0.01fF
C736 a_n29_109# a_n29_n389# 0.00fF
C737 a_n1217_n943# a_n327_n943# 0.01fF
C738 a_n327_553# a_n1039_553# 0.01fF
C739 a_n1039_n943# a_n505_n943# 0.02fF
C740 a_n1275_109# a_n1275_n389# 0.00fF
C741 a_n861_n943# a_741_n943# 0.01fF
C742 a_n149_553# a_1097_553# 0.01fF
C743 a_1217_n389# a_n29_n389# 0.01fF
C744 a_n29_607# a_n207_607# 0.06fF
C745 a_505_n887# a_n385_n887# 0.01fF
C746 a_n149_55# a_29_55# 0.10fF
C747 a_1217_n389# a_683_n389# 0.02fF
C748 a_n741_n389# a_149_n389# 0.01fF
C749 a_n29_607# a_n29_n887# 0.00fF
C750 a_149_n887# a_n741_n887# 0.01fF
C751 a_683_n887# a_n741_n887# 0.01fF
C752 a_1097_n943# a_n505_n943# 0.01fF
C753 a_n1217_n445# a_n683_n445# 0.02fF
C754 a_n1039_n943# a_n683_n943# 0.03fF
C755 a_n563_n887# a_n385_n887# 0.06fF
C756 a_505_109# a_327_109# 0.06fF
C757 a_29_553# a_919_553# 0.01fF
C758 a_n1275_n887# a_n1097_n887# 0.06fF
C759 a_n741_109# a_505_109# 0.01fF
C760 a_n385_109# a_n1097_109# 0.01fF
C761 a_505_607# a_n385_607# 0.01fF
C762 a_861_n389# a_n563_n389# 0.01fF
C763 a_n1097_n389# a_n1097_n887# 0.00fF
C764 a_n861_55# a_n683_55# 0.10fF
C765 a_861_n887# a_861_n389# 0.00fF
C766 a_149_607# a_149_n389# 0.00fF
C767 a_207_55# a_207_n943# 0.03fF
C768 a_n861_n943# a_385_n943# 0.01fF
C769 a_n207_n389# a_149_n389# 0.03fF
C770 a_n149_553# a_919_553# 0.01fF
C771 a_n563_n389# a_n919_n389# 0.03fF
C772 a_1097_553# a_207_553# 0.01fF
C773 a_327_n887# a_327_607# 0.00fF
C774 a_n1097_n389# a_n563_n389# 0.02fF
C775 a_n149_553# a_n149_n943# 0.01fF
C776 a_n385_109# a_n385_607# 0.00fF
C777 a_385_55# a_385_n943# 0.03fF
C778 a_505_607# a_n563_607# 0.01fF
C779 a_n861_55# a_29_55# 0.01fF
C780 a_n327_n445# a_n683_n445# 0.03fF
C781 a_n1097_n887# a_n385_n887# 0.01fF
C782 a_505_109# a_n919_109# 0.01fF
C783 a_149_109# a_683_109# 0.02fF
C784 a_n1097_109# a_327_109# 0.01fF
C785 a_n741_109# a_n1097_109# 0.03fF
C786 a_n505_55# a_207_55# 0.01fF
C787 a_n29_607# a_n385_607# 0.03fF
C788 a_861_607# a_505_607# 0.03fF
C789 a_n1217_n943# a_n1217_55# 0.03fF
C790 a_n29_109# a_1039_109# 0.01fF
C791 a_n505_n445# a_n149_n445# 0.03fF
C792 a_n1275_n887# a_n1275_607# 0.00fF
C793 a_741_n943# a_n327_n943# 0.01fF
C794 a_149_n389# a_505_n389# 0.03fF
C795 a_149_n887# a_n1275_n887# 0.01fF
C796 a_1097_55# a_29_55# 0.01fF
C797 a_n327_553# a_385_553# 0.01fF
C798 a_919_553# a_207_553# 0.01fF
C799 a_n385_n389# a_n29_n389# 0.03fF
C800 a_1039_607# a_683_607# 0.03fF
C801 a_505_607# a_n741_607# 0.01fF
C802 a_683_n389# a_n385_n389# 0.01fF
C803 a_741_553# a_741_n943# 0.01fF
C804 a_861_n887# a_n385_n887# 0.01fF
C805 a_1039_n887# a_1039_109# 0.00fF
C806 a_n505_n445# a_741_n445# 0.01fF
C807 a_n505_553# a_n505_n445# 0.03fF
C808 a_n505_55# a_n1217_55# 0.01fF
C809 a_149_607# a_1039_607# 0.01fF
C810 a_n1097_n389# a_n1097_607# 0.00fF
C811 a_n29_607# a_n563_607# 0.02fF
C812 a_919_n445# a_n505_n445# 0.01fF
C813 a_207_553# a_207_n943# 0.01fF
C814 a_919_55# a_741_55# 0.10fF
C815 a_385_55# a_n149_55# 0.02fF
C816 a_n1097_109# a_n919_109# 0.06fF
C817 a_563_553# a_n505_553# 0.01fF
C818 a_683_109# a_683_607# 0.00fF
C819 a_n1217_553# a_n683_553# 0.02fF
C820 a_n919_607# a_505_607# 0.01fF
C821 a_861_607# a_n29_607# 0.01fF
C822 a_563_55# a_n327_55# 0.01fF
C823 a_n327_n943# a_385_n943# 0.01fF
C824 a_563_n445# a_n149_n445# 0.01fF
C825 a_n563_n389# a_327_n389# 0.01fF
C826 a_919_553# a_1097_553# 0.10fF
C827 a_1217_n887# a_n29_n887# 0.01fF
C828 a_n683_553# a_n1039_553# 0.03fF
C829 a_n1275_n389# a_n29_n389# 0.01fF
C830 a_683_n887# a_n385_n887# 0.01fF
C831 a_149_n887# a_n385_n887# 0.02fF
C832 a_1217_n389# a_861_n389# 0.03fF
C833 a_327_n887# a_n741_n887# 0.01fF
C834 a_505_n887# a_505_607# 0.00fF
C835 a_n919_n887# a_n919_109# 0.00fF
C836 a_1039_607# a_n207_607# 0.01fF
C837 a_n29_607# a_n741_607# 0.01fF
C838 a_29_n445# a_n683_n445# 0.01fF
C839 a_563_n445# a_741_n445# 0.10fF
C840 a_149_109# a_149_607# 0.00fF
C841 a_n1039_n445# a_n505_n445# 0.02fF
C842 a_919_n445# a_563_n445# 0.03fF
C843 a_n861_55# a_n861_n943# 0.03fF
C844 a_683_109# a_505_109# 0.06fF
C845 a_1097_n943# a_1097_n445# 0.15fF
C846 a_563_n943# a_n149_n943# 0.01fF
C847 a_n683_n943# a_n683_n445# 0.15fF
C848 a_385_55# a_n861_55# 0.01fF
C849 a_n741_109# a_n741_607# 0.00fF
C850 a_149_109# a_505_109# 0.03fF
C851 a_563_n943# a_207_n943# 0.03fF
C852 a_n919_607# a_n29_607# 0.01fF
C853 a_741_553# a_n505_553# 0.01fF
C854 a_741_553# a_741_n445# 0.03fF
C855 a_385_n445# a_n861_n445# 0.01fF
C856 a_1039_n389# a_n563_n389# 0.01fF
C857 a_919_n943# a_29_n943# 0.01fF
C858 a_1217_n887# a_n1555_n1061# 0.10fF
C859 a_1039_n887# a_n1555_n1061# 0.05fF
C860 a_861_n887# a_n1555_n1061# 0.04fF
C861 a_683_n887# a_n1555_n1061# 0.03fF
C862 a_505_n887# a_n1555_n1061# 0.03fF
C863 a_327_n887# a_n1555_n1061# 0.03fF
C864 a_149_n887# a_n1555_n1061# 0.03fF
C865 a_n29_n887# a_n1555_n1061# 0.03fF
C866 a_n207_n887# a_n1555_n1061# 0.03fF
C867 a_n385_n887# a_n1555_n1061# 0.03fF
C868 a_n563_n887# a_n1555_n1061# 0.03fF
C869 a_n741_n887# a_n1555_n1061# 0.03fF
C870 a_n919_n887# a_n1555_n1061# 0.04fF
C871 a_n1097_n887# a_n1555_n1061# 0.05fF
C872 a_n1275_n887# a_n1555_n1061# 0.10fF
C873 a_1097_n943# a_n1555_n1061# 0.27fF
C874 a_919_n943# a_n1555_n1061# 0.23fF
C875 a_741_n943# a_n1555_n1061# 0.23fF
C876 a_563_n943# a_n1555_n1061# 0.24fF
C877 a_385_n943# a_n1555_n1061# 0.24fF
C878 a_207_n943# a_n1555_n1061# 0.25fF
C879 a_29_n943# a_n1555_n1061# 0.26fF
C880 a_n149_n943# a_n1555_n1061# 0.26fF
C881 a_n327_n943# a_n1555_n1061# 0.26fF
C882 a_n505_n943# a_n1555_n1061# 0.26fF
C883 a_n683_n943# a_n1555_n1061# 0.26fF
C884 a_n861_n943# a_n1555_n1061# 0.26fF
C885 a_n1039_n943# a_n1555_n1061# 0.27fF
C886 a_n1217_n943# a_n1555_n1061# 0.32fF
C887 a_1217_n389# a_n1555_n1061# 0.10fF
C888 a_1039_n389# a_n1555_n1061# 0.05fF
C889 a_861_n389# a_n1555_n1061# 0.04fF
C890 a_683_n389# a_n1555_n1061# 0.03fF
C891 a_505_n389# a_n1555_n1061# 0.03fF
C892 a_327_n389# a_n1555_n1061# 0.02fF
C893 a_149_n389# a_n1555_n1061# 0.03fF
C894 a_n29_n389# a_n1555_n1061# 0.03fF
C895 a_n207_n389# a_n1555_n1061# 0.03fF
C896 a_n385_n389# a_n1555_n1061# 0.02fF
C897 a_n563_n389# a_n1555_n1061# 0.03fF
C898 a_n741_n389# a_n1555_n1061# 0.03fF
C899 a_n919_n389# a_n1555_n1061# 0.04fF
C900 a_n1097_n389# a_n1555_n1061# 0.05fF
C901 a_n1275_n389# a_n1555_n1061# 0.10fF
C902 a_1097_n445# a_n1555_n1061# 0.22fF
C903 a_919_n445# a_n1555_n1061# 0.18fF
C904 a_741_n445# a_n1555_n1061# 0.18fF
C905 a_563_n445# a_n1555_n1061# 0.19fF
C906 a_385_n445# a_n1555_n1061# 0.19fF
C907 a_207_n445# a_n1555_n1061# 0.20fF
C908 a_29_n445# a_n1555_n1061# 0.21fF
C909 a_n149_n445# a_n1555_n1061# 0.21fF
C910 a_n327_n445# a_n1555_n1061# 0.21fF
C911 a_n505_n445# a_n1555_n1061# 0.21fF
C912 a_n683_n445# a_n1555_n1061# 0.21fF
C913 a_n861_n445# a_n1555_n1061# 0.21fF
C914 a_n1039_n445# a_n1555_n1061# 0.22fF
C915 a_n1217_n445# a_n1555_n1061# 0.27fF
C916 a_1217_109# a_n1555_n1061# 0.10fF
C917 a_1039_109# a_n1555_n1061# 0.05fF
C918 a_861_109# a_n1555_n1061# 0.04fF
C919 a_683_109# a_n1555_n1061# 0.03fF
C920 a_505_109# a_n1555_n1061# 0.03fF
C921 a_327_109# a_n1555_n1061# 0.03fF
C922 a_149_109# a_n1555_n1061# 0.03fF
C923 a_n29_109# a_n1555_n1061# 0.03fF
C924 a_n207_109# a_n1555_n1061# 0.03fF
C925 a_n385_109# a_n1555_n1061# 0.03fF
C926 a_n563_109# a_n1555_n1061# 0.03fF
C927 a_n741_109# a_n1555_n1061# 0.03fF
C928 a_n919_109# a_n1555_n1061# 0.04fF
C929 a_n1097_109# a_n1555_n1061# 0.06fF
C930 a_n1275_109# a_n1555_n1061# 0.10fF
C931 a_1097_55# a_n1555_n1061# 0.23fF
C932 a_919_55# a_n1555_n1061# 0.20fF
C933 a_741_55# a_n1555_n1061# 0.20fF
C934 a_563_55# a_n1555_n1061# 0.20fF
C935 a_385_55# a_n1555_n1061# 0.21fF
C936 a_207_55# a_n1555_n1061# 0.21fF
C937 a_29_55# a_n1555_n1061# 0.22fF
C938 a_n149_55# a_n1555_n1061# 0.22fF
C939 a_n327_55# a_n1555_n1061# 0.22fF
C940 a_n505_55# a_n1555_n1061# 0.22fF
C941 a_n683_55# a_n1555_n1061# 0.22fF
C942 a_n861_55# a_n1555_n1061# 0.23fF
C943 a_n1039_55# a_n1555_n1061# 0.23fF
C944 a_n1217_55# a_n1555_n1061# 0.28fF
C945 a_1217_607# a_n1555_n1061# 0.10fF
C946 a_1039_607# a_n1555_n1061# 0.06fF
C947 a_861_607# a_n1555_n1061# 0.05fF
C948 a_683_607# a_n1555_n1061# 0.04fF
C949 a_505_607# a_n1555_n1061# 0.03fF
C950 a_327_607# a_n1555_n1061# 0.03fF
C951 a_149_607# a_n1555_n1061# 0.03fF
C952 a_n29_607# a_n1555_n1061# 0.04fF
C953 a_n207_607# a_n1555_n1061# 0.03fF
C954 a_n385_607# a_n1555_n1061# 0.03fF
C955 a_n563_607# a_n1555_n1061# 0.03fF
C956 a_n741_607# a_n1555_n1061# 0.04fF
C957 a_n919_607# a_n1555_n1061# 0.05fF
C958 a_n1097_607# a_n1555_n1061# 0.06fF
C959 a_n1275_607# a_n1555_n1061# 0.10fF
C960 a_1097_553# a_n1555_n1061# 0.30fF
C961 a_919_553# a_n1555_n1061# 0.26fF
C962 a_741_553# a_n1555_n1061# 0.26fF
C963 a_563_553# a_n1555_n1061# 0.27fF
C964 a_385_553# a_n1555_n1061# 0.27fF
C965 a_207_553# a_n1555_n1061# 0.28fF
C966 a_29_553# a_n1555_n1061# 0.29fF
C967 a_n149_553# a_n1555_n1061# 0.29fF
C968 a_n327_553# a_n1555_n1061# 0.29fF
C969 a_n505_553# a_n1555_n1061# 0.29fF
C970 a_n683_553# a_n1555_n1061# 0.29fF
C971 a_n861_553# a_n1555_n1061# 0.29fF
C972 a_n1039_553# a_n1555_n1061# 0.30fF
C973 a_n1217_553# a_n1555_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EL6FQZ a_n1008_n140# a_1306_n140# a_n652_n140# a_652_n194#
+ a_n1662_n194# a_772_n140# a_n1720_n140# a_n60_n194# a_2076_n194# a_1008_n194# a_2196_n140#
+ a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194# a_594_n140# a_n1542_n140#
+ a_1720_n194# a_1840_n140# a_n238_n194# a_n296_n140# a_n1898_n140# a_296_n194# a_2018_n140#
+ a_60_n140# a_n1306_n194# a_n1364_n140# a_1542_n194# a_416_n140# a_n950_n194# a_n2432_n140#
+ a_1662_n140# a_1898_n194# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194# a_238_n140#
+ a_n1186_n140# a_n2254_n140# a_1364_n194# a_n772_n194# a_1484_n140# a_n830_n140#
+ a_830_n194# a_n1840_n194# a_950_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2254_n194# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2254_n140# a_n2432_n140# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_652_n194# a_n950_n194# 0.01fF
C1 a_1008_n194# a_1898_n194# 0.01fF
C2 a_2254_n194# a_950_n140# 0.01fF
C3 a_n594_n194# a_830_n194# 0.01fF
C4 a_2196_n140# a_1484_n140# 0.01fF
C5 a_296_n194# a_n60_n194# 0.03fF
C6 a_1008_n194# a_296_n194# 0.01fF
C7 a_n1542_n140# a_n296_n140# 0.01fF
C8 a_n1720_n140# a_n474_n140# 0.01fF
C9 a_n1186_n140# a_238_n140# 0.01fF
C10 a_1008_n194# a_n60_n194# 0.01fF
C11 a_1720_n194# a_652_n194# 0.01fF
C12 a_1484_n140# a_416_n140# 0.01fF
C13 a_416_n140# a_238_n140# 0.06fF
C14 a_n118_n140# a_1128_n140# 0.01fF
C15 a_2196_n140# a_594_n140# 0.01fF
C16 a_n1364_n140# a_n2076_n140# 0.01fF
C17 a_n1186_n140# a_n1364_n140# 0.06fF
C18 a_n2432_n140# a_n2076_n140# 0.03fF
C19 a_416_n140# a_594_n140# 0.06fF
C20 a_n1186_n140# a_n2432_n140# 0.01fF
C21 a_n830_n140# a_n1008_n140# 0.06fF
C22 a_772_n140# a_1484_n140# 0.01fF
C23 a_238_n140# a_n296_n140# 0.02fF
C24 a_1662_n140# a_1306_n140# 0.03fF
C25 a_772_n140# a_238_n140# 0.02fF
C26 a_n238_n194# a_n416_n194# 0.10fF
C27 a_n1128_n194# a_n238_n194# 0.01fF
C28 a_n2254_n140# a_n2076_n140# 0.06fF
C29 a_n416_n194# a_296_n194# 0.01fF
C30 a_n1364_n140# a_n296_n140# 0.01fF
C31 a_594_n140# a_n296_n140# 0.01fF
C32 a_772_n140# a_594_n140# 0.06fF
C33 a_n1186_n140# a_n2254_n140# 0.01fF
C34 a_n416_n194# a_n60_n194# 0.03fF
C35 a_n1128_n194# a_296_n194# 0.01fF
C36 a_830_n194# a_118_n194# 0.01fF
C37 a_1662_n140# a_2018_n140# 0.03fF
C38 a_1008_n194# a_n416_n194# 0.01fF
C39 a_n830_n140# a_n1898_n140# 0.01fF
C40 a_950_n140# a_238_n140# 0.01fF
C41 a_1484_n140# a_950_n140# 0.02fF
C42 a_n1128_n194# a_n60_n194# 0.01fF
C43 a_1128_n140# a_n474_n140# 0.01fF
C44 a_1186_n194# a_474_n194# 0.01fF
C45 a_1364_n194# a_118_n194# 0.01fF
C46 a_594_n140# a_950_n140# 0.03fF
C47 a_1364_n194# a_830_n194# 0.02fF
C48 a_2254_n194# a_1898_n194# 0.02fF
C49 a_n1542_n140# a_n652_n140# 0.01fF
C50 a_652_n194# a_474_n194# 0.10fF
C51 a_n1186_n140# a_60_n140# 0.01fF
C52 a_416_n140# a_60_n140# 0.03fF
C53 a_2076_n194# a_1898_n194# 0.10fF
C54 a_n118_n140# a_n1542_n140# 0.01fF
C55 a_1008_n194# a_2254_n194# 0.00fF
C56 a_n594_n194# a_n772_n194# 0.10fF
C57 a_1008_n194# a_2076_n194# 0.01fF
C58 a_1186_n194# a_1542_n194# 0.03fF
C59 a_n238_n194# a_n1306_n194# 0.01fF
C60 a_n1542_n140# a_n1720_n140# 0.06fF
C61 a_n1128_n194# a_n416_n194# 0.01fF
C62 a_n652_n140# a_238_n140# 0.01fF
C63 a_60_n140# a_n296_n140# 0.03fF
C64 a_772_n140# a_60_n140# 0.01fF
C65 a_n118_n140# a_1484_n140# 0.01fF
C66 a_n118_n140# a_238_n140# 0.03fF
C67 a_1542_n194# a_652_n194# 0.01fF
C68 a_2196_n140# a_1840_n140# 0.03fF
C69 a_n594_n194# a_n1484_n194# 0.01fF
C70 a_n1306_n194# a_296_n194# 0.01fF
C71 a_n652_n140# a_594_n140# 0.01fF
C72 a_n1364_n140# a_n652_n140# 0.01fF
C73 a_n1662_n194# a_n772_n194# 0.01fF
C74 a_n1306_n194# a_n60_n194# 0.01fF
C75 a_416_n140# a_1840_n140# 0.01fF
C76 a_2254_n194# a_1128_n140# 0.01fF
C77 a_n118_n140# a_n1364_n140# 0.01fF
C78 a_n118_n140# a_594_n140# 0.01fF
C79 a_n950_n194# a_n238_n194# 0.01fF
C80 a_60_n140# a_950_n140# 0.01fF
C81 a_n1542_n140# a_n474_n140# 0.01fF
C82 a_n950_n194# a_296_n194# 0.01fF
C83 a_n772_n194# a_118_n194# 0.01fF
C84 a_n1364_n140# a_n1720_n140# 0.03fF
C85 a_n2254_n140# a_n652_n140# 0.01fF
C86 a_772_n140# a_1840_n140# 0.01fF
C87 a_n1662_n194# a_n1484_n194# 0.10fF
C88 a_n950_n194# a_n60_n194# 0.01fF
C89 a_830_n194# a_n772_n194# 0.01fF
C90 a_n2432_n140# a_n1720_n140# 0.01fF
C91 a_1720_n194# a_1898_n194# 0.10fF
C92 a_1720_n194# a_296_n194# 0.01fF
C93 a_n474_n140# a_238_n140# 0.01fF
C94 a_1008_n194# a_1720_n194# 0.01fF
C95 a_n1840_n194# a_n238_n194# 0.01fF
C96 a_n2018_n194# a_n416_n194# 0.01fF
C97 a_n1484_n194# a_118_n194# 0.01fF
C98 a_n830_n140# a_n2076_n140# 0.01fF
C99 a_n416_n194# a_n1306_n194# 0.01fF
C100 a_n2254_n140# a_n1720_n140# 0.02fF
C101 a_1840_n140# a_950_n140# 0.01fF
C102 a_n2018_n194# a_n1128_n194# 0.01fF
C103 a_n1186_n140# a_n830_n140# 0.03fF
C104 a_2076_n194# a_2254_n194# 0.06fF
C105 a_n1364_n140# a_n474_n140# 0.01fF
C106 a_594_n140# a_n474_n140# 0.01fF
C107 a_n1128_n194# a_n1306_n194# 0.10fF
C108 a_n830_n140# a_416_n140# 0.01fF
C109 a_60_n140# a_n652_n140# 0.01fF
C110 a_n594_n194# a_652_n194# 0.01fF
C111 a_1484_n140# a_1128_n140# 0.03fF
C112 a_1128_n140# a_238_n140# 0.01fF
C113 a_n118_n140# a_60_n140# 0.06fF
C114 a_n1898_n140# a_n1008_n140# 0.01fF
C115 a_2196_n140# a_1306_n140# 0.01fF
C116 a_n950_n194# a_n416_n194# 0.02fF
C117 a_n830_n140# a_n296_n140# 0.02fF
C118 a_772_n140# a_n830_n140# 0.01fF
C119 a_594_n140# a_1128_n140# 0.02fF
C120 a_1306_n140# a_416_n140# 0.01fF
C121 a_n1128_n194# a_n950_n194# 0.10fF
C122 a_2196_n140# a_2018_n140# 0.06fF
C123 a_n238_n194# a_474_n194# 0.01fF
C124 a_1186_n194# a_118_n194# 0.01fF
C125 a_n2432_n140# a_n1128_n194# 0.00fF
C126 a_2018_n140# a_416_n140# 0.01fF
C127 a_474_n194# a_1898_n194# 0.01fF
C128 a_1186_n194# a_830_n194# 0.03fF
C129 a_1306_n140# a_n296_n140# 0.01fF
C130 a_772_n140# a_1306_n140# 0.02fF
C131 a_1484_n140# a_2254_n194# 0.01fF
C132 a_474_n194# a_296_n194# 0.10fF
C133 a_652_n194# a_118_n194# 0.02fF
C134 a_474_n194# a_n60_n194# 0.02fF
C135 a_n1840_n194# a_n416_n194# 0.01fF
C136 a_60_n140# a_n474_n140# 0.02fF
C137 a_1008_n194# a_474_n194# 0.02fF
C138 a_n2018_n194# a_n1306_n194# 0.01fF
C139 a_1186_n194# a_1364_n194# 0.10fF
C140 a_n1840_n194# a_n1128_n194# 0.01fF
C141 a_n2196_n194# a_n1128_n194# 0.01fF
C142 a_830_n194# a_652_n194# 0.10fF
C143 a_1720_n194# a_2254_n194# 0.01fF
C144 a_772_n140# a_2018_n140# 0.01fF
C145 a_1306_n140# a_950_n140# 0.03fF
C146 a_1720_n194# a_2076_n194# 0.03fF
C147 a_1364_n194# a_652_n194# 0.01fF
C148 a_1542_n194# a_1898_n194# 0.03fF
C149 a_60_n140# a_1128_n140# 0.01fF
C150 a_1542_n194# a_296_n194# 0.01fF
C151 a_n2018_n194# a_n950_n194# 0.01fF
C152 a_n772_n194# a_n1484_n194# 0.01fF
C153 a_n950_n194# a_n1306_n194# 0.03fF
C154 a_1542_n194# a_n60_n194# 0.01fF
C155 a_1542_n194# a_1008_n194# 0.02fF
C156 a_2018_n140# a_950_n140# 0.01fF
C157 a_n830_n140# a_n652_n140# 0.06fF
C158 a_n1542_n140# a_n1364_n140# 0.06fF
C159 a_2196_n140# a_1662_n140# 0.02fF
C160 a_n118_n140# a_n830_n140# 0.01fF
C161 a_n416_n194# a_474_n194# 0.01fF
C162 a_n2432_n140# a_n1542_n140# 0.01fF
C163 a_n2432_n140# a_n2018_n194# 0.02fF
C164 a_n2432_n140# a_n1306_n194# 0.01fF
C165 a_n1128_n194# a_474_n194# 0.01fF
C166 a_1484_n140# a_238_n140# 0.01fF
C167 a_1662_n140# a_416_n140# 0.01fF
C168 a_n830_n140# a_n1720_n140# 0.01fF
C169 a_1128_n140# a_1840_n140# 0.01fF
C170 a_n1542_n140# a_n2254_n140# 0.01fF
C171 a_1484_n140# a_594_n140# 0.01fF
C172 a_594_n140# a_238_n140# 0.03fF
C173 a_n2018_n194# a_n1840_n194# 0.10fF
C174 a_n1364_n140# a_238_n140# 0.01fF
C175 a_n2018_n194# a_n2196_n194# 0.10fF
C176 a_n2076_n140# a_n1008_n140# 0.01fF
C177 a_n118_n140# a_1306_n140# 0.01fF
C178 a_n1840_n194# a_n1306_n194# 0.02fF
C179 a_n2196_n194# a_n1306_n194# 0.01fF
C180 a_n1186_n140# a_n1008_n140# 0.06fF
C181 a_416_n140# a_n1008_n140# 0.01fF
C182 a_772_n140# a_1662_n140# 0.01fF
C183 a_n2432_n140# a_n950_n194# 0.00fF
C184 a_n594_n194# a_n238_n194# 0.03fF
C185 a_n2432_n140# a_n1364_n140# 0.01fF
C186 a_474_n194# a_2076_n194# 0.01fF
C187 a_n830_n140# a_n474_n140# 0.03fF
C188 a_n594_n194# a_296_n194# 0.01fF
C189 a_n2076_n140# a_n1898_n140# 0.06fF
C190 a_n1840_n194# a_n950_n194# 0.01fF
C191 a_n2196_n194# a_n950_n194# 0.01fF
C192 a_652_n194# a_n772_n194# 0.01fF
C193 a_n296_n140# a_n1008_n140# 0.01fF
C194 a_n594_n194# a_n60_n194# 0.02fF
C195 a_n1186_n140# a_n1898_n140# 0.01fF
C196 a_n1542_n140# a_60_n140# 0.01fF
C197 a_n594_n194# a_1008_n194# 0.01fF
C198 a_1662_n140# a_950_n140# 0.01fF
C199 a_2254_n194# a_1840_n140# 0.02fF
C200 a_n2254_n140# a_n1364_n140# 0.01fF
C201 a_n1662_n194# a_n238_n194# 0.01fF
C202 a_1542_n194# a_2254_n194# 0.01fF
C203 a_n2432_n140# a_n1840_n194# 0.01fF
C204 a_n2432_n140# a_n2254_n140# 0.06fF
C205 a_n2432_n140# a_n2196_n194# 0.06fF
C206 a_1542_n194# a_2076_n194# 0.02fF
C207 a_n296_n140# a_n1898_n140# 0.01fF
C208 a_1484_n140# a_60_n140# 0.01fF
C209 a_60_n140# a_238_n140# 0.06fF
C210 a_n1662_n194# a_n60_n194# 0.01fF
C211 a_n238_n194# a_118_n194# 0.03fF
C212 a_n2196_n194# a_n1840_n194# 0.03fF
C213 a_n1364_n140# a_60_n140# 0.01fF
C214 a_830_n194# a_n238_n194# 0.01fF
C215 a_60_n140# a_594_n140# 0.02fF
C216 a_n950_n194# a_474_n194# 0.01fF
C217 a_1306_n140# a_1128_n140# 0.06fF
C218 a_n594_n194# a_n416_n194# 0.10fF
C219 a_296_n194# a_118_n194# 0.10fF
C220 a_830_n194# a_1898_n194# 0.01fF
C221 a_n1128_n194# a_n594_n194# 0.02fF
C222 a_118_n194# a_n60_n194# 0.10fF
C223 a_1008_n194# a_118_n194# 0.01fF
C224 a_830_n194# a_296_n194# 0.02fF
C225 a_1720_n194# a_474_n194# 0.01fF
C226 a_1364_n194# a_n238_n194# 0.01fF
C227 a_830_n194# a_n60_n194# 0.01fF
C228 a_1008_n194# a_830_n194# 0.10fF
C229 a_2018_n140# a_1128_n140# 0.01fF
C230 a_1364_n194# a_1898_n194# 0.02fF
C231 a_1484_n140# a_1840_n140# 0.03fF
C232 a_1840_n140# a_238_n140# 0.01fF
C233 a_1364_n194# a_296_n194# 0.01fF
C234 a_1186_n194# a_652_n194# 0.02fF
C235 a_n652_n140# a_n1008_n140# 0.03fF
C236 a_1364_n194# a_n60_n194# 0.01fF
C237 a_1364_n194# a_1008_n194# 0.03fF
C238 a_n118_n140# a_n1008_n140# 0.01fF
C239 a_n1662_n194# a_n416_n194# 0.01fF
C240 a_594_n140# a_1840_n140# 0.01fF
C241 a_1306_n140# a_2254_n194# 0.01fF
C242 a_n1662_n194# a_n1128_n194# 0.02fF
C243 a_1542_n194# a_1720_n194# 0.10fF
C244 a_n830_n140# a_n1542_n140# 0.01fF
C245 a_n1720_n140# a_n1008_n140# 0.01fF
C246 a_n652_n140# a_n1898_n140# 0.01fF
C247 a_n416_n194# a_118_n194# 0.02fF
C248 a_2018_n140# a_2254_n194# 0.03fF
C249 a_n1128_n194# a_118_n194# 0.01fF
C250 a_830_n194# a_n416_n194# 0.01fF
C251 a_n1186_n140# a_n2076_n140# 0.01fF
C252 a_n2018_n194# a_n594_n194# 0.01fF
C253 a_n594_n194# a_n1306_n194# 0.01fF
C254 a_n1186_n140# a_416_n140# 0.01fF
C255 a_n830_n140# a_238_n140# 0.01fF
C256 a_n1720_n140# a_n1898_n140# 0.06fF
C257 a_n474_n140# a_n1008_n140# 0.02fF
C258 a_1662_n140# a_1128_n140# 0.02fF
C259 a_n772_n194# a_n238_n194# 0.02fF
C260 a_n830_n140# a_594_n140# 0.01fF
C261 a_n830_n140# a_n1364_n140# 0.02fF
C262 a_772_n140# a_2196_n140# 0.01fF
C263 a_n2432_n140# a_n830_n140# 0.01fF
C264 a_830_n194# a_2254_n194# 0.00fF
C265 a_n1186_n140# a_n296_n140# 0.01fF
C266 a_n594_n194# a_n950_n194# 0.03fF
C267 a_416_n140# a_n296_n140# 0.01fF
C268 a_1306_n140# a_1484_n140# 0.06fF
C269 a_1306_n140# a_238_n140# 0.01fF
C270 a_772_n140# a_416_n140# 0.03fF
C271 a_n772_n194# a_296_n194# 0.01fF
C272 a_n2018_n194# a_n1662_n194# 0.03fF
C273 a_830_n194# a_2076_n194# 0.01fF
C274 a_n1662_n194# a_n1306_n194# 0.03fF
C275 a_n772_n194# a_n60_n194# 0.01fF
C276 a_n474_n140# a_n1898_n140# 0.01fF
C277 a_1364_n194# a_2254_n194# 0.01fF
C278 a_n238_n194# a_n1484_n194# 0.01fF
C279 a_1306_n140# a_594_n140# 0.01fF
C280 a_n830_n140# a_n2254_n140# 0.01fF
C281 a_2196_n140# a_950_n140# 0.01fF
C282 a_1542_n194# a_474_n194# 0.01fF
C283 a_1484_n140# a_2018_n140# 0.02fF
C284 a_1364_n194# a_2076_n194# 0.01fF
C285 a_772_n140# a_n296_n140# 0.01fF
C286 a_n1306_n194# a_118_n194# 0.01fF
C287 a_1662_n140# a_2254_n194# 0.01fF
C288 a_416_n140# a_950_n140# 0.02fF
C289 a_n1662_n194# a_n950_n194# 0.01fF
C290 a_n1484_n194# a_n60_n194# 0.01fF
C291 a_2018_n140# a_594_n140# 0.01fF
C292 a_n1840_n194# a_n594_n194# 0.01fF
C293 a_n2196_n194# a_n594_n194# 0.01fF
C294 a_950_n140# a_n296_n140# 0.01fF
C295 a_n830_n140# a_60_n140# 0.01fF
C296 a_n2432_n140# a_n1662_n194# 0.01fF
C297 a_772_n140# a_950_n140# 0.06fF
C298 a_n950_n194# a_118_n194# 0.01fF
C299 a_n772_n194# a_n416_n194# 0.03fF
C300 a_n1128_n194# a_n772_n194# 0.03fF
C301 a_1186_n194# a_n238_n194# 0.01fF
C302 a_1720_n194# a_118_n194# 0.01fF
C303 a_n2076_n140# a_n652_n140# 0.01fF
C304 a_n1662_n194# a_n1840_n194# 0.10fF
C305 a_n2196_n194# a_n1662_n194# 0.02fF
C306 a_1186_n194# a_1898_n194# 0.01fF
C307 a_n1186_n140# a_n652_n140# 0.02fF
C308 a_830_n194# a_1720_n194# 0.01fF
C309 a_416_n140# a_n652_n140# 0.01fF
C310 a_1306_n140# a_60_n140# 0.01fF
C311 a_1186_n194# a_296_n194# 0.01fF
C312 a_652_n194# a_n238_n194# 0.01fF
C313 a_n118_n140# a_n1186_n140# 0.01fF
C314 a_n416_n194# a_n1484_n194# 0.01fF
C315 a_1186_n194# a_n60_n194# 0.01fF
C316 a_n118_n140# a_416_n140# 0.02fF
C317 a_1186_n194# a_1008_n194# 0.10fF
C318 a_n594_n194# a_474_n194# 0.01fF
C319 a_n1542_n140# a_n1008_n140# 0.02fF
C320 a_n1128_n194# a_n1484_n194# 0.03fF
C321 a_1662_n140# a_1484_n140# 0.06fF
C322 a_652_n194# a_1898_n194# 0.01fF
C323 a_1662_n140# a_238_n140# 0.01fF
C324 a_1364_n194# a_1720_n194# 0.03fF
C325 a_652_n194# a_296_n194# 0.03fF
C326 a_n2076_n140# a_n1720_n140# 0.03fF
C327 a_n652_n140# a_n296_n140# 0.03fF
C328 a_n1186_n140# a_n1720_n140# 0.02fF
C329 a_772_n140# a_n652_n140# 0.01fF
C330 a_652_n194# a_n60_n194# 0.01fF
C331 a_1008_n194# a_652_n194# 0.03fF
C332 a_1662_n140# a_594_n140# 0.01fF
C333 a_n118_n140# a_n296_n140# 0.06fF
C334 a_n118_n140# a_772_n140# 0.01fF
C335 a_n1542_n140# a_n1898_n140# 0.03fF
C336 a_238_n140# a_n1008_n140# 0.01fF
C337 a_1306_n140# a_1840_n140# 0.02fF
C338 a_n2076_n140# a_n474_n140# 0.01fF
C339 a_n1720_n140# a_n296_n140# 0.01fF
C340 a_n652_n140# a_950_n140# 0.01fF
C341 a_n2018_n194# a_n772_n194# 0.01fF
C342 a_594_n140# a_n1008_n140# 0.01fF
C343 a_n1364_n140# a_n1008_n140# 0.03fF
C344 a_n772_n194# a_n1306_n194# 0.02fF
C345 a_1186_n194# a_n416_n194# 0.01fF
C346 a_n1186_n140# a_n474_n140# 0.01fF
C347 a_n118_n140# a_950_n140# 0.01fF
C348 a_416_n140# a_n474_n140# 0.01fF
C349 a_n2432_n140# a_n1008_n140# 0.01fF
C350 a_2018_n140# a_1840_n140# 0.06fF
C351 a_474_n194# a_118_n194# 0.03fF
C352 a_830_n194# a_474_n194# 0.03fF
C353 a_2196_n140# a_1128_n140# 0.01fF
C354 a_652_n194# a_n416_n194# 0.01fF
C355 a_n2018_n194# a_n1484_n194# 0.02fF
C356 a_n1364_n140# a_n1898_n140# 0.02fF
C357 a_n1306_n194# a_n1484_n194# 0.10fF
C358 a_n2254_n140# a_n1008_n140# 0.01fF
C359 a_n474_n140# a_n296_n140# 0.06fF
C360 a_772_n140# a_n474_n140# 0.01fF
C361 a_n772_n194# a_n950_n194# 0.10fF
C362 a_416_n140# a_1128_n140# 0.01fF
C363 a_n2432_n140# a_n1898_n140# 0.02fF
C364 a_1364_n194# a_474_n194# 0.01fF
C365 a_1662_n140# a_60_n140# 0.01fF
C366 a_1186_n194# a_2254_n194# 0.01fF
C367 a_n2432_n140# a_n772_n194# 0.00fF
C368 a_1186_n194# a_2076_n194# 0.01fF
C369 a_1542_n194# a_118_n194# 0.01fF
C370 a_n2254_n140# a_n1898_n140# 0.03fF
C371 a_n950_n194# a_n1484_n194# 0.02fF
C372 a_n118_n140# a_n652_n140# 0.02fF
C373 a_n474_n140# a_950_n140# 0.01fF
C374 a_1128_n140# a_n296_n140# 0.01fF
C375 a_772_n140# a_1128_n140# 0.03fF
C376 a_1542_n194# a_830_n194# 0.01fF
C377 a_652_n194# a_2254_n194# 0.00fF
C378 a_60_n140# a_n1008_n140# 0.01fF
C379 a_2196_n140# a_2254_n194# 0.06fF
C380 a_652_n194# a_2076_n194# 0.01fF
C381 a_n1840_n194# a_n772_n194# 0.01fF
C382 a_n2196_n194# a_n772_n194# 0.01fF
C383 a_1364_n194# a_1542_n194# 0.10fF
C384 a_n2432_n140# a_n1484_n194# 0.01fF
C385 a_n1720_n140# a_n652_n140# 0.01fF
C386 a_1662_n140# a_1840_n140# 0.06fF
C387 a_1128_n140# a_950_n140# 0.06fF
C388 a_n118_n140# a_n1720_n140# 0.01fF
C389 a_1306_n140# a_2018_n140# 0.01fF
C390 a_n1840_n194# a_n1484_n194# 0.03fF
C391 a_n2196_n194# a_n1484_n194# 0.01fF
C392 a_n1662_n194# a_n594_n194# 0.01fF
C393 a_772_n140# a_2254_n194# 0.01fF
C394 a_n1542_n140# a_n2076_n140# 0.02fF
C395 a_n652_n140# a_n474_n140# 0.06fF
C396 a_n238_n194# a_296_n194# 0.02fF
C397 a_n1186_n140# a_n1542_n140# 0.03fF
C398 a_n238_n194# a_n60_n194# 0.10fF
C399 a_n118_n140# a_n474_n140# 0.03fF
C400 a_1008_n194# a_n238_n194# 0.01fF
C401 a_n772_n194# a_474_n194# 0.01fF
C402 a_1898_n194# a_296_n194# 0.01fF
C403 a_n594_n194# a_118_n194# 0.01fF
C404 a_1186_n194# a_1720_n194# 0.02fF
C405 a_2196_n140# VSUBS 0.01fF
C406 a_2018_n140# VSUBS 0.01fF
C407 a_1840_n140# VSUBS 0.02fF
C408 a_1662_n140# VSUBS 0.02fF
C409 a_1484_n140# VSUBS 0.02fF
C410 a_1306_n140# VSUBS 0.02fF
C411 a_1128_n140# VSUBS 0.02fF
C412 a_950_n140# VSUBS 0.02fF
C413 a_772_n140# VSUBS 0.02fF
C414 a_594_n140# VSUBS 0.02fF
C415 a_416_n140# VSUBS 0.02fF
C416 a_238_n140# VSUBS 0.02fF
C417 a_60_n140# VSUBS 0.02fF
C418 a_n118_n140# VSUBS 0.02fF
C419 a_n296_n140# VSUBS 0.02fF
C420 a_n474_n140# VSUBS 0.02fF
C421 a_n652_n140# VSUBS 0.02fF
C422 a_n830_n140# VSUBS 0.02fF
C423 a_n1008_n140# VSUBS 0.02fF
C424 a_n1186_n140# VSUBS 0.02fF
C425 a_n1364_n140# VSUBS 0.02fF
C426 a_n1542_n140# VSUBS 0.02fF
C427 a_n1720_n140# VSUBS 0.02fF
C428 a_n1898_n140# VSUBS 0.02fF
C429 a_n2076_n140# VSUBS 0.02fF
C430 a_n2254_n140# VSUBS 0.02fF
C431 a_2254_n194# VSUBS 0.31fF
C432 a_2076_n194# VSUBS 0.19fF
C433 a_1898_n194# VSUBS 0.20fF
C434 a_1720_n194# VSUBS 0.21fF
C435 a_1542_n194# VSUBS 0.22fF
C436 a_1364_n194# VSUBS 0.23fF
C437 a_1186_n194# VSUBS 0.23fF
C438 a_1008_n194# VSUBS 0.24fF
C439 a_830_n194# VSUBS 0.24fF
C440 a_652_n194# VSUBS 0.24fF
C441 a_474_n194# VSUBS 0.24fF
C442 a_296_n194# VSUBS 0.24fF
C443 a_118_n194# VSUBS 0.24fF
C444 a_n60_n194# VSUBS 0.24fF
C445 a_n238_n194# VSUBS 0.24fF
C446 a_n416_n194# VSUBS 0.24fF
C447 a_n594_n194# VSUBS 0.24fF
C448 a_n772_n194# VSUBS 0.24fF
C449 a_n950_n194# VSUBS 0.24fF
C450 a_n1128_n194# VSUBS 0.24fF
C451 a_n1306_n194# VSUBS 0.24fF
C452 a_n1484_n194# VSUBS 0.24fF
C453 a_n1662_n194# VSUBS 0.24fF
C454 a_n1840_n194# VSUBS 0.24fF
C455 a_n2018_n194# VSUBS 0.24fF
C456 a_n2196_n194# VSUBS 0.24fF
C457 a_n2432_n140# VSUBS 0.36fF
.ends

.subckt bias_circuit bias_c bias_e i_bias VDD m1_1243_5997# m1_3443_5997# bias_a m1_7347_1428#
+ m1_7639_1420# m1_7169_923# m1_7461_921# m1_7639_427# m1_7347_423# bias_b VSS m1_3551_3596#
+ m1_5643_5997# bias_d
Xsky130_fd_pr__nfet_01v8_6RUDQZ_0 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_1 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_2 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_3 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_SD55Q9_0 m1_7347_1428# m1_7639_1420# bias_e m1_7055_1417#
+ bias_e m1_6763_422# bias_e m1_6471_422# bias_e VSS VSS VSS m1_7639_427# m1_7347_423#
+ m1_7055_433# bias_e bias_e bias_e m1_6763_422# m1_6471_422# m1_7169_923# bias_e
+ m1_7461_921# bias_e bias_e m1_7639_427# m1_7347_423# m1_6877_922# m1_7055_433# VSS
+ bias_e VSS VSS bias_e bias_e bias_e m1_6877_922# m1_6585_923# VSS bias_e m1_6763_1422#
+ m1_6293_922# bias_e m1_6471_1426# m1_7347_1428# bias_e bias_e m1_7639_1420# m1_7169_923#
+ m1_7055_1417# bias_e bias_e m1_7461_921# bias_e bias_e bias_e m1_6585_923# bias_e
+ m1_6293_922# m1_6763_1422# bias_e m1_6471_1426# VSS sky130_fd_pr__nfet_01v8_SD55Q9
Xsky130_fd_pr__nfet_01v8_EZNTQN_0 bias_c VSS VSS i_bias i_bias i_bias i_bias VSS VSS
+ bias_c VSS VSS i_bias VSS bias_c i_bias i_bias i_bias i_bias VSS i_bias i_bias bias_c
+ i_bias VSS VSS i_bias i_bias i_bias bias_c VSS VSS i_bias bias_c VSS i_bias i_bias
+ VSS i_bias i_bias i_bias i_bias i_bias VSS i_bias i_bias i_bias i_bias i_bias i_bias
+ i_bias bias_c i_bias VSS i_bias i_bias bias_c i_bias i_bias i_bias i_bias VSS i_bias
+ VSS i_bias VSS VSS i_bias i_bias bias_c i_bias VSS i_bias i_bias i_bias i_bias bias_c
+ sky130_fd_pr__nfet_01v8_EZNTQN
Xsky130_fd_pr__pfet_01v8_JJWXCM_0 bias_b bias_c m1_1243_5997# m1_1243_5997# bias_b
+ bias_c VDD VDD bias_c bias_b bias_c VDD bias_c m1_1243_5997# bias_c bias_b VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_1 m1_3551_3596# bias_c m1_3443_5997# m1_3443_5997#
+ m1_3551_3596# bias_c VDD VDD bias_c m1_3551_3596# bias_c VDD bias_c m1_3443_5997#
+ bias_c m1_3551_3596# VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_2 bias_e bias_c m1_5643_5997# m1_5643_5997# bias_e
+ bias_c VDD VDD bias_c bias_e bias_c VDD bias_c m1_5643_5997# bias_c bias_e VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__nfet_01v8_LJREPQ_0 m1_3551_3596# bias_d VSS bias_a bias_d m1_3551_3596#
+ VSS VSS sky130_fd_pr__nfet_01v8_LJREPQ
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_0 m1_1243_5997# bias_b VDD VDD m1_1243_5997# bias_b
+ VDD VDD bias_b m1_1243_5997# bias_b VDD bias_b VDD bias_b m1_1243_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_1 m1_3443_5997# bias_b VDD VDD m1_3443_5997# bias_b
+ VDD VDD bias_b m1_3443_5997# bias_b VDD bias_b VDD bias_b m1_3443_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_2 m1_5643_5997# bias_b VDD VDD m1_5643_5997# bias_b
+ VDD VDD bias_b m1_5643_5997# bias_b VDD bias_b VDD bias_b m1_5643_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__nfet_01v8_lvt_28TRYY_0 bias_b bias_c bias_b bias_b bias_b bias_c bias_b
+ bias_b VSS bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_c bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_c bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_c bias_b bias_c bias_b bias_b bias_b
+ bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_c
+ bias_c bias_b bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_c
+ bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_c bias_c bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b
+ bias_b bias_b sky130_fd_pr__nfet_01v8_lvt_28TRYY
Xsky130_fd_pr__nfet_01v8_EL6FQZ_0 bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d VSS m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
Xsky130_fd_pr__nfet_01v8_EL6FQZ_1 bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d VSS m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
C0 i_bias bias_a 0.02fF
C1 m1_7639_427# bias_a 0.01fF
C2 m1_6763_1422# bias_d 0.00fF
C3 m1_7639_1420# bias_d 0.00fF
C4 m1_7055_1417# bias_a 0.00fF
C5 bias_e m1_7055_433# 0.26fF
C6 li_3433_399# m1_6471_1426# 0.01fF
C7 bias_e m1_7347_1428# 0.32fF
C8 m1_3551_3596# bias_a 0.26fF
C9 bias_e m1_6763_422# 0.26fF
C10 m1_6877_922# bias_a 0.00fF
C11 i_bias bias_d 0.00fF
C12 m1_6877_922# m1_7461_921# 0.01fF
C13 bias_c bias_a 0.02fF
C14 m1_3443_5997# bias_e 0.02fF
C15 m1_7055_433# m1_6471_422# 0.01fF
C16 m1_3443_5997# bias_b 0.65fF
C17 m1_6293_922# m1_6877_922# 0.01fF
C18 m1_7055_1417# bias_d 0.00fF
C19 m1_6877_922# m1_6585_923# 0.03fF
C20 bias_d VDD 0.07fF
C21 m1_7347_1428# m1_6763_1422# 0.01fF
C22 m1_7347_1428# m1_7639_1420# 0.03fF
C23 li_3433_399# bias_a 7.53fF
C24 bias_a m1_7347_423# 0.01fF
C25 m1_6763_1422# m1_6763_422# -0.00fF
C26 m1_5643_5997# bias_d 0.03fF
C27 m1_6763_422# m1_6471_422# 0.03fF
C28 m1_3551_3596# bias_d 18.83fF
C29 m1_6293_922# li_3433_399# 0.02fF
C30 li_3433_399# m1_6585_923# 0.01fF
C31 bias_a m1_6471_1426# 0.01fF
C32 bias_c bias_d 0.90fF
C33 m1_7639_427# m1_7055_433# 0.01fF
C34 m1_7055_1417# m1_7055_433# -0.00fF
C35 bias_e bias_b 0.07fF
C36 li_3433_399# bias_d 5.36fF
C37 m1_7347_1428# m1_7055_1417# 0.03fF
C38 m1_7639_427# m1_6763_422# 0.01fF
C39 bias_d m1_6471_1426# 0.01fF
C40 bias_a m1_7461_921# 0.00fF
C41 bias_e m1_7169_923# 0.22fF
C42 bias_e m1_6763_1422# 0.33fF
C43 bias_e m1_6471_422# 0.25fF
C44 bias_e m1_7639_1420# 0.18fF
C45 m1_3443_5997# VDD 0.84fF
C46 m1_6293_922# bias_a 0.01fF
C47 m1_6293_922# m1_7461_921# 0.01fF
C48 bias_a m1_6585_923# 0.00fF
C49 m1_6585_923# m1_7461_921# 0.01fF
C50 m1_3443_5997# m1_5643_5997# 0.11fF
C51 m1_3443_5997# m1_3551_3596# 0.98fF
C52 m1_3443_5997# m1_1243_5997# 0.07fF
C53 m1_7347_423# m1_7055_433# 0.03fF
C54 m1_6293_922# m1_6585_923# 0.03fF
C55 m1_3443_5997# bias_c 0.44fF
C56 m1_7347_1428# m1_7347_423# -0.00fF
C57 bias_e m1_7639_427# 0.18fF
C58 m1_7639_1420# m1_6763_1422# 0.01fF
C59 bias_a bias_d 7.33fF
C60 i_bias bias_b 0.60fF
C61 m1_6763_422# m1_7347_423# 0.01fF
C62 m1_7347_1428# m1_6471_1426# 0.01fF
C63 bias_e m1_7055_1417# 0.33fF
C64 bias_e VDD 0.26fF
C65 m1_6293_922# bias_d 0.00fF
C66 bias_d m1_6585_923# 0.00fF
C67 bias_b VDD 8.29fF
C68 m1_5643_5997# bias_e 0.71fF
C69 bias_e m1_3551_3596# 0.76fF
C70 m1_5643_5997# bias_b 0.63fF
C71 bias_e m1_6877_922# 0.22fF
C72 m1_3551_3596# bias_b 0.71fF
C73 m1_1243_5997# bias_b 0.77fF
C74 m1_7639_427# m1_6471_422# 0.01fF
C75 m1_7639_1420# m1_7639_427# -0.00fF
C76 bias_c bias_e 0.65fF
C77 bias_a m1_7055_433# 0.01fF
C78 m1_6763_1422# m1_7055_1417# 0.03fF
C79 bias_c bias_b 22.44fF
C80 m1_7639_1420# m1_7055_1417# 0.01fF
C81 m1_7347_1428# bias_a 0.00fF
C82 bias_e li_3433_399# 0.02fF
C83 m1_6763_422# bias_a 0.01fF
C84 bias_e m1_7347_423# 0.26fF
C85 m1_6877_922# m1_7169_923# 0.03fF
C86 bias_e m1_6471_1426# 0.34fF
C87 m1_7347_1428# bias_d 0.00fF
C88 li_3433_399# m1_6471_422# 0.01fF
C89 m1_7347_423# m1_6471_422# 0.01fF
C90 bias_c i_bias 5.62fF
C91 m1_5643_5997# VDD 1.16fF
C92 m1_3551_3596# VDD 0.64fF
C93 m1_1243_5997# VDD 1.50fF
C94 m1_6763_1422# m1_6471_1426# 0.03fF
C95 m1_6471_1426# m1_6471_422# -0.00fF
C96 m1_7639_1420# m1_6471_1426# 0.01fF
C97 m1_3443_5997# bias_d 0.03fF
C98 bias_e bias_a 0.24fF
C99 bias_e m1_7461_921# 0.21fF
C100 i_bias li_3433_399# 0.03fF
C101 bias_c VDD 4.90fF
C102 m1_5643_5997# m1_3551_3596# 0.08fF
C103 m1_1243_5997# m1_3551_3596# 0.03fF
C104 m1_7639_427# m1_7347_423# 0.03fF
C105 m1_6293_922# bias_e 0.18fF
C106 bias_e m1_6585_923# 0.22fF
C107 bias_c m1_5643_5997# 0.44fF
C108 bias_c m1_3551_3596# 2.13fF
C109 bias_c m1_1243_5997# 0.52fF
C110 m1_6763_422# m1_7055_433# 0.03fF
C111 m1_3551_3596# li_3433_399# 0.03fF
C112 bias_a m1_7169_923# 0.00fF
C113 m1_6763_1422# bias_a 0.00fF
C114 bias_a m1_6471_422# 0.01fF
C115 m1_7461_921# m1_7169_923# 0.03fF
C116 m1_7639_1420# bias_a 0.00fF
C117 m1_7055_1417# m1_6471_1426# 0.01fF
C118 bias_e bias_d 0.26fF
C119 bias_d bias_b 0.26fF
C120 m1_6293_922# m1_7169_923# 0.01fF
C121 m1_6585_923# m1_7169_923# 0.01fF
C122 m1_3551_3596# VSS -340.53fF
C123 bias_b VSS -284.38fF
C124 m1_5643_5997# VSS 38.06fF
C125 m1_3443_5997# VSS 35.86fF
C126 m1_1243_5997# VSS 25.05fF
C127 VDD VSS 131.75fF
C128 i_bias VSS -59.70fF
C129 bias_c VSS -50.79fF
C130 m1_7639_427# VSS 0.32fF
C131 m1_7347_423# VSS 0.26fF
C132 m1_7461_921# VSS 0.22fF
C133 m1_7169_923# VSS 0.19fF
C134 m1_7055_433# VSS 0.28fF
C135 m1_6763_422# VSS 0.34fF
C136 m1_6471_422# VSS 0.38fF
C137 m1_7639_1420# VSS 0.30fF
C138 m1_7347_1428# VSS 0.20fF
C139 m1_6877_922# VSS 0.21fF
C140 m1_6585_923# VSS 0.29fF
C141 m1_6293_922# VSS 0.32fF
C142 m1_7055_1417# VSS 0.19fF
C143 m1_6763_1422# VSS 0.28fF
C144 m1_6471_1426# VSS 0.29fF
C145 bias_e VSS 7.82fF
C146 bias_d VSS -76.92fF
C147 li_3433_399# VSS 5.57fF
C148 bias_a VSS -48.11fF
.ends

.subckt sky130_fd_pr__pfet_01v8_YVTMSC a_n207_n140# a_29_n205# a_327_n140# a_n683_n205#
+ a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_n505_n205# a_n741_n140# a_563_n205#
+ a_861_n140# a_919_n205# a_n327_n205# a_n563_n140# a_385_n205# a_683_n140# w_n1133_n241#
+ a_n919_n140# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n385_n140# a_n505_n205# a_n563_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n205# a_149_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n205# a_n29_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_861_n140# a_741_n205# a_683_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n205# a_n385_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n741_n140# a_n861_n205# a_n919_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_683_n140# a_563_n205# a_505_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_919_n205# a_919_n205# a_861_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_n29_n140# a_n149_n205# a_n207_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n563_n140# a_n683_n205# a_n741_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_n919_n140# a_n1097_n140# a_n1097_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_505_n140# a_385_n205# a_327_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1097_n140# a_385_n205# 0.00fF
C1 a_683_n140# a_n385_n140# 0.01fF
C2 a_683_n140# a_n563_n140# 0.01fF
C3 a_505_n140# a_683_n140# 0.06fF
C4 a_n741_n140# w_n1133_n241# 0.02fF
C5 a_207_n205# a_n683_n205# 0.01fF
C6 a_n207_n140# a_n919_n140# 0.01fF
C7 a_n1097_n140# a_149_n140# 0.01fF
C8 a_29_n205# a_n683_n205# 0.01fF
C9 a_n149_n205# a_385_n205# 0.02fF
C10 a_n1097_n140# a_n505_n205# 0.01fF
C11 a_385_n205# w_n1133_n241# 0.16fF
C12 a_683_n140# a_n29_n140# 0.01fF
C13 a_207_n205# a_741_n205# 0.02fF
C14 a_n327_n205# a_207_n205# 0.02fF
C15 w_n1133_n241# a_149_n140# 0.02fF
C16 a_29_n205# a_741_n205# 0.01fF
C17 a_n149_n205# a_n505_n205# 0.03fF
C18 a_n327_n205# a_29_n205# 0.03fF
C19 a_683_n140# a_327_n140# 0.03fF
C20 a_207_n205# a_563_n205# 0.03fF
C21 w_n1133_n241# a_n505_n205# 0.20fF
C22 a_29_n205# a_563_n205# 0.02fF
C23 a_207_n205# a_n861_n205# 0.01fF
C24 a_29_n205# a_n861_n205# 0.01fF
C25 a_n149_n205# a_919_n205# 0.01fF
C26 a_683_n140# a_n207_n140# 0.01fF
C27 a_n1097_n140# a_n683_n205# 0.02fF
C28 w_n1133_n241# a_861_n140# 0.01fF
C29 w_n1133_n241# a_919_n205# 0.28fF
C30 a_n1097_n140# a_n385_n140# 0.01fF
C31 a_n741_n140# a_149_n140# 0.01fF
C32 a_683_n140# a_n919_n140# 0.01fF
C33 a_n1097_n140# a_n563_n140# 0.02fF
C34 a_505_n140# a_n1097_n140# 0.01fF
C35 a_n149_n205# a_n683_n205# 0.02fF
C36 a_n683_n205# w_n1133_n241# 0.20fF
C37 a_n327_n205# a_n1097_n140# 0.01fF
C38 a_n741_n140# a_861_n140# 0.01fF
C39 a_385_n205# a_n505_n205# 0.01fF
C40 w_n1133_n241# a_n385_n140# 0.02fF
C41 a_n563_n140# w_n1133_n241# 0.02fF
C42 a_505_n140# w_n1133_n241# 0.02fF
C43 a_n1097_n140# a_n29_n140# 0.01fF
C44 a_n1097_n140# a_563_n205# 0.00fF
C45 a_n1097_n140# a_n861_n205# 0.07fF
C46 a_n149_n205# a_741_n205# 0.01fF
C47 a_n327_n205# a_n149_n205# 0.10fF
C48 a_385_n205# a_919_n205# 0.01fF
C49 a_n1097_n140# a_327_n140# 0.01fF
C50 a_741_n205# w_n1133_n241# 0.14fF
C51 a_n327_n205# w_n1133_n241# 0.19fF
C52 a_563_n205# a_n149_n205# 0.01fF
C53 a_149_n140# a_861_n140# 0.01fF
C54 a_n29_n140# w_n1133_n241# 0.02fF
C55 a_n741_n140# a_n385_n140# 0.03fF
C56 a_563_n205# w_n1133_n241# 0.15fF
C57 a_n149_n205# a_n861_n205# 0.01fF
C58 a_n741_n140# a_n563_n140# 0.06fF
C59 a_919_n205# a_149_n140# 0.01fF
C60 a_505_n140# a_n741_n140# 0.01fF
C61 a_n1097_n140# a_n207_n140# 0.01fF
C62 a_n683_n205# a_385_n205# 0.01fF
C63 a_n861_n205# w_n1133_n241# 0.20fF
C64 a_n505_n205# a_919_n205# 0.00fF
C65 a_n1097_n140# a_n919_n140# 0.06fF
C66 a_327_n140# w_n1133_n241# 0.02fF
C67 a_919_n205# a_861_n140# 0.06fF
C68 a_n741_n140# a_n29_n140# 0.01fF
C69 a_n207_n140# w_n1133_n241# 0.02fF
C70 a_29_n205# a_207_n205# 0.10fF
C71 a_n385_n140# a_149_n140# 0.02fF
C72 a_n563_n140# a_149_n140# 0.01fF
C73 a_505_n140# a_149_n140# 0.03fF
C74 a_n683_n205# a_n505_n205# 0.10fF
C75 a_741_n205# a_385_n205# 0.03fF
C76 a_n327_n205# a_385_n205# 0.01fF
C77 w_n1133_n241# a_n919_n140# 0.02fF
C78 a_n741_n140# a_327_n140# 0.01fF
C79 a_563_n205# a_385_n205# 0.10fF
C80 a_n683_n205# a_919_n205# 0.00fF
C81 a_n861_n205# a_385_n205# 0.01fF
C82 a_n385_n140# a_861_n140# 0.01fF
C83 a_n563_n140# a_861_n140# 0.01fF
C84 a_505_n140# a_861_n140# 0.03fF
C85 a_n385_n140# a_919_n205# 0.01fF
C86 a_n563_n140# a_919_n205# 0.01fF
C87 a_505_n140# a_919_n205# 0.02fF
C88 a_n741_n140# a_n207_n140# 0.02fF
C89 a_n29_n140# a_149_n140# 0.06fF
C90 a_741_n205# a_n505_n205# 0.01fF
C91 a_n327_n205# a_n505_n205# 0.10fF
C92 a_n741_n140# a_n919_n140# 0.06fF
C93 a_563_n205# a_n505_n205# 0.01fF
C94 a_327_n140# a_149_n140# 0.06fF
C95 a_741_n205# a_919_n205# 0.07fF
C96 a_207_n205# a_n1097_n140# 0.00fF
C97 a_n861_n205# a_n505_n205# 0.03fF
C98 a_n327_n205# a_919_n205# 0.00fF
C99 a_29_n205# a_n1097_n140# 0.01fF
C100 a_n29_n140# a_861_n140# 0.01fF
C101 a_n29_n140# a_919_n205# 0.01fF
C102 a_563_n205# a_919_n205# 0.02fF
C103 a_n563_n140# a_n385_n140# 0.06fF
C104 a_683_n140# w_n1133_n241# 0.01fF
C105 a_505_n140# a_n385_n140# 0.01fF
C106 a_505_n140# a_n563_n140# 0.01fF
C107 a_n207_n140# a_149_n140# 0.03fF
C108 a_327_n140# a_861_n140# 0.02fF
C109 a_207_n205# a_n149_n205# 0.03fF
C110 a_741_n205# a_n683_n205# 0.01fF
C111 a_327_n140# a_919_n205# 0.01fF
C112 a_149_n140# a_n919_n140# 0.01fF
C113 a_n327_n205# a_n683_n205# 0.03fF
C114 a_29_n205# a_n149_n205# 0.10fF
C115 a_207_n205# w_n1133_n241# 0.17fF
C116 a_563_n205# a_n683_n205# 0.01fF
C117 a_29_n205# w_n1133_n241# 0.18fF
C118 a_n207_n140# a_861_n140# 0.01fF
C119 a_n29_n140# a_n385_n140# 0.03fF
C120 a_n207_n140# a_919_n205# 0.01fF
C121 a_n861_n205# a_n683_n205# 0.10fF
C122 a_n563_n140# a_n29_n140# 0.02fF
C123 a_683_n140# a_n741_n140# 0.01fF
C124 a_505_n140# a_n29_n140# 0.02fF
C125 a_n327_n205# a_741_n205# 0.01fF
C126 a_327_n140# a_n385_n140# 0.01fF
C127 a_n563_n140# a_327_n140# 0.01fF
C128 a_505_n140# a_327_n140# 0.06fF
C129 a_563_n205# a_741_n205# 0.10fF
C130 a_n327_n205# a_563_n205# 0.01fF
C131 a_741_n205# a_n861_n205# 0.01fF
C132 a_n207_n140# a_n385_n140# 0.06fF
C133 a_n327_n205# a_n861_n205# 0.02fF
C134 a_n563_n140# a_n207_n140# 0.03fF
C135 a_505_n140# a_n207_n140# 0.01fF
C136 a_683_n140# a_149_n140# 0.02fF
C137 a_207_n205# a_385_n205# 0.10fF
C138 a_n1097_n140# a_n149_n205# 0.01fF
C139 a_29_n205# a_385_n205# 0.03fF
C140 a_563_n205# a_n861_n205# 0.01fF
C141 a_n385_n140# a_n919_n140# 0.02fF
C142 a_n1097_n140# w_n1133_n241# 0.33fF
C143 a_n563_n140# a_n919_n140# 0.03fF
C144 a_505_n140# a_n919_n140# 0.01fF
C145 a_n29_n140# a_327_n140# 0.03fF
C146 a_683_n140# a_861_n140# 0.06fF
C147 a_683_n140# a_919_n205# 0.03fF
C148 a_207_n205# a_n505_n205# 0.01fF
C149 a_n207_n140# a_n29_n140# 0.06fF
C150 a_n149_n205# w_n1133_n241# 0.19fF
C151 a_29_n205# a_n505_n205# 0.02fF
C152 a_n29_n140# a_n919_n140# 0.01fF
C153 a_n1097_n140# a_n741_n140# 0.03fF
C154 a_n207_n140# a_327_n140# 0.02fF
C155 a_207_n205# a_919_n205# 0.01fF
C156 a_29_n205# a_919_n205# 0.01fF
C157 a_327_n140# a_n919_n140# 0.01fF
C158 w_n1133_n241# VSUBS 3.28fF
.ends

.subckt ota_v2_without_cmfb in bias_c bias_e op on i_bias VDD bias_d VSS bias_circuit_0/m1_3551_3596#
+ li_11121_570# li_11122_5650# cmc li_14138_570# li_8434_570# li_8436_5651# bias_b
+ bias_circuit_0/m1_1243_5997# bias_circuit_0/m1_3443_5997# bias_a ip bias_circuit_0/m1_5643_5997#
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_0 VDD bias_b bias_b li_8436_5651# bias_b VDD bias_b
+ li_8436_5651# VDD li_8436_5651# VDD bias_b li_8436_5651# bias_b VDD VDD bias_b bias_b
+ VDD bias_b li_8436_5651# VDD bias_b li_8436_5651# li_8436_5651# bias_b VDD bias_b
+ VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_8 bias_d li_8434_570# bias_d on VSS bias_d on li_8434_570#
+ on bias_d bias_d bias_d on bias_d li_8434_570# VSS li_8434_570# bias_d bias_d on
+ li_8434_570# bias_d on on bias_d bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_1 VDD bias_b bias_b li_11122_5650# bias_b VDD
+ bias_b li_11122_5650# VDD li_11122_5650# VDD bias_b li_11122_5650# bias_b VDD VDD
+ bias_b bias_b VDD bias_b li_11122_5650# VDD bias_b li_11122_5650# li_11122_5650#
+ bias_b VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_9 bias_d li_11121_570# bias_d op VSS bias_d op li_11121_570#
+ op bias_d bias_d bias_d op bias_d li_11121_570# VSS li_11121_570# bias_d bias_d
+ op li_11121_570# bias_d op op bias_d bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_2 VDD bias_b bias_b li_8436_5651# bias_b VDD bias_b
+ li_8436_5651# VDD li_8436_5651# VDD bias_b li_8436_5651# bias_b VDD VDD bias_b bias_b
+ VDD bias_b li_8436_5651# VDD bias_b li_8436_5651# li_8436_5651# bias_b VDD bias_b
+ VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_3 VDD bias_b bias_b li_11122_5650# bias_b VDD
+ bias_b li_11122_5650# VDD li_11122_5650# VDD bias_b li_11122_5650# bias_b VDD VDD
+ bias_b bias_b VDD bias_b li_11122_5650# VDD bias_b li_11122_5650# li_11122_5650#
+ bias_b VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_0 VSS li_8436_5651# li_14138_570# ip li_8436_5651#
+ li_8436_5651# ip li_14138_570# li_8436_5651# li_14138_570# li_14138_570# li_8436_5651#
+ li_8436_5651# ip ip li_14138_570# ip li_14138_570# ip VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_1 VSS li_11122_5650# li_14138_570# in li_11122_5650#
+ li_11122_5650# in li_14138_570# li_11122_5650# li_14138_570# li_14138_570# li_11122_5650#
+ li_11122_5650# in in li_14138_570# in li_14138_570# in VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_AKSJZW_10 bias_d li_11121_570# bias_d op VSS bias_d op li_11121_570#
+ op bias_d bias_d bias_d op bias_d li_11121_570# VSS li_11121_570# bias_d bias_d
+ op li_11121_570# bias_d op op bias_d bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_0 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_AKSJZW_11 bias_d li_11121_570# bias_d op VSS bias_d op li_11121_570#
+ op bias_d bias_d bias_d op bias_d li_11121_570# VSS li_11121_570# bias_d bias_d
+ op li_11121_570# bias_d op op bias_d bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_1 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_2 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_3 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_4 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_5 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_6 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_7 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_8 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_9 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_10 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_11 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xbias_circuit_0 bias_c bias_e i_bias VDD bias_circuit_0/m1_1243_5997# bias_circuit_0/m1_3443_5997#
+ bias_a bias_circuit_0/m1_7347_1428# bias_circuit_0/m1_7639_1420# bias_circuit_0/m1_7169_923#
+ bias_circuit_0/m1_7461_921# bias_circuit_0/m1_7639_427# bias_circuit_0/m1_7347_423#
+ bias_b VSS bias_circuit_0/m1_3551_3596# bias_circuit_0/m1_5643_5997# bias_d bias_circuit
Xsky130_fd_pr__pfet_01v8_YVTMSC_0 on bias_c li_8436_5651# bias_c bias_c li_8436_5651#
+ on VDD bias_c li_8436_5651# bias_c on VDD bias_c on bias_c li_8436_5651# VDD on
+ bias_c li_8436_5651# bias_c on bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_1 on bias_c li_8436_5651# bias_c bias_c li_8436_5651#
+ on VDD bias_c li_8436_5651# bias_c on VDD bias_c on bias_c li_8436_5651# VDD on
+ bias_c li_8436_5651# bias_c on bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_0 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_YVTMSC_2 op bias_c li_11122_5650# bias_c bias_c li_11122_5650#
+ op VDD bias_c li_11122_5650# bias_c op VDD bias_c op bias_c li_11122_5650# VDD op
+ bias_c li_11122_5650# bias_c op bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_3 op bias_c li_11122_5650# bias_c bias_c li_11122_5650#
+ op VDD bias_c li_11122_5650# bias_c op VDD bias_c op bias_c li_11122_5650# VDD op
+ bias_c li_11122_5650# bias_c op bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_2 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_1 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_3 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_4 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_5 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_6 bias_d li_8434_570# bias_d on VSS bias_d on li_8434_570#
+ on bias_d bias_d bias_d on bias_d li_8434_570# VSS li_8434_570# bias_d bias_d on
+ li_8434_570# bias_d on on bias_d bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_7 bias_d li_8434_570# bias_d on VSS bias_d on li_8434_570#
+ on bias_d bias_d bias_d on bias_d li_8434_570# VSS li_8434_570# bias_d bias_d on
+ li_8434_570# bias_d on on bias_d bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
C0 bias_circuit_0/m1_3551_3596# VDD 0.15fF
C1 bias_circuit_0/m1_3551_3596# on 0.00fF
C2 in li_8436_5651# 0.01fF
C3 bias_c li_11122_5650# 3.17fF
C4 bias_c li_8434_570# 0.12fF
C5 m1_17097_3928# in 0.00fF
C6 cmc li_11122_5650# 0.13fF
C7 cmc li_14138_570# 26.78fF
C8 bias_circuit_0/m1_7639_1420# on 0.00fF
C9 bias_a bias_circuit_0/m1_7639_1420# 0.00fF
C10 m1_17393_3568# li_11122_5650# 0.00fF
C11 m1_17393_3568# li_14138_570# 0.01fF
C12 bias_a m1_15613_3568# 0.01fF
C13 li_8434_570# bias_e 0.00fF
C14 VDD li_11122_5650# 4.01fF
C15 on li_11122_5650# 0.12fF
C16 bias_b li_11122_5650# 4.74fF
C17 bias_a li_14138_570# 27.43fF
C18 li_8434_570# VDD 0.03fF
C19 li_8434_570# on 4.15fF
C20 bias_a li_8434_570# 10.56fF
C21 bias_d op 9.36fF
C22 bias_circuit_0/m1_5643_5997# VDD -0.00fF
C23 m1_18877_3928# in 0.01fF
C24 bias_c op 4.25fF
C25 m1_17393_3568# ip 0.00fF
C26 li_11121_570# li_11122_5650# 0.16fF
C27 li_11121_570# li_14138_570# 0.23fF
C28 bias_a ip 0.31fF
C29 li_11121_570# li_8434_570# 0.52fF
C30 bias_c bias_d 2.13fF
C31 op VDD 0.65fF
C32 li_8436_5651# li_11122_5650# 1.47fF
C33 on op 0.59fF
C34 in li_11122_5650# 1.14fF
C35 bias_b op 0.27fF
C36 bias_a op 0.52fF
C37 li_8436_5651# li_14138_570# 0.80fF
C38 in li_14138_570# 1.51fF
C39 li_8434_570# li_8436_5651# 0.16fF
C40 li_8434_570# bias_circuit_0/m1_7639_427# 0.01fF
C41 m1_17097_3928# li_14138_570# 0.00fF
C42 bias_d VDD 1.89fF
C43 bias_d on 10.13fF
C44 bias_d bias_b 0.02fF
C45 bias_a bias_d 2.86fF
C46 li_11121_570# op 4.14fF
C47 m1_18877_3928# li_14138_570# 0.00fF
C48 ip li_8436_5651# 1.22fF
C49 in ip 0.03fF
C50 bias_c VDD 6.20fF
C51 bias_c on 4.65fF
C52 bias_c bias_b 1.94fF
C53 bias_circuit_0/m1_7461_921# li_8434_570# 0.01fF
C54 m1_17097_3928# ip 0.01fF
C55 cmc bias_a 0.78fF
C56 op li_8436_5651# 0.12fF
C57 on bias_e 0.01fF
C58 li_11121_570# bias_d 6.30fF
C59 bias_a bias_e 0.00fF
C60 on VDD 0.63fF
C61 bias_b VDD 12.46fF
C62 on bias_b 0.27fF
C63 bias_a on 0.48fF
C64 li_8434_570# bias_circuit_0/m1_7639_1420# 0.01fF
C65 bias_d li_8436_5651# 0.66fF
C66 m1_15613_3568# li_14138_570# 0.01fF
C67 li_11122_5650# li_14138_570# 0.78fF
C68 li_11121_570# bias_c 0.12fF
C69 bias_c li_8436_5651# 4.18fF
C70 li_11121_570# VDD 0.02fF
C71 li_11121_570# on 0.17fF
C72 cmc in 0.31fF
C73 li_11121_570# bias_a 10.56fF
C74 m1_17393_3568# in 0.01fF
C75 ip m1_15613_3568# 0.01fF
C76 VDD li_8436_5651# 4.66fF
C77 on li_8436_5651# 2.52fF
C78 bias_b li_8436_5651# 4.47fF
C79 bias_a li_8436_5651# 0.14fF
C80 ip li_11122_5650# 0.01fF
C81 ip li_14138_570# 1.47fF
C82 bias_a bias_circuit_0/m1_7639_427# 0.01fF
C83 bias_circuit_0/m1_3551_3596# bias_d 0.03fF
C84 op li_11122_5650# 2.52fF
C85 op li_14138_570# 0.08fF
C86 li_8434_570# op 0.17fF
C87 bias_d bias_circuit_0/m1_7639_1420# 0.00fF
C88 cmc m1_18877_3928# 0.01fF
C89 bias_d li_11122_5650# 0.28fF
C90 bias_d li_14138_570# 0.02fF
C91 bias_c bias_circuit_0/m1_3551_3596# 0.00fF
C92 li_8434_570# bias_d 6.56fF
C93 m1_17393_3568# VSS 0.09fF $ **FLOATING
C94 m1_15613_3568# VSS 0.12fF $ **FLOATING
C95 m1_18877_3928# VSS 0.10fF $ **FLOATING
C96 m1_17097_3928# VSS 0.06fF $ **FLOATING
C97 on VSS 5.53fF
C98 li_11121_570# VSS 11.01fF
C99 li_11122_5650# VSS -32.46fF
C100 li_8434_570# VSS 10.89fF
C101 bias_a VSS -295.16fF
C102 li_8436_5651# VSS 5.93fF
C103 bias_circuit_0/m1_3551_3596# VSS -342.21fF
C104 bias_b VSS -361.08fF
C105 bias_circuit_0/m1_5643_5997# VSS 38.05fF
C106 bias_circuit_0/m1_3443_5997# VSS 35.85fF
C107 bias_circuit_0/m1_1243_5997# VSS 25.03fF
C108 VDD VSS 288.14fF
C109 i_bias VSS -60.67fF
C110 bias_c VSS -128.39fF
C111 bias_circuit_0/m1_7639_427# VSS 0.13fF
C112 bias_circuit_0/m1_7347_423# VSS 0.13fF
C113 bias_circuit_0/m1_7461_921# VSS 0.14fF
C114 bias_circuit_0/m1_7169_923# VSS 0.14fF
C115 bias_circuit_0/m1_7055_433# VSS 0.14fF
C116 bias_circuit_0/m1_6763_422# VSS 0.20fF
C117 bias_circuit_0/m1_6471_422# VSS 0.20fF
C118 bias_circuit_0/m1_7639_1420# VSS 0.13fF
C119 bias_circuit_0/m1_7347_1428# VSS 0.14fF
C120 bias_circuit_0/m1_6877_922# VSS 0.14fF
C121 bias_circuit_0/m1_6585_923# VSS 0.22fF
C122 bias_circuit_0/m1_6293_922# VSS 0.16fF
C123 bias_circuit_0/m1_7055_1417# VSS 0.13fF
C124 bias_circuit_0/m1_6763_1422# VSS 0.22fF
C125 bias_circuit_0/m1_6471_1426# VSS 0.22fF
C126 bias_e VSS 3.20fF
C127 bias_d VSS -235.00fF
C128 bias_circuit_0/li_3433_399# VSS 4.65fF
C129 li_14138_570# VSS 42.14fF
C130 cmc VSS -107.95fF
C131 op VSS 5.33fF
C132 in VSS -27.58fF
C133 ip VSS -28.74fF
.ends

.subckt pmos_tgate a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136# a_64_n136# a_160_n136#
+ a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136# a_n512_n234# a_256_n136#
+ VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_160_n136# a_64_n136# 0.33fF
C1 a_n224_n136# a_64_n136# 0.07fF
C2 a_448_n136# a_n508_n136# 0.02fF
C3 a_448_n136# a_352_n136# 0.33fF
C4 a_n32_n136# a_n416_n136# 0.05fF
C5 a_448_n136# a_n320_n136# 0.02fF
C6 a_256_n136# a_448_n136# 0.12fF
C7 a_n512_n234# a_n416_n136# 0.03fF
C8 a_n128_n136# a_n416_n136# 0.07fF
C9 a_n512_n234# a_n32_n136# 0.03fF
C10 a_n32_n136# a_n128_n136# 0.33fF
C11 a_448_n136# w_n646_n356# 0.13fF
C12 a_n512_n234# a_n128_n136# 0.03fF
C13 a_n508_n136# a_n416_n136# 0.33fF
C14 a_n508_n136# a_n32_n136# 0.04fF
C15 a_352_n136# a_n416_n136# 0.02fF
C16 a_n32_n136# a_352_n136# 0.05fF
C17 a_n508_n136# a_n512_n234# 0.03fF
C18 a_n508_n136# a_n128_n136# 0.05fF
C19 a_n320_n136# a_n416_n136# 0.33fF
C20 a_160_n136# a_448_n136# 0.07fF
C21 a_n32_n136# a_n320_n136# 0.07fF
C22 a_n512_n234# a_352_n136# 0.03fF
C23 a_352_n136# a_n128_n136# 0.04fF
C24 a_448_n136# a_n224_n136# 0.03fF
C25 a_256_n136# a_n416_n136# 0.03fF
C26 a_256_n136# a_n32_n136# 0.07fF
C27 a_n512_n234# a_n320_n136# 0.03fF
C28 a_n320_n136# a_n128_n136# 0.12fF
C29 a_256_n136# a_n512_n234# 0.03fF
C30 a_256_n136# a_n128_n136# 0.05fF
C31 w_n646_n356# a_n416_n136# 0.08fF
C32 a_n32_n136# w_n646_n356# 0.05fF
C33 a_n508_n136# a_352_n136# 0.02fF
C34 a_n512_n234# w_n646_n356# 1.47fF
C35 w_n646_n356# a_n128_n136# 0.05fF
C36 a_n508_n136# a_n320_n136# 0.12fF
C37 a_256_n136# a_n508_n136# 0.02fF
C38 a_n320_n136# a_352_n136# 0.03fF
C39 a_256_n136# a_352_n136# 0.33fF
C40 a_160_n136# a_n416_n136# 0.03fF
C41 a_160_n136# a_n32_n136# 0.12fF
C42 a_n224_n136# a_n416_n136# 0.12fF
C43 a_n224_n136# a_n32_n136# 0.12fF
C44 a_256_n136# a_n320_n136# 0.03fF
C45 a_n508_n136# w_n646_n356# 0.13fF
C46 a_160_n136# a_n512_n234# 0.03fF
C47 a_160_n136# a_n128_n136# 0.07fF
C48 w_n646_n356# a_352_n136# 0.08fF
C49 a_n224_n136# a_n512_n234# 0.03fF
C50 a_n224_n136# a_n128_n136# 0.33fF
C51 w_n646_n356# a_n320_n136# 0.06fF
C52 a_256_n136# w_n646_n356# 0.06fF
C53 a_448_n136# a_64_n136# 0.05fF
C54 a_160_n136# a_n508_n136# 0.03fF
C55 a_n508_n136# a_n224_n136# 0.07fF
C56 a_160_n136# a_352_n136# 0.12fF
C57 a_n224_n136# a_352_n136# 0.03fF
C58 a_160_n136# a_n320_n136# 0.04fF
C59 a_n224_n136# a_n320_n136# 0.33fF
C60 a_256_n136# a_160_n136# 0.33fF
C61 a_256_n136# a_n224_n136# 0.04fF
C62 a_160_n136# w_n646_n356# 0.06fF
C63 a_n224_n136# w_n646_n356# 0.06fF
C64 a_64_n136# a_n416_n136# 0.04fF
C65 a_n32_n136# a_64_n136# 0.33fF
C66 a_n512_n234# a_64_n136# 0.03fF
C67 a_64_n136# a_n128_n136# 0.12fF
C68 a_160_n136# a_n224_n136# 0.05fF
C69 a_n508_n136# a_64_n136# 0.03fF
C70 a_64_n136# a_352_n136# 0.07fF
C71 a_n320_n136# a_64_n136# 0.05fF
C72 a_256_n136# a_64_n136# 0.12fF
C73 w_n646_n356# a_64_n136# 0.05fF
C74 a_448_n136# a_n416_n136# 0.02fF
C75 a_448_n136# a_n32_n136# 0.04fF
C76 a_448_n136# a_n512_n234# 0.03fF
C77 a_448_n136# a_n128_n136# 0.03fF
C78 w_n646_n356# VSUBS 2.52fF
.ends

.subckt nmos_tgate a_256_n52# a_n32_n52# a_n224_n52# a_448_n52# a_n416_n52# a_160_n52#
+ a_n610_n226# a_n128_n52# a_352_n52# a_n320_n52# a_n508_n52# a_n512_n149# a_64_n52#
X0 a_n32_n52# a_n512_n149# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n149# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n149# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n149# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n149# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n149# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n149# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n149# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n149# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n149# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_352_n52# a_n320_n52# 0.01fF
C1 a_n416_n52# a_n508_n52# 0.13fF
C2 a_n416_n52# a_n128_n52# 0.03fF
C3 a_352_n52# a_448_n52# 0.13fF
C4 a_n32_n52# a_n416_n52# 0.02fF
C5 a_n224_n52# a_n508_n52# 0.03fF
C6 a_n224_n52# a_n128_n52# 0.13fF
C7 a_n224_n52# a_n32_n52# 0.05fF
C8 a_160_n52# a_256_n52# 0.13fF
C9 a_n416_n52# a_352_n52# 0.01fF
C10 a_n224_n52# a_352_n52# 0.01fF
C11 a_256_n52# a_n508_n52# 0.01fF
C12 a_256_n52# a_n128_n52# 0.02fF
C13 a_n512_n149# a_64_n52# 0.03fF
C14 a_n32_n52# a_256_n52# 0.03fF
C15 a_n320_n52# a_64_n52# 0.02fF
C16 a_n512_n149# a_n320_n52# 0.03fF
C17 a_64_n52# a_448_n52# 0.02fF
C18 a_n512_n149# a_448_n52# 0.03fF
C19 a_352_n52# a_256_n52# 0.13fF
C20 a_n320_n52# a_448_n52# 0.01fF
C21 a_n416_n52# a_64_n52# 0.02fF
C22 a_n512_n149# a_n416_n52# 0.03fF
C23 a_n416_n52# a_n320_n52# 0.13fF
C24 a_n224_n52# a_64_n52# 0.03fF
C25 a_n224_n52# a_n512_n149# 0.03fF
C26 a_n416_n52# a_448_n52# 0.01fF
C27 a_n224_n52# a_n320_n52# 0.13fF
C28 a_160_n52# a_n508_n52# 0.01fF
C29 a_160_n52# a_n128_n52# 0.03fF
C30 a_n224_n52# a_448_n52# 0.01fF
C31 a_n32_n52# a_160_n52# 0.05fF
C32 a_256_n52# a_64_n52# 0.05fF
C33 a_n512_n149# a_256_n52# 0.03fF
C34 a_n224_n52# a_n416_n52# 0.05fF
C35 a_n128_n52# a_n508_n52# 0.02fF
C36 a_160_n52# a_352_n52# 0.05fF
C37 a_256_n52# a_n320_n52# 0.01fF
C38 a_n32_n52# a_n508_n52# 0.02fF
C39 a_n32_n52# a_n128_n52# 0.13fF
C40 a_256_n52# a_448_n52# 0.05fF
C41 a_352_n52# a_n508_n52# 0.01fF
C42 a_352_n52# a_n128_n52# 0.02fF
C43 a_n416_n52# a_256_n52# 0.01fF
C44 a_n32_n52# a_352_n52# 0.02fF
C45 a_n224_n52# a_256_n52# 0.02fF
C46 a_160_n52# a_64_n52# 0.13fF
C47 a_n512_n149# a_160_n52# 0.03fF
C48 a_160_n52# a_n320_n52# 0.02fF
C49 a_160_n52# a_448_n52# 0.03fF
C50 a_n508_n52# a_64_n52# 0.01fF
C51 a_n512_n149# a_n508_n52# 0.03fF
C52 a_n128_n52# a_64_n52# 0.05fF
C53 a_n512_n149# a_n128_n52# 0.03fF
C54 a_n32_n52# a_64_n52# 0.13fF
C55 a_n512_n149# a_n32_n52# 0.03fF
C56 a_n508_n52# a_n320_n52# 0.05fF
C57 a_n128_n52# a_n320_n52# 0.05fF
C58 a_160_n52# a_n416_n52# 0.01fF
C59 a_n32_n52# a_n320_n52# 0.03fF
C60 a_n508_n52# a_448_n52# 0.01fF
C61 a_n128_n52# a_448_n52# 0.01fF
C62 a_n32_n52# a_448_n52# 0.02fF
C63 a_n224_n52# a_160_n52# 0.02fF
C64 a_352_n52# a_64_n52# 0.03fF
C65 a_n512_n149# a_352_n52# 0.03fF
C66 a_448_n52# a_n610_n226# 0.07fF
C67 a_352_n52# a_n610_n226# 0.05fF
C68 a_256_n52# a_n610_n226# 0.04fF
C69 a_160_n52# a_n610_n226# 0.04fF
C70 a_64_n52# a_n610_n226# 0.04fF
C71 a_n32_n52# a_n610_n226# 0.04fF
C72 a_n128_n52# a_n610_n226# 0.04fF
C73 a_n224_n52# a_n610_n226# 0.04fF
C74 a_n320_n52# a_n610_n226# 0.04fF
C75 a_n416_n52# a_n610_n226# 0.05fF
C76 a_n508_n52# a_n610_n226# 0.07fF
C77 a_n512_n149# a_n610_n226# 1.83fF
.ends

.subckt transmission_gate en en_b VDD in out VSS
Xpmos_tgate_0 in in out in out in out VDD in out out en_b out VSS pmos_tgate
Xnmos_tgate_0 out in in out in in VSS out in out out en out nmos_tgate
C0 VDD en_b -0.11fF
C1 VDD en 0.12fF
C2 en_b en 0.07fF
C3 out VDD 0.29fF
C4 VDD in 0.70fF
C5 out en_b 0.01fF
C6 en_b in 0.15fF
C7 out en 0.01fF
C8 in en 0.13fF
C9 out in 0.77fF
C10 en VSS 1.70fF
C11 out VSS 0.57fF
C12 in VSS 1.13fF
C13 en_b VSS 0.09fF
C14 VDD VSS 3.16fF
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580# VSUBS
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
C0 m3_n630_n580# c1_n530_n480# 2.88fF
C1 m3_n630_n580# VSUBS 1.37fF
.ends

.subckt sc_cmfb cm op cmc p2_b p2 p1 on unit_cap_mim_m3m4_30/m3_n630_n580# transmission_gate_8/in
+ transmission_gate_4/out bias_a VDD transmission_gate_7/in VSS p1_b
Xtransmission_gate_10 p1 p1_b VDD transmission_gate_3/out on VSS transmission_gate
Xtransmission_gate_11 p1 p1_b VDD transmission_gate_4/out op VSS transmission_gate
Xtransmission_gate_0 p1 p1_b VDD cm transmission_gate_7/in VSS transmission_gate
Xtransmission_gate_1 p1 p1_b VDD cm transmission_gate_6/in VSS transmission_gate
Xtransmission_gate_2 p1 p1_b VDD bias_a transmission_gate_8/in VSS transmission_gate
Xtransmission_gate_3 p2 p2_b VDD cm transmission_gate_3/out VSS transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xtransmission_gate_4 p2 p2_b VDD cm transmission_gate_4/out VSS transmission_gate
Xunit_cap_mim_m3m4_1 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_5 p2 p2_b VDD bias_a transmission_gate_9/in VSS transmission_gate
Xunit_cap_mim_m3m4_2 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_6 p2 p2_b VDD transmission_gate_6/in op VSS transmission_gate
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_7 p2 p2_b VDD transmission_gate_7/in on VSS transmission_gate
Xunit_cap_mim_m3m4_4 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_8 p2 p2_b VDD transmission_gate_8/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_9 p1 p1_b VDD transmission_gate_9/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
C0 unit_cap_mim_m3m4_24/m3_n630_n580# p1 0.08fF
C1 on transmission_gate_8/in 0.56fF
C2 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C3 unit_cap_mim_m3m4_29/m3_n630_n580# p1_b 0.05fF
C4 unit_cap_mim_m3m4_18/m3_n630_n580# cmc 0.17fF
C5 cm transmission_gate_4/out 0.07fF
C6 transmission_gate_8/in transmission_gate_4/out 0.27fF
C7 p2 unit_cap_mim_m3m4_17/m3_n630_n580# 0.04fF
C8 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C9 VDD cm 1.83fF
C10 VDD transmission_gate_8/in -0.07fF
C11 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580# -0.18fF
C12 unit_cap_mim_m3m4_19/m3_n630_n580# p1_b 0.06fF
C13 unit_cap_mim_m3m4_30/m3_n630_n580# p1_b 0.01fF
C14 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C15 cmc p1_b 0.53fF
C16 p1 on 0.49fF
C17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C18 transmission_gate_9/in unit_cap_mim_m3m4_16/m3_n630_n580# 0.17fF
C19 p1 transmission_gate_4/out 0.80fF
C20 unit_cap_mim_m3m4_22/c1_n530_n480# transmission_gate_9/in -0.37fF
C21 unit_cap_mim_m3m4_28/c1_n530_n480# transmission_gate_6/in 0.05fF
C22 VDD p1 1.10fF
C23 transmission_gate_6/in op 0.61fF
C24 unit_cap_mim_m3m4_23/m3_n630_n580# transmission_gate_9/in 0.17fF
C25 bias_a transmission_gate_6/in 0.07fF
C26 transmission_gate_7/in unit_cap_mim_m3m4_20/c1_n530_n480# -0.18fF
C27 p2 transmission_gate_6/in 0.61fF
C28 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C29 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C30 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.17fF
C31 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C32 transmission_gate_4/out unit_cap_mim_m3m4_31/c1_n530_n480# 0.05fF
C33 on cmc -0.58fF
C34 transmission_gate_3/out unit_cap_mim_m3m4_23/c1_n530_n480# -0.24fF
C35 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580# -0.33fF
C36 unit_cap_mim_m3m4_27/c1_n530_n480# p1_b 0.06fF
C37 unit_cap_mim_m3m4_30/m3_n630_n580# transmission_gate_4/out -0.80fF
C38 cmc transmission_gate_4/out 0.15fF
C39 unit_cap_mim_m3m4_28/m3_n630_n580# op 0.66fF
C40 p2_b transmission_gate_7/in 0.41fF
C41 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.17fF
C42 VDD cmc 1.23fF
C43 unit_cap_mim_m3m4_30/c1_n530_n480# op 0.18fF
C44 unit_cap_mim_m3m4_27/m3_n630_n580# cmc 0.10fF
C45 transmission_gate_3/out op 0.57fF
C46 transmission_gate_3/out bias_a 0.07fF
C47 p2 transmission_gate_3/out 0.15fF
C48 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C49 op unit_cap_mim_m3m4_31/m3_n630_n580# 0.03fF
C50 transmission_gate_7/in p1_b 0.40fF
C51 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580# -0.14fF
C52 unit_cap_mim_m3m4_22/m3_n630_n580# p1 0.06fF
C53 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_27/c1_n530_n480# -0.37fF
C54 transmission_gate_6/in unit_cap_mim_m3m4_29/c1_n530_n480# -0.37fF
C55 transmission_gate_8/in op 0.40fF
C56 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C57 transmission_gate_8/in bias_a 0.04fF
C58 cm bias_a 1.15fF
C59 p2 transmission_gate_8/in 0.63fF
C60 p2 cm 1.33fF
C61 unit_cap_mim_m3m4_34/m3_n630_n580# transmission_gate_8/in 0.38fF
C62 on transmission_gate_7/in 3.15fF
C63 unit_cap_mim_m3m4_28/c1_n530_n480# p1 0.11fF
C64 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580# -0.21fF
C65 unit_cap_mim_m3m4_22/m3_n630_n580# cmc 0.71fF
C66 transmission_gate_4/out transmission_gate_7/in 0.62fF
C67 p1 op 0.52fF
C68 unit_cap_mim_m3m4_25/c1_n530_n480# p1_b 0.06fF
C69 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.17fF
C70 transmission_gate_9/in transmission_gate_6/in 0.03fF
C71 p2_b p1_b 2.92fF
C72 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580# -0.19fF
C73 p1 bias_a 0.81fF
C74 VDD transmission_gate_7/in -0.16fF
C75 p2 p1 2.82fF
C76 unit_cap_mim_m3m4_24/c1_n530_n480# p1 0.11fF
C77 transmission_gate_3/out unit_cap_mim_m3m4_23/m3_n630_n580# -0.30fF
C78 unit_cap_mim_m3m4_29/m3_n630_n580# op 0.39fF
C79 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580# -0.35fF
C80 unit_cap_mim_m3m4_18/m3_n630_n580# p1_b 0.06fF
C81 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C82 on unit_cap_mim_m3m4_20/c1_n530_n480# 0.15fF
C83 unit_cap_mim_m3m4_31/c1_n530_n480# op 0.05fF
C84 unit_cap_mim_m3m4_30/m3_n630_n580# op 0.56fF
C85 cmc op -0.30fF
C86 transmission_gate_8/in unit_cap_mim_m3m4_21/c1_n530_n480# -0.41fF
C87 unit_cap_mim_m3m4_35/m3_n630_n580# p1_b 0.01fF
C88 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_35/c1_n530_n480# 0.06fF
C89 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_35/c1_n530_n480# 0.06fF
C90 p2_b on 0.34fF
C91 transmission_gate_4/out unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C92 unit_cap_mim_m3m4_26/c1_n530_n480# p1 0.11fF
C93 unit_cap_mim_m3m4_24/m3_n630_n580# p1_b 0.06fF
C94 transmission_gate_3/out transmission_gate_9/in 1.33fF
C95 p2 cmc 0.25fF
C96 p2_b transmission_gate_4/out 0.05fF
C97 p2_b VDD 1.67fF
C98 p1 unit_cap_mim_m3m4_16/m3_n630_n580# 0.08fF
C99 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.12fF
C100 transmission_gate_9/in unit_cap_mim_m3m4_31/m3_n630_n580# 0.12fF
C101 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C102 on p1_b 0.45fF
C103 unit_cap_mim_m3m4_27/c1_n530_n480# op 0.01fF
C104 p1 unit_cap_mim_m3m4_29/c1_n530_n480# 0.11fF
C105 transmission_gate_3/out unit_cap_mim_m3m4_17/m3_n630_n580# -0.23fF
C106 unit_cap_mim_m3m4_23/m3_n630_n580# p1 0.06fF
C107 transmission_gate_4/out p1_b 0.55fF
C108 p2 unit_cap_mim_m3m4_27/c1_n530_n480# 0.04fF
C109 VDD p1_b 1.01fF
C110 transmission_gate_9/in transmission_gate_8/in 0.93fF
C111 cm transmission_gate_9/in 0.04fF
C112 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C113 unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_29/c1_n530_n480# -0.29fF
C114 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.17fF
C115 cmc unit_cap_mim_m3m4_21/c1_n530_n480# 0.13fF
C116 unit_cap_mim_m3m4_22/c1_n530_n480# cmc 0.13fF
C117 unit_cap_mim_m3m4_28/m3_n630_n580# transmission_gate_6/in -0.13fF
C118 unit_cap_mim_m3m4_28/c1_n530_n480# transmission_gate_7/in 0.06fF
C119 p1 transmission_gate_9/in 0.70fF
C120 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.12fF
C121 transmission_gate_7/in op 2.65fF
C122 on transmission_gate_4/out 3.25fF
C123 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C124 transmission_gate_3/out transmission_gate_6/in 0.75fF
C125 bias_a transmission_gate_7/in 0.11fF
C126 VDD on 0.88fF
C127 p2 transmission_gate_7/in 0.60fF
C128 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_8/in 0.17fF
C129 VDD transmission_gate_4/out -0.06fF
C130 p1 unit_cap_mim_m3m4_17/m3_n630_n580# 0.08fF
C131 cmc unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C132 transmission_gate_9/in cmc 3.45fF
C133 unit_cap_mim_m3m4_20/m3_n630_n580# p1 0.06fF
C134 unit_cap_mim_m3m4_22/m3_n630_n580# p1_b 0.05fF
C135 cm transmission_gate_6/in 0.17fF
C136 transmission_gate_8/in transmission_gate_6/in -0.41fF
C137 p2_b op 0.40fF
C138 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.10fF
C139 p2_b bias_a 0.48fF
C140 p2 unit_cap_mim_m3m4_25/c1_n530_n480# 0.04fF
C141 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C142 p2 p2_b 6.58fF
C143 cmc unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C144 on unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C145 p1 transmission_gate_6/in 0.38fF
C146 transmission_gate_8/in unit_cap_mim_m3m4_28/m3_n630_n580# 0.10fF
C147 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_25/c1_n530_n480# -0.32fF
C148 unit_cap_mim_m3m4_28/c1_n530_n480# p1_b 0.06fF
C149 op p1_b 0.28fF
C150 unit_cap_mim_m3m4_29/m3_n630_n580# transmission_gate_6/in -0.80fF
C151 bias_a p1_b 0.52fF
C152 transmission_gate_3/out cm 0.17fF
C153 transmission_gate_3/out transmission_gate_8/in 0.16fF
C154 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C155 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480# 0.06fF
C156 p2 p1_b 5.94fF
C157 unit_cap_mim_m3m4_24/c1_n530_n480# p1_b 0.06fF
C158 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_34/m3_n630_n580# 0.17fF
C159 transmission_gate_8/in unit_cap_mim_m3m4_21/m3_n630_n580# -1.15fF
C160 on unit_cap_mim_m3m4_23/c1_n530_n480# 0.19fF
C161 unit_cap_mim_m3m4_24/m3_n630_n580# p2 0.05fF
C162 transmission_gate_4/out unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C163 cmc transmission_gate_6/in 0.96fF
C164 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_24/c1_n530_n480# -0.30fF
C165 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480# 0.06fF
C166 transmission_gate_3/out p1 0.72fF
C167 unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580# 0.17fF
C168 transmission_gate_9/in transmission_gate_7/in 0.04fF
C169 on op 2.09fF
C170 p1 unit_cap_mim_m3m4_21/m3_n630_n580# 0.06fF
C171 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C172 transmission_gate_4/out op 1.12fF
C173 cmc unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C174 unit_cap_mim_m3m4_26/c1_n530_n480# p1_b 0.06fF
C175 cm transmission_gate_8/in 0.03fF
C176 p2 on 0.24fF
C177 transmission_gate_4/out bias_a 0.10fF
C178 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_31/c1_n530_n480# 0.06fF
C179 VDD op 0.89fF
C180 unit_cap_mim_m3m4_27/m3_n630_n580# op 0.48fF
C181 p2 transmission_gate_4/out 0.15fF
C182 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_30/c1_n530_n480# -0.12fF
C183 VDD bias_a 0.99fF
C184 unit_cap_mim_m3m4_16/m3_n630_n580# p1_b 0.06fF
C185 p2 VDD 4.16fF
C186 unit_cap_mim_m3m4_27/c1_n530_n480# transmission_gate_6/in -0.13fF
C187 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C188 transmission_gate_3/out cmc 0.74fF
C189 cm p1 1.50fF
C190 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.10fF
C191 p1 transmission_gate_8/in 0.39fF
C192 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_7/in -0.56fF
C193 cmc unit_cap_mim_m3m4_21/m3_n630_n580# 0.69fF
C194 unit_cap_mim_m3m4_29/c1_n530_n480# p1_b 0.06fF
C195 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580# -0.25fF
C196 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580# -0.21fF
C197 unit_cap_mim_m3m4_23/m3_n630_n580# p1_b 0.05fF
C198 p2_b transmission_gate_9/in 0.01fF
C199 unit_cap_mim_m3m4_26/c1_n530_n480# on 0.06fF
C200 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.17fF
C201 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_35/c1_n530_n480# -0.13fF
C202 on unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C203 unit_cap_mim_m3m4_17/c1_n530_n480# op 0.06fF
C204 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_20/c1_n530_n480# -0.19fF
C205 cmc unit_cap_mim_m3m4_26/m3_n630_n580# 0.10fF
C206 transmission_gate_8/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.17fF
C207 unit_cap_mim_m3m4_16/m3_n630_n580# transmission_gate_4/out -0.28fF
C208 transmission_gate_7/in transmission_gate_6/in 0.47fF
C209 cmc transmission_gate_8/in 1.73fF
C210 p1 unit_cap_mim_m3m4_29/m3_n630_n580# 0.06fF
C211 transmission_gate_9/in p1_b 0.59fF
C212 unit_cap_mim_m3m4_23/m3_n630_n580# on 0.47fF
C213 unit_cap_mim_m3m4_33/c1_n530_n480# op 0.06fF
C214 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580# -0.20fF
C215 unit_cap_mim_m3m4_24/m3_n630_n580# transmission_gate_9/in 0.23fF
C216 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C217 p1 unit_cap_mim_m3m4_19/m3_n630_n580# 0.08fF
C218 unit_cap_mim_m3m4_30/m3_n630_n580# p1 0.06fF
C219 p1 cmc 0.49fF
C220 op unit_cap_mim_m3m4_23/c1_n530_n480# 0.13fF
C221 unit_cap_mim_m3m4_17/m3_n630_n580# p1_b 0.06fF
C222 transmission_gate_3/out transmission_gate_7/in 0.30fF
C223 transmission_gate_9/in on 0.82fF
C224 unit_cap_mim_m3m4_20/m3_n630_n580# p1_b 0.05fF
C225 p2_b transmission_gate_6/in 0.42fF
C226 unit_cap_mim_m3m4_28/c1_n530_n480# op 0.17fF
C227 transmission_gate_9/in transmission_gate_4/out -0.11fF
C228 unit_cap_mim_m3m4_34/c1_n530_n480# transmission_gate_7/in 0.06fF
C229 unit_cap_mim_m3m4_19/c1_n530_n480# transmission_gate_7/in 0.06fF
C230 VDD transmission_gate_9/in -0.11fF
C231 p2 unit_cap_mim_m3m4_28/c1_n530_n480# 0.04fF
C232 unit_cap_mim_m3m4_18/m3_n630_n580# transmission_gate_6/in 0.08fF
C233 p1 unit_cap_mim_m3m4_27/c1_n530_n480# 0.11fF
C234 p2 op 0.16fF
C235 unit_cap_mim_m3m4_18/c1_n530_n480# on 0.06fF
C236 p2 bias_a 0.60fF
C237 transmission_gate_6/in p1_b 0.41fF
C238 p2 unit_cap_mim_m3m4_24/c1_n530_n480# 0.04fF
C239 cm transmission_gate_7/in 0.10fF
C240 transmission_gate_8/in transmission_gate_7/in -0.35fF
C241 unit_cap_mim_m3m4_20/m3_n630_n580# on 0.61fF
C242 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580# -0.19fF
C243 p2_b transmission_gate_3/out 0.10fF
C244 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.12fF
C245 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C246 p1 transmission_gate_7/in 0.39fF
C247 p2 unit_cap_mim_m3m4_26/c1_n530_n480# 0.04fF
C248 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_32/c1_n530_n480# -0.20fF
C249 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_23/c1_n530_n480# -0.19fF
C250 on transmission_gate_6/in 0.41fF
C251 transmission_gate_3/out p1_b 0.59fF
C252 unit_cap_mim_m3m4_22/c1_n530_n480# op 0.07fF
C253 transmission_gate_4/out transmission_gate_6/in 0.48fF
C254 p2 unit_cap_mim_m3m4_16/m3_n630_n580# 0.05fF
C255 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C256 unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_9/in -0.80fF
C257 unit_cap_mim_m3m4_21/m3_n630_n580# p1_b 0.05fF
C258 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C259 p2_b transmission_gate_8/in 0.40fF
C260 p2_b cm 1.01fF
C261 VDD transmission_gate_6/in 0.03fF
C262 unit_cap_mim_m3m4_29/c1_n530_n480# op 0.03fF
C263 unit_cap_mim_m3m4_27/m3_n630_n580# transmission_gate_6/in 0.13fF
C264 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580# -0.20fF
C265 transmission_gate_7/in unit_cap_mim_m3m4_19/m3_n630_n580# -0.28fF
C266 cmc transmission_gate_7/in 0.11fF
C267 p2 unit_cap_mim_m3m4_29/c1_n530_n480# 0.04fF
C268 p1 unit_cap_mim_m3m4_25/c1_n530_n480# 0.11fF
C269 p2_b p1 2.16fF
C270 unit_cap_mim_m3m4_30/c1_n530_n480# transmission_gate_4/out -0.37fF
C271 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580# 0.12fF
C272 transmission_gate_3/out on 0.39fF
C273 transmission_gate_8/in p1_b 0.17fF
C274 cm p1_b 1.15fF
C275 unit_cap_mim_m3m4_35/m3_n630_n580# transmission_gate_8/in -0.10fF
C276 transmission_gate_3/out transmission_gate_4/out 0.38fF
C277 transmission_gate_9/in op 0.47fF
C278 unit_cap_mim_m3m4_16/c1_n530_n480# transmission_gate_4/out 0.06fF
C279 unit_cap_mim_m3m4_18/m3_n630_n580# p1 0.08fF
C280 transmission_gate_9/in bias_a 0.02fF
C281 transmission_gate_3/out VDD -0.05fF
C282 p2 transmission_gate_9/in 0.14fF
C283 transmission_gate_4/out unit_cap_mim_m3m4_31/m3_n630_n580# 0.32fF
C284 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C285 p1 p1_b 8.88fF
C286 unit_cap_mim_m3m4_35/m3_n630_n580# p1 0.07fF
C287 p2_b cmc 0.12fF
C288 unit_cap_mim_m3m4_25/m3_n630_n580# transmission_gate_9/in 0.27fF
C289 unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C290 unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.39fF
C291 unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C292 unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.51fF
C293 unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C294 unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.74fF
C295 unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C296 unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.51fF
C297 unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.51fF
C298 unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.82fF
C299 unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.60fF
C300 cmc VSS 7.45fF
C301 unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.61fF
C302 unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.61fF
C303 unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C304 unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C305 p2 VSS 148.24fF
C306 p2_b VSS 41.62fF
C307 unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.84fF
C308 unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C309 unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.39fF
C310 unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C311 unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.04fF
C312 transmission_gate_9/in VSS 2.27fF
C313 transmission_gate_4/out VSS -3.31fF
C314 transmission_gate_3/out VSS 2.40fF
C315 p1 VSS 111.99fF
C316 transmission_gate_8/in VSS -2.63fF
C317 bias_a VSS 11.61fF
C318 transmission_gate_6/in VSS -13.21fF
C319 transmission_gate_7/in VSS 8.85fF
C320 cm VSS 13.12fF
C321 op VSS 0.25fF
C322 p1_b VSS 173.74fF
C323 VDD VSS 71.01fF
C324 on VSS -22.35fF
.ends

.subckt ota_v2 ip in p1 p1_b p2 p2_b op on i_bias cm VDD VSS
Xota_v2_without_cmfb_0 in ota_v2_without_cmfb_0/bias_c cm op on i_bias VDD ota_v2_without_cmfb_0/bias_d
+ VSS ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# ota_v2_without_cmfb_0/li_11121_570#
+ ota_v2_without_cmfb_0/li_11122_5650# sc_cmfb_0/cmc ota_v2_without_cmfb_0/li_14138_570#
+ ota_v2_without_cmfb_0/li_8434_570# ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/bias_b
+ ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997#
+ sc_cmfb_0/bias_a ip ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# ota_v2_without_cmfb
Xsc_cmfb_0 cm op sc_cmfb_0/cmc p2_b p2 p1 on sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/bias_a
+ VDD sc_cmfb_0/transmission_gate_7/in VSS p1_b sc_cmfb
C0 op ota_v2_without_cmfb_0/bias_c 1.56fF
C1 op sc_cmfb_0/cmc 0.37fF
C2 cm ota_v2_without_cmfb_0/li_14138_570# 1.29fF
C3 VDD p1_b -0.00fF
C4 ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C5 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# 0.00fF
C6 p1 sc_cmfb_0/transmission_gate_4/out 0.05fF
C7 VDD op 3.19fF
C8 ota_v2_without_cmfb_0/li_14138_570# sc_cmfb_0/cmc 0.03fF
C9 ota_v2_without_cmfb_0/bias_b sc_cmfb_0/bias_a 0.15fF
C10 cm ota_v2_without_cmfb_0/li_11121_570# 0.39fF
C11 ota_v2_without_cmfb_0/li_8434_570# on 0.00fF
C12 VDD sc_cmfb_0/transmission_gate_7/in 0.01fF
C13 VDD sc_cmfb_0/transmission_gate_4/out 0.04fF
C14 ota_v2_without_cmfb_0/li_8436_5651# ip -0.00fF
C15 ota_v2_without_cmfb_0/li_11122_5650# op 0.36fF
C16 cm on 3.11fF
C17 cm sc_cmfb_0/bias_a 3.22fF
C18 op ota_v2_without_cmfb_0/li_8436_5651# 0.40fF
C19 ota_v2_without_cmfb_0/bias_d op -0.00fF
C20 ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# cm 0.23fF
C21 p1 on 0.01fF
C22 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.02fF
C23 p1 sc_cmfb_0/bias_a 0.00fF
C24 on ota_v2_without_cmfb_0/bias_c -0.00fF
C25 sc_cmfb_0/cmc on 0.31fF
C26 cm ota_v2_without_cmfb_0/bias_b 3.45fF
C27 sc_cmfb_0/bias_a ota_v2_without_cmfb_0/bias_c 2.52fF
C28 ota_v2_without_cmfb_0/li_14138_570# ota_v2_without_cmfb_0/li_8436_5651# 0.00fF
C29 ota_v2_without_cmfb_0/li_8434_570# cm 0.38fF
C30 op ip 0.01fF
C31 p1_b op 0.00fF
C32 VDD on 0.45fF
C33 ota_v2_without_cmfb_0/bias_b ota_v2_without_cmfb_0/bias_c 0.26fF
C34 VDD sc_cmfb_0/bias_a 0.02fF
C35 ota_v2_without_cmfb_0/li_14138_570# ip 0.00fF
C36 VDD ota_v2_without_cmfb_0/bias_b 0.16fF
C37 sc_cmfb_0/transmission_gate_4/out p1_b 0.00fF
C38 ota_v2_without_cmfb_0/bias_d ota_v2_without_cmfb_0/li_11121_570# -0.00fF
C39 cm ota_v2_without_cmfb_0/bias_c 2.51fF
C40 ota_v2_without_cmfb_0/li_14138_570# op 0.00fF
C41 cm sc_cmfb_0/cmc -2.78fF
C42 i_bias ota_v2_without_cmfb_0/bias_c 0.00fF
C43 ota_v2_without_cmfb_0/li_11122_5650# on 0.22fF
C44 sc_cmfb_0/transmission_gate_4/out op -0.00fF
C45 ota_v2_without_cmfb_0/li_8436_5651# on 0.37fF
C46 ota_v2_without_cmfb_0/bias_d on 7.34fF
C47 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/bias_a 0.00fF
C48 ota_v2_without_cmfb_0/bias_d sc_cmfb_0/bias_a -0.00fF
C49 VDD cm -0.07fF
C50 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# 0.00fF
C51 ota_v2_without_cmfb_0/bias_b ota_v2_without_cmfb_0/li_11122_5650# -0.00fF
C52 ota_v2_without_cmfb_0/li_11121_570# op 0.00fF
C53 VDD sc_cmfb_0/cmc -0.08fF
C54 ota_v2_without_cmfb_0/li_14138_570# in -0.00fF
C55 p1_b on 0.01fF
C56 ota_v2_without_cmfb_0/li_8434_570# ota_v2_without_cmfb_0/bias_d -0.00fF
C57 p1_b sc_cmfb_0/bias_a 0.00fF
C58 p1 p2_b 0.00fF
C59 op on 3.51fF
C60 ota_v2_without_cmfb_0/bias_d cm 4.24fF
C61 p1 sc_cmfb_0/transmission_gate_8/in 0.00fF
C62 ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/bias_c 0.00fF
C63 ota_v2_without_cmfb_0/li_14138_570# on 0.01fF
C64 ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/bias_c -0.00fF
C65 cm p1_b 0.01fF
C66 VDD ota_v2_without_cmfb_0/li_11122_5650# 0.23fF
C67 p1 p1_b 0.00fF
C68 ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VDD 0.00fF
C69 VDD sc_cmfb_0/transmission_gate_8/in 0.02fF
C70 VDD ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C71 cm op 1.43fF
C72 p1 op 0.01fF
C73 ota_v2_without_cmfb_0/li_11121_570# on 0.01fF
C74 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C75 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.37fF
C76 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C77 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C78 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C79 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C80 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C81 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C82 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C83 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.37fF
C84 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.37fF
C85 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C86 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C87 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C88 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C89 p2 VSS 147.98fF
C90 p2_b VSS 40.26fF
C91 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C92 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C93 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C94 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C95 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.86fF
C96 sc_cmfb_0/transmission_gate_9/in VSS 0.88fF
C97 sc_cmfb_0/transmission_gate_4/out VSS -4.45fF
C98 sc_cmfb_0/transmission_gate_3/out VSS 1.32fF
C99 p1 VSS 111.49fF
C100 sc_cmfb_0/transmission_gate_8/in VSS -3.90fF
C101 sc_cmfb_0/transmission_gate_6/in VSS -14.61fF
C102 sc_cmfb_0/transmission_gate_7/in VSS 7.44fF
C103 cm VSS 34.63fF
C104 op VSS 4.87fF
C105 p1_b VSS 173.22fF
C106 on VSS -20.35fF
C107 ota_v2_without_cmfb_0/m1_17393_3568# VSS 0.03fF $ **FLOATING
C108 ota_v2_without_cmfb_0/m1_15613_3568# VSS 0.05fF $ **FLOATING
C109 ota_v2_without_cmfb_0/m1_18877_3928# VSS 0.05fF $ **FLOATING
C110 ota_v2_without_cmfb_0/m1_17097_3928# VSS 0.04fF $ **FLOATING
C111 ota_v2_without_cmfb_0/li_11121_570# VSS 9.29fF
C112 ota_v2_without_cmfb_0/li_11122_5650# VSS -32.55fF
C113 ota_v2_without_cmfb_0/li_8434_570# VSS 9.00fF
C114 sc_cmfb_0/bias_a VSS -321.62fF
C115 ota_v2_without_cmfb_0/li_8436_5651# VSS 5.90fF
C116 ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VSS -342.20fF
C117 ota_v2_without_cmfb_0/bias_b VSS -361.14fF
C118 ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS 38.05fF
C119 ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VSS 35.85fF
C120 ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VSS 25.03fF
C121 VDD VSS 358.85fF
C122 i_bias VSS -61.81fF
C123 ota_v2_without_cmfb_0/bias_c VSS -128.72fF
C124 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_427# VSS 0.11fF
C125 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_423# VSS 0.11fF
C126 ota_v2_without_cmfb_0/bias_circuit_0/m1_7461_921# VSS 0.12fF
C127 ota_v2_without_cmfb_0/bias_circuit_0/m1_7169_923# VSS 0.13fF
C128 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_433# VSS 0.14fF
C129 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_422# VSS 0.20fF
C130 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_422# VSS 0.20fF
C131 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_1420# VSS 0.12fF
C132 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_1428# VSS 0.12fF
C133 ota_v2_without_cmfb_0/bias_circuit_0/m1_6877_922# VSS 0.14fF
C134 ota_v2_without_cmfb_0/bias_circuit_0/m1_6585_923# VSS 0.22fF
C135 ota_v2_without_cmfb_0/bias_circuit_0/m1_6293_922# VSS 0.16fF
C136 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_1417# VSS 0.13fF
C137 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_1422# VSS 0.22fF
C138 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_1426# VSS 0.22fF
C139 ota_v2_without_cmfb_0/bias_d VSS -236.30fF
C140 ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# VSS 4.65fF
C141 ota_v2_without_cmfb_0/li_14138_570# VSS 33.90fF
C142 sc_cmfb_0/cmc VSS -103.48fF
C143 in VSS -28.56fF
C144 ip VSS -29.73fF
.ends

