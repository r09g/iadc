magic
tech sky130A
magscale 1 2
timestamp 1654647308
<< pwell >>
rect -1146 -1097 1146 1097
<< nmos >>
rect -950 607 -830 887
rect -772 607 -652 887
rect -594 607 -474 887
rect -416 607 -296 887
rect -238 607 -118 887
rect -60 607 60 887
rect 118 607 238 887
rect 296 607 416 887
rect 474 607 594 887
rect 652 607 772 887
rect 830 607 950 887
rect -950 109 -830 389
rect -772 109 -652 389
rect -594 109 -474 389
rect -416 109 -296 389
rect -238 109 -118 389
rect -60 109 60 389
rect 118 109 238 389
rect 296 109 416 389
rect 474 109 594 389
rect 652 109 772 389
rect 830 109 950 389
rect -950 -389 -830 -109
rect -772 -389 -652 -109
rect -594 -389 -474 -109
rect -416 -389 -296 -109
rect -238 -389 -118 -109
rect -60 -389 60 -109
rect 118 -389 238 -109
rect 296 -389 416 -109
rect 474 -389 594 -109
rect 652 -389 772 -109
rect 830 -389 950 -109
rect -950 -887 -830 -607
rect -772 -887 -652 -607
rect -594 -887 -474 -607
rect -416 -887 -296 -607
rect -238 -887 -118 -607
rect -60 -887 60 -607
rect 118 -887 238 -607
rect 296 -887 416 -607
rect 474 -887 594 -607
rect 652 -887 772 -607
rect 830 -887 950 -607
<< ndiff >>
rect -1008 875 -950 887
rect -1008 619 -996 875
rect -962 619 -950 875
rect -1008 607 -950 619
rect -830 875 -772 887
rect -830 619 -818 875
rect -784 619 -772 875
rect -830 607 -772 619
rect -652 875 -594 887
rect -652 619 -640 875
rect -606 619 -594 875
rect -652 607 -594 619
rect -474 875 -416 887
rect -474 619 -462 875
rect -428 619 -416 875
rect -474 607 -416 619
rect -296 875 -238 887
rect -296 619 -284 875
rect -250 619 -238 875
rect -296 607 -238 619
rect -118 875 -60 887
rect -118 619 -106 875
rect -72 619 -60 875
rect -118 607 -60 619
rect 60 875 118 887
rect 60 619 72 875
rect 106 619 118 875
rect 60 607 118 619
rect 238 875 296 887
rect 238 619 250 875
rect 284 619 296 875
rect 238 607 296 619
rect 416 875 474 887
rect 416 619 428 875
rect 462 619 474 875
rect 416 607 474 619
rect 594 875 652 887
rect 594 619 606 875
rect 640 619 652 875
rect 594 607 652 619
rect 772 875 830 887
rect 772 619 784 875
rect 818 619 830 875
rect 772 607 830 619
rect 950 875 1008 887
rect 950 619 962 875
rect 996 619 1008 875
rect 950 607 1008 619
rect -1008 377 -950 389
rect -1008 121 -996 377
rect -962 121 -950 377
rect -1008 109 -950 121
rect -830 377 -772 389
rect -830 121 -818 377
rect -784 121 -772 377
rect -830 109 -772 121
rect -652 377 -594 389
rect -652 121 -640 377
rect -606 121 -594 377
rect -652 109 -594 121
rect -474 377 -416 389
rect -474 121 -462 377
rect -428 121 -416 377
rect -474 109 -416 121
rect -296 377 -238 389
rect -296 121 -284 377
rect -250 121 -238 377
rect -296 109 -238 121
rect -118 377 -60 389
rect -118 121 -106 377
rect -72 121 -60 377
rect -118 109 -60 121
rect 60 377 118 389
rect 60 121 72 377
rect 106 121 118 377
rect 60 109 118 121
rect 238 377 296 389
rect 238 121 250 377
rect 284 121 296 377
rect 238 109 296 121
rect 416 377 474 389
rect 416 121 428 377
rect 462 121 474 377
rect 416 109 474 121
rect 594 377 652 389
rect 594 121 606 377
rect 640 121 652 377
rect 594 109 652 121
rect 772 377 830 389
rect 772 121 784 377
rect 818 121 830 377
rect 772 109 830 121
rect 950 377 1008 389
rect 950 121 962 377
rect 996 121 1008 377
rect 950 109 1008 121
rect -1008 -121 -950 -109
rect -1008 -377 -996 -121
rect -962 -377 -950 -121
rect -1008 -389 -950 -377
rect -830 -121 -772 -109
rect -830 -377 -818 -121
rect -784 -377 -772 -121
rect -830 -389 -772 -377
rect -652 -121 -594 -109
rect -652 -377 -640 -121
rect -606 -377 -594 -121
rect -652 -389 -594 -377
rect -474 -121 -416 -109
rect -474 -377 -462 -121
rect -428 -377 -416 -121
rect -474 -389 -416 -377
rect -296 -121 -238 -109
rect -296 -377 -284 -121
rect -250 -377 -238 -121
rect -296 -389 -238 -377
rect -118 -121 -60 -109
rect -118 -377 -106 -121
rect -72 -377 -60 -121
rect -118 -389 -60 -377
rect 60 -121 118 -109
rect 60 -377 72 -121
rect 106 -377 118 -121
rect 60 -389 118 -377
rect 238 -121 296 -109
rect 238 -377 250 -121
rect 284 -377 296 -121
rect 238 -389 296 -377
rect 416 -121 474 -109
rect 416 -377 428 -121
rect 462 -377 474 -121
rect 416 -389 474 -377
rect 594 -121 652 -109
rect 594 -377 606 -121
rect 640 -377 652 -121
rect 594 -389 652 -377
rect 772 -121 830 -109
rect 772 -377 784 -121
rect 818 -377 830 -121
rect 772 -389 830 -377
rect 950 -121 1008 -109
rect 950 -377 962 -121
rect 996 -377 1008 -121
rect 950 -389 1008 -377
rect -1008 -619 -950 -607
rect -1008 -875 -996 -619
rect -962 -875 -950 -619
rect -1008 -887 -950 -875
rect -830 -619 -772 -607
rect -830 -875 -818 -619
rect -784 -875 -772 -619
rect -830 -887 -772 -875
rect -652 -619 -594 -607
rect -652 -875 -640 -619
rect -606 -875 -594 -619
rect -652 -887 -594 -875
rect -474 -619 -416 -607
rect -474 -875 -462 -619
rect -428 -875 -416 -619
rect -474 -887 -416 -875
rect -296 -619 -238 -607
rect -296 -875 -284 -619
rect -250 -875 -238 -619
rect -296 -887 -238 -875
rect -118 -619 -60 -607
rect -118 -875 -106 -619
rect -72 -875 -60 -619
rect -118 -887 -60 -875
rect 60 -619 118 -607
rect 60 -875 72 -619
rect 106 -875 118 -619
rect 60 -887 118 -875
rect 238 -619 296 -607
rect 238 -875 250 -619
rect 284 -875 296 -619
rect 238 -887 296 -875
rect 416 -619 474 -607
rect 416 -875 428 -619
rect 462 -875 474 -619
rect 416 -887 474 -875
rect 594 -619 652 -607
rect 594 -875 606 -619
rect 640 -875 652 -619
rect 594 -887 652 -875
rect 772 -619 830 -607
rect 772 -875 784 -619
rect 818 -875 830 -619
rect 772 -887 830 -875
rect 950 -619 1008 -607
rect 950 -875 962 -619
rect 996 -875 1008 -619
rect 950 -887 1008 -875
<< ndiffc >>
rect -996 619 -962 875
rect -818 619 -784 875
rect -640 619 -606 875
rect -462 619 -428 875
rect -284 619 -250 875
rect -106 619 -72 875
rect 72 619 106 875
rect 250 619 284 875
rect 428 619 462 875
rect 606 619 640 875
rect 784 619 818 875
rect 962 619 996 875
rect -996 121 -962 377
rect -818 121 -784 377
rect -640 121 -606 377
rect -462 121 -428 377
rect -284 121 -250 377
rect -106 121 -72 377
rect 72 121 106 377
rect 250 121 284 377
rect 428 121 462 377
rect 606 121 640 377
rect 784 121 818 377
rect 962 121 996 377
rect -996 -377 -962 -121
rect -818 -377 -784 -121
rect -640 -377 -606 -121
rect -462 -377 -428 -121
rect -284 -377 -250 -121
rect -106 -377 -72 -121
rect 72 -377 106 -121
rect 250 -377 284 -121
rect 428 -377 462 -121
rect 606 -377 640 -121
rect 784 -377 818 -121
rect 962 -377 996 -121
rect -996 -875 -962 -619
rect -818 -875 -784 -619
rect -640 -875 -606 -619
rect -462 -875 -428 -619
rect -284 -875 -250 -619
rect -106 -875 -72 -619
rect 72 -875 106 -619
rect 250 -875 284 -619
rect 428 -875 462 -619
rect 606 -875 640 -619
rect 784 -875 818 -619
rect 962 -875 996 -619
<< psubdiff >>
rect -1110 1027 -1014 1061
rect 1014 1027 1110 1061
rect -1110 965 -1076 1027
rect 1076 965 1110 1027
rect -1110 -1027 -1076 -965
rect 1076 -1027 1110 -965
rect -1110 -1061 -1014 -1027
rect 1014 -1061 1110 -1027
<< psubdiffcont >>
rect -1014 1027 1014 1061
rect -1110 -965 -1076 965
rect 1076 -965 1110 965
rect -1014 -1061 1014 -1027
<< poly >>
rect -932 959 -848 975
rect -932 942 -916 959
rect -950 925 -916 942
rect -864 942 -848 959
rect -754 959 -670 975
rect -754 942 -738 959
rect -864 925 -830 942
rect -950 887 -830 925
rect -772 925 -738 942
rect -686 942 -670 959
rect -576 959 -492 975
rect -576 942 -560 959
rect -686 925 -652 942
rect -772 887 -652 925
rect -594 925 -560 942
rect -508 942 -492 959
rect -398 959 -314 975
rect -398 942 -382 959
rect -508 925 -474 942
rect -594 887 -474 925
rect -416 925 -382 942
rect -330 942 -314 959
rect -220 959 -136 975
rect -220 942 -204 959
rect -330 925 -296 942
rect -416 887 -296 925
rect -238 925 -204 942
rect -152 942 -136 959
rect -42 959 42 975
rect -42 942 -26 959
rect -152 925 -118 942
rect -238 887 -118 925
rect -60 925 -26 942
rect 26 942 42 959
rect 136 959 220 975
rect 136 942 152 959
rect 26 925 60 942
rect -60 887 60 925
rect 118 925 152 942
rect 204 942 220 959
rect 314 959 398 975
rect 314 942 330 959
rect 204 925 238 942
rect 118 887 238 925
rect 296 925 330 942
rect 382 942 398 959
rect 492 959 576 975
rect 492 942 508 959
rect 382 925 416 942
rect 296 887 416 925
rect 474 925 508 942
rect 560 942 576 959
rect 670 959 754 975
rect 670 942 686 959
rect 560 925 594 942
rect 474 887 594 925
rect 652 925 686 942
rect 738 942 754 959
rect 848 959 932 975
rect 848 942 864 959
rect 738 925 772 942
rect 652 887 772 925
rect 830 925 864 942
rect 916 942 932 959
rect 916 925 950 942
rect 830 887 950 925
rect -950 569 -830 607
rect -950 552 -916 569
rect -932 535 -916 552
rect -864 552 -830 569
rect -772 569 -652 607
rect -772 552 -738 569
rect -864 535 -848 552
rect -932 519 -848 535
rect -754 535 -738 552
rect -686 552 -652 569
rect -594 569 -474 607
rect -594 552 -560 569
rect -686 535 -670 552
rect -754 519 -670 535
rect -576 535 -560 552
rect -508 552 -474 569
rect -416 569 -296 607
rect -416 552 -382 569
rect -508 535 -492 552
rect -576 519 -492 535
rect -398 535 -382 552
rect -330 552 -296 569
rect -238 569 -118 607
rect -238 552 -204 569
rect -330 535 -314 552
rect -398 519 -314 535
rect -220 535 -204 552
rect -152 552 -118 569
rect -60 569 60 607
rect -60 552 -26 569
rect -152 535 -136 552
rect -220 519 -136 535
rect -42 535 -26 552
rect 26 552 60 569
rect 118 569 238 607
rect 118 552 152 569
rect 26 535 42 552
rect -42 519 42 535
rect 136 535 152 552
rect 204 552 238 569
rect 296 569 416 607
rect 296 552 330 569
rect 204 535 220 552
rect 136 519 220 535
rect 314 535 330 552
rect 382 552 416 569
rect 474 569 594 607
rect 474 552 508 569
rect 382 535 398 552
rect 314 519 398 535
rect 492 535 508 552
rect 560 552 594 569
rect 652 569 772 607
rect 652 552 686 569
rect 560 535 576 552
rect 492 519 576 535
rect 670 535 686 552
rect 738 552 772 569
rect 830 569 950 607
rect 830 552 864 569
rect 738 535 754 552
rect 670 519 754 535
rect 848 535 864 552
rect 916 552 950 569
rect 916 535 932 552
rect 848 519 932 535
rect -932 461 -848 477
rect -932 444 -916 461
rect -950 427 -916 444
rect -864 444 -848 461
rect -754 461 -670 477
rect -754 444 -738 461
rect -864 427 -830 444
rect -950 389 -830 427
rect -772 427 -738 444
rect -686 444 -670 461
rect -576 461 -492 477
rect -576 444 -560 461
rect -686 427 -652 444
rect -772 389 -652 427
rect -594 427 -560 444
rect -508 444 -492 461
rect -398 461 -314 477
rect -398 444 -382 461
rect -508 427 -474 444
rect -594 389 -474 427
rect -416 427 -382 444
rect -330 444 -314 461
rect -220 461 -136 477
rect -220 444 -204 461
rect -330 427 -296 444
rect -416 389 -296 427
rect -238 427 -204 444
rect -152 444 -136 461
rect -42 461 42 477
rect -42 444 -26 461
rect -152 427 -118 444
rect -238 389 -118 427
rect -60 427 -26 444
rect 26 444 42 461
rect 136 461 220 477
rect 136 444 152 461
rect 26 427 60 444
rect -60 389 60 427
rect 118 427 152 444
rect 204 444 220 461
rect 314 461 398 477
rect 314 444 330 461
rect 204 427 238 444
rect 118 389 238 427
rect 296 427 330 444
rect 382 444 398 461
rect 492 461 576 477
rect 492 444 508 461
rect 382 427 416 444
rect 296 389 416 427
rect 474 427 508 444
rect 560 444 576 461
rect 670 461 754 477
rect 670 444 686 461
rect 560 427 594 444
rect 474 389 594 427
rect 652 427 686 444
rect 738 444 754 461
rect 848 461 932 477
rect 848 444 864 461
rect 738 427 772 444
rect 652 389 772 427
rect 830 427 864 444
rect 916 444 932 461
rect 916 427 950 444
rect 830 389 950 427
rect -950 71 -830 109
rect -950 54 -916 71
rect -932 37 -916 54
rect -864 54 -830 71
rect -772 71 -652 109
rect -772 54 -738 71
rect -864 37 -848 54
rect -932 21 -848 37
rect -754 37 -738 54
rect -686 54 -652 71
rect -594 71 -474 109
rect -594 54 -560 71
rect -686 37 -670 54
rect -754 21 -670 37
rect -576 37 -560 54
rect -508 54 -474 71
rect -416 71 -296 109
rect -416 54 -382 71
rect -508 37 -492 54
rect -576 21 -492 37
rect -398 37 -382 54
rect -330 54 -296 71
rect -238 71 -118 109
rect -238 54 -204 71
rect -330 37 -314 54
rect -398 21 -314 37
rect -220 37 -204 54
rect -152 54 -118 71
rect -60 71 60 109
rect -60 54 -26 71
rect -152 37 -136 54
rect -220 21 -136 37
rect -42 37 -26 54
rect 26 54 60 71
rect 118 71 238 109
rect 118 54 152 71
rect 26 37 42 54
rect -42 21 42 37
rect 136 37 152 54
rect 204 54 238 71
rect 296 71 416 109
rect 296 54 330 71
rect 204 37 220 54
rect 136 21 220 37
rect 314 37 330 54
rect 382 54 416 71
rect 474 71 594 109
rect 474 54 508 71
rect 382 37 398 54
rect 314 21 398 37
rect 492 37 508 54
rect 560 54 594 71
rect 652 71 772 109
rect 652 54 686 71
rect 560 37 576 54
rect 492 21 576 37
rect 670 37 686 54
rect 738 54 772 71
rect 830 71 950 109
rect 830 54 864 71
rect 738 37 754 54
rect 670 21 754 37
rect 848 37 864 54
rect 916 54 950 71
rect 916 37 932 54
rect 848 21 932 37
rect -932 -37 -848 -21
rect -932 -54 -916 -37
rect -950 -71 -916 -54
rect -864 -54 -848 -37
rect -754 -37 -670 -21
rect -754 -54 -738 -37
rect -864 -71 -830 -54
rect -950 -109 -830 -71
rect -772 -71 -738 -54
rect -686 -54 -670 -37
rect -576 -37 -492 -21
rect -576 -54 -560 -37
rect -686 -71 -652 -54
rect -772 -109 -652 -71
rect -594 -71 -560 -54
rect -508 -54 -492 -37
rect -398 -37 -314 -21
rect -398 -54 -382 -37
rect -508 -71 -474 -54
rect -594 -109 -474 -71
rect -416 -71 -382 -54
rect -330 -54 -314 -37
rect -220 -37 -136 -21
rect -220 -54 -204 -37
rect -330 -71 -296 -54
rect -416 -109 -296 -71
rect -238 -71 -204 -54
rect -152 -54 -136 -37
rect -42 -37 42 -21
rect -42 -54 -26 -37
rect -152 -71 -118 -54
rect -238 -109 -118 -71
rect -60 -71 -26 -54
rect 26 -54 42 -37
rect 136 -37 220 -21
rect 136 -54 152 -37
rect 26 -71 60 -54
rect -60 -109 60 -71
rect 118 -71 152 -54
rect 204 -54 220 -37
rect 314 -37 398 -21
rect 314 -54 330 -37
rect 204 -71 238 -54
rect 118 -109 238 -71
rect 296 -71 330 -54
rect 382 -54 398 -37
rect 492 -37 576 -21
rect 492 -54 508 -37
rect 382 -71 416 -54
rect 296 -109 416 -71
rect 474 -71 508 -54
rect 560 -54 576 -37
rect 670 -37 754 -21
rect 670 -54 686 -37
rect 560 -71 594 -54
rect 474 -109 594 -71
rect 652 -71 686 -54
rect 738 -54 754 -37
rect 848 -37 932 -21
rect 848 -54 864 -37
rect 738 -71 772 -54
rect 652 -109 772 -71
rect 830 -71 864 -54
rect 916 -54 932 -37
rect 916 -71 950 -54
rect 830 -109 950 -71
rect -950 -427 -830 -389
rect -950 -444 -916 -427
rect -932 -461 -916 -444
rect -864 -444 -830 -427
rect -772 -427 -652 -389
rect -772 -444 -738 -427
rect -864 -461 -848 -444
rect -932 -477 -848 -461
rect -754 -461 -738 -444
rect -686 -444 -652 -427
rect -594 -427 -474 -389
rect -594 -444 -560 -427
rect -686 -461 -670 -444
rect -754 -477 -670 -461
rect -576 -461 -560 -444
rect -508 -444 -474 -427
rect -416 -427 -296 -389
rect -416 -444 -382 -427
rect -508 -461 -492 -444
rect -576 -477 -492 -461
rect -398 -461 -382 -444
rect -330 -444 -296 -427
rect -238 -427 -118 -389
rect -238 -444 -204 -427
rect -330 -461 -314 -444
rect -398 -477 -314 -461
rect -220 -461 -204 -444
rect -152 -444 -118 -427
rect -60 -427 60 -389
rect -60 -444 -26 -427
rect -152 -461 -136 -444
rect -220 -477 -136 -461
rect -42 -461 -26 -444
rect 26 -444 60 -427
rect 118 -427 238 -389
rect 118 -444 152 -427
rect 26 -461 42 -444
rect -42 -477 42 -461
rect 136 -461 152 -444
rect 204 -444 238 -427
rect 296 -427 416 -389
rect 296 -444 330 -427
rect 204 -461 220 -444
rect 136 -477 220 -461
rect 314 -461 330 -444
rect 382 -444 416 -427
rect 474 -427 594 -389
rect 474 -444 508 -427
rect 382 -461 398 -444
rect 314 -477 398 -461
rect 492 -461 508 -444
rect 560 -444 594 -427
rect 652 -427 772 -389
rect 652 -444 686 -427
rect 560 -461 576 -444
rect 492 -477 576 -461
rect 670 -461 686 -444
rect 738 -444 772 -427
rect 830 -427 950 -389
rect 830 -444 864 -427
rect 738 -461 754 -444
rect 670 -477 754 -461
rect 848 -461 864 -444
rect 916 -444 950 -427
rect 916 -461 932 -444
rect 848 -477 932 -461
rect -932 -535 -848 -519
rect -932 -552 -916 -535
rect -950 -569 -916 -552
rect -864 -552 -848 -535
rect -754 -535 -670 -519
rect -754 -552 -738 -535
rect -864 -569 -830 -552
rect -950 -607 -830 -569
rect -772 -569 -738 -552
rect -686 -552 -670 -535
rect -576 -535 -492 -519
rect -576 -552 -560 -535
rect -686 -569 -652 -552
rect -772 -607 -652 -569
rect -594 -569 -560 -552
rect -508 -552 -492 -535
rect -398 -535 -314 -519
rect -398 -552 -382 -535
rect -508 -569 -474 -552
rect -594 -607 -474 -569
rect -416 -569 -382 -552
rect -330 -552 -314 -535
rect -220 -535 -136 -519
rect -220 -552 -204 -535
rect -330 -569 -296 -552
rect -416 -607 -296 -569
rect -238 -569 -204 -552
rect -152 -552 -136 -535
rect -42 -535 42 -519
rect -42 -552 -26 -535
rect -152 -569 -118 -552
rect -238 -607 -118 -569
rect -60 -569 -26 -552
rect 26 -552 42 -535
rect 136 -535 220 -519
rect 136 -552 152 -535
rect 26 -569 60 -552
rect -60 -607 60 -569
rect 118 -569 152 -552
rect 204 -552 220 -535
rect 314 -535 398 -519
rect 314 -552 330 -535
rect 204 -569 238 -552
rect 118 -607 238 -569
rect 296 -569 330 -552
rect 382 -552 398 -535
rect 492 -535 576 -519
rect 492 -552 508 -535
rect 382 -569 416 -552
rect 296 -607 416 -569
rect 474 -569 508 -552
rect 560 -552 576 -535
rect 670 -535 754 -519
rect 670 -552 686 -535
rect 560 -569 594 -552
rect 474 -607 594 -569
rect 652 -569 686 -552
rect 738 -552 754 -535
rect 848 -535 932 -519
rect 848 -552 864 -535
rect 738 -569 772 -552
rect 652 -607 772 -569
rect 830 -569 864 -552
rect 916 -552 932 -535
rect 916 -569 950 -552
rect 830 -607 950 -569
rect -950 -925 -830 -887
rect -950 -942 -916 -925
rect -932 -959 -916 -942
rect -864 -942 -830 -925
rect -772 -925 -652 -887
rect -772 -942 -738 -925
rect -864 -959 -848 -942
rect -932 -975 -848 -959
rect -754 -959 -738 -942
rect -686 -942 -652 -925
rect -594 -925 -474 -887
rect -594 -942 -560 -925
rect -686 -959 -670 -942
rect -754 -975 -670 -959
rect -576 -959 -560 -942
rect -508 -942 -474 -925
rect -416 -925 -296 -887
rect -416 -942 -382 -925
rect -508 -959 -492 -942
rect -576 -975 -492 -959
rect -398 -959 -382 -942
rect -330 -942 -296 -925
rect -238 -925 -118 -887
rect -238 -942 -204 -925
rect -330 -959 -314 -942
rect -398 -975 -314 -959
rect -220 -959 -204 -942
rect -152 -942 -118 -925
rect -60 -925 60 -887
rect -60 -942 -26 -925
rect -152 -959 -136 -942
rect -220 -975 -136 -959
rect -42 -959 -26 -942
rect 26 -942 60 -925
rect 118 -925 238 -887
rect 118 -942 152 -925
rect 26 -959 42 -942
rect -42 -975 42 -959
rect 136 -959 152 -942
rect 204 -942 238 -925
rect 296 -925 416 -887
rect 296 -942 330 -925
rect 204 -959 220 -942
rect 136 -975 220 -959
rect 314 -959 330 -942
rect 382 -942 416 -925
rect 474 -925 594 -887
rect 474 -942 508 -925
rect 382 -959 398 -942
rect 314 -975 398 -959
rect 492 -959 508 -942
rect 560 -942 594 -925
rect 652 -925 772 -887
rect 652 -942 686 -925
rect 560 -959 576 -942
rect 492 -975 576 -959
rect 670 -959 686 -942
rect 738 -942 772 -925
rect 830 -925 950 -887
rect 830 -942 864 -925
rect 738 -959 754 -942
rect 670 -975 754 -959
rect 848 -959 864 -942
rect 916 -942 950 -925
rect 916 -959 932 -942
rect 848 -975 932 -959
<< polycont >>
rect -916 925 -864 959
rect -738 925 -686 959
rect -560 925 -508 959
rect -382 925 -330 959
rect -204 925 -152 959
rect -26 925 26 959
rect 152 925 204 959
rect 330 925 382 959
rect 508 925 560 959
rect 686 925 738 959
rect 864 925 916 959
rect -916 535 -864 569
rect -738 535 -686 569
rect -560 535 -508 569
rect -382 535 -330 569
rect -204 535 -152 569
rect -26 535 26 569
rect 152 535 204 569
rect 330 535 382 569
rect 508 535 560 569
rect 686 535 738 569
rect 864 535 916 569
rect -916 427 -864 461
rect -738 427 -686 461
rect -560 427 -508 461
rect -382 427 -330 461
rect -204 427 -152 461
rect -26 427 26 461
rect 152 427 204 461
rect 330 427 382 461
rect 508 427 560 461
rect 686 427 738 461
rect 864 427 916 461
rect -916 37 -864 71
rect -738 37 -686 71
rect -560 37 -508 71
rect -382 37 -330 71
rect -204 37 -152 71
rect -26 37 26 71
rect 152 37 204 71
rect 330 37 382 71
rect 508 37 560 71
rect 686 37 738 71
rect 864 37 916 71
rect -916 -71 -864 -37
rect -738 -71 -686 -37
rect -560 -71 -508 -37
rect -382 -71 -330 -37
rect -204 -71 -152 -37
rect -26 -71 26 -37
rect 152 -71 204 -37
rect 330 -71 382 -37
rect 508 -71 560 -37
rect 686 -71 738 -37
rect 864 -71 916 -37
rect -916 -461 -864 -427
rect -738 -461 -686 -427
rect -560 -461 -508 -427
rect -382 -461 -330 -427
rect -204 -461 -152 -427
rect -26 -461 26 -427
rect 152 -461 204 -427
rect 330 -461 382 -427
rect 508 -461 560 -427
rect 686 -461 738 -427
rect 864 -461 916 -427
rect -916 -569 -864 -535
rect -738 -569 -686 -535
rect -560 -569 -508 -535
rect -382 -569 -330 -535
rect -204 -569 -152 -535
rect -26 -569 26 -535
rect 152 -569 204 -535
rect 330 -569 382 -535
rect 508 -569 560 -535
rect 686 -569 738 -535
rect 864 -569 916 -535
rect -916 -959 -864 -925
rect -738 -959 -686 -925
rect -560 -959 -508 -925
rect -382 -959 -330 -925
rect -204 -959 -152 -925
rect -26 -959 26 -925
rect 152 -959 204 -925
rect 330 -959 382 -925
rect 508 -959 560 -925
rect 686 -959 738 -925
rect 864 -959 916 -925
<< locali >>
rect -1110 1027 -1014 1061
rect 1014 1027 1110 1061
rect -1110 965 -1076 1027
rect 1076 965 1110 1027
rect -1076 925 -916 959
rect -864 925 -848 959
rect -754 925 -738 959
rect -686 925 -670 959
rect -576 925 -560 959
rect -508 925 -492 959
rect -398 925 -382 959
rect -330 925 -314 959
rect -220 925 -204 959
rect -152 925 -136 959
rect -42 925 -26 959
rect 26 925 42 959
rect 136 925 152 959
rect 204 925 220 959
rect 314 925 330 959
rect 382 925 398 959
rect 492 925 508 959
rect 560 925 576 959
rect 670 925 686 959
rect 738 925 754 959
rect 848 925 864 959
rect 916 925 1076 959
rect -996 875 -962 925
rect -996 569 -962 619
rect -818 875 -784 891
rect -818 603 -784 619
rect -640 875 -606 891
rect -640 603 -606 619
rect -462 875 -428 891
rect -462 603 -428 619
rect -284 875 -250 891
rect -284 603 -250 619
rect -106 875 -72 891
rect -106 603 -72 619
rect 72 875 106 891
rect 72 603 106 619
rect 250 875 284 891
rect 250 603 284 619
rect 428 875 462 891
rect 428 603 462 619
rect 606 875 640 891
rect 606 603 640 619
rect 784 875 818 891
rect 784 603 818 619
rect 962 875 996 925
rect 962 569 996 619
rect -1076 535 -916 569
rect -864 535 -848 569
rect -754 535 -738 569
rect -686 535 -670 569
rect -576 535 -560 569
rect -508 535 -492 569
rect -398 535 -382 569
rect -330 535 -314 569
rect -220 535 -204 569
rect -152 535 -136 569
rect -42 535 -26 569
rect 26 535 42 569
rect 136 535 152 569
rect 204 535 220 569
rect 314 535 330 569
rect 382 535 398 569
rect 492 535 508 569
rect 560 535 576 569
rect 670 535 686 569
rect 738 535 754 569
rect 848 535 864 569
rect 916 535 1076 569
rect -1076 427 -916 461
rect -864 427 -848 461
rect -754 427 -738 461
rect -686 427 -670 461
rect -576 427 -560 461
rect -508 427 -492 461
rect -398 427 -382 461
rect -330 427 -314 461
rect -220 427 -204 461
rect -152 427 -136 461
rect -42 427 -26 461
rect 26 427 42 461
rect 136 427 152 461
rect 204 427 220 461
rect 314 427 330 461
rect 382 427 398 461
rect 492 427 508 461
rect 560 427 576 461
rect 670 427 686 461
rect 738 427 754 461
rect 848 427 864 461
rect 916 427 1076 461
rect -996 377 -962 427
rect -996 71 -962 121
rect -818 377 -784 393
rect -818 105 -784 121
rect -640 377 -606 393
rect -640 105 -606 121
rect -462 377 -428 393
rect -462 105 -428 121
rect -284 377 -250 393
rect -284 105 -250 121
rect -106 377 -72 393
rect -106 105 -72 121
rect 72 377 106 393
rect 72 105 106 121
rect 250 377 284 393
rect 250 105 284 121
rect 428 377 462 393
rect 428 105 462 121
rect 606 377 640 393
rect 606 105 640 121
rect 784 377 818 393
rect 784 105 818 121
rect 962 377 996 427
rect 962 71 996 121
rect -1076 37 -916 71
rect -864 37 -848 71
rect -754 37 -738 71
rect -686 37 -670 71
rect -576 37 -560 71
rect -508 37 -492 71
rect -398 37 -382 71
rect -330 37 -314 71
rect -220 37 -204 71
rect -152 37 -136 71
rect -42 37 -26 71
rect 26 37 42 71
rect 136 37 152 71
rect 204 37 220 71
rect 314 37 330 71
rect 382 37 398 71
rect 492 37 508 71
rect 560 37 576 71
rect 670 37 686 71
rect 738 37 754 71
rect 848 37 864 71
rect 916 37 1076 71
rect -1076 -71 -916 -37
rect -864 -71 -848 -37
rect -754 -71 -738 -37
rect -686 -71 -670 -37
rect -576 -71 -560 -37
rect -508 -71 -492 -37
rect -398 -71 -382 -37
rect -330 -71 -314 -37
rect -220 -71 -204 -37
rect -152 -71 -136 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 136 -71 152 -37
rect 204 -71 220 -37
rect 314 -71 330 -37
rect 382 -71 398 -37
rect 492 -71 508 -37
rect 560 -71 576 -37
rect 670 -71 686 -37
rect 738 -71 754 -37
rect 848 -71 864 -37
rect 916 -71 1076 -37
rect -996 -121 -962 -71
rect -996 -427 -962 -377
rect -818 -121 -784 -105
rect -818 -393 -784 -377
rect -640 -121 -606 -105
rect -640 -393 -606 -377
rect -462 -121 -428 -105
rect -462 -393 -428 -377
rect -284 -121 -250 -105
rect -284 -393 -250 -377
rect -106 -121 -72 -105
rect -106 -393 -72 -377
rect 72 -121 106 -105
rect 72 -393 106 -377
rect 250 -121 284 -105
rect 250 -393 284 -377
rect 428 -121 462 -105
rect 428 -393 462 -377
rect 606 -121 640 -105
rect 606 -393 640 -377
rect 784 -121 818 -105
rect 784 -393 818 -377
rect 962 -121 996 -71
rect 962 -427 996 -377
rect -1076 -461 -916 -427
rect -864 -461 -848 -427
rect -754 -461 -738 -427
rect -686 -461 -670 -427
rect -576 -461 -560 -427
rect -508 -461 -492 -427
rect -398 -461 -382 -427
rect -330 -461 -314 -427
rect -220 -461 -204 -427
rect -152 -461 -136 -427
rect -42 -461 -26 -427
rect 26 -461 42 -427
rect 136 -461 152 -427
rect 204 -461 220 -427
rect 314 -461 330 -427
rect 382 -461 398 -427
rect 492 -461 508 -427
rect 560 -461 576 -427
rect 670 -461 686 -427
rect 738 -461 754 -427
rect 848 -461 864 -427
rect 916 -461 1076 -427
rect -1076 -569 -916 -535
rect -864 -569 -848 -535
rect -754 -569 -738 -535
rect -686 -569 -670 -535
rect -576 -569 -560 -535
rect -508 -569 -492 -535
rect -398 -569 -382 -535
rect -330 -569 -314 -535
rect -220 -569 -204 -535
rect -152 -569 -136 -535
rect -42 -569 -26 -535
rect 26 -569 42 -535
rect 136 -569 152 -535
rect 204 -569 220 -535
rect 314 -569 330 -535
rect 382 -569 398 -535
rect 492 -569 508 -535
rect 560 -569 576 -535
rect 670 -569 686 -535
rect 738 -569 754 -535
rect 848 -569 864 -535
rect 916 -569 1076 -535
rect -996 -619 -962 -569
rect -996 -925 -962 -875
rect -818 -619 -784 -603
rect -818 -891 -784 -875
rect -640 -619 -606 -603
rect -640 -891 -606 -875
rect -462 -619 -428 -603
rect -462 -891 -428 -875
rect -284 -619 -250 -603
rect -284 -891 -250 -875
rect -106 -619 -72 -603
rect -106 -891 -72 -875
rect 72 -619 106 -603
rect 72 -891 106 -875
rect 250 -619 284 -603
rect 250 -891 284 -875
rect 428 -619 462 -603
rect 428 -891 462 -875
rect 606 -619 640 -603
rect 606 -891 640 -875
rect 784 -619 818 -603
rect 784 -891 818 -875
rect 962 -619 996 -569
rect 962 -925 996 -875
rect -1076 -959 -916 -925
rect -864 -959 -848 -925
rect -754 -959 -738 -925
rect -686 -959 -670 -925
rect -576 -959 -560 -925
rect -508 -959 -492 -925
rect -398 -959 -382 -925
rect -330 -959 -314 -925
rect -220 -959 -204 -925
rect -152 -959 -136 -925
rect -42 -959 -26 -925
rect 26 -959 42 -925
rect 136 -959 152 -925
rect 204 -959 220 -925
rect 314 -959 330 -925
rect 382 -959 398 -925
rect 492 -959 508 -925
rect 560 -959 576 -925
rect 670 -959 686 -925
rect 738 -959 754 -925
rect 848 -959 864 -925
rect 916 -959 1076 -925
rect -1110 -1027 -1076 -965
rect 1076 -1027 1110 -965
rect -1110 -1061 -1014 -1027
rect 1014 -1061 1110 -1027
<< viali >>
rect -738 925 -686 959
rect -560 925 -508 959
rect -382 925 -330 959
rect -204 925 -152 959
rect -26 925 26 959
rect 152 925 204 959
rect 330 925 382 959
rect 508 925 560 959
rect 686 925 738 959
rect -738 535 -686 569
rect -560 535 -508 569
rect -382 535 -330 569
rect -204 535 -152 569
rect -26 535 26 569
rect 152 535 204 569
rect 330 535 382 569
rect 508 535 560 569
rect 686 535 738 569
rect -738 427 -686 461
rect -560 427 -508 461
rect -382 427 -330 461
rect -204 427 -152 461
rect -26 427 26 461
rect 152 427 204 461
rect 330 427 382 461
rect 508 427 560 461
rect 686 427 738 461
rect -738 37 -686 71
rect -560 37 -508 71
rect -382 37 -330 71
rect -204 37 -152 71
rect -26 37 26 71
rect 152 37 204 71
rect 330 37 382 71
rect 508 37 560 71
rect 686 37 738 71
rect -738 -71 -686 -37
rect -560 -71 -508 -37
rect -382 -71 -330 -37
rect -204 -71 -152 -37
rect -26 -71 26 -37
rect 152 -71 204 -37
rect 330 -71 382 -37
rect 508 -71 560 -37
rect 686 -71 738 -37
rect -738 -461 -686 -427
rect -560 -461 -508 -427
rect -382 -461 -330 -427
rect -204 -461 -152 -427
rect -26 -461 26 -427
rect 152 -461 204 -427
rect 330 -461 382 -427
rect 508 -461 560 -427
rect 686 -461 738 -427
rect -738 -569 -686 -535
rect -560 -569 -508 -535
rect -382 -569 -330 -535
rect -204 -569 -152 -535
rect -26 -569 26 -535
rect 152 -569 204 -535
rect 330 -569 382 -535
rect 508 -569 560 -535
rect 686 -569 738 -535
rect -738 -959 -686 -925
rect -560 -959 -508 -925
rect -382 -959 -330 -925
rect -204 -959 -152 -925
rect -26 -959 26 -925
rect 152 -959 204 -925
rect 330 -959 382 -925
rect 508 -959 560 -925
rect 686 -959 738 -925
<< metal1 >>
rect -750 959 -674 965
rect -750 925 -738 959
rect -686 925 -674 959
rect -750 919 -674 925
rect -572 959 -496 965
rect -572 925 -560 959
rect -508 925 -496 959
rect -572 919 -496 925
rect -394 959 -318 965
rect -394 925 -382 959
rect -330 925 -318 959
rect -394 919 -318 925
rect -216 959 -140 965
rect -216 925 -204 959
rect -152 925 -140 959
rect -216 919 -140 925
rect -38 959 38 965
rect -38 925 -26 959
rect 26 925 38 959
rect -38 919 38 925
rect 140 959 216 965
rect 140 925 152 959
rect 204 925 216 959
rect 140 919 216 925
rect 318 959 394 965
rect 318 925 330 959
rect 382 925 394 959
rect 318 919 394 925
rect 496 959 572 965
rect 496 925 508 959
rect 560 925 572 959
rect 496 919 572 925
rect 674 959 750 965
rect 674 925 686 959
rect 738 925 750 959
rect 674 919 750 925
rect -750 569 -674 575
rect -750 535 -738 569
rect -686 535 -674 569
rect -750 529 -674 535
rect -572 569 -496 575
rect -572 535 -560 569
rect -508 535 -496 569
rect -572 529 -496 535
rect -394 569 -318 575
rect -394 535 -382 569
rect -330 535 -318 569
rect -394 529 -318 535
rect -216 569 -140 575
rect -216 535 -204 569
rect -152 535 -140 569
rect -216 529 -140 535
rect -38 569 38 575
rect -38 535 -26 569
rect 26 535 38 569
rect -38 529 38 535
rect 140 569 216 575
rect 140 535 152 569
rect 204 535 216 569
rect 140 529 216 535
rect 318 569 394 575
rect 318 535 330 569
rect 382 535 394 569
rect 318 529 394 535
rect 496 569 572 575
rect 496 535 508 569
rect 560 535 572 569
rect 496 529 572 535
rect 674 569 750 575
rect 674 535 686 569
rect 738 535 750 569
rect 674 529 750 535
rect -750 461 -674 467
rect -750 427 -738 461
rect -686 427 -674 461
rect -750 421 -674 427
rect -572 461 -496 467
rect -572 427 -560 461
rect -508 427 -496 461
rect -572 421 -496 427
rect -394 461 -318 467
rect -394 427 -382 461
rect -330 427 -318 461
rect -394 421 -318 427
rect -216 461 -140 467
rect -216 427 -204 461
rect -152 427 -140 461
rect -216 421 -140 427
rect -38 461 38 467
rect -38 427 -26 461
rect 26 427 38 461
rect -38 421 38 427
rect 140 461 216 467
rect 140 427 152 461
rect 204 427 216 461
rect 140 421 216 427
rect 318 461 394 467
rect 318 427 330 461
rect 382 427 394 461
rect 318 421 394 427
rect 496 461 572 467
rect 496 427 508 461
rect 560 427 572 461
rect 496 421 572 427
rect 674 461 750 467
rect 674 427 686 461
rect 738 427 750 461
rect 674 421 750 427
rect -750 71 -674 77
rect -750 37 -738 71
rect -686 37 -674 71
rect -750 31 -674 37
rect -572 71 -496 77
rect -572 37 -560 71
rect -508 37 -496 71
rect -572 31 -496 37
rect -394 71 -318 77
rect -394 37 -382 71
rect -330 37 -318 71
rect -394 31 -318 37
rect -216 71 -140 77
rect -216 37 -204 71
rect -152 37 -140 71
rect -216 31 -140 37
rect -38 71 38 77
rect -38 37 -26 71
rect 26 37 38 71
rect -38 31 38 37
rect 140 71 216 77
rect 140 37 152 71
rect 204 37 216 71
rect 140 31 216 37
rect 318 71 394 77
rect 318 37 330 71
rect 382 37 394 71
rect 318 31 394 37
rect 496 71 572 77
rect 496 37 508 71
rect 560 37 572 71
rect 496 31 572 37
rect 674 71 750 77
rect 674 37 686 71
rect 738 37 750 71
rect 674 31 750 37
rect -750 -37 -674 -31
rect -750 -71 -738 -37
rect -686 -71 -674 -37
rect -750 -77 -674 -71
rect -572 -37 -496 -31
rect -572 -71 -560 -37
rect -508 -71 -496 -37
rect -572 -77 -496 -71
rect -394 -37 -318 -31
rect -394 -71 -382 -37
rect -330 -71 -318 -37
rect -394 -77 -318 -71
rect -216 -37 -140 -31
rect -216 -71 -204 -37
rect -152 -71 -140 -37
rect -216 -77 -140 -71
rect -38 -37 38 -31
rect -38 -71 -26 -37
rect 26 -71 38 -37
rect -38 -77 38 -71
rect 140 -37 216 -31
rect 140 -71 152 -37
rect 204 -71 216 -37
rect 140 -77 216 -71
rect 318 -37 394 -31
rect 318 -71 330 -37
rect 382 -71 394 -37
rect 318 -77 394 -71
rect 496 -37 572 -31
rect 496 -71 508 -37
rect 560 -71 572 -37
rect 496 -77 572 -71
rect 674 -37 750 -31
rect 674 -71 686 -37
rect 738 -71 750 -37
rect 674 -77 750 -71
rect -750 -427 -674 -421
rect -750 -461 -738 -427
rect -686 -461 -674 -427
rect -750 -467 -674 -461
rect -572 -427 -496 -421
rect -572 -461 -560 -427
rect -508 -461 -496 -427
rect -572 -467 -496 -461
rect -394 -427 -318 -421
rect -394 -461 -382 -427
rect -330 -461 -318 -427
rect -394 -467 -318 -461
rect -216 -427 -140 -421
rect -216 -461 -204 -427
rect -152 -461 -140 -427
rect -216 -467 -140 -461
rect -38 -427 38 -421
rect -38 -461 -26 -427
rect 26 -461 38 -427
rect -38 -467 38 -461
rect 140 -427 216 -421
rect 140 -461 152 -427
rect 204 -461 216 -427
rect 140 -467 216 -461
rect 318 -427 394 -421
rect 318 -461 330 -427
rect 382 -461 394 -427
rect 318 -467 394 -461
rect 496 -427 572 -421
rect 496 -461 508 -427
rect 560 -461 572 -427
rect 496 -467 572 -461
rect 674 -427 750 -421
rect 674 -461 686 -427
rect 738 -461 750 -427
rect 674 -467 750 -461
rect -750 -535 -674 -529
rect -750 -569 -738 -535
rect -686 -569 -674 -535
rect -750 -575 -674 -569
rect -572 -535 -496 -529
rect -572 -569 -560 -535
rect -508 -569 -496 -535
rect -572 -575 -496 -569
rect -394 -535 -318 -529
rect -394 -569 -382 -535
rect -330 -569 -318 -535
rect -394 -575 -318 -569
rect -216 -535 -140 -529
rect -216 -569 -204 -535
rect -152 -569 -140 -535
rect -216 -575 -140 -569
rect -38 -535 38 -529
rect -38 -569 -26 -535
rect 26 -569 38 -535
rect -38 -575 38 -569
rect 140 -535 216 -529
rect 140 -569 152 -535
rect 204 -569 216 -535
rect 140 -575 216 -569
rect 318 -535 394 -529
rect 318 -569 330 -535
rect 382 -569 394 -535
rect 318 -575 394 -569
rect 496 -535 572 -529
rect 496 -569 508 -535
rect 560 -569 572 -535
rect 496 -575 572 -569
rect 674 -535 750 -529
rect 674 -569 686 -535
rect 738 -569 750 -535
rect 674 -575 750 -569
rect -750 -925 -674 -919
rect -750 -959 -738 -925
rect -686 -959 -674 -925
rect -750 -965 -674 -959
rect -572 -925 -496 -919
rect -572 -959 -560 -925
rect -508 -959 -496 -925
rect -572 -965 -496 -959
rect -394 -925 -318 -919
rect -394 -959 -382 -925
rect -330 -959 -318 -925
rect -394 -965 -318 -959
rect -216 -925 -140 -919
rect -216 -959 -204 -925
rect -152 -959 -140 -925
rect -216 -965 -140 -959
rect -38 -925 38 -919
rect -38 -959 -26 -925
rect 26 -959 38 -925
rect -38 -965 38 -959
rect 140 -925 216 -919
rect 140 -959 152 -925
rect 204 -959 216 -925
rect 140 -965 216 -959
rect 318 -925 394 -919
rect 318 -959 330 -925
rect 382 -959 394 -925
rect 318 -965 394 -959
rect 496 -925 572 -919
rect 496 -959 508 -925
rect 560 -959 572 -925
rect 496 -965 572 -959
rect 674 -925 750 -919
rect 674 -959 686 -925
rect 738 -959 750 -925
rect 674 -965 750 -959
<< properties >>
string FIXED_BBOX -1093 -1044 1093 1044
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 4 nf 11 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
