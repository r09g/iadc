magic
tech sky130A
magscale 1 2
timestamp 1654727055
<< nwell >>
rect -3788 8059 -3150 8060
rect 1443 8059 2009 10671
rect 6612 8059 7250 8060
rect -3788 6889 7250 8059
rect -3788 6888 6246 6889
rect -3788 6887 -2673 6888
rect -3788 5650 -3150 6887
rect -3788 5635 -3148 5650
rect -3786 3588 -3148 5635
rect 6612 3588 7250 6889
<< pwell >>
rect 1203 10604 1385 10632
rect 1165 10570 1385 10604
rect 1203 9530 1385 10570
rect 1230 9526 1385 9530
rect 1220 9440 1385 9526
rect 1230 9436 1385 9440
rect 1203 9407 1385 9436
rect 1165 9373 1385 9407
rect 1203 9003 1385 9373
rect 1203 8939 1393 9003
rect 1203 8304 1385 8939
rect 1165 8270 1385 8304
rect 1203 8242 1385 8270
rect 2067 9592 2249 10632
rect 2067 9558 2287 9592
rect 2067 9407 2249 9558
rect 2067 9373 2287 9407
rect 2067 8304 2249 9373
rect 2067 8270 2287 8304
rect 2067 8242 2249 8270
rect -2789 -193 6262 6567
<< nmos >>
rect -2580 6157 -2550 6357
rect -2370 6157 -2340 6357
rect -2160 6157 -2130 6357
rect -1950 6157 -1920 6357
rect -1740 6157 -1710 6357
rect -1530 6157 -1500 6357
rect -1320 6157 -1290 6357
rect -1110 6157 -1080 6357
rect -900 6157 -870 6357
rect -690 6157 -660 6357
rect -480 6157 -450 6357
rect -270 6157 -240 6357
rect -60 6157 -30 6357
rect 150 6157 180 6357
rect 360 6157 390 6357
rect 570 6157 600 6357
rect 780 6157 810 6357
rect 990 6157 1020 6357
rect 1200 6157 1230 6357
rect 1410 6157 1440 6357
rect 1620 6157 1650 6357
rect 1830 6157 1860 6357
rect 2040 6157 2070 6357
rect 2250 6157 2280 6357
rect 2460 6157 2490 6357
rect 2670 6157 2700 6357
rect 2880 6157 2910 6357
rect 3090 6157 3120 6357
rect 3300 6157 3330 6357
rect 3510 6157 3540 6357
rect 3720 6157 3750 6357
rect 3930 6157 3960 6357
rect 4140 6157 4170 6357
rect 4350 6157 4380 6357
rect 4560 6157 4590 6357
rect 4770 6157 4800 6357
rect 4980 6157 5010 6357
rect 5190 6157 5220 6357
rect 5400 6157 5430 6357
rect 5610 6157 5640 6357
rect 5820 6157 5850 6357
rect 6030 6157 6060 6357
rect -2580 5717 -2550 5917
rect -2370 5717 -2340 5917
rect -2160 5717 -2130 5917
rect -1950 5717 -1920 5917
rect -1740 5717 -1710 5917
rect -1530 5717 -1500 5917
rect -1320 5717 -1290 5917
rect -1110 5717 -1080 5917
rect -900 5717 -870 5917
rect -690 5717 -660 5917
rect -480 5717 -450 5917
rect -270 5717 -240 5917
rect -60 5717 -30 5917
rect 150 5717 180 5917
rect 360 5717 390 5917
rect 570 5717 600 5917
rect 780 5717 810 5917
rect 990 5717 1020 5917
rect 1200 5717 1230 5917
rect 1410 5717 1440 5917
rect 1620 5717 1650 5917
rect 1830 5717 1860 5917
rect 2040 5717 2070 5917
rect 2250 5717 2280 5917
rect 2460 5717 2490 5917
rect 2670 5717 2700 5917
rect 2880 5717 2910 5917
rect 3090 5717 3120 5917
rect 3300 5717 3330 5917
rect 3510 5717 3540 5917
rect 3720 5717 3750 5917
rect 3930 5717 3960 5917
rect 4140 5717 4170 5917
rect 4350 5717 4380 5917
rect 4560 5717 4590 5917
rect 4770 5717 4800 5917
rect 4980 5717 5010 5917
rect 5190 5717 5220 5917
rect 5400 5717 5430 5917
rect 5610 5717 5640 5917
rect 5820 5717 5850 5917
rect 6030 5717 6060 5917
rect -2580 5277 -2550 5477
rect -2370 5277 -2340 5477
rect -2160 5277 -2130 5477
rect -1950 5277 -1920 5477
rect -1740 5277 -1710 5477
rect -1530 5277 -1500 5477
rect -1320 5277 -1290 5477
rect -1110 5277 -1080 5477
rect -900 5277 -870 5477
rect -690 5277 -660 5477
rect -480 5277 -450 5477
rect -270 5277 -240 5477
rect -60 5277 -30 5477
rect 150 5277 180 5477
rect 360 5277 390 5477
rect 570 5277 600 5477
rect 780 5277 810 5477
rect 990 5277 1020 5477
rect 1200 5277 1230 5477
rect 1410 5277 1440 5477
rect 1620 5277 1650 5477
rect 1830 5277 1860 5477
rect 2040 5277 2070 5477
rect 2250 5277 2280 5477
rect 2460 5277 2490 5477
rect 2670 5277 2700 5477
rect 2880 5277 2910 5477
rect 3090 5277 3120 5477
rect 3300 5277 3330 5477
rect 3510 5277 3540 5477
rect 3720 5277 3750 5477
rect 3930 5277 3960 5477
rect 4140 5277 4170 5477
rect 4350 5277 4380 5477
rect 4560 5277 4590 5477
rect 4770 5277 4800 5477
rect 4980 5277 5010 5477
rect 5190 5277 5220 5477
rect 5400 5277 5430 5477
rect 5610 5277 5640 5477
rect 5820 5277 5850 5477
rect 6030 5277 6060 5477
rect -2580 4837 -2550 5037
rect -2370 4837 -2340 5037
rect -2160 4837 -2130 5037
rect -1950 4837 -1920 5037
rect -1740 4837 -1710 5037
rect -1530 4837 -1500 5037
rect -1320 4837 -1290 5037
rect -1110 4837 -1080 5037
rect -900 4837 -870 5037
rect -690 4837 -660 5037
rect -480 4837 -450 5037
rect -270 4837 -240 5037
rect -60 4837 -30 5037
rect 150 4837 180 5037
rect 360 4837 390 5037
rect 570 4837 600 5037
rect 780 4837 810 5037
rect 990 4837 1020 5037
rect 1200 4837 1230 5037
rect 1410 4837 1440 5037
rect 1620 4837 1650 5037
rect 1830 4837 1860 5037
rect 2040 4837 2070 5037
rect 2250 4837 2280 5037
rect 2460 4837 2490 5037
rect 2670 4837 2700 5037
rect 2880 4837 2910 5037
rect 3090 4837 3120 5037
rect 3300 4837 3330 5037
rect 3510 4837 3540 5037
rect 3720 4837 3750 5037
rect 3930 4837 3960 5037
rect 4140 4837 4170 5037
rect 4350 4837 4380 5037
rect 4560 4837 4590 5037
rect 4770 4837 4800 5037
rect 4980 4837 5010 5037
rect 5190 4837 5220 5037
rect 5400 4837 5430 5037
rect 5610 4837 5640 5037
rect 5820 4837 5850 5037
rect 6030 4837 6060 5037
rect -2580 3902 -2550 4102
rect -2370 3902 -2340 4102
rect -2160 3902 -2130 4102
rect -1950 3902 -1920 4102
rect -1740 3902 -1710 4102
rect -1530 3902 -1500 4102
rect -1320 3902 -1290 4102
rect -1110 3902 -1080 4102
rect -900 3902 -870 4102
rect -690 3902 -660 4102
rect -480 3902 -450 4102
rect -270 3902 -240 4102
rect -60 3902 -30 4102
rect 150 3902 180 4102
rect 360 3902 390 4102
rect 570 3902 600 4102
rect 780 3902 810 4102
rect 990 3902 1020 4102
rect 1200 3902 1230 4102
rect 1410 3902 1440 4102
rect 1620 3902 1650 4102
rect 1830 3902 1860 4102
rect 2040 3902 2070 4102
rect 2250 3902 2280 4102
rect 2460 3902 2490 4102
rect 2670 3902 2700 4102
rect 2880 3902 2910 4102
rect 3090 3902 3120 4102
rect 3300 3902 3330 4102
rect 3510 3902 3540 4102
rect 3720 3902 3750 4102
rect 3930 3902 3960 4102
rect 4140 3902 4170 4102
rect 4350 3902 4380 4102
rect 4560 3902 4590 4102
rect 4770 3902 4800 4102
rect 4980 3902 5010 4102
rect 5190 3902 5220 4102
rect 5400 3902 5430 4102
rect 5610 3902 5640 4102
rect 5820 3902 5850 4102
rect 6030 3902 6060 4102
rect -2580 3462 -2550 3662
rect -2370 3462 -2340 3662
rect -2160 3462 -2130 3662
rect -1950 3462 -1920 3662
rect -1740 3462 -1710 3662
rect -1530 3462 -1500 3662
rect -1320 3462 -1290 3662
rect -1110 3462 -1080 3662
rect -900 3462 -870 3662
rect -690 3462 -660 3662
rect -480 3462 -450 3662
rect -270 3462 -240 3662
rect -60 3462 -30 3662
rect 150 3462 180 3662
rect 360 3462 390 3662
rect 570 3462 600 3662
rect 780 3462 810 3662
rect 990 3462 1020 3662
rect 1200 3462 1230 3662
rect 1410 3462 1440 3662
rect 1620 3462 1650 3662
rect 1830 3462 1860 3662
rect 2040 3462 2070 3662
rect 2250 3462 2280 3662
rect 2460 3462 2490 3662
rect 2670 3462 2700 3662
rect 2880 3462 2910 3662
rect 3090 3462 3120 3662
rect 3300 3462 3330 3662
rect 3510 3462 3540 3662
rect 3720 3462 3750 3662
rect 3930 3462 3960 3662
rect 4140 3462 4170 3662
rect 4350 3462 4380 3662
rect 4560 3462 4590 3662
rect 4770 3462 4800 3662
rect 4980 3462 5010 3662
rect 5190 3462 5220 3662
rect 5400 3462 5430 3662
rect 5610 3462 5640 3662
rect 5820 3462 5850 3662
rect 6030 3462 6060 3662
rect -2580 3022 -2550 3222
rect -2370 3022 -2340 3222
rect -2160 3022 -2130 3222
rect -1950 3022 -1920 3222
rect -1740 3022 -1710 3222
rect -1530 3022 -1500 3222
rect -1320 3022 -1290 3222
rect -1110 3022 -1080 3222
rect -900 3022 -870 3222
rect -690 3022 -660 3222
rect -480 3022 -450 3222
rect -270 3022 -240 3222
rect -60 3022 -30 3222
rect 150 3022 180 3222
rect 360 3022 390 3222
rect 570 3022 600 3222
rect 780 3022 810 3222
rect 990 3022 1020 3222
rect 1200 3022 1230 3222
rect 1410 3022 1440 3222
rect 1620 3022 1650 3222
rect 1830 3022 1860 3222
rect 2040 3022 2070 3222
rect 2250 3022 2280 3222
rect 2460 3022 2490 3222
rect 2670 3022 2700 3222
rect 2880 3022 2910 3222
rect 3090 3022 3120 3222
rect 3300 3022 3330 3222
rect 3510 3022 3540 3222
rect 3720 3022 3750 3222
rect 3930 3022 3960 3222
rect 4140 3022 4170 3222
rect 4350 3022 4380 3222
rect 4560 3022 4590 3222
rect 4770 3022 4800 3222
rect 4980 3022 5010 3222
rect 5190 3022 5220 3222
rect 5400 3022 5430 3222
rect 5610 3022 5640 3222
rect 5820 3022 5850 3222
rect 6030 3022 6060 3222
rect -2580 2582 -2550 2782
rect -2370 2582 -2340 2782
rect -2160 2582 -2130 2782
rect -1950 2582 -1920 2782
rect -1740 2582 -1710 2782
rect -1530 2582 -1500 2782
rect -1320 2582 -1290 2782
rect -1110 2582 -1080 2782
rect -900 2582 -870 2782
rect -690 2582 -660 2782
rect -480 2582 -450 2782
rect -270 2582 -240 2782
rect -60 2582 -30 2782
rect 150 2582 180 2782
rect 360 2582 390 2782
rect 570 2582 600 2782
rect 780 2582 810 2782
rect 990 2582 1020 2782
rect 1200 2582 1230 2782
rect 1410 2582 1440 2782
rect 1620 2582 1650 2782
rect 1830 2582 1860 2782
rect 2040 2582 2070 2782
rect 2250 2582 2280 2782
rect 2460 2582 2490 2782
rect 2670 2582 2700 2782
rect 2880 2582 2910 2782
rect 3090 2582 3120 2782
rect 3300 2582 3330 2782
rect 3510 2582 3540 2782
rect 3720 2582 3750 2782
rect 3930 2582 3960 2782
rect 4140 2582 4170 2782
rect 4350 2582 4380 2782
rect 4560 2582 4590 2782
rect 4770 2582 4800 2782
rect 4980 2582 5010 2782
rect 5190 2582 5220 2782
rect 5400 2582 5430 2782
rect 5610 2582 5640 2782
rect 5820 2582 5850 2782
rect 6030 2582 6060 2782
rect -2580 2142 -2550 2342
rect -2370 2142 -2340 2342
rect -2160 2142 -2130 2342
rect -1950 2142 -1920 2342
rect -1740 2142 -1710 2342
rect -1530 2142 -1500 2342
rect -1320 2142 -1290 2342
rect -1110 2142 -1080 2342
rect -900 2142 -870 2342
rect -690 2142 -660 2342
rect -480 2142 -450 2342
rect -270 2142 -240 2342
rect -60 2142 -30 2342
rect 150 2142 180 2342
rect 360 2142 390 2342
rect 570 2142 600 2342
rect 780 2142 810 2342
rect 990 2142 1020 2342
rect 1200 2142 1230 2342
rect 1410 2142 1440 2342
rect 1620 2142 1650 2342
rect 1830 2142 1860 2342
rect 2040 2142 2070 2342
rect 2250 2142 2280 2342
rect 2460 2142 2490 2342
rect 2670 2142 2700 2342
rect 2880 2142 2910 2342
rect 3090 2142 3120 2342
rect 3300 2142 3330 2342
rect 3510 2142 3540 2342
rect 3720 2142 3750 2342
rect 3930 2142 3960 2342
rect 4140 2142 4170 2342
rect 4350 2142 4380 2342
rect 4560 2142 4590 2342
rect 4770 2142 4800 2342
rect 4980 2142 5010 2342
rect 5190 2142 5220 2342
rect 5400 2142 5430 2342
rect 5610 2142 5640 2342
rect 5820 2142 5850 2342
rect 6030 2142 6060 2342
rect -2580 1702 -2550 1902
rect -2370 1702 -2340 1902
rect -2160 1702 -2130 1902
rect -1950 1702 -1920 1902
rect -1740 1702 -1710 1902
rect -1530 1702 -1500 1902
rect -1320 1702 -1290 1902
rect -1110 1702 -1080 1902
rect -900 1702 -870 1902
rect -690 1702 -660 1902
rect -480 1702 -450 1902
rect -270 1702 -240 1902
rect -60 1702 -30 1902
rect 150 1702 180 1902
rect 360 1702 390 1902
rect 570 1702 600 1902
rect 780 1702 810 1902
rect 990 1702 1020 1902
rect 1200 1702 1230 1902
rect 1410 1702 1440 1902
rect 1620 1702 1650 1902
rect 1830 1702 1860 1902
rect 2040 1702 2070 1902
rect 2250 1702 2280 1902
rect 2460 1702 2490 1902
rect 2670 1702 2700 1902
rect 2880 1702 2910 1902
rect 3090 1702 3120 1902
rect 3300 1702 3330 1902
rect 3510 1702 3540 1902
rect 3720 1702 3750 1902
rect 3930 1702 3960 1902
rect 4140 1702 4170 1902
rect 4350 1702 4380 1902
rect 4560 1702 4590 1902
rect 4770 1702 4800 1902
rect 4980 1702 5010 1902
rect 5190 1702 5220 1902
rect 5400 1702 5430 1902
rect 5610 1702 5640 1902
rect 5820 1702 5850 1902
rect 6030 1702 6060 1902
rect -2580 1262 -2550 1462
rect -2370 1262 -2340 1462
rect -2160 1262 -2130 1462
rect -1950 1262 -1920 1462
rect -1740 1262 -1710 1462
rect -1530 1262 -1500 1462
rect -1320 1262 -1290 1462
rect -1110 1262 -1080 1462
rect -900 1262 -870 1462
rect -690 1262 -660 1462
rect -480 1262 -450 1462
rect -270 1262 -240 1462
rect -60 1262 -30 1462
rect 150 1262 180 1462
rect 360 1262 390 1462
rect 570 1262 600 1462
rect 780 1262 810 1462
rect 990 1262 1020 1462
rect 1200 1262 1230 1462
rect 1410 1262 1440 1462
rect 1620 1262 1650 1462
rect 1830 1262 1860 1462
rect 2040 1262 2070 1462
rect 2250 1262 2280 1462
rect 2460 1262 2490 1462
rect 2670 1262 2700 1462
rect 2880 1262 2910 1462
rect 3090 1262 3120 1462
rect 3300 1262 3330 1462
rect 3510 1262 3540 1462
rect 3720 1262 3750 1462
rect 3930 1262 3960 1462
rect 4140 1262 4170 1462
rect 4350 1262 4380 1462
rect 4560 1262 4590 1462
rect 4770 1262 4800 1462
rect 4980 1262 5010 1462
rect 5190 1262 5220 1462
rect 5400 1262 5430 1462
rect 5610 1262 5640 1462
rect 5820 1262 5850 1462
rect 6030 1262 6060 1462
rect -2580 822 -2550 1022
rect -2370 822 -2340 1022
rect -2160 822 -2130 1022
rect -1950 822 -1920 1022
rect -1740 822 -1710 1022
rect -1530 822 -1500 1022
rect -1320 822 -1290 1022
rect -1110 822 -1080 1022
rect -900 822 -870 1022
rect -690 822 -660 1022
rect -480 822 -450 1022
rect -270 822 -240 1022
rect -60 822 -30 1022
rect 150 822 180 1022
rect 360 822 390 1022
rect 570 822 600 1022
rect 780 822 810 1022
rect 990 822 1020 1022
rect 1200 822 1230 1022
rect 1410 822 1440 1022
rect 1620 822 1650 1022
rect 1830 822 1860 1022
rect 2040 822 2070 1022
rect 2250 822 2280 1022
rect 2460 822 2490 1022
rect 2670 822 2700 1022
rect 2880 822 2910 1022
rect 3090 822 3120 1022
rect 3300 822 3330 1022
rect 3510 822 3540 1022
rect 3720 822 3750 1022
rect 3930 822 3960 1022
rect 4140 822 4170 1022
rect 4350 822 4380 1022
rect 4560 822 4590 1022
rect 4770 822 4800 1022
rect 4980 822 5010 1022
rect 5190 822 5220 1022
rect 5400 822 5430 1022
rect 5610 822 5640 1022
rect 5820 822 5850 1022
rect 6030 822 6060 1022
rect 140 18 170 218
rect 236 18 266 218
rect 332 18 362 218
rect 428 18 458 218
rect 524 18 554 218
rect 620 18 650 218
rect 716 18 746 218
rect 812 18 842 218
rect 908 18 938 218
rect 1004 18 1034 218
rect 1100 18 1130 218
rect 1196 18 1226 218
rect 1292 18 1322 218
rect 1388 18 1418 218
rect 1484 18 1514 218
rect 1580 18 1610 218
rect 1676 18 1706 218
rect 1772 18 1802 218
rect 1868 18 1898 218
rect 1964 18 1994 218
rect 2060 18 2090 218
rect 2156 18 2186 218
rect 2252 18 2282 218
rect 2348 18 2378 218
rect 2444 18 2474 218
rect 2540 18 2570 218
rect 2636 18 2666 218
rect 2732 18 2762 218
rect 2828 18 2858 218
rect 2924 18 2954 218
rect 3020 18 3050 218
rect 3116 18 3146 218
rect 3212 18 3242 218
rect 3308 18 3338 218
<< scnmos >>
rect 1229 9608 1339 10554
rect 2113 9608 2223 10554
rect 1229 9328 1359 9358
rect 2093 9328 2223 9358
rect 1229 9244 1359 9274
rect 2093 9244 2223 9274
rect 1229 9160 1359 9190
rect 2093 9160 2223 9190
rect 1229 9076 1359 9106
rect 2093 9076 2223 9106
rect 1229 8992 1359 9022
rect 2093 8992 2223 9022
rect 1229 8908 1359 8938
rect 2093 8908 2223 8938
rect 1229 8824 1359 8854
rect 2093 8824 2223 8854
rect 1229 8740 1359 8770
rect 2093 8740 2223 8770
rect 1229 8499 1359 8529
rect 2093 8499 2223 8529
rect 1229 8415 1359 8445
rect 2093 8415 2223 8445
rect 1229 8320 1313 8350
rect 2139 8320 2223 8350
<< pmos >>
rect -3569 7830 -3369 7860
rect -3569 7734 -3369 7764
rect -3569 7638 -3369 7668
rect -3569 7542 -3369 7572
rect -3569 7446 -3369 7476
rect -3569 7350 -3369 7380
rect -3569 7254 -3369 7284
rect -3569 7158 -3369 7188
rect -3569 7062 -3369 7092
rect -3569 6966 -3369 6996
rect -3569 6870 -3369 6900
rect -3569 6774 -3369 6804
rect -3569 6678 -3369 6708
rect -3569 6582 -3369 6612
rect -3569 6486 -3369 6516
rect -3569 6390 -3369 6420
rect -3569 6294 -3369 6324
rect -3569 6198 -3369 6228
rect -2594 7640 -2564 7840
rect -2384 7640 -2354 7840
rect -2174 7640 -2144 7840
rect -1964 7640 -1934 7840
rect -1754 7640 -1724 7840
rect -1544 7640 -1514 7840
rect -1334 7640 -1304 7840
rect -1124 7640 -1094 7840
rect -914 7640 -884 7840
rect -704 7640 -674 7840
rect -494 7640 -464 7840
rect -284 7640 -254 7840
rect -74 7640 -44 7840
rect 136 7640 166 7840
rect 346 7640 376 7840
rect 556 7640 586 7840
rect 766 7640 796 7840
rect 976 7640 1006 7840
rect 1186 7640 1216 7840
rect 1396 7640 1426 7840
rect 1606 7640 1636 7840
rect 1816 7640 1846 7840
rect 2026 7640 2056 7840
rect 2236 7640 2266 7840
rect 2446 7640 2476 7840
rect 2656 7640 2686 7840
rect 2866 7640 2896 7840
rect 3076 7640 3106 7840
rect 3286 7640 3316 7840
rect 3496 7640 3526 7840
rect 3706 7640 3736 7840
rect 3916 7640 3946 7840
rect 4126 7640 4156 7840
rect 4336 7640 4366 7840
rect 4546 7640 4576 7840
rect 4756 7640 4786 7840
rect 4966 7640 4996 7840
rect 5176 7640 5206 7840
rect 5386 7640 5416 7840
rect 5596 7640 5626 7840
rect 5806 7640 5836 7840
rect 6016 7640 6046 7840
rect -2592 7107 -2562 7307
rect -2382 7107 -2352 7307
rect -2172 7107 -2142 7307
rect -1962 7107 -1932 7307
rect -1752 7107 -1722 7307
rect -1542 7107 -1512 7307
rect -1332 7107 -1302 7307
rect -1122 7107 -1092 7307
rect -912 7107 -882 7307
rect -702 7107 -672 7307
rect -492 7107 -462 7307
rect -282 7107 -252 7307
rect -72 7107 -42 7307
rect 138 7107 168 7307
rect 348 7107 378 7307
rect 558 7107 588 7307
rect 768 7107 798 7307
rect 978 7107 1008 7307
rect 1188 7107 1218 7307
rect 1398 7107 1428 7307
rect 1608 7107 1638 7307
rect 1818 7107 1848 7307
rect 2028 7107 2058 7307
rect 2238 7107 2268 7307
rect 2448 7107 2478 7307
rect 2658 7107 2688 7307
rect 2868 7107 2898 7307
rect 3078 7107 3108 7307
rect 3288 7107 3318 7307
rect 3498 7107 3528 7307
rect 3708 7107 3738 7307
rect 3918 7107 3948 7307
rect 4128 7107 4158 7307
rect 4338 7107 4368 7307
rect 4548 7107 4578 7307
rect 4758 7107 4788 7307
rect 4968 7107 4998 7307
rect 5178 7107 5208 7307
rect 5388 7107 5418 7307
rect 5598 7107 5628 7307
rect 5808 7107 5838 7307
rect 6018 7107 6048 7307
rect -3567 5420 -3367 5450
rect -3567 5324 -3367 5354
rect -3567 5228 -3367 5258
rect -3567 5132 -3367 5162
rect -3567 5036 -3367 5066
rect -3567 4940 -3367 4970
rect -3567 4844 -3367 4874
rect -3567 4748 -3367 4778
rect -3567 4652 -3367 4682
rect -3567 4556 -3367 4586
rect -3567 4460 -3367 4490
rect -3567 4364 -3367 4394
rect -3567 4268 -3367 4298
rect -3567 4172 -3367 4202
rect -3567 4076 -3367 4106
rect -3567 3980 -3367 4010
rect -3567 3884 -3367 3914
rect -3567 3788 -3367 3818
rect 6831 7830 7031 7860
rect 6831 7734 7031 7764
rect 6831 7638 7031 7668
rect 6831 7542 7031 7572
rect 6831 7446 7031 7476
rect 6831 7350 7031 7380
rect 6831 7254 7031 7284
rect 6831 7158 7031 7188
rect 6831 7062 7031 7092
rect 6831 6966 7031 6996
rect 6831 6870 7031 6900
rect 6831 6774 7031 6804
rect 6831 6678 7031 6708
rect 6831 6582 7031 6612
rect 6831 6486 7031 6516
rect 6831 6390 7031 6420
rect 6831 6294 7031 6324
rect 6831 6198 7031 6228
rect 6831 5420 7031 5450
rect 6831 5324 7031 5354
rect 6831 5228 7031 5258
rect 6831 5132 7031 5162
rect 6831 5036 7031 5066
rect 6831 4940 7031 4970
rect 6831 4844 7031 4874
rect 6831 4748 7031 4778
rect 6831 4652 7031 4682
rect 6831 4556 7031 4586
rect 6831 4460 7031 4490
rect 6831 4364 7031 4394
rect 6831 4268 7031 4298
rect 6831 4172 7031 4202
rect 6831 4076 7031 4106
rect 6831 3980 7031 4010
rect 6831 3884 7031 3914
rect 6831 3788 7031 3818
<< scpmoshvt >>
rect 1505 9608 1679 10554
rect 1773 9608 1947 10554
rect 1479 9328 1679 9358
rect 1773 9328 1973 9358
rect 1479 9244 1679 9274
rect 1773 9244 1973 9274
rect 1479 9160 1679 9190
rect 1773 9160 1973 9190
rect 1479 9076 1679 9106
rect 1773 9076 1973 9106
rect 1479 8992 1679 9022
rect 1773 8992 1973 9022
rect 1479 8908 1679 8938
rect 1773 8908 1973 8938
rect 1479 8824 1679 8854
rect 1773 8824 1973 8854
rect 1479 8740 1679 8770
rect 1773 8740 1973 8770
rect 1479 8499 1679 8529
rect 1773 8499 1973 8529
rect 1479 8415 1679 8445
rect 1773 8415 1973 8445
rect 1543 8320 1671 8350
rect 1781 8320 1909 8350
<< ndiff >>
rect 1229 10598 1339 10606
rect 1229 10564 1260 10598
rect 1294 10564 1339 10598
rect 1229 10554 1339 10564
rect 2113 10598 2223 10606
rect 2113 10564 2158 10598
rect 2192 10564 2223 10598
rect 2113 10554 2223 10564
rect 1229 9598 1339 9608
rect 1229 9564 1260 9598
rect 1294 9564 1339 9598
rect 1229 9556 1339 9564
rect 2113 9598 2223 9608
rect 2113 9564 2158 9598
rect 2192 9564 2223 9598
rect 2113 9556 2223 9564
rect 1229 9402 1359 9410
rect 1229 9368 1241 9402
rect 1275 9368 1309 9402
rect 1343 9368 1359 9402
rect 1229 9358 1359 9368
rect 2093 9402 2223 9410
rect 2093 9368 2109 9402
rect 2143 9368 2177 9402
rect 2211 9368 2223 9402
rect 2093 9358 2223 9368
rect 1229 9318 1359 9328
rect 1229 9284 1241 9318
rect 1275 9284 1359 9318
rect 1229 9274 1359 9284
rect 2093 9318 2223 9328
rect 2093 9284 2177 9318
rect 2211 9284 2223 9318
rect 2093 9274 2223 9284
rect 1229 9234 1359 9244
rect 1229 9200 1241 9234
rect 1275 9200 1309 9234
rect 1343 9200 1359 9234
rect 1229 9190 1359 9200
rect 2093 9234 2223 9244
rect 2093 9200 2109 9234
rect 2143 9200 2177 9234
rect 2211 9200 2223 9234
rect 2093 9190 2223 9200
rect 1229 9150 1359 9160
rect 1229 9116 1241 9150
rect 1275 9116 1359 9150
rect 1229 9106 1359 9116
rect 2093 9150 2223 9160
rect 2093 9116 2177 9150
rect 2211 9116 2223 9150
rect 2093 9106 2223 9116
rect 1229 9066 1359 9076
rect 1229 9032 1241 9066
rect 1275 9032 1309 9066
rect 1343 9032 1359 9066
rect 1229 9022 1359 9032
rect 2093 9066 2223 9076
rect 2093 9032 2109 9066
rect 2143 9032 2177 9066
rect 2211 9032 2223 9066
rect 2093 9022 2223 9032
rect 1229 8982 1359 8992
rect 1229 8948 1309 8982
rect 1343 8948 1359 8982
rect 1229 8938 1359 8948
rect 2093 8982 2223 8992
rect 2093 8948 2109 8982
rect 2143 8948 2223 8982
rect 2093 8938 2223 8948
rect 1229 8898 1359 8908
rect 1229 8864 1241 8898
rect 1275 8864 1359 8898
rect 1229 8854 1359 8864
rect 2093 8898 2223 8908
rect 2093 8864 2177 8898
rect 2211 8864 2223 8898
rect 2093 8854 2223 8864
rect 1229 8814 1359 8824
rect 1229 8780 1309 8814
rect 1343 8780 1359 8814
rect 1229 8770 1359 8780
rect 2093 8814 2223 8824
rect 2093 8780 2109 8814
rect 2143 8780 2223 8814
rect 2093 8770 2223 8780
rect 1229 8730 1359 8740
rect 1229 8696 1241 8730
rect 1275 8696 1309 8730
rect 1343 8696 1359 8730
rect 1229 8688 1359 8696
rect 2093 8730 2223 8740
rect 2093 8696 2109 8730
rect 2143 8696 2177 8730
rect 2211 8696 2223 8730
rect 2093 8688 2223 8696
rect 1229 8573 1359 8582
rect 1229 8539 1245 8573
rect 1279 8539 1313 8573
rect 1347 8539 1359 8573
rect 1229 8529 1359 8539
rect 2093 8573 2223 8582
rect 2093 8539 2105 8573
rect 2139 8539 2173 8573
rect 2207 8539 2223 8573
rect 2093 8529 2223 8539
rect 1229 8489 1359 8499
rect 1229 8455 1271 8489
rect 1305 8455 1359 8489
rect 1229 8445 1359 8455
rect 2093 8489 2223 8499
rect 2093 8455 2147 8489
rect 2181 8455 2223 8489
rect 2093 8445 2223 8455
rect 1229 8403 1359 8415
rect 1229 8369 1241 8403
rect 1275 8369 1359 8403
rect 1229 8365 1359 8369
rect 2093 8403 2223 8415
rect 2093 8369 2177 8403
rect 2211 8369 2223 8403
rect 2093 8365 2223 8369
rect 1229 8350 1313 8365
rect 2139 8350 2223 8365
rect 1229 8310 1313 8320
rect 1229 8276 1254 8310
rect 1288 8276 1313 8310
rect 1229 8268 1313 8276
rect 2139 8310 2223 8320
rect 2139 8276 2164 8310
rect 2198 8276 2223 8310
rect 2139 8268 2223 8276
rect -2642 6345 -2580 6357
rect -2642 6169 -2630 6345
rect -2596 6169 -2580 6345
rect -2642 6157 -2580 6169
rect -2550 6345 -2488 6357
rect -2550 6169 -2534 6345
rect -2500 6169 -2488 6345
rect -2550 6157 -2488 6169
rect -2432 6345 -2370 6357
rect -2432 6169 -2420 6345
rect -2386 6169 -2370 6345
rect -2432 6157 -2370 6169
rect -2340 6345 -2278 6357
rect -2340 6169 -2324 6345
rect -2290 6169 -2278 6345
rect -2340 6157 -2278 6169
rect -2222 6345 -2160 6357
rect -2222 6169 -2210 6345
rect -2176 6169 -2160 6345
rect -2222 6157 -2160 6169
rect -2130 6345 -2068 6357
rect -2130 6169 -2114 6345
rect -2080 6169 -2068 6345
rect -2130 6157 -2068 6169
rect -2012 6345 -1950 6357
rect -2012 6169 -2000 6345
rect -1966 6169 -1950 6345
rect -2012 6157 -1950 6169
rect -1920 6345 -1858 6357
rect -1920 6169 -1904 6345
rect -1870 6169 -1858 6345
rect -1920 6157 -1858 6169
rect -1802 6345 -1740 6357
rect -1802 6169 -1790 6345
rect -1756 6169 -1740 6345
rect -1802 6157 -1740 6169
rect -1710 6345 -1648 6357
rect -1710 6169 -1694 6345
rect -1660 6169 -1648 6345
rect -1710 6157 -1648 6169
rect -1592 6345 -1530 6357
rect -1592 6169 -1580 6345
rect -1546 6169 -1530 6345
rect -1592 6157 -1530 6169
rect -1500 6345 -1438 6357
rect -1500 6169 -1484 6345
rect -1450 6169 -1438 6345
rect -1500 6157 -1438 6169
rect -1382 6345 -1320 6357
rect -1382 6169 -1370 6345
rect -1336 6169 -1320 6345
rect -1382 6157 -1320 6169
rect -1290 6345 -1228 6357
rect -1290 6169 -1274 6345
rect -1240 6169 -1228 6345
rect -1290 6157 -1228 6169
rect -1172 6345 -1110 6357
rect -1172 6169 -1160 6345
rect -1126 6169 -1110 6345
rect -1172 6157 -1110 6169
rect -1080 6345 -1018 6357
rect -1080 6169 -1064 6345
rect -1030 6169 -1018 6345
rect -1080 6157 -1018 6169
rect -962 6345 -900 6357
rect -962 6169 -950 6345
rect -916 6169 -900 6345
rect -962 6157 -900 6169
rect -870 6345 -808 6357
rect -870 6169 -854 6345
rect -820 6169 -808 6345
rect -870 6157 -808 6169
rect -752 6345 -690 6357
rect -752 6169 -740 6345
rect -706 6169 -690 6345
rect -752 6157 -690 6169
rect -660 6345 -598 6357
rect -660 6169 -644 6345
rect -610 6169 -598 6345
rect -660 6157 -598 6169
rect -542 6345 -480 6357
rect -542 6169 -530 6345
rect -496 6169 -480 6345
rect -542 6157 -480 6169
rect -450 6345 -388 6357
rect -450 6169 -434 6345
rect -400 6169 -388 6345
rect -450 6157 -388 6169
rect -332 6345 -270 6357
rect -332 6169 -320 6345
rect -286 6169 -270 6345
rect -332 6157 -270 6169
rect -240 6345 -178 6357
rect -240 6169 -224 6345
rect -190 6169 -178 6345
rect -240 6157 -178 6169
rect -122 6345 -60 6357
rect -122 6169 -110 6345
rect -76 6169 -60 6345
rect -122 6157 -60 6169
rect -30 6345 32 6357
rect -30 6169 -14 6345
rect 20 6169 32 6345
rect -30 6157 32 6169
rect 88 6345 150 6357
rect 88 6169 100 6345
rect 134 6169 150 6345
rect 88 6157 150 6169
rect 180 6345 242 6357
rect 180 6169 196 6345
rect 230 6169 242 6345
rect 180 6157 242 6169
rect 298 6345 360 6357
rect 298 6169 310 6345
rect 344 6169 360 6345
rect 298 6157 360 6169
rect 390 6345 452 6357
rect 390 6169 406 6345
rect 440 6169 452 6345
rect 390 6157 452 6169
rect 508 6345 570 6357
rect 508 6169 520 6345
rect 554 6169 570 6345
rect 508 6157 570 6169
rect 600 6345 662 6357
rect 600 6169 616 6345
rect 650 6169 662 6345
rect 600 6157 662 6169
rect 718 6345 780 6357
rect 718 6169 730 6345
rect 764 6169 780 6345
rect 718 6157 780 6169
rect 810 6345 872 6357
rect 810 6169 826 6345
rect 860 6169 872 6345
rect 810 6157 872 6169
rect 928 6345 990 6357
rect 928 6169 940 6345
rect 974 6169 990 6345
rect 928 6157 990 6169
rect 1020 6345 1082 6357
rect 1020 6169 1036 6345
rect 1070 6169 1082 6345
rect 1020 6157 1082 6169
rect 1138 6345 1200 6357
rect 1138 6169 1150 6345
rect 1184 6169 1200 6345
rect 1138 6157 1200 6169
rect 1230 6345 1292 6357
rect 1230 6169 1246 6345
rect 1280 6169 1292 6345
rect 1230 6157 1292 6169
rect 1348 6345 1410 6357
rect 1348 6169 1360 6345
rect 1394 6169 1410 6345
rect 1348 6157 1410 6169
rect 1440 6345 1502 6357
rect 1440 6169 1456 6345
rect 1490 6169 1502 6345
rect 1440 6157 1502 6169
rect 1558 6345 1620 6357
rect 1558 6169 1570 6345
rect 1604 6169 1620 6345
rect 1558 6157 1620 6169
rect 1650 6345 1712 6357
rect 1650 6169 1666 6345
rect 1700 6169 1712 6345
rect 1650 6157 1712 6169
rect 1768 6345 1830 6357
rect 1768 6169 1780 6345
rect 1814 6169 1830 6345
rect 1768 6157 1830 6169
rect 1860 6345 1922 6357
rect 1860 6169 1876 6345
rect 1910 6169 1922 6345
rect 1860 6157 1922 6169
rect 1978 6345 2040 6357
rect 1978 6169 1990 6345
rect 2024 6169 2040 6345
rect 1978 6157 2040 6169
rect 2070 6345 2132 6357
rect 2070 6169 2086 6345
rect 2120 6169 2132 6345
rect 2070 6157 2132 6169
rect 2188 6345 2250 6357
rect 2188 6169 2200 6345
rect 2234 6169 2250 6345
rect 2188 6157 2250 6169
rect 2280 6345 2342 6357
rect 2280 6169 2296 6345
rect 2330 6169 2342 6345
rect 2280 6157 2342 6169
rect 2398 6345 2460 6357
rect 2398 6169 2410 6345
rect 2444 6169 2460 6345
rect 2398 6157 2460 6169
rect 2490 6345 2552 6357
rect 2490 6169 2506 6345
rect 2540 6169 2552 6345
rect 2490 6157 2552 6169
rect 2608 6345 2670 6357
rect 2608 6169 2620 6345
rect 2654 6169 2670 6345
rect 2608 6157 2670 6169
rect 2700 6345 2762 6357
rect 2700 6169 2716 6345
rect 2750 6169 2762 6345
rect 2700 6157 2762 6169
rect 2818 6345 2880 6357
rect 2818 6169 2830 6345
rect 2864 6169 2880 6345
rect 2818 6157 2880 6169
rect 2910 6345 2972 6357
rect 2910 6169 2926 6345
rect 2960 6169 2972 6345
rect 2910 6157 2972 6169
rect 3028 6345 3090 6357
rect 3028 6169 3040 6345
rect 3074 6169 3090 6345
rect 3028 6157 3090 6169
rect 3120 6345 3182 6357
rect 3120 6169 3136 6345
rect 3170 6169 3182 6345
rect 3120 6157 3182 6169
rect 3238 6345 3300 6357
rect 3238 6169 3250 6345
rect 3284 6169 3300 6345
rect 3238 6157 3300 6169
rect 3330 6345 3392 6357
rect 3330 6169 3346 6345
rect 3380 6169 3392 6345
rect 3330 6157 3392 6169
rect 3448 6345 3510 6357
rect 3448 6169 3460 6345
rect 3494 6169 3510 6345
rect 3448 6157 3510 6169
rect 3540 6345 3602 6357
rect 3540 6169 3556 6345
rect 3590 6169 3602 6345
rect 3540 6157 3602 6169
rect 3658 6345 3720 6357
rect 3658 6169 3670 6345
rect 3704 6169 3720 6345
rect 3658 6157 3720 6169
rect 3750 6345 3812 6357
rect 3750 6169 3766 6345
rect 3800 6169 3812 6345
rect 3750 6157 3812 6169
rect 3868 6345 3930 6357
rect 3868 6169 3880 6345
rect 3914 6169 3930 6345
rect 3868 6157 3930 6169
rect 3960 6345 4022 6357
rect 3960 6169 3976 6345
rect 4010 6169 4022 6345
rect 3960 6157 4022 6169
rect 4078 6345 4140 6357
rect 4078 6169 4090 6345
rect 4124 6169 4140 6345
rect 4078 6157 4140 6169
rect 4170 6345 4232 6357
rect 4170 6169 4186 6345
rect 4220 6169 4232 6345
rect 4170 6157 4232 6169
rect 4288 6345 4350 6357
rect 4288 6169 4300 6345
rect 4334 6169 4350 6345
rect 4288 6157 4350 6169
rect 4380 6345 4442 6357
rect 4380 6169 4396 6345
rect 4430 6169 4442 6345
rect 4380 6157 4442 6169
rect 4498 6345 4560 6357
rect 4498 6169 4510 6345
rect 4544 6169 4560 6345
rect 4498 6157 4560 6169
rect 4590 6345 4652 6357
rect 4590 6169 4606 6345
rect 4640 6169 4652 6345
rect 4590 6157 4652 6169
rect 4708 6345 4770 6357
rect 4708 6169 4720 6345
rect 4754 6169 4770 6345
rect 4708 6157 4770 6169
rect 4800 6345 4862 6357
rect 4800 6169 4816 6345
rect 4850 6169 4862 6345
rect 4800 6157 4862 6169
rect 4918 6345 4980 6357
rect 4918 6169 4930 6345
rect 4964 6169 4980 6345
rect 4918 6157 4980 6169
rect 5010 6345 5072 6357
rect 5010 6169 5026 6345
rect 5060 6169 5072 6345
rect 5010 6157 5072 6169
rect 5128 6345 5190 6357
rect 5128 6169 5140 6345
rect 5174 6169 5190 6345
rect 5128 6157 5190 6169
rect 5220 6345 5282 6357
rect 5220 6169 5236 6345
rect 5270 6169 5282 6345
rect 5220 6157 5282 6169
rect 5338 6345 5400 6357
rect 5338 6169 5350 6345
rect 5384 6169 5400 6345
rect 5338 6157 5400 6169
rect 5430 6345 5492 6357
rect 5430 6169 5446 6345
rect 5480 6169 5492 6345
rect 5430 6157 5492 6169
rect 5548 6345 5610 6357
rect 5548 6169 5560 6345
rect 5594 6169 5610 6345
rect 5548 6157 5610 6169
rect 5640 6345 5702 6357
rect 5640 6169 5656 6345
rect 5690 6169 5702 6345
rect 5640 6157 5702 6169
rect 5758 6345 5820 6357
rect 5758 6169 5770 6345
rect 5804 6169 5820 6345
rect 5758 6157 5820 6169
rect 5850 6345 5912 6357
rect 5850 6169 5866 6345
rect 5900 6169 5912 6345
rect 5850 6157 5912 6169
rect 5968 6345 6030 6357
rect 5968 6169 5980 6345
rect 6014 6169 6030 6345
rect 5968 6157 6030 6169
rect 6060 6345 6122 6357
rect 6060 6169 6076 6345
rect 6110 6169 6122 6345
rect 6060 6157 6122 6169
rect -2642 5905 -2580 5917
rect -2642 5729 -2630 5905
rect -2596 5729 -2580 5905
rect -2642 5717 -2580 5729
rect -2550 5905 -2488 5917
rect -2550 5729 -2534 5905
rect -2500 5729 -2488 5905
rect -2550 5717 -2488 5729
rect -2432 5905 -2370 5917
rect -2432 5729 -2420 5905
rect -2386 5729 -2370 5905
rect -2432 5717 -2370 5729
rect -2340 5905 -2278 5917
rect -2340 5729 -2324 5905
rect -2290 5729 -2278 5905
rect -2340 5717 -2278 5729
rect -2222 5905 -2160 5917
rect -2222 5729 -2210 5905
rect -2176 5729 -2160 5905
rect -2222 5717 -2160 5729
rect -2130 5905 -2068 5917
rect -2130 5729 -2114 5905
rect -2080 5729 -2068 5905
rect -2130 5717 -2068 5729
rect -2012 5905 -1950 5917
rect -2012 5729 -2000 5905
rect -1966 5729 -1950 5905
rect -2012 5717 -1950 5729
rect -1920 5905 -1858 5917
rect -1920 5729 -1904 5905
rect -1870 5729 -1858 5905
rect -1920 5717 -1858 5729
rect -1802 5905 -1740 5917
rect -1802 5729 -1790 5905
rect -1756 5729 -1740 5905
rect -1802 5717 -1740 5729
rect -1710 5905 -1648 5917
rect -1710 5729 -1694 5905
rect -1660 5729 -1648 5905
rect -1710 5717 -1648 5729
rect -1592 5905 -1530 5917
rect -1592 5729 -1580 5905
rect -1546 5729 -1530 5905
rect -1592 5717 -1530 5729
rect -1500 5905 -1438 5917
rect -1500 5729 -1484 5905
rect -1450 5729 -1438 5905
rect -1500 5717 -1438 5729
rect -1382 5905 -1320 5917
rect -1382 5729 -1370 5905
rect -1336 5729 -1320 5905
rect -1382 5717 -1320 5729
rect -1290 5905 -1228 5917
rect -1290 5729 -1274 5905
rect -1240 5729 -1228 5905
rect -1290 5717 -1228 5729
rect -1172 5905 -1110 5917
rect -1172 5729 -1160 5905
rect -1126 5729 -1110 5905
rect -1172 5717 -1110 5729
rect -1080 5905 -1018 5917
rect -1080 5729 -1064 5905
rect -1030 5729 -1018 5905
rect -1080 5717 -1018 5729
rect -962 5905 -900 5917
rect -962 5729 -950 5905
rect -916 5729 -900 5905
rect -962 5717 -900 5729
rect -870 5905 -808 5917
rect -870 5729 -854 5905
rect -820 5729 -808 5905
rect -870 5717 -808 5729
rect -752 5905 -690 5917
rect -752 5729 -740 5905
rect -706 5729 -690 5905
rect -752 5717 -690 5729
rect -660 5905 -598 5917
rect -660 5729 -644 5905
rect -610 5729 -598 5905
rect -660 5717 -598 5729
rect -542 5905 -480 5917
rect -542 5729 -530 5905
rect -496 5729 -480 5905
rect -542 5717 -480 5729
rect -450 5905 -388 5917
rect -450 5729 -434 5905
rect -400 5729 -388 5905
rect -450 5717 -388 5729
rect -332 5905 -270 5917
rect -332 5729 -320 5905
rect -286 5729 -270 5905
rect -332 5717 -270 5729
rect -240 5905 -178 5917
rect -240 5729 -224 5905
rect -190 5729 -178 5905
rect -240 5717 -178 5729
rect -122 5905 -60 5917
rect -122 5729 -110 5905
rect -76 5729 -60 5905
rect -122 5717 -60 5729
rect -30 5905 32 5917
rect -30 5729 -14 5905
rect 20 5729 32 5905
rect -30 5717 32 5729
rect 88 5905 150 5917
rect 88 5729 100 5905
rect 134 5729 150 5905
rect 88 5717 150 5729
rect 180 5905 242 5917
rect 180 5729 196 5905
rect 230 5729 242 5905
rect 180 5717 242 5729
rect 298 5905 360 5917
rect 298 5729 310 5905
rect 344 5729 360 5905
rect 298 5717 360 5729
rect 390 5905 452 5917
rect 390 5729 406 5905
rect 440 5729 452 5905
rect 390 5717 452 5729
rect 508 5905 570 5917
rect 508 5729 520 5905
rect 554 5729 570 5905
rect 508 5717 570 5729
rect 600 5905 662 5917
rect 600 5729 616 5905
rect 650 5729 662 5905
rect 600 5717 662 5729
rect 718 5905 780 5917
rect 718 5729 730 5905
rect 764 5729 780 5905
rect 718 5717 780 5729
rect 810 5905 872 5917
rect 810 5729 826 5905
rect 860 5729 872 5905
rect 810 5717 872 5729
rect 928 5905 990 5917
rect 928 5729 940 5905
rect 974 5729 990 5905
rect 928 5717 990 5729
rect 1020 5905 1082 5917
rect 1020 5729 1036 5905
rect 1070 5729 1082 5905
rect 1020 5717 1082 5729
rect 1138 5905 1200 5917
rect 1138 5729 1150 5905
rect 1184 5729 1200 5905
rect 1138 5717 1200 5729
rect 1230 5905 1292 5917
rect 1230 5729 1246 5905
rect 1280 5729 1292 5905
rect 1230 5717 1292 5729
rect 1348 5905 1410 5917
rect 1348 5729 1360 5905
rect 1394 5729 1410 5905
rect 1348 5717 1410 5729
rect 1440 5905 1502 5917
rect 1440 5729 1456 5905
rect 1490 5729 1502 5905
rect 1440 5717 1502 5729
rect 1558 5905 1620 5917
rect 1558 5729 1570 5905
rect 1604 5729 1620 5905
rect 1558 5717 1620 5729
rect 1650 5905 1712 5917
rect 1650 5729 1666 5905
rect 1700 5729 1712 5905
rect 1650 5717 1712 5729
rect 1768 5905 1830 5917
rect 1768 5729 1780 5905
rect 1814 5729 1830 5905
rect 1768 5717 1830 5729
rect 1860 5905 1922 5917
rect 1860 5729 1876 5905
rect 1910 5729 1922 5905
rect 1860 5717 1922 5729
rect 1978 5905 2040 5917
rect 1978 5729 1990 5905
rect 2024 5729 2040 5905
rect 1978 5717 2040 5729
rect 2070 5905 2132 5917
rect 2070 5729 2086 5905
rect 2120 5729 2132 5905
rect 2070 5717 2132 5729
rect 2188 5905 2250 5917
rect 2188 5729 2200 5905
rect 2234 5729 2250 5905
rect 2188 5717 2250 5729
rect 2280 5905 2342 5917
rect 2280 5729 2296 5905
rect 2330 5729 2342 5905
rect 2280 5717 2342 5729
rect 2398 5905 2460 5917
rect 2398 5729 2410 5905
rect 2444 5729 2460 5905
rect 2398 5717 2460 5729
rect 2490 5905 2552 5917
rect 2490 5729 2506 5905
rect 2540 5729 2552 5905
rect 2490 5717 2552 5729
rect 2608 5905 2670 5917
rect 2608 5729 2620 5905
rect 2654 5729 2670 5905
rect 2608 5717 2670 5729
rect 2700 5905 2762 5917
rect 2700 5729 2716 5905
rect 2750 5729 2762 5905
rect 2700 5717 2762 5729
rect 2818 5905 2880 5917
rect 2818 5729 2830 5905
rect 2864 5729 2880 5905
rect 2818 5717 2880 5729
rect 2910 5905 2972 5917
rect 2910 5729 2926 5905
rect 2960 5729 2972 5905
rect 2910 5717 2972 5729
rect 3028 5905 3090 5917
rect 3028 5729 3040 5905
rect 3074 5729 3090 5905
rect 3028 5717 3090 5729
rect 3120 5905 3182 5917
rect 3120 5729 3136 5905
rect 3170 5729 3182 5905
rect 3120 5717 3182 5729
rect 3238 5905 3300 5917
rect 3238 5729 3250 5905
rect 3284 5729 3300 5905
rect 3238 5717 3300 5729
rect 3330 5905 3392 5917
rect 3330 5729 3346 5905
rect 3380 5729 3392 5905
rect 3330 5717 3392 5729
rect 3448 5905 3510 5917
rect 3448 5729 3460 5905
rect 3494 5729 3510 5905
rect 3448 5717 3510 5729
rect 3540 5905 3602 5917
rect 3540 5729 3556 5905
rect 3590 5729 3602 5905
rect 3540 5717 3602 5729
rect 3658 5905 3720 5917
rect 3658 5729 3670 5905
rect 3704 5729 3720 5905
rect 3658 5717 3720 5729
rect 3750 5905 3812 5917
rect 3750 5729 3766 5905
rect 3800 5729 3812 5905
rect 3750 5717 3812 5729
rect 3868 5905 3930 5917
rect 3868 5729 3880 5905
rect 3914 5729 3930 5905
rect 3868 5717 3930 5729
rect 3960 5905 4022 5917
rect 3960 5729 3976 5905
rect 4010 5729 4022 5905
rect 3960 5717 4022 5729
rect 4078 5905 4140 5917
rect 4078 5729 4090 5905
rect 4124 5729 4140 5905
rect 4078 5717 4140 5729
rect 4170 5905 4232 5917
rect 4170 5729 4186 5905
rect 4220 5729 4232 5905
rect 4170 5717 4232 5729
rect 4288 5905 4350 5917
rect 4288 5729 4300 5905
rect 4334 5729 4350 5905
rect 4288 5717 4350 5729
rect 4380 5905 4442 5917
rect 4380 5729 4396 5905
rect 4430 5729 4442 5905
rect 4380 5717 4442 5729
rect 4498 5905 4560 5917
rect 4498 5729 4510 5905
rect 4544 5729 4560 5905
rect 4498 5717 4560 5729
rect 4590 5905 4652 5917
rect 4590 5729 4606 5905
rect 4640 5729 4652 5905
rect 4590 5717 4652 5729
rect 4708 5905 4770 5917
rect 4708 5729 4720 5905
rect 4754 5729 4770 5905
rect 4708 5717 4770 5729
rect 4800 5905 4862 5917
rect 4800 5729 4816 5905
rect 4850 5729 4862 5905
rect 4800 5717 4862 5729
rect 4918 5905 4980 5917
rect 4918 5729 4930 5905
rect 4964 5729 4980 5905
rect 4918 5717 4980 5729
rect 5010 5905 5072 5917
rect 5010 5729 5026 5905
rect 5060 5729 5072 5905
rect 5010 5717 5072 5729
rect 5128 5905 5190 5917
rect 5128 5729 5140 5905
rect 5174 5729 5190 5905
rect 5128 5717 5190 5729
rect 5220 5905 5282 5917
rect 5220 5729 5236 5905
rect 5270 5729 5282 5905
rect 5220 5717 5282 5729
rect 5338 5905 5400 5917
rect 5338 5729 5350 5905
rect 5384 5729 5400 5905
rect 5338 5717 5400 5729
rect 5430 5905 5492 5917
rect 5430 5729 5446 5905
rect 5480 5729 5492 5905
rect 5430 5717 5492 5729
rect 5548 5905 5610 5917
rect 5548 5729 5560 5905
rect 5594 5729 5610 5905
rect 5548 5717 5610 5729
rect 5640 5905 5702 5917
rect 5640 5729 5656 5905
rect 5690 5729 5702 5905
rect 5640 5717 5702 5729
rect 5758 5905 5820 5917
rect 5758 5729 5770 5905
rect 5804 5729 5820 5905
rect 5758 5717 5820 5729
rect 5850 5905 5912 5917
rect 5850 5729 5866 5905
rect 5900 5729 5912 5905
rect 5850 5717 5912 5729
rect 5968 5905 6030 5917
rect 5968 5729 5980 5905
rect 6014 5729 6030 5905
rect 5968 5717 6030 5729
rect 6060 5905 6122 5917
rect 6060 5729 6076 5905
rect 6110 5729 6122 5905
rect 6060 5717 6122 5729
rect -2642 5465 -2580 5477
rect -2642 5289 -2630 5465
rect -2596 5289 -2580 5465
rect -2642 5277 -2580 5289
rect -2550 5465 -2488 5477
rect -2550 5289 -2534 5465
rect -2500 5289 -2488 5465
rect -2550 5277 -2488 5289
rect -2432 5465 -2370 5477
rect -2432 5289 -2420 5465
rect -2386 5289 -2370 5465
rect -2432 5277 -2370 5289
rect -2340 5465 -2278 5477
rect -2340 5289 -2324 5465
rect -2290 5289 -2278 5465
rect -2340 5277 -2278 5289
rect -2222 5465 -2160 5477
rect -2222 5289 -2210 5465
rect -2176 5289 -2160 5465
rect -2222 5277 -2160 5289
rect -2130 5465 -2068 5477
rect -2130 5289 -2114 5465
rect -2080 5289 -2068 5465
rect -2130 5277 -2068 5289
rect -2012 5465 -1950 5477
rect -2012 5289 -2000 5465
rect -1966 5289 -1950 5465
rect -2012 5277 -1950 5289
rect -1920 5465 -1858 5477
rect -1920 5289 -1904 5465
rect -1870 5289 -1858 5465
rect -1920 5277 -1858 5289
rect -1802 5465 -1740 5477
rect -1802 5289 -1790 5465
rect -1756 5289 -1740 5465
rect -1802 5277 -1740 5289
rect -1710 5465 -1648 5477
rect -1710 5289 -1694 5465
rect -1660 5289 -1648 5465
rect -1710 5277 -1648 5289
rect -1592 5465 -1530 5477
rect -1592 5289 -1580 5465
rect -1546 5289 -1530 5465
rect -1592 5277 -1530 5289
rect -1500 5465 -1438 5477
rect -1500 5289 -1484 5465
rect -1450 5289 -1438 5465
rect -1500 5277 -1438 5289
rect -1382 5465 -1320 5477
rect -1382 5289 -1370 5465
rect -1336 5289 -1320 5465
rect -1382 5277 -1320 5289
rect -1290 5465 -1228 5477
rect -1290 5289 -1274 5465
rect -1240 5289 -1228 5465
rect -1290 5277 -1228 5289
rect -1172 5465 -1110 5477
rect -1172 5289 -1160 5465
rect -1126 5289 -1110 5465
rect -1172 5277 -1110 5289
rect -1080 5465 -1018 5477
rect -1080 5289 -1064 5465
rect -1030 5289 -1018 5465
rect -1080 5277 -1018 5289
rect -962 5465 -900 5477
rect -962 5289 -950 5465
rect -916 5289 -900 5465
rect -962 5277 -900 5289
rect -870 5465 -808 5477
rect -870 5289 -854 5465
rect -820 5289 -808 5465
rect -870 5277 -808 5289
rect -752 5465 -690 5477
rect -752 5289 -740 5465
rect -706 5289 -690 5465
rect -752 5277 -690 5289
rect -660 5465 -598 5477
rect -660 5289 -644 5465
rect -610 5289 -598 5465
rect -660 5277 -598 5289
rect -542 5465 -480 5477
rect -542 5289 -530 5465
rect -496 5289 -480 5465
rect -542 5277 -480 5289
rect -450 5465 -388 5477
rect -450 5289 -434 5465
rect -400 5289 -388 5465
rect -450 5277 -388 5289
rect -332 5465 -270 5477
rect -332 5289 -320 5465
rect -286 5289 -270 5465
rect -332 5277 -270 5289
rect -240 5465 -178 5477
rect -240 5289 -224 5465
rect -190 5289 -178 5465
rect -240 5277 -178 5289
rect -122 5465 -60 5477
rect -122 5289 -110 5465
rect -76 5289 -60 5465
rect -122 5277 -60 5289
rect -30 5465 32 5477
rect -30 5289 -14 5465
rect 20 5289 32 5465
rect -30 5277 32 5289
rect 88 5465 150 5477
rect 88 5289 100 5465
rect 134 5289 150 5465
rect 88 5277 150 5289
rect 180 5465 242 5477
rect 180 5289 196 5465
rect 230 5289 242 5465
rect 180 5277 242 5289
rect 298 5465 360 5477
rect 298 5289 310 5465
rect 344 5289 360 5465
rect 298 5277 360 5289
rect 390 5465 452 5477
rect 390 5289 406 5465
rect 440 5289 452 5465
rect 390 5277 452 5289
rect 508 5465 570 5477
rect 508 5289 520 5465
rect 554 5289 570 5465
rect 508 5277 570 5289
rect 600 5465 662 5477
rect 600 5289 616 5465
rect 650 5289 662 5465
rect 600 5277 662 5289
rect 718 5465 780 5477
rect 718 5289 730 5465
rect 764 5289 780 5465
rect 718 5277 780 5289
rect 810 5465 872 5477
rect 810 5289 826 5465
rect 860 5289 872 5465
rect 810 5277 872 5289
rect 928 5465 990 5477
rect 928 5289 940 5465
rect 974 5289 990 5465
rect 928 5277 990 5289
rect 1020 5465 1082 5477
rect 1020 5289 1036 5465
rect 1070 5289 1082 5465
rect 1020 5277 1082 5289
rect 1138 5465 1200 5477
rect 1138 5289 1150 5465
rect 1184 5289 1200 5465
rect 1138 5277 1200 5289
rect 1230 5465 1292 5477
rect 1230 5289 1246 5465
rect 1280 5289 1292 5465
rect 1230 5277 1292 5289
rect 1348 5465 1410 5477
rect 1348 5289 1360 5465
rect 1394 5289 1410 5465
rect 1348 5277 1410 5289
rect 1440 5465 1502 5477
rect 1440 5289 1456 5465
rect 1490 5289 1502 5465
rect 1440 5277 1502 5289
rect 1558 5465 1620 5477
rect 1558 5289 1570 5465
rect 1604 5289 1620 5465
rect 1558 5277 1620 5289
rect 1650 5465 1712 5477
rect 1650 5289 1666 5465
rect 1700 5289 1712 5465
rect 1650 5277 1712 5289
rect 1768 5465 1830 5477
rect 1768 5289 1780 5465
rect 1814 5289 1830 5465
rect 1768 5277 1830 5289
rect 1860 5465 1922 5477
rect 1860 5289 1876 5465
rect 1910 5289 1922 5465
rect 1860 5277 1922 5289
rect 1978 5465 2040 5477
rect 1978 5289 1990 5465
rect 2024 5289 2040 5465
rect 1978 5277 2040 5289
rect 2070 5465 2132 5477
rect 2070 5289 2086 5465
rect 2120 5289 2132 5465
rect 2070 5277 2132 5289
rect 2188 5465 2250 5477
rect 2188 5289 2200 5465
rect 2234 5289 2250 5465
rect 2188 5277 2250 5289
rect 2280 5465 2342 5477
rect 2280 5289 2296 5465
rect 2330 5289 2342 5465
rect 2280 5277 2342 5289
rect 2398 5465 2460 5477
rect 2398 5289 2410 5465
rect 2444 5289 2460 5465
rect 2398 5277 2460 5289
rect 2490 5465 2552 5477
rect 2490 5289 2506 5465
rect 2540 5289 2552 5465
rect 2490 5277 2552 5289
rect 2608 5465 2670 5477
rect 2608 5289 2620 5465
rect 2654 5289 2670 5465
rect 2608 5277 2670 5289
rect 2700 5465 2762 5477
rect 2700 5289 2716 5465
rect 2750 5289 2762 5465
rect 2700 5277 2762 5289
rect 2818 5465 2880 5477
rect 2818 5289 2830 5465
rect 2864 5289 2880 5465
rect 2818 5277 2880 5289
rect 2910 5465 2972 5477
rect 2910 5289 2926 5465
rect 2960 5289 2972 5465
rect 2910 5277 2972 5289
rect 3028 5465 3090 5477
rect 3028 5289 3040 5465
rect 3074 5289 3090 5465
rect 3028 5277 3090 5289
rect 3120 5465 3182 5477
rect 3120 5289 3136 5465
rect 3170 5289 3182 5465
rect 3120 5277 3182 5289
rect 3238 5465 3300 5477
rect 3238 5289 3250 5465
rect 3284 5289 3300 5465
rect 3238 5277 3300 5289
rect 3330 5465 3392 5477
rect 3330 5289 3346 5465
rect 3380 5289 3392 5465
rect 3330 5277 3392 5289
rect 3448 5465 3510 5477
rect 3448 5289 3460 5465
rect 3494 5289 3510 5465
rect 3448 5277 3510 5289
rect 3540 5465 3602 5477
rect 3540 5289 3556 5465
rect 3590 5289 3602 5465
rect 3540 5277 3602 5289
rect 3658 5465 3720 5477
rect 3658 5289 3670 5465
rect 3704 5289 3720 5465
rect 3658 5277 3720 5289
rect 3750 5465 3812 5477
rect 3750 5289 3766 5465
rect 3800 5289 3812 5465
rect 3750 5277 3812 5289
rect 3868 5465 3930 5477
rect 3868 5289 3880 5465
rect 3914 5289 3930 5465
rect 3868 5277 3930 5289
rect 3960 5465 4022 5477
rect 3960 5289 3976 5465
rect 4010 5289 4022 5465
rect 3960 5277 4022 5289
rect 4078 5465 4140 5477
rect 4078 5289 4090 5465
rect 4124 5289 4140 5465
rect 4078 5277 4140 5289
rect 4170 5465 4232 5477
rect 4170 5289 4186 5465
rect 4220 5289 4232 5465
rect 4170 5277 4232 5289
rect 4288 5465 4350 5477
rect 4288 5289 4300 5465
rect 4334 5289 4350 5465
rect 4288 5277 4350 5289
rect 4380 5465 4442 5477
rect 4380 5289 4396 5465
rect 4430 5289 4442 5465
rect 4380 5277 4442 5289
rect 4498 5465 4560 5477
rect 4498 5289 4510 5465
rect 4544 5289 4560 5465
rect 4498 5277 4560 5289
rect 4590 5465 4652 5477
rect 4590 5289 4606 5465
rect 4640 5289 4652 5465
rect 4590 5277 4652 5289
rect 4708 5465 4770 5477
rect 4708 5289 4720 5465
rect 4754 5289 4770 5465
rect 4708 5277 4770 5289
rect 4800 5465 4862 5477
rect 4800 5289 4816 5465
rect 4850 5289 4862 5465
rect 4800 5277 4862 5289
rect 4918 5465 4980 5477
rect 4918 5289 4930 5465
rect 4964 5289 4980 5465
rect 4918 5277 4980 5289
rect 5010 5465 5072 5477
rect 5010 5289 5026 5465
rect 5060 5289 5072 5465
rect 5010 5277 5072 5289
rect 5128 5465 5190 5477
rect 5128 5289 5140 5465
rect 5174 5289 5190 5465
rect 5128 5277 5190 5289
rect 5220 5465 5282 5477
rect 5220 5289 5236 5465
rect 5270 5289 5282 5465
rect 5220 5277 5282 5289
rect 5338 5465 5400 5477
rect 5338 5289 5350 5465
rect 5384 5289 5400 5465
rect 5338 5277 5400 5289
rect 5430 5465 5492 5477
rect 5430 5289 5446 5465
rect 5480 5289 5492 5465
rect 5430 5277 5492 5289
rect 5548 5465 5610 5477
rect 5548 5289 5560 5465
rect 5594 5289 5610 5465
rect 5548 5277 5610 5289
rect 5640 5465 5702 5477
rect 5640 5289 5656 5465
rect 5690 5289 5702 5465
rect 5640 5277 5702 5289
rect 5758 5465 5820 5477
rect 5758 5289 5770 5465
rect 5804 5289 5820 5465
rect 5758 5277 5820 5289
rect 5850 5465 5912 5477
rect 5850 5289 5866 5465
rect 5900 5289 5912 5465
rect 5850 5277 5912 5289
rect 5968 5465 6030 5477
rect 5968 5289 5980 5465
rect 6014 5289 6030 5465
rect 5968 5277 6030 5289
rect 6060 5465 6122 5477
rect 6060 5289 6076 5465
rect 6110 5289 6122 5465
rect 6060 5277 6122 5289
rect -2642 5025 -2580 5037
rect -2642 4849 -2630 5025
rect -2596 4849 -2580 5025
rect -2642 4837 -2580 4849
rect -2550 5025 -2488 5037
rect -2550 4849 -2534 5025
rect -2500 4849 -2488 5025
rect -2550 4837 -2488 4849
rect -2432 5025 -2370 5037
rect -2432 4849 -2420 5025
rect -2386 4849 -2370 5025
rect -2432 4837 -2370 4849
rect -2340 5025 -2278 5037
rect -2340 4849 -2324 5025
rect -2290 4849 -2278 5025
rect -2340 4837 -2278 4849
rect -2222 5025 -2160 5037
rect -2222 4849 -2210 5025
rect -2176 4849 -2160 5025
rect -2222 4837 -2160 4849
rect -2130 5025 -2068 5037
rect -2130 4849 -2114 5025
rect -2080 4849 -2068 5025
rect -2130 4837 -2068 4849
rect -2012 5025 -1950 5037
rect -2012 4849 -2000 5025
rect -1966 4849 -1950 5025
rect -2012 4837 -1950 4849
rect -1920 5025 -1858 5037
rect -1920 4849 -1904 5025
rect -1870 4849 -1858 5025
rect -1920 4837 -1858 4849
rect -1802 5025 -1740 5037
rect -1802 4849 -1790 5025
rect -1756 4849 -1740 5025
rect -1802 4837 -1740 4849
rect -1710 5025 -1648 5037
rect -1710 4849 -1694 5025
rect -1660 4849 -1648 5025
rect -1710 4837 -1648 4849
rect -1592 5025 -1530 5037
rect -1592 4849 -1580 5025
rect -1546 4849 -1530 5025
rect -1592 4837 -1530 4849
rect -1500 5025 -1438 5037
rect -1500 4849 -1484 5025
rect -1450 4849 -1438 5025
rect -1500 4837 -1438 4849
rect -1382 5025 -1320 5037
rect -1382 4849 -1370 5025
rect -1336 4849 -1320 5025
rect -1382 4837 -1320 4849
rect -1290 5025 -1228 5037
rect -1290 4849 -1274 5025
rect -1240 4849 -1228 5025
rect -1290 4837 -1228 4849
rect -1172 5025 -1110 5037
rect -1172 4849 -1160 5025
rect -1126 4849 -1110 5025
rect -1172 4837 -1110 4849
rect -1080 5025 -1018 5037
rect -1080 4849 -1064 5025
rect -1030 4849 -1018 5025
rect -1080 4837 -1018 4849
rect -962 5025 -900 5037
rect -962 4849 -950 5025
rect -916 4849 -900 5025
rect -962 4837 -900 4849
rect -870 5025 -808 5037
rect -870 4849 -854 5025
rect -820 4849 -808 5025
rect -870 4837 -808 4849
rect -752 5025 -690 5037
rect -752 4849 -740 5025
rect -706 4849 -690 5025
rect -752 4837 -690 4849
rect -660 5025 -598 5037
rect -660 4849 -644 5025
rect -610 4849 -598 5025
rect -660 4837 -598 4849
rect -542 5025 -480 5037
rect -542 4849 -530 5025
rect -496 4849 -480 5025
rect -542 4837 -480 4849
rect -450 5025 -388 5037
rect -450 4849 -434 5025
rect -400 4849 -388 5025
rect -450 4837 -388 4849
rect -332 5025 -270 5037
rect -332 4849 -320 5025
rect -286 4849 -270 5025
rect -332 4837 -270 4849
rect -240 5025 -178 5037
rect -240 4849 -224 5025
rect -190 4849 -178 5025
rect -240 4837 -178 4849
rect -122 5025 -60 5037
rect -122 4849 -110 5025
rect -76 4849 -60 5025
rect -122 4837 -60 4849
rect -30 5025 32 5037
rect -30 4849 -14 5025
rect 20 4849 32 5025
rect -30 4837 32 4849
rect 88 5025 150 5037
rect 88 4849 100 5025
rect 134 4849 150 5025
rect 88 4837 150 4849
rect 180 5025 242 5037
rect 180 4849 196 5025
rect 230 4849 242 5025
rect 180 4837 242 4849
rect 298 5025 360 5037
rect 298 4849 310 5025
rect 344 4849 360 5025
rect 298 4837 360 4849
rect 390 5025 452 5037
rect 390 4849 406 5025
rect 440 4849 452 5025
rect 390 4837 452 4849
rect 508 5025 570 5037
rect 508 4849 520 5025
rect 554 4849 570 5025
rect 508 4837 570 4849
rect 600 5025 662 5037
rect 600 4849 616 5025
rect 650 4849 662 5025
rect 600 4837 662 4849
rect 718 5025 780 5037
rect 718 4849 730 5025
rect 764 4849 780 5025
rect 718 4837 780 4849
rect 810 5025 872 5037
rect 810 4849 826 5025
rect 860 4849 872 5025
rect 810 4837 872 4849
rect 928 5025 990 5037
rect 928 4849 940 5025
rect 974 4849 990 5025
rect 928 4837 990 4849
rect 1020 5025 1082 5037
rect 1020 4849 1036 5025
rect 1070 4849 1082 5025
rect 1020 4837 1082 4849
rect 1138 5025 1200 5037
rect 1138 4849 1150 5025
rect 1184 4849 1200 5025
rect 1138 4837 1200 4849
rect 1230 5025 1292 5037
rect 1230 4849 1246 5025
rect 1280 4849 1292 5025
rect 1230 4837 1292 4849
rect 1348 5025 1410 5037
rect 1348 4849 1360 5025
rect 1394 4849 1410 5025
rect 1348 4837 1410 4849
rect 1440 5025 1502 5037
rect 1440 4849 1456 5025
rect 1490 4849 1502 5025
rect 1440 4837 1502 4849
rect 1558 5025 1620 5037
rect 1558 4849 1570 5025
rect 1604 4849 1620 5025
rect 1558 4837 1620 4849
rect 1650 5025 1712 5037
rect 1650 4849 1666 5025
rect 1700 4849 1712 5025
rect 1650 4837 1712 4849
rect 1768 5025 1830 5037
rect 1768 4849 1780 5025
rect 1814 4849 1830 5025
rect 1768 4837 1830 4849
rect 1860 5025 1922 5037
rect 1860 4849 1876 5025
rect 1910 4849 1922 5025
rect 1860 4837 1922 4849
rect 1978 5025 2040 5037
rect 1978 4849 1990 5025
rect 2024 4849 2040 5025
rect 1978 4837 2040 4849
rect 2070 5025 2132 5037
rect 2070 4849 2086 5025
rect 2120 4849 2132 5025
rect 2070 4837 2132 4849
rect 2188 5025 2250 5037
rect 2188 4849 2200 5025
rect 2234 4849 2250 5025
rect 2188 4837 2250 4849
rect 2280 5025 2342 5037
rect 2280 4849 2296 5025
rect 2330 4849 2342 5025
rect 2280 4837 2342 4849
rect 2398 5025 2460 5037
rect 2398 4849 2410 5025
rect 2444 4849 2460 5025
rect 2398 4837 2460 4849
rect 2490 5025 2552 5037
rect 2490 4849 2506 5025
rect 2540 4849 2552 5025
rect 2490 4837 2552 4849
rect 2608 5025 2670 5037
rect 2608 4849 2620 5025
rect 2654 4849 2670 5025
rect 2608 4837 2670 4849
rect 2700 5025 2762 5037
rect 2700 4849 2716 5025
rect 2750 4849 2762 5025
rect 2700 4837 2762 4849
rect 2818 5025 2880 5037
rect 2818 4849 2830 5025
rect 2864 4849 2880 5025
rect 2818 4837 2880 4849
rect 2910 5025 2972 5037
rect 2910 4849 2926 5025
rect 2960 4849 2972 5025
rect 2910 4837 2972 4849
rect 3028 5025 3090 5037
rect 3028 4849 3040 5025
rect 3074 4849 3090 5025
rect 3028 4837 3090 4849
rect 3120 5025 3182 5037
rect 3120 4849 3136 5025
rect 3170 4849 3182 5025
rect 3120 4837 3182 4849
rect 3238 5025 3300 5037
rect 3238 4849 3250 5025
rect 3284 4849 3300 5025
rect 3238 4837 3300 4849
rect 3330 5025 3392 5037
rect 3330 4849 3346 5025
rect 3380 4849 3392 5025
rect 3330 4837 3392 4849
rect 3448 5025 3510 5037
rect 3448 4849 3460 5025
rect 3494 4849 3510 5025
rect 3448 4837 3510 4849
rect 3540 5025 3602 5037
rect 3540 4849 3556 5025
rect 3590 4849 3602 5025
rect 3540 4837 3602 4849
rect 3658 5025 3720 5037
rect 3658 4849 3670 5025
rect 3704 4849 3720 5025
rect 3658 4837 3720 4849
rect 3750 5025 3812 5037
rect 3750 4849 3766 5025
rect 3800 4849 3812 5025
rect 3750 4837 3812 4849
rect 3868 5025 3930 5037
rect 3868 4849 3880 5025
rect 3914 4849 3930 5025
rect 3868 4837 3930 4849
rect 3960 5025 4022 5037
rect 3960 4849 3976 5025
rect 4010 4849 4022 5025
rect 3960 4837 4022 4849
rect 4078 5025 4140 5037
rect 4078 4849 4090 5025
rect 4124 4849 4140 5025
rect 4078 4837 4140 4849
rect 4170 5025 4232 5037
rect 4170 4849 4186 5025
rect 4220 4849 4232 5025
rect 4170 4837 4232 4849
rect 4288 5025 4350 5037
rect 4288 4849 4300 5025
rect 4334 4849 4350 5025
rect 4288 4837 4350 4849
rect 4380 5025 4442 5037
rect 4380 4849 4396 5025
rect 4430 4849 4442 5025
rect 4380 4837 4442 4849
rect 4498 5025 4560 5037
rect 4498 4849 4510 5025
rect 4544 4849 4560 5025
rect 4498 4837 4560 4849
rect 4590 5025 4652 5037
rect 4590 4849 4606 5025
rect 4640 4849 4652 5025
rect 4590 4837 4652 4849
rect 4708 5025 4770 5037
rect 4708 4849 4720 5025
rect 4754 4849 4770 5025
rect 4708 4837 4770 4849
rect 4800 5025 4862 5037
rect 4800 4849 4816 5025
rect 4850 4849 4862 5025
rect 4800 4837 4862 4849
rect 4918 5025 4980 5037
rect 4918 4849 4930 5025
rect 4964 4849 4980 5025
rect 4918 4837 4980 4849
rect 5010 5025 5072 5037
rect 5010 4849 5026 5025
rect 5060 4849 5072 5025
rect 5010 4837 5072 4849
rect 5128 5025 5190 5037
rect 5128 4849 5140 5025
rect 5174 4849 5190 5025
rect 5128 4837 5190 4849
rect 5220 5025 5282 5037
rect 5220 4849 5236 5025
rect 5270 4849 5282 5025
rect 5220 4837 5282 4849
rect 5338 5025 5400 5037
rect 5338 4849 5350 5025
rect 5384 4849 5400 5025
rect 5338 4837 5400 4849
rect 5430 5025 5492 5037
rect 5430 4849 5446 5025
rect 5480 4849 5492 5025
rect 5430 4837 5492 4849
rect 5548 5025 5610 5037
rect 5548 4849 5560 5025
rect 5594 4849 5610 5025
rect 5548 4837 5610 4849
rect 5640 5025 5702 5037
rect 5640 4849 5656 5025
rect 5690 4849 5702 5025
rect 5640 4837 5702 4849
rect 5758 5025 5820 5037
rect 5758 4849 5770 5025
rect 5804 4849 5820 5025
rect 5758 4837 5820 4849
rect 5850 5025 5912 5037
rect 5850 4849 5866 5025
rect 5900 4849 5912 5025
rect 5850 4837 5912 4849
rect 5968 5025 6030 5037
rect 5968 4849 5980 5025
rect 6014 4849 6030 5025
rect 5968 4837 6030 4849
rect 6060 5025 6122 5037
rect 6060 4849 6076 5025
rect 6110 4849 6122 5025
rect 6060 4837 6122 4849
rect -2642 4090 -2580 4102
rect -2642 3914 -2630 4090
rect -2596 3914 -2580 4090
rect -2642 3902 -2580 3914
rect -2550 4090 -2488 4102
rect -2550 3914 -2534 4090
rect -2500 3914 -2488 4090
rect -2550 3902 -2488 3914
rect -2432 4090 -2370 4102
rect -2432 3914 -2420 4090
rect -2386 3914 -2370 4090
rect -2432 3902 -2370 3914
rect -2340 4090 -2278 4102
rect -2340 3914 -2324 4090
rect -2290 3914 -2278 4090
rect -2340 3902 -2278 3914
rect -2222 4090 -2160 4102
rect -2222 3914 -2210 4090
rect -2176 3914 -2160 4090
rect -2222 3902 -2160 3914
rect -2130 4090 -2068 4102
rect -2130 3914 -2114 4090
rect -2080 3914 -2068 4090
rect -2130 3902 -2068 3914
rect -2012 4090 -1950 4102
rect -2012 3914 -2000 4090
rect -1966 3914 -1950 4090
rect -2012 3902 -1950 3914
rect -1920 4090 -1858 4102
rect -1920 3914 -1904 4090
rect -1870 3914 -1858 4090
rect -1920 3902 -1858 3914
rect -1802 4090 -1740 4102
rect -1802 3914 -1790 4090
rect -1756 3914 -1740 4090
rect -1802 3902 -1740 3914
rect -1710 4090 -1648 4102
rect -1710 3914 -1694 4090
rect -1660 3914 -1648 4090
rect -1710 3902 -1648 3914
rect -1592 4090 -1530 4102
rect -1592 3914 -1580 4090
rect -1546 3914 -1530 4090
rect -1592 3902 -1530 3914
rect -1500 4090 -1438 4102
rect -1500 3914 -1484 4090
rect -1450 3914 -1438 4090
rect -1500 3902 -1438 3914
rect -1382 4090 -1320 4102
rect -1382 3914 -1370 4090
rect -1336 3914 -1320 4090
rect -1382 3902 -1320 3914
rect -1290 4090 -1228 4102
rect -1290 3914 -1274 4090
rect -1240 3914 -1228 4090
rect -1290 3902 -1228 3914
rect -1172 4090 -1110 4102
rect -1172 3914 -1160 4090
rect -1126 3914 -1110 4090
rect -1172 3902 -1110 3914
rect -1080 4090 -1018 4102
rect -1080 3914 -1064 4090
rect -1030 3914 -1018 4090
rect -1080 3902 -1018 3914
rect -962 4090 -900 4102
rect -962 3914 -950 4090
rect -916 3914 -900 4090
rect -962 3902 -900 3914
rect -870 4090 -808 4102
rect -870 3914 -854 4090
rect -820 3914 -808 4090
rect -870 3902 -808 3914
rect -752 4090 -690 4102
rect -752 3914 -740 4090
rect -706 3914 -690 4090
rect -752 3902 -690 3914
rect -660 4090 -598 4102
rect -660 3914 -644 4090
rect -610 3914 -598 4090
rect -660 3902 -598 3914
rect -542 4090 -480 4102
rect -542 3914 -530 4090
rect -496 3914 -480 4090
rect -542 3902 -480 3914
rect -450 4090 -388 4102
rect -450 3914 -434 4090
rect -400 3914 -388 4090
rect -450 3902 -388 3914
rect -332 4090 -270 4102
rect -332 3914 -320 4090
rect -286 3914 -270 4090
rect -332 3902 -270 3914
rect -240 4090 -178 4102
rect -240 3914 -224 4090
rect -190 3914 -178 4090
rect -240 3902 -178 3914
rect -122 4090 -60 4102
rect -122 3914 -110 4090
rect -76 3914 -60 4090
rect -122 3902 -60 3914
rect -30 4090 32 4102
rect -30 3914 -14 4090
rect 20 3914 32 4090
rect -30 3902 32 3914
rect 88 4090 150 4102
rect 88 3914 100 4090
rect 134 3914 150 4090
rect 88 3902 150 3914
rect 180 4090 242 4102
rect 180 3914 196 4090
rect 230 3914 242 4090
rect 180 3902 242 3914
rect 298 4090 360 4102
rect 298 3914 310 4090
rect 344 3914 360 4090
rect 298 3902 360 3914
rect 390 4090 452 4102
rect 390 3914 406 4090
rect 440 3914 452 4090
rect 390 3902 452 3914
rect 508 4090 570 4102
rect 508 3914 520 4090
rect 554 3914 570 4090
rect 508 3902 570 3914
rect 600 4090 662 4102
rect 600 3914 616 4090
rect 650 3914 662 4090
rect 600 3902 662 3914
rect 718 4090 780 4102
rect 718 3914 730 4090
rect 764 3914 780 4090
rect 718 3902 780 3914
rect 810 4090 872 4102
rect 810 3914 826 4090
rect 860 3914 872 4090
rect 810 3902 872 3914
rect 928 4090 990 4102
rect 928 3914 940 4090
rect 974 3914 990 4090
rect 928 3902 990 3914
rect 1020 4090 1082 4102
rect 1020 3914 1036 4090
rect 1070 3914 1082 4090
rect 1020 3902 1082 3914
rect 1138 4090 1200 4102
rect 1138 3914 1150 4090
rect 1184 3914 1200 4090
rect 1138 3902 1200 3914
rect 1230 4090 1292 4102
rect 1230 3914 1246 4090
rect 1280 3914 1292 4090
rect 1230 3902 1292 3914
rect 1348 4090 1410 4102
rect 1348 3914 1360 4090
rect 1394 3914 1410 4090
rect 1348 3902 1410 3914
rect 1440 4090 1502 4102
rect 1440 3914 1456 4090
rect 1490 3914 1502 4090
rect 1440 3902 1502 3914
rect 1558 4090 1620 4102
rect 1558 3914 1570 4090
rect 1604 3914 1620 4090
rect 1558 3902 1620 3914
rect 1650 4090 1712 4102
rect 1650 3914 1666 4090
rect 1700 3914 1712 4090
rect 1650 3902 1712 3914
rect 1768 4090 1830 4102
rect 1768 3914 1780 4090
rect 1814 3914 1830 4090
rect 1768 3902 1830 3914
rect 1860 4090 1922 4102
rect 1860 3914 1876 4090
rect 1910 3914 1922 4090
rect 1860 3902 1922 3914
rect 1978 4090 2040 4102
rect 1978 3914 1990 4090
rect 2024 3914 2040 4090
rect 1978 3902 2040 3914
rect 2070 4090 2132 4102
rect 2070 3914 2086 4090
rect 2120 3914 2132 4090
rect 2070 3902 2132 3914
rect 2188 4090 2250 4102
rect 2188 3914 2200 4090
rect 2234 3914 2250 4090
rect 2188 3902 2250 3914
rect 2280 4090 2342 4102
rect 2280 3914 2296 4090
rect 2330 3914 2342 4090
rect 2280 3902 2342 3914
rect 2398 4090 2460 4102
rect 2398 3914 2410 4090
rect 2444 3914 2460 4090
rect 2398 3902 2460 3914
rect 2490 4090 2552 4102
rect 2490 3914 2506 4090
rect 2540 3914 2552 4090
rect 2490 3902 2552 3914
rect 2608 4090 2670 4102
rect 2608 3914 2620 4090
rect 2654 3914 2670 4090
rect 2608 3902 2670 3914
rect 2700 4090 2762 4102
rect 2700 3914 2716 4090
rect 2750 3914 2762 4090
rect 2700 3902 2762 3914
rect 2818 4090 2880 4102
rect 2818 3914 2830 4090
rect 2864 3914 2880 4090
rect 2818 3902 2880 3914
rect 2910 4090 2972 4102
rect 2910 3914 2926 4090
rect 2960 3914 2972 4090
rect 2910 3902 2972 3914
rect 3028 4090 3090 4102
rect 3028 3914 3040 4090
rect 3074 3914 3090 4090
rect 3028 3902 3090 3914
rect 3120 4090 3182 4102
rect 3120 3914 3136 4090
rect 3170 3914 3182 4090
rect 3120 3902 3182 3914
rect 3238 4090 3300 4102
rect 3238 3914 3250 4090
rect 3284 3914 3300 4090
rect 3238 3902 3300 3914
rect 3330 4090 3392 4102
rect 3330 3914 3346 4090
rect 3380 3914 3392 4090
rect 3330 3902 3392 3914
rect 3448 4090 3510 4102
rect 3448 3914 3460 4090
rect 3494 3914 3510 4090
rect 3448 3902 3510 3914
rect 3540 4090 3602 4102
rect 3540 3914 3556 4090
rect 3590 3914 3602 4090
rect 3540 3902 3602 3914
rect 3658 4090 3720 4102
rect 3658 3914 3670 4090
rect 3704 3914 3720 4090
rect 3658 3902 3720 3914
rect 3750 4090 3812 4102
rect 3750 3914 3766 4090
rect 3800 3914 3812 4090
rect 3750 3902 3812 3914
rect 3868 4090 3930 4102
rect 3868 3914 3880 4090
rect 3914 3914 3930 4090
rect 3868 3902 3930 3914
rect 3960 4090 4022 4102
rect 3960 3914 3976 4090
rect 4010 3914 4022 4090
rect 3960 3902 4022 3914
rect 4078 4090 4140 4102
rect 4078 3914 4090 4090
rect 4124 3914 4140 4090
rect 4078 3902 4140 3914
rect 4170 4090 4232 4102
rect 4170 3914 4186 4090
rect 4220 3914 4232 4090
rect 4170 3902 4232 3914
rect 4288 4090 4350 4102
rect 4288 3914 4300 4090
rect 4334 3914 4350 4090
rect 4288 3902 4350 3914
rect 4380 4090 4442 4102
rect 4380 3914 4396 4090
rect 4430 3914 4442 4090
rect 4380 3902 4442 3914
rect 4498 4090 4560 4102
rect 4498 3914 4510 4090
rect 4544 3914 4560 4090
rect 4498 3902 4560 3914
rect 4590 4090 4652 4102
rect 4590 3914 4606 4090
rect 4640 3914 4652 4090
rect 4590 3902 4652 3914
rect 4708 4090 4770 4102
rect 4708 3914 4720 4090
rect 4754 3914 4770 4090
rect 4708 3902 4770 3914
rect 4800 4090 4862 4102
rect 4800 3914 4816 4090
rect 4850 3914 4862 4090
rect 4800 3902 4862 3914
rect 4918 4090 4980 4102
rect 4918 3914 4930 4090
rect 4964 3914 4980 4090
rect 4918 3902 4980 3914
rect 5010 4090 5072 4102
rect 5010 3914 5026 4090
rect 5060 3914 5072 4090
rect 5010 3902 5072 3914
rect 5128 4090 5190 4102
rect 5128 3914 5140 4090
rect 5174 3914 5190 4090
rect 5128 3902 5190 3914
rect 5220 4090 5282 4102
rect 5220 3914 5236 4090
rect 5270 3914 5282 4090
rect 5220 3902 5282 3914
rect 5338 4090 5400 4102
rect 5338 3914 5350 4090
rect 5384 3914 5400 4090
rect 5338 3902 5400 3914
rect 5430 4090 5492 4102
rect 5430 3914 5446 4090
rect 5480 3914 5492 4090
rect 5430 3902 5492 3914
rect 5548 4090 5610 4102
rect 5548 3914 5560 4090
rect 5594 3914 5610 4090
rect 5548 3902 5610 3914
rect 5640 4090 5702 4102
rect 5640 3914 5656 4090
rect 5690 3914 5702 4090
rect 5640 3902 5702 3914
rect 5758 4090 5820 4102
rect 5758 3914 5770 4090
rect 5804 3914 5820 4090
rect 5758 3902 5820 3914
rect 5850 4090 5912 4102
rect 5850 3914 5866 4090
rect 5900 3914 5912 4090
rect 5850 3902 5912 3914
rect 5968 4090 6030 4102
rect 5968 3914 5980 4090
rect 6014 3914 6030 4090
rect 5968 3902 6030 3914
rect 6060 4090 6122 4102
rect 6060 3914 6076 4090
rect 6110 3914 6122 4090
rect 6060 3902 6122 3914
rect -2642 3650 -2580 3662
rect -2642 3474 -2630 3650
rect -2596 3474 -2580 3650
rect -2642 3462 -2580 3474
rect -2550 3650 -2488 3662
rect -2550 3474 -2534 3650
rect -2500 3474 -2488 3650
rect -2550 3462 -2488 3474
rect -2432 3650 -2370 3662
rect -2432 3474 -2420 3650
rect -2386 3474 -2370 3650
rect -2432 3462 -2370 3474
rect -2340 3650 -2278 3662
rect -2340 3474 -2324 3650
rect -2290 3474 -2278 3650
rect -2340 3462 -2278 3474
rect -2222 3650 -2160 3662
rect -2222 3474 -2210 3650
rect -2176 3474 -2160 3650
rect -2222 3462 -2160 3474
rect -2130 3650 -2068 3662
rect -2130 3474 -2114 3650
rect -2080 3474 -2068 3650
rect -2130 3462 -2068 3474
rect -2012 3650 -1950 3662
rect -2012 3474 -2000 3650
rect -1966 3474 -1950 3650
rect -2012 3462 -1950 3474
rect -1920 3650 -1858 3662
rect -1920 3474 -1904 3650
rect -1870 3474 -1858 3650
rect -1920 3462 -1858 3474
rect -1802 3650 -1740 3662
rect -1802 3474 -1790 3650
rect -1756 3474 -1740 3650
rect -1802 3462 -1740 3474
rect -1710 3650 -1648 3662
rect -1710 3474 -1694 3650
rect -1660 3474 -1648 3650
rect -1710 3462 -1648 3474
rect -1592 3650 -1530 3662
rect -1592 3474 -1580 3650
rect -1546 3474 -1530 3650
rect -1592 3462 -1530 3474
rect -1500 3650 -1438 3662
rect -1500 3474 -1484 3650
rect -1450 3474 -1438 3650
rect -1500 3462 -1438 3474
rect -1382 3650 -1320 3662
rect -1382 3474 -1370 3650
rect -1336 3474 -1320 3650
rect -1382 3462 -1320 3474
rect -1290 3650 -1228 3662
rect -1290 3474 -1274 3650
rect -1240 3474 -1228 3650
rect -1290 3462 -1228 3474
rect -1172 3650 -1110 3662
rect -1172 3474 -1160 3650
rect -1126 3474 -1110 3650
rect -1172 3462 -1110 3474
rect -1080 3650 -1018 3662
rect -1080 3474 -1064 3650
rect -1030 3474 -1018 3650
rect -1080 3462 -1018 3474
rect -962 3650 -900 3662
rect -962 3474 -950 3650
rect -916 3474 -900 3650
rect -962 3462 -900 3474
rect -870 3650 -808 3662
rect -870 3474 -854 3650
rect -820 3474 -808 3650
rect -870 3462 -808 3474
rect -752 3650 -690 3662
rect -752 3474 -740 3650
rect -706 3474 -690 3650
rect -752 3462 -690 3474
rect -660 3650 -598 3662
rect -660 3474 -644 3650
rect -610 3474 -598 3650
rect -660 3462 -598 3474
rect -542 3650 -480 3662
rect -542 3474 -530 3650
rect -496 3474 -480 3650
rect -542 3462 -480 3474
rect -450 3650 -388 3662
rect -450 3474 -434 3650
rect -400 3474 -388 3650
rect -450 3462 -388 3474
rect -332 3650 -270 3662
rect -332 3474 -320 3650
rect -286 3474 -270 3650
rect -332 3462 -270 3474
rect -240 3650 -178 3662
rect -240 3474 -224 3650
rect -190 3474 -178 3650
rect -240 3462 -178 3474
rect -122 3650 -60 3662
rect -122 3474 -110 3650
rect -76 3474 -60 3650
rect -122 3462 -60 3474
rect -30 3650 32 3662
rect -30 3474 -14 3650
rect 20 3474 32 3650
rect -30 3462 32 3474
rect 88 3650 150 3662
rect 88 3474 100 3650
rect 134 3474 150 3650
rect 88 3462 150 3474
rect 180 3650 242 3662
rect 180 3474 196 3650
rect 230 3474 242 3650
rect 180 3462 242 3474
rect 298 3650 360 3662
rect 298 3474 310 3650
rect 344 3474 360 3650
rect 298 3462 360 3474
rect 390 3650 452 3662
rect 390 3474 406 3650
rect 440 3474 452 3650
rect 390 3462 452 3474
rect 508 3650 570 3662
rect 508 3474 520 3650
rect 554 3474 570 3650
rect 508 3462 570 3474
rect 600 3650 662 3662
rect 600 3474 616 3650
rect 650 3474 662 3650
rect 600 3462 662 3474
rect 718 3650 780 3662
rect 718 3474 730 3650
rect 764 3474 780 3650
rect 718 3462 780 3474
rect 810 3650 872 3662
rect 810 3474 826 3650
rect 860 3474 872 3650
rect 810 3462 872 3474
rect 928 3650 990 3662
rect 928 3474 940 3650
rect 974 3474 990 3650
rect 928 3462 990 3474
rect 1020 3650 1082 3662
rect 1020 3474 1036 3650
rect 1070 3474 1082 3650
rect 1020 3462 1082 3474
rect 1138 3650 1200 3662
rect 1138 3474 1150 3650
rect 1184 3474 1200 3650
rect 1138 3462 1200 3474
rect 1230 3650 1292 3662
rect 1230 3474 1246 3650
rect 1280 3474 1292 3650
rect 1230 3462 1292 3474
rect 1348 3650 1410 3662
rect 1348 3474 1360 3650
rect 1394 3474 1410 3650
rect 1348 3462 1410 3474
rect 1440 3650 1502 3662
rect 1440 3474 1456 3650
rect 1490 3474 1502 3650
rect 1440 3462 1502 3474
rect 1558 3650 1620 3662
rect 1558 3474 1570 3650
rect 1604 3474 1620 3650
rect 1558 3462 1620 3474
rect 1650 3650 1712 3662
rect 1650 3474 1666 3650
rect 1700 3474 1712 3650
rect 1650 3462 1712 3474
rect 1768 3650 1830 3662
rect 1768 3474 1780 3650
rect 1814 3474 1830 3650
rect 1768 3462 1830 3474
rect 1860 3650 1922 3662
rect 1860 3474 1876 3650
rect 1910 3474 1922 3650
rect 1860 3462 1922 3474
rect 1978 3650 2040 3662
rect 1978 3474 1990 3650
rect 2024 3474 2040 3650
rect 1978 3462 2040 3474
rect 2070 3650 2132 3662
rect 2070 3474 2086 3650
rect 2120 3474 2132 3650
rect 2070 3462 2132 3474
rect 2188 3650 2250 3662
rect 2188 3474 2200 3650
rect 2234 3474 2250 3650
rect 2188 3462 2250 3474
rect 2280 3650 2342 3662
rect 2280 3474 2296 3650
rect 2330 3474 2342 3650
rect 2280 3462 2342 3474
rect 2398 3650 2460 3662
rect 2398 3474 2410 3650
rect 2444 3474 2460 3650
rect 2398 3462 2460 3474
rect 2490 3650 2552 3662
rect 2490 3474 2506 3650
rect 2540 3474 2552 3650
rect 2490 3462 2552 3474
rect 2608 3650 2670 3662
rect 2608 3474 2620 3650
rect 2654 3474 2670 3650
rect 2608 3462 2670 3474
rect 2700 3650 2762 3662
rect 2700 3474 2716 3650
rect 2750 3474 2762 3650
rect 2700 3462 2762 3474
rect 2818 3650 2880 3662
rect 2818 3474 2830 3650
rect 2864 3474 2880 3650
rect 2818 3462 2880 3474
rect 2910 3650 2972 3662
rect 2910 3474 2926 3650
rect 2960 3474 2972 3650
rect 2910 3462 2972 3474
rect 3028 3650 3090 3662
rect 3028 3474 3040 3650
rect 3074 3474 3090 3650
rect 3028 3462 3090 3474
rect 3120 3650 3182 3662
rect 3120 3474 3136 3650
rect 3170 3474 3182 3650
rect 3120 3462 3182 3474
rect 3238 3650 3300 3662
rect 3238 3474 3250 3650
rect 3284 3474 3300 3650
rect 3238 3462 3300 3474
rect 3330 3650 3392 3662
rect 3330 3474 3346 3650
rect 3380 3474 3392 3650
rect 3330 3462 3392 3474
rect 3448 3650 3510 3662
rect 3448 3474 3460 3650
rect 3494 3474 3510 3650
rect 3448 3462 3510 3474
rect 3540 3650 3602 3662
rect 3540 3474 3556 3650
rect 3590 3474 3602 3650
rect 3540 3462 3602 3474
rect 3658 3650 3720 3662
rect 3658 3474 3670 3650
rect 3704 3474 3720 3650
rect 3658 3462 3720 3474
rect 3750 3650 3812 3662
rect 3750 3474 3766 3650
rect 3800 3474 3812 3650
rect 3750 3462 3812 3474
rect 3868 3650 3930 3662
rect 3868 3474 3880 3650
rect 3914 3474 3930 3650
rect 3868 3462 3930 3474
rect 3960 3650 4022 3662
rect 3960 3474 3976 3650
rect 4010 3474 4022 3650
rect 3960 3462 4022 3474
rect 4078 3650 4140 3662
rect 4078 3474 4090 3650
rect 4124 3474 4140 3650
rect 4078 3462 4140 3474
rect 4170 3650 4232 3662
rect 4170 3474 4186 3650
rect 4220 3474 4232 3650
rect 4170 3462 4232 3474
rect 4288 3650 4350 3662
rect 4288 3474 4300 3650
rect 4334 3474 4350 3650
rect 4288 3462 4350 3474
rect 4380 3650 4442 3662
rect 4380 3474 4396 3650
rect 4430 3474 4442 3650
rect 4380 3462 4442 3474
rect 4498 3650 4560 3662
rect 4498 3474 4510 3650
rect 4544 3474 4560 3650
rect 4498 3462 4560 3474
rect 4590 3650 4652 3662
rect 4590 3474 4606 3650
rect 4640 3474 4652 3650
rect 4590 3462 4652 3474
rect 4708 3650 4770 3662
rect 4708 3474 4720 3650
rect 4754 3474 4770 3650
rect 4708 3462 4770 3474
rect 4800 3650 4862 3662
rect 4800 3474 4816 3650
rect 4850 3474 4862 3650
rect 4800 3462 4862 3474
rect 4918 3650 4980 3662
rect 4918 3474 4930 3650
rect 4964 3474 4980 3650
rect 4918 3462 4980 3474
rect 5010 3650 5072 3662
rect 5010 3474 5026 3650
rect 5060 3474 5072 3650
rect 5010 3462 5072 3474
rect 5128 3650 5190 3662
rect 5128 3474 5140 3650
rect 5174 3474 5190 3650
rect 5128 3462 5190 3474
rect 5220 3650 5282 3662
rect 5220 3474 5236 3650
rect 5270 3474 5282 3650
rect 5220 3462 5282 3474
rect 5338 3650 5400 3662
rect 5338 3474 5350 3650
rect 5384 3474 5400 3650
rect 5338 3462 5400 3474
rect 5430 3650 5492 3662
rect 5430 3474 5446 3650
rect 5480 3474 5492 3650
rect 5430 3462 5492 3474
rect 5548 3650 5610 3662
rect 5548 3474 5560 3650
rect 5594 3474 5610 3650
rect 5548 3462 5610 3474
rect 5640 3650 5702 3662
rect 5640 3474 5656 3650
rect 5690 3474 5702 3650
rect 5640 3462 5702 3474
rect 5758 3650 5820 3662
rect 5758 3474 5770 3650
rect 5804 3474 5820 3650
rect 5758 3462 5820 3474
rect 5850 3650 5912 3662
rect 5850 3474 5866 3650
rect 5900 3474 5912 3650
rect 5850 3462 5912 3474
rect 5968 3650 6030 3662
rect 5968 3474 5980 3650
rect 6014 3474 6030 3650
rect 5968 3462 6030 3474
rect 6060 3650 6122 3662
rect 6060 3474 6076 3650
rect 6110 3474 6122 3650
rect 6060 3462 6122 3474
rect -2642 3210 -2580 3222
rect -2642 3034 -2630 3210
rect -2596 3034 -2580 3210
rect -2642 3022 -2580 3034
rect -2550 3210 -2488 3222
rect -2550 3034 -2534 3210
rect -2500 3034 -2488 3210
rect -2550 3022 -2488 3034
rect -2432 3210 -2370 3222
rect -2432 3034 -2420 3210
rect -2386 3034 -2370 3210
rect -2432 3022 -2370 3034
rect -2340 3210 -2278 3222
rect -2340 3034 -2324 3210
rect -2290 3034 -2278 3210
rect -2340 3022 -2278 3034
rect -2222 3210 -2160 3222
rect -2222 3034 -2210 3210
rect -2176 3034 -2160 3210
rect -2222 3022 -2160 3034
rect -2130 3210 -2068 3222
rect -2130 3034 -2114 3210
rect -2080 3034 -2068 3210
rect -2130 3022 -2068 3034
rect -2012 3210 -1950 3222
rect -2012 3034 -2000 3210
rect -1966 3034 -1950 3210
rect -2012 3022 -1950 3034
rect -1920 3210 -1858 3222
rect -1920 3034 -1904 3210
rect -1870 3034 -1858 3210
rect -1920 3022 -1858 3034
rect -1802 3210 -1740 3222
rect -1802 3034 -1790 3210
rect -1756 3034 -1740 3210
rect -1802 3022 -1740 3034
rect -1710 3210 -1648 3222
rect -1710 3034 -1694 3210
rect -1660 3034 -1648 3210
rect -1710 3022 -1648 3034
rect -1592 3210 -1530 3222
rect -1592 3034 -1580 3210
rect -1546 3034 -1530 3210
rect -1592 3022 -1530 3034
rect -1500 3210 -1438 3222
rect -1500 3034 -1484 3210
rect -1450 3034 -1438 3210
rect -1500 3022 -1438 3034
rect -1382 3210 -1320 3222
rect -1382 3034 -1370 3210
rect -1336 3034 -1320 3210
rect -1382 3022 -1320 3034
rect -1290 3210 -1228 3222
rect -1290 3034 -1274 3210
rect -1240 3034 -1228 3210
rect -1290 3022 -1228 3034
rect -1172 3210 -1110 3222
rect -1172 3034 -1160 3210
rect -1126 3034 -1110 3210
rect -1172 3022 -1110 3034
rect -1080 3210 -1018 3222
rect -1080 3034 -1064 3210
rect -1030 3034 -1018 3210
rect -1080 3022 -1018 3034
rect -962 3210 -900 3222
rect -962 3034 -950 3210
rect -916 3034 -900 3210
rect -962 3022 -900 3034
rect -870 3210 -808 3222
rect -870 3034 -854 3210
rect -820 3034 -808 3210
rect -870 3022 -808 3034
rect -752 3210 -690 3222
rect -752 3034 -740 3210
rect -706 3034 -690 3210
rect -752 3022 -690 3034
rect -660 3210 -598 3222
rect -660 3034 -644 3210
rect -610 3034 -598 3210
rect -660 3022 -598 3034
rect -542 3210 -480 3222
rect -542 3034 -530 3210
rect -496 3034 -480 3210
rect -542 3022 -480 3034
rect -450 3210 -388 3222
rect -450 3034 -434 3210
rect -400 3034 -388 3210
rect -450 3022 -388 3034
rect -332 3210 -270 3222
rect -332 3034 -320 3210
rect -286 3034 -270 3210
rect -332 3022 -270 3034
rect -240 3210 -178 3222
rect -240 3034 -224 3210
rect -190 3034 -178 3210
rect -240 3022 -178 3034
rect -122 3210 -60 3222
rect -122 3034 -110 3210
rect -76 3034 -60 3210
rect -122 3022 -60 3034
rect -30 3210 32 3222
rect -30 3034 -14 3210
rect 20 3034 32 3210
rect -30 3022 32 3034
rect 88 3210 150 3222
rect 88 3034 100 3210
rect 134 3034 150 3210
rect 88 3022 150 3034
rect 180 3210 242 3222
rect 180 3034 196 3210
rect 230 3034 242 3210
rect 180 3022 242 3034
rect 298 3210 360 3222
rect 298 3034 310 3210
rect 344 3034 360 3210
rect 298 3022 360 3034
rect 390 3210 452 3222
rect 390 3034 406 3210
rect 440 3034 452 3210
rect 390 3022 452 3034
rect 508 3210 570 3222
rect 508 3034 520 3210
rect 554 3034 570 3210
rect 508 3022 570 3034
rect 600 3210 662 3222
rect 600 3034 616 3210
rect 650 3034 662 3210
rect 600 3022 662 3034
rect 718 3210 780 3222
rect 718 3034 730 3210
rect 764 3034 780 3210
rect 718 3022 780 3034
rect 810 3210 872 3222
rect 810 3034 826 3210
rect 860 3034 872 3210
rect 810 3022 872 3034
rect 928 3210 990 3222
rect 928 3034 940 3210
rect 974 3034 990 3210
rect 928 3022 990 3034
rect 1020 3210 1082 3222
rect 1020 3034 1036 3210
rect 1070 3034 1082 3210
rect 1020 3022 1082 3034
rect 1138 3210 1200 3222
rect 1138 3034 1150 3210
rect 1184 3034 1200 3210
rect 1138 3022 1200 3034
rect 1230 3210 1292 3222
rect 1230 3034 1246 3210
rect 1280 3034 1292 3210
rect 1230 3022 1292 3034
rect 1348 3210 1410 3222
rect 1348 3034 1360 3210
rect 1394 3034 1410 3210
rect 1348 3022 1410 3034
rect 1440 3210 1502 3222
rect 1440 3034 1456 3210
rect 1490 3034 1502 3210
rect 1440 3022 1502 3034
rect 1558 3210 1620 3222
rect 1558 3034 1570 3210
rect 1604 3034 1620 3210
rect 1558 3022 1620 3034
rect 1650 3210 1712 3222
rect 1650 3034 1666 3210
rect 1700 3034 1712 3210
rect 1650 3022 1712 3034
rect 1768 3210 1830 3222
rect 1768 3034 1780 3210
rect 1814 3034 1830 3210
rect 1768 3022 1830 3034
rect 1860 3210 1922 3222
rect 1860 3034 1876 3210
rect 1910 3034 1922 3210
rect 1860 3022 1922 3034
rect 1978 3210 2040 3222
rect 1978 3034 1990 3210
rect 2024 3034 2040 3210
rect 1978 3022 2040 3034
rect 2070 3210 2132 3222
rect 2070 3034 2086 3210
rect 2120 3034 2132 3210
rect 2070 3022 2132 3034
rect 2188 3210 2250 3222
rect 2188 3034 2200 3210
rect 2234 3034 2250 3210
rect 2188 3022 2250 3034
rect 2280 3210 2342 3222
rect 2280 3034 2296 3210
rect 2330 3034 2342 3210
rect 2280 3022 2342 3034
rect 2398 3210 2460 3222
rect 2398 3034 2410 3210
rect 2444 3034 2460 3210
rect 2398 3022 2460 3034
rect 2490 3210 2552 3222
rect 2490 3034 2506 3210
rect 2540 3034 2552 3210
rect 2490 3022 2552 3034
rect 2608 3210 2670 3222
rect 2608 3034 2620 3210
rect 2654 3034 2670 3210
rect 2608 3022 2670 3034
rect 2700 3210 2762 3222
rect 2700 3034 2716 3210
rect 2750 3034 2762 3210
rect 2700 3022 2762 3034
rect 2818 3210 2880 3222
rect 2818 3034 2830 3210
rect 2864 3034 2880 3210
rect 2818 3022 2880 3034
rect 2910 3210 2972 3222
rect 2910 3034 2926 3210
rect 2960 3034 2972 3210
rect 2910 3022 2972 3034
rect 3028 3210 3090 3222
rect 3028 3034 3040 3210
rect 3074 3034 3090 3210
rect 3028 3022 3090 3034
rect 3120 3210 3182 3222
rect 3120 3034 3136 3210
rect 3170 3034 3182 3210
rect 3120 3022 3182 3034
rect 3238 3210 3300 3222
rect 3238 3034 3250 3210
rect 3284 3034 3300 3210
rect 3238 3022 3300 3034
rect 3330 3210 3392 3222
rect 3330 3034 3346 3210
rect 3380 3034 3392 3210
rect 3330 3022 3392 3034
rect 3448 3210 3510 3222
rect 3448 3034 3460 3210
rect 3494 3034 3510 3210
rect 3448 3022 3510 3034
rect 3540 3210 3602 3222
rect 3540 3034 3556 3210
rect 3590 3034 3602 3210
rect 3540 3022 3602 3034
rect 3658 3210 3720 3222
rect 3658 3034 3670 3210
rect 3704 3034 3720 3210
rect 3658 3022 3720 3034
rect 3750 3210 3812 3222
rect 3750 3034 3766 3210
rect 3800 3034 3812 3210
rect 3750 3022 3812 3034
rect 3868 3210 3930 3222
rect 3868 3034 3880 3210
rect 3914 3034 3930 3210
rect 3868 3022 3930 3034
rect 3960 3210 4022 3222
rect 3960 3034 3976 3210
rect 4010 3034 4022 3210
rect 3960 3022 4022 3034
rect 4078 3210 4140 3222
rect 4078 3034 4090 3210
rect 4124 3034 4140 3210
rect 4078 3022 4140 3034
rect 4170 3210 4232 3222
rect 4170 3034 4186 3210
rect 4220 3034 4232 3210
rect 4170 3022 4232 3034
rect 4288 3210 4350 3222
rect 4288 3034 4300 3210
rect 4334 3034 4350 3210
rect 4288 3022 4350 3034
rect 4380 3210 4442 3222
rect 4380 3034 4396 3210
rect 4430 3034 4442 3210
rect 4380 3022 4442 3034
rect 4498 3210 4560 3222
rect 4498 3034 4510 3210
rect 4544 3034 4560 3210
rect 4498 3022 4560 3034
rect 4590 3210 4652 3222
rect 4590 3034 4606 3210
rect 4640 3034 4652 3210
rect 4590 3022 4652 3034
rect 4708 3210 4770 3222
rect 4708 3034 4720 3210
rect 4754 3034 4770 3210
rect 4708 3022 4770 3034
rect 4800 3210 4862 3222
rect 4800 3034 4816 3210
rect 4850 3034 4862 3210
rect 4800 3022 4862 3034
rect 4918 3210 4980 3222
rect 4918 3034 4930 3210
rect 4964 3034 4980 3210
rect 4918 3022 4980 3034
rect 5010 3210 5072 3222
rect 5010 3034 5026 3210
rect 5060 3034 5072 3210
rect 5010 3022 5072 3034
rect 5128 3210 5190 3222
rect 5128 3034 5140 3210
rect 5174 3034 5190 3210
rect 5128 3022 5190 3034
rect 5220 3210 5282 3222
rect 5220 3034 5236 3210
rect 5270 3034 5282 3210
rect 5220 3022 5282 3034
rect 5338 3210 5400 3222
rect 5338 3034 5350 3210
rect 5384 3034 5400 3210
rect 5338 3022 5400 3034
rect 5430 3210 5492 3222
rect 5430 3034 5446 3210
rect 5480 3034 5492 3210
rect 5430 3022 5492 3034
rect 5548 3210 5610 3222
rect 5548 3034 5560 3210
rect 5594 3034 5610 3210
rect 5548 3022 5610 3034
rect 5640 3210 5702 3222
rect 5640 3034 5656 3210
rect 5690 3034 5702 3210
rect 5640 3022 5702 3034
rect 5758 3210 5820 3222
rect 5758 3034 5770 3210
rect 5804 3034 5820 3210
rect 5758 3022 5820 3034
rect 5850 3210 5912 3222
rect 5850 3034 5866 3210
rect 5900 3034 5912 3210
rect 5850 3022 5912 3034
rect 5968 3210 6030 3222
rect 5968 3034 5980 3210
rect 6014 3034 6030 3210
rect 5968 3022 6030 3034
rect 6060 3210 6122 3222
rect 6060 3034 6076 3210
rect 6110 3034 6122 3210
rect 6060 3022 6122 3034
rect -2642 2770 -2580 2782
rect -2642 2594 -2630 2770
rect -2596 2594 -2580 2770
rect -2642 2582 -2580 2594
rect -2550 2770 -2488 2782
rect -2550 2594 -2534 2770
rect -2500 2594 -2488 2770
rect -2550 2582 -2488 2594
rect -2432 2770 -2370 2782
rect -2432 2594 -2420 2770
rect -2386 2594 -2370 2770
rect -2432 2582 -2370 2594
rect -2340 2770 -2278 2782
rect -2340 2594 -2324 2770
rect -2290 2594 -2278 2770
rect -2340 2582 -2278 2594
rect -2222 2770 -2160 2782
rect -2222 2594 -2210 2770
rect -2176 2594 -2160 2770
rect -2222 2582 -2160 2594
rect -2130 2770 -2068 2782
rect -2130 2594 -2114 2770
rect -2080 2594 -2068 2770
rect -2130 2582 -2068 2594
rect -2012 2770 -1950 2782
rect -2012 2594 -2000 2770
rect -1966 2594 -1950 2770
rect -2012 2582 -1950 2594
rect -1920 2770 -1858 2782
rect -1920 2594 -1904 2770
rect -1870 2594 -1858 2770
rect -1920 2582 -1858 2594
rect -1802 2770 -1740 2782
rect -1802 2594 -1790 2770
rect -1756 2594 -1740 2770
rect -1802 2582 -1740 2594
rect -1710 2770 -1648 2782
rect -1710 2594 -1694 2770
rect -1660 2594 -1648 2770
rect -1710 2582 -1648 2594
rect -1592 2770 -1530 2782
rect -1592 2594 -1580 2770
rect -1546 2594 -1530 2770
rect -1592 2582 -1530 2594
rect -1500 2770 -1438 2782
rect -1500 2594 -1484 2770
rect -1450 2594 -1438 2770
rect -1500 2582 -1438 2594
rect -1382 2770 -1320 2782
rect -1382 2594 -1370 2770
rect -1336 2594 -1320 2770
rect -1382 2582 -1320 2594
rect -1290 2770 -1228 2782
rect -1290 2594 -1274 2770
rect -1240 2594 -1228 2770
rect -1290 2582 -1228 2594
rect -1172 2770 -1110 2782
rect -1172 2594 -1160 2770
rect -1126 2594 -1110 2770
rect -1172 2582 -1110 2594
rect -1080 2770 -1018 2782
rect -1080 2594 -1064 2770
rect -1030 2594 -1018 2770
rect -1080 2582 -1018 2594
rect -962 2770 -900 2782
rect -962 2594 -950 2770
rect -916 2594 -900 2770
rect -962 2582 -900 2594
rect -870 2770 -808 2782
rect -870 2594 -854 2770
rect -820 2594 -808 2770
rect -870 2582 -808 2594
rect -752 2770 -690 2782
rect -752 2594 -740 2770
rect -706 2594 -690 2770
rect -752 2582 -690 2594
rect -660 2770 -598 2782
rect -660 2594 -644 2770
rect -610 2594 -598 2770
rect -660 2582 -598 2594
rect -542 2770 -480 2782
rect -542 2594 -530 2770
rect -496 2594 -480 2770
rect -542 2582 -480 2594
rect -450 2770 -388 2782
rect -450 2594 -434 2770
rect -400 2594 -388 2770
rect -450 2582 -388 2594
rect -332 2770 -270 2782
rect -332 2594 -320 2770
rect -286 2594 -270 2770
rect -332 2582 -270 2594
rect -240 2770 -178 2782
rect -240 2594 -224 2770
rect -190 2594 -178 2770
rect -240 2582 -178 2594
rect -122 2770 -60 2782
rect -122 2594 -110 2770
rect -76 2594 -60 2770
rect -122 2582 -60 2594
rect -30 2770 32 2782
rect -30 2594 -14 2770
rect 20 2594 32 2770
rect -30 2582 32 2594
rect 88 2770 150 2782
rect 88 2594 100 2770
rect 134 2594 150 2770
rect 88 2582 150 2594
rect 180 2770 242 2782
rect 180 2594 196 2770
rect 230 2594 242 2770
rect 180 2582 242 2594
rect 298 2770 360 2782
rect 298 2594 310 2770
rect 344 2594 360 2770
rect 298 2582 360 2594
rect 390 2770 452 2782
rect 390 2594 406 2770
rect 440 2594 452 2770
rect 390 2582 452 2594
rect 508 2770 570 2782
rect 508 2594 520 2770
rect 554 2594 570 2770
rect 508 2582 570 2594
rect 600 2770 662 2782
rect 600 2594 616 2770
rect 650 2594 662 2770
rect 600 2582 662 2594
rect 718 2770 780 2782
rect 718 2594 730 2770
rect 764 2594 780 2770
rect 718 2582 780 2594
rect 810 2770 872 2782
rect 810 2594 826 2770
rect 860 2594 872 2770
rect 810 2582 872 2594
rect 928 2770 990 2782
rect 928 2594 940 2770
rect 974 2594 990 2770
rect 928 2582 990 2594
rect 1020 2770 1082 2782
rect 1020 2594 1036 2770
rect 1070 2594 1082 2770
rect 1020 2582 1082 2594
rect 1138 2770 1200 2782
rect 1138 2594 1150 2770
rect 1184 2594 1200 2770
rect 1138 2582 1200 2594
rect 1230 2770 1292 2782
rect 1230 2594 1246 2770
rect 1280 2594 1292 2770
rect 1230 2582 1292 2594
rect 1348 2770 1410 2782
rect 1348 2594 1360 2770
rect 1394 2594 1410 2770
rect 1348 2582 1410 2594
rect 1440 2770 1502 2782
rect 1440 2594 1456 2770
rect 1490 2594 1502 2770
rect 1440 2582 1502 2594
rect 1558 2770 1620 2782
rect 1558 2594 1570 2770
rect 1604 2594 1620 2770
rect 1558 2582 1620 2594
rect 1650 2770 1712 2782
rect 1650 2594 1666 2770
rect 1700 2594 1712 2770
rect 1650 2582 1712 2594
rect 1768 2770 1830 2782
rect 1768 2594 1780 2770
rect 1814 2594 1830 2770
rect 1768 2582 1830 2594
rect 1860 2770 1922 2782
rect 1860 2594 1876 2770
rect 1910 2594 1922 2770
rect 1860 2582 1922 2594
rect 1978 2770 2040 2782
rect 1978 2594 1990 2770
rect 2024 2594 2040 2770
rect 1978 2582 2040 2594
rect 2070 2770 2132 2782
rect 2070 2594 2086 2770
rect 2120 2594 2132 2770
rect 2070 2582 2132 2594
rect 2188 2770 2250 2782
rect 2188 2594 2200 2770
rect 2234 2594 2250 2770
rect 2188 2582 2250 2594
rect 2280 2770 2342 2782
rect 2280 2594 2296 2770
rect 2330 2594 2342 2770
rect 2280 2582 2342 2594
rect 2398 2770 2460 2782
rect 2398 2594 2410 2770
rect 2444 2594 2460 2770
rect 2398 2582 2460 2594
rect 2490 2770 2552 2782
rect 2490 2594 2506 2770
rect 2540 2594 2552 2770
rect 2490 2582 2552 2594
rect 2608 2770 2670 2782
rect 2608 2594 2620 2770
rect 2654 2594 2670 2770
rect 2608 2582 2670 2594
rect 2700 2770 2762 2782
rect 2700 2594 2716 2770
rect 2750 2594 2762 2770
rect 2700 2582 2762 2594
rect 2818 2770 2880 2782
rect 2818 2594 2830 2770
rect 2864 2594 2880 2770
rect 2818 2582 2880 2594
rect 2910 2770 2972 2782
rect 2910 2594 2926 2770
rect 2960 2594 2972 2770
rect 2910 2582 2972 2594
rect 3028 2770 3090 2782
rect 3028 2594 3040 2770
rect 3074 2594 3090 2770
rect 3028 2582 3090 2594
rect 3120 2770 3182 2782
rect 3120 2594 3136 2770
rect 3170 2594 3182 2770
rect 3120 2582 3182 2594
rect 3238 2770 3300 2782
rect 3238 2594 3250 2770
rect 3284 2594 3300 2770
rect 3238 2582 3300 2594
rect 3330 2770 3392 2782
rect 3330 2594 3346 2770
rect 3380 2594 3392 2770
rect 3330 2582 3392 2594
rect 3448 2770 3510 2782
rect 3448 2594 3460 2770
rect 3494 2594 3510 2770
rect 3448 2582 3510 2594
rect 3540 2770 3602 2782
rect 3540 2594 3556 2770
rect 3590 2594 3602 2770
rect 3540 2582 3602 2594
rect 3658 2770 3720 2782
rect 3658 2594 3670 2770
rect 3704 2594 3720 2770
rect 3658 2582 3720 2594
rect 3750 2770 3812 2782
rect 3750 2594 3766 2770
rect 3800 2594 3812 2770
rect 3750 2582 3812 2594
rect 3868 2770 3930 2782
rect 3868 2594 3880 2770
rect 3914 2594 3930 2770
rect 3868 2582 3930 2594
rect 3960 2770 4022 2782
rect 3960 2594 3976 2770
rect 4010 2594 4022 2770
rect 3960 2582 4022 2594
rect 4078 2770 4140 2782
rect 4078 2594 4090 2770
rect 4124 2594 4140 2770
rect 4078 2582 4140 2594
rect 4170 2770 4232 2782
rect 4170 2594 4186 2770
rect 4220 2594 4232 2770
rect 4170 2582 4232 2594
rect 4288 2770 4350 2782
rect 4288 2594 4300 2770
rect 4334 2594 4350 2770
rect 4288 2582 4350 2594
rect 4380 2770 4442 2782
rect 4380 2594 4396 2770
rect 4430 2594 4442 2770
rect 4380 2582 4442 2594
rect 4498 2770 4560 2782
rect 4498 2594 4510 2770
rect 4544 2594 4560 2770
rect 4498 2582 4560 2594
rect 4590 2770 4652 2782
rect 4590 2594 4606 2770
rect 4640 2594 4652 2770
rect 4590 2582 4652 2594
rect 4708 2770 4770 2782
rect 4708 2594 4720 2770
rect 4754 2594 4770 2770
rect 4708 2582 4770 2594
rect 4800 2770 4862 2782
rect 4800 2594 4816 2770
rect 4850 2594 4862 2770
rect 4800 2582 4862 2594
rect 4918 2770 4980 2782
rect 4918 2594 4930 2770
rect 4964 2594 4980 2770
rect 4918 2582 4980 2594
rect 5010 2770 5072 2782
rect 5010 2594 5026 2770
rect 5060 2594 5072 2770
rect 5010 2582 5072 2594
rect 5128 2770 5190 2782
rect 5128 2594 5140 2770
rect 5174 2594 5190 2770
rect 5128 2582 5190 2594
rect 5220 2770 5282 2782
rect 5220 2594 5236 2770
rect 5270 2594 5282 2770
rect 5220 2582 5282 2594
rect 5338 2770 5400 2782
rect 5338 2594 5350 2770
rect 5384 2594 5400 2770
rect 5338 2582 5400 2594
rect 5430 2770 5492 2782
rect 5430 2594 5446 2770
rect 5480 2594 5492 2770
rect 5430 2582 5492 2594
rect 5548 2770 5610 2782
rect 5548 2594 5560 2770
rect 5594 2594 5610 2770
rect 5548 2582 5610 2594
rect 5640 2770 5702 2782
rect 5640 2594 5656 2770
rect 5690 2594 5702 2770
rect 5640 2582 5702 2594
rect 5758 2770 5820 2782
rect 5758 2594 5770 2770
rect 5804 2594 5820 2770
rect 5758 2582 5820 2594
rect 5850 2770 5912 2782
rect 5850 2594 5866 2770
rect 5900 2594 5912 2770
rect 5850 2582 5912 2594
rect 5968 2770 6030 2782
rect 5968 2594 5980 2770
rect 6014 2594 6030 2770
rect 5968 2582 6030 2594
rect 6060 2770 6122 2782
rect 6060 2594 6076 2770
rect 6110 2594 6122 2770
rect 6060 2582 6122 2594
rect -2642 2330 -2580 2342
rect -2642 2154 -2630 2330
rect -2596 2154 -2580 2330
rect -2642 2142 -2580 2154
rect -2550 2330 -2488 2342
rect -2550 2154 -2534 2330
rect -2500 2154 -2488 2330
rect -2550 2142 -2488 2154
rect -2432 2330 -2370 2342
rect -2432 2154 -2420 2330
rect -2386 2154 -2370 2330
rect -2432 2142 -2370 2154
rect -2340 2330 -2278 2342
rect -2340 2154 -2324 2330
rect -2290 2154 -2278 2330
rect -2340 2142 -2278 2154
rect -2222 2330 -2160 2342
rect -2222 2154 -2210 2330
rect -2176 2154 -2160 2330
rect -2222 2142 -2160 2154
rect -2130 2330 -2068 2342
rect -2130 2154 -2114 2330
rect -2080 2154 -2068 2330
rect -2130 2142 -2068 2154
rect -2012 2330 -1950 2342
rect -2012 2154 -2000 2330
rect -1966 2154 -1950 2330
rect -2012 2142 -1950 2154
rect -1920 2330 -1858 2342
rect -1920 2154 -1904 2330
rect -1870 2154 -1858 2330
rect -1920 2142 -1858 2154
rect -1802 2330 -1740 2342
rect -1802 2154 -1790 2330
rect -1756 2154 -1740 2330
rect -1802 2142 -1740 2154
rect -1710 2330 -1648 2342
rect -1710 2154 -1694 2330
rect -1660 2154 -1648 2330
rect -1710 2142 -1648 2154
rect -1592 2330 -1530 2342
rect -1592 2154 -1580 2330
rect -1546 2154 -1530 2330
rect -1592 2142 -1530 2154
rect -1500 2330 -1438 2342
rect -1500 2154 -1484 2330
rect -1450 2154 -1438 2330
rect -1500 2142 -1438 2154
rect -1382 2330 -1320 2342
rect -1382 2154 -1370 2330
rect -1336 2154 -1320 2330
rect -1382 2142 -1320 2154
rect -1290 2330 -1228 2342
rect -1290 2154 -1274 2330
rect -1240 2154 -1228 2330
rect -1290 2142 -1228 2154
rect -1172 2330 -1110 2342
rect -1172 2154 -1160 2330
rect -1126 2154 -1110 2330
rect -1172 2142 -1110 2154
rect -1080 2330 -1018 2342
rect -1080 2154 -1064 2330
rect -1030 2154 -1018 2330
rect -1080 2142 -1018 2154
rect -962 2330 -900 2342
rect -962 2154 -950 2330
rect -916 2154 -900 2330
rect -962 2142 -900 2154
rect -870 2330 -808 2342
rect -870 2154 -854 2330
rect -820 2154 -808 2330
rect -870 2142 -808 2154
rect -752 2330 -690 2342
rect -752 2154 -740 2330
rect -706 2154 -690 2330
rect -752 2142 -690 2154
rect -660 2330 -598 2342
rect -660 2154 -644 2330
rect -610 2154 -598 2330
rect -660 2142 -598 2154
rect -542 2330 -480 2342
rect -542 2154 -530 2330
rect -496 2154 -480 2330
rect -542 2142 -480 2154
rect -450 2330 -388 2342
rect -450 2154 -434 2330
rect -400 2154 -388 2330
rect -450 2142 -388 2154
rect -332 2330 -270 2342
rect -332 2154 -320 2330
rect -286 2154 -270 2330
rect -332 2142 -270 2154
rect -240 2330 -178 2342
rect -240 2154 -224 2330
rect -190 2154 -178 2330
rect -240 2142 -178 2154
rect -122 2330 -60 2342
rect -122 2154 -110 2330
rect -76 2154 -60 2330
rect -122 2142 -60 2154
rect -30 2330 32 2342
rect -30 2154 -14 2330
rect 20 2154 32 2330
rect -30 2142 32 2154
rect 88 2330 150 2342
rect 88 2154 100 2330
rect 134 2154 150 2330
rect 88 2142 150 2154
rect 180 2330 242 2342
rect 180 2154 196 2330
rect 230 2154 242 2330
rect 180 2142 242 2154
rect 298 2330 360 2342
rect 298 2154 310 2330
rect 344 2154 360 2330
rect 298 2142 360 2154
rect 390 2330 452 2342
rect 390 2154 406 2330
rect 440 2154 452 2330
rect 390 2142 452 2154
rect 508 2330 570 2342
rect 508 2154 520 2330
rect 554 2154 570 2330
rect 508 2142 570 2154
rect 600 2330 662 2342
rect 600 2154 616 2330
rect 650 2154 662 2330
rect 600 2142 662 2154
rect 718 2330 780 2342
rect 718 2154 730 2330
rect 764 2154 780 2330
rect 718 2142 780 2154
rect 810 2330 872 2342
rect 810 2154 826 2330
rect 860 2154 872 2330
rect 810 2142 872 2154
rect 928 2330 990 2342
rect 928 2154 940 2330
rect 974 2154 990 2330
rect 928 2142 990 2154
rect 1020 2330 1082 2342
rect 1020 2154 1036 2330
rect 1070 2154 1082 2330
rect 1020 2142 1082 2154
rect 1138 2330 1200 2342
rect 1138 2154 1150 2330
rect 1184 2154 1200 2330
rect 1138 2142 1200 2154
rect 1230 2330 1292 2342
rect 1230 2154 1246 2330
rect 1280 2154 1292 2330
rect 1230 2142 1292 2154
rect 1348 2330 1410 2342
rect 1348 2154 1360 2330
rect 1394 2154 1410 2330
rect 1348 2142 1410 2154
rect 1440 2330 1502 2342
rect 1440 2154 1456 2330
rect 1490 2154 1502 2330
rect 1440 2142 1502 2154
rect 1558 2330 1620 2342
rect 1558 2154 1570 2330
rect 1604 2154 1620 2330
rect 1558 2142 1620 2154
rect 1650 2330 1712 2342
rect 1650 2154 1666 2330
rect 1700 2154 1712 2330
rect 1650 2142 1712 2154
rect 1768 2330 1830 2342
rect 1768 2154 1780 2330
rect 1814 2154 1830 2330
rect 1768 2142 1830 2154
rect 1860 2330 1922 2342
rect 1860 2154 1876 2330
rect 1910 2154 1922 2330
rect 1860 2142 1922 2154
rect 1978 2330 2040 2342
rect 1978 2154 1990 2330
rect 2024 2154 2040 2330
rect 1978 2142 2040 2154
rect 2070 2330 2132 2342
rect 2070 2154 2086 2330
rect 2120 2154 2132 2330
rect 2070 2142 2132 2154
rect 2188 2330 2250 2342
rect 2188 2154 2200 2330
rect 2234 2154 2250 2330
rect 2188 2142 2250 2154
rect 2280 2330 2342 2342
rect 2280 2154 2296 2330
rect 2330 2154 2342 2330
rect 2280 2142 2342 2154
rect 2398 2330 2460 2342
rect 2398 2154 2410 2330
rect 2444 2154 2460 2330
rect 2398 2142 2460 2154
rect 2490 2330 2552 2342
rect 2490 2154 2506 2330
rect 2540 2154 2552 2330
rect 2490 2142 2552 2154
rect 2608 2330 2670 2342
rect 2608 2154 2620 2330
rect 2654 2154 2670 2330
rect 2608 2142 2670 2154
rect 2700 2330 2762 2342
rect 2700 2154 2716 2330
rect 2750 2154 2762 2330
rect 2700 2142 2762 2154
rect 2818 2330 2880 2342
rect 2818 2154 2830 2330
rect 2864 2154 2880 2330
rect 2818 2142 2880 2154
rect 2910 2330 2972 2342
rect 2910 2154 2926 2330
rect 2960 2154 2972 2330
rect 2910 2142 2972 2154
rect 3028 2330 3090 2342
rect 3028 2154 3040 2330
rect 3074 2154 3090 2330
rect 3028 2142 3090 2154
rect 3120 2330 3182 2342
rect 3120 2154 3136 2330
rect 3170 2154 3182 2330
rect 3120 2142 3182 2154
rect 3238 2330 3300 2342
rect 3238 2154 3250 2330
rect 3284 2154 3300 2330
rect 3238 2142 3300 2154
rect 3330 2330 3392 2342
rect 3330 2154 3346 2330
rect 3380 2154 3392 2330
rect 3330 2142 3392 2154
rect 3448 2330 3510 2342
rect 3448 2154 3460 2330
rect 3494 2154 3510 2330
rect 3448 2142 3510 2154
rect 3540 2330 3602 2342
rect 3540 2154 3556 2330
rect 3590 2154 3602 2330
rect 3540 2142 3602 2154
rect 3658 2330 3720 2342
rect 3658 2154 3670 2330
rect 3704 2154 3720 2330
rect 3658 2142 3720 2154
rect 3750 2330 3812 2342
rect 3750 2154 3766 2330
rect 3800 2154 3812 2330
rect 3750 2142 3812 2154
rect 3868 2330 3930 2342
rect 3868 2154 3880 2330
rect 3914 2154 3930 2330
rect 3868 2142 3930 2154
rect 3960 2330 4022 2342
rect 3960 2154 3976 2330
rect 4010 2154 4022 2330
rect 3960 2142 4022 2154
rect 4078 2330 4140 2342
rect 4078 2154 4090 2330
rect 4124 2154 4140 2330
rect 4078 2142 4140 2154
rect 4170 2330 4232 2342
rect 4170 2154 4186 2330
rect 4220 2154 4232 2330
rect 4170 2142 4232 2154
rect 4288 2330 4350 2342
rect 4288 2154 4300 2330
rect 4334 2154 4350 2330
rect 4288 2142 4350 2154
rect 4380 2330 4442 2342
rect 4380 2154 4396 2330
rect 4430 2154 4442 2330
rect 4380 2142 4442 2154
rect 4498 2330 4560 2342
rect 4498 2154 4510 2330
rect 4544 2154 4560 2330
rect 4498 2142 4560 2154
rect 4590 2330 4652 2342
rect 4590 2154 4606 2330
rect 4640 2154 4652 2330
rect 4590 2142 4652 2154
rect 4708 2330 4770 2342
rect 4708 2154 4720 2330
rect 4754 2154 4770 2330
rect 4708 2142 4770 2154
rect 4800 2330 4862 2342
rect 4800 2154 4816 2330
rect 4850 2154 4862 2330
rect 4800 2142 4862 2154
rect 4918 2330 4980 2342
rect 4918 2154 4930 2330
rect 4964 2154 4980 2330
rect 4918 2142 4980 2154
rect 5010 2330 5072 2342
rect 5010 2154 5026 2330
rect 5060 2154 5072 2330
rect 5010 2142 5072 2154
rect 5128 2330 5190 2342
rect 5128 2154 5140 2330
rect 5174 2154 5190 2330
rect 5128 2142 5190 2154
rect 5220 2330 5282 2342
rect 5220 2154 5236 2330
rect 5270 2154 5282 2330
rect 5220 2142 5282 2154
rect 5338 2330 5400 2342
rect 5338 2154 5350 2330
rect 5384 2154 5400 2330
rect 5338 2142 5400 2154
rect 5430 2330 5492 2342
rect 5430 2154 5446 2330
rect 5480 2154 5492 2330
rect 5430 2142 5492 2154
rect 5548 2330 5610 2342
rect 5548 2154 5560 2330
rect 5594 2154 5610 2330
rect 5548 2142 5610 2154
rect 5640 2330 5702 2342
rect 5640 2154 5656 2330
rect 5690 2154 5702 2330
rect 5640 2142 5702 2154
rect 5758 2330 5820 2342
rect 5758 2154 5770 2330
rect 5804 2154 5820 2330
rect 5758 2142 5820 2154
rect 5850 2330 5912 2342
rect 5850 2154 5866 2330
rect 5900 2154 5912 2330
rect 5850 2142 5912 2154
rect 5968 2330 6030 2342
rect 5968 2154 5980 2330
rect 6014 2154 6030 2330
rect 5968 2142 6030 2154
rect 6060 2330 6122 2342
rect 6060 2154 6076 2330
rect 6110 2154 6122 2330
rect 6060 2142 6122 2154
rect -2642 1890 -2580 1902
rect -2642 1714 -2630 1890
rect -2596 1714 -2580 1890
rect -2642 1702 -2580 1714
rect -2550 1890 -2488 1902
rect -2550 1714 -2534 1890
rect -2500 1714 -2488 1890
rect -2550 1702 -2488 1714
rect -2432 1890 -2370 1902
rect -2432 1714 -2420 1890
rect -2386 1714 -2370 1890
rect -2432 1702 -2370 1714
rect -2340 1890 -2278 1902
rect -2340 1714 -2324 1890
rect -2290 1714 -2278 1890
rect -2340 1702 -2278 1714
rect -2222 1890 -2160 1902
rect -2222 1714 -2210 1890
rect -2176 1714 -2160 1890
rect -2222 1702 -2160 1714
rect -2130 1890 -2068 1902
rect -2130 1714 -2114 1890
rect -2080 1714 -2068 1890
rect -2130 1702 -2068 1714
rect -2012 1890 -1950 1902
rect -2012 1714 -2000 1890
rect -1966 1714 -1950 1890
rect -2012 1702 -1950 1714
rect -1920 1890 -1858 1902
rect -1920 1714 -1904 1890
rect -1870 1714 -1858 1890
rect -1920 1702 -1858 1714
rect -1802 1890 -1740 1902
rect -1802 1714 -1790 1890
rect -1756 1714 -1740 1890
rect -1802 1702 -1740 1714
rect -1710 1890 -1648 1902
rect -1710 1714 -1694 1890
rect -1660 1714 -1648 1890
rect -1710 1702 -1648 1714
rect -1592 1890 -1530 1902
rect -1592 1714 -1580 1890
rect -1546 1714 -1530 1890
rect -1592 1702 -1530 1714
rect -1500 1890 -1438 1902
rect -1500 1714 -1484 1890
rect -1450 1714 -1438 1890
rect -1500 1702 -1438 1714
rect -1382 1890 -1320 1902
rect -1382 1714 -1370 1890
rect -1336 1714 -1320 1890
rect -1382 1702 -1320 1714
rect -1290 1890 -1228 1902
rect -1290 1714 -1274 1890
rect -1240 1714 -1228 1890
rect -1290 1702 -1228 1714
rect -1172 1890 -1110 1902
rect -1172 1714 -1160 1890
rect -1126 1714 -1110 1890
rect -1172 1702 -1110 1714
rect -1080 1890 -1018 1902
rect -1080 1714 -1064 1890
rect -1030 1714 -1018 1890
rect -1080 1702 -1018 1714
rect -962 1890 -900 1902
rect -962 1714 -950 1890
rect -916 1714 -900 1890
rect -962 1702 -900 1714
rect -870 1890 -808 1902
rect -870 1714 -854 1890
rect -820 1714 -808 1890
rect -870 1702 -808 1714
rect -752 1890 -690 1902
rect -752 1714 -740 1890
rect -706 1714 -690 1890
rect -752 1702 -690 1714
rect -660 1890 -598 1902
rect -660 1714 -644 1890
rect -610 1714 -598 1890
rect -660 1702 -598 1714
rect -542 1890 -480 1902
rect -542 1714 -530 1890
rect -496 1714 -480 1890
rect -542 1702 -480 1714
rect -450 1890 -388 1902
rect -450 1714 -434 1890
rect -400 1714 -388 1890
rect -450 1702 -388 1714
rect -332 1890 -270 1902
rect -332 1714 -320 1890
rect -286 1714 -270 1890
rect -332 1702 -270 1714
rect -240 1890 -178 1902
rect -240 1714 -224 1890
rect -190 1714 -178 1890
rect -240 1702 -178 1714
rect -122 1890 -60 1902
rect -122 1714 -110 1890
rect -76 1714 -60 1890
rect -122 1702 -60 1714
rect -30 1890 32 1902
rect -30 1714 -14 1890
rect 20 1714 32 1890
rect -30 1702 32 1714
rect 88 1890 150 1902
rect 88 1714 100 1890
rect 134 1714 150 1890
rect 88 1702 150 1714
rect 180 1890 242 1902
rect 180 1714 196 1890
rect 230 1714 242 1890
rect 180 1702 242 1714
rect 298 1890 360 1902
rect 298 1714 310 1890
rect 344 1714 360 1890
rect 298 1702 360 1714
rect 390 1890 452 1902
rect 390 1714 406 1890
rect 440 1714 452 1890
rect 390 1702 452 1714
rect 508 1890 570 1902
rect 508 1714 520 1890
rect 554 1714 570 1890
rect 508 1702 570 1714
rect 600 1890 662 1902
rect 600 1714 616 1890
rect 650 1714 662 1890
rect 600 1702 662 1714
rect 718 1890 780 1902
rect 718 1714 730 1890
rect 764 1714 780 1890
rect 718 1702 780 1714
rect 810 1890 872 1902
rect 810 1714 826 1890
rect 860 1714 872 1890
rect 810 1702 872 1714
rect 928 1890 990 1902
rect 928 1714 940 1890
rect 974 1714 990 1890
rect 928 1702 990 1714
rect 1020 1890 1082 1902
rect 1020 1714 1036 1890
rect 1070 1714 1082 1890
rect 1020 1702 1082 1714
rect 1138 1890 1200 1902
rect 1138 1714 1150 1890
rect 1184 1714 1200 1890
rect 1138 1702 1200 1714
rect 1230 1890 1292 1902
rect 1230 1714 1246 1890
rect 1280 1714 1292 1890
rect 1230 1702 1292 1714
rect 1348 1890 1410 1902
rect 1348 1714 1360 1890
rect 1394 1714 1410 1890
rect 1348 1702 1410 1714
rect 1440 1890 1502 1902
rect 1440 1714 1456 1890
rect 1490 1714 1502 1890
rect 1440 1702 1502 1714
rect 1558 1890 1620 1902
rect 1558 1714 1570 1890
rect 1604 1714 1620 1890
rect 1558 1702 1620 1714
rect 1650 1890 1712 1902
rect 1650 1714 1666 1890
rect 1700 1714 1712 1890
rect 1650 1702 1712 1714
rect 1768 1890 1830 1902
rect 1768 1714 1780 1890
rect 1814 1714 1830 1890
rect 1768 1702 1830 1714
rect 1860 1890 1922 1902
rect 1860 1714 1876 1890
rect 1910 1714 1922 1890
rect 1860 1702 1922 1714
rect 1978 1890 2040 1902
rect 1978 1714 1990 1890
rect 2024 1714 2040 1890
rect 1978 1702 2040 1714
rect 2070 1890 2132 1902
rect 2070 1714 2086 1890
rect 2120 1714 2132 1890
rect 2070 1702 2132 1714
rect 2188 1890 2250 1902
rect 2188 1714 2200 1890
rect 2234 1714 2250 1890
rect 2188 1702 2250 1714
rect 2280 1890 2342 1902
rect 2280 1714 2296 1890
rect 2330 1714 2342 1890
rect 2280 1702 2342 1714
rect 2398 1890 2460 1902
rect 2398 1714 2410 1890
rect 2444 1714 2460 1890
rect 2398 1702 2460 1714
rect 2490 1890 2552 1902
rect 2490 1714 2506 1890
rect 2540 1714 2552 1890
rect 2490 1702 2552 1714
rect 2608 1890 2670 1902
rect 2608 1714 2620 1890
rect 2654 1714 2670 1890
rect 2608 1702 2670 1714
rect 2700 1890 2762 1902
rect 2700 1714 2716 1890
rect 2750 1714 2762 1890
rect 2700 1702 2762 1714
rect 2818 1890 2880 1902
rect 2818 1714 2830 1890
rect 2864 1714 2880 1890
rect 2818 1702 2880 1714
rect 2910 1890 2972 1902
rect 2910 1714 2926 1890
rect 2960 1714 2972 1890
rect 2910 1702 2972 1714
rect 3028 1890 3090 1902
rect 3028 1714 3040 1890
rect 3074 1714 3090 1890
rect 3028 1702 3090 1714
rect 3120 1890 3182 1902
rect 3120 1714 3136 1890
rect 3170 1714 3182 1890
rect 3120 1702 3182 1714
rect 3238 1890 3300 1902
rect 3238 1714 3250 1890
rect 3284 1714 3300 1890
rect 3238 1702 3300 1714
rect 3330 1890 3392 1902
rect 3330 1714 3346 1890
rect 3380 1714 3392 1890
rect 3330 1702 3392 1714
rect 3448 1890 3510 1902
rect 3448 1714 3460 1890
rect 3494 1714 3510 1890
rect 3448 1702 3510 1714
rect 3540 1890 3602 1902
rect 3540 1714 3556 1890
rect 3590 1714 3602 1890
rect 3540 1702 3602 1714
rect 3658 1890 3720 1902
rect 3658 1714 3670 1890
rect 3704 1714 3720 1890
rect 3658 1702 3720 1714
rect 3750 1890 3812 1902
rect 3750 1714 3766 1890
rect 3800 1714 3812 1890
rect 3750 1702 3812 1714
rect 3868 1890 3930 1902
rect 3868 1714 3880 1890
rect 3914 1714 3930 1890
rect 3868 1702 3930 1714
rect 3960 1890 4022 1902
rect 3960 1714 3976 1890
rect 4010 1714 4022 1890
rect 3960 1702 4022 1714
rect 4078 1890 4140 1902
rect 4078 1714 4090 1890
rect 4124 1714 4140 1890
rect 4078 1702 4140 1714
rect 4170 1890 4232 1902
rect 4170 1714 4186 1890
rect 4220 1714 4232 1890
rect 4170 1702 4232 1714
rect 4288 1890 4350 1902
rect 4288 1714 4300 1890
rect 4334 1714 4350 1890
rect 4288 1702 4350 1714
rect 4380 1890 4442 1902
rect 4380 1714 4396 1890
rect 4430 1714 4442 1890
rect 4380 1702 4442 1714
rect 4498 1890 4560 1902
rect 4498 1714 4510 1890
rect 4544 1714 4560 1890
rect 4498 1702 4560 1714
rect 4590 1890 4652 1902
rect 4590 1714 4606 1890
rect 4640 1714 4652 1890
rect 4590 1702 4652 1714
rect 4708 1890 4770 1902
rect 4708 1714 4720 1890
rect 4754 1714 4770 1890
rect 4708 1702 4770 1714
rect 4800 1890 4862 1902
rect 4800 1714 4816 1890
rect 4850 1714 4862 1890
rect 4800 1702 4862 1714
rect 4918 1890 4980 1902
rect 4918 1714 4930 1890
rect 4964 1714 4980 1890
rect 4918 1702 4980 1714
rect 5010 1890 5072 1902
rect 5010 1714 5026 1890
rect 5060 1714 5072 1890
rect 5010 1702 5072 1714
rect 5128 1890 5190 1902
rect 5128 1714 5140 1890
rect 5174 1714 5190 1890
rect 5128 1702 5190 1714
rect 5220 1890 5282 1902
rect 5220 1714 5236 1890
rect 5270 1714 5282 1890
rect 5220 1702 5282 1714
rect 5338 1890 5400 1902
rect 5338 1714 5350 1890
rect 5384 1714 5400 1890
rect 5338 1702 5400 1714
rect 5430 1890 5492 1902
rect 5430 1714 5446 1890
rect 5480 1714 5492 1890
rect 5430 1702 5492 1714
rect 5548 1890 5610 1902
rect 5548 1714 5560 1890
rect 5594 1714 5610 1890
rect 5548 1702 5610 1714
rect 5640 1890 5702 1902
rect 5640 1714 5656 1890
rect 5690 1714 5702 1890
rect 5640 1702 5702 1714
rect 5758 1890 5820 1902
rect 5758 1714 5770 1890
rect 5804 1714 5820 1890
rect 5758 1702 5820 1714
rect 5850 1890 5912 1902
rect 5850 1714 5866 1890
rect 5900 1714 5912 1890
rect 5850 1702 5912 1714
rect 5968 1890 6030 1902
rect 5968 1714 5980 1890
rect 6014 1714 6030 1890
rect 5968 1702 6030 1714
rect 6060 1890 6122 1902
rect 6060 1714 6076 1890
rect 6110 1714 6122 1890
rect 6060 1702 6122 1714
rect -2642 1450 -2580 1462
rect -2642 1274 -2630 1450
rect -2596 1274 -2580 1450
rect -2642 1262 -2580 1274
rect -2550 1450 -2488 1462
rect -2550 1274 -2534 1450
rect -2500 1274 -2488 1450
rect -2550 1262 -2488 1274
rect -2432 1450 -2370 1462
rect -2432 1274 -2420 1450
rect -2386 1274 -2370 1450
rect -2432 1262 -2370 1274
rect -2340 1450 -2278 1462
rect -2340 1274 -2324 1450
rect -2290 1274 -2278 1450
rect -2340 1262 -2278 1274
rect -2222 1450 -2160 1462
rect -2222 1274 -2210 1450
rect -2176 1274 -2160 1450
rect -2222 1262 -2160 1274
rect -2130 1450 -2068 1462
rect -2130 1274 -2114 1450
rect -2080 1274 -2068 1450
rect -2130 1262 -2068 1274
rect -2012 1450 -1950 1462
rect -2012 1274 -2000 1450
rect -1966 1274 -1950 1450
rect -2012 1262 -1950 1274
rect -1920 1450 -1858 1462
rect -1920 1274 -1904 1450
rect -1870 1274 -1858 1450
rect -1920 1262 -1858 1274
rect -1802 1450 -1740 1462
rect -1802 1274 -1790 1450
rect -1756 1274 -1740 1450
rect -1802 1262 -1740 1274
rect -1710 1450 -1648 1462
rect -1710 1274 -1694 1450
rect -1660 1274 -1648 1450
rect -1710 1262 -1648 1274
rect -1592 1450 -1530 1462
rect -1592 1274 -1580 1450
rect -1546 1274 -1530 1450
rect -1592 1262 -1530 1274
rect -1500 1450 -1438 1462
rect -1500 1274 -1484 1450
rect -1450 1274 -1438 1450
rect -1500 1262 -1438 1274
rect -1382 1450 -1320 1462
rect -1382 1274 -1370 1450
rect -1336 1274 -1320 1450
rect -1382 1262 -1320 1274
rect -1290 1450 -1228 1462
rect -1290 1274 -1274 1450
rect -1240 1274 -1228 1450
rect -1290 1262 -1228 1274
rect -1172 1450 -1110 1462
rect -1172 1274 -1160 1450
rect -1126 1274 -1110 1450
rect -1172 1262 -1110 1274
rect -1080 1450 -1018 1462
rect -1080 1274 -1064 1450
rect -1030 1274 -1018 1450
rect -1080 1262 -1018 1274
rect -962 1450 -900 1462
rect -962 1274 -950 1450
rect -916 1274 -900 1450
rect -962 1262 -900 1274
rect -870 1450 -808 1462
rect -870 1274 -854 1450
rect -820 1274 -808 1450
rect -870 1262 -808 1274
rect -752 1450 -690 1462
rect -752 1274 -740 1450
rect -706 1274 -690 1450
rect -752 1262 -690 1274
rect -660 1450 -598 1462
rect -660 1274 -644 1450
rect -610 1274 -598 1450
rect -660 1262 -598 1274
rect -542 1450 -480 1462
rect -542 1274 -530 1450
rect -496 1274 -480 1450
rect -542 1262 -480 1274
rect -450 1450 -388 1462
rect -450 1274 -434 1450
rect -400 1274 -388 1450
rect -450 1262 -388 1274
rect -332 1450 -270 1462
rect -332 1274 -320 1450
rect -286 1274 -270 1450
rect -332 1262 -270 1274
rect -240 1450 -178 1462
rect -240 1274 -224 1450
rect -190 1274 -178 1450
rect -240 1262 -178 1274
rect -122 1450 -60 1462
rect -122 1274 -110 1450
rect -76 1274 -60 1450
rect -122 1262 -60 1274
rect -30 1450 32 1462
rect -30 1274 -14 1450
rect 20 1274 32 1450
rect -30 1262 32 1274
rect 88 1450 150 1462
rect 88 1274 100 1450
rect 134 1274 150 1450
rect 88 1262 150 1274
rect 180 1450 242 1462
rect 180 1274 196 1450
rect 230 1274 242 1450
rect 180 1262 242 1274
rect 298 1450 360 1462
rect 298 1274 310 1450
rect 344 1274 360 1450
rect 298 1262 360 1274
rect 390 1450 452 1462
rect 390 1274 406 1450
rect 440 1274 452 1450
rect 390 1262 452 1274
rect 508 1450 570 1462
rect 508 1274 520 1450
rect 554 1274 570 1450
rect 508 1262 570 1274
rect 600 1450 662 1462
rect 600 1274 616 1450
rect 650 1274 662 1450
rect 600 1262 662 1274
rect 718 1450 780 1462
rect 718 1274 730 1450
rect 764 1274 780 1450
rect 718 1262 780 1274
rect 810 1450 872 1462
rect 810 1274 826 1450
rect 860 1274 872 1450
rect 810 1262 872 1274
rect 928 1450 990 1462
rect 928 1274 940 1450
rect 974 1274 990 1450
rect 928 1262 990 1274
rect 1020 1450 1082 1462
rect 1020 1274 1036 1450
rect 1070 1274 1082 1450
rect 1020 1262 1082 1274
rect 1138 1450 1200 1462
rect 1138 1274 1150 1450
rect 1184 1274 1200 1450
rect 1138 1262 1200 1274
rect 1230 1450 1292 1462
rect 1230 1274 1246 1450
rect 1280 1274 1292 1450
rect 1230 1262 1292 1274
rect 1348 1450 1410 1462
rect 1348 1274 1360 1450
rect 1394 1274 1410 1450
rect 1348 1262 1410 1274
rect 1440 1450 1502 1462
rect 1440 1274 1456 1450
rect 1490 1274 1502 1450
rect 1440 1262 1502 1274
rect 1558 1450 1620 1462
rect 1558 1274 1570 1450
rect 1604 1274 1620 1450
rect 1558 1262 1620 1274
rect 1650 1450 1712 1462
rect 1650 1274 1666 1450
rect 1700 1274 1712 1450
rect 1650 1262 1712 1274
rect 1768 1450 1830 1462
rect 1768 1274 1780 1450
rect 1814 1274 1830 1450
rect 1768 1262 1830 1274
rect 1860 1450 1922 1462
rect 1860 1274 1876 1450
rect 1910 1274 1922 1450
rect 1860 1262 1922 1274
rect 1978 1450 2040 1462
rect 1978 1274 1990 1450
rect 2024 1274 2040 1450
rect 1978 1262 2040 1274
rect 2070 1450 2132 1462
rect 2070 1274 2086 1450
rect 2120 1274 2132 1450
rect 2070 1262 2132 1274
rect 2188 1450 2250 1462
rect 2188 1274 2200 1450
rect 2234 1274 2250 1450
rect 2188 1262 2250 1274
rect 2280 1450 2342 1462
rect 2280 1274 2296 1450
rect 2330 1274 2342 1450
rect 2280 1262 2342 1274
rect 2398 1450 2460 1462
rect 2398 1274 2410 1450
rect 2444 1274 2460 1450
rect 2398 1262 2460 1274
rect 2490 1450 2552 1462
rect 2490 1274 2506 1450
rect 2540 1274 2552 1450
rect 2490 1262 2552 1274
rect 2608 1450 2670 1462
rect 2608 1274 2620 1450
rect 2654 1274 2670 1450
rect 2608 1262 2670 1274
rect 2700 1450 2762 1462
rect 2700 1274 2716 1450
rect 2750 1274 2762 1450
rect 2700 1262 2762 1274
rect 2818 1450 2880 1462
rect 2818 1274 2830 1450
rect 2864 1274 2880 1450
rect 2818 1262 2880 1274
rect 2910 1450 2972 1462
rect 2910 1274 2926 1450
rect 2960 1274 2972 1450
rect 2910 1262 2972 1274
rect 3028 1450 3090 1462
rect 3028 1274 3040 1450
rect 3074 1274 3090 1450
rect 3028 1262 3090 1274
rect 3120 1450 3182 1462
rect 3120 1274 3136 1450
rect 3170 1274 3182 1450
rect 3120 1262 3182 1274
rect 3238 1450 3300 1462
rect 3238 1274 3250 1450
rect 3284 1274 3300 1450
rect 3238 1262 3300 1274
rect 3330 1450 3392 1462
rect 3330 1274 3346 1450
rect 3380 1274 3392 1450
rect 3330 1262 3392 1274
rect 3448 1450 3510 1462
rect 3448 1274 3460 1450
rect 3494 1274 3510 1450
rect 3448 1262 3510 1274
rect 3540 1450 3602 1462
rect 3540 1274 3556 1450
rect 3590 1274 3602 1450
rect 3540 1262 3602 1274
rect 3658 1450 3720 1462
rect 3658 1274 3670 1450
rect 3704 1274 3720 1450
rect 3658 1262 3720 1274
rect 3750 1450 3812 1462
rect 3750 1274 3766 1450
rect 3800 1274 3812 1450
rect 3750 1262 3812 1274
rect 3868 1450 3930 1462
rect 3868 1274 3880 1450
rect 3914 1274 3930 1450
rect 3868 1262 3930 1274
rect 3960 1450 4022 1462
rect 3960 1274 3976 1450
rect 4010 1274 4022 1450
rect 3960 1262 4022 1274
rect 4078 1450 4140 1462
rect 4078 1274 4090 1450
rect 4124 1274 4140 1450
rect 4078 1262 4140 1274
rect 4170 1450 4232 1462
rect 4170 1274 4186 1450
rect 4220 1274 4232 1450
rect 4170 1262 4232 1274
rect 4288 1450 4350 1462
rect 4288 1274 4300 1450
rect 4334 1274 4350 1450
rect 4288 1262 4350 1274
rect 4380 1450 4442 1462
rect 4380 1274 4396 1450
rect 4430 1274 4442 1450
rect 4380 1262 4442 1274
rect 4498 1450 4560 1462
rect 4498 1274 4510 1450
rect 4544 1274 4560 1450
rect 4498 1262 4560 1274
rect 4590 1450 4652 1462
rect 4590 1274 4606 1450
rect 4640 1274 4652 1450
rect 4590 1262 4652 1274
rect 4708 1450 4770 1462
rect 4708 1274 4720 1450
rect 4754 1274 4770 1450
rect 4708 1262 4770 1274
rect 4800 1450 4862 1462
rect 4800 1274 4816 1450
rect 4850 1274 4862 1450
rect 4800 1262 4862 1274
rect 4918 1450 4980 1462
rect 4918 1274 4930 1450
rect 4964 1274 4980 1450
rect 4918 1262 4980 1274
rect 5010 1450 5072 1462
rect 5010 1274 5026 1450
rect 5060 1274 5072 1450
rect 5010 1262 5072 1274
rect 5128 1450 5190 1462
rect 5128 1274 5140 1450
rect 5174 1274 5190 1450
rect 5128 1262 5190 1274
rect 5220 1450 5282 1462
rect 5220 1274 5236 1450
rect 5270 1274 5282 1450
rect 5220 1262 5282 1274
rect 5338 1450 5400 1462
rect 5338 1274 5350 1450
rect 5384 1274 5400 1450
rect 5338 1262 5400 1274
rect 5430 1450 5492 1462
rect 5430 1274 5446 1450
rect 5480 1274 5492 1450
rect 5430 1262 5492 1274
rect 5548 1450 5610 1462
rect 5548 1274 5560 1450
rect 5594 1274 5610 1450
rect 5548 1262 5610 1274
rect 5640 1450 5702 1462
rect 5640 1274 5656 1450
rect 5690 1274 5702 1450
rect 5640 1262 5702 1274
rect 5758 1450 5820 1462
rect 5758 1274 5770 1450
rect 5804 1274 5820 1450
rect 5758 1262 5820 1274
rect 5850 1450 5912 1462
rect 5850 1274 5866 1450
rect 5900 1274 5912 1450
rect 5850 1262 5912 1274
rect 5968 1450 6030 1462
rect 5968 1274 5980 1450
rect 6014 1274 6030 1450
rect 5968 1262 6030 1274
rect 6060 1450 6122 1462
rect 6060 1274 6076 1450
rect 6110 1274 6122 1450
rect 6060 1262 6122 1274
rect -2642 1010 -2580 1022
rect -2642 834 -2630 1010
rect -2596 834 -2580 1010
rect -2642 822 -2580 834
rect -2550 1010 -2488 1022
rect -2550 834 -2534 1010
rect -2500 834 -2488 1010
rect -2550 822 -2488 834
rect -2432 1010 -2370 1022
rect -2432 834 -2420 1010
rect -2386 834 -2370 1010
rect -2432 822 -2370 834
rect -2340 1010 -2278 1022
rect -2340 834 -2324 1010
rect -2290 834 -2278 1010
rect -2340 822 -2278 834
rect -2222 1010 -2160 1022
rect -2222 834 -2210 1010
rect -2176 834 -2160 1010
rect -2222 822 -2160 834
rect -2130 1010 -2068 1022
rect -2130 834 -2114 1010
rect -2080 834 -2068 1010
rect -2130 822 -2068 834
rect -2012 1010 -1950 1022
rect -2012 834 -2000 1010
rect -1966 834 -1950 1010
rect -2012 822 -1950 834
rect -1920 1010 -1858 1022
rect -1920 834 -1904 1010
rect -1870 834 -1858 1010
rect -1920 822 -1858 834
rect -1802 1010 -1740 1022
rect -1802 834 -1790 1010
rect -1756 834 -1740 1010
rect -1802 822 -1740 834
rect -1710 1010 -1648 1022
rect -1710 834 -1694 1010
rect -1660 834 -1648 1010
rect -1710 822 -1648 834
rect -1592 1010 -1530 1022
rect -1592 834 -1580 1010
rect -1546 834 -1530 1010
rect -1592 822 -1530 834
rect -1500 1010 -1438 1022
rect -1500 834 -1484 1010
rect -1450 834 -1438 1010
rect -1500 822 -1438 834
rect -1382 1010 -1320 1022
rect -1382 834 -1370 1010
rect -1336 834 -1320 1010
rect -1382 822 -1320 834
rect -1290 1010 -1228 1022
rect -1290 834 -1274 1010
rect -1240 834 -1228 1010
rect -1290 822 -1228 834
rect -1172 1010 -1110 1022
rect -1172 834 -1160 1010
rect -1126 834 -1110 1010
rect -1172 822 -1110 834
rect -1080 1010 -1018 1022
rect -1080 834 -1064 1010
rect -1030 834 -1018 1010
rect -1080 822 -1018 834
rect -962 1010 -900 1022
rect -962 834 -950 1010
rect -916 834 -900 1010
rect -962 822 -900 834
rect -870 1010 -808 1022
rect -870 834 -854 1010
rect -820 834 -808 1010
rect -870 822 -808 834
rect -752 1010 -690 1022
rect -752 834 -740 1010
rect -706 834 -690 1010
rect -752 822 -690 834
rect -660 1010 -598 1022
rect -660 834 -644 1010
rect -610 834 -598 1010
rect -660 822 -598 834
rect -542 1010 -480 1022
rect -542 834 -530 1010
rect -496 834 -480 1010
rect -542 822 -480 834
rect -450 1010 -388 1022
rect -450 834 -434 1010
rect -400 834 -388 1010
rect -450 822 -388 834
rect -332 1010 -270 1022
rect -332 834 -320 1010
rect -286 834 -270 1010
rect -332 822 -270 834
rect -240 1010 -178 1022
rect -240 834 -224 1010
rect -190 834 -178 1010
rect -240 822 -178 834
rect -122 1010 -60 1022
rect -122 834 -110 1010
rect -76 834 -60 1010
rect -122 822 -60 834
rect -30 1010 32 1022
rect -30 834 -14 1010
rect 20 834 32 1010
rect -30 822 32 834
rect 88 1010 150 1022
rect 88 834 100 1010
rect 134 834 150 1010
rect 88 822 150 834
rect 180 1010 242 1022
rect 180 834 196 1010
rect 230 834 242 1010
rect 180 822 242 834
rect 298 1010 360 1022
rect 298 834 310 1010
rect 344 834 360 1010
rect 298 822 360 834
rect 390 1010 452 1022
rect 390 834 406 1010
rect 440 834 452 1010
rect 390 822 452 834
rect 508 1010 570 1022
rect 508 834 520 1010
rect 554 834 570 1010
rect 508 822 570 834
rect 600 1010 662 1022
rect 600 834 616 1010
rect 650 834 662 1010
rect 600 822 662 834
rect 718 1010 780 1022
rect 718 834 730 1010
rect 764 834 780 1010
rect 718 822 780 834
rect 810 1010 872 1022
rect 810 834 826 1010
rect 860 834 872 1010
rect 810 822 872 834
rect 928 1010 990 1022
rect 928 834 940 1010
rect 974 834 990 1010
rect 928 822 990 834
rect 1020 1010 1082 1022
rect 1020 834 1036 1010
rect 1070 834 1082 1010
rect 1020 822 1082 834
rect 1138 1010 1200 1022
rect 1138 834 1150 1010
rect 1184 834 1200 1010
rect 1138 822 1200 834
rect 1230 1010 1292 1022
rect 1230 834 1246 1010
rect 1280 834 1292 1010
rect 1230 822 1292 834
rect 1348 1010 1410 1022
rect 1348 834 1360 1010
rect 1394 834 1410 1010
rect 1348 822 1410 834
rect 1440 1010 1502 1022
rect 1440 834 1456 1010
rect 1490 834 1502 1010
rect 1440 822 1502 834
rect 1558 1010 1620 1022
rect 1558 834 1570 1010
rect 1604 834 1620 1010
rect 1558 822 1620 834
rect 1650 1010 1712 1022
rect 1650 834 1666 1010
rect 1700 834 1712 1010
rect 1650 822 1712 834
rect 1768 1010 1830 1022
rect 1768 834 1780 1010
rect 1814 834 1830 1010
rect 1768 822 1830 834
rect 1860 1010 1922 1022
rect 1860 834 1876 1010
rect 1910 834 1922 1010
rect 1860 822 1922 834
rect 1978 1010 2040 1022
rect 1978 834 1990 1010
rect 2024 834 2040 1010
rect 1978 822 2040 834
rect 2070 1010 2132 1022
rect 2070 834 2086 1010
rect 2120 834 2132 1010
rect 2070 822 2132 834
rect 2188 1010 2250 1022
rect 2188 834 2200 1010
rect 2234 834 2250 1010
rect 2188 822 2250 834
rect 2280 1010 2342 1022
rect 2280 834 2296 1010
rect 2330 834 2342 1010
rect 2280 822 2342 834
rect 2398 1010 2460 1022
rect 2398 834 2410 1010
rect 2444 834 2460 1010
rect 2398 822 2460 834
rect 2490 1010 2552 1022
rect 2490 834 2506 1010
rect 2540 834 2552 1010
rect 2490 822 2552 834
rect 2608 1010 2670 1022
rect 2608 834 2620 1010
rect 2654 834 2670 1010
rect 2608 822 2670 834
rect 2700 1010 2762 1022
rect 2700 834 2716 1010
rect 2750 834 2762 1010
rect 2700 822 2762 834
rect 2818 1010 2880 1022
rect 2818 834 2830 1010
rect 2864 834 2880 1010
rect 2818 822 2880 834
rect 2910 1010 2972 1022
rect 2910 834 2926 1010
rect 2960 834 2972 1010
rect 2910 822 2972 834
rect 3028 1010 3090 1022
rect 3028 834 3040 1010
rect 3074 834 3090 1010
rect 3028 822 3090 834
rect 3120 1010 3182 1022
rect 3120 834 3136 1010
rect 3170 834 3182 1010
rect 3120 822 3182 834
rect 3238 1010 3300 1022
rect 3238 834 3250 1010
rect 3284 834 3300 1010
rect 3238 822 3300 834
rect 3330 1010 3392 1022
rect 3330 834 3346 1010
rect 3380 834 3392 1010
rect 3330 822 3392 834
rect 3448 1010 3510 1022
rect 3448 834 3460 1010
rect 3494 834 3510 1010
rect 3448 822 3510 834
rect 3540 1010 3602 1022
rect 3540 834 3556 1010
rect 3590 834 3602 1010
rect 3540 822 3602 834
rect 3658 1010 3720 1022
rect 3658 834 3670 1010
rect 3704 834 3720 1010
rect 3658 822 3720 834
rect 3750 1010 3812 1022
rect 3750 834 3766 1010
rect 3800 834 3812 1010
rect 3750 822 3812 834
rect 3868 1010 3930 1022
rect 3868 834 3880 1010
rect 3914 834 3930 1010
rect 3868 822 3930 834
rect 3960 1010 4022 1022
rect 3960 834 3976 1010
rect 4010 834 4022 1010
rect 3960 822 4022 834
rect 4078 1010 4140 1022
rect 4078 834 4090 1010
rect 4124 834 4140 1010
rect 4078 822 4140 834
rect 4170 1010 4232 1022
rect 4170 834 4186 1010
rect 4220 834 4232 1010
rect 4170 822 4232 834
rect 4288 1010 4350 1022
rect 4288 834 4300 1010
rect 4334 834 4350 1010
rect 4288 822 4350 834
rect 4380 1010 4442 1022
rect 4380 834 4396 1010
rect 4430 834 4442 1010
rect 4380 822 4442 834
rect 4498 1010 4560 1022
rect 4498 834 4510 1010
rect 4544 834 4560 1010
rect 4498 822 4560 834
rect 4590 1010 4652 1022
rect 4590 834 4606 1010
rect 4640 834 4652 1010
rect 4590 822 4652 834
rect 4708 1010 4770 1022
rect 4708 834 4720 1010
rect 4754 834 4770 1010
rect 4708 822 4770 834
rect 4800 1010 4862 1022
rect 4800 834 4816 1010
rect 4850 834 4862 1010
rect 4800 822 4862 834
rect 4918 1010 4980 1022
rect 4918 834 4930 1010
rect 4964 834 4980 1010
rect 4918 822 4980 834
rect 5010 1010 5072 1022
rect 5010 834 5026 1010
rect 5060 834 5072 1010
rect 5010 822 5072 834
rect 5128 1010 5190 1022
rect 5128 834 5140 1010
rect 5174 834 5190 1010
rect 5128 822 5190 834
rect 5220 1010 5282 1022
rect 5220 834 5236 1010
rect 5270 834 5282 1010
rect 5220 822 5282 834
rect 5338 1010 5400 1022
rect 5338 834 5350 1010
rect 5384 834 5400 1010
rect 5338 822 5400 834
rect 5430 1010 5492 1022
rect 5430 834 5446 1010
rect 5480 834 5492 1010
rect 5430 822 5492 834
rect 5548 1010 5610 1022
rect 5548 834 5560 1010
rect 5594 834 5610 1010
rect 5548 822 5610 834
rect 5640 1010 5702 1022
rect 5640 834 5656 1010
rect 5690 834 5702 1010
rect 5640 822 5702 834
rect 5758 1010 5820 1022
rect 5758 834 5770 1010
rect 5804 834 5820 1010
rect 5758 822 5820 834
rect 5850 1010 5912 1022
rect 5850 834 5866 1010
rect 5900 834 5912 1010
rect 5850 822 5912 834
rect 5968 1010 6030 1022
rect 5968 834 5980 1010
rect 6014 834 6030 1010
rect 5968 822 6030 834
rect 6060 1010 6122 1022
rect 6060 834 6076 1010
rect 6110 834 6122 1010
rect 6060 822 6122 834
rect 78 206 140 218
rect 78 30 90 206
rect 124 30 140 206
rect 78 18 140 30
rect 170 206 236 218
rect 170 30 186 206
rect 220 30 236 206
rect 170 18 236 30
rect 266 206 332 218
rect 266 30 282 206
rect 316 30 332 206
rect 266 18 332 30
rect 362 206 428 218
rect 362 30 378 206
rect 412 30 428 206
rect 362 18 428 30
rect 458 206 524 218
rect 458 30 474 206
rect 508 30 524 206
rect 458 18 524 30
rect 554 206 620 218
rect 554 30 570 206
rect 604 30 620 206
rect 554 18 620 30
rect 650 206 716 218
rect 650 30 666 206
rect 700 30 716 206
rect 650 18 716 30
rect 746 206 812 218
rect 746 30 762 206
rect 796 30 812 206
rect 746 18 812 30
rect 842 206 908 218
rect 842 30 858 206
rect 892 30 908 206
rect 842 18 908 30
rect 938 206 1004 218
rect 938 30 954 206
rect 988 30 1004 206
rect 938 18 1004 30
rect 1034 206 1100 218
rect 1034 30 1050 206
rect 1084 30 1100 206
rect 1034 18 1100 30
rect 1130 206 1196 218
rect 1130 30 1146 206
rect 1180 30 1196 206
rect 1130 18 1196 30
rect 1226 206 1292 218
rect 1226 30 1242 206
rect 1276 30 1292 206
rect 1226 18 1292 30
rect 1322 206 1388 218
rect 1322 30 1338 206
rect 1372 30 1388 206
rect 1322 18 1388 30
rect 1418 206 1484 218
rect 1418 30 1434 206
rect 1468 30 1484 206
rect 1418 18 1484 30
rect 1514 206 1580 218
rect 1514 30 1530 206
rect 1564 30 1580 206
rect 1514 18 1580 30
rect 1610 206 1676 218
rect 1610 30 1626 206
rect 1660 30 1676 206
rect 1610 18 1676 30
rect 1706 206 1772 218
rect 1706 30 1722 206
rect 1756 30 1772 206
rect 1706 18 1772 30
rect 1802 206 1868 218
rect 1802 30 1818 206
rect 1852 30 1868 206
rect 1802 18 1868 30
rect 1898 206 1964 218
rect 1898 30 1914 206
rect 1948 30 1964 206
rect 1898 18 1964 30
rect 1994 206 2060 218
rect 1994 30 2010 206
rect 2044 30 2060 206
rect 1994 18 2060 30
rect 2090 206 2156 218
rect 2090 30 2106 206
rect 2140 30 2156 206
rect 2090 18 2156 30
rect 2186 206 2252 218
rect 2186 30 2202 206
rect 2236 30 2252 206
rect 2186 18 2252 30
rect 2282 206 2348 218
rect 2282 30 2298 206
rect 2332 30 2348 206
rect 2282 18 2348 30
rect 2378 206 2444 218
rect 2378 30 2394 206
rect 2428 30 2444 206
rect 2378 18 2444 30
rect 2474 206 2540 218
rect 2474 30 2490 206
rect 2524 30 2540 206
rect 2474 18 2540 30
rect 2570 206 2636 218
rect 2570 30 2586 206
rect 2620 30 2636 206
rect 2570 18 2636 30
rect 2666 206 2732 218
rect 2666 30 2682 206
rect 2716 30 2732 206
rect 2666 18 2732 30
rect 2762 206 2828 218
rect 2762 30 2778 206
rect 2812 30 2828 206
rect 2762 18 2828 30
rect 2858 206 2924 218
rect 2858 30 2874 206
rect 2908 30 2924 206
rect 2858 18 2924 30
rect 2954 206 3020 218
rect 2954 30 2970 206
rect 3004 30 3020 206
rect 2954 18 3020 30
rect 3050 206 3116 218
rect 3050 30 3066 206
rect 3100 30 3116 206
rect 3050 18 3116 30
rect 3146 206 3212 218
rect 3146 30 3162 206
rect 3196 30 3212 206
rect 3146 18 3212 30
rect 3242 206 3308 218
rect 3242 30 3258 206
rect 3292 30 3308 206
rect 3242 18 3308 30
rect 3338 206 3400 218
rect 3338 30 3354 206
rect 3388 30 3400 206
rect 3338 18 3400 30
<< pdiff >>
rect 1505 10598 1679 10606
rect 1505 10564 1531 10598
rect 1565 10564 1633 10598
rect 1667 10564 1679 10598
rect 1505 10554 1679 10564
rect 1773 10598 1947 10606
rect 1773 10564 1785 10598
rect 1819 10564 1887 10598
rect 1921 10564 1947 10598
rect 1773 10554 1947 10564
rect 1505 9598 1679 9608
rect 1505 9564 1531 9598
rect 1565 9564 1633 9598
rect 1667 9564 1679 9598
rect 1505 9556 1679 9564
rect 1773 9598 1947 9608
rect 1773 9564 1785 9598
rect 1819 9564 1887 9598
rect 1921 9564 1947 9598
rect 1773 9556 1947 9564
rect 1479 9402 1679 9410
rect 1479 9368 1497 9402
rect 1531 9368 1565 9402
rect 1599 9368 1633 9402
rect 1667 9368 1679 9402
rect 1479 9358 1679 9368
rect 1773 9402 1973 9410
rect 1773 9368 1785 9402
rect 1819 9368 1853 9402
rect 1887 9368 1921 9402
rect 1955 9368 1973 9402
rect 1773 9358 1973 9368
rect 1479 9318 1679 9328
rect 1479 9284 1497 9318
rect 1531 9284 1565 9318
rect 1599 9284 1633 9318
rect 1667 9284 1679 9318
rect 1479 9274 1679 9284
rect 1773 9318 1973 9328
rect 1773 9284 1785 9318
rect 1819 9284 1853 9318
rect 1887 9284 1921 9318
rect 1955 9284 1973 9318
rect 1773 9274 1973 9284
rect 1479 9234 1679 9244
rect 1479 9200 1565 9234
rect 1599 9200 1633 9234
rect 1667 9200 1679 9234
rect 1479 9190 1679 9200
rect 1773 9234 1973 9244
rect 1773 9200 1785 9234
rect 1819 9200 1853 9234
rect 1887 9200 1973 9234
rect 1773 9190 1973 9200
rect 1479 9150 1679 9160
rect 1479 9116 1497 9150
rect 1531 9116 1565 9150
rect 1599 9116 1633 9150
rect 1667 9116 1679 9150
rect 1479 9106 1679 9116
rect 1773 9150 1973 9160
rect 1773 9116 1785 9150
rect 1819 9116 1853 9150
rect 1887 9116 1921 9150
rect 1955 9116 1973 9150
rect 1773 9106 1973 9116
rect 1479 9066 1679 9076
rect 1479 9032 1565 9066
rect 1599 9032 1633 9066
rect 1667 9032 1679 9066
rect 1479 9022 1679 9032
rect 1773 9066 1973 9076
rect 1773 9032 1785 9066
rect 1819 9032 1853 9066
rect 1887 9032 1973 9066
rect 1773 9022 1973 9032
rect 1479 8982 1679 8992
rect 1479 8948 1497 8982
rect 1531 8948 1565 8982
rect 1599 8948 1633 8982
rect 1667 8948 1679 8982
rect 1479 8938 1679 8948
rect 1773 8982 1973 8992
rect 1773 8948 1785 8982
rect 1819 8948 1853 8982
rect 1887 8948 1921 8982
rect 1955 8948 1973 8982
rect 1773 8938 1973 8948
rect 1479 8898 1679 8908
rect 1479 8864 1565 8898
rect 1599 8864 1633 8898
rect 1667 8864 1679 8898
rect 1479 8854 1679 8864
rect 1773 8898 1973 8908
rect 1773 8864 1785 8898
rect 1819 8864 1853 8898
rect 1887 8864 1973 8898
rect 1773 8854 1973 8864
rect 1479 8814 1679 8824
rect 1479 8780 1497 8814
rect 1531 8780 1565 8814
rect 1599 8780 1633 8814
rect 1667 8780 1679 8814
rect 1479 8770 1679 8780
rect 1773 8814 1973 8824
rect 1773 8780 1785 8814
rect 1819 8780 1853 8814
rect 1887 8780 1921 8814
rect 1955 8780 1973 8814
rect 1773 8770 1973 8780
rect 1479 8730 1679 8740
rect 1479 8696 1565 8730
rect 1599 8696 1633 8730
rect 1667 8696 1679 8730
rect 1479 8688 1679 8696
rect 1773 8730 1973 8740
rect 1773 8696 1785 8730
rect 1819 8696 1853 8730
rect 1887 8696 1973 8730
rect 1773 8688 1973 8696
rect 1479 8573 1679 8582
rect 1479 8539 1497 8573
rect 1531 8539 1565 8573
rect 1599 8539 1633 8573
rect 1667 8539 1679 8573
rect 1479 8529 1679 8539
rect 1773 8573 1973 8582
rect 1773 8539 1785 8573
rect 1819 8539 1853 8573
rect 1887 8539 1921 8573
rect 1955 8539 1973 8573
rect 1773 8529 1973 8539
rect 1479 8489 1679 8499
rect 1479 8455 1528 8489
rect 1562 8455 1609 8489
rect 1643 8455 1679 8489
rect 1479 8445 1679 8455
rect 1773 8489 1973 8499
rect 1773 8455 1809 8489
rect 1843 8455 1890 8489
rect 1924 8455 1973 8489
rect 1773 8445 1973 8455
rect 1479 8403 1679 8415
rect 1479 8369 1557 8403
rect 1591 8369 1625 8403
rect 1659 8369 1679 8403
rect 1479 8365 1679 8369
rect 1773 8403 1973 8415
rect 1773 8369 1793 8403
rect 1827 8369 1861 8403
rect 1895 8369 1973 8403
rect 1773 8365 1973 8369
rect 1543 8350 1671 8365
rect 1781 8350 1909 8365
rect 1543 8310 1671 8320
rect 1543 8276 1557 8310
rect 1591 8276 1625 8310
rect 1659 8276 1671 8310
rect 1543 8268 1671 8276
rect 1781 8310 1909 8320
rect 1781 8276 1793 8310
rect 1827 8276 1861 8310
rect 1895 8276 1909 8310
rect 1781 8268 1909 8276
rect -3569 7910 -3369 7922
rect -3569 7876 -3557 7910
rect -3381 7876 -3369 7910
rect -3569 7860 -3369 7876
rect -3569 7814 -3369 7830
rect -3569 7780 -3557 7814
rect -3381 7780 -3369 7814
rect -3569 7764 -3369 7780
rect -3569 7718 -3369 7734
rect -3569 7684 -3557 7718
rect -3381 7684 -3369 7718
rect -3569 7668 -3369 7684
rect -3569 7622 -3369 7638
rect -3569 7588 -3557 7622
rect -3381 7588 -3369 7622
rect -3569 7572 -3369 7588
rect -3569 7526 -3369 7542
rect -3569 7492 -3557 7526
rect -3381 7492 -3369 7526
rect -3569 7476 -3369 7492
rect -3569 7430 -3369 7446
rect -3569 7396 -3557 7430
rect -3381 7396 -3369 7430
rect -3569 7380 -3369 7396
rect -3569 7334 -3369 7350
rect -3569 7300 -3557 7334
rect -3381 7300 -3369 7334
rect -3569 7284 -3369 7300
rect -3569 7238 -3369 7254
rect -3569 7204 -3557 7238
rect -3381 7204 -3369 7238
rect -3569 7188 -3369 7204
rect -3569 7142 -3369 7158
rect -3569 7108 -3557 7142
rect -3381 7108 -3369 7142
rect -3569 7092 -3369 7108
rect -3569 7046 -3369 7062
rect -3569 7012 -3557 7046
rect -3381 7012 -3369 7046
rect -3569 6996 -3369 7012
rect -3569 6950 -3369 6966
rect -3569 6916 -3557 6950
rect -3381 6916 -3369 6950
rect -3569 6900 -3369 6916
rect -3569 6854 -3369 6870
rect -3569 6820 -3557 6854
rect -3381 6820 -3369 6854
rect -3569 6804 -3369 6820
rect -3569 6758 -3369 6774
rect -3569 6724 -3557 6758
rect -3381 6724 -3369 6758
rect -3569 6708 -3369 6724
rect -3569 6662 -3369 6678
rect -3569 6628 -3557 6662
rect -3381 6628 -3369 6662
rect -3569 6612 -3369 6628
rect -3569 6566 -3369 6582
rect -3569 6532 -3557 6566
rect -3381 6532 -3369 6566
rect -3569 6516 -3369 6532
rect -3569 6470 -3369 6486
rect -3569 6436 -3557 6470
rect -3381 6436 -3369 6470
rect -3569 6420 -3369 6436
rect -3569 6374 -3369 6390
rect -3569 6340 -3557 6374
rect -3381 6340 -3369 6374
rect -3569 6324 -3369 6340
rect -3569 6278 -3369 6294
rect -3569 6244 -3557 6278
rect -3381 6244 -3369 6278
rect -3569 6228 -3369 6244
rect -3569 6182 -3369 6198
rect -3569 6148 -3557 6182
rect -3381 6148 -3369 6182
rect -3569 6136 -3369 6148
rect -2656 7828 -2594 7840
rect -2656 7652 -2644 7828
rect -2610 7652 -2594 7828
rect -2656 7640 -2594 7652
rect -2564 7828 -2502 7840
rect -2564 7652 -2548 7828
rect -2514 7652 -2502 7828
rect -2564 7640 -2502 7652
rect -2446 7828 -2384 7840
rect -2446 7652 -2434 7828
rect -2400 7652 -2384 7828
rect -2446 7640 -2384 7652
rect -2354 7828 -2292 7840
rect -2354 7652 -2338 7828
rect -2304 7652 -2292 7828
rect -2354 7640 -2292 7652
rect -2236 7828 -2174 7840
rect -2236 7652 -2224 7828
rect -2190 7652 -2174 7828
rect -2236 7640 -2174 7652
rect -2144 7828 -2082 7840
rect -2144 7652 -2128 7828
rect -2094 7652 -2082 7828
rect -2144 7640 -2082 7652
rect -2026 7828 -1964 7840
rect -2026 7652 -2014 7828
rect -1980 7652 -1964 7828
rect -2026 7640 -1964 7652
rect -1934 7828 -1872 7840
rect -1934 7652 -1918 7828
rect -1884 7652 -1872 7828
rect -1934 7640 -1872 7652
rect -1816 7828 -1754 7840
rect -1816 7652 -1804 7828
rect -1770 7652 -1754 7828
rect -1816 7640 -1754 7652
rect -1724 7828 -1662 7840
rect -1724 7652 -1708 7828
rect -1674 7652 -1662 7828
rect -1724 7640 -1662 7652
rect -1606 7828 -1544 7840
rect -1606 7652 -1594 7828
rect -1560 7652 -1544 7828
rect -1606 7640 -1544 7652
rect -1514 7828 -1452 7840
rect -1514 7652 -1498 7828
rect -1464 7652 -1452 7828
rect -1514 7640 -1452 7652
rect -1396 7828 -1334 7840
rect -1396 7652 -1384 7828
rect -1350 7652 -1334 7828
rect -1396 7640 -1334 7652
rect -1304 7828 -1242 7840
rect -1304 7652 -1288 7828
rect -1254 7652 -1242 7828
rect -1304 7640 -1242 7652
rect -1186 7828 -1124 7840
rect -1186 7652 -1174 7828
rect -1140 7652 -1124 7828
rect -1186 7640 -1124 7652
rect -1094 7828 -1032 7840
rect -1094 7652 -1078 7828
rect -1044 7652 -1032 7828
rect -1094 7640 -1032 7652
rect -976 7828 -914 7840
rect -976 7652 -964 7828
rect -930 7652 -914 7828
rect -976 7640 -914 7652
rect -884 7828 -822 7840
rect -884 7652 -868 7828
rect -834 7652 -822 7828
rect -884 7640 -822 7652
rect -766 7828 -704 7840
rect -766 7652 -754 7828
rect -720 7652 -704 7828
rect -766 7640 -704 7652
rect -674 7828 -612 7840
rect -674 7652 -658 7828
rect -624 7652 -612 7828
rect -674 7640 -612 7652
rect -556 7828 -494 7840
rect -556 7652 -544 7828
rect -510 7652 -494 7828
rect -556 7640 -494 7652
rect -464 7828 -402 7840
rect -464 7652 -448 7828
rect -414 7652 -402 7828
rect -464 7640 -402 7652
rect -346 7828 -284 7840
rect -346 7652 -334 7828
rect -300 7652 -284 7828
rect -346 7640 -284 7652
rect -254 7828 -192 7840
rect -254 7652 -238 7828
rect -204 7652 -192 7828
rect -254 7640 -192 7652
rect -136 7828 -74 7840
rect -136 7652 -124 7828
rect -90 7652 -74 7828
rect -136 7640 -74 7652
rect -44 7828 18 7840
rect -44 7652 -28 7828
rect 6 7652 18 7828
rect -44 7640 18 7652
rect 74 7828 136 7840
rect 74 7652 86 7828
rect 120 7652 136 7828
rect 74 7640 136 7652
rect 166 7828 228 7840
rect 166 7652 182 7828
rect 216 7652 228 7828
rect 166 7640 228 7652
rect 284 7828 346 7840
rect 284 7652 296 7828
rect 330 7652 346 7828
rect 284 7640 346 7652
rect 376 7828 438 7840
rect 376 7652 392 7828
rect 426 7652 438 7828
rect 376 7640 438 7652
rect 494 7828 556 7840
rect 494 7652 506 7828
rect 540 7652 556 7828
rect 494 7640 556 7652
rect 586 7828 648 7840
rect 586 7652 602 7828
rect 636 7652 648 7828
rect 586 7640 648 7652
rect 704 7828 766 7840
rect 704 7652 716 7828
rect 750 7652 766 7828
rect 704 7640 766 7652
rect 796 7828 858 7840
rect 796 7652 812 7828
rect 846 7652 858 7828
rect 796 7640 858 7652
rect 914 7828 976 7840
rect 914 7652 926 7828
rect 960 7652 976 7828
rect 914 7640 976 7652
rect 1006 7828 1068 7840
rect 1006 7652 1022 7828
rect 1056 7652 1068 7828
rect 1006 7640 1068 7652
rect 1124 7828 1186 7840
rect 1124 7652 1136 7828
rect 1170 7652 1186 7828
rect 1124 7640 1186 7652
rect 1216 7828 1278 7840
rect 1216 7652 1232 7828
rect 1266 7652 1278 7828
rect 1216 7640 1278 7652
rect 1334 7828 1396 7840
rect 1334 7652 1346 7828
rect 1380 7652 1396 7828
rect 1334 7640 1396 7652
rect 1426 7828 1488 7840
rect 1426 7652 1442 7828
rect 1476 7652 1488 7828
rect 1426 7640 1488 7652
rect 1544 7828 1606 7840
rect 1544 7652 1556 7828
rect 1590 7652 1606 7828
rect 1544 7640 1606 7652
rect 1636 7828 1698 7840
rect 1636 7652 1652 7828
rect 1686 7652 1698 7828
rect 1636 7640 1698 7652
rect 1754 7828 1816 7840
rect 1754 7652 1766 7828
rect 1800 7652 1816 7828
rect 1754 7640 1816 7652
rect 1846 7828 1908 7840
rect 1846 7652 1862 7828
rect 1896 7652 1908 7828
rect 1846 7640 1908 7652
rect 1964 7828 2026 7840
rect 1964 7652 1976 7828
rect 2010 7652 2026 7828
rect 1964 7640 2026 7652
rect 2056 7828 2118 7840
rect 2056 7652 2072 7828
rect 2106 7652 2118 7828
rect 2056 7640 2118 7652
rect 2174 7828 2236 7840
rect 2174 7652 2186 7828
rect 2220 7652 2236 7828
rect 2174 7640 2236 7652
rect 2266 7828 2328 7840
rect 2266 7652 2282 7828
rect 2316 7652 2328 7828
rect 2266 7640 2328 7652
rect 2384 7828 2446 7840
rect 2384 7652 2396 7828
rect 2430 7652 2446 7828
rect 2384 7640 2446 7652
rect 2476 7828 2538 7840
rect 2476 7652 2492 7828
rect 2526 7652 2538 7828
rect 2476 7640 2538 7652
rect 2594 7828 2656 7840
rect 2594 7652 2606 7828
rect 2640 7652 2656 7828
rect 2594 7640 2656 7652
rect 2686 7828 2748 7840
rect 2686 7652 2702 7828
rect 2736 7652 2748 7828
rect 2686 7640 2748 7652
rect 2804 7828 2866 7840
rect 2804 7652 2816 7828
rect 2850 7652 2866 7828
rect 2804 7640 2866 7652
rect 2896 7828 2958 7840
rect 2896 7652 2912 7828
rect 2946 7652 2958 7828
rect 2896 7640 2958 7652
rect 3014 7828 3076 7840
rect 3014 7652 3026 7828
rect 3060 7652 3076 7828
rect 3014 7640 3076 7652
rect 3106 7828 3168 7840
rect 3106 7652 3122 7828
rect 3156 7652 3168 7828
rect 3106 7640 3168 7652
rect 3224 7828 3286 7840
rect 3224 7652 3236 7828
rect 3270 7652 3286 7828
rect 3224 7640 3286 7652
rect 3316 7828 3378 7840
rect 3316 7652 3332 7828
rect 3366 7652 3378 7828
rect 3316 7640 3378 7652
rect 3434 7828 3496 7840
rect 3434 7652 3446 7828
rect 3480 7652 3496 7828
rect 3434 7640 3496 7652
rect 3526 7828 3588 7840
rect 3526 7652 3542 7828
rect 3576 7652 3588 7828
rect 3526 7640 3588 7652
rect 3644 7828 3706 7840
rect 3644 7652 3656 7828
rect 3690 7652 3706 7828
rect 3644 7640 3706 7652
rect 3736 7828 3798 7840
rect 3736 7652 3752 7828
rect 3786 7652 3798 7828
rect 3736 7640 3798 7652
rect 3854 7828 3916 7840
rect 3854 7652 3866 7828
rect 3900 7652 3916 7828
rect 3854 7640 3916 7652
rect 3946 7828 4008 7840
rect 3946 7652 3962 7828
rect 3996 7652 4008 7828
rect 3946 7640 4008 7652
rect 4064 7828 4126 7840
rect 4064 7652 4076 7828
rect 4110 7652 4126 7828
rect 4064 7640 4126 7652
rect 4156 7828 4218 7840
rect 4156 7652 4172 7828
rect 4206 7652 4218 7828
rect 4156 7640 4218 7652
rect 4274 7828 4336 7840
rect 4274 7652 4286 7828
rect 4320 7652 4336 7828
rect 4274 7640 4336 7652
rect 4366 7828 4428 7840
rect 4366 7652 4382 7828
rect 4416 7652 4428 7828
rect 4366 7640 4428 7652
rect 4484 7828 4546 7840
rect 4484 7652 4496 7828
rect 4530 7652 4546 7828
rect 4484 7640 4546 7652
rect 4576 7828 4638 7840
rect 4576 7652 4592 7828
rect 4626 7652 4638 7828
rect 4576 7640 4638 7652
rect 4694 7828 4756 7840
rect 4694 7652 4706 7828
rect 4740 7652 4756 7828
rect 4694 7640 4756 7652
rect 4786 7828 4848 7840
rect 4786 7652 4802 7828
rect 4836 7652 4848 7828
rect 4786 7640 4848 7652
rect 4904 7828 4966 7840
rect 4904 7652 4916 7828
rect 4950 7652 4966 7828
rect 4904 7640 4966 7652
rect 4996 7828 5058 7840
rect 4996 7652 5012 7828
rect 5046 7652 5058 7828
rect 4996 7640 5058 7652
rect 5114 7828 5176 7840
rect 5114 7652 5126 7828
rect 5160 7652 5176 7828
rect 5114 7640 5176 7652
rect 5206 7828 5268 7840
rect 5206 7652 5222 7828
rect 5256 7652 5268 7828
rect 5206 7640 5268 7652
rect 5324 7828 5386 7840
rect 5324 7652 5336 7828
rect 5370 7652 5386 7828
rect 5324 7640 5386 7652
rect 5416 7828 5478 7840
rect 5416 7652 5432 7828
rect 5466 7652 5478 7828
rect 5416 7640 5478 7652
rect 5534 7828 5596 7840
rect 5534 7652 5546 7828
rect 5580 7652 5596 7828
rect 5534 7640 5596 7652
rect 5626 7828 5688 7840
rect 5626 7652 5642 7828
rect 5676 7652 5688 7828
rect 5626 7640 5688 7652
rect 5744 7828 5806 7840
rect 5744 7652 5756 7828
rect 5790 7652 5806 7828
rect 5744 7640 5806 7652
rect 5836 7828 5898 7840
rect 5836 7652 5852 7828
rect 5886 7652 5898 7828
rect 5836 7640 5898 7652
rect 5954 7828 6016 7840
rect 5954 7652 5966 7828
rect 6000 7652 6016 7828
rect 5954 7640 6016 7652
rect 6046 7828 6108 7840
rect 6046 7652 6062 7828
rect 6096 7652 6108 7828
rect 6046 7640 6108 7652
rect -2654 7295 -2592 7307
rect -2654 7119 -2642 7295
rect -2608 7119 -2592 7295
rect -2654 7107 -2592 7119
rect -2562 7295 -2500 7307
rect -2562 7119 -2546 7295
rect -2512 7119 -2500 7295
rect -2562 7107 -2500 7119
rect -2444 7295 -2382 7307
rect -2444 7119 -2432 7295
rect -2398 7119 -2382 7295
rect -2444 7107 -2382 7119
rect -2352 7295 -2290 7307
rect -2352 7119 -2336 7295
rect -2302 7119 -2290 7295
rect -2352 7107 -2290 7119
rect -2234 7295 -2172 7307
rect -2234 7119 -2222 7295
rect -2188 7119 -2172 7295
rect -2234 7107 -2172 7119
rect -2142 7295 -2080 7307
rect -2142 7119 -2126 7295
rect -2092 7119 -2080 7295
rect -2142 7107 -2080 7119
rect -2024 7295 -1962 7307
rect -2024 7119 -2012 7295
rect -1978 7119 -1962 7295
rect -2024 7107 -1962 7119
rect -1932 7295 -1870 7307
rect -1932 7119 -1916 7295
rect -1882 7119 -1870 7295
rect -1932 7107 -1870 7119
rect -1814 7295 -1752 7307
rect -1814 7119 -1802 7295
rect -1768 7119 -1752 7295
rect -1814 7107 -1752 7119
rect -1722 7295 -1660 7307
rect -1722 7119 -1706 7295
rect -1672 7119 -1660 7295
rect -1722 7107 -1660 7119
rect -1604 7295 -1542 7307
rect -1604 7119 -1592 7295
rect -1558 7119 -1542 7295
rect -1604 7107 -1542 7119
rect -1512 7295 -1450 7307
rect -1512 7119 -1496 7295
rect -1462 7119 -1450 7295
rect -1512 7107 -1450 7119
rect -1394 7295 -1332 7307
rect -1394 7119 -1382 7295
rect -1348 7119 -1332 7295
rect -1394 7107 -1332 7119
rect -1302 7295 -1240 7307
rect -1302 7119 -1286 7295
rect -1252 7119 -1240 7295
rect -1302 7107 -1240 7119
rect -1184 7295 -1122 7307
rect -1184 7119 -1172 7295
rect -1138 7119 -1122 7295
rect -1184 7107 -1122 7119
rect -1092 7295 -1030 7307
rect -1092 7119 -1076 7295
rect -1042 7119 -1030 7295
rect -1092 7107 -1030 7119
rect -974 7295 -912 7307
rect -974 7119 -962 7295
rect -928 7119 -912 7295
rect -974 7107 -912 7119
rect -882 7295 -820 7307
rect -882 7119 -866 7295
rect -832 7119 -820 7295
rect -882 7107 -820 7119
rect -764 7295 -702 7307
rect -764 7119 -752 7295
rect -718 7119 -702 7295
rect -764 7107 -702 7119
rect -672 7295 -610 7307
rect -672 7119 -656 7295
rect -622 7119 -610 7295
rect -672 7107 -610 7119
rect -554 7295 -492 7307
rect -554 7119 -542 7295
rect -508 7119 -492 7295
rect -554 7107 -492 7119
rect -462 7295 -400 7307
rect -462 7119 -446 7295
rect -412 7119 -400 7295
rect -462 7107 -400 7119
rect -344 7295 -282 7307
rect -344 7119 -332 7295
rect -298 7119 -282 7295
rect -344 7107 -282 7119
rect -252 7295 -190 7307
rect -252 7119 -236 7295
rect -202 7119 -190 7295
rect -252 7107 -190 7119
rect -134 7295 -72 7307
rect -134 7119 -122 7295
rect -88 7119 -72 7295
rect -134 7107 -72 7119
rect -42 7295 20 7307
rect -42 7119 -26 7295
rect 8 7119 20 7295
rect -42 7107 20 7119
rect 76 7295 138 7307
rect 76 7119 88 7295
rect 122 7119 138 7295
rect 76 7107 138 7119
rect 168 7295 230 7307
rect 168 7119 184 7295
rect 218 7119 230 7295
rect 168 7107 230 7119
rect 286 7295 348 7307
rect 286 7119 298 7295
rect 332 7119 348 7295
rect 286 7107 348 7119
rect 378 7295 440 7307
rect 378 7119 394 7295
rect 428 7119 440 7295
rect 378 7107 440 7119
rect 496 7295 558 7307
rect 496 7119 508 7295
rect 542 7119 558 7295
rect 496 7107 558 7119
rect 588 7295 650 7307
rect 588 7119 604 7295
rect 638 7119 650 7295
rect 588 7107 650 7119
rect 706 7295 768 7307
rect 706 7119 718 7295
rect 752 7119 768 7295
rect 706 7107 768 7119
rect 798 7295 860 7307
rect 798 7119 814 7295
rect 848 7119 860 7295
rect 798 7107 860 7119
rect 916 7295 978 7307
rect 916 7119 928 7295
rect 962 7119 978 7295
rect 916 7107 978 7119
rect 1008 7295 1070 7307
rect 1008 7119 1024 7295
rect 1058 7119 1070 7295
rect 1008 7107 1070 7119
rect 1126 7295 1188 7307
rect 1126 7119 1138 7295
rect 1172 7119 1188 7295
rect 1126 7107 1188 7119
rect 1218 7295 1280 7307
rect 1218 7119 1234 7295
rect 1268 7119 1280 7295
rect 1218 7107 1280 7119
rect 1336 7295 1398 7307
rect 1336 7119 1348 7295
rect 1382 7119 1398 7295
rect 1336 7107 1398 7119
rect 1428 7295 1490 7307
rect 1428 7119 1444 7295
rect 1478 7119 1490 7295
rect 1428 7107 1490 7119
rect 1546 7295 1608 7307
rect 1546 7119 1558 7295
rect 1592 7119 1608 7295
rect 1546 7107 1608 7119
rect 1638 7295 1700 7307
rect 1638 7119 1654 7295
rect 1688 7119 1700 7295
rect 1638 7107 1700 7119
rect 1756 7295 1818 7307
rect 1756 7119 1768 7295
rect 1802 7119 1818 7295
rect 1756 7107 1818 7119
rect 1848 7295 1910 7307
rect 1848 7119 1864 7295
rect 1898 7119 1910 7295
rect 1848 7107 1910 7119
rect 1966 7295 2028 7307
rect 1966 7119 1978 7295
rect 2012 7119 2028 7295
rect 1966 7107 2028 7119
rect 2058 7295 2120 7307
rect 2058 7119 2074 7295
rect 2108 7119 2120 7295
rect 2058 7107 2120 7119
rect 2176 7295 2238 7307
rect 2176 7119 2188 7295
rect 2222 7119 2238 7295
rect 2176 7107 2238 7119
rect 2268 7295 2330 7307
rect 2268 7119 2284 7295
rect 2318 7119 2330 7295
rect 2268 7107 2330 7119
rect 2386 7295 2448 7307
rect 2386 7119 2398 7295
rect 2432 7119 2448 7295
rect 2386 7107 2448 7119
rect 2478 7295 2540 7307
rect 2478 7119 2494 7295
rect 2528 7119 2540 7295
rect 2478 7107 2540 7119
rect 2596 7295 2658 7307
rect 2596 7119 2608 7295
rect 2642 7119 2658 7295
rect 2596 7107 2658 7119
rect 2688 7295 2750 7307
rect 2688 7119 2704 7295
rect 2738 7119 2750 7295
rect 2688 7107 2750 7119
rect 2806 7295 2868 7307
rect 2806 7119 2818 7295
rect 2852 7119 2868 7295
rect 2806 7107 2868 7119
rect 2898 7295 2960 7307
rect 2898 7119 2914 7295
rect 2948 7119 2960 7295
rect 2898 7107 2960 7119
rect 3016 7295 3078 7307
rect 3016 7119 3028 7295
rect 3062 7119 3078 7295
rect 3016 7107 3078 7119
rect 3108 7295 3170 7307
rect 3108 7119 3124 7295
rect 3158 7119 3170 7295
rect 3108 7107 3170 7119
rect 3226 7295 3288 7307
rect 3226 7119 3238 7295
rect 3272 7119 3288 7295
rect 3226 7107 3288 7119
rect 3318 7295 3380 7307
rect 3318 7119 3334 7295
rect 3368 7119 3380 7295
rect 3318 7107 3380 7119
rect 3436 7295 3498 7307
rect 3436 7119 3448 7295
rect 3482 7119 3498 7295
rect 3436 7107 3498 7119
rect 3528 7295 3590 7307
rect 3528 7119 3544 7295
rect 3578 7119 3590 7295
rect 3528 7107 3590 7119
rect 3646 7295 3708 7307
rect 3646 7119 3658 7295
rect 3692 7119 3708 7295
rect 3646 7107 3708 7119
rect 3738 7295 3800 7307
rect 3738 7119 3754 7295
rect 3788 7119 3800 7295
rect 3738 7107 3800 7119
rect 3856 7295 3918 7307
rect 3856 7119 3868 7295
rect 3902 7119 3918 7295
rect 3856 7107 3918 7119
rect 3948 7295 4010 7307
rect 3948 7119 3964 7295
rect 3998 7119 4010 7295
rect 3948 7107 4010 7119
rect 4066 7295 4128 7307
rect 4066 7119 4078 7295
rect 4112 7119 4128 7295
rect 4066 7107 4128 7119
rect 4158 7295 4220 7307
rect 4158 7119 4174 7295
rect 4208 7119 4220 7295
rect 4158 7107 4220 7119
rect 4276 7295 4338 7307
rect 4276 7119 4288 7295
rect 4322 7119 4338 7295
rect 4276 7107 4338 7119
rect 4368 7295 4430 7307
rect 4368 7119 4384 7295
rect 4418 7119 4430 7295
rect 4368 7107 4430 7119
rect 4486 7295 4548 7307
rect 4486 7119 4498 7295
rect 4532 7119 4548 7295
rect 4486 7107 4548 7119
rect 4578 7295 4640 7307
rect 4578 7119 4594 7295
rect 4628 7119 4640 7295
rect 4578 7107 4640 7119
rect 4696 7295 4758 7307
rect 4696 7119 4708 7295
rect 4742 7119 4758 7295
rect 4696 7107 4758 7119
rect 4788 7295 4850 7307
rect 4788 7119 4804 7295
rect 4838 7119 4850 7295
rect 4788 7107 4850 7119
rect 4906 7295 4968 7307
rect 4906 7119 4918 7295
rect 4952 7119 4968 7295
rect 4906 7107 4968 7119
rect 4998 7295 5060 7307
rect 4998 7119 5014 7295
rect 5048 7119 5060 7295
rect 4998 7107 5060 7119
rect 5116 7295 5178 7307
rect 5116 7119 5128 7295
rect 5162 7119 5178 7295
rect 5116 7107 5178 7119
rect 5208 7295 5270 7307
rect 5208 7119 5224 7295
rect 5258 7119 5270 7295
rect 5208 7107 5270 7119
rect 5326 7295 5388 7307
rect 5326 7119 5338 7295
rect 5372 7119 5388 7295
rect 5326 7107 5388 7119
rect 5418 7295 5480 7307
rect 5418 7119 5434 7295
rect 5468 7119 5480 7295
rect 5418 7107 5480 7119
rect 5536 7295 5598 7307
rect 5536 7119 5548 7295
rect 5582 7119 5598 7295
rect 5536 7107 5598 7119
rect 5628 7295 5690 7307
rect 5628 7119 5644 7295
rect 5678 7119 5690 7295
rect 5628 7107 5690 7119
rect 5746 7295 5808 7307
rect 5746 7119 5758 7295
rect 5792 7119 5808 7295
rect 5746 7107 5808 7119
rect 5838 7295 5900 7307
rect 5838 7119 5854 7295
rect 5888 7119 5900 7295
rect 5838 7107 5900 7119
rect 5956 7295 6018 7307
rect 5956 7119 5968 7295
rect 6002 7119 6018 7295
rect 5956 7107 6018 7119
rect 6048 7295 6110 7307
rect 6048 7119 6064 7295
rect 6098 7119 6110 7295
rect 6048 7107 6110 7119
rect -3567 5500 -3367 5512
rect -3567 5466 -3555 5500
rect -3379 5466 -3367 5500
rect -3567 5450 -3367 5466
rect -3567 5404 -3367 5420
rect -3567 5370 -3555 5404
rect -3379 5370 -3367 5404
rect -3567 5354 -3367 5370
rect -3567 5308 -3367 5324
rect -3567 5274 -3555 5308
rect -3379 5274 -3367 5308
rect -3567 5258 -3367 5274
rect -3567 5212 -3367 5228
rect -3567 5178 -3555 5212
rect -3379 5178 -3367 5212
rect -3567 5162 -3367 5178
rect -3567 5116 -3367 5132
rect -3567 5082 -3555 5116
rect -3379 5082 -3367 5116
rect -3567 5066 -3367 5082
rect -3567 5020 -3367 5036
rect -3567 4986 -3555 5020
rect -3379 4986 -3367 5020
rect -3567 4970 -3367 4986
rect -3567 4924 -3367 4940
rect -3567 4890 -3555 4924
rect -3379 4890 -3367 4924
rect -3567 4874 -3367 4890
rect -3567 4828 -3367 4844
rect -3567 4794 -3555 4828
rect -3379 4794 -3367 4828
rect -3567 4778 -3367 4794
rect -3567 4732 -3367 4748
rect -3567 4698 -3555 4732
rect -3379 4698 -3367 4732
rect -3567 4682 -3367 4698
rect -3567 4636 -3367 4652
rect -3567 4602 -3555 4636
rect -3379 4602 -3367 4636
rect -3567 4586 -3367 4602
rect -3567 4540 -3367 4556
rect -3567 4506 -3555 4540
rect -3379 4506 -3367 4540
rect -3567 4490 -3367 4506
rect -3567 4444 -3367 4460
rect -3567 4410 -3555 4444
rect -3379 4410 -3367 4444
rect -3567 4394 -3367 4410
rect -3567 4348 -3367 4364
rect -3567 4314 -3555 4348
rect -3379 4314 -3367 4348
rect -3567 4298 -3367 4314
rect -3567 4252 -3367 4268
rect -3567 4218 -3555 4252
rect -3379 4218 -3367 4252
rect -3567 4202 -3367 4218
rect -3567 4156 -3367 4172
rect -3567 4122 -3555 4156
rect -3379 4122 -3367 4156
rect -3567 4106 -3367 4122
rect -3567 4060 -3367 4076
rect -3567 4026 -3555 4060
rect -3379 4026 -3367 4060
rect -3567 4010 -3367 4026
rect -3567 3964 -3367 3980
rect -3567 3930 -3555 3964
rect -3379 3930 -3367 3964
rect -3567 3914 -3367 3930
rect -3567 3868 -3367 3884
rect -3567 3834 -3555 3868
rect -3379 3834 -3367 3868
rect -3567 3818 -3367 3834
rect -3567 3772 -3367 3788
rect -3567 3738 -3555 3772
rect -3379 3738 -3367 3772
rect -3567 3726 -3367 3738
rect 6831 7910 7031 7922
rect 6831 7876 6843 7910
rect 7019 7876 7031 7910
rect 6831 7860 7031 7876
rect 6831 7814 7031 7830
rect 6831 7780 6843 7814
rect 7019 7780 7031 7814
rect 6831 7764 7031 7780
rect 6831 7718 7031 7734
rect 6831 7684 6843 7718
rect 7019 7684 7031 7718
rect 6831 7668 7031 7684
rect 6831 7622 7031 7638
rect 6831 7588 6843 7622
rect 7019 7588 7031 7622
rect 6831 7572 7031 7588
rect 6831 7526 7031 7542
rect 6831 7492 6843 7526
rect 7019 7492 7031 7526
rect 6831 7476 7031 7492
rect 6831 7430 7031 7446
rect 6831 7396 6843 7430
rect 7019 7396 7031 7430
rect 6831 7380 7031 7396
rect 6831 7334 7031 7350
rect 6831 7300 6843 7334
rect 7019 7300 7031 7334
rect 6831 7284 7031 7300
rect 6831 7238 7031 7254
rect 6831 7204 6843 7238
rect 7019 7204 7031 7238
rect 6831 7188 7031 7204
rect 6831 7142 7031 7158
rect 6831 7108 6843 7142
rect 7019 7108 7031 7142
rect 6831 7092 7031 7108
rect 6831 7046 7031 7062
rect 6831 7012 6843 7046
rect 7019 7012 7031 7046
rect 6831 6996 7031 7012
rect 6831 6950 7031 6966
rect 6831 6916 6843 6950
rect 7019 6916 7031 6950
rect 6831 6900 7031 6916
rect 6831 6854 7031 6870
rect 6831 6820 6843 6854
rect 7019 6820 7031 6854
rect 6831 6804 7031 6820
rect 6831 6758 7031 6774
rect 6831 6724 6843 6758
rect 7019 6724 7031 6758
rect 6831 6708 7031 6724
rect 6831 6662 7031 6678
rect 6831 6628 6843 6662
rect 7019 6628 7031 6662
rect 6831 6612 7031 6628
rect 6831 6566 7031 6582
rect 6831 6532 6843 6566
rect 7019 6532 7031 6566
rect 6831 6516 7031 6532
rect 6831 6470 7031 6486
rect 6831 6436 6843 6470
rect 7019 6436 7031 6470
rect 6831 6420 7031 6436
rect 6831 6374 7031 6390
rect 6831 6340 6843 6374
rect 7019 6340 7031 6374
rect 6831 6324 7031 6340
rect 6831 6278 7031 6294
rect 6831 6244 6843 6278
rect 7019 6244 7031 6278
rect 6831 6228 7031 6244
rect 6831 6182 7031 6198
rect 6831 6148 6843 6182
rect 7019 6148 7031 6182
rect 6831 6136 7031 6148
rect 6831 5500 7031 5512
rect 6831 5466 6843 5500
rect 7019 5466 7031 5500
rect 6831 5450 7031 5466
rect 6831 5404 7031 5420
rect 6831 5370 6843 5404
rect 7019 5370 7031 5404
rect 6831 5354 7031 5370
rect 6831 5308 7031 5324
rect 6831 5274 6843 5308
rect 7019 5274 7031 5308
rect 6831 5258 7031 5274
rect 6831 5212 7031 5228
rect 6831 5178 6843 5212
rect 7019 5178 7031 5212
rect 6831 5162 7031 5178
rect 6831 5116 7031 5132
rect 6831 5082 6843 5116
rect 7019 5082 7031 5116
rect 6831 5066 7031 5082
rect 6831 5020 7031 5036
rect 6831 4986 6843 5020
rect 7019 4986 7031 5020
rect 6831 4970 7031 4986
rect 6831 4924 7031 4940
rect 6831 4890 6843 4924
rect 7019 4890 7031 4924
rect 6831 4874 7031 4890
rect 6831 4828 7031 4844
rect 6831 4794 6843 4828
rect 7019 4794 7031 4828
rect 6831 4778 7031 4794
rect 6831 4732 7031 4748
rect 6831 4698 6843 4732
rect 7019 4698 7031 4732
rect 6831 4682 7031 4698
rect 6831 4636 7031 4652
rect 6831 4602 6843 4636
rect 7019 4602 7031 4636
rect 6831 4586 7031 4602
rect 6831 4540 7031 4556
rect 6831 4506 6843 4540
rect 7019 4506 7031 4540
rect 6831 4490 7031 4506
rect 6831 4444 7031 4460
rect 6831 4410 6843 4444
rect 7019 4410 7031 4444
rect 6831 4394 7031 4410
rect 6831 4348 7031 4364
rect 6831 4314 6843 4348
rect 7019 4314 7031 4348
rect 6831 4298 7031 4314
rect 6831 4252 7031 4268
rect 6831 4218 6843 4252
rect 7019 4218 7031 4252
rect 6831 4202 7031 4218
rect 6831 4156 7031 4172
rect 6831 4122 6843 4156
rect 7019 4122 7031 4156
rect 6831 4106 7031 4122
rect 6831 4060 7031 4076
rect 6831 4026 6843 4060
rect 7019 4026 7031 4060
rect 6831 4010 7031 4026
rect 6831 3964 7031 3980
rect 6831 3930 6843 3964
rect 7019 3930 7031 3964
rect 6831 3914 7031 3930
rect 6831 3868 7031 3884
rect 6831 3834 6843 3868
rect 7019 3834 7031 3868
rect 6831 3818 7031 3834
rect 6831 3772 7031 3788
rect 6831 3738 6843 3772
rect 7019 3738 7031 3772
rect 6831 3726 7031 3738
<< ndiffc >>
rect 1260 10564 1294 10598
rect 2158 10564 2192 10598
rect 1260 9564 1294 9598
rect 2158 9564 2192 9598
rect 1241 9368 1275 9402
rect 1309 9368 1343 9402
rect 2109 9368 2143 9402
rect 2177 9368 2211 9402
rect 1241 9284 1275 9318
rect 2177 9284 2211 9318
rect 1241 9200 1275 9234
rect 1309 9200 1343 9234
rect 2109 9200 2143 9234
rect 2177 9200 2211 9234
rect 1241 9116 1275 9150
rect 2177 9116 2211 9150
rect 1241 9032 1275 9066
rect 1309 9032 1343 9066
rect 2109 9032 2143 9066
rect 2177 9032 2211 9066
rect 1309 8948 1343 8982
rect 2109 8948 2143 8982
rect 1241 8864 1275 8898
rect 2177 8864 2211 8898
rect 1309 8780 1343 8814
rect 2109 8780 2143 8814
rect 1241 8696 1275 8730
rect 1309 8696 1343 8730
rect 2109 8696 2143 8730
rect 2177 8696 2211 8730
rect 1245 8539 1279 8573
rect 1313 8539 1347 8573
rect 2105 8539 2139 8573
rect 2173 8539 2207 8573
rect 1271 8455 1305 8489
rect 2147 8455 2181 8489
rect 1241 8369 1275 8403
rect 2177 8369 2211 8403
rect 1254 8276 1288 8310
rect 2164 8276 2198 8310
rect -2630 6169 -2596 6345
rect -2534 6169 -2500 6345
rect -2420 6169 -2386 6345
rect -2324 6169 -2290 6345
rect -2210 6169 -2176 6345
rect -2114 6169 -2080 6345
rect -2000 6169 -1966 6345
rect -1904 6169 -1870 6345
rect -1790 6169 -1756 6345
rect -1694 6169 -1660 6345
rect -1580 6169 -1546 6345
rect -1484 6169 -1450 6345
rect -1370 6169 -1336 6345
rect -1274 6169 -1240 6345
rect -1160 6169 -1126 6345
rect -1064 6169 -1030 6345
rect -950 6169 -916 6345
rect -854 6169 -820 6345
rect -740 6169 -706 6345
rect -644 6169 -610 6345
rect -530 6169 -496 6345
rect -434 6169 -400 6345
rect -320 6169 -286 6345
rect -224 6169 -190 6345
rect -110 6169 -76 6345
rect -14 6169 20 6345
rect 100 6169 134 6345
rect 196 6169 230 6345
rect 310 6169 344 6345
rect 406 6169 440 6345
rect 520 6169 554 6345
rect 616 6169 650 6345
rect 730 6169 764 6345
rect 826 6169 860 6345
rect 940 6169 974 6345
rect 1036 6169 1070 6345
rect 1150 6169 1184 6345
rect 1246 6169 1280 6345
rect 1360 6169 1394 6345
rect 1456 6169 1490 6345
rect 1570 6169 1604 6345
rect 1666 6169 1700 6345
rect 1780 6169 1814 6345
rect 1876 6169 1910 6345
rect 1990 6169 2024 6345
rect 2086 6169 2120 6345
rect 2200 6169 2234 6345
rect 2296 6169 2330 6345
rect 2410 6169 2444 6345
rect 2506 6169 2540 6345
rect 2620 6169 2654 6345
rect 2716 6169 2750 6345
rect 2830 6169 2864 6345
rect 2926 6169 2960 6345
rect 3040 6169 3074 6345
rect 3136 6169 3170 6345
rect 3250 6169 3284 6345
rect 3346 6169 3380 6345
rect 3460 6169 3494 6345
rect 3556 6169 3590 6345
rect 3670 6169 3704 6345
rect 3766 6169 3800 6345
rect 3880 6169 3914 6345
rect 3976 6169 4010 6345
rect 4090 6169 4124 6345
rect 4186 6169 4220 6345
rect 4300 6169 4334 6345
rect 4396 6169 4430 6345
rect 4510 6169 4544 6345
rect 4606 6169 4640 6345
rect 4720 6169 4754 6345
rect 4816 6169 4850 6345
rect 4930 6169 4964 6345
rect 5026 6169 5060 6345
rect 5140 6169 5174 6345
rect 5236 6169 5270 6345
rect 5350 6169 5384 6345
rect 5446 6169 5480 6345
rect 5560 6169 5594 6345
rect 5656 6169 5690 6345
rect 5770 6169 5804 6345
rect 5866 6169 5900 6345
rect 5980 6169 6014 6345
rect 6076 6169 6110 6345
rect -2630 5729 -2596 5905
rect -2534 5729 -2500 5905
rect -2420 5729 -2386 5905
rect -2324 5729 -2290 5905
rect -2210 5729 -2176 5905
rect -2114 5729 -2080 5905
rect -2000 5729 -1966 5905
rect -1904 5729 -1870 5905
rect -1790 5729 -1756 5905
rect -1694 5729 -1660 5905
rect -1580 5729 -1546 5905
rect -1484 5729 -1450 5905
rect -1370 5729 -1336 5905
rect -1274 5729 -1240 5905
rect -1160 5729 -1126 5905
rect -1064 5729 -1030 5905
rect -950 5729 -916 5905
rect -854 5729 -820 5905
rect -740 5729 -706 5905
rect -644 5729 -610 5905
rect -530 5729 -496 5905
rect -434 5729 -400 5905
rect -320 5729 -286 5905
rect -224 5729 -190 5905
rect -110 5729 -76 5905
rect -14 5729 20 5905
rect 100 5729 134 5905
rect 196 5729 230 5905
rect 310 5729 344 5905
rect 406 5729 440 5905
rect 520 5729 554 5905
rect 616 5729 650 5905
rect 730 5729 764 5905
rect 826 5729 860 5905
rect 940 5729 974 5905
rect 1036 5729 1070 5905
rect 1150 5729 1184 5905
rect 1246 5729 1280 5905
rect 1360 5729 1394 5905
rect 1456 5729 1490 5905
rect 1570 5729 1604 5905
rect 1666 5729 1700 5905
rect 1780 5729 1814 5905
rect 1876 5729 1910 5905
rect 1990 5729 2024 5905
rect 2086 5729 2120 5905
rect 2200 5729 2234 5905
rect 2296 5729 2330 5905
rect 2410 5729 2444 5905
rect 2506 5729 2540 5905
rect 2620 5729 2654 5905
rect 2716 5729 2750 5905
rect 2830 5729 2864 5905
rect 2926 5729 2960 5905
rect 3040 5729 3074 5905
rect 3136 5729 3170 5905
rect 3250 5729 3284 5905
rect 3346 5729 3380 5905
rect 3460 5729 3494 5905
rect 3556 5729 3590 5905
rect 3670 5729 3704 5905
rect 3766 5729 3800 5905
rect 3880 5729 3914 5905
rect 3976 5729 4010 5905
rect 4090 5729 4124 5905
rect 4186 5729 4220 5905
rect 4300 5729 4334 5905
rect 4396 5729 4430 5905
rect 4510 5729 4544 5905
rect 4606 5729 4640 5905
rect 4720 5729 4754 5905
rect 4816 5729 4850 5905
rect 4930 5729 4964 5905
rect 5026 5729 5060 5905
rect 5140 5729 5174 5905
rect 5236 5729 5270 5905
rect 5350 5729 5384 5905
rect 5446 5729 5480 5905
rect 5560 5729 5594 5905
rect 5656 5729 5690 5905
rect 5770 5729 5804 5905
rect 5866 5729 5900 5905
rect 5980 5729 6014 5905
rect 6076 5729 6110 5905
rect -2630 5289 -2596 5465
rect -2534 5289 -2500 5465
rect -2420 5289 -2386 5465
rect -2324 5289 -2290 5465
rect -2210 5289 -2176 5465
rect -2114 5289 -2080 5465
rect -2000 5289 -1966 5465
rect -1904 5289 -1870 5465
rect -1790 5289 -1756 5465
rect -1694 5289 -1660 5465
rect -1580 5289 -1546 5465
rect -1484 5289 -1450 5465
rect -1370 5289 -1336 5465
rect -1274 5289 -1240 5465
rect -1160 5289 -1126 5465
rect -1064 5289 -1030 5465
rect -950 5289 -916 5465
rect -854 5289 -820 5465
rect -740 5289 -706 5465
rect -644 5289 -610 5465
rect -530 5289 -496 5465
rect -434 5289 -400 5465
rect -320 5289 -286 5465
rect -224 5289 -190 5465
rect -110 5289 -76 5465
rect -14 5289 20 5465
rect 100 5289 134 5465
rect 196 5289 230 5465
rect 310 5289 344 5465
rect 406 5289 440 5465
rect 520 5289 554 5465
rect 616 5289 650 5465
rect 730 5289 764 5465
rect 826 5289 860 5465
rect 940 5289 974 5465
rect 1036 5289 1070 5465
rect 1150 5289 1184 5465
rect 1246 5289 1280 5465
rect 1360 5289 1394 5465
rect 1456 5289 1490 5465
rect 1570 5289 1604 5465
rect 1666 5289 1700 5465
rect 1780 5289 1814 5465
rect 1876 5289 1910 5465
rect 1990 5289 2024 5465
rect 2086 5289 2120 5465
rect 2200 5289 2234 5465
rect 2296 5289 2330 5465
rect 2410 5289 2444 5465
rect 2506 5289 2540 5465
rect 2620 5289 2654 5465
rect 2716 5289 2750 5465
rect 2830 5289 2864 5465
rect 2926 5289 2960 5465
rect 3040 5289 3074 5465
rect 3136 5289 3170 5465
rect 3250 5289 3284 5465
rect 3346 5289 3380 5465
rect 3460 5289 3494 5465
rect 3556 5289 3590 5465
rect 3670 5289 3704 5465
rect 3766 5289 3800 5465
rect 3880 5289 3914 5465
rect 3976 5289 4010 5465
rect 4090 5289 4124 5465
rect 4186 5289 4220 5465
rect 4300 5289 4334 5465
rect 4396 5289 4430 5465
rect 4510 5289 4544 5465
rect 4606 5289 4640 5465
rect 4720 5289 4754 5465
rect 4816 5289 4850 5465
rect 4930 5289 4964 5465
rect 5026 5289 5060 5465
rect 5140 5289 5174 5465
rect 5236 5289 5270 5465
rect 5350 5289 5384 5465
rect 5446 5289 5480 5465
rect 5560 5289 5594 5465
rect 5656 5289 5690 5465
rect 5770 5289 5804 5465
rect 5866 5289 5900 5465
rect 5980 5289 6014 5465
rect 6076 5289 6110 5465
rect -2630 4849 -2596 5025
rect -2534 4849 -2500 5025
rect -2420 4849 -2386 5025
rect -2324 4849 -2290 5025
rect -2210 4849 -2176 5025
rect -2114 4849 -2080 5025
rect -2000 4849 -1966 5025
rect -1904 4849 -1870 5025
rect -1790 4849 -1756 5025
rect -1694 4849 -1660 5025
rect -1580 4849 -1546 5025
rect -1484 4849 -1450 5025
rect -1370 4849 -1336 5025
rect -1274 4849 -1240 5025
rect -1160 4849 -1126 5025
rect -1064 4849 -1030 5025
rect -950 4849 -916 5025
rect -854 4849 -820 5025
rect -740 4849 -706 5025
rect -644 4849 -610 5025
rect -530 4849 -496 5025
rect -434 4849 -400 5025
rect -320 4849 -286 5025
rect -224 4849 -190 5025
rect -110 4849 -76 5025
rect -14 4849 20 5025
rect 100 4849 134 5025
rect 196 4849 230 5025
rect 310 4849 344 5025
rect 406 4849 440 5025
rect 520 4849 554 5025
rect 616 4849 650 5025
rect 730 4849 764 5025
rect 826 4849 860 5025
rect 940 4849 974 5025
rect 1036 4849 1070 5025
rect 1150 4849 1184 5025
rect 1246 4849 1280 5025
rect 1360 4849 1394 5025
rect 1456 4849 1490 5025
rect 1570 4849 1604 5025
rect 1666 4849 1700 5025
rect 1780 4849 1814 5025
rect 1876 4849 1910 5025
rect 1990 4849 2024 5025
rect 2086 4849 2120 5025
rect 2200 4849 2234 5025
rect 2296 4849 2330 5025
rect 2410 4849 2444 5025
rect 2506 4849 2540 5025
rect 2620 4849 2654 5025
rect 2716 4849 2750 5025
rect 2830 4849 2864 5025
rect 2926 4849 2960 5025
rect 3040 4849 3074 5025
rect 3136 4849 3170 5025
rect 3250 4849 3284 5025
rect 3346 4849 3380 5025
rect 3460 4849 3494 5025
rect 3556 4849 3590 5025
rect 3670 4849 3704 5025
rect 3766 4849 3800 5025
rect 3880 4849 3914 5025
rect 3976 4849 4010 5025
rect 4090 4849 4124 5025
rect 4186 4849 4220 5025
rect 4300 4849 4334 5025
rect 4396 4849 4430 5025
rect 4510 4849 4544 5025
rect 4606 4849 4640 5025
rect 4720 4849 4754 5025
rect 4816 4849 4850 5025
rect 4930 4849 4964 5025
rect 5026 4849 5060 5025
rect 5140 4849 5174 5025
rect 5236 4849 5270 5025
rect 5350 4849 5384 5025
rect 5446 4849 5480 5025
rect 5560 4849 5594 5025
rect 5656 4849 5690 5025
rect 5770 4849 5804 5025
rect 5866 4849 5900 5025
rect 5980 4849 6014 5025
rect 6076 4849 6110 5025
rect -2630 3914 -2596 4090
rect -2534 3914 -2500 4090
rect -2420 3914 -2386 4090
rect -2324 3914 -2290 4090
rect -2210 3914 -2176 4090
rect -2114 3914 -2080 4090
rect -2000 3914 -1966 4090
rect -1904 3914 -1870 4090
rect -1790 3914 -1756 4090
rect -1694 3914 -1660 4090
rect -1580 3914 -1546 4090
rect -1484 3914 -1450 4090
rect -1370 3914 -1336 4090
rect -1274 3914 -1240 4090
rect -1160 3914 -1126 4090
rect -1064 3914 -1030 4090
rect -950 3914 -916 4090
rect -854 3914 -820 4090
rect -740 3914 -706 4090
rect -644 3914 -610 4090
rect -530 3914 -496 4090
rect -434 3914 -400 4090
rect -320 3914 -286 4090
rect -224 3914 -190 4090
rect -110 3914 -76 4090
rect -14 3914 20 4090
rect 100 3914 134 4090
rect 196 3914 230 4090
rect 310 3914 344 4090
rect 406 3914 440 4090
rect 520 3914 554 4090
rect 616 3914 650 4090
rect 730 3914 764 4090
rect 826 3914 860 4090
rect 940 3914 974 4090
rect 1036 3914 1070 4090
rect 1150 3914 1184 4090
rect 1246 3914 1280 4090
rect 1360 3914 1394 4090
rect 1456 3914 1490 4090
rect 1570 3914 1604 4090
rect 1666 3914 1700 4090
rect 1780 3914 1814 4090
rect 1876 3914 1910 4090
rect 1990 3914 2024 4090
rect 2086 3914 2120 4090
rect 2200 3914 2234 4090
rect 2296 3914 2330 4090
rect 2410 3914 2444 4090
rect 2506 3914 2540 4090
rect 2620 3914 2654 4090
rect 2716 3914 2750 4090
rect 2830 3914 2864 4090
rect 2926 3914 2960 4090
rect 3040 3914 3074 4090
rect 3136 3914 3170 4090
rect 3250 3914 3284 4090
rect 3346 3914 3380 4090
rect 3460 3914 3494 4090
rect 3556 3914 3590 4090
rect 3670 3914 3704 4090
rect 3766 3914 3800 4090
rect 3880 3914 3914 4090
rect 3976 3914 4010 4090
rect 4090 3914 4124 4090
rect 4186 3914 4220 4090
rect 4300 3914 4334 4090
rect 4396 3914 4430 4090
rect 4510 3914 4544 4090
rect 4606 3914 4640 4090
rect 4720 3914 4754 4090
rect 4816 3914 4850 4090
rect 4930 3914 4964 4090
rect 5026 3914 5060 4090
rect 5140 3914 5174 4090
rect 5236 3914 5270 4090
rect 5350 3914 5384 4090
rect 5446 3914 5480 4090
rect 5560 3914 5594 4090
rect 5656 3914 5690 4090
rect 5770 3914 5804 4090
rect 5866 3914 5900 4090
rect 5980 3914 6014 4090
rect 6076 3914 6110 4090
rect -2630 3474 -2596 3650
rect -2534 3474 -2500 3650
rect -2420 3474 -2386 3650
rect -2324 3474 -2290 3650
rect -2210 3474 -2176 3650
rect -2114 3474 -2080 3650
rect -2000 3474 -1966 3650
rect -1904 3474 -1870 3650
rect -1790 3474 -1756 3650
rect -1694 3474 -1660 3650
rect -1580 3474 -1546 3650
rect -1484 3474 -1450 3650
rect -1370 3474 -1336 3650
rect -1274 3474 -1240 3650
rect -1160 3474 -1126 3650
rect -1064 3474 -1030 3650
rect -950 3474 -916 3650
rect -854 3474 -820 3650
rect -740 3474 -706 3650
rect -644 3474 -610 3650
rect -530 3474 -496 3650
rect -434 3474 -400 3650
rect -320 3474 -286 3650
rect -224 3474 -190 3650
rect -110 3474 -76 3650
rect -14 3474 20 3650
rect 100 3474 134 3650
rect 196 3474 230 3650
rect 310 3474 344 3650
rect 406 3474 440 3650
rect 520 3474 554 3650
rect 616 3474 650 3650
rect 730 3474 764 3650
rect 826 3474 860 3650
rect 940 3474 974 3650
rect 1036 3474 1070 3650
rect 1150 3474 1184 3650
rect 1246 3474 1280 3650
rect 1360 3474 1394 3650
rect 1456 3474 1490 3650
rect 1570 3474 1604 3650
rect 1666 3474 1700 3650
rect 1780 3474 1814 3650
rect 1876 3474 1910 3650
rect 1990 3474 2024 3650
rect 2086 3474 2120 3650
rect 2200 3474 2234 3650
rect 2296 3474 2330 3650
rect 2410 3474 2444 3650
rect 2506 3474 2540 3650
rect 2620 3474 2654 3650
rect 2716 3474 2750 3650
rect 2830 3474 2864 3650
rect 2926 3474 2960 3650
rect 3040 3474 3074 3650
rect 3136 3474 3170 3650
rect 3250 3474 3284 3650
rect 3346 3474 3380 3650
rect 3460 3474 3494 3650
rect 3556 3474 3590 3650
rect 3670 3474 3704 3650
rect 3766 3474 3800 3650
rect 3880 3474 3914 3650
rect 3976 3474 4010 3650
rect 4090 3474 4124 3650
rect 4186 3474 4220 3650
rect 4300 3474 4334 3650
rect 4396 3474 4430 3650
rect 4510 3474 4544 3650
rect 4606 3474 4640 3650
rect 4720 3474 4754 3650
rect 4816 3474 4850 3650
rect 4930 3474 4964 3650
rect 5026 3474 5060 3650
rect 5140 3474 5174 3650
rect 5236 3474 5270 3650
rect 5350 3474 5384 3650
rect 5446 3474 5480 3650
rect 5560 3474 5594 3650
rect 5656 3474 5690 3650
rect 5770 3474 5804 3650
rect 5866 3474 5900 3650
rect 5980 3474 6014 3650
rect 6076 3474 6110 3650
rect -2630 3034 -2596 3210
rect -2534 3034 -2500 3210
rect -2420 3034 -2386 3210
rect -2324 3034 -2290 3210
rect -2210 3034 -2176 3210
rect -2114 3034 -2080 3210
rect -2000 3034 -1966 3210
rect -1904 3034 -1870 3210
rect -1790 3034 -1756 3210
rect -1694 3034 -1660 3210
rect -1580 3034 -1546 3210
rect -1484 3034 -1450 3210
rect -1370 3034 -1336 3210
rect -1274 3034 -1240 3210
rect -1160 3034 -1126 3210
rect -1064 3034 -1030 3210
rect -950 3034 -916 3210
rect -854 3034 -820 3210
rect -740 3034 -706 3210
rect -644 3034 -610 3210
rect -530 3034 -496 3210
rect -434 3034 -400 3210
rect -320 3034 -286 3210
rect -224 3034 -190 3210
rect -110 3034 -76 3210
rect -14 3034 20 3210
rect 100 3034 134 3210
rect 196 3034 230 3210
rect 310 3034 344 3210
rect 406 3034 440 3210
rect 520 3034 554 3210
rect 616 3034 650 3210
rect 730 3034 764 3210
rect 826 3034 860 3210
rect 940 3034 974 3210
rect 1036 3034 1070 3210
rect 1150 3034 1184 3210
rect 1246 3034 1280 3210
rect 1360 3034 1394 3210
rect 1456 3034 1490 3210
rect 1570 3034 1604 3210
rect 1666 3034 1700 3210
rect 1780 3034 1814 3210
rect 1876 3034 1910 3210
rect 1990 3034 2024 3210
rect 2086 3034 2120 3210
rect 2200 3034 2234 3210
rect 2296 3034 2330 3210
rect 2410 3034 2444 3210
rect 2506 3034 2540 3210
rect 2620 3034 2654 3210
rect 2716 3034 2750 3210
rect 2830 3034 2864 3210
rect 2926 3034 2960 3210
rect 3040 3034 3074 3210
rect 3136 3034 3170 3210
rect 3250 3034 3284 3210
rect 3346 3034 3380 3210
rect 3460 3034 3494 3210
rect 3556 3034 3590 3210
rect 3670 3034 3704 3210
rect 3766 3034 3800 3210
rect 3880 3034 3914 3210
rect 3976 3034 4010 3210
rect 4090 3034 4124 3210
rect 4186 3034 4220 3210
rect 4300 3034 4334 3210
rect 4396 3034 4430 3210
rect 4510 3034 4544 3210
rect 4606 3034 4640 3210
rect 4720 3034 4754 3210
rect 4816 3034 4850 3210
rect 4930 3034 4964 3210
rect 5026 3034 5060 3210
rect 5140 3034 5174 3210
rect 5236 3034 5270 3210
rect 5350 3034 5384 3210
rect 5446 3034 5480 3210
rect 5560 3034 5594 3210
rect 5656 3034 5690 3210
rect 5770 3034 5804 3210
rect 5866 3034 5900 3210
rect 5980 3034 6014 3210
rect 6076 3034 6110 3210
rect -2630 2594 -2596 2770
rect -2534 2594 -2500 2770
rect -2420 2594 -2386 2770
rect -2324 2594 -2290 2770
rect -2210 2594 -2176 2770
rect -2114 2594 -2080 2770
rect -2000 2594 -1966 2770
rect -1904 2594 -1870 2770
rect -1790 2594 -1756 2770
rect -1694 2594 -1660 2770
rect -1580 2594 -1546 2770
rect -1484 2594 -1450 2770
rect -1370 2594 -1336 2770
rect -1274 2594 -1240 2770
rect -1160 2594 -1126 2770
rect -1064 2594 -1030 2770
rect -950 2594 -916 2770
rect -854 2594 -820 2770
rect -740 2594 -706 2770
rect -644 2594 -610 2770
rect -530 2594 -496 2770
rect -434 2594 -400 2770
rect -320 2594 -286 2770
rect -224 2594 -190 2770
rect -110 2594 -76 2770
rect -14 2594 20 2770
rect 100 2594 134 2770
rect 196 2594 230 2770
rect 310 2594 344 2770
rect 406 2594 440 2770
rect 520 2594 554 2770
rect 616 2594 650 2770
rect 730 2594 764 2770
rect 826 2594 860 2770
rect 940 2594 974 2770
rect 1036 2594 1070 2770
rect 1150 2594 1184 2770
rect 1246 2594 1280 2770
rect 1360 2594 1394 2770
rect 1456 2594 1490 2770
rect 1570 2594 1604 2770
rect 1666 2594 1700 2770
rect 1780 2594 1814 2770
rect 1876 2594 1910 2770
rect 1990 2594 2024 2770
rect 2086 2594 2120 2770
rect 2200 2594 2234 2770
rect 2296 2594 2330 2770
rect 2410 2594 2444 2770
rect 2506 2594 2540 2770
rect 2620 2594 2654 2770
rect 2716 2594 2750 2770
rect 2830 2594 2864 2770
rect 2926 2594 2960 2770
rect 3040 2594 3074 2770
rect 3136 2594 3170 2770
rect 3250 2594 3284 2770
rect 3346 2594 3380 2770
rect 3460 2594 3494 2770
rect 3556 2594 3590 2770
rect 3670 2594 3704 2770
rect 3766 2594 3800 2770
rect 3880 2594 3914 2770
rect 3976 2594 4010 2770
rect 4090 2594 4124 2770
rect 4186 2594 4220 2770
rect 4300 2594 4334 2770
rect 4396 2594 4430 2770
rect 4510 2594 4544 2770
rect 4606 2594 4640 2770
rect 4720 2594 4754 2770
rect 4816 2594 4850 2770
rect 4930 2594 4964 2770
rect 5026 2594 5060 2770
rect 5140 2594 5174 2770
rect 5236 2594 5270 2770
rect 5350 2594 5384 2770
rect 5446 2594 5480 2770
rect 5560 2594 5594 2770
rect 5656 2594 5690 2770
rect 5770 2594 5804 2770
rect 5866 2594 5900 2770
rect 5980 2594 6014 2770
rect 6076 2594 6110 2770
rect -2630 2154 -2596 2330
rect -2534 2154 -2500 2330
rect -2420 2154 -2386 2330
rect -2324 2154 -2290 2330
rect -2210 2154 -2176 2330
rect -2114 2154 -2080 2330
rect -2000 2154 -1966 2330
rect -1904 2154 -1870 2330
rect -1790 2154 -1756 2330
rect -1694 2154 -1660 2330
rect -1580 2154 -1546 2330
rect -1484 2154 -1450 2330
rect -1370 2154 -1336 2330
rect -1274 2154 -1240 2330
rect -1160 2154 -1126 2330
rect -1064 2154 -1030 2330
rect -950 2154 -916 2330
rect -854 2154 -820 2330
rect -740 2154 -706 2330
rect -644 2154 -610 2330
rect -530 2154 -496 2330
rect -434 2154 -400 2330
rect -320 2154 -286 2330
rect -224 2154 -190 2330
rect -110 2154 -76 2330
rect -14 2154 20 2330
rect 100 2154 134 2330
rect 196 2154 230 2330
rect 310 2154 344 2330
rect 406 2154 440 2330
rect 520 2154 554 2330
rect 616 2154 650 2330
rect 730 2154 764 2330
rect 826 2154 860 2330
rect 940 2154 974 2330
rect 1036 2154 1070 2330
rect 1150 2154 1184 2330
rect 1246 2154 1280 2330
rect 1360 2154 1394 2330
rect 1456 2154 1490 2330
rect 1570 2154 1604 2330
rect 1666 2154 1700 2330
rect 1780 2154 1814 2330
rect 1876 2154 1910 2330
rect 1990 2154 2024 2330
rect 2086 2154 2120 2330
rect 2200 2154 2234 2330
rect 2296 2154 2330 2330
rect 2410 2154 2444 2330
rect 2506 2154 2540 2330
rect 2620 2154 2654 2330
rect 2716 2154 2750 2330
rect 2830 2154 2864 2330
rect 2926 2154 2960 2330
rect 3040 2154 3074 2330
rect 3136 2154 3170 2330
rect 3250 2154 3284 2330
rect 3346 2154 3380 2330
rect 3460 2154 3494 2330
rect 3556 2154 3590 2330
rect 3670 2154 3704 2330
rect 3766 2154 3800 2330
rect 3880 2154 3914 2330
rect 3976 2154 4010 2330
rect 4090 2154 4124 2330
rect 4186 2154 4220 2330
rect 4300 2154 4334 2330
rect 4396 2154 4430 2330
rect 4510 2154 4544 2330
rect 4606 2154 4640 2330
rect 4720 2154 4754 2330
rect 4816 2154 4850 2330
rect 4930 2154 4964 2330
rect 5026 2154 5060 2330
rect 5140 2154 5174 2330
rect 5236 2154 5270 2330
rect 5350 2154 5384 2330
rect 5446 2154 5480 2330
rect 5560 2154 5594 2330
rect 5656 2154 5690 2330
rect 5770 2154 5804 2330
rect 5866 2154 5900 2330
rect 5980 2154 6014 2330
rect 6076 2154 6110 2330
rect -2630 1714 -2596 1890
rect -2534 1714 -2500 1890
rect -2420 1714 -2386 1890
rect -2324 1714 -2290 1890
rect -2210 1714 -2176 1890
rect -2114 1714 -2080 1890
rect -2000 1714 -1966 1890
rect -1904 1714 -1870 1890
rect -1790 1714 -1756 1890
rect -1694 1714 -1660 1890
rect -1580 1714 -1546 1890
rect -1484 1714 -1450 1890
rect -1370 1714 -1336 1890
rect -1274 1714 -1240 1890
rect -1160 1714 -1126 1890
rect -1064 1714 -1030 1890
rect -950 1714 -916 1890
rect -854 1714 -820 1890
rect -740 1714 -706 1890
rect -644 1714 -610 1890
rect -530 1714 -496 1890
rect -434 1714 -400 1890
rect -320 1714 -286 1890
rect -224 1714 -190 1890
rect -110 1714 -76 1890
rect -14 1714 20 1890
rect 100 1714 134 1890
rect 196 1714 230 1890
rect 310 1714 344 1890
rect 406 1714 440 1890
rect 520 1714 554 1890
rect 616 1714 650 1890
rect 730 1714 764 1890
rect 826 1714 860 1890
rect 940 1714 974 1890
rect 1036 1714 1070 1890
rect 1150 1714 1184 1890
rect 1246 1714 1280 1890
rect 1360 1714 1394 1890
rect 1456 1714 1490 1890
rect 1570 1714 1604 1890
rect 1666 1714 1700 1890
rect 1780 1714 1814 1890
rect 1876 1714 1910 1890
rect 1990 1714 2024 1890
rect 2086 1714 2120 1890
rect 2200 1714 2234 1890
rect 2296 1714 2330 1890
rect 2410 1714 2444 1890
rect 2506 1714 2540 1890
rect 2620 1714 2654 1890
rect 2716 1714 2750 1890
rect 2830 1714 2864 1890
rect 2926 1714 2960 1890
rect 3040 1714 3074 1890
rect 3136 1714 3170 1890
rect 3250 1714 3284 1890
rect 3346 1714 3380 1890
rect 3460 1714 3494 1890
rect 3556 1714 3590 1890
rect 3670 1714 3704 1890
rect 3766 1714 3800 1890
rect 3880 1714 3914 1890
rect 3976 1714 4010 1890
rect 4090 1714 4124 1890
rect 4186 1714 4220 1890
rect 4300 1714 4334 1890
rect 4396 1714 4430 1890
rect 4510 1714 4544 1890
rect 4606 1714 4640 1890
rect 4720 1714 4754 1890
rect 4816 1714 4850 1890
rect 4930 1714 4964 1890
rect 5026 1714 5060 1890
rect 5140 1714 5174 1890
rect 5236 1714 5270 1890
rect 5350 1714 5384 1890
rect 5446 1714 5480 1890
rect 5560 1714 5594 1890
rect 5656 1714 5690 1890
rect 5770 1714 5804 1890
rect 5866 1714 5900 1890
rect 5980 1714 6014 1890
rect 6076 1714 6110 1890
rect -2630 1274 -2596 1450
rect -2534 1274 -2500 1450
rect -2420 1274 -2386 1450
rect -2324 1274 -2290 1450
rect -2210 1274 -2176 1450
rect -2114 1274 -2080 1450
rect -2000 1274 -1966 1450
rect -1904 1274 -1870 1450
rect -1790 1274 -1756 1450
rect -1694 1274 -1660 1450
rect -1580 1274 -1546 1450
rect -1484 1274 -1450 1450
rect -1370 1274 -1336 1450
rect -1274 1274 -1240 1450
rect -1160 1274 -1126 1450
rect -1064 1274 -1030 1450
rect -950 1274 -916 1450
rect -854 1274 -820 1450
rect -740 1274 -706 1450
rect -644 1274 -610 1450
rect -530 1274 -496 1450
rect -434 1274 -400 1450
rect -320 1274 -286 1450
rect -224 1274 -190 1450
rect -110 1274 -76 1450
rect -14 1274 20 1450
rect 100 1274 134 1450
rect 196 1274 230 1450
rect 310 1274 344 1450
rect 406 1274 440 1450
rect 520 1274 554 1450
rect 616 1274 650 1450
rect 730 1274 764 1450
rect 826 1274 860 1450
rect 940 1274 974 1450
rect 1036 1274 1070 1450
rect 1150 1274 1184 1450
rect 1246 1274 1280 1450
rect 1360 1274 1394 1450
rect 1456 1274 1490 1450
rect 1570 1274 1604 1450
rect 1666 1274 1700 1450
rect 1780 1274 1814 1450
rect 1876 1274 1910 1450
rect 1990 1274 2024 1450
rect 2086 1274 2120 1450
rect 2200 1274 2234 1450
rect 2296 1274 2330 1450
rect 2410 1274 2444 1450
rect 2506 1274 2540 1450
rect 2620 1274 2654 1450
rect 2716 1274 2750 1450
rect 2830 1274 2864 1450
rect 2926 1274 2960 1450
rect 3040 1274 3074 1450
rect 3136 1274 3170 1450
rect 3250 1274 3284 1450
rect 3346 1274 3380 1450
rect 3460 1274 3494 1450
rect 3556 1274 3590 1450
rect 3670 1274 3704 1450
rect 3766 1274 3800 1450
rect 3880 1274 3914 1450
rect 3976 1274 4010 1450
rect 4090 1274 4124 1450
rect 4186 1274 4220 1450
rect 4300 1274 4334 1450
rect 4396 1274 4430 1450
rect 4510 1274 4544 1450
rect 4606 1274 4640 1450
rect 4720 1274 4754 1450
rect 4816 1274 4850 1450
rect 4930 1274 4964 1450
rect 5026 1274 5060 1450
rect 5140 1274 5174 1450
rect 5236 1274 5270 1450
rect 5350 1274 5384 1450
rect 5446 1274 5480 1450
rect 5560 1274 5594 1450
rect 5656 1274 5690 1450
rect 5770 1274 5804 1450
rect 5866 1274 5900 1450
rect 5980 1274 6014 1450
rect 6076 1274 6110 1450
rect -2630 834 -2596 1010
rect -2534 834 -2500 1010
rect -2420 834 -2386 1010
rect -2324 834 -2290 1010
rect -2210 834 -2176 1010
rect -2114 834 -2080 1010
rect -2000 834 -1966 1010
rect -1904 834 -1870 1010
rect -1790 834 -1756 1010
rect -1694 834 -1660 1010
rect -1580 834 -1546 1010
rect -1484 834 -1450 1010
rect -1370 834 -1336 1010
rect -1274 834 -1240 1010
rect -1160 834 -1126 1010
rect -1064 834 -1030 1010
rect -950 834 -916 1010
rect -854 834 -820 1010
rect -740 834 -706 1010
rect -644 834 -610 1010
rect -530 834 -496 1010
rect -434 834 -400 1010
rect -320 834 -286 1010
rect -224 834 -190 1010
rect -110 834 -76 1010
rect -14 834 20 1010
rect 100 834 134 1010
rect 196 834 230 1010
rect 310 834 344 1010
rect 406 834 440 1010
rect 520 834 554 1010
rect 616 834 650 1010
rect 730 834 764 1010
rect 826 834 860 1010
rect 940 834 974 1010
rect 1036 834 1070 1010
rect 1150 834 1184 1010
rect 1246 834 1280 1010
rect 1360 834 1394 1010
rect 1456 834 1490 1010
rect 1570 834 1604 1010
rect 1666 834 1700 1010
rect 1780 834 1814 1010
rect 1876 834 1910 1010
rect 1990 834 2024 1010
rect 2086 834 2120 1010
rect 2200 834 2234 1010
rect 2296 834 2330 1010
rect 2410 834 2444 1010
rect 2506 834 2540 1010
rect 2620 834 2654 1010
rect 2716 834 2750 1010
rect 2830 834 2864 1010
rect 2926 834 2960 1010
rect 3040 834 3074 1010
rect 3136 834 3170 1010
rect 3250 834 3284 1010
rect 3346 834 3380 1010
rect 3460 834 3494 1010
rect 3556 834 3590 1010
rect 3670 834 3704 1010
rect 3766 834 3800 1010
rect 3880 834 3914 1010
rect 3976 834 4010 1010
rect 4090 834 4124 1010
rect 4186 834 4220 1010
rect 4300 834 4334 1010
rect 4396 834 4430 1010
rect 4510 834 4544 1010
rect 4606 834 4640 1010
rect 4720 834 4754 1010
rect 4816 834 4850 1010
rect 4930 834 4964 1010
rect 5026 834 5060 1010
rect 5140 834 5174 1010
rect 5236 834 5270 1010
rect 5350 834 5384 1010
rect 5446 834 5480 1010
rect 5560 834 5594 1010
rect 5656 834 5690 1010
rect 5770 834 5804 1010
rect 5866 834 5900 1010
rect 5980 834 6014 1010
rect 6076 834 6110 1010
rect 90 30 124 206
rect 186 30 220 206
rect 282 30 316 206
rect 378 30 412 206
rect 474 30 508 206
rect 570 30 604 206
rect 666 30 700 206
rect 762 30 796 206
rect 858 30 892 206
rect 954 30 988 206
rect 1050 30 1084 206
rect 1146 30 1180 206
rect 1242 30 1276 206
rect 1338 30 1372 206
rect 1434 30 1468 206
rect 1530 30 1564 206
rect 1626 30 1660 206
rect 1722 30 1756 206
rect 1818 30 1852 206
rect 1914 30 1948 206
rect 2010 30 2044 206
rect 2106 30 2140 206
rect 2202 30 2236 206
rect 2298 30 2332 206
rect 2394 30 2428 206
rect 2490 30 2524 206
rect 2586 30 2620 206
rect 2682 30 2716 206
rect 2778 30 2812 206
rect 2874 30 2908 206
rect 2970 30 3004 206
rect 3066 30 3100 206
rect 3162 30 3196 206
rect 3258 30 3292 206
rect 3354 30 3388 206
<< pdiffc >>
rect 1531 10564 1565 10598
rect 1633 10564 1667 10598
rect 1785 10564 1819 10598
rect 1887 10564 1921 10598
rect 1531 9564 1565 9598
rect 1633 9564 1667 9598
rect 1785 9564 1819 9598
rect 1887 9564 1921 9598
rect 1497 9368 1531 9402
rect 1565 9368 1599 9402
rect 1633 9368 1667 9402
rect 1785 9368 1819 9402
rect 1853 9368 1887 9402
rect 1921 9368 1955 9402
rect 1497 9284 1531 9318
rect 1565 9284 1599 9318
rect 1633 9284 1667 9318
rect 1785 9284 1819 9318
rect 1853 9284 1887 9318
rect 1921 9284 1955 9318
rect 1565 9200 1599 9234
rect 1633 9200 1667 9234
rect 1785 9200 1819 9234
rect 1853 9200 1887 9234
rect 1497 9116 1531 9150
rect 1565 9116 1599 9150
rect 1633 9116 1667 9150
rect 1785 9116 1819 9150
rect 1853 9116 1887 9150
rect 1921 9116 1955 9150
rect 1565 9032 1599 9066
rect 1633 9032 1667 9066
rect 1785 9032 1819 9066
rect 1853 9032 1887 9066
rect 1497 8948 1531 8982
rect 1565 8948 1599 8982
rect 1633 8948 1667 8982
rect 1785 8948 1819 8982
rect 1853 8948 1887 8982
rect 1921 8948 1955 8982
rect 1565 8864 1599 8898
rect 1633 8864 1667 8898
rect 1785 8864 1819 8898
rect 1853 8864 1887 8898
rect 1497 8780 1531 8814
rect 1565 8780 1599 8814
rect 1633 8780 1667 8814
rect 1785 8780 1819 8814
rect 1853 8780 1887 8814
rect 1921 8780 1955 8814
rect 1565 8696 1599 8730
rect 1633 8696 1667 8730
rect 1785 8696 1819 8730
rect 1853 8696 1887 8730
rect 1497 8539 1531 8573
rect 1565 8539 1599 8573
rect 1633 8539 1667 8573
rect 1785 8539 1819 8573
rect 1853 8539 1887 8573
rect 1921 8539 1955 8573
rect 1528 8455 1562 8489
rect 1609 8455 1643 8489
rect 1809 8455 1843 8489
rect 1890 8455 1924 8489
rect 1557 8369 1591 8403
rect 1625 8369 1659 8403
rect 1793 8369 1827 8403
rect 1861 8369 1895 8403
rect 1557 8276 1591 8310
rect 1625 8276 1659 8310
rect 1793 8276 1827 8310
rect 1861 8276 1895 8310
rect -3557 7876 -3381 7910
rect -3557 7780 -3381 7814
rect -3557 7684 -3381 7718
rect -3557 7588 -3381 7622
rect -3557 7492 -3381 7526
rect -3557 7396 -3381 7430
rect -3557 7300 -3381 7334
rect -3557 7204 -3381 7238
rect -3557 7108 -3381 7142
rect -3557 7012 -3381 7046
rect -3557 6916 -3381 6950
rect -3557 6820 -3381 6854
rect -3557 6724 -3381 6758
rect -3557 6628 -3381 6662
rect -3557 6532 -3381 6566
rect -3557 6436 -3381 6470
rect -3557 6340 -3381 6374
rect -3557 6244 -3381 6278
rect -3557 6148 -3381 6182
rect -2644 7652 -2610 7828
rect -2548 7652 -2514 7828
rect -2434 7652 -2400 7828
rect -2338 7652 -2304 7828
rect -2224 7652 -2190 7828
rect -2128 7652 -2094 7828
rect -2014 7652 -1980 7828
rect -1918 7652 -1884 7828
rect -1804 7652 -1770 7828
rect -1708 7652 -1674 7828
rect -1594 7652 -1560 7828
rect -1498 7652 -1464 7828
rect -1384 7652 -1350 7828
rect -1288 7652 -1254 7828
rect -1174 7652 -1140 7828
rect -1078 7652 -1044 7828
rect -964 7652 -930 7828
rect -868 7652 -834 7828
rect -754 7652 -720 7828
rect -658 7652 -624 7828
rect -544 7652 -510 7828
rect -448 7652 -414 7828
rect -334 7652 -300 7828
rect -238 7652 -204 7828
rect -124 7652 -90 7828
rect -28 7652 6 7828
rect 86 7652 120 7828
rect 182 7652 216 7828
rect 296 7652 330 7828
rect 392 7652 426 7828
rect 506 7652 540 7828
rect 602 7652 636 7828
rect 716 7652 750 7828
rect 812 7652 846 7828
rect 926 7652 960 7828
rect 1022 7652 1056 7828
rect 1136 7652 1170 7828
rect 1232 7652 1266 7828
rect 1346 7652 1380 7828
rect 1442 7652 1476 7828
rect 1556 7652 1590 7828
rect 1652 7652 1686 7828
rect 1766 7652 1800 7828
rect 1862 7652 1896 7828
rect 1976 7652 2010 7828
rect 2072 7652 2106 7828
rect 2186 7652 2220 7828
rect 2282 7652 2316 7828
rect 2396 7652 2430 7828
rect 2492 7652 2526 7828
rect 2606 7652 2640 7828
rect 2702 7652 2736 7828
rect 2816 7652 2850 7828
rect 2912 7652 2946 7828
rect 3026 7652 3060 7828
rect 3122 7652 3156 7828
rect 3236 7652 3270 7828
rect 3332 7652 3366 7828
rect 3446 7652 3480 7828
rect 3542 7652 3576 7828
rect 3656 7652 3690 7828
rect 3752 7652 3786 7828
rect 3866 7652 3900 7828
rect 3962 7652 3996 7828
rect 4076 7652 4110 7828
rect 4172 7652 4206 7828
rect 4286 7652 4320 7828
rect 4382 7652 4416 7828
rect 4496 7652 4530 7828
rect 4592 7652 4626 7828
rect 4706 7652 4740 7828
rect 4802 7652 4836 7828
rect 4916 7652 4950 7828
rect 5012 7652 5046 7828
rect 5126 7652 5160 7828
rect 5222 7652 5256 7828
rect 5336 7652 5370 7828
rect 5432 7652 5466 7828
rect 5546 7652 5580 7828
rect 5642 7652 5676 7828
rect 5756 7652 5790 7828
rect 5852 7652 5886 7828
rect 5966 7652 6000 7828
rect 6062 7652 6096 7828
rect -2642 7119 -2608 7295
rect -2546 7119 -2512 7295
rect -2432 7119 -2398 7295
rect -2336 7119 -2302 7295
rect -2222 7119 -2188 7295
rect -2126 7119 -2092 7295
rect -2012 7119 -1978 7295
rect -1916 7119 -1882 7295
rect -1802 7119 -1768 7295
rect -1706 7119 -1672 7295
rect -1592 7119 -1558 7295
rect -1496 7119 -1462 7295
rect -1382 7119 -1348 7295
rect -1286 7119 -1252 7295
rect -1172 7119 -1138 7295
rect -1076 7119 -1042 7295
rect -962 7119 -928 7295
rect -866 7119 -832 7295
rect -752 7119 -718 7295
rect -656 7119 -622 7295
rect -542 7119 -508 7295
rect -446 7119 -412 7295
rect -332 7119 -298 7295
rect -236 7119 -202 7295
rect -122 7119 -88 7295
rect -26 7119 8 7295
rect 88 7119 122 7295
rect 184 7119 218 7295
rect 298 7119 332 7295
rect 394 7119 428 7295
rect 508 7119 542 7295
rect 604 7119 638 7295
rect 718 7119 752 7295
rect 814 7119 848 7295
rect 928 7119 962 7295
rect 1024 7119 1058 7295
rect 1138 7119 1172 7295
rect 1234 7119 1268 7295
rect 1348 7119 1382 7295
rect 1444 7119 1478 7295
rect 1558 7119 1592 7295
rect 1654 7119 1688 7295
rect 1768 7119 1802 7295
rect 1864 7119 1898 7295
rect 1978 7119 2012 7295
rect 2074 7119 2108 7295
rect 2188 7119 2222 7295
rect 2284 7119 2318 7295
rect 2398 7119 2432 7295
rect 2494 7119 2528 7295
rect 2608 7119 2642 7295
rect 2704 7119 2738 7295
rect 2818 7119 2852 7295
rect 2914 7119 2948 7295
rect 3028 7119 3062 7295
rect 3124 7119 3158 7295
rect 3238 7119 3272 7295
rect 3334 7119 3368 7295
rect 3448 7119 3482 7295
rect 3544 7119 3578 7295
rect 3658 7119 3692 7295
rect 3754 7119 3788 7295
rect 3868 7119 3902 7295
rect 3964 7119 3998 7295
rect 4078 7119 4112 7295
rect 4174 7119 4208 7295
rect 4288 7119 4322 7295
rect 4384 7119 4418 7295
rect 4498 7119 4532 7295
rect 4594 7119 4628 7295
rect 4708 7119 4742 7295
rect 4804 7119 4838 7295
rect 4918 7119 4952 7295
rect 5014 7119 5048 7295
rect 5128 7119 5162 7295
rect 5224 7119 5258 7295
rect 5338 7119 5372 7295
rect 5434 7119 5468 7295
rect 5548 7119 5582 7295
rect 5644 7119 5678 7295
rect 5758 7119 5792 7295
rect 5854 7119 5888 7295
rect 5968 7119 6002 7295
rect 6064 7119 6098 7295
rect -3555 5466 -3379 5500
rect -3555 5370 -3379 5404
rect -3555 5274 -3379 5308
rect -3555 5178 -3379 5212
rect -3555 5082 -3379 5116
rect -3555 4986 -3379 5020
rect -3555 4890 -3379 4924
rect -3555 4794 -3379 4828
rect -3555 4698 -3379 4732
rect -3555 4602 -3379 4636
rect -3555 4506 -3379 4540
rect -3555 4410 -3379 4444
rect -3555 4314 -3379 4348
rect -3555 4218 -3379 4252
rect -3555 4122 -3379 4156
rect -3555 4026 -3379 4060
rect -3555 3930 -3379 3964
rect -3555 3834 -3379 3868
rect -3555 3738 -3379 3772
rect 6843 7876 7019 7910
rect 6843 7780 7019 7814
rect 6843 7684 7019 7718
rect 6843 7588 7019 7622
rect 6843 7492 7019 7526
rect 6843 7396 7019 7430
rect 6843 7300 7019 7334
rect 6843 7204 7019 7238
rect 6843 7108 7019 7142
rect 6843 7012 7019 7046
rect 6843 6916 7019 6950
rect 6843 6820 7019 6854
rect 6843 6724 7019 6758
rect 6843 6628 7019 6662
rect 6843 6532 7019 6566
rect 6843 6436 7019 6470
rect 6843 6340 7019 6374
rect 6843 6244 7019 6278
rect 6843 6148 7019 6182
rect 6843 5466 7019 5500
rect 6843 5370 7019 5404
rect 6843 5274 7019 5308
rect 6843 5178 7019 5212
rect 6843 5082 7019 5116
rect 6843 4986 7019 5020
rect 6843 4890 7019 4924
rect 6843 4794 7019 4828
rect 6843 4698 7019 4732
rect 6843 4602 7019 4636
rect 6843 4506 7019 4540
rect 6843 4410 7019 4444
rect 6843 4314 7019 4348
rect 6843 4218 7019 4252
rect 6843 4122 7019 4156
rect 6843 4026 7019 4060
rect 6843 3930 7019 3964
rect 6843 3834 7019 3868
rect 6843 3738 7019 3772
<< psubdiff >>
rect 1246 9466 1293 9500
rect 1327 9466 1351 9500
rect 2101 9466 2125 9500
rect 2159 9466 2206 9500
rect -2744 6497 -2648 6531
rect 6130 6497 6226 6531
rect -2744 6435 -2710 6497
rect 6192 6435 6226 6497
rect -2744 4697 -2710 4759
rect 6192 4697 6226 4759
rect -2744 4663 -2648 4697
rect 6130 4663 6226 4697
rect -2744 4242 -2648 4276
rect 6130 4242 6226 4276
rect -2744 4180 -2710 4242
rect 6192 4180 6226 4242
rect -2744 682 -2710 745
rect 6192 682 6226 745
rect -2744 648 -2647 682
rect 6129 648 6226 682
rect -24 358 72 392
rect 3406 358 3502 392
rect -24 296 10 358
rect 3468 296 3502 358
rect -24 -122 10 -60
rect 3468 -122 3502 -60
rect -24 -156 72 -122
rect 3406 -156 3502 -122
<< nsubdiff >>
rect 1487 9466 1511 9500
rect 1545 9466 1604 9500
rect 1638 9466 1662 9500
rect 1790 9466 1814 9500
rect 1848 9466 1907 9500
rect 1941 9466 1965 9500
rect -3752 7990 -3656 8024
rect -3282 7990 -3186 8024
rect -3752 7928 -3718 7990
rect -3220 7928 -3186 7990
rect -3752 6068 -3718 6130
rect -2758 7989 -2662 8023
rect 6114 7989 6210 8023
rect -2758 7927 -2724 7989
rect 6176 7927 6210 7989
rect -2758 7395 -2724 7553
rect 6176 7395 6210 7553
rect -2758 6958 -2724 7020
rect 6176 6958 6210 7020
rect -2758 6924 -2662 6958
rect 6114 6924 6210 6958
rect 6648 7990 6744 8024
rect 7118 7990 7214 8024
rect 6648 7928 6682 7990
rect -3220 6068 -3186 6130
rect -3752 6034 -3656 6068
rect -3282 6034 -3186 6068
rect -3750 5580 -3654 5614
rect -3280 5580 -3184 5614
rect -3750 5518 -3716 5580
rect -3218 5518 -3184 5580
rect -3750 3658 -3716 3720
rect 7180 7928 7214 7990
rect 6648 6068 6682 6130
rect 7180 6068 7214 6130
rect 6648 6034 6744 6068
rect 7118 6034 7214 6068
rect 6648 5580 6744 5614
rect 7118 5580 7214 5614
rect 6648 5518 6682 5580
rect -3218 3658 -3184 3720
rect -3750 3624 -3654 3658
rect -3280 3624 -3184 3658
rect 7180 5518 7214 5580
rect 6648 3658 6682 3720
rect 7180 3658 7214 3720
rect 6648 3624 6744 3658
rect 7118 3624 7214 3658
<< psubdiffcont >>
rect 1293 9466 1327 9500
rect 2125 9466 2159 9500
rect -2648 6497 6130 6531
rect -2744 4759 -2710 6435
rect 6192 4759 6226 6435
rect -2648 4663 6130 4697
rect -2648 4242 6130 4276
rect -2744 745 -2710 4180
rect 6192 745 6226 4180
rect -2647 648 6129 682
rect 72 358 3406 392
rect -24 -60 10 296
rect 3468 -60 3502 296
rect 72 -156 3406 -122
<< nsubdiffcont >>
rect 1511 9466 1545 9500
rect 1604 9466 1638 9500
rect 1814 9466 1848 9500
rect 1907 9466 1941 9500
rect -3656 7990 -3282 8024
rect -3752 6130 -3718 7928
rect -3220 6130 -3186 7928
rect -2662 7989 6114 8023
rect -2758 7553 -2724 7927
rect 6176 7553 6210 7927
rect -2758 7020 -2724 7395
rect 6176 7020 6210 7395
rect -2662 6924 6114 6958
rect 6744 7990 7118 8024
rect -3656 6034 -3282 6068
rect -3654 5580 -3280 5614
rect -3750 3720 -3716 5518
rect -3218 3720 -3184 5518
rect 6648 6130 6682 7928
rect 7180 6130 7214 7928
rect 6744 6034 7118 6068
rect 6744 5580 7118 5614
rect -3654 3624 -3280 3658
rect 6648 3720 6682 5518
rect 7180 3720 7214 5518
rect 6744 3624 7118 3658
<< poly >>
rect 1203 9608 1229 10554
rect 1339 10062 1365 10554
rect 1407 10538 1505 10554
rect 1407 10504 1423 10538
rect 1457 10504 1505 10538
rect 1407 10410 1505 10504
rect 1407 10376 1423 10410
rect 1457 10376 1505 10410
rect 1407 10282 1505 10376
rect 1407 10248 1423 10282
rect 1457 10248 1505 10282
rect 1407 10154 1505 10248
rect 1407 10120 1423 10154
rect 1457 10120 1505 10154
rect 1407 10104 1505 10120
rect 1339 10046 1437 10062
rect 1339 10012 1387 10046
rect 1421 10012 1437 10046
rect 1339 9918 1437 10012
rect 1339 9884 1387 9918
rect 1421 9884 1437 9918
rect 1339 9790 1437 9884
rect 1339 9756 1387 9790
rect 1421 9756 1437 9790
rect 1339 9662 1437 9756
rect 1339 9628 1387 9662
rect 1421 9628 1437 9662
rect 1339 9608 1437 9628
rect 1479 9608 1505 10104
rect 1679 9608 1705 10554
rect 1747 9608 1773 10554
rect 1947 10058 1973 10554
rect 2015 10534 2113 10554
rect 2015 10500 2031 10534
rect 2065 10500 2113 10534
rect 2015 10406 2113 10500
rect 2015 10372 2031 10406
rect 2065 10372 2113 10406
rect 2015 10278 2113 10372
rect 2015 10244 2031 10278
rect 2065 10244 2113 10278
rect 2015 10150 2113 10244
rect 2015 10116 2031 10150
rect 2065 10116 2113 10150
rect 2015 10100 2113 10116
rect 1947 10042 2045 10058
rect 1947 10008 1995 10042
rect 2029 10008 2045 10042
rect 1947 9914 2045 10008
rect 1947 9880 1995 9914
rect 2029 9880 2045 9914
rect 1947 9786 2045 9880
rect 1947 9752 1995 9786
rect 2029 9752 2045 9786
rect 1947 9658 2045 9752
rect 1947 9624 1995 9658
rect 2029 9624 2045 9658
rect 1947 9608 2045 9624
rect 2087 9608 2113 10100
rect 2223 9608 2249 10554
rect 1381 9399 1447 9415
rect 1381 9365 1397 9399
rect 1431 9365 1447 9399
rect 1381 9358 1447 9365
rect 2005 9399 2071 9415
rect 2005 9365 2021 9399
rect 2055 9365 2071 9399
rect 2005 9358 2071 9365
rect 1203 9328 1229 9358
rect 1359 9328 1479 9358
rect 1679 9328 1705 9358
rect 1747 9328 1773 9358
rect 1973 9328 2093 9358
rect 2223 9328 2249 9358
rect 1381 9318 1447 9328
rect 1381 9284 1397 9318
rect 1431 9284 1447 9318
rect 1381 9274 1447 9284
rect 2005 9318 2071 9328
rect 2005 9284 2021 9318
rect 2055 9284 2071 9318
rect 2005 9274 2071 9284
rect 1203 9244 1229 9274
rect 1359 9244 1479 9274
rect 1679 9244 1705 9274
rect 1747 9244 1773 9274
rect 1973 9244 2093 9274
rect 2223 9244 2249 9274
rect 1381 9234 1447 9244
rect 1381 9200 1397 9234
rect 1431 9200 1447 9234
rect 1381 9190 1447 9200
rect 2005 9234 2071 9244
rect 2005 9200 2021 9234
rect 2055 9200 2071 9234
rect 2005 9190 2071 9200
rect 1203 9160 1229 9190
rect 1359 9160 1479 9190
rect 1679 9160 1705 9190
rect 1747 9160 1773 9190
rect 1973 9160 2093 9190
rect 2223 9160 2249 9190
rect 1381 9150 1447 9160
rect 1381 9116 1397 9150
rect 1431 9116 1447 9150
rect 1381 9106 1447 9116
rect 2005 9150 2071 9160
rect 2005 9116 2021 9150
rect 2055 9116 2071 9150
rect 2005 9106 2071 9116
rect 1203 9076 1229 9106
rect 1359 9076 1479 9106
rect 1679 9076 1705 9106
rect 1747 9076 1773 9106
rect 1973 9076 2093 9106
rect 2223 9076 2249 9106
rect 1203 8992 1229 9022
rect 1359 8992 1479 9022
rect 1679 8992 1705 9022
rect 1747 8992 1773 9022
rect 1973 8992 2093 9022
rect 2223 8992 2249 9022
rect 1381 8938 1447 8992
rect 2005 8938 2071 8992
rect 1203 8908 1229 8938
rect 1359 8908 1479 8938
rect 1679 8908 1705 8938
rect 1747 8908 1773 8938
rect 1973 8908 2093 8938
rect 2223 8908 2249 8938
rect 1381 8898 1447 8908
rect 1381 8864 1397 8898
rect 1431 8864 1447 8898
rect 1381 8854 1447 8864
rect 2005 8898 2071 8908
rect 2005 8864 2021 8898
rect 2055 8864 2071 8898
rect 2005 8854 2071 8864
rect 1203 8824 1229 8854
rect 1359 8824 1479 8854
rect 1679 8824 1705 8854
rect 1747 8824 1773 8854
rect 1973 8824 2093 8854
rect 2223 8824 2249 8854
rect 1381 8814 1447 8824
rect 1381 8780 1397 8814
rect 1431 8780 1447 8814
rect 1381 8770 1447 8780
rect 2005 8814 2071 8824
rect 2005 8780 2021 8814
rect 2055 8780 2071 8814
rect 2005 8770 2071 8780
rect 1203 8740 1229 8770
rect 1359 8740 1479 8770
rect 1679 8740 1705 8770
rect 1747 8740 1773 8770
rect 1973 8740 2093 8770
rect 2223 8740 2249 8770
rect 1203 8499 1229 8529
rect 1359 8499 1479 8529
rect 1679 8499 1705 8529
rect 1747 8499 1773 8529
rect 1973 8499 2093 8529
rect 2223 8499 2249 8529
rect 1381 8445 1447 8499
rect 2005 8445 2071 8499
rect 1203 8415 1229 8445
rect 1359 8436 1479 8445
rect 1359 8415 1397 8436
rect 1381 8402 1397 8415
rect 1431 8415 1479 8436
rect 1679 8415 1705 8445
rect 1747 8415 1773 8445
rect 1973 8436 2093 8445
rect 1973 8415 2021 8436
rect 1431 8402 1447 8415
rect 1381 8392 1447 8402
rect 2005 8402 2021 8415
rect 2055 8415 2093 8436
rect 2223 8415 2249 8445
rect 2055 8402 2071 8415
rect 2005 8392 2071 8402
rect 1203 8320 1229 8350
rect 1313 8320 1543 8350
rect 1671 8320 1697 8350
rect 1755 8320 1781 8350
rect 1909 8320 2139 8350
rect 2223 8320 2249 8350
rect 1381 8312 1447 8320
rect 1381 8278 1397 8312
rect 1431 8278 1447 8312
rect 1381 8268 1447 8278
rect 2005 8312 2071 8320
rect 2005 8278 2021 8312
rect 2055 8278 2071 8312
rect 2005 8268 2071 8278
rect -3666 7862 -3600 7878
rect -3666 7828 -3650 7862
rect -3616 7860 -3600 7862
rect -3616 7830 -3569 7860
rect -3369 7830 -3342 7860
rect -3616 7828 -3600 7830
rect -3666 7812 -3600 7828
rect -3338 7766 -3272 7782
rect -3338 7764 -3322 7766
rect -3596 7734 -3569 7764
rect -3369 7734 -3322 7764
rect -3666 7670 -3600 7686
rect -3666 7636 -3650 7670
rect -3616 7668 -3600 7670
rect -3338 7732 -3322 7734
rect -3288 7732 -3272 7766
rect -3338 7716 -3272 7732
rect -3616 7638 -3569 7668
rect -3369 7638 -3342 7668
rect -3616 7636 -3600 7638
rect -3666 7620 -3600 7636
rect -3338 7574 -3272 7590
rect -3338 7572 -3322 7574
rect -3596 7542 -3569 7572
rect -3369 7542 -3322 7572
rect -3666 7478 -3600 7494
rect -3666 7444 -3650 7478
rect -3616 7476 -3600 7478
rect -3338 7540 -3322 7542
rect -3288 7540 -3272 7574
rect -3338 7524 -3272 7540
rect -3616 7446 -3569 7476
rect -3369 7446 -3342 7476
rect -3616 7444 -3600 7446
rect -3666 7428 -3600 7444
rect -3338 7382 -3272 7398
rect -3338 7380 -3322 7382
rect -3596 7350 -3569 7380
rect -3369 7350 -3322 7380
rect -3666 7286 -3600 7302
rect -3666 7252 -3650 7286
rect -3616 7284 -3600 7286
rect -3338 7348 -3322 7350
rect -3288 7348 -3272 7382
rect -3338 7332 -3272 7348
rect -3616 7254 -3569 7284
rect -3369 7254 -3342 7284
rect -3616 7252 -3600 7254
rect -3666 7236 -3600 7252
rect -3338 7190 -3272 7206
rect -3338 7188 -3322 7190
rect -3596 7158 -3569 7188
rect -3369 7158 -3322 7188
rect -3666 7094 -3600 7110
rect -3666 7060 -3650 7094
rect -3616 7092 -3600 7094
rect -3338 7156 -3322 7158
rect -3288 7156 -3272 7190
rect -3338 7140 -3272 7156
rect -3616 7062 -3569 7092
rect -3369 7062 -3342 7092
rect -3616 7060 -3600 7062
rect -3666 7044 -3600 7060
rect -3338 6998 -3272 7014
rect -3338 6996 -3322 6998
rect -3596 6966 -3569 6996
rect -3369 6966 -3322 6996
rect -3666 6902 -3600 6918
rect -3666 6868 -3650 6902
rect -3616 6900 -3600 6902
rect -3338 6964 -3322 6966
rect -3288 6964 -3272 6998
rect -3338 6948 -3272 6964
rect -3616 6870 -3569 6900
rect -3369 6870 -3342 6900
rect -3616 6868 -3600 6870
rect -3666 6852 -3600 6868
rect -3338 6806 -3272 6822
rect -3338 6804 -3322 6806
rect -3596 6774 -3569 6804
rect -3369 6774 -3322 6804
rect -3666 6710 -3600 6726
rect -3666 6676 -3650 6710
rect -3616 6708 -3600 6710
rect -3338 6772 -3322 6774
rect -3288 6772 -3272 6806
rect -3338 6756 -3272 6772
rect -3616 6678 -3569 6708
rect -3369 6678 -3342 6708
rect -3616 6676 -3600 6678
rect -3666 6660 -3600 6676
rect -3338 6614 -3272 6630
rect -3338 6612 -3322 6614
rect -3596 6582 -3569 6612
rect -3369 6582 -3322 6612
rect -3666 6518 -3600 6534
rect -3666 6484 -3650 6518
rect -3616 6516 -3600 6518
rect -3338 6580 -3322 6582
rect -3288 6580 -3272 6614
rect -3338 6564 -3272 6580
rect -3616 6486 -3569 6516
rect -3369 6486 -3342 6516
rect -3616 6484 -3600 6486
rect -3666 6468 -3600 6484
rect -3338 6422 -3272 6438
rect -3338 6420 -3322 6422
rect -3596 6390 -3569 6420
rect -3369 6390 -3322 6420
rect -3666 6326 -3600 6342
rect -3666 6292 -3650 6326
rect -3616 6324 -3600 6326
rect -3338 6388 -3322 6390
rect -3288 6388 -3272 6422
rect -3338 6372 -3272 6388
rect -3616 6294 -3569 6324
rect -3369 6294 -3342 6324
rect -3616 6292 -3600 6294
rect -3666 6276 -3600 6292
rect -3338 6230 -3272 6246
rect -3338 6228 -3322 6230
rect -3596 6198 -3569 6228
rect -3369 6198 -3322 6228
rect -3338 6196 -3322 6198
rect -3288 6196 -3272 6230
rect -3338 6180 -3272 6196
rect -2402 7921 -2336 7937
rect -2402 7887 -2386 7921
rect -2352 7887 -2336 7921
rect -2402 7871 -2336 7887
rect -1982 7921 -1916 7937
rect -1982 7887 -1966 7921
rect -1932 7887 -1916 7921
rect -1982 7871 -1916 7887
rect -1562 7921 -1496 7937
rect -1562 7887 -1546 7921
rect -1512 7887 -1496 7921
rect -1562 7871 -1496 7887
rect -1142 7921 -1076 7937
rect -1142 7887 -1126 7921
rect -1092 7887 -1076 7921
rect -1142 7871 -1076 7887
rect -722 7921 -656 7937
rect -722 7887 -706 7921
rect -672 7887 -656 7921
rect -722 7871 -656 7887
rect -302 7921 -236 7937
rect -302 7887 -286 7921
rect -252 7887 -236 7921
rect -302 7871 -236 7887
rect 118 7921 184 7937
rect 118 7887 134 7921
rect 168 7887 184 7921
rect 118 7871 184 7887
rect 538 7921 604 7937
rect 538 7887 554 7921
rect 588 7887 604 7921
rect 538 7871 604 7887
rect 958 7921 1024 7937
rect 958 7887 974 7921
rect 1008 7887 1024 7921
rect 958 7871 1024 7887
rect 1378 7921 1444 7937
rect 1378 7887 1394 7921
rect 1428 7887 1444 7921
rect 1378 7871 1444 7887
rect 1798 7921 1864 7937
rect 1798 7887 1814 7921
rect 1848 7887 1864 7921
rect 1798 7871 1864 7887
rect 2218 7921 2284 7937
rect 2218 7887 2234 7921
rect 2268 7887 2284 7921
rect 2218 7871 2284 7887
rect 2638 7921 2704 7937
rect 2638 7887 2654 7921
rect 2688 7887 2704 7921
rect 2638 7871 2704 7887
rect 3058 7921 3124 7937
rect 3058 7887 3074 7921
rect 3108 7887 3124 7921
rect 3058 7871 3124 7887
rect 3478 7921 3544 7937
rect 3478 7887 3494 7921
rect 3528 7887 3544 7921
rect 3478 7871 3544 7887
rect 3898 7921 3964 7937
rect 3898 7887 3914 7921
rect 3948 7887 3964 7921
rect 3898 7871 3964 7887
rect 4318 7921 4384 7937
rect 4318 7887 4334 7921
rect 4368 7887 4384 7921
rect 4318 7871 4384 7887
rect 4738 7921 4804 7937
rect 4738 7887 4754 7921
rect 4788 7887 4804 7921
rect 4738 7871 4804 7887
rect 5158 7921 5224 7937
rect 5158 7887 5174 7921
rect 5208 7887 5224 7921
rect 5158 7871 5224 7887
rect 5578 7921 5644 7937
rect 5578 7887 5594 7921
rect 5628 7887 5644 7921
rect 5578 7871 5644 7887
rect 5998 7921 6064 7937
rect 5998 7887 6014 7921
rect 6048 7887 6064 7921
rect 5998 7871 6064 7887
rect -2594 7840 -2564 7867
rect -2384 7840 -2354 7871
rect -2174 7840 -2144 7867
rect -1964 7840 -1934 7871
rect -1754 7840 -1724 7867
rect -1544 7840 -1514 7871
rect -1334 7840 -1304 7867
rect -1124 7840 -1094 7871
rect -914 7840 -884 7867
rect -704 7840 -674 7871
rect -494 7840 -464 7867
rect -284 7840 -254 7871
rect -74 7840 -44 7867
rect 136 7840 166 7871
rect 346 7840 376 7867
rect 556 7840 586 7871
rect 766 7840 796 7867
rect 976 7840 1006 7871
rect 1186 7840 1216 7867
rect 1396 7840 1426 7871
rect 1606 7840 1636 7867
rect 1816 7840 1846 7871
rect 2026 7840 2056 7867
rect 2236 7840 2266 7871
rect 2446 7840 2476 7867
rect 2656 7840 2686 7871
rect 2866 7840 2896 7867
rect 3076 7840 3106 7871
rect 3286 7840 3316 7867
rect 3496 7840 3526 7871
rect 3706 7840 3736 7867
rect 3916 7840 3946 7871
rect 4126 7840 4156 7867
rect 4336 7840 4366 7871
rect 4546 7840 4576 7867
rect 4756 7840 4786 7871
rect 4966 7840 4996 7867
rect 5176 7840 5206 7871
rect 5386 7840 5416 7867
rect 5596 7840 5626 7871
rect 5806 7840 5836 7867
rect 6016 7840 6046 7871
rect -2594 7609 -2564 7640
rect -2384 7613 -2354 7640
rect -2174 7609 -2144 7640
rect -1964 7613 -1934 7640
rect -1754 7609 -1724 7640
rect -1544 7613 -1514 7640
rect -1334 7609 -1304 7640
rect -1124 7613 -1094 7640
rect -914 7609 -884 7640
rect -704 7613 -674 7640
rect -494 7609 -464 7640
rect -284 7613 -254 7640
rect -74 7609 -44 7640
rect 136 7613 166 7640
rect 346 7609 376 7640
rect 556 7613 586 7640
rect 766 7609 796 7640
rect 976 7613 1006 7640
rect 1186 7609 1216 7640
rect 1396 7613 1426 7640
rect 1606 7609 1636 7640
rect 1816 7613 1846 7640
rect 2026 7609 2056 7640
rect 2236 7613 2266 7640
rect 2446 7609 2476 7640
rect 2656 7613 2686 7640
rect 2866 7609 2896 7640
rect 3076 7613 3106 7640
rect 3286 7609 3316 7640
rect 3496 7613 3526 7640
rect 3706 7609 3736 7640
rect 3916 7613 3946 7640
rect 4126 7609 4156 7640
rect 4336 7613 4366 7640
rect 4546 7609 4576 7640
rect 4756 7613 4786 7640
rect 4966 7609 4996 7640
rect 5176 7613 5206 7640
rect 5386 7609 5416 7640
rect 5596 7613 5626 7640
rect 5806 7609 5836 7640
rect 6016 7613 6046 7640
rect -2612 7593 -2546 7609
rect -2612 7559 -2596 7593
rect -2562 7559 -2546 7593
rect -2612 7543 -2546 7559
rect -2192 7593 -2126 7609
rect -2192 7559 -2176 7593
rect -2142 7559 -2126 7593
rect -2192 7543 -2126 7559
rect -1772 7593 -1706 7609
rect -1772 7559 -1756 7593
rect -1722 7559 -1706 7593
rect -1772 7543 -1706 7559
rect -1352 7593 -1286 7609
rect -1352 7559 -1336 7593
rect -1302 7559 -1286 7593
rect -1352 7543 -1286 7559
rect -932 7593 -866 7609
rect -932 7559 -916 7593
rect -882 7559 -866 7593
rect -932 7543 -866 7559
rect -512 7593 -446 7609
rect -512 7559 -496 7593
rect -462 7559 -446 7593
rect -512 7543 -446 7559
rect -92 7593 -26 7609
rect -92 7559 -76 7593
rect -42 7559 -26 7593
rect -92 7543 -26 7559
rect 328 7593 394 7609
rect 328 7559 344 7593
rect 378 7559 394 7593
rect 328 7543 394 7559
rect 748 7593 814 7609
rect 748 7559 764 7593
rect 798 7559 814 7593
rect 748 7543 814 7559
rect 1168 7593 1234 7609
rect 1168 7559 1184 7593
rect 1218 7559 1234 7593
rect 1168 7543 1234 7559
rect 1588 7593 1654 7609
rect 1588 7559 1604 7593
rect 1638 7559 1654 7593
rect 1588 7543 1654 7559
rect 2008 7593 2074 7609
rect 2008 7559 2024 7593
rect 2058 7559 2074 7593
rect 2008 7543 2074 7559
rect 2428 7593 2494 7609
rect 2428 7559 2444 7593
rect 2478 7559 2494 7593
rect 2428 7543 2494 7559
rect 2848 7593 2914 7609
rect 2848 7559 2864 7593
rect 2898 7559 2914 7593
rect 2848 7543 2914 7559
rect 3268 7593 3334 7609
rect 3268 7559 3284 7593
rect 3318 7559 3334 7593
rect 3268 7543 3334 7559
rect 3688 7593 3754 7609
rect 3688 7559 3704 7593
rect 3738 7559 3754 7593
rect 3688 7543 3754 7559
rect 4108 7593 4174 7609
rect 4108 7559 4124 7593
rect 4158 7559 4174 7593
rect 4108 7543 4174 7559
rect 4528 7593 4594 7609
rect 4528 7559 4544 7593
rect 4578 7559 4594 7593
rect 4528 7543 4594 7559
rect 4948 7593 5014 7609
rect 4948 7559 4964 7593
rect 4998 7559 5014 7593
rect 4948 7543 5014 7559
rect 5368 7593 5434 7609
rect 5368 7559 5384 7593
rect 5418 7559 5434 7593
rect 5368 7543 5434 7559
rect 5788 7593 5854 7609
rect 5788 7559 5804 7593
rect 5838 7559 5854 7593
rect 5788 7543 5854 7559
rect -2400 7389 -2334 7405
rect -2400 7355 -2384 7389
rect -2350 7355 -2334 7389
rect -2400 7339 -2334 7355
rect -1980 7389 -1914 7405
rect -1980 7355 -1964 7389
rect -1930 7355 -1914 7389
rect -1980 7339 -1914 7355
rect -1560 7389 -1494 7405
rect -1560 7355 -1544 7389
rect -1510 7355 -1494 7389
rect -1560 7339 -1494 7355
rect -1140 7389 -1074 7405
rect -1140 7355 -1124 7389
rect -1090 7355 -1074 7389
rect -1140 7339 -1074 7355
rect -720 7389 -654 7405
rect -720 7355 -704 7389
rect -670 7355 -654 7389
rect -720 7339 -654 7355
rect -300 7389 -234 7405
rect -300 7355 -284 7389
rect -250 7355 -234 7389
rect -300 7339 -234 7355
rect 120 7389 186 7405
rect 120 7355 136 7389
rect 170 7355 186 7389
rect 120 7339 186 7355
rect 540 7389 606 7405
rect 540 7355 556 7389
rect 590 7355 606 7389
rect 540 7339 606 7355
rect 960 7389 1026 7405
rect 960 7355 976 7389
rect 1010 7355 1026 7389
rect 960 7339 1026 7355
rect 1380 7389 1446 7405
rect 1380 7355 1396 7389
rect 1430 7355 1446 7389
rect 1380 7339 1446 7355
rect 1800 7389 1866 7405
rect 1800 7355 1816 7389
rect 1850 7355 1866 7389
rect 1800 7339 1866 7355
rect 2220 7389 2286 7405
rect 2220 7355 2236 7389
rect 2270 7355 2286 7389
rect 2220 7339 2286 7355
rect 2640 7389 2706 7405
rect 2640 7355 2656 7389
rect 2690 7355 2706 7389
rect 2640 7339 2706 7355
rect 3060 7389 3126 7405
rect 3060 7355 3076 7389
rect 3110 7355 3126 7389
rect 3060 7339 3126 7355
rect 3480 7389 3546 7405
rect 3480 7355 3496 7389
rect 3530 7355 3546 7389
rect 3480 7339 3546 7355
rect 3900 7389 3966 7405
rect 3900 7355 3916 7389
rect 3950 7355 3966 7389
rect 3900 7339 3966 7355
rect 4320 7389 4386 7405
rect 4320 7355 4336 7389
rect 4370 7355 4386 7389
rect 4320 7339 4386 7355
rect 4740 7389 4806 7405
rect 4740 7355 4756 7389
rect 4790 7355 4806 7389
rect 4740 7339 4806 7355
rect 5160 7389 5226 7405
rect 5160 7355 5176 7389
rect 5210 7355 5226 7389
rect 5160 7339 5226 7355
rect 5580 7389 5646 7405
rect 5580 7355 5596 7389
rect 5630 7355 5646 7389
rect 5580 7339 5646 7355
rect 6000 7389 6066 7405
rect 6000 7355 6016 7389
rect 6050 7355 6066 7389
rect 6000 7339 6066 7355
rect -2592 7307 -2562 7333
rect -2382 7307 -2352 7339
rect -2172 7307 -2142 7333
rect -1962 7307 -1932 7339
rect -1752 7307 -1722 7333
rect -1542 7307 -1512 7339
rect -1332 7307 -1302 7333
rect -1122 7307 -1092 7339
rect -912 7307 -882 7333
rect -702 7307 -672 7339
rect -492 7307 -462 7333
rect -282 7307 -252 7339
rect -72 7307 -42 7333
rect 138 7307 168 7339
rect 348 7307 378 7333
rect 558 7307 588 7339
rect 768 7307 798 7333
rect 978 7307 1008 7339
rect 1188 7307 1218 7333
rect 1398 7307 1428 7339
rect 1608 7307 1638 7333
rect 1818 7307 1848 7339
rect 2028 7307 2058 7333
rect 2238 7307 2268 7339
rect 2448 7307 2478 7333
rect 2658 7307 2688 7339
rect 2868 7307 2898 7333
rect 3078 7307 3108 7339
rect 3288 7307 3318 7333
rect 3498 7307 3528 7339
rect 3708 7307 3738 7333
rect 3918 7307 3948 7339
rect 4128 7307 4158 7333
rect 4338 7307 4368 7339
rect 4548 7307 4578 7333
rect 4758 7307 4788 7339
rect 4968 7307 4998 7333
rect 5178 7307 5208 7339
rect 5388 7307 5418 7333
rect 5598 7307 5628 7339
rect 5808 7307 5838 7333
rect 6018 7307 6048 7339
rect -2592 7076 -2562 7107
rect -2382 7080 -2352 7107
rect -2172 7076 -2142 7107
rect -1962 7080 -1932 7107
rect -1752 7076 -1722 7107
rect -1542 7080 -1512 7107
rect -1332 7076 -1302 7107
rect -1122 7080 -1092 7107
rect -912 7076 -882 7107
rect -702 7080 -672 7107
rect -492 7076 -462 7107
rect -282 7080 -252 7107
rect -72 7076 -42 7107
rect 138 7080 168 7107
rect 348 7076 378 7107
rect 558 7080 588 7107
rect 768 7076 798 7107
rect 978 7080 1008 7107
rect 1188 7076 1218 7107
rect 1398 7080 1428 7107
rect 1608 7076 1638 7107
rect 1818 7080 1848 7107
rect 2028 7076 2058 7107
rect 2238 7080 2268 7107
rect 2448 7076 2478 7107
rect 2658 7080 2688 7107
rect 2868 7076 2898 7107
rect 3078 7080 3108 7107
rect 3288 7076 3318 7107
rect 3498 7080 3528 7107
rect 3708 7076 3738 7107
rect 3918 7080 3948 7107
rect 4128 7076 4158 7107
rect 4338 7080 4368 7107
rect 4548 7076 4578 7107
rect 4758 7080 4788 7107
rect 4968 7076 4998 7107
rect 5178 7080 5208 7107
rect 5388 7076 5418 7107
rect 5598 7080 5628 7107
rect 5808 7076 5838 7107
rect 6018 7080 6048 7107
rect -2610 7060 -2544 7076
rect -2610 7026 -2594 7060
rect -2560 7026 -2544 7060
rect -2610 7010 -2544 7026
rect -2190 7060 -2124 7076
rect -2190 7026 -2174 7060
rect -2140 7026 -2124 7060
rect -2190 7010 -2124 7026
rect -1770 7060 -1704 7076
rect -1770 7026 -1754 7060
rect -1720 7026 -1704 7060
rect -1770 7010 -1704 7026
rect -1350 7060 -1284 7076
rect -1350 7026 -1334 7060
rect -1300 7026 -1284 7060
rect -1350 7010 -1284 7026
rect -930 7060 -864 7076
rect -930 7026 -914 7060
rect -880 7026 -864 7060
rect -930 7010 -864 7026
rect -510 7060 -444 7076
rect -510 7026 -494 7060
rect -460 7026 -444 7060
rect -510 7010 -444 7026
rect -90 7060 -24 7076
rect -90 7026 -74 7060
rect -40 7026 -24 7060
rect -90 7010 -24 7026
rect 330 7060 396 7076
rect 330 7026 346 7060
rect 380 7026 396 7060
rect 330 7010 396 7026
rect 750 7060 816 7076
rect 750 7026 766 7060
rect 800 7026 816 7060
rect 750 7010 816 7026
rect 1170 7060 1236 7076
rect 1170 7026 1186 7060
rect 1220 7026 1236 7060
rect 1170 7010 1236 7026
rect 1590 7060 1656 7076
rect 1590 7026 1606 7060
rect 1640 7026 1656 7060
rect 1590 7010 1656 7026
rect 2010 7060 2076 7076
rect 2010 7026 2026 7060
rect 2060 7026 2076 7060
rect 2010 7010 2076 7026
rect 2430 7060 2496 7076
rect 2430 7026 2446 7060
rect 2480 7026 2496 7060
rect 2430 7010 2496 7026
rect 2850 7060 2916 7076
rect 2850 7026 2866 7060
rect 2900 7026 2916 7060
rect 2850 7010 2916 7026
rect 3270 7060 3336 7076
rect 3270 7026 3286 7060
rect 3320 7026 3336 7060
rect 3270 7010 3336 7026
rect 3690 7060 3756 7076
rect 3690 7026 3706 7060
rect 3740 7026 3756 7060
rect 3690 7010 3756 7026
rect 4110 7060 4176 7076
rect 4110 7026 4126 7060
rect 4160 7026 4176 7060
rect 4110 7010 4176 7026
rect 4530 7060 4596 7076
rect 4530 7026 4546 7060
rect 4580 7026 4596 7060
rect 4530 7010 4596 7026
rect 4950 7060 5016 7076
rect 4950 7026 4966 7060
rect 5000 7026 5016 7060
rect 4950 7010 5016 7026
rect 5370 7060 5436 7076
rect 5370 7026 5386 7060
rect 5420 7026 5436 7060
rect 5370 7010 5436 7026
rect 5790 7060 5856 7076
rect 5790 7026 5806 7060
rect 5840 7026 5856 7060
rect 5790 7010 5856 7026
rect -3664 5452 -3598 5468
rect -3664 5418 -3648 5452
rect -3614 5450 -3598 5452
rect -3614 5420 -3567 5450
rect -3367 5420 -3340 5450
rect -3614 5418 -3598 5420
rect -3664 5402 -3598 5418
rect -3336 5356 -3270 5372
rect -3336 5354 -3320 5356
rect -3594 5324 -3567 5354
rect -3367 5324 -3320 5354
rect -3664 5260 -3598 5276
rect -3664 5226 -3648 5260
rect -3614 5258 -3598 5260
rect -3336 5322 -3320 5324
rect -3286 5322 -3270 5356
rect -3336 5306 -3270 5322
rect -3614 5228 -3567 5258
rect -3367 5228 -3340 5258
rect -3614 5226 -3598 5228
rect -3664 5210 -3598 5226
rect -3336 5164 -3270 5180
rect -3336 5162 -3320 5164
rect -3594 5132 -3567 5162
rect -3367 5132 -3320 5162
rect -3664 5068 -3598 5084
rect -3664 5034 -3648 5068
rect -3614 5066 -3598 5068
rect -3336 5130 -3320 5132
rect -3286 5130 -3270 5164
rect -3336 5114 -3270 5130
rect -3614 5036 -3567 5066
rect -3367 5036 -3340 5066
rect -3614 5034 -3598 5036
rect -3664 5018 -3598 5034
rect -3336 4972 -3270 4988
rect -3336 4970 -3320 4972
rect -3594 4940 -3567 4970
rect -3367 4940 -3320 4970
rect -3664 4876 -3598 4892
rect -3664 4842 -3648 4876
rect -3614 4874 -3598 4876
rect -3336 4938 -3320 4940
rect -3286 4938 -3270 4972
rect -3336 4922 -3270 4938
rect -3614 4844 -3567 4874
rect -3367 4844 -3340 4874
rect -3614 4842 -3598 4844
rect -3664 4826 -3598 4842
rect -3336 4780 -3270 4796
rect -3336 4778 -3320 4780
rect -3594 4748 -3567 4778
rect -3367 4748 -3320 4778
rect -3664 4684 -3598 4700
rect -3664 4650 -3648 4684
rect -3614 4682 -3598 4684
rect -3336 4746 -3320 4748
rect -3286 4746 -3270 4780
rect -3336 4730 -3270 4746
rect -3614 4652 -3567 4682
rect -3367 4652 -3340 4682
rect -3614 4650 -3598 4652
rect -3664 4634 -3598 4650
rect -3336 4588 -3270 4604
rect -3336 4586 -3320 4588
rect -3594 4556 -3567 4586
rect -3367 4556 -3320 4586
rect -3664 4492 -3598 4508
rect -3664 4458 -3648 4492
rect -3614 4490 -3598 4492
rect -3336 4554 -3320 4556
rect -3286 4554 -3270 4588
rect -3336 4538 -3270 4554
rect -3614 4460 -3567 4490
rect -3367 4460 -3340 4490
rect -3614 4458 -3598 4460
rect -3664 4442 -3598 4458
rect -3336 4396 -3270 4412
rect -3336 4394 -3320 4396
rect -3594 4364 -3567 4394
rect -3367 4364 -3320 4394
rect -3664 4300 -3598 4316
rect -3664 4266 -3648 4300
rect -3614 4298 -3598 4300
rect -3336 4362 -3320 4364
rect -3286 4362 -3270 4396
rect -3336 4346 -3270 4362
rect -3614 4268 -3567 4298
rect -3367 4268 -3340 4298
rect -3614 4266 -3598 4268
rect -3664 4250 -3598 4266
rect -3336 4204 -3270 4220
rect -3336 4202 -3320 4204
rect -3594 4172 -3567 4202
rect -3367 4172 -3320 4202
rect -3664 4108 -3598 4124
rect -3664 4074 -3648 4108
rect -3614 4106 -3598 4108
rect -3336 4170 -3320 4172
rect -3286 4170 -3270 4204
rect -3336 4154 -3270 4170
rect -3614 4076 -3567 4106
rect -3367 4076 -3340 4106
rect -3614 4074 -3598 4076
rect -3664 4058 -3598 4074
rect -3336 4012 -3270 4028
rect -3336 4010 -3320 4012
rect -3594 3980 -3567 4010
rect -3367 3980 -3320 4010
rect -3664 3916 -3598 3932
rect -3664 3882 -3648 3916
rect -3614 3914 -3598 3916
rect -3336 3978 -3320 3980
rect -3286 3978 -3270 4012
rect -3336 3962 -3270 3978
rect -3614 3884 -3567 3914
rect -3367 3884 -3340 3914
rect -3614 3882 -3598 3884
rect -3664 3866 -3598 3882
rect -3336 3820 -3270 3836
rect -3336 3818 -3320 3820
rect -3594 3788 -3567 3818
rect -3367 3788 -3320 3818
rect -3336 3786 -3320 3788
rect -3286 3786 -3270 3820
rect -3336 3770 -3270 3786
rect -2388 6429 -2322 6445
rect -2388 6395 -2372 6429
rect -2338 6395 -2322 6429
rect -2580 6357 -2550 6383
rect -2388 6379 -2322 6395
rect -1968 6429 -1902 6445
rect -1968 6395 -1952 6429
rect -1918 6395 -1902 6429
rect -2370 6357 -2340 6379
rect -2160 6357 -2130 6383
rect -1968 6379 -1902 6395
rect -1548 6429 -1482 6445
rect -1548 6395 -1532 6429
rect -1498 6395 -1482 6429
rect -1950 6357 -1920 6379
rect -1740 6357 -1710 6383
rect -1548 6379 -1482 6395
rect -1128 6429 -1062 6445
rect -1128 6395 -1112 6429
rect -1078 6395 -1062 6429
rect -1530 6357 -1500 6379
rect -1320 6357 -1290 6383
rect -1128 6379 -1062 6395
rect -708 6429 -642 6445
rect -708 6395 -692 6429
rect -658 6395 -642 6429
rect -1110 6357 -1080 6379
rect -900 6357 -870 6383
rect -708 6379 -642 6395
rect -288 6429 -222 6445
rect -288 6395 -272 6429
rect -238 6395 -222 6429
rect -690 6357 -660 6379
rect -480 6357 -450 6383
rect -288 6379 -222 6395
rect 132 6429 198 6445
rect 132 6395 148 6429
rect 182 6395 198 6429
rect -270 6357 -240 6379
rect -60 6357 -30 6383
rect 132 6379 198 6395
rect 552 6429 618 6445
rect 552 6395 568 6429
rect 602 6395 618 6429
rect 150 6357 180 6379
rect 360 6357 390 6383
rect 552 6379 618 6395
rect 972 6429 1038 6445
rect 972 6395 988 6429
rect 1022 6395 1038 6429
rect 570 6357 600 6379
rect 780 6357 810 6383
rect 972 6379 1038 6395
rect 1392 6429 1458 6445
rect 1392 6395 1408 6429
rect 1442 6395 1458 6429
rect 990 6357 1020 6379
rect 1200 6357 1230 6383
rect 1392 6379 1458 6395
rect 1812 6429 1878 6445
rect 1812 6395 1828 6429
rect 1862 6395 1878 6429
rect 1410 6357 1440 6379
rect 1620 6357 1650 6383
rect 1812 6379 1878 6395
rect 2232 6429 2298 6445
rect 2232 6395 2248 6429
rect 2282 6395 2298 6429
rect 1830 6357 1860 6379
rect 2040 6357 2070 6383
rect 2232 6379 2298 6395
rect 2652 6429 2718 6445
rect 2652 6395 2668 6429
rect 2702 6395 2718 6429
rect 2250 6357 2280 6379
rect 2460 6357 2490 6383
rect 2652 6379 2718 6395
rect 3072 6429 3138 6445
rect 3072 6395 3088 6429
rect 3122 6395 3138 6429
rect 2670 6357 2700 6379
rect 2880 6357 2910 6383
rect 3072 6379 3138 6395
rect 3492 6429 3558 6445
rect 3492 6395 3508 6429
rect 3542 6395 3558 6429
rect 3090 6357 3120 6379
rect 3300 6357 3330 6383
rect 3492 6379 3558 6395
rect 3912 6429 3978 6445
rect 3912 6395 3928 6429
rect 3962 6395 3978 6429
rect 3510 6357 3540 6379
rect 3720 6357 3750 6383
rect 3912 6379 3978 6395
rect 4332 6429 4398 6445
rect 4332 6395 4348 6429
rect 4382 6395 4398 6429
rect 3930 6357 3960 6379
rect 4140 6357 4170 6383
rect 4332 6379 4398 6395
rect 4752 6429 4818 6445
rect 4752 6395 4768 6429
rect 4802 6395 4818 6429
rect 4350 6357 4380 6379
rect 4560 6357 4590 6383
rect 4752 6379 4818 6395
rect 5172 6429 5238 6445
rect 5172 6395 5188 6429
rect 5222 6395 5238 6429
rect 4770 6357 4800 6379
rect 4980 6357 5010 6383
rect 5172 6379 5238 6395
rect 5592 6429 5658 6445
rect 5592 6395 5608 6429
rect 5642 6395 5658 6429
rect 5190 6357 5220 6379
rect 5400 6357 5430 6383
rect 5592 6379 5658 6395
rect 6012 6429 6078 6445
rect 6012 6395 6028 6429
rect 6062 6395 6078 6429
rect 5610 6357 5640 6379
rect 5820 6357 5850 6383
rect 6012 6379 6078 6395
rect 6030 6357 6060 6379
rect -2580 6135 -2550 6157
rect -2598 6119 -2532 6135
rect -2370 6131 -2340 6157
rect -2160 6135 -2130 6157
rect -2598 6085 -2582 6119
rect -2548 6085 -2532 6119
rect -2598 6069 -2532 6085
rect -2178 6119 -2112 6135
rect -1950 6131 -1920 6157
rect -1740 6135 -1710 6157
rect -2178 6085 -2162 6119
rect -2128 6085 -2112 6119
rect -2178 6069 -2112 6085
rect -1758 6119 -1692 6135
rect -1530 6131 -1500 6157
rect -1320 6135 -1290 6157
rect -1758 6085 -1742 6119
rect -1708 6085 -1692 6119
rect -1758 6069 -1692 6085
rect -1338 6119 -1272 6135
rect -1110 6131 -1080 6157
rect -900 6135 -870 6157
rect -1338 6085 -1322 6119
rect -1288 6085 -1272 6119
rect -1338 6069 -1272 6085
rect -918 6119 -852 6135
rect -690 6131 -660 6157
rect -480 6135 -450 6157
rect -918 6085 -902 6119
rect -868 6085 -852 6119
rect -918 6069 -852 6085
rect -498 6119 -432 6135
rect -270 6131 -240 6157
rect -60 6135 -30 6157
rect -498 6085 -482 6119
rect -448 6085 -432 6119
rect -498 6069 -432 6085
rect -78 6119 -12 6135
rect 150 6131 180 6157
rect 360 6135 390 6157
rect -78 6085 -62 6119
rect -28 6085 -12 6119
rect -78 6069 -12 6085
rect 342 6119 408 6135
rect 570 6131 600 6157
rect 780 6135 810 6157
rect 342 6085 358 6119
rect 392 6085 408 6119
rect 342 6069 408 6085
rect 762 6119 828 6135
rect 990 6131 1020 6157
rect 1200 6135 1230 6157
rect 762 6085 778 6119
rect 812 6085 828 6119
rect 762 6069 828 6085
rect 1182 6119 1248 6135
rect 1410 6131 1440 6157
rect 1620 6135 1650 6157
rect 1182 6085 1198 6119
rect 1232 6085 1248 6119
rect 1182 6069 1248 6085
rect 1602 6119 1668 6135
rect 1830 6131 1860 6157
rect 2040 6135 2070 6157
rect 1602 6085 1618 6119
rect 1652 6085 1668 6119
rect 1602 6069 1668 6085
rect 2022 6119 2088 6135
rect 2250 6131 2280 6157
rect 2460 6135 2490 6157
rect 2022 6085 2038 6119
rect 2072 6085 2088 6119
rect 2022 6069 2088 6085
rect 2442 6119 2508 6135
rect 2670 6131 2700 6157
rect 2880 6135 2910 6157
rect 2442 6085 2458 6119
rect 2492 6085 2508 6119
rect 2442 6069 2508 6085
rect 2862 6119 2928 6135
rect 3090 6131 3120 6157
rect 3300 6135 3330 6157
rect 2862 6085 2878 6119
rect 2912 6085 2928 6119
rect 2862 6069 2928 6085
rect 3282 6119 3348 6135
rect 3510 6131 3540 6157
rect 3720 6135 3750 6157
rect 3282 6085 3298 6119
rect 3332 6085 3348 6119
rect 3282 6069 3348 6085
rect 3702 6119 3768 6135
rect 3930 6131 3960 6157
rect 4140 6135 4170 6157
rect 3702 6085 3718 6119
rect 3752 6085 3768 6119
rect 3702 6069 3768 6085
rect 4122 6119 4188 6135
rect 4350 6131 4380 6157
rect 4560 6135 4590 6157
rect 4122 6085 4138 6119
rect 4172 6085 4188 6119
rect 4122 6069 4188 6085
rect 4542 6119 4608 6135
rect 4770 6131 4800 6157
rect 4980 6135 5010 6157
rect 4542 6085 4558 6119
rect 4592 6085 4608 6119
rect 4542 6069 4608 6085
rect 4962 6119 5028 6135
rect 5190 6131 5220 6157
rect 5400 6135 5430 6157
rect 4962 6085 4978 6119
rect 5012 6085 5028 6119
rect 4962 6069 5028 6085
rect 5382 6119 5448 6135
rect 5610 6131 5640 6157
rect 5820 6135 5850 6157
rect 5382 6085 5398 6119
rect 5432 6085 5448 6119
rect 5382 6069 5448 6085
rect 5802 6119 5868 6135
rect 6030 6131 6060 6157
rect 5802 6085 5818 6119
rect 5852 6085 5868 6119
rect 5802 6069 5868 6085
rect -2388 5989 -2322 6005
rect -2388 5955 -2372 5989
rect -2338 5955 -2322 5989
rect -2580 5917 -2550 5943
rect -2388 5939 -2322 5955
rect -1968 5989 -1902 6005
rect -1968 5955 -1952 5989
rect -1918 5955 -1902 5989
rect -2370 5917 -2340 5939
rect -2160 5917 -2130 5943
rect -1968 5939 -1902 5955
rect -1548 5989 -1482 6005
rect -1548 5955 -1532 5989
rect -1498 5955 -1482 5989
rect -1950 5917 -1920 5939
rect -1740 5917 -1710 5943
rect -1548 5939 -1482 5955
rect -1128 5989 -1062 6005
rect -1128 5955 -1112 5989
rect -1078 5955 -1062 5989
rect -1530 5917 -1500 5939
rect -1320 5917 -1290 5943
rect -1128 5939 -1062 5955
rect -708 5989 -642 6005
rect -708 5955 -692 5989
rect -658 5955 -642 5989
rect -1110 5917 -1080 5939
rect -900 5917 -870 5943
rect -708 5939 -642 5955
rect -288 5989 -222 6005
rect -288 5955 -272 5989
rect -238 5955 -222 5989
rect -690 5917 -660 5939
rect -480 5917 -450 5943
rect -288 5939 -222 5955
rect 132 5989 198 6005
rect 132 5955 148 5989
rect 182 5955 198 5989
rect -270 5917 -240 5939
rect -60 5917 -30 5943
rect 132 5939 198 5955
rect 552 5989 618 6005
rect 552 5955 568 5989
rect 602 5955 618 5989
rect 150 5917 180 5939
rect 360 5917 390 5943
rect 552 5939 618 5955
rect 972 5989 1038 6005
rect 972 5955 988 5989
rect 1022 5955 1038 5989
rect 570 5917 600 5939
rect 780 5917 810 5943
rect 972 5939 1038 5955
rect 1392 5989 1458 6005
rect 1392 5955 1408 5989
rect 1442 5955 1458 5989
rect 990 5917 1020 5939
rect 1200 5917 1230 5943
rect 1392 5939 1458 5955
rect 1812 5989 1878 6005
rect 1812 5955 1828 5989
rect 1862 5955 1878 5989
rect 1410 5917 1440 5939
rect 1620 5917 1650 5943
rect 1812 5939 1878 5955
rect 2232 5989 2298 6005
rect 2232 5955 2248 5989
rect 2282 5955 2298 5989
rect 1830 5917 1860 5939
rect 2040 5917 2070 5943
rect 2232 5939 2298 5955
rect 2652 5989 2718 6005
rect 2652 5955 2668 5989
rect 2702 5955 2718 5989
rect 2250 5917 2280 5939
rect 2460 5917 2490 5943
rect 2652 5939 2718 5955
rect 3072 5989 3138 6005
rect 3072 5955 3088 5989
rect 3122 5955 3138 5989
rect 2670 5917 2700 5939
rect 2880 5917 2910 5943
rect 3072 5939 3138 5955
rect 3492 5989 3558 6005
rect 3492 5955 3508 5989
rect 3542 5955 3558 5989
rect 3090 5917 3120 5939
rect 3300 5917 3330 5943
rect 3492 5939 3558 5955
rect 3912 5989 3978 6005
rect 3912 5955 3928 5989
rect 3962 5955 3978 5989
rect 3510 5917 3540 5939
rect 3720 5917 3750 5943
rect 3912 5939 3978 5955
rect 4332 5989 4398 6005
rect 4332 5955 4348 5989
rect 4382 5955 4398 5989
rect 3930 5917 3960 5939
rect 4140 5917 4170 5943
rect 4332 5939 4398 5955
rect 4752 5989 4818 6005
rect 4752 5955 4768 5989
rect 4802 5955 4818 5989
rect 4350 5917 4380 5939
rect 4560 5917 4590 5943
rect 4752 5939 4818 5955
rect 5172 5989 5238 6005
rect 5172 5955 5188 5989
rect 5222 5955 5238 5989
rect 4770 5917 4800 5939
rect 4980 5917 5010 5943
rect 5172 5939 5238 5955
rect 5592 5989 5658 6005
rect 5592 5955 5608 5989
rect 5642 5955 5658 5989
rect 5190 5917 5220 5939
rect 5400 5917 5430 5943
rect 5592 5939 5658 5955
rect 6012 5989 6078 6005
rect 6012 5955 6028 5989
rect 6062 5955 6078 5989
rect 5610 5917 5640 5939
rect 5820 5917 5850 5943
rect 6012 5939 6078 5955
rect 6030 5917 6060 5939
rect -2580 5695 -2550 5717
rect -2598 5679 -2532 5695
rect -2370 5691 -2340 5717
rect -2160 5695 -2130 5717
rect -2598 5645 -2582 5679
rect -2548 5645 -2532 5679
rect -2598 5629 -2532 5645
rect -2178 5679 -2112 5695
rect -1950 5691 -1920 5717
rect -1740 5695 -1710 5717
rect -2178 5645 -2162 5679
rect -2128 5645 -2112 5679
rect -2178 5629 -2112 5645
rect -1758 5679 -1692 5695
rect -1530 5691 -1500 5717
rect -1320 5695 -1290 5717
rect -1758 5645 -1742 5679
rect -1708 5645 -1692 5679
rect -1758 5629 -1692 5645
rect -1338 5679 -1272 5695
rect -1110 5691 -1080 5717
rect -900 5695 -870 5717
rect -1338 5645 -1322 5679
rect -1288 5645 -1272 5679
rect -1338 5629 -1272 5645
rect -918 5679 -852 5695
rect -690 5691 -660 5717
rect -480 5695 -450 5717
rect -918 5645 -902 5679
rect -868 5645 -852 5679
rect -918 5629 -852 5645
rect -498 5679 -432 5695
rect -270 5691 -240 5717
rect -60 5695 -30 5717
rect -498 5645 -482 5679
rect -448 5645 -432 5679
rect -498 5629 -432 5645
rect -78 5679 -12 5695
rect 150 5691 180 5717
rect 360 5695 390 5717
rect -78 5645 -62 5679
rect -28 5645 -12 5679
rect -78 5629 -12 5645
rect 342 5679 408 5695
rect 570 5691 600 5717
rect 780 5695 810 5717
rect 342 5645 358 5679
rect 392 5645 408 5679
rect 342 5629 408 5645
rect 762 5679 828 5695
rect 990 5691 1020 5717
rect 1200 5695 1230 5717
rect 762 5645 778 5679
rect 812 5645 828 5679
rect 762 5629 828 5645
rect 1182 5679 1248 5695
rect 1410 5691 1440 5717
rect 1620 5695 1650 5717
rect 1182 5645 1198 5679
rect 1232 5645 1248 5679
rect 1182 5629 1248 5645
rect 1602 5679 1668 5695
rect 1830 5691 1860 5717
rect 2040 5695 2070 5717
rect 1602 5645 1618 5679
rect 1652 5645 1668 5679
rect 1602 5629 1668 5645
rect 2022 5679 2088 5695
rect 2250 5691 2280 5717
rect 2460 5695 2490 5717
rect 2022 5645 2038 5679
rect 2072 5645 2088 5679
rect 2022 5629 2088 5645
rect 2442 5679 2508 5695
rect 2670 5691 2700 5717
rect 2880 5695 2910 5717
rect 2442 5645 2458 5679
rect 2492 5645 2508 5679
rect 2442 5629 2508 5645
rect 2862 5679 2928 5695
rect 3090 5691 3120 5717
rect 3300 5695 3330 5717
rect 2862 5645 2878 5679
rect 2912 5645 2928 5679
rect 2862 5629 2928 5645
rect 3282 5679 3348 5695
rect 3510 5691 3540 5717
rect 3720 5695 3750 5717
rect 3282 5645 3298 5679
rect 3332 5645 3348 5679
rect 3282 5629 3348 5645
rect 3702 5679 3768 5695
rect 3930 5691 3960 5717
rect 4140 5695 4170 5717
rect 3702 5645 3718 5679
rect 3752 5645 3768 5679
rect 3702 5629 3768 5645
rect 4122 5679 4188 5695
rect 4350 5691 4380 5717
rect 4560 5695 4590 5717
rect 4122 5645 4138 5679
rect 4172 5645 4188 5679
rect 4122 5629 4188 5645
rect 4542 5679 4608 5695
rect 4770 5691 4800 5717
rect 4980 5695 5010 5717
rect 4542 5645 4558 5679
rect 4592 5645 4608 5679
rect 4542 5629 4608 5645
rect 4962 5679 5028 5695
rect 5190 5691 5220 5717
rect 5400 5695 5430 5717
rect 4962 5645 4978 5679
rect 5012 5645 5028 5679
rect 4962 5629 5028 5645
rect 5382 5679 5448 5695
rect 5610 5691 5640 5717
rect 5820 5695 5850 5717
rect 5382 5645 5398 5679
rect 5432 5645 5448 5679
rect 5382 5629 5448 5645
rect 5802 5679 5868 5695
rect 6030 5691 6060 5717
rect 5802 5645 5818 5679
rect 5852 5645 5868 5679
rect 5802 5629 5868 5645
rect -2388 5549 -2322 5565
rect -2388 5515 -2372 5549
rect -2338 5515 -2322 5549
rect -2580 5477 -2550 5503
rect -2388 5499 -2322 5515
rect -1968 5549 -1902 5565
rect -1968 5515 -1952 5549
rect -1918 5515 -1902 5549
rect -2370 5477 -2340 5499
rect -2160 5477 -2130 5503
rect -1968 5499 -1902 5515
rect -1548 5549 -1482 5565
rect -1548 5515 -1532 5549
rect -1498 5515 -1482 5549
rect -1950 5477 -1920 5499
rect -1740 5477 -1710 5503
rect -1548 5499 -1482 5515
rect -1128 5549 -1062 5565
rect -1128 5515 -1112 5549
rect -1078 5515 -1062 5549
rect -1530 5477 -1500 5499
rect -1320 5477 -1290 5503
rect -1128 5499 -1062 5515
rect -708 5549 -642 5565
rect -708 5515 -692 5549
rect -658 5515 -642 5549
rect -1110 5477 -1080 5499
rect -900 5477 -870 5503
rect -708 5499 -642 5515
rect -288 5549 -222 5565
rect -288 5515 -272 5549
rect -238 5515 -222 5549
rect -690 5477 -660 5499
rect -480 5477 -450 5503
rect -288 5499 -222 5515
rect 132 5549 198 5565
rect 132 5515 148 5549
rect 182 5515 198 5549
rect -270 5477 -240 5499
rect -60 5477 -30 5503
rect 132 5499 198 5515
rect 552 5549 618 5565
rect 552 5515 568 5549
rect 602 5515 618 5549
rect 150 5477 180 5499
rect 360 5477 390 5503
rect 552 5499 618 5515
rect 972 5549 1038 5565
rect 972 5515 988 5549
rect 1022 5515 1038 5549
rect 570 5477 600 5499
rect 780 5477 810 5503
rect 972 5499 1038 5515
rect 1392 5549 1458 5565
rect 1392 5515 1408 5549
rect 1442 5515 1458 5549
rect 990 5477 1020 5499
rect 1200 5477 1230 5503
rect 1392 5499 1458 5515
rect 1812 5549 1878 5565
rect 1812 5515 1828 5549
rect 1862 5515 1878 5549
rect 1410 5477 1440 5499
rect 1620 5477 1650 5503
rect 1812 5499 1878 5515
rect 2232 5549 2298 5565
rect 2232 5515 2248 5549
rect 2282 5515 2298 5549
rect 1830 5477 1860 5499
rect 2040 5477 2070 5503
rect 2232 5499 2298 5515
rect 2652 5549 2718 5565
rect 2652 5515 2668 5549
rect 2702 5515 2718 5549
rect 2250 5477 2280 5499
rect 2460 5477 2490 5503
rect 2652 5499 2718 5515
rect 3072 5549 3138 5565
rect 3072 5515 3088 5549
rect 3122 5515 3138 5549
rect 2670 5477 2700 5499
rect 2880 5477 2910 5503
rect 3072 5499 3138 5515
rect 3492 5549 3558 5565
rect 3492 5515 3508 5549
rect 3542 5515 3558 5549
rect 3090 5477 3120 5499
rect 3300 5477 3330 5503
rect 3492 5499 3558 5515
rect 3912 5549 3978 5565
rect 3912 5515 3928 5549
rect 3962 5515 3978 5549
rect 3510 5477 3540 5499
rect 3720 5477 3750 5503
rect 3912 5499 3978 5515
rect 4332 5549 4398 5565
rect 4332 5515 4348 5549
rect 4382 5515 4398 5549
rect 3930 5477 3960 5499
rect 4140 5477 4170 5503
rect 4332 5499 4398 5515
rect 4752 5549 4818 5565
rect 4752 5515 4768 5549
rect 4802 5515 4818 5549
rect 4350 5477 4380 5499
rect 4560 5477 4590 5503
rect 4752 5499 4818 5515
rect 5172 5549 5238 5565
rect 5172 5515 5188 5549
rect 5222 5515 5238 5549
rect 4770 5477 4800 5499
rect 4980 5477 5010 5503
rect 5172 5499 5238 5515
rect 5592 5549 5658 5565
rect 5592 5515 5608 5549
rect 5642 5515 5658 5549
rect 5190 5477 5220 5499
rect 5400 5477 5430 5503
rect 5592 5499 5658 5515
rect 6012 5549 6078 5565
rect 6012 5515 6028 5549
rect 6062 5515 6078 5549
rect 5610 5477 5640 5499
rect 5820 5477 5850 5503
rect 6012 5499 6078 5515
rect 6030 5477 6060 5499
rect -2580 5255 -2550 5277
rect -2598 5239 -2532 5255
rect -2370 5251 -2340 5277
rect -2160 5255 -2130 5277
rect -2598 5205 -2582 5239
rect -2548 5205 -2532 5239
rect -2598 5189 -2532 5205
rect -2178 5239 -2112 5255
rect -1950 5251 -1920 5277
rect -1740 5255 -1710 5277
rect -2178 5205 -2162 5239
rect -2128 5205 -2112 5239
rect -2178 5189 -2112 5205
rect -1758 5239 -1692 5255
rect -1530 5251 -1500 5277
rect -1320 5255 -1290 5277
rect -1758 5205 -1742 5239
rect -1708 5205 -1692 5239
rect -1758 5189 -1692 5205
rect -1338 5239 -1272 5255
rect -1110 5251 -1080 5277
rect -900 5255 -870 5277
rect -1338 5205 -1322 5239
rect -1288 5205 -1272 5239
rect -1338 5189 -1272 5205
rect -918 5239 -852 5255
rect -690 5251 -660 5277
rect -480 5255 -450 5277
rect -918 5205 -902 5239
rect -868 5205 -852 5239
rect -918 5189 -852 5205
rect -498 5239 -432 5255
rect -270 5251 -240 5277
rect -60 5255 -30 5277
rect -498 5205 -482 5239
rect -448 5205 -432 5239
rect -498 5189 -432 5205
rect -78 5239 -12 5255
rect 150 5251 180 5277
rect 360 5255 390 5277
rect -78 5205 -62 5239
rect -28 5205 -12 5239
rect -78 5189 -12 5205
rect 342 5239 408 5255
rect 570 5251 600 5277
rect 780 5255 810 5277
rect 342 5205 358 5239
rect 392 5205 408 5239
rect 342 5189 408 5205
rect 762 5239 828 5255
rect 990 5251 1020 5277
rect 1200 5255 1230 5277
rect 762 5205 778 5239
rect 812 5205 828 5239
rect 762 5189 828 5205
rect 1182 5239 1248 5255
rect 1410 5251 1440 5277
rect 1620 5255 1650 5277
rect 1182 5205 1198 5239
rect 1232 5205 1248 5239
rect 1182 5189 1248 5205
rect 1602 5239 1668 5255
rect 1830 5251 1860 5277
rect 2040 5255 2070 5277
rect 1602 5205 1618 5239
rect 1652 5205 1668 5239
rect 1602 5189 1668 5205
rect 2022 5239 2088 5255
rect 2250 5251 2280 5277
rect 2460 5255 2490 5277
rect 2022 5205 2038 5239
rect 2072 5205 2088 5239
rect 2022 5189 2088 5205
rect 2442 5239 2508 5255
rect 2670 5251 2700 5277
rect 2880 5255 2910 5277
rect 2442 5205 2458 5239
rect 2492 5205 2508 5239
rect 2442 5189 2508 5205
rect 2862 5239 2928 5255
rect 3090 5251 3120 5277
rect 3300 5255 3330 5277
rect 2862 5205 2878 5239
rect 2912 5205 2928 5239
rect 2862 5189 2928 5205
rect 3282 5239 3348 5255
rect 3510 5251 3540 5277
rect 3720 5255 3750 5277
rect 3282 5205 3298 5239
rect 3332 5205 3348 5239
rect 3282 5189 3348 5205
rect 3702 5239 3768 5255
rect 3930 5251 3960 5277
rect 4140 5255 4170 5277
rect 3702 5205 3718 5239
rect 3752 5205 3768 5239
rect 3702 5189 3768 5205
rect 4122 5239 4188 5255
rect 4350 5251 4380 5277
rect 4560 5255 4590 5277
rect 4122 5205 4138 5239
rect 4172 5205 4188 5239
rect 4122 5189 4188 5205
rect 4542 5239 4608 5255
rect 4770 5251 4800 5277
rect 4980 5255 5010 5277
rect 4542 5205 4558 5239
rect 4592 5205 4608 5239
rect 4542 5189 4608 5205
rect 4962 5239 5028 5255
rect 5190 5251 5220 5277
rect 5400 5255 5430 5277
rect 4962 5205 4978 5239
rect 5012 5205 5028 5239
rect 4962 5189 5028 5205
rect 5382 5239 5448 5255
rect 5610 5251 5640 5277
rect 5820 5255 5850 5277
rect 5382 5205 5398 5239
rect 5432 5205 5448 5239
rect 5382 5189 5448 5205
rect 5802 5239 5868 5255
rect 6030 5251 6060 5277
rect 5802 5205 5818 5239
rect 5852 5205 5868 5239
rect 5802 5189 5868 5205
rect -2388 5109 -2322 5125
rect -2388 5075 -2372 5109
rect -2338 5075 -2322 5109
rect -2580 5037 -2550 5063
rect -2388 5059 -2322 5075
rect -1968 5109 -1902 5125
rect -1968 5075 -1952 5109
rect -1918 5075 -1902 5109
rect -2370 5037 -2340 5059
rect -2160 5037 -2130 5063
rect -1968 5059 -1902 5075
rect -1548 5109 -1482 5125
rect -1548 5075 -1532 5109
rect -1498 5075 -1482 5109
rect -1950 5037 -1920 5059
rect -1740 5037 -1710 5063
rect -1548 5059 -1482 5075
rect -1128 5109 -1062 5125
rect -1128 5075 -1112 5109
rect -1078 5075 -1062 5109
rect -1530 5037 -1500 5059
rect -1320 5037 -1290 5063
rect -1128 5059 -1062 5075
rect -708 5109 -642 5125
rect -708 5075 -692 5109
rect -658 5075 -642 5109
rect -1110 5037 -1080 5059
rect -900 5037 -870 5063
rect -708 5059 -642 5075
rect -288 5109 -222 5125
rect -288 5075 -272 5109
rect -238 5075 -222 5109
rect -690 5037 -660 5059
rect -480 5037 -450 5063
rect -288 5059 -222 5075
rect 132 5109 198 5125
rect 132 5075 148 5109
rect 182 5075 198 5109
rect -270 5037 -240 5059
rect -60 5037 -30 5063
rect 132 5059 198 5075
rect 552 5109 618 5125
rect 552 5075 568 5109
rect 602 5075 618 5109
rect 150 5037 180 5059
rect 360 5037 390 5063
rect 552 5059 618 5075
rect 972 5109 1038 5125
rect 972 5075 988 5109
rect 1022 5075 1038 5109
rect 570 5037 600 5059
rect 780 5037 810 5063
rect 972 5059 1038 5075
rect 1392 5109 1458 5125
rect 1392 5075 1408 5109
rect 1442 5075 1458 5109
rect 990 5037 1020 5059
rect 1200 5037 1230 5063
rect 1392 5059 1458 5075
rect 1812 5109 1878 5125
rect 1812 5075 1828 5109
rect 1862 5075 1878 5109
rect 1410 5037 1440 5059
rect 1620 5037 1650 5063
rect 1812 5059 1878 5075
rect 2232 5109 2298 5125
rect 2232 5075 2248 5109
rect 2282 5075 2298 5109
rect 1830 5037 1860 5059
rect 2040 5037 2070 5063
rect 2232 5059 2298 5075
rect 2652 5109 2718 5125
rect 2652 5075 2668 5109
rect 2702 5075 2718 5109
rect 2250 5037 2280 5059
rect 2460 5037 2490 5063
rect 2652 5059 2718 5075
rect 3072 5109 3138 5125
rect 3072 5075 3088 5109
rect 3122 5075 3138 5109
rect 2670 5037 2700 5059
rect 2880 5037 2910 5063
rect 3072 5059 3138 5075
rect 3492 5109 3558 5125
rect 3492 5075 3508 5109
rect 3542 5075 3558 5109
rect 3090 5037 3120 5059
rect 3300 5037 3330 5063
rect 3492 5059 3558 5075
rect 3912 5109 3978 5125
rect 3912 5075 3928 5109
rect 3962 5075 3978 5109
rect 3510 5037 3540 5059
rect 3720 5037 3750 5063
rect 3912 5059 3978 5075
rect 4332 5109 4398 5125
rect 4332 5075 4348 5109
rect 4382 5075 4398 5109
rect 3930 5037 3960 5059
rect 4140 5037 4170 5063
rect 4332 5059 4398 5075
rect 4752 5109 4818 5125
rect 4752 5075 4768 5109
rect 4802 5075 4818 5109
rect 4350 5037 4380 5059
rect 4560 5037 4590 5063
rect 4752 5059 4818 5075
rect 5172 5109 5238 5125
rect 5172 5075 5188 5109
rect 5222 5075 5238 5109
rect 4770 5037 4800 5059
rect 4980 5037 5010 5063
rect 5172 5059 5238 5075
rect 5592 5109 5658 5125
rect 5592 5075 5608 5109
rect 5642 5075 5658 5109
rect 5190 5037 5220 5059
rect 5400 5037 5430 5063
rect 5592 5059 5658 5075
rect 6012 5109 6078 5125
rect 6012 5075 6028 5109
rect 6062 5075 6078 5109
rect 5610 5037 5640 5059
rect 5820 5037 5850 5063
rect 6012 5059 6078 5075
rect 6030 5037 6060 5059
rect -2580 4815 -2550 4837
rect -2598 4799 -2532 4815
rect -2370 4811 -2340 4837
rect -2160 4815 -2130 4837
rect -2598 4765 -2582 4799
rect -2548 4765 -2532 4799
rect -2598 4749 -2532 4765
rect -2178 4799 -2112 4815
rect -1950 4811 -1920 4837
rect -1740 4815 -1710 4837
rect -2178 4765 -2162 4799
rect -2128 4765 -2112 4799
rect -2178 4749 -2112 4765
rect -1758 4799 -1692 4815
rect -1530 4811 -1500 4837
rect -1320 4815 -1290 4837
rect -1758 4765 -1742 4799
rect -1708 4765 -1692 4799
rect -1758 4749 -1692 4765
rect -1338 4799 -1272 4815
rect -1110 4811 -1080 4837
rect -900 4815 -870 4837
rect -1338 4765 -1322 4799
rect -1288 4765 -1272 4799
rect -1338 4749 -1272 4765
rect -918 4799 -852 4815
rect -690 4811 -660 4837
rect -480 4815 -450 4837
rect -918 4765 -902 4799
rect -868 4765 -852 4799
rect -918 4749 -852 4765
rect -498 4799 -432 4815
rect -270 4811 -240 4837
rect -60 4815 -30 4837
rect -498 4765 -482 4799
rect -448 4765 -432 4799
rect -498 4749 -432 4765
rect -78 4799 -12 4815
rect 150 4811 180 4837
rect 360 4815 390 4837
rect -78 4765 -62 4799
rect -28 4765 -12 4799
rect -78 4749 -12 4765
rect 342 4799 408 4815
rect 570 4811 600 4837
rect 780 4815 810 4837
rect 342 4765 358 4799
rect 392 4765 408 4799
rect 342 4749 408 4765
rect 762 4799 828 4815
rect 990 4811 1020 4837
rect 1200 4815 1230 4837
rect 762 4765 778 4799
rect 812 4765 828 4799
rect 762 4749 828 4765
rect 1182 4799 1248 4815
rect 1410 4811 1440 4837
rect 1620 4815 1650 4837
rect 1182 4765 1198 4799
rect 1232 4765 1248 4799
rect 1182 4749 1248 4765
rect 1602 4799 1668 4815
rect 1830 4811 1860 4837
rect 2040 4815 2070 4837
rect 1602 4765 1618 4799
rect 1652 4765 1668 4799
rect 1602 4749 1668 4765
rect 2022 4799 2088 4815
rect 2250 4811 2280 4837
rect 2460 4815 2490 4837
rect 2022 4765 2038 4799
rect 2072 4765 2088 4799
rect 2022 4749 2088 4765
rect 2442 4799 2508 4815
rect 2670 4811 2700 4837
rect 2880 4815 2910 4837
rect 2442 4765 2458 4799
rect 2492 4765 2508 4799
rect 2442 4749 2508 4765
rect 2862 4799 2928 4815
rect 3090 4811 3120 4837
rect 3300 4815 3330 4837
rect 2862 4765 2878 4799
rect 2912 4765 2928 4799
rect 2862 4749 2928 4765
rect 3282 4799 3348 4815
rect 3510 4811 3540 4837
rect 3720 4815 3750 4837
rect 3282 4765 3298 4799
rect 3332 4765 3348 4799
rect 3282 4749 3348 4765
rect 3702 4799 3768 4815
rect 3930 4811 3960 4837
rect 4140 4815 4170 4837
rect 3702 4765 3718 4799
rect 3752 4765 3768 4799
rect 3702 4749 3768 4765
rect 4122 4799 4188 4815
rect 4350 4811 4380 4837
rect 4560 4815 4590 4837
rect 4122 4765 4138 4799
rect 4172 4765 4188 4799
rect 4122 4749 4188 4765
rect 4542 4799 4608 4815
rect 4770 4811 4800 4837
rect 4980 4815 5010 4837
rect 4542 4765 4558 4799
rect 4592 4765 4608 4799
rect 4542 4749 4608 4765
rect 4962 4799 5028 4815
rect 5190 4811 5220 4837
rect 5400 4815 5430 4837
rect 4962 4765 4978 4799
rect 5012 4765 5028 4799
rect 4962 4749 5028 4765
rect 5382 4799 5448 4815
rect 5610 4811 5640 4837
rect 5820 4815 5850 4837
rect 5382 4765 5398 4799
rect 5432 4765 5448 4799
rect 5382 4749 5448 4765
rect 5802 4799 5868 4815
rect 6030 4811 6060 4837
rect 5802 4765 5818 4799
rect 5852 4765 5868 4799
rect 5802 4749 5868 4765
rect 7062 7862 7128 7878
rect 7062 7860 7078 7862
rect 6804 7830 6831 7860
rect 7031 7830 7078 7860
rect 6734 7766 6800 7782
rect 6734 7732 6750 7766
rect 6784 7764 6800 7766
rect 7062 7828 7078 7830
rect 7112 7828 7128 7862
rect 7062 7812 7128 7828
rect 6784 7734 6831 7764
rect 7031 7734 7058 7764
rect 6784 7732 6800 7734
rect 6734 7716 6800 7732
rect 7062 7670 7128 7686
rect 7062 7668 7078 7670
rect 6804 7638 6831 7668
rect 7031 7638 7078 7668
rect 6734 7574 6800 7590
rect 6734 7540 6750 7574
rect 6784 7572 6800 7574
rect 7062 7636 7078 7638
rect 7112 7636 7128 7670
rect 7062 7620 7128 7636
rect 6784 7542 6831 7572
rect 7031 7542 7058 7572
rect 6784 7540 6800 7542
rect 6734 7524 6800 7540
rect 7062 7478 7128 7494
rect 7062 7476 7078 7478
rect 6804 7446 6831 7476
rect 7031 7446 7078 7476
rect 6734 7382 6800 7398
rect 6734 7348 6750 7382
rect 6784 7380 6800 7382
rect 7062 7444 7078 7446
rect 7112 7444 7128 7478
rect 7062 7428 7128 7444
rect 6784 7350 6831 7380
rect 7031 7350 7058 7380
rect 6784 7348 6800 7350
rect 6734 7332 6800 7348
rect 7062 7286 7128 7302
rect 7062 7284 7078 7286
rect 6804 7254 6831 7284
rect 7031 7254 7078 7284
rect 6734 7190 6800 7206
rect 6734 7156 6750 7190
rect 6784 7188 6800 7190
rect 7062 7252 7078 7254
rect 7112 7252 7128 7286
rect 7062 7236 7128 7252
rect 6784 7158 6831 7188
rect 7031 7158 7058 7188
rect 6784 7156 6800 7158
rect 6734 7140 6800 7156
rect 7062 7094 7128 7110
rect 7062 7092 7078 7094
rect 6804 7062 6831 7092
rect 7031 7062 7078 7092
rect 6734 6998 6800 7014
rect 6734 6964 6750 6998
rect 6784 6996 6800 6998
rect 7062 7060 7078 7062
rect 7112 7060 7128 7094
rect 7062 7044 7128 7060
rect 6784 6966 6831 6996
rect 7031 6966 7058 6996
rect 6784 6964 6800 6966
rect 6734 6948 6800 6964
rect 7062 6902 7128 6918
rect 7062 6900 7078 6902
rect 6804 6870 6831 6900
rect 7031 6870 7078 6900
rect 6734 6806 6800 6822
rect 6734 6772 6750 6806
rect 6784 6804 6800 6806
rect 7062 6868 7078 6870
rect 7112 6868 7128 6902
rect 7062 6852 7128 6868
rect 6784 6774 6831 6804
rect 7031 6774 7058 6804
rect 6784 6772 6800 6774
rect 6734 6756 6800 6772
rect 7062 6710 7128 6726
rect 7062 6708 7078 6710
rect 6804 6678 6831 6708
rect 7031 6678 7078 6708
rect 6734 6614 6800 6630
rect 6734 6580 6750 6614
rect 6784 6612 6800 6614
rect 7062 6676 7078 6678
rect 7112 6676 7128 6710
rect 7062 6660 7128 6676
rect 6784 6582 6831 6612
rect 7031 6582 7058 6612
rect 6784 6580 6800 6582
rect 6734 6564 6800 6580
rect 7062 6518 7128 6534
rect 7062 6516 7078 6518
rect 6804 6486 6831 6516
rect 7031 6486 7078 6516
rect 6734 6422 6800 6438
rect 6734 6388 6750 6422
rect 6784 6420 6800 6422
rect 7062 6484 7078 6486
rect 7112 6484 7128 6518
rect 7062 6468 7128 6484
rect 6784 6390 6831 6420
rect 7031 6390 7058 6420
rect 6784 6388 6800 6390
rect 6734 6372 6800 6388
rect 7062 6326 7128 6342
rect 7062 6324 7078 6326
rect 6804 6294 6831 6324
rect 7031 6294 7078 6324
rect 6734 6230 6800 6246
rect 6734 6196 6750 6230
rect 6784 6228 6800 6230
rect 7062 6292 7078 6294
rect 7112 6292 7128 6326
rect 7062 6276 7128 6292
rect 6784 6198 6831 6228
rect 7031 6198 7058 6228
rect 6784 6196 6800 6198
rect 6734 6180 6800 6196
rect -2388 4174 -2322 4190
rect -2388 4140 -2372 4174
rect -2338 4140 -2322 4174
rect -2580 4102 -2550 4128
rect -2388 4124 -2322 4140
rect -1968 4174 -1902 4190
rect -1968 4140 -1952 4174
rect -1918 4140 -1902 4174
rect -2370 4102 -2340 4124
rect -2160 4102 -2130 4128
rect -1968 4124 -1902 4140
rect -1548 4174 -1482 4190
rect -1548 4140 -1532 4174
rect -1498 4140 -1482 4174
rect -1950 4102 -1920 4124
rect -1740 4102 -1710 4128
rect -1548 4124 -1482 4140
rect -1128 4174 -1062 4190
rect -1128 4140 -1112 4174
rect -1078 4140 -1062 4174
rect -1530 4102 -1500 4124
rect -1320 4102 -1290 4128
rect -1128 4124 -1062 4140
rect -708 4174 -642 4190
rect -708 4140 -692 4174
rect -658 4140 -642 4174
rect -1110 4102 -1080 4124
rect -900 4102 -870 4128
rect -708 4124 -642 4140
rect -288 4174 -222 4190
rect -288 4140 -272 4174
rect -238 4140 -222 4174
rect -690 4102 -660 4124
rect -480 4102 -450 4128
rect -288 4124 -222 4140
rect 132 4174 198 4190
rect 132 4140 148 4174
rect 182 4140 198 4174
rect -270 4102 -240 4124
rect -60 4102 -30 4128
rect 132 4124 198 4140
rect 552 4174 618 4190
rect 552 4140 568 4174
rect 602 4140 618 4174
rect 150 4102 180 4124
rect 360 4102 390 4128
rect 552 4124 618 4140
rect 972 4174 1038 4190
rect 972 4140 988 4174
rect 1022 4140 1038 4174
rect 570 4102 600 4124
rect 780 4102 810 4128
rect 972 4124 1038 4140
rect 1392 4174 1458 4190
rect 1392 4140 1408 4174
rect 1442 4140 1458 4174
rect 990 4102 1020 4124
rect 1200 4102 1230 4128
rect 1392 4124 1458 4140
rect 1812 4174 1878 4190
rect 1812 4140 1828 4174
rect 1862 4140 1878 4174
rect 1410 4102 1440 4124
rect 1620 4102 1650 4128
rect 1812 4124 1878 4140
rect 2232 4174 2298 4190
rect 2232 4140 2248 4174
rect 2282 4140 2298 4174
rect 1830 4102 1860 4124
rect 2040 4102 2070 4128
rect 2232 4124 2298 4140
rect 2652 4174 2718 4190
rect 2652 4140 2668 4174
rect 2702 4140 2718 4174
rect 2250 4102 2280 4124
rect 2460 4102 2490 4128
rect 2652 4124 2718 4140
rect 3072 4174 3138 4190
rect 3072 4140 3088 4174
rect 3122 4140 3138 4174
rect 2670 4102 2700 4124
rect 2880 4102 2910 4128
rect 3072 4124 3138 4140
rect 3492 4174 3558 4190
rect 3492 4140 3508 4174
rect 3542 4140 3558 4174
rect 3090 4102 3120 4124
rect 3300 4102 3330 4128
rect 3492 4124 3558 4140
rect 3912 4174 3978 4190
rect 3912 4140 3928 4174
rect 3962 4140 3978 4174
rect 3510 4102 3540 4124
rect 3720 4102 3750 4128
rect 3912 4124 3978 4140
rect 4332 4174 4398 4190
rect 4332 4140 4348 4174
rect 4382 4140 4398 4174
rect 3930 4102 3960 4124
rect 4140 4102 4170 4128
rect 4332 4124 4398 4140
rect 4752 4174 4818 4190
rect 4752 4140 4768 4174
rect 4802 4140 4818 4174
rect 4350 4102 4380 4124
rect 4560 4102 4590 4128
rect 4752 4124 4818 4140
rect 5172 4174 5238 4190
rect 5172 4140 5188 4174
rect 5222 4140 5238 4174
rect 4770 4102 4800 4124
rect 4980 4102 5010 4128
rect 5172 4124 5238 4140
rect 5592 4174 5658 4190
rect 5592 4140 5608 4174
rect 5642 4140 5658 4174
rect 5190 4102 5220 4124
rect 5400 4102 5430 4128
rect 5592 4124 5658 4140
rect 6012 4174 6078 4190
rect 6012 4140 6028 4174
rect 6062 4140 6078 4174
rect 5610 4102 5640 4124
rect 5820 4102 5850 4128
rect 6012 4124 6078 4140
rect 6030 4102 6060 4124
rect -2580 3880 -2550 3902
rect -2598 3864 -2532 3880
rect -2370 3876 -2340 3902
rect -2160 3880 -2130 3902
rect -2598 3830 -2582 3864
rect -2548 3830 -2532 3864
rect -2598 3814 -2532 3830
rect -2178 3864 -2112 3880
rect -1950 3876 -1920 3902
rect -1740 3880 -1710 3902
rect -2178 3830 -2162 3864
rect -2128 3830 -2112 3864
rect -2178 3814 -2112 3830
rect -1758 3864 -1692 3880
rect -1530 3876 -1500 3902
rect -1320 3880 -1290 3902
rect -1758 3830 -1742 3864
rect -1708 3830 -1692 3864
rect -1758 3814 -1692 3830
rect -1338 3864 -1272 3880
rect -1110 3876 -1080 3902
rect -900 3880 -870 3902
rect -1338 3830 -1322 3864
rect -1288 3830 -1272 3864
rect -1338 3814 -1272 3830
rect -918 3864 -852 3880
rect -690 3876 -660 3902
rect -480 3880 -450 3902
rect -918 3830 -902 3864
rect -868 3830 -852 3864
rect -918 3814 -852 3830
rect -498 3864 -432 3880
rect -270 3876 -240 3902
rect -60 3880 -30 3902
rect -498 3830 -482 3864
rect -448 3830 -432 3864
rect -498 3814 -432 3830
rect -78 3864 -12 3880
rect 150 3876 180 3902
rect 360 3880 390 3902
rect -78 3830 -62 3864
rect -28 3830 -12 3864
rect -78 3814 -12 3830
rect 342 3864 408 3880
rect 570 3876 600 3902
rect 780 3880 810 3902
rect 342 3830 358 3864
rect 392 3830 408 3864
rect 342 3814 408 3830
rect 762 3864 828 3880
rect 990 3876 1020 3902
rect 1200 3880 1230 3902
rect 762 3830 778 3864
rect 812 3830 828 3864
rect 762 3814 828 3830
rect 1182 3864 1248 3880
rect 1410 3876 1440 3902
rect 1620 3880 1650 3902
rect 1182 3830 1198 3864
rect 1232 3830 1248 3864
rect 1182 3814 1248 3830
rect 1602 3864 1668 3880
rect 1830 3876 1860 3902
rect 2040 3880 2070 3902
rect 1602 3830 1618 3864
rect 1652 3830 1668 3864
rect 1602 3814 1668 3830
rect 2022 3864 2088 3880
rect 2250 3876 2280 3902
rect 2460 3880 2490 3902
rect 2022 3830 2038 3864
rect 2072 3830 2088 3864
rect 2022 3814 2088 3830
rect 2442 3864 2508 3880
rect 2670 3876 2700 3902
rect 2880 3880 2910 3902
rect 2442 3830 2458 3864
rect 2492 3830 2508 3864
rect 2442 3814 2508 3830
rect 2862 3864 2928 3880
rect 3090 3876 3120 3902
rect 3300 3880 3330 3902
rect 2862 3830 2878 3864
rect 2912 3830 2928 3864
rect 2862 3814 2928 3830
rect 3282 3864 3348 3880
rect 3510 3876 3540 3902
rect 3720 3880 3750 3902
rect 3282 3830 3298 3864
rect 3332 3830 3348 3864
rect 3282 3814 3348 3830
rect 3702 3864 3768 3880
rect 3930 3876 3960 3902
rect 4140 3880 4170 3902
rect 3702 3830 3718 3864
rect 3752 3830 3768 3864
rect 3702 3814 3768 3830
rect 4122 3864 4188 3880
rect 4350 3876 4380 3902
rect 4560 3880 4590 3902
rect 4122 3830 4138 3864
rect 4172 3830 4188 3864
rect 4122 3814 4188 3830
rect 4542 3864 4608 3880
rect 4770 3876 4800 3902
rect 4980 3880 5010 3902
rect 4542 3830 4558 3864
rect 4592 3830 4608 3864
rect 4542 3814 4608 3830
rect 4962 3864 5028 3880
rect 5190 3876 5220 3902
rect 5400 3880 5430 3902
rect 4962 3830 4978 3864
rect 5012 3830 5028 3864
rect 4962 3814 5028 3830
rect 5382 3864 5448 3880
rect 5610 3876 5640 3902
rect 5820 3880 5850 3902
rect 5382 3830 5398 3864
rect 5432 3830 5448 3864
rect 5382 3814 5448 3830
rect 5802 3864 5868 3880
rect 6030 3876 6060 3902
rect 5802 3830 5818 3864
rect 5852 3830 5868 3864
rect 5802 3814 5868 3830
rect -2388 3734 -2322 3750
rect -2388 3700 -2372 3734
rect -2338 3700 -2322 3734
rect -2580 3662 -2550 3688
rect -2388 3684 -2322 3700
rect -1968 3734 -1902 3750
rect -1968 3700 -1952 3734
rect -1918 3700 -1902 3734
rect -2370 3662 -2340 3684
rect -2160 3662 -2130 3688
rect -1968 3684 -1902 3700
rect -1548 3734 -1482 3750
rect -1548 3700 -1532 3734
rect -1498 3700 -1482 3734
rect -1950 3662 -1920 3684
rect -1740 3662 -1710 3688
rect -1548 3684 -1482 3700
rect -1128 3734 -1062 3750
rect -1128 3700 -1112 3734
rect -1078 3700 -1062 3734
rect -1530 3662 -1500 3684
rect -1320 3662 -1290 3688
rect -1128 3684 -1062 3700
rect -708 3734 -642 3750
rect -708 3700 -692 3734
rect -658 3700 -642 3734
rect -1110 3662 -1080 3684
rect -900 3662 -870 3688
rect -708 3684 -642 3700
rect -288 3734 -222 3750
rect -288 3700 -272 3734
rect -238 3700 -222 3734
rect -690 3662 -660 3684
rect -480 3662 -450 3688
rect -288 3684 -222 3700
rect 132 3734 198 3750
rect 132 3700 148 3734
rect 182 3700 198 3734
rect -270 3662 -240 3684
rect -60 3662 -30 3688
rect 132 3684 198 3700
rect 552 3734 618 3750
rect 552 3700 568 3734
rect 602 3700 618 3734
rect 150 3662 180 3684
rect 360 3662 390 3688
rect 552 3684 618 3700
rect 972 3734 1038 3750
rect 972 3700 988 3734
rect 1022 3700 1038 3734
rect 570 3662 600 3684
rect 780 3662 810 3688
rect 972 3684 1038 3700
rect 1392 3734 1458 3750
rect 1392 3700 1408 3734
rect 1442 3700 1458 3734
rect 990 3662 1020 3684
rect 1200 3662 1230 3688
rect 1392 3684 1458 3700
rect 1812 3734 1878 3750
rect 1812 3700 1828 3734
rect 1862 3700 1878 3734
rect 1410 3662 1440 3684
rect 1620 3662 1650 3688
rect 1812 3684 1878 3700
rect 2232 3734 2298 3750
rect 2232 3700 2248 3734
rect 2282 3700 2298 3734
rect 1830 3662 1860 3684
rect 2040 3662 2070 3688
rect 2232 3684 2298 3700
rect 2652 3734 2718 3750
rect 2652 3700 2668 3734
rect 2702 3700 2718 3734
rect 2250 3662 2280 3684
rect 2460 3662 2490 3688
rect 2652 3684 2718 3700
rect 3072 3734 3138 3750
rect 3072 3700 3088 3734
rect 3122 3700 3138 3734
rect 2670 3662 2700 3684
rect 2880 3662 2910 3688
rect 3072 3684 3138 3700
rect 3492 3734 3558 3750
rect 3492 3700 3508 3734
rect 3542 3700 3558 3734
rect 3090 3662 3120 3684
rect 3300 3662 3330 3688
rect 3492 3684 3558 3700
rect 3912 3734 3978 3750
rect 3912 3700 3928 3734
rect 3962 3700 3978 3734
rect 3510 3662 3540 3684
rect 3720 3662 3750 3688
rect 3912 3684 3978 3700
rect 4332 3734 4398 3750
rect 4332 3700 4348 3734
rect 4382 3700 4398 3734
rect 3930 3662 3960 3684
rect 4140 3662 4170 3688
rect 4332 3684 4398 3700
rect 4752 3734 4818 3750
rect 4752 3700 4768 3734
rect 4802 3700 4818 3734
rect 4350 3662 4380 3684
rect 4560 3662 4590 3688
rect 4752 3684 4818 3700
rect 5172 3734 5238 3750
rect 5172 3700 5188 3734
rect 5222 3700 5238 3734
rect 4770 3662 4800 3684
rect 4980 3662 5010 3688
rect 5172 3684 5238 3700
rect 5592 3734 5658 3750
rect 5592 3700 5608 3734
rect 5642 3700 5658 3734
rect 5190 3662 5220 3684
rect 5400 3662 5430 3688
rect 5592 3684 5658 3700
rect 6012 3734 6078 3750
rect 6012 3700 6028 3734
rect 6062 3700 6078 3734
rect 5610 3662 5640 3684
rect 5820 3662 5850 3688
rect 6012 3684 6078 3700
rect 6030 3662 6060 3684
rect -2580 3440 -2550 3462
rect -2598 3424 -2532 3440
rect -2370 3436 -2340 3462
rect -2160 3440 -2130 3462
rect -2598 3390 -2582 3424
rect -2548 3390 -2532 3424
rect -2598 3374 -2532 3390
rect -2178 3424 -2112 3440
rect -1950 3436 -1920 3462
rect -1740 3440 -1710 3462
rect -2178 3390 -2162 3424
rect -2128 3390 -2112 3424
rect -2178 3374 -2112 3390
rect -1758 3424 -1692 3440
rect -1530 3436 -1500 3462
rect -1320 3440 -1290 3462
rect -1758 3390 -1742 3424
rect -1708 3390 -1692 3424
rect -1758 3374 -1692 3390
rect -1338 3424 -1272 3440
rect -1110 3436 -1080 3462
rect -900 3440 -870 3462
rect -1338 3390 -1322 3424
rect -1288 3390 -1272 3424
rect -1338 3374 -1272 3390
rect -918 3424 -852 3440
rect -690 3436 -660 3462
rect -480 3440 -450 3462
rect -918 3390 -902 3424
rect -868 3390 -852 3424
rect -918 3374 -852 3390
rect -498 3424 -432 3440
rect -270 3436 -240 3462
rect -60 3440 -30 3462
rect -498 3390 -482 3424
rect -448 3390 -432 3424
rect -498 3374 -432 3390
rect -78 3424 -12 3440
rect 150 3436 180 3462
rect 360 3440 390 3462
rect -78 3390 -62 3424
rect -28 3390 -12 3424
rect -78 3374 -12 3390
rect 342 3424 408 3440
rect 570 3436 600 3462
rect 780 3440 810 3462
rect 342 3390 358 3424
rect 392 3390 408 3424
rect 342 3374 408 3390
rect 762 3424 828 3440
rect 990 3436 1020 3462
rect 1200 3440 1230 3462
rect 762 3390 778 3424
rect 812 3390 828 3424
rect 762 3374 828 3390
rect 1182 3424 1248 3440
rect 1410 3436 1440 3462
rect 1620 3440 1650 3462
rect 1182 3390 1198 3424
rect 1232 3390 1248 3424
rect 1182 3374 1248 3390
rect 1602 3424 1668 3440
rect 1830 3436 1860 3462
rect 2040 3440 2070 3462
rect 1602 3390 1618 3424
rect 1652 3390 1668 3424
rect 1602 3374 1668 3390
rect 2022 3424 2088 3440
rect 2250 3436 2280 3462
rect 2460 3440 2490 3462
rect 2022 3390 2038 3424
rect 2072 3390 2088 3424
rect 2022 3374 2088 3390
rect 2442 3424 2508 3440
rect 2670 3436 2700 3462
rect 2880 3440 2910 3462
rect 2442 3390 2458 3424
rect 2492 3390 2508 3424
rect 2442 3374 2508 3390
rect 2862 3424 2928 3440
rect 3090 3436 3120 3462
rect 3300 3440 3330 3462
rect 2862 3390 2878 3424
rect 2912 3390 2928 3424
rect 2862 3374 2928 3390
rect 3282 3424 3348 3440
rect 3510 3436 3540 3462
rect 3720 3440 3750 3462
rect 3282 3390 3298 3424
rect 3332 3390 3348 3424
rect 3282 3374 3348 3390
rect 3702 3424 3768 3440
rect 3930 3436 3960 3462
rect 4140 3440 4170 3462
rect 3702 3390 3718 3424
rect 3752 3390 3768 3424
rect 3702 3374 3768 3390
rect 4122 3424 4188 3440
rect 4350 3436 4380 3462
rect 4560 3440 4590 3462
rect 4122 3390 4138 3424
rect 4172 3390 4188 3424
rect 4122 3374 4188 3390
rect 4542 3424 4608 3440
rect 4770 3436 4800 3462
rect 4980 3440 5010 3462
rect 4542 3390 4558 3424
rect 4592 3390 4608 3424
rect 4542 3374 4608 3390
rect 4962 3424 5028 3440
rect 5190 3436 5220 3462
rect 5400 3440 5430 3462
rect 4962 3390 4978 3424
rect 5012 3390 5028 3424
rect 4962 3374 5028 3390
rect 5382 3424 5448 3440
rect 5610 3436 5640 3462
rect 5820 3440 5850 3462
rect 5382 3390 5398 3424
rect 5432 3390 5448 3424
rect 5382 3374 5448 3390
rect 5802 3424 5868 3440
rect 6030 3436 6060 3462
rect 5802 3390 5818 3424
rect 5852 3390 5868 3424
rect 5802 3374 5868 3390
rect -2388 3294 -2322 3310
rect -2388 3260 -2372 3294
rect -2338 3260 -2322 3294
rect -2580 3222 -2550 3248
rect -2388 3244 -2322 3260
rect -1968 3294 -1902 3310
rect -1968 3260 -1952 3294
rect -1918 3260 -1902 3294
rect -2370 3222 -2340 3244
rect -2160 3222 -2130 3248
rect -1968 3244 -1902 3260
rect -1548 3294 -1482 3310
rect -1548 3260 -1532 3294
rect -1498 3260 -1482 3294
rect -1950 3222 -1920 3244
rect -1740 3222 -1710 3248
rect -1548 3244 -1482 3260
rect -1128 3294 -1062 3310
rect -1128 3260 -1112 3294
rect -1078 3260 -1062 3294
rect -1530 3222 -1500 3244
rect -1320 3222 -1290 3248
rect -1128 3244 -1062 3260
rect -708 3294 -642 3310
rect -708 3260 -692 3294
rect -658 3260 -642 3294
rect -1110 3222 -1080 3244
rect -900 3222 -870 3248
rect -708 3244 -642 3260
rect -288 3294 -222 3310
rect -288 3260 -272 3294
rect -238 3260 -222 3294
rect -690 3222 -660 3244
rect -480 3222 -450 3248
rect -288 3244 -222 3260
rect 132 3294 198 3310
rect 132 3260 148 3294
rect 182 3260 198 3294
rect -270 3222 -240 3244
rect -60 3222 -30 3248
rect 132 3244 198 3260
rect 552 3294 618 3310
rect 552 3260 568 3294
rect 602 3260 618 3294
rect 150 3222 180 3244
rect 360 3222 390 3248
rect 552 3244 618 3260
rect 972 3294 1038 3310
rect 972 3260 988 3294
rect 1022 3260 1038 3294
rect 570 3222 600 3244
rect 780 3222 810 3248
rect 972 3244 1038 3260
rect 1392 3294 1458 3310
rect 1392 3260 1408 3294
rect 1442 3260 1458 3294
rect 990 3222 1020 3244
rect 1200 3222 1230 3248
rect 1392 3244 1458 3260
rect 1812 3294 1878 3310
rect 1812 3260 1828 3294
rect 1862 3260 1878 3294
rect 1410 3222 1440 3244
rect 1620 3222 1650 3248
rect 1812 3244 1878 3260
rect 2232 3294 2298 3310
rect 2232 3260 2248 3294
rect 2282 3260 2298 3294
rect 1830 3222 1860 3244
rect 2040 3222 2070 3248
rect 2232 3244 2298 3260
rect 2652 3294 2718 3310
rect 2652 3260 2668 3294
rect 2702 3260 2718 3294
rect 2250 3222 2280 3244
rect 2460 3222 2490 3248
rect 2652 3244 2718 3260
rect 3072 3294 3138 3310
rect 3072 3260 3088 3294
rect 3122 3260 3138 3294
rect 2670 3222 2700 3244
rect 2880 3222 2910 3248
rect 3072 3244 3138 3260
rect 3492 3294 3558 3310
rect 3492 3260 3508 3294
rect 3542 3260 3558 3294
rect 3090 3222 3120 3244
rect 3300 3222 3330 3248
rect 3492 3244 3558 3260
rect 3912 3294 3978 3310
rect 3912 3260 3928 3294
rect 3962 3260 3978 3294
rect 3510 3222 3540 3244
rect 3720 3222 3750 3248
rect 3912 3244 3978 3260
rect 4332 3294 4398 3310
rect 4332 3260 4348 3294
rect 4382 3260 4398 3294
rect 3930 3222 3960 3244
rect 4140 3222 4170 3248
rect 4332 3244 4398 3260
rect 4752 3294 4818 3310
rect 4752 3260 4768 3294
rect 4802 3260 4818 3294
rect 4350 3222 4380 3244
rect 4560 3222 4590 3248
rect 4752 3244 4818 3260
rect 5172 3294 5238 3310
rect 5172 3260 5188 3294
rect 5222 3260 5238 3294
rect 4770 3222 4800 3244
rect 4980 3222 5010 3248
rect 5172 3244 5238 3260
rect 5592 3294 5658 3310
rect 5592 3260 5608 3294
rect 5642 3260 5658 3294
rect 5190 3222 5220 3244
rect 5400 3222 5430 3248
rect 5592 3244 5658 3260
rect 6012 3294 6078 3310
rect 6012 3260 6028 3294
rect 6062 3260 6078 3294
rect 5610 3222 5640 3244
rect 5820 3222 5850 3248
rect 6012 3244 6078 3260
rect 6030 3222 6060 3244
rect -2580 3000 -2550 3022
rect -2598 2984 -2532 3000
rect -2370 2996 -2340 3022
rect -2160 3000 -2130 3022
rect -2598 2950 -2582 2984
rect -2548 2950 -2532 2984
rect -2598 2934 -2532 2950
rect -2178 2984 -2112 3000
rect -1950 2996 -1920 3022
rect -1740 3000 -1710 3022
rect -2178 2950 -2162 2984
rect -2128 2950 -2112 2984
rect -2178 2934 -2112 2950
rect -1758 2984 -1692 3000
rect -1530 2996 -1500 3022
rect -1320 3000 -1290 3022
rect -1758 2950 -1742 2984
rect -1708 2950 -1692 2984
rect -1758 2934 -1692 2950
rect -1338 2984 -1272 3000
rect -1110 2996 -1080 3022
rect -900 3000 -870 3022
rect -1338 2950 -1322 2984
rect -1288 2950 -1272 2984
rect -1338 2934 -1272 2950
rect -918 2984 -852 3000
rect -690 2996 -660 3022
rect -480 3000 -450 3022
rect -918 2950 -902 2984
rect -868 2950 -852 2984
rect -918 2934 -852 2950
rect -498 2984 -432 3000
rect -270 2996 -240 3022
rect -60 3000 -30 3022
rect -498 2950 -482 2984
rect -448 2950 -432 2984
rect -498 2934 -432 2950
rect -78 2984 -12 3000
rect 150 2996 180 3022
rect 360 3000 390 3022
rect -78 2950 -62 2984
rect -28 2950 -12 2984
rect -78 2934 -12 2950
rect 342 2984 408 3000
rect 570 2996 600 3022
rect 780 3000 810 3022
rect 342 2950 358 2984
rect 392 2950 408 2984
rect 342 2934 408 2950
rect 762 2984 828 3000
rect 990 2996 1020 3022
rect 1200 3000 1230 3022
rect 762 2950 778 2984
rect 812 2950 828 2984
rect 762 2934 828 2950
rect 1182 2984 1248 3000
rect 1410 2996 1440 3022
rect 1620 3000 1650 3022
rect 1182 2950 1198 2984
rect 1232 2950 1248 2984
rect 1182 2934 1248 2950
rect 1602 2984 1668 3000
rect 1830 2996 1860 3022
rect 2040 3000 2070 3022
rect 1602 2950 1618 2984
rect 1652 2950 1668 2984
rect 1602 2934 1668 2950
rect 2022 2984 2088 3000
rect 2250 2996 2280 3022
rect 2460 3000 2490 3022
rect 2022 2950 2038 2984
rect 2072 2950 2088 2984
rect 2022 2934 2088 2950
rect 2442 2984 2508 3000
rect 2670 2996 2700 3022
rect 2880 3000 2910 3022
rect 2442 2950 2458 2984
rect 2492 2950 2508 2984
rect 2442 2934 2508 2950
rect 2862 2984 2928 3000
rect 3090 2996 3120 3022
rect 3300 3000 3330 3022
rect 2862 2950 2878 2984
rect 2912 2950 2928 2984
rect 2862 2934 2928 2950
rect 3282 2984 3348 3000
rect 3510 2996 3540 3022
rect 3720 3000 3750 3022
rect 3282 2950 3298 2984
rect 3332 2950 3348 2984
rect 3282 2934 3348 2950
rect 3702 2984 3768 3000
rect 3930 2996 3960 3022
rect 4140 3000 4170 3022
rect 3702 2950 3718 2984
rect 3752 2950 3768 2984
rect 3702 2934 3768 2950
rect 4122 2984 4188 3000
rect 4350 2996 4380 3022
rect 4560 3000 4590 3022
rect 4122 2950 4138 2984
rect 4172 2950 4188 2984
rect 4122 2934 4188 2950
rect 4542 2984 4608 3000
rect 4770 2996 4800 3022
rect 4980 3000 5010 3022
rect 4542 2950 4558 2984
rect 4592 2950 4608 2984
rect 4542 2934 4608 2950
rect 4962 2984 5028 3000
rect 5190 2996 5220 3022
rect 5400 3000 5430 3022
rect 4962 2950 4978 2984
rect 5012 2950 5028 2984
rect 4962 2934 5028 2950
rect 5382 2984 5448 3000
rect 5610 2996 5640 3022
rect 5820 3000 5850 3022
rect 5382 2950 5398 2984
rect 5432 2950 5448 2984
rect 5382 2934 5448 2950
rect 5802 2984 5868 3000
rect 6030 2996 6060 3022
rect 5802 2950 5818 2984
rect 5852 2950 5868 2984
rect 5802 2934 5868 2950
rect -2388 2854 -2322 2870
rect -2388 2820 -2372 2854
rect -2338 2820 -2322 2854
rect -2580 2782 -2550 2808
rect -2388 2804 -2322 2820
rect -1968 2854 -1902 2870
rect -1968 2820 -1952 2854
rect -1918 2820 -1902 2854
rect -2370 2782 -2340 2804
rect -2160 2782 -2130 2808
rect -1968 2804 -1902 2820
rect -1548 2854 -1482 2870
rect -1548 2820 -1532 2854
rect -1498 2820 -1482 2854
rect -1950 2782 -1920 2804
rect -1740 2782 -1710 2808
rect -1548 2804 -1482 2820
rect -1128 2854 -1062 2870
rect -1128 2820 -1112 2854
rect -1078 2820 -1062 2854
rect -1530 2782 -1500 2804
rect -1320 2782 -1290 2808
rect -1128 2804 -1062 2820
rect -708 2854 -642 2870
rect -708 2820 -692 2854
rect -658 2820 -642 2854
rect -1110 2782 -1080 2804
rect -900 2782 -870 2808
rect -708 2804 -642 2820
rect -288 2854 -222 2870
rect -288 2820 -272 2854
rect -238 2820 -222 2854
rect -690 2782 -660 2804
rect -480 2782 -450 2808
rect -288 2804 -222 2820
rect 132 2854 198 2870
rect 132 2820 148 2854
rect 182 2820 198 2854
rect -270 2782 -240 2804
rect -60 2782 -30 2808
rect 132 2804 198 2820
rect 552 2854 618 2870
rect 552 2820 568 2854
rect 602 2820 618 2854
rect 150 2782 180 2804
rect 360 2782 390 2808
rect 552 2804 618 2820
rect 972 2854 1038 2870
rect 972 2820 988 2854
rect 1022 2820 1038 2854
rect 570 2782 600 2804
rect 780 2782 810 2808
rect 972 2804 1038 2820
rect 1392 2854 1458 2870
rect 1392 2820 1408 2854
rect 1442 2820 1458 2854
rect 990 2782 1020 2804
rect 1200 2782 1230 2808
rect 1392 2804 1458 2820
rect 1812 2854 1878 2870
rect 1812 2820 1828 2854
rect 1862 2820 1878 2854
rect 1410 2782 1440 2804
rect 1620 2782 1650 2808
rect 1812 2804 1878 2820
rect 2232 2854 2298 2870
rect 2232 2820 2248 2854
rect 2282 2820 2298 2854
rect 1830 2782 1860 2804
rect 2040 2782 2070 2808
rect 2232 2804 2298 2820
rect 2652 2854 2718 2870
rect 2652 2820 2668 2854
rect 2702 2820 2718 2854
rect 2250 2782 2280 2804
rect 2460 2782 2490 2808
rect 2652 2804 2718 2820
rect 3072 2854 3138 2870
rect 3072 2820 3088 2854
rect 3122 2820 3138 2854
rect 2670 2782 2700 2804
rect 2880 2782 2910 2808
rect 3072 2804 3138 2820
rect 3492 2854 3558 2870
rect 3492 2820 3508 2854
rect 3542 2820 3558 2854
rect 3090 2782 3120 2804
rect 3300 2782 3330 2808
rect 3492 2804 3558 2820
rect 3912 2854 3978 2870
rect 3912 2820 3928 2854
rect 3962 2820 3978 2854
rect 3510 2782 3540 2804
rect 3720 2782 3750 2808
rect 3912 2804 3978 2820
rect 4332 2854 4398 2870
rect 4332 2820 4348 2854
rect 4382 2820 4398 2854
rect 3930 2782 3960 2804
rect 4140 2782 4170 2808
rect 4332 2804 4398 2820
rect 4752 2854 4818 2870
rect 4752 2820 4768 2854
rect 4802 2820 4818 2854
rect 4350 2782 4380 2804
rect 4560 2782 4590 2808
rect 4752 2804 4818 2820
rect 5172 2854 5238 2870
rect 5172 2820 5188 2854
rect 5222 2820 5238 2854
rect 4770 2782 4800 2804
rect 4980 2782 5010 2808
rect 5172 2804 5238 2820
rect 5592 2854 5658 2870
rect 5592 2820 5608 2854
rect 5642 2820 5658 2854
rect 5190 2782 5220 2804
rect 5400 2782 5430 2808
rect 5592 2804 5658 2820
rect 6012 2854 6078 2870
rect 6012 2820 6028 2854
rect 6062 2820 6078 2854
rect 5610 2782 5640 2804
rect 5820 2782 5850 2808
rect 6012 2804 6078 2820
rect 6030 2782 6060 2804
rect -2580 2560 -2550 2582
rect -2598 2544 -2532 2560
rect -2370 2556 -2340 2582
rect -2160 2560 -2130 2582
rect -2598 2510 -2582 2544
rect -2548 2510 -2532 2544
rect -2598 2494 -2532 2510
rect -2178 2544 -2112 2560
rect -1950 2556 -1920 2582
rect -1740 2560 -1710 2582
rect -2178 2510 -2162 2544
rect -2128 2510 -2112 2544
rect -2178 2494 -2112 2510
rect -1758 2544 -1692 2560
rect -1530 2556 -1500 2582
rect -1320 2560 -1290 2582
rect -1758 2510 -1742 2544
rect -1708 2510 -1692 2544
rect -1758 2494 -1692 2510
rect -1338 2544 -1272 2560
rect -1110 2556 -1080 2582
rect -900 2560 -870 2582
rect -1338 2510 -1322 2544
rect -1288 2510 -1272 2544
rect -1338 2494 -1272 2510
rect -918 2544 -852 2560
rect -690 2556 -660 2582
rect -480 2560 -450 2582
rect -918 2510 -902 2544
rect -868 2510 -852 2544
rect -918 2494 -852 2510
rect -498 2544 -432 2560
rect -270 2556 -240 2582
rect -60 2560 -30 2582
rect -498 2510 -482 2544
rect -448 2510 -432 2544
rect -498 2494 -432 2510
rect -78 2544 -12 2560
rect 150 2556 180 2582
rect 360 2560 390 2582
rect -78 2510 -62 2544
rect -28 2510 -12 2544
rect -78 2494 -12 2510
rect 342 2544 408 2560
rect 570 2556 600 2582
rect 780 2560 810 2582
rect 342 2510 358 2544
rect 392 2510 408 2544
rect 342 2494 408 2510
rect 762 2544 828 2560
rect 990 2556 1020 2582
rect 1200 2560 1230 2582
rect 762 2510 778 2544
rect 812 2510 828 2544
rect 762 2494 828 2510
rect 1182 2544 1248 2560
rect 1410 2556 1440 2582
rect 1620 2560 1650 2582
rect 1182 2510 1198 2544
rect 1232 2510 1248 2544
rect 1182 2494 1248 2510
rect 1602 2544 1668 2560
rect 1830 2556 1860 2582
rect 2040 2560 2070 2582
rect 1602 2510 1618 2544
rect 1652 2510 1668 2544
rect 1602 2494 1668 2510
rect 2022 2544 2088 2560
rect 2250 2556 2280 2582
rect 2460 2560 2490 2582
rect 2022 2510 2038 2544
rect 2072 2510 2088 2544
rect 2022 2494 2088 2510
rect 2442 2544 2508 2560
rect 2670 2556 2700 2582
rect 2880 2560 2910 2582
rect 2442 2510 2458 2544
rect 2492 2510 2508 2544
rect 2442 2494 2508 2510
rect 2862 2544 2928 2560
rect 3090 2556 3120 2582
rect 3300 2560 3330 2582
rect 2862 2510 2878 2544
rect 2912 2510 2928 2544
rect 2862 2494 2928 2510
rect 3282 2544 3348 2560
rect 3510 2556 3540 2582
rect 3720 2560 3750 2582
rect 3282 2510 3298 2544
rect 3332 2510 3348 2544
rect 3282 2494 3348 2510
rect 3702 2544 3768 2560
rect 3930 2556 3960 2582
rect 4140 2560 4170 2582
rect 3702 2510 3718 2544
rect 3752 2510 3768 2544
rect 3702 2494 3768 2510
rect 4122 2544 4188 2560
rect 4350 2556 4380 2582
rect 4560 2560 4590 2582
rect 4122 2510 4138 2544
rect 4172 2510 4188 2544
rect 4122 2494 4188 2510
rect 4542 2544 4608 2560
rect 4770 2556 4800 2582
rect 4980 2560 5010 2582
rect 4542 2510 4558 2544
rect 4592 2510 4608 2544
rect 4542 2494 4608 2510
rect 4962 2544 5028 2560
rect 5190 2556 5220 2582
rect 5400 2560 5430 2582
rect 4962 2510 4978 2544
rect 5012 2510 5028 2544
rect 4962 2494 5028 2510
rect 5382 2544 5448 2560
rect 5610 2556 5640 2582
rect 5820 2560 5850 2582
rect 5382 2510 5398 2544
rect 5432 2510 5448 2544
rect 5382 2494 5448 2510
rect 5802 2544 5868 2560
rect 6030 2556 6060 2582
rect 5802 2510 5818 2544
rect 5852 2510 5868 2544
rect 5802 2494 5868 2510
rect -2388 2414 -2322 2430
rect -2388 2380 -2372 2414
rect -2338 2380 -2322 2414
rect -2580 2342 -2550 2368
rect -2388 2364 -2322 2380
rect -1968 2414 -1902 2430
rect -1968 2380 -1952 2414
rect -1918 2380 -1902 2414
rect -2370 2342 -2340 2364
rect -2160 2342 -2130 2368
rect -1968 2364 -1902 2380
rect -1548 2414 -1482 2430
rect -1548 2380 -1532 2414
rect -1498 2380 -1482 2414
rect -1950 2342 -1920 2364
rect -1740 2342 -1710 2368
rect -1548 2364 -1482 2380
rect -1128 2414 -1062 2430
rect -1128 2380 -1112 2414
rect -1078 2380 -1062 2414
rect -1530 2342 -1500 2364
rect -1320 2342 -1290 2368
rect -1128 2364 -1062 2380
rect -708 2414 -642 2430
rect -708 2380 -692 2414
rect -658 2380 -642 2414
rect -1110 2342 -1080 2364
rect -900 2342 -870 2368
rect -708 2364 -642 2380
rect -288 2414 -222 2430
rect -288 2380 -272 2414
rect -238 2380 -222 2414
rect -690 2342 -660 2364
rect -480 2342 -450 2368
rect -288 2364 -222 2380
rect 132 2414 198 2430
rect 132 2380 148 2414
rect 182 2380 198 2414
rect -270 2342 -240 2364
rect -60 2342 -30 2368
rect 132 2364 198 2380
rect 552 2414 618 2430
rect 552 2380 568 2414
rect 602 2380 618 2414
rect 150 2342 180 2364
rect 360 2342 390 2368
rect 552 2364 618 2380
rect 972 2414 1038 2430
rect 972 2380 988 2414
rect 1022 2380 1038 2414
rect 570 2342 600 2364
rect 780 2342 810 2368
rect 972 2364 1038 2380
rect 1392 2414 1458 2430
rect 1392 2380 1408 2414
rect 1442 2380 1458 2414
rect 990 2342 1020 2364
rect 1200 2342 1230 2368
rect 1392 2364 1458 2380
rect 1812 2414 1878 2430
rect 1812 2380 1828 2414
rect 1862 2380 1878 2414
rect 1410 2342 1440 2364
rect 1620 2342 1650 2368
rect 1812 2364 1878 2380
rect 2232 2414 2298 2430
rect 2232 2380 2248 2414
rect 2282 2380 2298 2414
rect 1830 2342 1860 2364
rect 2040 2342 2070 2368
rect 2232 2364 2298 2380
rect 2652 2414 2718 2430
rect 2652 2380 2668 2414
rect 2702 2380 2718 2414
rect 2250 2342 2280 2364
rect 2460 2342 2490 2368
rect 2652 2364 2718 2380
rect 3072 2414 3138 2430
rect 3072 2380 3088 2414
rect 3122 2380 3138 2414
rect 2670 2342 2700 2364
rect 2880 2342 2910 2368
rect 3072 2364 3138 2380
rect 3492 2414 3558 2430
rect 3492 2380 3508 2414
rect 3542 2380 3558 2414
rect 3090 2342 3120 2364
rect 3300 2342 3330 2368
rect 3492 2364 3558 2380
rect 3912 2414 3978 2430
rect 3912 2380 3928 2414
rect 3962 2380 3978 2414
rect 3510 2342 3540 2364
rect 3720 2342 3750 2368
rect 3912 2364 3978 2380
rect 4332 2414 4398 2430
rect 4332 2380 4348 2414
rect 4382 2380 4398 2414
rect 3930 2342 3960 2364
rect 4140 2342 4170 2368
rect 4332 2364 4398 2380
rect 4752 2414 4818 2430
rect 4752 2380 4768 2414
rect 4802 2380 4818 2414
rect 4350 2342 4380 2364
rect 4560 2342 4590 2368
rect 4752 2364 4818 2380
rect 5172 2414 5238 2430
rect 5172 2380 5188 2414
rect 5222 2380 5238 2414
rect 4770 2342 4800 2364
rect 4980 2342 5010 2368
rect 5172 2364 5238 2380
rect 5592 2414 5658 2430
rect 5592 2380 5608 2414
rect 5642 2380 5658 2414
rect 5190 2342 5220 2364
rect 5400 2342 5430 2368
rect 5592 2364 5658 2380
rect 6012 2414 6078 2430
rect 6012 2380 6028 2414
rect 6062 2380 6078 2414
rect 5610 2342 5640 2364
rect 5820 2342 5850 2368
rect 6012 2364 6078 2380
rect 6030 2342 6060 2364
rect -2580 2120 -2550 2142
rect -2598 2104 -2532 2120
rect -2370 2116 -2340 2142
rect -2160 2120 -2130 2142
rect -2598 2070 -2582 2104
rect -2548 2070 -2532 2104
rect -2598 2054 -2532 2070
rect -2178 2104 -2112 2120
rect -1950 2116 -1920 2142
rect -1740 2120 -1710 2142
rect -2178 2070 -2162 2104
rect -2128 2070 -2112 2104
rect -2178 2054 -2112 2070
rect -1758 2104 -1692 2120
rect -1530 2116 -1500 2142
rect -1320 2120 -1290 2142
rect -1758 2070 -1742 2104
rect -1708 2070 -1692 2104
rect -1758 2054 -1692 2070
rect -1338 2104 -1272 2120
rect -1110 2116 -1080 2142
rect -900 2120 -870 2142
rect -1338 2070 -1322 2104
rect -1288 2070 -1272 2104
rect -1338 2054 -1272 2070
rect -918 2104 -852 2120
rect -690 2116 -660 2142
rect -480 2120 -450 2142
rect -918 2070 -902 2104
rect -868 2070 -852 2104
rect -918 2054 -852 2070
rect -498 2104 -432 2120
rect -270 2116 -240 2142
rect -60 2120 -30 2142
rect -498 2070 -482 2104
rect -448 2070 -432 2104
rect -498 2054 -432 2070
rect -78 2104 -12 2120
rect 150 2116 180 2142
rect 360 2120 390 2142
rect -78 2070 -62 2104
rect -28 2070 -12 2104
rect -78 2054 -12 2070
rect 342 2104 408 2120
rect 570 2116 600 2142
rect 780 2120 810 2142
rect 342 2070 358 2104
rect 392 2070 408 2104
rect 342 2054 408 2070
rect 762 2104 828 2120
rect 990 2116 1020 2142
rect 1200 2120 1230 2142
rect 762 2070 778 2104
rect 812 2070 828 2104
rect 762 2054 828 2070
rect 1182 2104 1248 2120
rect 1410 2116 1440 2142
rect 1620 2120 1650 2142
rect 1182 2070 1198 2104
rect 1232 2070 1248 2104
rect 1182 2054 1248 2070
rect 1602 2104 1668 2120
rect 1830 2116 1860 2142
rect 2040 2120 2070 2142
rect 1602 2070 1618 2104
rect 1652 2070 1668 2104
rect 1602 2054 1668 2070
rect 2022 2104 2088 2120
rect 2250 2116 2280 2142
rect 2460 2120 2490 2142
rect 2022 2070 2038 2104
rect 2072 2070 2088 2104
rect 2022 2054 2088 2070
rect 2442 2104 2508 2120
rect 2670 2116 2700 2142
rect 2880 2120 2910 2142
rect 2442 2070 2458 2104
rect 2492 2070 2508 2104
rect 2442 2054 2508 2070
rect 2862 2104 2928 2120
rect 3090 2116 3120 2142
rect 3300 2120 3330 2142
rect 2862 2070 2878 2104
rect 2912 2070 2928 2104
rect 2862 2054 2928 2070
rect 3282 2104 3348 2120
rect 3510 2116 3540 2142
rect 3720 2120 3750 2142
rect 3282 2070 3298 2104
rect 3332 2070 3348 2104
rect 3282 2054 3348 2070
rect 3702 2104 3768 2120
rect 3930 2116 3960 2142
rect 4140 2120 4170 2142
rect 3702 2070 3718 2104
rect 3752 2070 3768 2104
rect 3702 2054 3768 2070
rect 4122 2104 4188 2120
rect 4350 2116 4380 2142
rect 4560 2120 4590 2142
rect 4122 2070 4138 2104
rect 4172 2070 4188 2104
rect 4122 2054 4188 2070
rect 4542 2104 4608 2120
rect 4770 2116 4800 2142
rect 4980 2120 5010 2142
rect 4542 2070 4558 2104
rect 4592 2070 4608 2104
rect 4542 2054 4608 2070
rect 4962 2104 5028 2120
rect 5190 2116 5220 2142
rect 5400 2120 5430 2142
rect 4962 2070 4978 2104
rect 5012 2070 5028 2104
rect 4962 2054 5028 2070
rect 5382 2104 5448 2120
rect 5610 2116 5640 2142
rect 5820 2120 5850 2142
rect 5382 2070 5398 2104
rect 5432 2070 5448 2104
rect 5382 2054 5448 2070
rect 5802 2104 5868 2120
rect 6030 2116 6060 2142
rect 5802 2070 5818 2104
rect 5852 2070 5868 2104
rect 5802 2054 5868 2070
rect -2388 1974 -2322 1990
rect -2388 1940 -2372 1974
rect -2338 1940 -2322 1974
rect -2580 1902 -2550 1928
rect -2388 1924 -2322 1940
rect -1968 1974 -1902 1990
rect -1968 1940 -1952 1974
rect -1918 1940 -1902 1974
rect -2370 1902 -2340 1924
rect -2160 1902 -2130 1928
rect -1968 1924 -1902 1940
rect -1548 1974 -1482 1990
rect -1548 1940 -1532 1974
rect -1498 1940 -1482 1974
rect -1950 1902 -1920 1924
rect -1740 1902 -1710 1928
rect -1548 1924 -1482 1940
rect -1128 1974 -1062 1990
rect -1128 1940 -1112 1974
rect -1078 1940 -1062 1974
rect -1530 1902 -1500 1924
rect -1320 1902 -1290 1928
rect -1128 1924 -1062 1940
rect -708 1974 -642 1990
rect -708 1940 -692 1974
rect -658 1940 -642 1974
rect -1110 1902 -1080 1924
rect -900 1902 -870 1928
rect -708 1924 -642 1940
rect -288 1974 -222 1990
rect -288 1940 -272 1974
rect -238 1940 -222 1974
rect -690 1902 -660 1924
rect -480 1902 -450 1928
rect -288 1924 -222 1940
rect 132 1974 198 1990
rect 132 1940 148 1974
rect 182 1940 198 1974
rect -270 1902 -240 1924
rect -60 1902 -30 1928
rect 132 1924 198 1940
rect 552 1974 618 1990
rect 552 1940 568 1974
rect 602 1940 618 1974
rect 150 1902 180 1924
rect 360 1902 390 1928
rect 552 1924 618 1940
rect 972 1974 1038 1990
rect 972 1940 988 1974
rect 1022 1940 1038 1974
rect 570 1902 600 1924
rect 780 1902 810 1928
rect 972 1924 1038 1940
rect 1392 1974 1458 1990
rect 1392 1940 1408 1974
rect 1442 1940 1458 1974
rect 990 1902 1020 1924
rect 1200 1902 1230 1928
rect 1392 1924 1458 1940
rect 1812 1974 1878 1990
rect 1812 1940 1828 1974
rect 1862 1940 1878 1974
rect 1410 1902 1440 1924
rect 1620 1902 1650 1928
rect 1812 1924 1878 1940
rect 2232 1974 2298 1990
rect 2232 1940 2248 1974
rect 2282 1940 2298 1974
rect 1830 1902 1860 1924
rect 2040 1902 2070 1928
rect 2232 1924 2298 1940
rect 2652 1974 2718 1990
rect 2652 1940 2668 1974
rect 2702 1940 2718 1974
rect 2250 1902 2280 1924
rect 2460 1902 2490 1928
rect 2652 1924 2718 1940
rect 3072 1974 3138 1990
rect 3072 1940 3088 1974
rect 3122 1940 3138 1974
rect 2670 1902 2700 1924
rect 2880 1902 2910 1928
rect 3072 1924 3138 1940
rect 3492 1974 3558 1990
rect 3492 1940 3508 1974
rect 3542 1940 3558 1974
rect 3090 1902 3120 1924
rect 3300 1902 3330 1928
rect 3492 1924 3558 1940
rect 3912 1974 3978 1990
rect 3912 1940 3928 1974
rect 3962 1940 3978 1974
rect 3510 1902 3540 1924
rect 3720 1902 3750 1928
rect 3912 1924 3978 1940
rect 4332 1974 4398 1990
rect 4332 1940 4348 1974
rect 4382 1940 4398 1974
rect 3930 1902 3960 1924
rect 4140 1902 4170 1928
rect 4332 1924 4398 1940
rect 4752 1974 4818 1990
rect 4752 1940 4768 1974
rect 4802 1940 4818 1974
rect 4350 1902 4380 1924
rect 4560 1902 4590 1928
rect 4752 1924 4818 1940
rect 5172 1974 5238 1990
rect 5172 1940 5188 1974
rect 5222 1940 5238 1974
rect 4770 1902 4800 1924
rect 4980 1902 5010 1928
rect 5172 1924 5238 1940
rect 5592 1974 5658 1990
rect 5592 1940 5608 1974
rect 5642 1940 5658 1974
rect 5190 1902 5220 1924
rect 5400 1902 5430 1928
rect 5592 1924 5658 1940
rect 6012 1974 6078 1990
rect 6012 1940 6028 1974
rect 6062 1940 6078 1974
rect 5610 1902 5640 1924
rect 5820 1902 5850 1928
rect 6012 1924 6078 1940
rect 6030 1902 6060 1924
rect -2580 1680 -2550 1702
rect -2598 1664 -2532 1680
rect -2370 1676 -2340 1702
rect -2160 1680 -2130 1702
rect -2598 1630 -2582 1664
rect -2548 1630 -2532 1664
rect -2598 1614 -2532 1630
rect -2178 1664 -2112 1680
rect -1950 1676 -1920 1702
rect -1740 1680 -1710 1702
rect -2178 1630 -2162 1664
rect -2128 1630 -2112 1664
rect -2178 1614 -2112 1630
rect -1758 1664 -1692 1680
rect -1530 1676 -1500 1702
rect -1320 1680 -1290 1702
rect -1758 1630 -1742 1664
rect -1708 1630 -1692 1664
rect -1758 1614 -1692 1630
rect -1338 1664 -1272 1680
rect -1110 1676 -1080 1702
rect -900 1680 -870 1702
rect -1338 1630 -1322 1664
rect -1288 1630 -1272 1664
rect -1338 1614 -1272 1630
rect -918 1664 -852 1680
rect -690 1676 -660 1702
rect -480 1680 -450 1702
rect -918 1630 -902 1664
rect -868 1630 -852 1664
rect -918 1614 -852 1630
rect -498 1664 -432 1680
rect -270 1676 -240 1702
rect -60 1680 -30 1702
rect -498 1630 -482 1664
rect -448 1630 -432 1664
rect -498 1614 -432 1630
rect -78 1664 -12 1680
rect 150 1676 180 1702
rect 360 1680 390 1702
rect -78 1630 -62 1664
rect -28 1630 -12 1664
rect -78 1614 -12 1630
rect 342 1664 408 1680
rect 570 1676 600 1702
rect 780 1680 810 1702
rect 342 1630 358 1664
rect 392 1630 408 1664
rect 342 1614 408 1630
rect 762 1664 828 1680
rect 990 1676 1020 1702
rect 1200 1680 1230 1702
rect 762 1630 778 1664
rect 812 1630 828 1664
rect 762 1614 828 1630
rect 1182 1664 1248 1680
rect 1410 1676 1440 1702
rect 1620 1680 1650 1702
rect 1182 1630 1198 1664
rect 1232 1630 1248 1664
rect 1182 1614 1248 1630
rect 1602 1664 1668 1680
rect 1830 1676 1860 1702
rect 2040 1680 2070 1702
rect 1602 1630 1618 1664
rect 1652 1630 1668 1664
rect 1602 1614 1668 1630
rect 2022 1664 2088 1680
rect 2250 1676 2280 1702
rect 2460 1680 2490 1702
rect 2022 1630 2038 1664
rect 2072 1630 2088 1664
rect 2022 1614 2088 1630
rect 2442 1664 2508 1680
rect 2670 1676 2700 1702
rect 2880 1680 2910 1702
rect 2442 1630 2458 1664
rect 2492 1630 2508 1664
rect 2442 1614 2508 1630
rect 2862 1664 2928 1680
rect 3090 1676 3120 1702
rect 3300 1680 3330 1702
rect 2862 1630 2878 1664
rect 2912 1630 2928 1664
rect 2862 1614 2928 1630
rect 3282 1664 3348 1680
rect 3510 1676 3540 1702
rect 3720 1680 3750 1702
rect 3282 1630 3298 1664
rect 3332 1630 3348 1664
rect 3282 1614 3348 1630
rect 3702 1664 3768 1680
rect 3930 1676 3960 1702
rect 4140 1680 4170 1702
rect 3702 1630 3718 1664
rect 3752 1630 3768 1664
rect 3702 1614 3768 1630
rect 4122 1664 4188 1680
rect 4350 1676 4380 1702
rect 4560 1680 4590 1702
rect 4122 1630 4138 1664
rect 4172 1630 4188 1664
rect 4122 1614 4188 1630
rect 4542 1664 4608 1680
rect 4770 1676 4800 1702
rect 4980 1680 5010 1702
rect 4542 1630 4558 1664
rect 4592 1630 4608 1664
rect 4542 1614 4608 1630
rect 4962 1664 5028 1680
rect 5190 1676 5220 1702
rect 5400 1680 5430 1702
rect 4962 1630 4978 1664
rect 5012 1630 5028 1664
rect 4962 1614 5028 1630
rect 5382 1664 5448 1680
rect 5610 1676 5640 1702
rect 5820 1680 5850 1702
rect 5382 1630 5398 1664
rect 5432 1630 5448 1664
rect 5382 1614 5448 1630
rect 5802 1664 5868 1680
rect 6030 1676 6060 1702
rect 5802 1630 5818 1664
rect 5852 1630 5868 1664
rect 5802 1614 5868 1630
rect -2388 1534 -2322 1550
rect -2388 1500 -2372 1534
rect -2338 1500 -2322 1534
rect -2580 1462 -2550 1488
rect -2388 1484 -2322 1500
rect -1968 1534 -1902 1550
rect -1968 1500 -1952 1534
rect -1918 1500 -1902 1534
rect -2370 1462 -2340 1484
rect -2160 1462 -2130 1488
rect -1968 1484 -1902 1500
rect -1548 1534 -1482 1550
rect -1548 1500 -1532 1534
rect -1498 1500 -1482 1534
rect -1950 1462 -1920 1484
rect -1740 1462 -1710 1488
rect -1548 1484 -1482 1500
rect -1128 1534 -1062 1550
rect -1128 1500 -1112 1534
rect -1078 1500 -1062 1534
rect -1530 1462 -1500 1484
rect -1320 1462 -1290 1488
rect -1128 1484 -1062 1500
rect -708 1534 -642 1550
rect -708 1500 -692 1534
rect -658 1500 -642 1534
rect -1110 1462 -1080 1484
rect -900 1462 -870 1488
rect -708 1484 -642 1500
rect -288 1534 -222 1550
rect -288 1500 -272 1534
rect -238 1500 -222 1534
rect -690 1462 -660 1484
rect -480 1462 -450 1488
rect -288 1484 -222 1500
rect 132 1534 198 1550
rect 132 1500 148 1534
rect 182 1500 198 1534
rect -270 1462 -240 1484
rect -60 1462 -30 1488
rect 132 1484 198 1500
rect 552 1534 618 1550
rect 552 1500 568 1534
rect 602 1500 618 1534
rect 150 1462 180 1484
rect 360 1462 390 1488
rect 552 1484 618 1500
rect 972 1534 1038 1550
rect 972 1500 988 1534
rect 1022 1500 1038 1534
rect 570 1462 600 1484
rect 780 1462 810 1488
rect 972 1484 1038 1500
rect 1392 1534 1458 1550
rect 1392 1500 1408 1534
rect 1442 1500 1458 1534
rect 990 1462 1020 1484
rect 1200 1462 1230 1488
rect 1392 1484 1458 1500
rect 1812 1534 1878 1550
rect 1812 1500 1828 1534
rect 1862 1500 1878 1534
rect 1410 1462 1440 1484
rect 1620 1462 1650 1488
rect 1812 1484 1878 1500
rect 2232 1534 2298 1550
rect 2232 1500 2248 1534
rect 2282 1500 2298 1534
rect 1830 1462 1860 1484
rect 2040 1462 2070 1488
rect 2232 1484 2298 1500
rect 2652 1534 2718 1550
rect 2652 1500 2668 1534
rect 2702 1500 2718 1534
rect 2250 1462 2280 1484
rect 2460 1462 2490 1488
rect 2652 1484 2718 1500
rect 3072 1534 3138 1550
rect 3072 1500 3088 1534
rect 3122 1500 3138 1534
rect 2670 1462 2700 1484
rect 2880 1462 2910 1488
rect 3072 1484 3138 1500
rect 3492 1534 3558 1550
rect 3492 1500 3508 1534
rect 3542 1500 3558 1534
rect 3090 1462 3120 1484
rect 3300 1462 3330 1488
rect 3492 1484 3558 1500
rect 3912 1534 3978 1550
rect 3912 1500 3928 1534
rect 3962 1500 3978 1534
rect 3510 1462 3540 1484
rect 3720 1462 3750 1488
rect 3912 1484 3978 1500
rect 4332 1534 4398 1550
rect 4332 1500 4348 1534
rect 4382 1500 4398 1534
rect 3930 1462 3960 1484
rect 4140 1462 4170 1488
rect 4332 1484 4398 1500
rect 4752 1534 4818 1550
rect 4752 1500 4768 1534
rect 4802 1500 4818 1534
rect 4350 1462 4380 1484
rect 4560 1462 4590 1488
rect 4752 1484 4818 1500
rect 5172 1534 5238 1550
rect 5172 1500 5188 1534
rect 5222 1500 5238 1534
rect 4770 1462 4800 1484
rect 4980 1462 5010 1488
rect 5172 1484 5238 1500
rect 5592 1534 5658 1550
rect 5592 1500 5608 1534
rect 5642 1500 5658 1534
rect 5190 1462 5220 1484
rect 5400 1462 5430 1488
rect 5592 1484 5658 1500
rect 6012 1534 6078 1550
rect 6012 1500 6028 1534
rect 6062 1500 6078 1534
rect 5610 1462 5640 1484
rect 5820 1462 5850 1488
rect 6012 1484 6078 1500
rect 6030 1462 6060 1484
rect -2580 1240 -2550 1262
rect -2598 1224 -2532 1240
rect -2370 1236 -2340 1262
rect -2160 1240 -2130 1262
rect -2598 1190 -2582 1224
rect -2548 1190 -2532 1224
rect -2598 1174 -2532 1190
rect -2178 1224 -2112 1240
rect -1950 1236 -1920 1262
rect -1740 1240 -1710 1262
rect -2178 1190 -2162 1224
rect -2128 1190 -2112 1224
rect -2178 1174 -2112 1190
rect -1758 1224 -1692 1240
rect -1530 1236 -1500 1262
rect -1320 1240 -1290 1262
rect -1758 1190 -1742 1224
rect -1708 1190 -1692 1224
rect -1758 1174 -1692 1190
rect -1338 1224 -1272 1240
rect -1110 1236 -1080 1262
rect -900 1240 -870 1262
rect -1338 1190 -1322 1224
rect -1288 1190 -1272 1224
rect -1338 1174 -1272 1190
rect -918 1224 -852 1240
rect -690 1236 -660 1262
rect -480 1240 -450 1262
rect -918 1190 -902 1224
rect -868 1190 -852 1224
rect -918 1174 -852 1190
rect -498 1224 -432 1240
rect -270 1236 -240 1262
rect -60 1240 -30 1262
rect -498 1190 -482 1224
rect -448 1190 -432 1224
rect -498 1174 -432 1190
rect -78 1224 -12 1240
rect 150 1236 180 1262
rect 360 1240 390 1262
rect -78 1190 -62 1224
rect -28 1190 -12 1224
rect -78 1174 -12 1190
rect 342 1224 408 1240
rect 570 1236 600 1262
rect 780 1240 810 1262
rect 342 1190 358 1224
rect 392 1190 408 1224
rect 342 1174 408 1190
rect 762 1224 828 1240
rect 990 1236 1020 1262
rect 1200 1240 1230 1262
rect 762 1190 778 1224
rect 812 1190 828 1224
rect 762 1174 828 1190
rect 1182 1224 1248 1240
rect 1410 1236 1440 1262
rect 1620 1240 1650 1262
rect 1182 1190 1198 1224
rect 1232 1190 1248 1224
rect 1182 1174 1248 1190
rect 1602 1224 1668 1240
rect 1830 1236 1860 1262
rect 2040 1240 2070 1262
rect 1602 1190 1618 1224
rect 1652 1190 1668 1224
rect 1602 1174 1668 1190
rect 2022 1224 2088 1240
rect 2250 1236 2280 1262
rect 2460 1240 2490 1262
rect 2022 1190 2038 1224
rect 2072 1190 2088 1224
rect 2022 1174 2088 1190
rect 2442 1224 2508 1240
rect 2670 1236 2700 1262
rect 2880 1240 2910 1262
rect 2442 1190 2458 1224
rect 2492 1190 2508 1224
rect 2442 1174 2508 1190
rect 2862 1224 2928 1240
rect 3090 1236 3120 1262
rect 3300 1240 3330 1262
rect 2862 1190 2878 1224
rect 2912 1190 2928 1224
rect 2862 1174 2928 1190
rect 3282 1224 3348 1240
rect 3510 1236 3540 1262
rect 3720 1240 3750 1262
rect 3282 1190 3298 1224
rect 3332 1190 3348 1224
rect 3282 1174 3348 1190
rect 3702 1224 3768 1240
rect 3930 1236 3960 1262
rect 4140 1240 4170 1262
rect 3702 1190 3718 1224
rect 3752 1190 3768 1224
rect 3702 1174 3768 1190
rect 4122 1224 4188 1240
rect 4350 1236 4380 1262
rect 4560 1240 4590 1262
rect 4122 1190 4138 1224
rect 4172 1190 4188 1224
rect 4122 1174 4188 1190
rect 4542 1224 4608 1240
rect 4770 1236 4800 1262
rect 4980 1240 5010 1262
rect 4542 1190 4558 1224
rect 4592 1190 4608 1224
rect 4542 1174 4608 1190
rect 4962 1224 5028 1240
rect 5190 1236 5220 1262
rect 5400 1240 5430 1262
rect 4962 1190 4978 1224
rect 5012 1190 5028 1224
rect 4962 1174 5028 1190
rect 5382 1224 5448 1240
rect 5610 1236 5640 1262
rect 5820 1240 5850 1262
rect 5382 1190 5398 1224
rect 5432 1190 5448 1224
rect 5382 1174 5448 1190
rect 5802 1224 5868 1240
rect 6030 1236 6060 1262
rect 5802 1190 5818 1224
rect 5852 1190 5868 1224
rect 5802 1174 5868 1190
rect -2388 1094 -2322 1110
rect -2388 1060 -2372 1094
rect -2338 1060 -2322 1094
rect -2580 1022 -2550 1048
rect -2388 1044 -2322 1060
rect -1968 1094 -1902 1110
rect -1968 1060 -1952 1094
rect -1918 1060 -1902 1094
rect -2370 1022 -2340 1044
rect -2160 1022 -2130 1048
rect -1968 1044 -1902 1060
rect -1548 1094 -1482 1110
rect -1548 1060 -1532 1094
rect -1498 1060 -1482 1094
rect -1950 1022 -1920 1044
rect -1740 1022 -1710 1048
rect -1548 1044 -1482 1060
rect -1128 1094 -1062 1110
rect -1128 1060 -1112 1094
rect -1078 1060 -1062 1094
rect -1530 1022 -1500 1044
rect -1320 1022 -1290 1048
rect -1128 1044 -1062 1060
rect -708 1094 -642 1110
rect -708 1060 -692 1094
rect -658 1060 -642 1094
rect -1110 1022 -1080 1044
rect -900 1022 -870 1048
rect -708 1044 -642 1060
rect -288 1094 -222 1110
rect -288 1060 -272 1094
rect -238 1060 -222 1094
rect -690 1022 -660 1044
rect -480 1022 -450 1048
rect -288 1044 -222 1060
rect 132 1094 198 1110
rect 132 1060 148 1094
rect 182 1060 198 1094
rect -270 1022 -240 1044
rect -60 1022 -30 1048
rect 132 1044 198 1060
rect 552 1094 618 1110
rect 552 1060 568 1094
rect 602 1060 618 1094
rect 150 1022 180 1044
rect 360 1022 390 1048
rect 552 1044 618 1060
rect 972 1094 1038 1110
rect 972 1060 988 1094
rect 1022 1060 1038 1094
rect 570 1022 600 1044
rect 780 1022 810 1048
rect 972 1044 1038 1060
rect 1392 1094 1458 1110
rect 1392 1060 1408 1094
rect 1442 1060 1458 1094
rect 990 1022 1020 1044
rect 1200 1022 1230 1048
rect 1392 1044 1458 1060
rect 1812 1094 1878 1110
rect 1812 1060 1828 1094
rect 1862 1060 1878 1094
rect 1410 1022 1440 1044
rect 1620 1022 1650 1048
rect 1812 1044 1878 1060
rect 2232 1094 2298 1110
rect 2232 1060 2248 1094
rect 2282 1060 2298 1094
rect 1830 1022 1860 1044
rect 2040 1022 2070 1048
rect 2232 1044 2298 1060
rect 2652 1094 2718 1110
rect 2652 1060 2668 1094
rect 2702 1060 2718 1094
rect 2250 1022 2280 1044
rect 2460 1022 2490 1048
rect 2652 1044 2718 1060
rect 3072 1094 3138 1110
rect 3072 1060 3088 1094
rect 3122 1060 3138 1094
rect 2670 1022 2700 1044
rect 2880 1022 2910 1048
rect 3072 1044 3138 1060
rect 3492 1094 3558 1110
rect 3492 1060 3508 1094
rect 3542 1060 3558 1094
rect 3090 1022 3120 1044
rect 3300 1022 3330 1048
rect 3492 1044 3558 1060
rect 3912 1094 3978 1110
rect 3912 1060 3928 1094
rect 3962 1060 3978 1094
rect 3510 1022 3540 1044
rect 3720 1022 3750 1048
rect 3912 1044 3978 1060
rect 4332 1094 4398 1110
rect 4332 1060 4348 1094
rect 4382 1060 4398 1094
rect 3930 1022 3960 1044
rect 4140 1022 4170 1048
rect 4332 1044 4398 1060
rect 4752 1094 4818 1110
rect 4752 1060 4768 1094
rect 4802 1060 4818 1094
rect 4350 1022 4380 1044
rect 4560 1022 4590 1048
rect 4752 1044 4818 1060
rect 5172 1094 5238 1110
rect 5172 1060 5188 1094
rect 5222 1060 5238 1094
rect 4770 1022 4800 1044
rect 4980 1022 5010 1048
rect 5172 1044 5238 1060
rect 5592 1094 5658 1110
rect 5592 1060 5608 1094
rect 5642 1060 5658 1094
rect 5190 1022 5220 1044
rect 5400 1022 5430 1048
rect 5592 1044 5658 1060
rect 6012 1094 6078 1110
rect 6012 1060 6028 1094
rect 6062 1060 6078 1094
rect 5610 1022 5640 1044
rect 5820 1022 5850 1048
rect 6012 1044 6078 1060
rect 6030 1022 6060 1044
rect -2580 800 -2550 822
rect -2598 784 -2532 800
rect -2370 796 -2340 822
rect -2160 800 -2130 822
rect -2598 750 -2582 784
rect -2548 750 -2532 784
rect -2598 734 -2532 750
rect -2178 784 -2112 800
rect -1950 796 -1920 822
rect -1740 800 -1710 822
rect -2178 750 -2162 784
rect -2128 750 -2112 784
rect -2178 734 -2112 750
rect -1758 784 -1692 800
rect -1530 796 -1500 822
rect -1320 800 -1290 822
rect -1758 750 -1742 784
rect -1708 750 -1692 784
rect -1758 734 -1692 750
rect -1338 784 -1272 800
rect -1110 796 -1080 822
rect -900 800 -870 822
rect -1338 750 -1322 784
rect -1288 750 -1272 784
rect -1338 734 -1272 750
rect -918 784 -852 800
rect -690 796 -660 822
rect -480 800 -450 822
rect -918 750 -902 784
rect -868 750 -852 784
rect -918 734 -852 750
rect -498 784 -432 800
rect -270 796 -240 822
rect -60 800 -30 822
rect -498 750 -482 784
rect -448 750 -432 784
rect -498 734 -432 750
rect -78 784 -12 800
rect 150 796 180 822
rect 360 800 390 822
rect -78 750 -62 784
rect -28 750 -12 784
rect -78 734 -12 750
rect 342 784 408 800
rect 570 796 600 822
rect 780 800 810 822
rect 342 750 358 784
rect 392 750 408 784
rect 342 734 408 750
rect 762 784 828 800
rect 990 796 1020 822
rect 1200 800 1230 822
rect 762 750 778 784
rect 812 750 828 784
rect 762 734 828 750
rect 1182 784 1248 800
rect 1410 796 1440 822
rect 1620 800 1650 822
rect 1182 750 1198 784
rect 1232 750 1248 784
rect 1182 734 1248 750
rect 1602 784 1668 800
rect 1830 796 1860 822
rect 2040 800 2070 822
rect 1602 750 1618 784
rect 1652 750 1668 784
rect 1602 734 1668 750
rect 2022 784 2088 800
rect 2250 796 2280 822
rect 2460 800 2490 822
rect 2022 750 2038 784
rect 2072 750 2088 784
rect 2022 734 2088 750
rect 2442 784 2508 800
rect 2670 796 2700 822
rect 2880 800 2910 822
rect 2442 750 2458 784
rect 2492 750 2508 784
rect 2442 734 2508 750
rect 2862 784 2928 800
rect 3090 796 3120 822
rect 3300 800 3330 822
rect 2862 750 2878 784
rect 2912 750 2928 784
rect 2862 734 2928 750
rect 3282 784 3348 800
rect 3510 796 3540 822
rect 3720 800 3750 822
rect 3282 750 3298 784
rect 3332 750 3348 784
rect 3282 734 3348 750
rect 3702 784 3768 800
rect 3930 796 3960 822
rect 4140 800 4170 822
rect 3702 750 3718 784
rect 3752 750 3768 784
rect 3702 734 3768 750
rect 4122 784 4188 800
rect 4350 796 4380 822
rect 4560 800 4590 822
rect 4122 750 4138 784
rect 4172 750 4188 784
rect 4122 734 4188 750
rect 4542 784 4608 800
rect 4770 796 4800 822
rect 4980 800 5010 822
rect 4542 750 4558 784
rect 4592 750 4608 784
rect 4542 734 4608 750
rect 4962 784 5028 800
rect 5190 796 5220 822
rect 5400 800 5430 822
rect 4962 750 4978 784
rect 5012 750 5028 784
rect 4962 734 5028 750
rect 5382 784 5448 800
rect 5610 796 5640 822
rect 5820 800 5850 822
rect 5382 750 5398 784
rect 5432 750 5448 784
rect 5382 734 5448 750
rect 5802 784 5868 800
rect 6030 796 6060 822
rect 5802 750 5818 784
rect 5852 750 5868 784
rect 5802 734 5868 750
rect 7062 5452 7128 5468
rect 7062 5450 7078 5452
rect 6804 5420 6831 5450
rect 7031 5420 7078 5450
rect 6734 5356 6800 5372
rect 6734 5322 6750 5356
rect 6784 5354 6800 5356
rect 7062 5418 7078 5420
rect 7112 5418 7128 5452
rect 7062 5402 7128 5418
rect 6784 5324 6831 5354
rect 7031 5324 7058 5354
rect 6784 5322 6800 5324
rect 6734 5306 6800 5322
rect 7062 5260 7128 5276
rect 7062 5258 7078 5260
rect 6804 5228 6831 5258
rect 7031 5228 7078 5258
rect 6734 5164 6800 5180
rect 6734 5130 6750 5164
rect 6784 5162 6800 5164
rect 7062 5226 7078 5228
rect 7112 5226 7128 5260
rect 7062 5210 7128 5226
rect 6784 5132 6831 5162
rect 7031 5132 7058 5162
rect 6784 5130 6800 5132
rect 6734 5114 6800 5130
rect 7062 5068 7128 5084
rect 7062 5066 7078 5068
rect 6804 5036 6831 5066
rect 7031 5036 7078 5066
rect 6734 4972 6800 4988
rect 6734 4938 6750 4972
rect 6784 4970 6800 4972
rect 7062 5034 7078 5036
rect 7112 5034 7128 5068
rect 7062 5018 7128 5034
rect 6784 4940 6831 4970
rect 7031 4940 7058 4970
rect 6784 4938 6800 4940
rect 6734 4922 6800 4938
rect 7062 4876 7128 4892
rect 7062 4874 7078 4876
rect 6804 4844 6831 4874
rect 7031 4844 7078 4874
rect 6734 4780 6800 4796
rect 6734 4746 6750 4780
rect 6784 4778 6800 4780
rect 7062 4842 7078 4844
rect 7112 4842 7128 4876
rect 7062 4826 7128 4842
rect 6784 4748 6831 4778
rect 7031 4748 7058 4778
rect 6784 4746 6800 4748
rect 6734 4730 6800 4746
rect 7062 4684 7128 4700
rect 7062 4682 7078 4684
rect 6804 4652 6831 4682
rect 7031 4652 7078 4682
rect 6734 4588 6800 4604
rect 6734 4554 6750 4588
rect 6784 4586 6800 4588
rect 7062 4650 7078 4652
rect 7112 4650 7128 4684
rect 7062 4634 7128 4650
rect 6784 4556 6831 4586
rect 7031 4556 7058 4586
rect 6784 4554 6800 4556
rect 6734 4538 6800 4554
rect 7062 4492 7128 4508
rect 7062 4490 7078 4492
rect 6804 4460 6831 4490
rect 7031 4460 7078 4490
rect 6734 4396 6800 4412
rect 6734 4362 6750 4396
rect 6784 4394 6800 4396
rect 7062 4458 7078 4460
rect 7112 4458 7128 4492
rect 7062 4442 7128 4458
rect 6784 4364 6831 4394
rect 7031 4364 7058 4394
rect 6784 4362 6800 4364
rect 6734 4346 6800 4362
rect 7062 4300 7128 4316
rect 7062 4298 7078 4300
rect 6804 4268 6831 4298
rect 7031 4268 7078 4298
rect 6734 4204 6800 4220
rect 6734 4170 6750 4204
rect 6784 4202 6800 4204
rect 7062 4266 7078 4268
rect 7112 4266 7128 4300
rect 7062 4250 7128 4266
rect 6784 4172 6831 4202
rect 7031 4172 7058 4202
rect 6784 4170 6800 4172
rect 6734 4154 6800 4170
rect 7062 4108 7128 4124
rect 7062 4106 7078 4108
rect 6804 4076 6831 4106
rect 7031 4076 7078 4106
rect 6734 4012 6800 4028
rect 6734 3978 6750 4012
rect 6784 4010 6800 4012
rect 7062 4074 7078 4076
rect 7112 4074 7128 4108
rect 7062 4058 7128 4074
rect 6784 3980 6831 4010
rect 7031 3980 7058 4010
rect 6784 3978 6800 3980
rect 6734 3962 6800 3978
rect 7062 3916 7128 3932
rect 7062 3914 7078 3916
rect 6804 3884 6831 3914
rect 7031 3884 7078 3914
rect 6734 3820 6800 3836
rect 6734 3786 6750 3820
rect 6784 3818 6800 3820
rect 7062 3882 7078 3884
rect 7112 3882 7128 3916
rect 7062 3866 7128 3882
rect 6784 3788 6831 3818
rect 7031 3788 7058 3818
rect 6784 3786 6800 3788
rect 6734 3770 6800 3786
rect 218 290 3260 306
rect 218 256 282 290
rect 316 256 474 290
rect 508 256 666 290
rect 700 256 858 290
rect 892 256 1050 290
rect 1084 256 1242 290
rect 1276 256 1434 290
rect 1468 256 1626 290
rect 1660 256 1818 290
rect 1852 256 2010 290
rect 2044 256 2202 290
rect 2236 256 2394 290
rect 2428 256 2586 290
rect 2620 256 2778 290
rect 2812 256 2970 290
rect 3004 256 3162 290
rect 3196 256 3260 290
rect 140 218 170 244
rect 218 240 3260 256
rect 236 218 266 240
rect 332 218 362 240
rect 428 218 458 240
rect 524 218 554 240
rect 620 218 650 240
rect 716 218 746 240
rect 812 218 842 240
rect 908 218 938 240
rect 1004 218 1034 240
rect 1100 218 1130 240
rect 1196 218 1226 240
rect 1292 218 1322 240
rect 1388 218 1418 240
rect 1484 218 1514 240
rect 1580 218 1610 240
rect 1676 218 1706 240
rect 1772 218 1802 240
rect 1868 218 1898 240
rect 1964 218 1994 240
rect 2060 218 2090 240
rect 2156 218 2186 240
rect 2252 218 2282 240
rect 2348 218 2378 240
rect 2444 218 2474 240
rect 2540 218 2570 240
rect 2636 218 2666 240
rect 2732 218 2762 240
rect 2828 218 2858 240
rect 2924 218 2954 240
rect 3020 218 3050 240
rect 3116 218 3146 240
rect 3212 218 3242 240
rect 3308 218 3338 244
rect 140 -4 170 18
rect 122 -20 188 -4
rect 236 -8 266 18
rect 332 -8 362 18
rect 428 -8 458 18
rect 524 -8 554 18
rect 620 -8 650 18
rect 716 -8 746 18
rect 812 -8 842 18
rect 908 -8 938 18
rect 1004 -8 1034 18
rect 1100 -8 1130 18
rect 1196 -8 1226 18
rect 1292 -8 1322 18
rect 1388 -8 1418 18
rect 1484 -8 1514 18
rect 1580 -8 1610 18
rect 1676 -8 1706 18
rect 1772 -8 1802 18
rect 1868 -8 1898 18
rect 1964 -8 1994 18
rect 2060 -8 2090 18
rect 2156 -8 2186 18
rect 2252 -8 2282 18
rect 2348 -8 2378 18
rect 2444 -8 2474 18
rect 2540 -8 2570 18
rect 2636 -8 2666 18
rect 2732 -8 2762 18
rect 2828 -8 2858 18
rect 2924 -8 2954 18
rect 3020 -8 3050 18
rect 3116 -8 3146 18
rect 3212 -8 3242 18
rect 3308 -8 3338 18
rect 122 -54 138 -20
rect 172 -54 188 -20
rect 122 -70 188 -54
rect 3290 -24 3356 -8
rect 3290 -58 3306 -24
rect 3340 -58 3356 -24
rect 3290 -74 3356 -58
<< polycont >>
rect 1423 10504 1457 10538
rect 1423 10376 1457 10410
rect 1423 10248 1457 10282
rect 1423 10120 1457 10154
rect 1387 10012 1421 10046
rect 1387 9884 1421 9918
rect 1387 9756 1421 9790
rect 1387 9628 1421 9662
rect 2031 10500 2065 10534
rect 2031 10372 2065 10406
rect 2031 10244 2065 10278
rect 2031 10116 2065 10150
rect 1995 10008 2029 10042
rect 1995 9880 2029 9914
rect 1995 9752 2029 9786
rect 1995 9624 2029 9658
rect 1397 9365 1431 9399
rect 2021 9365 2055 9399
rect 1397 9284 1431 9318
rect 2021 9284 2055 9318
rect 1397 9200 1431 9234
rect 2021 9200 2055 9234
rect 1397 9116 1431 9150
rect 2021 9116 2055 9150
rect 1397 8864 1431 8898
rect 2021 8864 2055 8898
rect 1397 8780 1431 8814
rect 2021 8780 2055 8814
rect 1397 8402 1431 8436
rect 2021 8402 2055 8436
rect 1397 8278 1431 8312
rect 2021 8278 2055 8312
rect -3650 7828 -3616 7862
rect -3650 7636 -3616 7670
rect -3322 7732 -3288 7766
rect -3650 7444 -3616 7478
rect -3322 7540 -3288 7574
rect -3650 7252 -3616 7286
rect -3322 7348 -3288 7382
rect -3650 7060 -3616 7094
rect -3322 7156 -3288 7190
rect -3650 6868 -3616 6902
rect -3322 6964 -3288 6998
rect -3650 6676 -3616 6710
rect -3322 6772 -3288 6806
rect -3650 6484 -3616 6518
rect -3322 6580 -3288 6614
rect -3650 6292 -3616 6326
rect -3322 6388 -3288 6422
rect -3322 6196 -3288 6230
rect -2386 7887 -2352 7921
rect -1966 7887 -1932 7921
rect -1546 7887 -1512 7921
rect -1126 7887 -1092 7921
rect -706 7887 -672 7921
rect -286 7887 -252 7921
rect 134 7887 168 7921
rect 554 7887 588 7921
rect 974 7887 1008 7921
rect 1394 7887 1428 7921
rect 1814 7887 1848 7921
rect 2234 7887 2268 7921
rect 2654 7887 2688 7921
rect 3074 7887 3108 7921
rect 3494 7887 3528 7921
rect 3914 7887 3948 7921
rect 4334 7887 4368 7921
rect 4754 7887 4788 7921
rect 5174 7887 5208 7921
rect 5594 7887 5628 7921
rect 6014 7887 6048 7921
rect -2596 7559 -2562 7593
rect -2176 7559 -2142 7593
rect -1756 7559 -1722 7593
rect -1336 7559 -1302 7593
rect -916 7559 -882 7593
rect -496 7559 -462 7593
rect -76 7559 -42 7593
rect 344 7559 378 7593
rect 764 7559 798 7593
rect 1184 7559 1218 7593
rect 1604 7559 1638 7593
rect 2024 7559 2058 7593
rect 2444 7559 2478 7593
rect 2864 7559 2898 7593
rect 3284 7559 3318 7593
rect 3704 7559 3738 7593
rect 4124 7559 4158 7593
rect 4544 7559 4578 7593
rect 4964 7559 4998 7593
rect 5384 7559 5418 7593
rect 5804 7559 5838 7593
rect -2384 7355 -2350 7389
rect -1964 7355 -1930 7389
rect -1544 7355 -1510 7389
rect -1124 7355 -1090 7389
rect -704 7355 -670 7389
rect -284 7355 -250 7389
rect 136 7355 170 7389
rect 556 7355 590 7389
rect 976 7355 1010 7389
rect 1396 7355 1430 7389
rect 1816 7355 1850 7389
rect 2236 7355 2270 7389
rect 2656 7355 2690 7389
rect 3076 7355 3110 7389
rect 3496 7355 3530 7389
rect 3916 7355 3950 7389
rect 4336 7355 4370 7389
rect 4756 7355 4790 7389
rect 5176 7355 5210 7389
rect 5596 7355 5630 7389
rect 6016 7355 6050 7389
rect -2594 7026 -2560 7060
rect -2174 7026 -2140 7060
rect -1754 7026 -1720 7060
rect -1334 7026 -1300 7060
rect -914 7026 -880 7060
rect -494 7026 -460 7060
rect -74 7026 -40 7060
rect 346 7026 380 7060
rect 766 7026 800 7060
rect 1186 7026 1220 7060
rect 1606 7026 1640 7060
rect 2026 7026 2060 7060
rect 2446 7026 2480 7060
rect 2866 7026 2900 7060
rect 3286 7026 3320 7060
rect 3706 7026 3740 7060
rect 4126 7026 4160 7060
rect 4546 7026 4580 7060
rect 4966 7026 5000 7060
rect 5386 7026 5420 7060
rect 5806 7026 5840 7060
rect -3648 5418 -3614 5452
rect -3648 5226 -3614 5260
rect -3320 5322 -3286 5356
rect -3648 5034 -3614 5068
rect -3320 5130 -3286 5164
rect -3648 4842 -3614 4876
rect -3320 4938 -3286 4972
rect -3648 4650 -3614 4684
rect -3320 4746 -3286 4780
rect -3648 4458 -3614 4492
rect -3320 4554 -3286 4588
rect -3648 4266 -3614 4300
rect -3320 4362 -3286 4396
rect -3648 4074 -3614 4108
rect -3320 4170 -3286 4204
rect -3648 3882 -3614 3916
rect -3320 3978 -3286 4012
rect -3320 3786 -3286 3820
rect -2372 6395 -2338 6429
rect -1952 6395 -1918 6429
rect -1532 6395 -1498 6429
rect -1112 6395 -1078 6429
rect -692 6395 -658 6429
rect -272 6395 -238 6429
rect 148 6395 182 6429
rect 568 6395 602 6429
rect 988 6395 1022 6429
rect 1408 6395 1442 6429
rect 1828 6395 1862 6429
rect 2248 6395 2282 6429
rect 2668 6395 2702 6429
rect 3088 6395 3122 6429
rect 3508 6395 3542 6429
rect 3928 6395 3962 6429
rect 4348 6395 4382 6429
rect 4768 6395 4802 6429
rect 5188 6395 5222 6429
rect 5608 6395 5642 6429
rect 6028 6395 6062 6429
rect -2582 6085 -2548 6119
rect -2162 6085 -2128 6119
rect -1742 6085 -1708 6119
rect -1322 6085 -1288 6119
rect -902 6085 -868 6119
rect -482 6085 -448 6119
rect -62 6085 -28 6119
rect 358 6085 392 6119
rect 778 6085 812 6119
rect 1198 6085 1232 6119
rect 1618 6085 1652 6119
rect 2038 6085 2072 6119
rect 2458 6085 2492 6119
rect 2878 6085 2912 6119
rect 3298 6085 3332 6119
rect 3718 6085 3752 6119
rect 4138 6085 4172 6119
rect 4558 6085 4592 6119
rect 4978 6085 5012 6119
rect 5398 6085 5432 6119
rect 5818 6085 5852 6119
rect -2372 5955 -2338 5989
rect -1952 5955 -1918 5989
rect -1532 5955 -1498 5989
rect -1112 5955 -1078 5989
rect -692 5955 -658 5989
rect -272 5955 -238 5989
rect 148 5955 182 5989
rect 568 5955 602 5989
rect 988 5955 1022 5989
rect 1408 5955 1442 5989
rect 1828 5955 1862 5989
rect 2248 5955 2282 5989
rect 2668 5955 2702 5989
rect 3088 5955 3122 5989
rect 3508 5955 3542 5989
rect 3928 5955 3962 5989
rect 4348 5955 4382 5989
rect 4768 5955 4802 5989
rect 5188 5955 5222 5989
rect 5608 5955 5642 5989
rect 6028 5955 6062 5989
rect -2582 5645 -2548 5679
rect -2162 5645 -2128 5679
rect -1742 5645 -1708 5679
rect -1322 5645 -1288 5679
rect -902 5645 -868 5679
rect -482 5645 -448 5679
rect -62 5645 -28 5679
rect 358 5645 392 5679
rect 778 5645 812 5679
rect 1198 5645 1232 5679
rect 1618 5645 1652 5679
rect 2038 5645 2072 5679
rect 2458 5645 2492 5679
rect 2878 5645 2912 5679
rect 3298 5645 3332 5679
rect 3718 5645 3752 5679
rect 4138 5645 4172 5679
rect 4558 5645 4592 5679
rect 4978 5645 5012 5679
rect 5398 5645 5432 5679
rect 5818 5645 5852 5679
rect -2372 5515 -2338 5549
rect -1952 5515 -1918 5549
rect -1532 5515 -1498 5549
rect -1112 5515 -1078 5549
rect -692 5515 -658 5549
rect -272 5515 -238 5549
rect 148 5515 182 5549
rect 568 5515 602 5549
rect 988 5515 1022 5549
rect 1408 5515 1442 5549
rect 1828 5515 1862 5549
rect 2248 5515 2282 5549
rect 2668 5515 2702 5549
rect 3088 5515 3122 5549
rect 3508 5515 3542 5549
rect 3928 5515 3962 5549
rect 4348 5515 4382 5549
rect 4768 5515 4802 5549
rect 5188 5515 5222 5549
rect 5608 5515 5642 5549
rect 6028 5515 6062 5549
rect -2582 5205 -2548 5239
rect -2162 5205 -2128 5239
rect -1742 5205 -1708 5239
rect -1322 5205 -1288 5239
rect -902 5205 -868 5239
rect -482 5205 -448 5239
rect -62 5205 -28 5239
rect 358 5205 392 5239
rect 778 5205 812 5239
rect 1198 5205 1232 5239
rect 1618 5205 1652 5239
rect 2038 5205 2072 5239
rect 2458 5205 2492 5239
rect 2878 5205 2912 5239
rect 3298 5205 3332 5239
rect 3718 5205 3752 5239
rect 4138 5205 4172 5239
rect 4558 5205 4592 5239
rect 4978 5205 5012 5239
rect 5398 5205 5432 5239
rect 5818 5205 5852 5239
rect -2372 5075 -2338 5109
rect -1952 5075 -1918 5109
rect -1532 5075 -1498 5109
rect -1112 5075 -1078 5109
rect -692 5075 -658 5109
rect -272 5075 -238 5109
rect 148 5075 182 5109
rect 568 5075 602 5109
rect 988 5075 1022 5109
rect 1408 5075 1442 5109
rect 1828 5075 1862 5109
rect 2248 5075 2282 5109
rect 2668 5075 2702 5109
rect 3088 5075 3122 5109
rect 3508 5075 3542 5109
rect 3928 5075 3962 5109
rect 4348 5075 4382 5109
rect 4768 5075 4802 5109
rect 5188 5075 5222 5109
rect 5608 5075 5642 5109
rect 6028 5075 6062 5109
rect -2582 4765 -2548 4799
rect -2162 4765 -2128 4799
rect -1742 4765 -1708 4799
rect -1322 4765 -1288 4799
rect -902 4765 -868 4799
rect -482 4765 -448 4799
rect -62 4765 -28 4799
rect 358 4765 392 4799
rect 778 4765 812 4799
rect 1198 4765 1232 4799
rect 1618 4765 1652 4799
rect 2038 4765 2072 4799
rect 2458 4765 2492 4799
rect 2878 4765 2912 4799
rect 3298 4765 3332 4799
rect 3718 4765 3752 4799
rect 4138 4765 4172 4799
rect 4558 4765 4592 4799
rect 4978 4765 5012 4799
rect 5398 4765 5432 4799
rect 5818 4765 5852 4799
rect 6750 7732 6784 7766
rect 7078 7828 7112 7862
rect 6750 7540 6784 7574
rect 7078 7636 7112 7670
rect 6750 7348 6784 7382
rect 7078 7444 7112 7478
rect 6750 7156 6784 7190
rect 7078 7252 7112 7286
rect 6750 6964 6784 6998
rect 7078 7060 7112 7094
rect 6750 6772 6784 6806
rect 7078 6868 7112 6902
rect 6750 6580 6784 6614
rect 7078 6676 7112 6710
rect 6750 6388 6784 6422
rect 7078 6484 7112 6518
rect 6750 6196 6784 6230
rect 7078 6292 7112 6326
rect -2372 4140 -2338 4174
rect -1952 4140 -1918 4174
rect -1532 4140 -1498 4174
rect -1112 4140 -1078 4174
rect -692 4140 -658 4174
rect -272 4140 -238 4174
rect 148 4140 182 4174
rect 568 4140 602 4174
rect 988 4140 1022 4174
rect 1408 4140 1442 4174
rect 1828 4140 1862 4174
rect 2248 4140 2282 4174
rect 2668 4140 2702 4174
rect 3088 4140 3122 4174
rect 3508 4140 3542 4174
rect 3928 4140 3962 4174
rect 4348 4140 4382 4174
rect 4768 4140 4802 4174
rect 5188 4140 5222 4174
rect 5608 4140 5642 4174
rect 6028 4140 6062 4174
rect -2582 3830 -2548 3864
rect -2162 3830 -2128 3864
rect -1742 3830 -1708 3864
rect -1322 3830 -1288 3864
rect -902 3830 -868 3864
rect -482 3830 -448 3864
rect -62 3830 -28 3864
rect 358 3830 392 3864
rect 778 3830 812 3864
rect 1198 3830 1232 3864
rect 1618 3830 1652 3864
rect 2038 3830 2072 3864
rect 2458 3830 2492 3864
rect 2878 3830 2912 3864
rect 3298 3830 3332 3864
rect 3718 3830 3752 3864
rect 4138 3830 4172 3864
rect 4558 3830 4592 3864
rect 4978 3830 5012 3864
rect 5398 3830 5432 3864
rect 5818 3830 5852 3864
rect -2372 3700 -2338 3734
rect -1952 3700 -1918 3734
rect -1532 3700 -1498 3734
rect -1112 3700 -1078 3734
rect -692 3700 -658 3734
rect -272 3700 -238 3734
rect 148 3700 182 3734
rect 568 3700 602 3734
rect 988 3700 1022 3734
rect 1408 3700 1442 3734
rect 1828 3700 1862 3734
rect 2248 3700 2282 3734
rect 2668 3700 2702 3734
rect 3088 3700 3122 3734
rect 3508 3700 3542 3734
rect 3928 3700 3962 3734
rect 4348 3700 4382 3734
rect 4768 3700 4802 3734
rect 5188 3700 5222 3734
rect 5608 3700 5642 3734
rect 6028 3700 6062 3734
rect -2582 3390 -2548 3424
rect -2162 3390 -2128 3424
rect -1742 3390 -1708 3424
rect -1322 3390 -1288 3424
rect -902 3390 -868 3424
rect -482 3390 -448 3424
rect -62 3390 -28 3424
rect 358 3390 392 3424
rect 778 3390 812 3424
rect 1198 3390 1232 3424
rect 1618 3390 1652 3424
rect 2038 3390 2072 3424
rect 2458 3390 2492 3424
rect 2878 3390 2912 3424
rect 3298 3390 3332 3424
rect 3718 3390 3752 3424
rect 4138 3390 4172 3424
rect 4558 3390 4592 3424
rect 4978 3390 5012 3424
rect 5398 3390 5432 3424
rect 5818 3390 5852 3424
rect -2372 3260 -2338 3294
rect -1952 3260 -1918 3294
rect -1532 3260 -1498 3294
rect -1112 3260 -1078 3294
rect -692 3260 -658 3294
rect -272 3260 -238 3294
rect 148 3260 182 3294
rect 568 3260 602 3294
rect 988 3260 1022 3294
rect 1408 3260 1442 3294
rect 1828 3260 1862 3294
rect 2248 3260 2282 3294
rect 2668 3260 2702 3294
rect 3088 3260 3122 3294
rect 3508 3260 3542 3294
rect 3928 3260 3962 3294
rect 4348 3260 4382 3294
rect 4768 3260 4802 3294
rect 5188 3260 5222 3294
rect 5608 3260 5642 3294
rect 6028 3260 6062 3294
rect -2582 2950 -2548 2984
rect -2162 2950 -2128 2984
rect -1742 2950 -1708 2984
rect -1322 2950 -1288 2984
rect -902 2950 -868 2984
rect -482 2950 -448 2984
rect -62 2950 -28 2984
rect 358 2950 392 2984
rect 778 2950 812 2984
rect 1198 2950 1232 2984
rect 1618 2950 1652 2984
rect 2038 2950 2072 2984
rect 2458 2950 2492 2984
rect 2878 2950 2912 2984
rect 3298 2950 3332 2984
rect 3718 2950 3752 2984
rect 4138 2950 4172 2984
rect 4558 2950 4592 2984
rect 4978 2950 5012 2984
rect 5398 2950 5432 2984
rect 5818 2950 5852 2984
rect -2372 2820 -2338 2854
rect -1952 2820 -1918 2854
rect -1532 2820 -1498 2854
rect -1112 2820 -1078 2854
rect -692 2820 -658 2854
rect -272 2820 -238 2854
rect 148 2820 182 2854
rect 568 2820 602 2854
rect 988 2820 1022 2854
rect 1408 2820 1442 2854
rect 1828 2820 1862 2854
rect 2248 2820 2282 2854
rect 2668 2820 2702 2854
rect 3088 2820 3122 2854
rect 3508 2820 3542 2854
rect 3928 2820 3962 2854
rect 4348 2820 4382 2854
rect 4768 2820 4802 2854
rect 5188 2820 5222 2854
rect 5608 2820 5642 2854
rect 6028 2820 6062 2854
rect -2582 2510 -2548 2544
rect -2162 2510 -2128 2544
rect -1742 2510 -1708 2544
rect -1322 2510 -1288 2544
rect -902 2510 -868 2544
rect -482 2510 -448 2544
rect -62 2510 -28 2544
rect 358 2510 392 2544
rect 778 2510 812 2544
rect 1198 2510 1232 2544
rect 1618 2510 1652 2544
rect 2038 2510 2072 2544
rect 2458 2510 2492 2544
rect 2878 2510 2912 2544
rect 3298 2510 3332 2544
rect 3718 2510 3752 2544
rect 4138 2510 4172 2544
rect 4558 2510 4592 2544
rect 4978 2510 5012 2544
rect 5398 2510 5432 2544
rect 5818 2510 5852 2544
rect -2372 2380 -2338 2414
rect -1952 2380 -1918 2414
rect -1532 2380 -1498 2414
rect -1112 2380 -1078 2414
rect -692 2380 -658 2414
rect -272 2380 -238 2414
rect 148 2380 182 2414
rect 568 2380 602 2414
rect 988 2380 1022 2414
rect 1408 2380 1442 2414
rect 1828 2380 1862 2414
rect 2248 2380 2282 2414
rect 2668 2380 2702 2414
rect 3088 2380 3122 2414
rect 3508 2380 3542 2414
rect 3928 2380 3962 2414
rect 4348 2380 4382 2414
rect 4768 2380 4802 2414
rect 5188 2380 5222 2414
rect 5608 2380 5642 2414
rect 6028 2380 6062 2414
rect -2582 2070 -2548 2104
rect -2162 2070 -2128 2104
rect -1742 2070 -1708 2104
rect -1322 2070 -1288 2104
rect -902 2070 -868 2104
rect -482 2070 -448 2104
rect -62 2070 -28 2104
rect 358 2070 392 2104
rect 778 2070 812 2104
rect 1198 2070 1232 2104
rect 1618 2070 1652 2104
rect 2038 2070 2072 2104
rect 2458 2070 2492 2104
rect 2878 2070 2912 2104
rect 3298 2070 3332 2104
rect 3718 2070 3752 2104
rect 4138 2070 4172 2104
rect 4558 2070 4592 2104
rect 4978 2070 5012 2104
rect 5398 2070 5432 2104
rect 5818 2070 5852 2104
rect -2372 1940 -2338 1974
rect -1952 1940 -1918 1974
rect -1532 1940 -1498 1974
rect -1112 1940 -1078 1974
rect -692 1940 -658 1974
rect -272 1940 -238 1974
rect 148 1940 182 1974
rect 568 1940 602 1974
rect 988 1940 1022 1974
rect 1408 1940 1442 1974
rect 1828 1940 1862 1974
rect 2248 1940 2282 1974
rect 2668 1940 2702 1974
rect 3088 1940 3122 1974
rect 3508 1940 3542 1974
rect 3928 1940 3962 1974
rect 4348 1940 4382 1974
rect 4768 1940 4802 1974
rect 5188 1940 5222 1974
rect 5608 1940 5642 1974
rect 6028 1940 6062 1974
rect -2582 1630 -2548 1664
rect -2162 1630 -2128 1664
rect -1742 1630 -1708 1664
rect -1322 1630 -1288 1664
rect -902 1630 -868 1664
rect -482 1630 -448 1664
rect -62 1630 -28 1664
rect 358 1630 392 1664
rect 778 1630 812 1664
rect 1198 1630 1232 1664
rect 1618 1630 1652 1664
rect 2038 1630 2072 1664
rect 2458 1630 2492 1664
rect 2878 1630 2912 1664
rect 3298 1630 3332 1664
rect 3718 1630 3752 1664
rect 4138 1630 4172 1664
rect 4558 1630 4592 1664
rect 4978 1630 5012 1664
rect 5398 1630 5432 1664
rect 5818 1630 5852 1664
rect -2372 1500 -2338 1534
rect -1952 1500 -1918 1534
rect -1532 1500 -1498 1534
rect -1112 1500 -1078 1534
rect -692 1500 -658 1534
rect -272 1500 -238 1534
rect 148 1500 182 1534
rect 568 1500 602 1534
rect 988 1500 1022 1534
rect 1408 1500 1442 1534
rect 1828 1500 1862 1534
rect 2248 1500 2282 1534
rect 2668 1500 2702 1534
rect 3088 1500 3122 1534
rect 3508 1500 3542 1534
rect 3928 1500 3962 1534
rect 4348 1500 4382 1534
rect 4768 1500 4802 1534
rect 5188 1500 5222 1534
rect 5608 1500 5642 1534
rect 6028 1500 6062 1534
rect -2582 1190 -2548 1224
rect -2162 1190 -2128 1224
rect -1742 1190 -1708 1224
rect -1322 1190 -1288 1224
rect -902 1190 -868 1224
rect -482 1190 -448 1224
rect -62 1190 -28 1224
rect 358 1190 392 1224
rect 778 1190 812 1224
rect 1198 1190 1232 1224
rect 1618 1190 1652 1224
rect 2038 1190 2072 1224
rect 2458 1190 2492 1224
rect 2878 1190 2912 1224
rect 3298 1190 3332 1224
rect 3718 1190 3752 1224
rect 4138 1190 4172 1224
rect 4558 1190 4592 1224
rect 4978 1190 5012 1224
rect 5398 1190 5432 1224
rect 5818 1190 5852 1224
rect -2372 1060 -2338 1094
rect -1952 1060 -1918 1094
rect -1532 1060 -1498 1094
rect -1112 1060 -1078 1094
rect -692 1060 -658 1094
rect -272 1060 -238 1094
rect 148 1060 182 1094
rect 568 1060 602 1094
rect 988 1060 1022 1094
rect 1408 1060 1442 1094
rect 1828 1060 1862 1094
rect 2248 1060 2282 1094
rect 2668 1060 2702 1094
rect 3088 1060 3122 1094
rect 3508 1060 3542 1094
rect 3928 1060 3962 1094
rect 4348 1060 4382 1094
rect 4768 1060 4802 1094
rect 5188 1060 5222 1094
rect 5608 1060 5642 1094
rect 6028 1060 6062 1094
rect -2582 750 -2548 784
rect -2162 750 -2128 784
rect -1742 750 -1708 784
rect -1322 750 -1288 784
rect -902 750 -868 784
rect -482 750 -448 784
rect -62 750 -28 784
rect 358 750 392 784
rect 778 750 812 784
rect 1198 750 1232 784
rect 1618 750 1652 784
rect 2038 750 2072 784
rect 2458 750 2492 784
rect 2878 750 2912 784
rect 3298 750 3332 784
rect 3718 750 3752 784
rect 4138 750 4172 784
rect 4558 750 4592 784
rect 4978 750 5012 784
rect 5398 750 5432 784
rect 5818 750 5852 784
rect 6750 5322 6784 5356
rect 7078 5418 7112 5452
rect 6750 5130 6784 5164
rect 7078 5226 7112 5260
rect 6750 4938 6784 4972
rect 7078 5034 7112 5068
rect 6750 4746 6784 4780
rect 7078 4842 7112 4876
rect 6750 4554 6784 4588
rect 7078 4650 7112 4684
rect 6750 4362 6784 4396
rect 7078 4458 7112 4492
rect 6750 4170 6784 4204
rect 7078 4266 7112 4300
rect 6750 3978 6784 4012
rect 7078 4074 7112 4108
rect 6750 3786 6784 3820
rect 7078 3882 7112 3916
rect 282 256 316 290
rect 474 256 508 290
rect 666 256 700 290
rect 858 256 892 290
rect 1050 256 1084 290
rect 1242 256 1276 290
rect 1434 256 1468 290
rect 1626 256 1660 290
rect 1818 256 1852 290
rect 2010 256 2044 290
rect 2202 256 2236 290
rect 2394 256 2428 290
rect 2586 256 2620 290
rect 2778 256 2812 290
rect 2970 256 3004 290
rect 3162 256 3196 290
rect 138 -54 172 -20
rect 3306 -58 3340 -24
<< locali >>
rect 1165 10616 1199 10633
rect 1709 10616 1743 10633
rect 1165 10604 1457 10616
rect 1199 10598 1457 10604
rect 1199 10570 1260 10598
rect 1165 10564 1260 10570
rect 1294 10564 1457 10598
rect 1165 10538 1457 10564
rect 1165 10512 1423 10538
rect 1199 10504 1423 10512
rect 1199 10478 1457 10504
rect 1165 10420 1457 10478
rect 1199 10410 1457 10420
rect 1199 10386 1423 10410
rect 1165 10376 1423 10386
rect 1165 10328 1457 10376
rect 1199 10294 1457 10328
rect 1165 10282 1457 10294
rect 1165 10248 1423 10282
rect 1165 10236 1457 10248
rect 1199 10202 1457 10236
rect 1165 10154 1457 10202
rect 1165 10144 1423 10154
rect 1199 10120 1423 10144
rect 1199 10110 1457 10120
rect 1165 10100 1457 10110
rect 1491 10615 1743 10616
rect 2253 10615 2287 10633
rect 1491 10604 2065 10615
rect 1491 10598 1709 10604
rect 1491 10564 1531 10598
rect 1565 10564 1633 10598
rect 1667 10570 1709 10598
rect 1743 10598 2065 10604
rect 1743 10570 1785 10598
rect 1667 10564 1785 10570
rect 1819 10564 1887 10598
rect 1921 10564 2065 10598
rect 1491 10534 2065 10564
rect 1491 10512 2031 10534
rect 1491 10478 1709 10512
rect 1743 10500 2031 10512
rect 1743 10478 2065 10500
rect 1491 10420 2065 10478
rect 1491 10386 1709 10420
rect 1743 10406 2065 10420
rect 1743 10386 2031 10406
rect 1491 10372 2031 10386
rect 1491 10328 2065 10372
rect 1491 10294 1709 10328
rect 1743 10294 2065 10328
rect 1491 10278 2065 10294
rect 1491 10244 2031 10278
rect 1491 10236 2065 10244
rect 1491 10202 1709 10236
rect 1743 10202 2065 10236
rect 1491 10150 2065 10202
rect 1491 10144 2031 10150
rect 1491 10110 1709 10144
rect 1743 10116 2031 10144
rect 1743 10110 2065 10116
rect 1165 10052 1353 10100
rect 1491 10096 2065 10110
rect 2099 10604 2287 10615
rect 2099 10598 2253 10604
rect 2099 10564 2158 10598
rect 2192 10570 2253 10598
rect 2192 10564 2287 10570
rect 2099 10512 2287 10564
rect 2099 10478 2253 10512
rect 2099 10420 2287 10478
rect 2099 10386 2253 10420
rect 2099 10328 2287 10386
rect 2099 10294 2253 10328
rect 2099 10236 2287 10294
rect 2099 10202 2253 10236
rect 2099 10144 2287 10202
rect 2099 10110 2253 10144
rect 1491 10066 1961 10096
rect 1199 10018 1353 10052
rect 1165 9960 1353 10018
rect 1199 9926 1353 9960
rect 1165 9868 1353 9926
rect 1199 9834 1353 9868
rect 1165 9776 1353 9834
rect 1199 9742 1353 9776
rect 1165 9684 1353 9742
rect 1199 9650 1353 9684
rect 1165 9598 1353 9650
rect 1165 9592 1260 9598
rect 1199 9564 1260 9592
rect 1294 9564 1353 9598
rect 1199 9558 1353 9564
rect 1165 9547 1353 9558
rect 1387 10052 1961 10066
rect 2099 10062 2287 10110
rect 1387 10046 1709 10052
rect 1421 10018 1709 10046
rect 1743 10018 1961 10052
rect 1421 10012 1961 10018
rect 1387 9960 1961 10012
rect 1387 9926 1709 9960
rect 1743 9926 1961 9960
rect 1387 9918 1961 9926
rect 1421 9884 1961 9918
rect 1387 9868 1961 9884
rect 1387 9834 1709 9868
rect 1743 9834 1961 9868
rect 1387 9790 1961 9834
rect 1421 9776 1961 9790
rect 1421 9756 1709 9776
rect 1387 9742 1709 9756
rect 1743 9742 1961 9776
rect 1387 9684 1961 9742
rect 1387 9662 1709 9684
rect 1421 9650 1709 9662
rect 1743 9650 1961 9684
rect 1421 9628 1961 9650
rect 1387 9598 1961 9628
rect 1387 9564 1531 9598
rect 1565 9564 1633 9598
rect 1667 9592 1785 9598
rect 1667 9564 1709 9592
rect 1387 9558 1709 9564
rect 1743 9564 1785 9592
rect 1819 9564 1887 9598
rect 1921 9564 1961 9598
rect 1743 9558 1961 9564
rect 1387 9547 1961 9558
rect 1165 9512 1199 9547
rect 1709 9546 1961 9547
rect 1995 10052 2287 10062
rect 1995 10042 2253 10052
rect 2029 10018 2253 10042
rect 2029 10008 2287 10018
rect 1995 9960 2287 10008
rect 1995 9926 2253 9960
rect 1995 9914 2287 9926
rect 2029 9880 2287 9914
rect 1995 9868 2287 9880
rect 1995 9834 2253 9868
rect 1995 9786 2287 9834
rect 2029 9776 2287 9786
rect 2029 9752 2253 9776
rect 1995 9742 2253 9752
rect 1995 9684 2287 9742
rect 1995 9658 2253 9684
rect 2029 9650 2253 9658
rect 2029 9624 2287 9650
rect 1995 9598 2287 9624
rect 1995 9564 2158 9598
rect 2192 9592 2287 9598
rect 2192 9564 2253 9592
rect 1995 9558 2253 9564
rect 1995 9546 2287 9558
rect 1709 9512 1743 9546
rect 2253 9512 2287 9546
rect 1165 9500 1344 9512
rect 1199 9466 1293 9500
rect 1327 9466 1344 9500
rect 1165 9454 1344 9466
rect 1476 9500 1976 9512
rect 1476 9466 1511 9500
rect 1545 9466 1604 9500
rect 1638 9466 1709 9500
rect 1743 9466 1814 9500
rect 1848 9466 1907 9500
rect 1941 9466 1976 9500
rect 1476 9454 1976 9466
rect 2108 9500 2287 9512
rect 2108 9466 2125 9500
rect 2159 9466 2253 9500
rect 2108 9454 2287 9466
rect 1165 9408 1199 9454
rect 1709 9419 1743 9454
rect 1165 9318 1199 9374
rect 1233 9402 1363 9419
rect 1233 9368 1241 9402
rect 1275 9368 1309 9402
rect 1343 9368 1363 9402
rect 1233 9352 1363 9368
rect 1165 9316 1241 9318
rect 1199 9284 1241 9316
rect 1275 9284 1291 9318
rect 1165 9224 1199 9282
rect 1325 9250 1363 9352
rect 1165 9150 1199 9190
rect 1233 9234 1363 9250
rect 1233 9200 1241 9234
rect 1275 9200 1309 9234
rect 1343 9200 1363 9234
rect 1233 9184 1363 9200
rect 1165 9132 1241 9150
rect 1199 9116 1241 9132
rect 1275 9116 1291 9150
rect 1165 9040 1199 9098
rect 1325 9082 1363 9184
rect 1397 9399 1447 9415
rect 1431 9365 1447 9399
rect 1481 9408 1971 9419
rect 1481 9402 1709 9408
rect 1481 9368 1497 9402
rect 1531 9368 1565 9402
rect 1599 9368 1633 9402
rect 1667 9374 1709 9402
rect 1743 9402 1971 9408
rect 1743 9374 1785 9402
rect 1667 9368 1785 9374
rect 1819 9368 1853 9402
rect 1887 9368 1921 9402
rect 1955 9368 1971 9402
rect 2005 9399 2055 9415
rect 1397 9356 1447 9365
rect 1397 9322 1404 9356
rect 1438 9322 1447 9356
rect 1397 9318 1447 9322
rect 1431 9284 1447 9318
rect 1397 9265 1447 9284
rect 1397 9234 1404 9265
rect 1438 9231 1447 9265
rect 1431 9200 1447 9231
rect 1397 9150 1447 9200
rect 1431 9116 1447 9150
rect 1397 9091 1447 9116
rect 1481 9318 1675 9334
rect 1481 9284 1497 9318
rect 1531 9284 1565 9318
rect 1599 9284 1633 9318
rect 1667 9284 1675 9318
rect 1481 9268 1675 9284
rect 1709 9316 1743 9368
rect 2005 9365 2021 9399
rect 2005 9364 2055 9365
rect 1481 9166 1515 9268
rect 1709 9234 1743 9282
rect 1777 9318 1971 9334
rect 1777 9284 1785 9318
rect 1819 9284 1853 9318
rect 1887 9284 1921 9318
rect 1955 9284 1971 9318
rect 1777 9268 1971 9284
rect 1549 9200 1565 9234
rect 1599 9200 1633 9234
rect 1667 9224 1785 9234
rect 1667 9200 1709 9224
rect 1743 9200 1785 9224
rect 1819 9200 1853 9234
rect 1887 9200 1903 9234
rect 1481 9150 1675 9166
rect 1481 9116 1497 9150
rect 1531 9116 1565 9150
rect 1599 9116 1633 9150
rect 1667 9116 1675 9150
rect 1481 9100 1675 9116
rect 1709 9132 1743 9190
rect 1937 9166 1971 9268
rect 1165 8948 1199 9006
rect 1165 8856 1199 8914
rect 1165 8764 1199 8822
rect 1165 8672 1199 8730
rect 1233 9066 1363 9082
rect 1233 9032 1241 9066
rect 1275 9032 1309 9066
rect 1343 9032 1363 9066
rect 1481 9055 1515 9100
rect 1777 9150 1971 9166
rect 1777 9116 1785 9150
rect 1819 9116 1853 9150
rect 1887 9116 1921 9150
rect 1955 9116 1971 9150
rect 1777 9100 1971 9116
rect 1709 9066 1743 9098
rect 1233 8898 1275 9032
rect 1397 8998 1515 9055
rect 1549 9032 1565 9066
rect 1599 9032 1633 9066
rect 1667 9040 1785 9066
rect 1667 9032 1709 9040
rect 1743 9032 1785 9040
rect 1819 9032 1853 9066
rect 1887 9032 1903 9066
rect 1937 9055 1971 9100
rect 2005 9330 2016 9364
rect 2050 9330 2055 9364
rect 2005 9318 2055 9330
rect 2005 9284 2021 9318
rect 2005 9258 2055 9284
rect 2005 9224 2015 9258
rect 2049 9234 2055 9258
rect 2005 9200 2021 9224
rect 2005 9150 2055 9200
rect 2005 9116 2021 9150
rect 2005 9091 2055 9116
rect 2089 9402 2219 9419
rect 2089 9368 2109 9402
rect 2143 9368 2177 9402
rect 2211 9368 2219 9402
rect 2089 9352 2219 9368
rect 2253 9408 2287 9454
rect 2089 9250 2127 9352
rect 2253 9318 2287 9374
rect 2161 9284 2177 9318
rect 2211 9316 2287 9318
rect 2211 9284 2253 9316
rect 2089 9234 2219 9250
rect 2089 9200 2109 9234
rect 2143 9200 2177 9234
rect 2211 9200 2219 9234
rect 2089 9184 2219 9200
rect 2253 9224 2287 9282
rect 2089 9082 2127 9184
rect 2253 9150 2287 9190
rect 2161 9116 2177 9150
rect 2211 9132 2287 9150
rect 2211 9116 2253 9132
rect 2089 9066 2219 9082
rect 1233 8864 1241 8898
rect 1233 8730 1275 8864
rect 1309 8989 1675 8998
rect 1309 8982 1317 8989
rect 1351 8955 1403 8989
rect 1437 8982 1675 8989
rect 1437 8955 1497 8982
rect 1343 8948 1497 8955
rect 1531 8948 1565 8982
rect 1667 8948 1675 8982
rect 1309 8814 1343 8948
rect 1481 8932 1675 8948
rect 1709 8948 1743 9006
rect 1937 8998 2055 9055
rect 2089 9032 2109 9066
rect 2143 9032 2177 9066
rect 2211 9032 2219 9066
rect 1309 8764 1343 8780
rect 1397 8898 1447 8914
rect 1431 8864 1447 8898
rect 1397 8814 1447 8864
rect 1431 8780 1447 8814
rect 1397 8746 1404 8780
rect 1438 8746 1447 8780
rect 1481 8830 1515 8932
rect 1777 8989 2143 8998
rect 1777 8982 2016 8989
rect 1777 8948 1785 8982
rect 1819 8948 1820 8982
rect 1887 8948 1921 8982
rect 1955 8955 2016 8982
rect 2050 8955 2102 8989
rect 2136 8982 2143 8989
rect 1955 8948 2109 8955
rect 1777 8932 1971 8948
rect 1709 8898 1743 8914
rect 1549 8864 1565 8898
rect 1599 8864 1633 8898
rect 1667 8864 1785 8898
rect 1819 8864 1853 8898
rect 1887 8864 1903 8898
rect 1709 8856 1743 8864
rect 1481 8814 1675 8830
rect 1481 8780 1497 8814
rect 1531 8780 1565 8814
rect 1599 8780 1633 8814
rect 1667 8780 1675 8814
rect 1481 8764 1675 8780
rect 1937 8830 1971 8932
rect 1709 8764 1743 8822
rect 1777 8814 1971 8830
rect 1777 8780 1785 8814
rect 1819 8780 1853 8814
rect 1887 8780 1921 8814
rect 1955 8780 1971 8814
rect 1777 8764 1971 8780
rect 2005 8898 2055 8914
rect 2005 8864 2021 8898
rect 2005 8814 2055 8864
rect 2005 8780 2021 8814
rect 2005 8779 2055 8780
rect 1233 8696 1241 8730
rect 1275 8696 1309 8730
rect 1343 8696 1359 8730
rect 1233 8680 1359 8696
rect 1397 8694 1447 8746
rect 2005 8745 2012 8779
rect 2046 8745 2055 8779
rect 2109 8814 2143 8948
rect 2109 8764 2143 8780
rect 2177 8898 2219 9032
rect 2211 8864 2219 8898
rect 1165 8591 1199 8638
rect 1397 8660 1404 8694
rect 1438 8660 1447 8694
rect 1549 8696 1565 8730
rect 1599 8696 1633 8730
rect 1667 8696 1785 8730
rect 1819 8696 1853 8730
rect 1887 8696 1903 8730
rect 1549 8680 1903 8696
rect 2005 8693 2055 8745
rect 2177 8730 2219 8864
rect 1397 8626 1447 8660
rect 1709 8672 1743 8680
rect 1709 8591 1743 8638
rect 2005 8659 2012 8693
rect 2046 8659 2055 8693
rect 2093 8696 2109 8730
rect 2143 8696 2177 8730
rect 2211 8696 2219 8730
rect 2093 8680 2219 8696
rect 2253 9040 2287 9098
rect 2253 8948 2287 9006
rect 2253 8856 2287 8914
rect 2253 8764 2287 8822
rect 2005 8626 2055 8659
rect 2253 8672 2287 8730
rect 2253 8591 2287 8638
rect 1165 8580 1367 8591
rect 1199 8573 1367 8580
rect 1199 8546 1245 8573
rect 1165 8539 1245 8546
rect 1279 8539 1313 8573
rect 1347 8539 1367 8573
rect 1479 8580 1973 8591
rect 1479 8573 1709 8580
rect 1479 8539 1497 8573
rect 1531 8539 1565 8573
rect 1599 8539 1633 8573
rect 1667 8546 1709 8573
rect 1743 8573 1973 8580
rect 1743 8546 1785 8573
rect 1667 8539 1785 8546
rect 1819 8539 1853 8573
rect 1887 8539 1921 8573
rect 1955 8539 1973 8573
rect 2085 8580 2287 8591
rect 2085 8573 2253 8580
rect 2085 8539 2105 8573
rect 2139 8539 2173 8573
rect 2207 8546 2253 8573
rect 2207 8539 2287 8546
rect 1165 8488 1199 8539
rect 1165 8419 1199 8454
rect 1233 8498 1675 8504
rect 1233 8489 1306 8498
rect 1233 8455 1271 8489
rect 1305 8463 1306 8489
rect 1341 8497 1675 8498
rect 1341 8470 1518 8497
rect 1552 8489 1675 8497
rect 1341 8463 1348 8470
rect 1305 8455 1348 8463
rect 1233 8453 1348 8455
rect 1494 8463 1518 8470
rect 1494 8455 1528 8463
rect 1562 8455 1609 8489
rect 1643 8455 1675 8489
rect 1494 8453 1675 8455
rect 1709 8488 1743 8539
rect 1381 8419 1397 8436
rect 1165 8403 1275 8419
rect 1165 8396 1241 8403
rect 1199 8369 1241 8396
rect 1199 8362 1275 8369
rect 1165 8353 1275 8362
rect 1309 8402 1397 8419
rect 1431 8419 1447 8436
rect 1709 8419 1743 8454
rect 1777 8497 2219 8504
rect 1777 8496 2109 8497
rect 1777 8489 1898 8496
rect 1777 8455 1809 8489
rect 1843 8455 1890 8489
rect 1932 8470 2109 8496
rect 1932 8462 1958 8470
rect 1924 8455 1958 8462
rect 1777 8453 1958 8455
rect 2104 8462 2109 8470
rect 2144 8489 2219 8497
rect 2144 8462 2147 8489
rect 2104 8455 2147 8462
rect 2181 8455 2219 8489
rect 2104 8453 2219 8455
rect 2253 8488 2287 8539
rect 2005 8419 2021 8436
rect 1431 8402 1523 8419
rect 1309 8385 1523 8402
rect 1165 8304 1199 8353
rect 1309 8310 1343 8385
rect 1233 8276 1254 8310
rect 1288 8276 1343 8310
rect 1379 8312 1453 8329
rect 1379 8278 1397 8312
rect 1431 8278 1453 8312
rect 1165 8241 1199 8270
rect 1379 8258 1453 8278
rect 1489 8310 1523 8385
rect 1557 8403 1895 8419
rect 1591 8369 1625 8403
rect 1659 8396 1793 8403
rect 1659 8369 1709 8396
rect 1557 8362 1709 8369
rect 1743 8369 1793 8396
rect 1827 8369 1861 8403
rect 1743 8362 1895 8369
rect 1557 8353 1895 8362
rect 1929 8402 2021 8419
rect 2055 8419 2071 8436
rect 2253 8419 2287 8454
rect 2055 8402 2143 8419
rect 1929 8385 2143 8402
rect 1489 8276 1557 8310
rect 1591 8276 1625 8310
rect 1659 8276 1675 8310
rect 1709 8304 1743 8353
rect 1929 8310 1963 8385
rect 1777 8276 1793 8310
rect 1827 8276 1861 8310
rect 1895 8276 1963 8310
rect 1999 8313 2073 8329
rect 1999 8312 2022 8313
rect 1999 8278 2021 8312
rect 2056 8279 2073 8313
rect 2055 8278 2073 8279
rect 1709 8241 1743 8270
rect 1999 8258 2073 8278
rect 2109 8310 2143 8385
rect 2177 8403 2287 8419
rect 2211 8396 2287 8403
rect 2211 8369 2253 8396
rect 2177 8362 2253 8369
rect 2177 8353 2287 8362
rect 2109 8276 2164 8310
rect 2198 8276 2219 8310
rect 2253 8304 2287 8353
rect 2253 8241 2287 8270
rect -3752 7990 -3656 8024
rect -3282 7990 -3186 8024
rect -3752 7928 -3718 7990
rect -3220 7928 -3186 7990
rect -3718 7876 -3557 7910
rect -3381 7876 -3365 7910
rect -3650 7862 -3616 7876
rect -3650 7812 -3616 7828
rect -3573 7780 -3557 7814
rect -3381 7780 -3365 7814
rect -3322 7766 -3288 7782
rect -3650 7670 -3616 7686
rect -3573 7684 -3557 7718
rect -3381 7684 -3365 7718
rect -3322 7716 -3288 7732
rect -3650 7620 -3616 7636
rect -3573 7588 -3557 7622
rect -3381 7588 -3365 7622
rect -3322 7574 -3288 7590
rect -3650 7478 -3616 7494
rect -3573 7492 -3557 7526
rect -3381 7492 -3365 7526
rect -3322 7524 -3288 7540
rect -3650 7428 -3616 7444
rect -3573 7396 -3557 7430
rect -3381 7396 -3365 7430
rect -3322 7382 -3288 7398
rect -3650 7286 -3616 7302
rect -3573 7300 -3557 7334
rect -3381 7300 -3365 7334
rect -3322 7332 -3288 7348
rect -3650 7236 -3616 7252
rect -3573 7204 -3557 7238
rect -3381 7204 -3365 7238
rect -3322 7190 -3288 7206
rect -3650 7094 -3616 7110
rect -3573 7108 -3557 7142
rect -3381 7108 -3365 7142
rect -3322 7140 -3288 7156
rect -3650 7044 -3616 7060
rect -3573 7012 -3557 7046
rect -3381 7012 -3365 7046
rect -3322 6998 -3288 7014
rect -3650 6902 -3616 6918
rect -3573 6916 -3557 6950
rect -3381 6916 -3365 6950
rect -3322 6948 -3288 6964
rect -3650 6852 -3616 6868
rect -3573 6820 -3557 6854
rect -3381 6820 -3365 6854
rect -3322 6806 -3288 6822
rect -3650 6710 -3616 6726
rect -3573 6724 -3557 6758
rect -3381 6724 -3365 6758
rect -3322 6756 -3288 6772
rect -3650 6660 -3616 6676
rect -3573 6628 -3557 6662
rect -3381 6628 -3365 6662
rect -3322 6614 -3288 6630
rect -3650 6518 -3616 6534
rect -3573 6532 -3557 6566
rect -3381 6532 -3365 6566
rect -3322 6564 -3288 6580
rect -3650 6468 -3616 6484
rect -3573 6436 -3557 6470
rect -3381 6436 -3365 6470
rect -3322 6422 -3288 6438
rect -3650 6326 -3616 6342
rect -3573 6340 -3557 6374
rect -3381 6340 -3365 6374
rect -3322 6372 -3288 6388
rect -3650 6276 -3616 6292
rect -3573 6244 -3557 6278
rect -3381 6244 -3365 6278
rect -3322 6230 -3288 6246
rect -3322 6182 -3288 6196
rect -3573 6148 -3557 6182
rect -3381 6148 -3220 6182
rect -3752 6068 -3718 6130
rect -2758 7989 -2662 8023
rect 6114 7989 6210 8023
rect -2758 7927 -2724 7989
rect 6176 7927 6210 7989
rect -2402 7887 -2386 7921
rect -2352 7887 -2336 7921
rect -1982 7887 -1966 7921
rect -1932 7887 -1916 7921
rect -1562 7887 -1546 7921
rect -1512 7887 -1496 7921
rect -1142 7887 -1126 7921
rect -1092 7887 -1076 7921
rect -722 7887 -706 7921
rect -672 7887 -656 7921
rect -302 7887 -286 7921
rect -252 7887 -236 7921
rect 118 7887 134 7921
rect 168 7887 184 7921
rect 538 7887 554 7921
rect 588 7887 604 7921
rect 958 7887 974 7921
rect 1008 7887 1024 7921
rect 1378 7887 1394 7921
rect 1428 7887 1444 7921
rect 1798 7887 1814 7921
rect 1848 7887 1864 7921
rect 2218 7887 2234 7921
rect 2268 7887 2284 7921
rect 2638 7887 2654 7921
rect 2688 7887 2704 7921
rect 3058 7887 3074 7921
rect 3108 7887 3124 7921
rect 3478 7887 3494 7921
rect 3528 7887 3544 7921
rect 3898 7887 3914 7921
rect 3948 7887 3964 7921
rect 4318 7887 4334 7921
rect 4368 7887 4384 7921
rect 4738 7887 4754 7921
rect 4788 7887 4804 7921
rect 5158 7887 5174 7921
rect 5208 7887 5224 7921
rect 5578 7887 5594 7921
rect 5628 7887 5644 7921
rect 5966 7887 6014 7921
rect 6048 7887 6176 7921
rect -2644 7828 -2610 7844
rect -2644 7593 -2610 7652
rect -2548 7828 -2514 7844
rect -2548 7593 -2514 7652
rect -2434 7828 -2400 7844
rect -2434 7636 -2400 7652
rect -2338 7828 -2304 7844
rect -2338 7636 -2304 7652
rect -2224 7828 -2190 7844
rect -2224 7636 -2190 7652
rect -2128 7828 -2094 7844
rect -2128 7636 -2094 7652
rect -2014 7828 -1980 7844
rect -2014 7636 -1980 7652
rect -1918 7828 -1884 7844
rect -1918 7636 -1884 7652
rect -1804 7828 -1770 7844
rect -1804 7636 -1770 7652
rect -1708 7828 -1674 7844
rect -1708 7636 -1674 7652
rect -1594 7828 -1560 7844
rect -1594 7636 -1560 7652
rect -1498 7828 -1464 7844
rect -1498 7636 -1464 7652
rect -1384 7828 -1350 7844
rect -1384 7636 -1350 7652
rect -1288 7828 -1254 7844
rect -1288 7636 -1254 7652
rect -1174 7828 -1140 7844
rect -1174 7636 -1140 7652
rect -1078 7828 -1044 7844
rect -1078 7636 -1044 7652
rect -964 7828 -930 7844
rect -964 7636 -930 7652
rect -868 7828 -834 7844
rect -868 7636 -834 7652
rect -754 7828 -720 7844
rect -754 7636 -720 7652
rect -658 7828 -624 7844
rect -658 7636 -624 7652
rect -544 7828 -510 7844
rect -544 7636 -510 7652
rect -448 7828 -414 7844
rect -448 7636 -414 7652
rect -334 7828 -300 7844
rect -334 7636 -300 7652
rect -238 7828 -204 7844
rect -238 7636 -204 7652
rect -124 7828 -90 7844
rect -124 7636 -90 7652
rect -28 7828 6 7844
rect -28 7636 6 7652
rect 86 7828 120 7844
rect 86 7636 120 7652
rect 182 7828 216 7844
rect 182 7636 216 7652
rect 296 7828 330 7844
rect 296 7636 330 7652
rect 392 7828 426 7844
rect 392 7636 426 7652
rect 506 7828 540 7844
rect 506 7636 540 7652
rect 602 7828 636 7844
rect 602 7636 636 7652
rect 716 7828 750 7844
rect 716 7636 750 7652
rect 812 7828 846 7844
rect 812 7636 846 7652
rect 926 7828 960 7844
rect 926 7636 960 7652
rect 1022 7828 1056 7844
rect 1022 7636 1056 7652
rect 1136 7828 1170 7844
rect 1136 7636 1170 7652
rect 1232 7828 1266 7844
rect 1232 7636 1266 7652
rect 1346 7828 1380 7844
rect 1346 7636 1380 7652
rect 1442 7828 1476 7844
rect 1442 7636 1476 7652
rect 1556 7828 1590 7844
rect 1556 7636 1590 7652
rect 1652 7828 1686 7844
rect 1652 7636 1686 7652
rect 1766 7828 1800 7844
rect 1766 7636 1800 7652
rect 1862 7828 1896 7844
rect 1862 7636 1896 7652
rect 1976 7828 2010 7844
rect 1976 7636 2010 7652
rect 2072 7828 2106 7844
rect 2072 7636 2106 7652
rect 2186 7828 2220 7844
rect 2186 7636 2220 7652
rect 2282 7828 2316 7844
rect 2282 7636 2316 7652
rect 2396 7828 2430 7844
rect 2396 7636 2430 7652
rect 2492 7828 2526 7844
rect 2492 7636 2526 7652
rect 2606 7828 2640 7844
rect 2606 7636 2640 7652
rect 2702 7828 2736 7844
rect 2702 7636 2736 7652
rect 2816 7828 2850 7844
rect 2816 7636 2850 7652
rect 2912 7828 2946 7844
rect 2912 7636 2946 7652
rect 3026 7828 3060 7844
rect 3026 7636 3060 7652
rect 3122 7828 3156 7844
rect 3122 7636 3156 7652
rect 3236 7828 3270 7844
rect 3236 7636 3270 7652
rect 3332 7828 3366 7844
rect 3332 7636 3366 7652
rect 3446 7828 3480 7844
rect 3446 7636 3480 7652
rect 3542 7828 3576 7844
rect 3542 7636 3576 7652
rect 3656 7828 3690 7844
rect 3656 7636 3690 7652
rect 3752 7828 3786 7844
rect 3752 7636 3786 7652
rect 3866 7828 3900 7844
rect 3866 7636 3900 7652
rect 3962 7828 3996 7844
rect 3962 7636 3996 7652
rect 4076 7828 4110 7844
rect 4076 7636 4110 7652
rect 4172 7828 4206 7844
rect 4172 7636 4206 7652
rect 4286 7828 4320 7844
rect 4286 7636 4320 7652
rect 4382 7828 4416 7844
rect 4382 7636 4416 7652
rect 4496 7828 4530 7844
rect 4496 7636 4530 7652
rect 4592 7828 4626 7844
rect 4592 7636 4626 7652
rect 4706 7828 4740 7844
rect 4706 7636 4740 7652
rect 4802 7828 4836 7844
rect 4802 7636 4836 7652
rect 4916 7828 4950 7844
rect 4916 7636 4950 7652
rect 5012 7828 5046 7844
rect 5012 7636 5046 7652
rect 5126 7828 5160 7844
rect 5126 7636 5160 7652
rect 5222 7828 5256 7844
rect 5222 7636 5256 7652
rect 5336 7828 5370 7844
rect 5336 7636 5370 7652
rect 5432 7828 5466 7844
rect 5432 7636 5466 7652
rect 5546 7828 5580 7844
rect 5546 7636 5580 7652
rect 5642 7828 5676 7844
rect 5642 7636 5676 7652
rect 5756 7828 5790 7844
rect 5756 7636 5790 7652
rect 5852 7828 5886 7844
rect 5852 7636 5886 7652
rect 5966 7828 6000 7887
rect 5966 7636 6000 7652
rect 6062 7828 6096 7887
rect 6062 7636 6096 7652
rect -2724 7559 -2596 7593
rect -2562 7559 -2514 7593
rect -2192 7559 -2176 7593
rect -2142 7559 -2126 7593
rect -1772 7559 -1756 7593
rect -1722 7559 -1706 7593
rect -1352 7559 -1336 7593
rect -1302 7559 -1286 7593
rect -932 7559 -916 7593
rect -882 7559 -866 7593
rect -512 7559 -496 7593
rect -462 7559 -446 7593
rect -92 7559 -76 7593
rect -42 7559 -26 7593
rect 328 7559 344 7593
rect 378 7559 394 7593
rect 748 7559 764 7593
rect 798 7559 814 7593
rect 1168 7559 1184 7593
rect 1218 7559 1234 7593
rect 1588 7559 1604 7593
rect 1638 7559 1654 7593
rect 2008 7559 2024 7593
rect 2058 7559 2074 7593
rect 2428 7559 2444 7593
rect 2478 7559 2494 7593
rect 2848 7559 2864 7593
rect 2898 7559 2914 7593
rect 3268 7559 3284 7593
rect 3318 7559 3334 7593
rect 3688 7559 3704 7593
rect 3738 7559 3754 7593
rect 4108 7559 4124 7593
rect 4158 7559 4174 7593
rect 4528 7559 4544 7593
rect 4578 7559 4594 7593
rect 4948 7559 4964 7593
rect 4998 7559 5014 7593
rect 5368 7559 5384 7593
rect 5418 7559 5434 7593
rect 5788 7559 5804 7593
rect 5838 7559 5854 7593
rect -2758 7395 -2724 7553
rect 6176 7395 6210 7553
rect -2400 7355 -2384 7389
rect -2350 7355 -2334 7389
rect -1980 7355 -1964 7389
rect -1930 7355 -1914 7389
rect -1560 7355 -1544 7389
rect -1510 7355 -1494 7389
rect -1140 7355 -1124 7389
rect -1090 7355 -1074 7389
rect -720 7355 -704 7389
rect -670 7355 -654 7389
rect -300 7355 -284 7389
rect -250 7355 -234 7389
rect 120 7355 136 7389
rect 170 7355 186 7389
rect 540 7355 556 7389
rect 590 7355 606 7389
rect 960 7355 976 7389
rect 1010 7355 1026 7389
rect 1380 7355 1396 7389
rect 1430 7355 1446 7389
rect 1800 7355 1816 7389
rect 1850 7355 1866 7389
rect 2220 7355 2236 7389
rect 2270 7355 2286 7389
rect 2640 7355 2656 7389
rect 2690 7355 2706 7389
rect 3060 7355 3076 7389
rect 3110 7355 3126 7389
rect 3480 7355 3496 7389
rect 3530 7355 3546 7389
rect 3900 7355 3916 7389
rect 3950 7355 3966 7389
rect 4320 7355 4336 7389
rect 4370 7355 4386 7389
rect 4740 7355 4756 7389
rect 4790 7355 4806 7389
rect 5160 7355 5176 7389
rect 5210 7355 5226 7389
rect 5580 7355 5596 7389
rect 5630 7355 5646 7389
rect 5968 7355 6016 7389
rect 6050 7355 6176 7389
rect -2642 7295 -2608 7311
rect -2642 7060 -2608 7119
rect -2546 7295 -2512 7311
rect -2546 7060 -2512 7119
rect -2432 7296 -2398 7311
rect -2432 7103 -2398 7119
rect -2336 7295 -2302 7311
rect -2336 7103 -2302 7119
rect -2222 7296 -2188 7311
rect -2222 7103 -2188 7119
rect -2126 7295 -2092 7311
rect -2126 7103 -2092 7119
rect -2012 7296 -1978 7311
rect -2012 7103 -1978 7119
rect -1916 7295 -1882 7311
rect -1916 7103 -1882 7119
rect -1802 7296 -1768 7311
rect -1802 7103 -1768 7119
rect -1706 7295 -1672 7311
rect -1706 7103 -1672 7119
rect -1592 7296 -1558 7311
rect -1592 7103 -1558 7119
rect -1496 7295 -1462 7311
rect -1496 7103 -1462 7119
rect -1382 7296 -1348 7311
rect -1382 7103 -1348 7119
rect -1286 7295 -1252 7311
rect -1286 7103 -1252 7119
rect -1172 7296 -1138 7311
rect -1172 7103 -1138 7119
rect -1076 7295 -1042 7311
rect -1076 7103 -1042 7119
rect -962 7296 -928 7311
rect -962 7103 -928 7119
rect -866 7295 -832 7311
rect -866 7103 -832 7119
rect -752 7296 -718 7311
rect -752 7103 -718 7119
rect -656 7295 -622 7311
rect -656 7103 -622 7119
rect -542 7296 -508 7311
rect -542 7103 -508 7119
rect -446 7295 -412 7311
rect -446 7103 -412 7119
rect -332 7296 -298 7311
rect -332 7103 -298 7119
rect -236 7295 -202 7311
rect -236 7103 -202 7119
rect -122 7296 -88 7311
rect -122 7103 -88 7119
rect -26 7295 8 7311
rect -26 7103 8 7119
rect 88 7296 122 7311
rect 88 7103 122 7119
rect 184 7295 218 7311
rect 184 7103 218 7119
rect 298 7296 332 7311
rect 298 7103 332 7119
rect 394 7295 428 7311
rect 394 7103 428 7119
rect 508 7296 542 7311
rect 508 7103 542 7119
rect 604 7295 638 7311
rect 604 7103 638 7119
rect 718 7296 752 7311
rect 718 7103 752 7119
rect 814 7295 848 7311
rect 814 7103 848 7119
rect 928 7296 962 7311
rect 928 7103 962 7119
rect 1024 7295 1058 7311
rect 1024 7103 1058 7119
rect 1138 7296 1172 7311
rect 1138 7103 1172 7119
rect 1234 7295 1268 7311
rect 1234 7103 1268 7119
rect 1348 7296 1382 7311
rect 1348 7103 1382 7119
rect 1444 7295 1478 7311
rect 1444 7103 1478 7119
rect 1558 7296 1592 7311
rect 1558 7103 1592 7119
rect 1654 7295 1688 7311
rect 1654 7103 1688 7119
rect 1768 7296 1802 7311
rect 1768 7103 1802 7119
rect 1864 7295 1898 7311
rect 1864 7103 1898 7119
rect 1978 7296 2012 7311
rect 1978 7103 2012 7119
rect 2074 7295 2108 7311
rect 2074 7103 2108 7119
rect 2188 7296 2222 7311
rect 2188 7103 2222 7119
rect 2284 7295 2318 7311
rect 2284 7103 2318 7119
rect 2398 7296 2432 7311
rect 2398 7103 2432 7119
rect 2494 7295 2528 7311
rect 2494 7103 2528 7119
rect 2608 7296 2642 7311
rect 2608 7103 2642 7119
rect 2704 7295 2738 7311
rect 2704 7103 2738 7119
rect 2818 7296 2852 7311
rect 2818 7103 2852 7119
rect 2914 7295 2948 7311
rect 2914 7103 2948 7119
rect 3028 7296 3062 7311
rect 3028 7103 3062 7119
rect 3124 7295 3158 7311
rect 3124 7103 3158 7119
rect 3238 7296 3272 7311
rect 3238 7103 3272 7119
rect 3334 7295 3368 7311
rect 3334 7103 3368 7119
rect 3448 7296 3482 7311
rect 3448 7103 3482 7119
rect 3544 7295 3578 7311
rect 3544 7103 3578 7119
rect 3658 7296 3692 7311
rect 3658 7103 3692 7119
rect 3754 7295 3788 7311
rect 3754 7103 3788 7119
rect 3868 7296 3902 7311
rect 3868 7103 3902 7119
rect 3964 7295 3998 7311
rect 3964 7103 3998 7119
rect 4078 7296 4112 7311
rect 4078 7103 4112 7119
rect 4174 7295 4208 7311
rect 4174 7103 4208 7119
rect 4288 7296 4322 7311
rect 4288 7103 4322 7119
rect 4384 7295 4418 7311
rect 4384 7103 4418 7119
rect 4498 7296 4532 7311
rect 4498 7103 4532 7119
rect 4594 7295 4628 7311
rect 4594 7103 4628 7119
rect 4708 7296 4742 7311
rect 4708 7103 4742 7119
rect 4804 7295 4838 7311
rect 4804 7103 4838 7119
rect 4918 7296 4952 7311
rect 4918 7103 4952 7119
rect 5014 7295 5048 7311
rect 5014 7103 5048 7119
rect 5128 7296 5162 7311
rect 5128 7103 5162 7119
rect 5224 7295 5258 7311
rect 5224 7103 5258 7119
rect 5338 7296 5372 7311
rect 5338 7103 5372 7119
rect 5434 7295 5468 7311
rect 5434 7103 5468 7119
rect 5548 7296 5582 7311
rect 5548 7103 5582 7119
rect 5644 7295 5678 7311
rect 5644 7103 5678 7119
rect 5758 7296 5792 7311
rect 5758 7103 5792 7119
rect 5854 7295 5888 7311
rect 5854 7103 5888 7119
rect 5968 7295 6002 7355
rect 5968 7103 6002 7119
rect 6064 7295 6098 7355
rect 6064 7103 6098 7119
rect -2724 7026 -2594 7060
rect -2560 7026 -2512 7060
rect -2190 7026 -2174 7060
rect -2140 7026 -2124 7060
rect -1770 7026 -1754 7060
rect -1720 7026 -1704 7060
rect -1350 7026 -1334 7060
rect -1300 7026 -1284 7060
rect -930 7026 -914 7060
rect -880 7026 -864 7060
rect -510 7026 -494 7060
rect -460 7026 -444 7060
rect -90 7026 -74 7060
rect -40 7026 -24 7060
rect 330 7026 346 7060
rect 380 7026 396 7060
rect 750 7026 766 7060
rect 800 7026 816 7060
rect 1170 7026 1186 7060
rect 1220 7026 1236 7060
rect 1590 7026 1606 7060
rect 1640 7026 1656 7060
rect 2010 7026 2026 7060
rect 2060 7026 2076 7060
rect 2430 7026 2446 7060
rect 2480 7026 2496 7060
rect 2850 7026 2866 7060
rect 2900 7026 2916 7060
rect 3270 7026 3286 7060
rect 3320 7026 3336 7060
rect 3690 7026 3706 7060
rect 3740 7026 3756 7060
rect 4110 7026 4126 7060
rect 4160 7026 4176 7060
rect 4530 7026 4546 7060
rect 4580 7026 4596 7060
rect 4950 7026 4966 7060
rect 5000 7026 5016 7060
rect 5370 7026 5386 7060
rect 5420 7026 5436 7060
rect 5790 7026 5806 7060
rect 5840 7026 5856 7060
rect -2758 6958 -2724 7020
rect 6176 6958 6210 7020
rect -2758 6924 -2662 6958
rect 6114 6924 6210 6958
rect 6648 7990 6744 8024
rect 7118 7990 7214 8024
rect 6648 7928 6682 7990
rect -3220 6068 -3186 6130
rect -3752 6034 -3656 6068
rect -3282 6034 -3186 6068
rect -2744 6497 -2648 6531
rect 6130 6497 6226 6531
rect -2744 6435 -2710 6497
rect -3750 5613 -3654 5614
rect -3750 5580 -3656 5613
rect -3280 5580 -3184 5614
rect -3750 5518 -3716 5580
rect -3218 5518 -3184 5580
rect -3716 5466 -3555 5500
rect -3379 5466 -3363 5500
rect -3648 5452 -3614 5466
rect -3648 5402 -3614 5418
rect -3571 5370 -3555 5404
rect -3379 5370 -3363 5404
rect -3320 5356 -3286 5372
rect -3571 5307 -3555 5308
rect -3648 5260 -3614 5276
rect -3571 5274 -3557 5307
rect -3379 5274 -3363 5308
rect -3320 5306 -3286 5322
rect -3648 5210 -3614 5226
rect -3571 5178 -3555 5212
rect -3379 5178 -3363 5212
rect -3320 5164 -3286 5180
rect -3571 5115 -3555 5116
rect -3648 5068 -3614 5084
rect -3571 5082 -3557 5115
rect -3379 5082 -3363 5116
rect -3320 5114 -3286 5130
rect -3648 5018 -3614 5034
rect -3571 4986 -3555 5020
rect -3379 4986 -3363 5020
rect -3320 4972 -3286 4988
rect -3571 4923 -3555 4924
rect -3648 4876 -3614 4892
rect -3571 4890 -3557 4923
rect -3379 4890 -3363 4924
rect -3320 4922 -3286 4938
rect -3648 4826 -3614 4842
rect -3571 4794 -3555 4828
rect -3379 4794 -3363 4828
rect -3320 4780 -3286 4796
rect -3571 4731 -3555 4732
rect -3648 4684 -3614 4700
rect -3571 4698 -3557 4731
rect -3379 4698 -3363 4732
rect -3320 4730 -3286 4746
rect -3648 4634 -3614 4650
rect -3571 4602 -3555 4636
rect -3379 4602 -3363 4636
rect -3320 4588 -3286 4604
rect -3571 4539 -3555 4540
rect -3648 4492 -3614 4508
rect -3571 4506 -3557 4539
rect -3379 4506 -3363 4540
rect -3320 4538 -3286 4554
rect -3648 4442 -3614 4458
rect -3571 4410 -3555 4444
rect -3379 4410 -3363 4444
rect -3320 4396 -3286 4412
rect -3571 4347 -3555 4348
rect -3648 4300 -3614 4316
rect -3571 4314 -3557 4347
rect -3379 4314 -3363 4348
rect -3320 4346 -3286 4362
rect -3648 4250 -3614 4266
rect -3571 4218 -3555 4252
rect -3379 4218 -3363 4252
rect -3320 4204 -3286 4220
rect -3571 4155 -3555 4156
rect -3648 4108 -3614 4124
rect -3571 4122 -3557 4155
rect -3379 4122 -3363 4156
rect -3320 4154 -3286 4170
rect -3648 4058 -3614 4074
rect -3571 4026 -3555 4060
rect -3379 4026 -3363 4060
rect -3320 4012 -3286 4028
rect -3571 3963 -3555 3964
rect -3648 3916 -3614 3932
rect -3571 3930 -3557 3963
rect -3379 3930 -3363 3964
rect -3320 3962 -3286 3978
rect -3648 3866 -3614 3882
rect -3571 3834 -3555 3868
rect -3379 3834 -3363 3868
rect -3320 3820 -3286 3836
rect -3320 3772 -3286 3786
rect -3571 3738 -3555 3772
rect -3379 3738 -3218 3772
rect -3750 3658 -3716 3720
rect 6192 6435 6226 6497
rect -2388 6395 -2372 6429
rect -2338 6395 -2322 6429
rect -1968 6395 -1952 6429
rect -1918 6395 -1902 6429
rect -1548 6395 -1532 6429
rect -1498 6395 -1482 6429
rect -1128 6395 -1112 6429
rect -1078 6395 -1062 6429
rect -708 6395 -692 6429
rect -658 6395 -642 6429
rect -288 6395 -272 6429
rect -238 6395 -222 6429
rect 132 6395 148 6429
rect 182 6395 198 6429
rect 552 6395 568 6429
rect 602 6395 618 6429
rect 972 6395 988 6429
rect 1022 6395 1038 6429
rect 1392 6395 1408 6429
rect 1442 6395 1458 6429
rect 1812 6395 1828 6429
rect 1862 6395 1878 6429
rect 2232 6395 2248 6429
rect 2282 6395 2298 6429
rect 2652 6395 2668 6429
rect 2702 6395 2718 6429
rect 3072 6395 3088 6429
rect 3122 6395 3138 6429
rect 3492 6395 3508 6429
rect 3542 6395 3558 6429
rect 3912 6395 3928 6429
rect 3962 6395 3978 6429
rect 4332 6395 4348 6429
rect 4382 6395 4398 6429
rect 4752 6395 4768 6429
rect 4802 6395 4818 6429
rect 5172 6395 5188 6429
rect 5222 6395 5238 6429
rect 5592 6395 5608 6429
rect 5642 6395 5658 6429
rect 5980 6395 6028 6429
rect 6062 6395 6192 6429
rect -2630 6345 -2596 6361
rect -2630 6119 -2596 6169
rect -2534 6345 -2500 6361
rect -2534 6119 -2500 6169
rect -2420 6345 -2386 6361
rect -2420 6153 -2386 6169
rect -2324 6345 -2290 6361
rect -2324 6153 -2290 6169
rect -2210 6345 -2176 6361
rect -2210 6153 -2176 6169
rect -2114 6345 -2080 6361
rect -2114 6153 -2080 6169
rect -2000 6345 -1966 6361
rect -2000 6153 -1966 6169
rect -1904 6345 -1870 6361
rect -1904 6153 -1870 6169
rect -1790 6345 -1756 6361
rect -1790 6153 -1756 6169
rect -1694 6345 -1660 6361
rect -1694 6153 -1660 6169
rect -1580 6345 -1546 6361
rect -1580 6153 -1546 6169
rect -1484 6345 -1450 6361
rect -1484 6153 -1450 6169
rect -1370 6345 -1336 6361
rect -1370 6153 -1336 6169
rect -1274 6345 -1240 6361
rect -1274 6153 -1240 6169
rect -1160 6345 -1126 6361
rect -1160 6153 -1126 6169
rect -1064 6345 -1030 6361
rect -1064 6153 -1030 6169
rect -950 6345 -916 6361
rect -950 6153 -916 6169
rect -854 6345 -820 6361
rect -854 6153 -820 6169
rect -740 6345 -706 6361
rect -740 6153 -706 6169
rect -644 6345 -610 6361
rect -644 6153 -610 6169
rect -530 6345 -496 6361
rect -530 6153 -496 6169
rect -434 6345 -400 6361
rect -434 6153 -400 6169
rect -320 6345 -286 6361
rect -320 6153 -286 6169
rect -224 6345 -190 6361
rect -224 6153 -190 6169
rect -110 6345 -76 6361
rect -110 6153 -76 6169
rect -14 6345 20 6361
rect -14 6153 20 6169
rect 100 6345 134 6361
rect 100 6153 134 6169
rect 196 6345 230 6361
rect 196 6153 230 6169
rect 310 6345 344 6361
rect 310 6153 344 6169
rect 406 6345 440 6361
rect 406 6153 440 6169
rect 520 6345 554 6361
rect 520 6153 554 6169
rect 616 6345 650 6361
rect 616 6153 650 6169
rect 730 6345 764 6361
rect 730 6153 764 6169
rect 826 6345 860 6361
rect 826 6153 860 6169
rect 940 6345 974 6361
rect 940 6153 974 6169
rect 1036 6345 1070 6361
rect 1036 6153 1070 6169
rect 1150 6345 1184 6361
rect 1150 6153 1184 6169
rect 1246 6345 1280 6361
rect 1246 6153 1280 6169
rect 1360 6345 1394 6361
rect 1360 6153 1394 6169
rect 1456 6345 1490 6361
rect 1456 6153 1490 6169
rect 1570 6345 1604 6361
rect 1570 6153 1604 6169
rect 1666 6345 1700 6361
rect 1666 6153 1700 6169
rect 1780 6345 1814 6361
rect 1780 6153 1814 6169
rect 1876 6345 1910 6361
rect 1876 6153 1910 6169
rect 1990 6345 2024 6361
rect 1990 6153 2024 6169
rect 2086 6345 2120 6361
rect 2086 6153 2120 6169
rect 2200 6345 2234 6361
rect 2200 6153 2234 6169
rect 2296 6345 2330 6361
rect 2296 6153 2330 6169
rect 2410 6345 2444 6361
rect 2410 6153 2444 6169
rect 2506 6345 2540 6361
rect 2506 6153 2540 6169
rect 2620 6345 2654 6361
rect 2620 6153 2654 6169
rect 2716 6345 2750 6361
rect 2716 6153 2750 6169
rect 2830 6345 2864 6361
rect 2830 6153 2864 6169
rect 2926 6345 2960 6361
rect 2926 6153 2960 6169
rect 3040 6345 3074 6361
rect 3040 6153 3074 6169
rect 3136 6345 3170 6361
rect 3136 6153 3170 6169
rect 3250 6345 3284 6361
rect 3250 6153 3284 6169
rect 3346 6345 3380 6361
rect 3346 6153 3380 6169
rect 3460 6345 3494 6361
rect 3460 6153 3494 6169
rect 3556 6345 3590 6361
rect 3556 6153 3590 6169
rect 3670 6345 3704 6361
rect 3670 6153 3704 6169
rect 3766 6345 3800 6361
rect 3766 6153 3800 6169
rect 3880 6345 3914 6361
rect 3880 6153 3914 6169
rect 3976 6345 4010 6361
rect 3976 6153 4010 6169
rect 4090 6345 4124 6361
rect 4090 6153 4124 6169
rect 4186 6345 4220 6361
rect 4186 6153 4220 6169
rect 4300 6345 4334 6361
rect 4300 6153 4334 6169
rect 4396 6345 4430 6361
rect 4396 6153 4430 6169
rect 4510 6345 4544 6361
rect 4510 6153 4544 6169
rect 4606 6345 4640 6361
rect 4606 6153 4640 6169
rect 4720 6345 4754 6361
rect 4720 6153 4754 6169
rect 4816 6345 4850 6361
rect 4816 6153 4850 6169
rect 4930 6345 4964 6361
rect 4930 6153 4964 6169
rect 5026 6345 5060 6361
rect 5026 6153 5060 6169
rect 5140 6345 5174 6361
rect 5140 6153 5174 6169
rect 5236 6345 5270 6361
rect 5236 6153 5270 6169
rect 5350 6345 5384 6361
rect 5350 6153 5384 6169
rect 5446 6345 5480 6361
rect 5446 6153 5480 6169
rect 5560 6345 5594 6361
rect 5560 6153 5594 6169
rect 5656 6345 5690 6361
rect 5656 6153 5690 6169
rect 5770 6345 5804 6361
rect 5770 6153 5804 6169
rect 5866 6345 5900 6361
rect 5866 6153 5900 6169
rect 5980 6345 6014 6395
rect 5980 6153 6014 6169
rect 6076 6345 6110 6395
rect 6076 6153 6110 6169
rect -2710 6085 -2582 6119
rect -2548 6085 -2500 6119
rect -2178 6085 -2162 6119
rect -2128 6085 -2112 6119
rect -1758 6085 -1742 6119
rect -1708 6085 -1692 6119
rect -1338 6085 -1322 6119
rect -1288 6085 -1272 6119
rect -918 6085 -902 6119
rect -868 6085 -852 6119
rect -498 6085 -482 6119
rect -448 6085 -432 6119
rect -78 6085 -62 6119
rect -28 6085 -12 6119
rect 342 6085 358 6119
rect 392 6085 408 6119
rect 762 6085 778 6119
rect 812 6085 828 6119
rect 1182 6085 1198 6119
rect 1232 6085 1248 6119
rect 1602 6085 1618 6119
rect 1652 6085 1668 6119
rect 2022 6085 2038 6119
rect 2072 6085 2088 6119
rect 2442 6085 2458 6119
rect 2492 6085 2508 6119
rect 2862 6085 2878 6119
rect 2912 6085 2928 6119
rect 3282 6085 3298 6119
rect 3332 6085 3348 6119
rect 3702 6085 3718 6119
rect 3752 6085 3768 6119
rect 4122 6085 4138 6119
rect 4172 6085 4188 6119
rect 4542 6085 4558 6119
rect 4592 6085 4608 6119
rect 4962 6085 4978 6119
rect 5012 6085 5028 6119
rect 5382 6085 5398 6119
rect 5432 6085 5448 6119
rect 5802 6085 5818 6119
rect 5852 6085 5868 6119
rect -2388 5955 -2372 5989
rect -2338 5955 -2322 5989
rect -1968 5955 -1952 5989
rect -1918 5955 -1902 5989
rect -1548 5955 -1532 5989
rect -1498 5955 -1482 5989
rect -1128 5955 -1112 5989
rect -1078 5955 -1062 5989
rect -708 5955 -692 5989
rect -658 5955 -642 5989
rect -288 5955 -272 5989
rect -238 5955 -222 5989
rect 132 5955 148 5989
rect 182 5955 198 5989
rect 552 5955 568 5989
rect 602 5955 618 5989
rect 972 5955 988 5989
rect 1022 5955 1038 5989
rect 1392 5955 1408 5989
rect 1442 5955 1458 5989
rect 1812 5955 1828 5989
rect 1862 5955 1878 5989
rect 2232 5955 2248 5989
rect 2282 5955 2298 5989
rect 2652 5955 2668 5989
rect 2702 5955 2718 5989
rect 3072 5955 3088 5989
rect 3122 5955 3138 5989
rect 3492 5955 3508 5989
rect 3542 5955 3558 5989
rect 3912 5955 3928 5989
rect 3962 5955 3978 5989
rect 4332 5955 4348 5989
rect 4382 5955 4398 5989
rect 4752 5955 4768 5989
rect 4802 5955 4818 5989
rect 5172 5955 5188 5989
rect 5222 5955 5238 5989
rect 5592 5955 5608 5989
rect 5642 5955 5658 5989
rect 5980 5955 6028 5989
rect 6062 5955 6192 5989
rect -2630 5905 -2596 5921
rect -2630 5683 -2596 5729
rect -2710 5679 -2596 5683
rect -2534 5905 -2500 5921
rect -2534 5679 -2500 5729
rect -2420 5905 -2386 5921
rect -2420 5713 -2386 5729
rect -2324 5905 -2290 5921
rect -2324 5713 -2290 5729
rect -2210 5905 -2176 5921
rect -2210 5713 -2176 5729
rect -2114 5905 -2080 5921
rect -2114 5713 -2080 5729
rect -2000 5905 -1966 5921
rect -2000 5713 -1966 5729
rect -1904 5905 -1870 5921
rect -1904 5713 -1870 5729
rect -1790 5905 -1756 5921
rect -1790 5713 -1756 5729
rect -1694 5905 -1660 5921
rect -1694 5713 -1660 5729
rect -1580 5905 -1546 5921
rect -1580 5713 -1546 5729
rect -1484 5905 -1450 5921
rect -1484 5713 -1450 5729
rect -1370 5905 -1336 5921
rect -1370 5713 -1336 5729
rect -1274 5905 -1240 5921
rect -1274 5713 -1240 5729
rect -1160 5905 -1126 5921
rect -1160 5713 -1126 5729
rect -1064 5905 -1030 5921
rect -1064 5713 -1030 5729
rect -950 5905 -916 5921
rect -950 5713 -916 5729
rect -854 5905 -820 5921
rect -854 5713 -820 5729
rect -740 5905 -706 5921
rect -740 5713 -706 5729
rect -644 5905 -610 5921
rect -644 5713 -610 5729
rect -530 5905 -496 5921
rect -530 5713 -496 5729
rect -434 5905 -400 5921
rect -434 5713 -400 5729
rect -320 5905 -286 5921
rect -320 5713 -286 5729
rect -224 5905 -190 5921
rect -224 5713 -190 5729
rect -110 5905 -76 5921
rect -110 5713 -76 5729
rect -14 5905 20 5921
rect -14 5713 20 5729
rect 100 5905 134 5921
rect 100 5713 134 5729
rect 196 5905 230 5921
rect 196 5713 230 5729
rect 310 5905 344 5921
rect 310 5713 344 5729
rect 406 5905 440 5921
rect 406 5713 440 5729
rect 520 5905 554 5921
rect 520 5713 554 5729
rect 616 5905 650 5921
rect 616 5713 650 5729
rect 730 5905 764 5921
rect 730 5713 764 5729
rect 826 5905 860 5921
rect 826 5713 860 5729
rect 940 5905 974 5921
rect 940 5713 974 5729
rect 1036 5905 1070 5921
rect 1036 5713 1070 5729
rect 1150 5905 1184 5921
rect 1150 5713 1184 5729
rect 1246 5905 1280 5921
rect 1246 5713 1280 5729
rect 1360 5905 1394 5921
rect 1360 5713 1394 5729
rect 1456 5905 1490 5921
rect 1456 5713 1490 5729
rect 1570 5905 1604 5921
rect 1570 5713 1604 5729
rect 1666 5905 1700 5921
rect 1666 5713 1700 5729
rect 1780 5905 1814 5921
rect 1780 5713 1814 5729
rect 1876 5905 1910 5921
rect 1876 5713 1910 5729
rect 1990 5905 2024 5921
rect 1990 5713 2024 5729
rect 2086 5905 2120 5921
rect 2086 5713 2120 5729
rect 2200 5905 2234 5921
rect 2200 5713 2234 5729
rect 2296 5905 2330 5921
rect 2296 5713 2330 5729
rect 2410 5905 2444 5921
rect 2410 5713 2444 5729
rect 2506 5905 2540 5921
rect 2506 5713 2540 5729
rect 2620 5905 2654 5921
rect 2620 5713 2654 5729
rect 2716 5905 2750 5921
rect 2716 5713 2750 5729
rect 2830 5905 2864 5921
rect 2830 5713 2864 5729
rect 2926 5905 2960 5921
rect 2926 5713 2960 5729
rect 3040 5905 3074 5921
rect 3040 5713 3074 5729
rect 3136 5905 3170 5921
rect 3136 5713 3170 5729
rect 3250 5905 3284 5921
rect 3250 5713 3284 5729
rect 3346 5905 3380 5921
rect 3346 5713 3380 5729
rect 3460 5905 3494 5921
rect 3460 5713 3494 5729
rect 3556 5905 3590 5921
rect 3556 5713 3590 5729
rect 3670 5905 3704 5921
rect 3670 5713 3704 5729
rect 3766 5905 3800 5921
rect 3766 5713 3800 5729
rect 3880 5905 3914 5921
rect 3880 5713 3914 5729
rect 3976 5905 4010 5921
rect 3976 5713 4010 5729
rect 4090 5905 4124 5921
rect 4090 5713 4124 5729
rect 4186 5905 4220 5921
rect 4186 5713 4220 5729
rect 4300 5905 4334 5921
rect 4300 5713 4334 5729
rect 4396 5905 4430 5921
rect 4396 5713 4430 5729
rect 4510 5905 4544 5921
rect 4510 5713 4544 5729
rect 4606 5905 4640 5921
rect 4606 5713 4640 5729
rect 4720 5905 4754 5921
rect 4720 5713 4754 5729
rect 4816 5905 4850 5921
rect 4816 5713 4850 5729
rect 4930 5905 4964 5921
rect 4930 5713 4964 5729
rect 5026 5905 5060 5921
rect 5026 5713 5060 5729
rect 5140 5905 5174 5921
rect 5140 5713 5174 5729
rect 5236 5905 5270 5921
rect 5236 5713 5270 5729
rect 5350 5905 5384 5921
rect 5350 5713 5384 5729
rect 5446 5905 5480 5921
rect 5446 5713 5480 5729
rect 5560 5905 5594 5921
rect 5560 5713 5594 5729
rect 5656 5905 5690 5921
rect 5656 5713 5690 5729
rect 5770 5905 5804 5921
rect 5770 5713 5804 5729
rect 5866 5905 5900 5921
rect 5866 5713 5900 5729
rect 5980 5905 6014 5955
rect 5980 5713 6014 5729
rect 6076 5905 6110 5955
rect 6076 5713 6110 5729
rect -2710 5649 -2582 5679
rect -2630 5645 -2582 5649
rect -2548 5645 -2500 5679
rect -2178 5645 -2162 5679
rect -2128 5645 -2112 5679
rect -1758 5645 -1742 5679
rect -1708 5645 -1692 5679
rect -1338 5645 -1322 5679
rect -1288 5645 -1272 5679
rect -918 5645 -902 5679
rect -868 5645 -852 5679
rect -498 5645 -482 5679
rect -448 5645 -432 5679
rect -78 5645 -62 5679
rect -28 5645 -12 5679
rect 342 5645 358 5679
rect 392 5645 408 5679
rect 762 5645 778 5679
rect 812 5645 828 5679
rect 1182 5645 1198 5679
rect 1232 5645 1248 5679
rect 1602 5645 1618 5679
rect 1652 5645 1668 5679
rect 2022 5645 2038 5679
rect 2072 5645 2088 5679
rect 2442 5645 2458 5679
rect 2492 5645 2508 5679
rect 2862 5645 2878 5679
rect 2912 5645 2928 5679
rect 3282 5645 3298 5679
rect 3332 5645 3348 5679
rect 3702 5645 3718 5679
rect 3752 5645 3768 5679
rect 4122 5645 4138 5679
rect 4172 5645 4188 5679
rect 4542 5645 4558 5679
rect 4592 5645 4608 5679
rect 4962 5645 4978 5679
rect 5012 5645 5028 5679
rect 5382 5645 5398 5679
rect 5432 5645 5448 5679
rect 5802 5645 5818 5679
rect 5852 5645 5868 5679
rect -2388 5515 -2372 5549
rect -2338 5515 -2322 5549
rect -1968 5515 -1952 5549
rect -1918 5515 -1902 5549
rect -1548 5515 -1532 5549
rect -1498 5515 -1482 5549
rect -1128 5515 -1112 5549
rect -1078 5515 -1062 5549
rect -708 5515 -692 5549
rect -658 5515 -642 5549
rect -288 5515 -272 5549
rect -238 5515 -222 5549
rect 132 5515 148 5549
rect 182 5515 198 5549
rect 552 5515 568 5549
rect 602 5515 618 5549
rect 972 5515 988 5549
rect 1022 5515 1038 5549
rect 1392 5515 1408 5549
rect 1442 5515 1458 5549
rect 1812 5515 1828 5549
rect 1862 5515 1878 5549
rect 2232 5515 2248 5549
rect 2282 5515 2298 5549
rect 2652 5515 2668 5549
rect 2702 5515 2718 5549
rect 3072 5515 3088 5549
rect 3122 5515 3138 5549
rect 3492 5515 3508 5549
rect 3542 5515 3558 5549
rect 3912 5515 3928 5549
rect 3962 5515 3978 5549
rect 4332 5515 4348 5549
rect 4382 5515 4398 5549
rect 4752 5515 4768 5549
rect 4802 5515 4818 5549
rect 5172 5515 5188 5549
rect 5222 5515 5238 5549
rect 5592 5515 5608 5549
rect 5642 5515 5658 5549
rect 5980 5515 6028 5549
rect 6062 5515 6192 5549
rect -2630 5465 -2596 5481
rect -2630 5239 -2596 5289
rect -2534 5465 -2500 5481
rect -2534 5239 -2500 5289
rect -2420 5465 -2386 5481
rect -2420 5273 -2386 5289
rect -2324 5465 -2290 5481
rect -2324 5273 -2290 5289
rect -2210 5465 -2176 5481
rect -2210 5273 -2176 5289
rect -2114 5465 -2080 5481
rect -2114 5273 -2080 5289
rect -2000 5465 -1966 5481
rect -2000 5273 -1966 5289
rect -1904 5465 -1870 5481
rect -1904 5273 -1870 5289
rect -1790 5465 -1756 5481
rect -1790 5273 -1756 5289
rect -1694 5465 -1660 5481
rect -1694 5273 -1660 5289
rect -1580 5465 -1546 5481
rect -1580 5273 -1546 5289
rect -1484 5465 -1450 5481
rect -1484 5273 -1450 5289
rect -1370 5465 -1336 5481
rect -1370 5273 -1336 5289
rect -1274 5465 -1240 5481
rect -1274 5273 -1240 5289
rect -1160 5465 -1126 5481
rect -1160 5273 -1126 5289
rect -1064 5465 -1030 5481
rect -1064 5273 -1030 5289
rect -950 5465 -916 5481
rect -950 5273 -916 5289
rect -854 5465 -820 5481
rect -854 5273 -820 5289
rect -740 5465 -706 5481
rect -740 5273 -706 5289
rect -644 5465 -610 5481
rect -644 5273 -610 5289
rect -530 5465 -496 5481
rect -530 5273 -496 5289
rect -434 5465 -400 5481
rect -434 5273 -400 5289
rect -320 5465 -286 5481
rect -320 5273 -286 5289
rect -224 5465 -190 5481
rect -224 5273 -190 5289
rect -110 5465 -76 5481
rect -110 5273 -76 5289
rect -14 5465 20 5481
rect -14 5273 20 5289
rect 100 5465 134 5481
rect 100 5273 134 5289
rect 196 5465 230 5481
rect 196 5273 230 5289
rect 310 5465 344 5481
rect 310 5273 344 5289
rect 406 5465 440 5481
rect 406 5273 440 5289
rect 520 5465 554 5481
rect 520 5273 554 5289
rect 616 5465 650 5481
rect 616 5273 650 5289
rect 730 5465 764 5481
rect 730 5273 764 5289
rect 826 5465 860 5481
rect 826 5273 860 5289
rect 940 5465 974 5481
rect 940 5273 974 5289
rect 1036 5465 1070 5481
rect 1036 5273 1070 5289
rect 1150 5465 1184 5481
rect 1150 5273 1184 5289
rect 1246 5465 1280 5481
rect 1246 5273 1280 5289
rect 1360 5465 1394 5481
rect 1360 5273 1394 5289
rect 1456 5465 1490 5481
rect 1456 5273 1490 5289
rect 1570 5465 1604 5481
rect 1570 5273 1604 5289
rect 1666 5465 1700 5481
rect 1666 5273 1700 5289
rect 1780 5465 1814 5481
rect 1780 5273 1814 5289
rect 1876 5465 1910 5481
rect 1876 5273 1910 5289
rect 1990 5465 2024 5481
rect 1990 5273 2024 5289
rect 2086 5465 2120 5481
rect 2086 5273 2120 5289
rect 2200 5465 2234 5481
rect 2200 5273 2234 5289
rect 2296 5465 2330 5481
rect 2296 5273 2330 5289
rect 2410 5465 2444 5481
rect 2410 5273 2444 5289
rect 2506 5465 2540 5481
rect 2506 5273 2540 5289
rect 2620 5465 2654 5481
rect 2620 5273 2654 5289
rect 2716 5465 2750 5481
rect 2716 5273 2750 5289
rect 2830 5465 2864 5481
rect 2830 5273 2864 5289
rect 2926 5465 2960 5481
rect 2926 5273 2960 5289
rect 3040 5465 3074 5481
rect 3040 5273 3074 5289
rect 3136 5465 3170 5481
rect 3136 5273 3170 5289
rect 3250 5465 3284 5481
rect 3250 5273 3284 5289
rect 3346 5465 3380 5481
rect 3346 5273 3380 5289
rect 3460 5465 3494 5481
rect 3460 5273 3494 5289
rect 3556 5465 3590 5481
rect 3556 5273 3590 5289
rect 3670 5465 3704 5481
rect 3670 5273 3704 5289
rect 3766 5465 3800 5481
rect 3766 5273 3800 5289
rect 3880 5465 3914 5481
rect 3880 5273 3914 5289
rect 3976 5465 4010 5481
rect 3976 5273 4010 5289
rect 4090 5465 4124 5481
rect 4090 5273 4124 5289
rect 4186 5465 4220 5481
rect 4186 5273 4220 5289
rect 4300 5465 4334 5481
rect 4300 5273 4334 5289
rect 4396 5465 4430 5481
rect 4396 5273 4430 5289
rect 4510 5465 4544 5481
rect 4510 5273 4544 5289
rect 4606 5465 4640 5481
rect 4606 5273 4640 5289
rect 4720 5465 4754 5481
rect 4720 5273 4754 5289
rect 4816 5465 4850 5481
rect 4816 5273 4850 5289
rect 4930 5465 4964 5481
rect 4930 5273 4964 5289
rect 5026 5465 5060 5481
rect 5026 5273 5060 5289
rect 5140 5465 5174 5481
rect 5140 5273 5174 5289
rect 5236 5465 5270 5481
rect 5236 5273 5270 5289
rect 5350 5465 5384 5481
rect 5350 5273 5384 5289
rect 5446 5465 5480 5481
rect 5446 5273 5480 5289
rect 5560 5465 5594 5481
rect 5560 5273 5594 5289
rect 5656 5465 5690 5481
rect 5656 5273 5690 5289
rect 5770 5465 5804 5481
rect 5770 5273 5804 5289
rect 5866 5465 5900 5481
rect 5866 5273 5900 5289
rect 5980 5465 6014 5515
rect 5980 5273 6014 5289
rect 6076 5465 6110 5515
rect 6076 5273 6110 5289
rect -2710 5205 -2582 5239
rect -2548 5205 -2500 5239
rect -2178 5205 -2162 5239
rect -2128 5205 -2112 5239
rect -1758 5205 -1742 5239
rect -1708 5205 -1692 5239
rect -1338 5205 -1322 5239
rect -1288 5205 -1272 5239
rect -918 5205 -902 5239
rect -868 5205 -852 5239
rect -498 5205 -482 5239
rect -448 5205 -432 5239
rect -78 5205 -62 5239
rect -28 5205 -12 5239
rect 342 5205 358 5239
rect 392 5205 408 5239
rect 762 5205 778 5239
rect 812 5205 828 5239
rect 1182 5205 1198 5239
rect 1232 5205 1248 5239
rect 1602 5205 1618 5239
rect 1652 5205 1668 5239
rect 2022 5205 2038 5239
rect 2072 5205 2088 5239
rect 2442 5205 2458 5239
rect 2492 5205 2508 5239
rect 2862 5205 2878 5239
rect 2912 5205 2928 5239
rect 3282 5205 3298 5239
rect 3332 5205 3348 5239
rect 3702 5205 3718 5239
rect 3752 5205 3768 5239
rect 4122 5205 4138 5239
rect 4172 5205 4188 5239
rect 4542 5205 4558 5239
rect 4592 5205 4608 5239
rect 4962 5205 4978 5239
rect 5012 5205 5028 5239
rect 5382 5205 5398 5239
rect 5432 5205 5448 5239
rect 5802 5205 5818 5239
rect 5852 5205 5868 5239
rect -2388 5075 -2372 5109
rect -2338 5075 -2322 5109
rect -1968 5075 -1952 5109
rect -1918 5075 -1902 5109
rect -1548 5075 -1532 5109
rect -1498 5075 -1482 5109
rect -1128 5075 -1112 5109
rect -1078 5075 -1062 5109
rect -708 5075 -692 5109
rect -658 5075 -642 5109
rect -288 5075 -272 5109
rect -238 5075 -222 5109
rect 132 5075 148 5109
rect 182 5075 198 5109
rect 552 5075 568 5109
rect 602 5075 618 5109
rect 972 5075 988 5109
rect 1022 5075 1038 5109
rect 1392 5075 1408 5109
rect 1442 5075 1458 5109
rect 1812 5075 1828 5109
rect 1862 5075 1878 5109
rect 2232 5075 2248 5109
rect 2282 5075 2298 5109
rect 2652 5075 2668 5109
rect 2702 5075 2718 5109
rect 3072 5075 3088 5109
rect 3122 5075 3138 5109
rect 3492 5075 3508 5109
rect 3542 5075 3558 5109
rect 3912 5075 3928 5109
rect 3962 5075 3978 5109
rect 4332 5075 4348 5109
rect 4382 5075 4398 5109
rect 4752 5075 4768 5109
rect 4802 5075 4818 5109
rect 5172 5075 5188 5109
rect 5222 5075 5238 5109
rect 5592 5075 5608 5109
rect 5642 5075 5658 5109
rect 5980 5075 6028 5109
rect 6062 5075 6192 5109
rect -2630 5025 -2596 5041
rect -2630 4799 -2596 4849
rect -2534 5025 -2500 5041
rect -2534 4799 -2500 4849
rect -2420 5025 -2386 5041
rect -2420 4833 -2386 4849
rect -2324 5025 -2290 5041
rect -2324 4833 -2290 4849
rect -2210 5025 -2176 5041
rect -2210 4833 -2176 4849
rect -2114 5025 -2080 5041
rect -2114 4833 -2080 4849
rect -2000 5025 -1966 5041
rect -2000 4833 -1966 4849
rect -1904 5025 -1870 5041
rect -1904 4833 -1870 4849
rect -1790 5025 -1756 5041
rect -1790 4833 -1756 4849
rect -1694 5025 -1660 5041
rect -1694 4833 -1660 4849
rect -1580 5025 -1546 5041
rect -1580 4833 -1546 4849
rect -1484 5025 -1450 5041
rect -1484 4833 -1450 4849
rect -1370 5025 -1336 5041
rect -1370 4833 -1336 4849
rect -1274 5025 -1240 5041
rect -1274 4833 -1240 4849
rect -1160 5025 -1126 5041
rect -1160 4833 -1126 4849
rect -1064 5025 -1030 5041
rect -1064 4833 -1030 4849
rect -950 5025 -916 5041
rect -950 4833 -916 4849
rect -854 5025 -820 5041
rect -854 4833 -820 4849
rect -740 5025 -706 5041
rect -740 4833 -706 4849
rect -644 5025 -610 5041
rect -644 4833 -610 4849
rect -530 5025 -496 5041
rect -530 4833 -496 4849
rect -434 5025 -400 5041
rect -434 4833 -400 4849
rect -320 5025 -286 5041
rect -320 4833 -286 4849
rect -224 5025 -190 5041
rect -224 4833 -190 4849
rect -110 5025 -76 5041
rect -110 4833 -76 4849
rect -14 5025 20 5041
rect -14 4833 20 4849
rect 100 5025 134 5041
rect 100 4833 134 4849
rect 196 5025 230 5041
rect 196 4833 230 4849
rect 310 5025 344 5041
rect 310 4833 344 4849
rect 406 5025 440 5041
rect 406 4833 440 4849
rect 520 5025 554 5041
rect 520 4833 554 4849
rect 616 5025 650 5041
rect 616 4833 650 4849
rect 730 5025 764 5041
rect 730 4833 764 4849
rect 826 5025 860 5041
rect 826 4833 860 4849
rect 940 5025 974 5041
rect 940 4833 974 4849
rect 1036 5025 1070 5041
rect 1036 4833 1070 4849
rect 1150 5025 1184 5041
rect 1150 4833 1184 4849
rect 1246 5025 1280 5041
rect 1246 4833 1280 4849
rect 1360 5025 1394 5041
rect 1360 4833 1394 4849
rect 1456 5025 1490 5041
rect 1456 4833 1490 4849
rect 1570 5025 1604 5041
rect 1570 4833 1604 4849
rect 1666 5025 1700 5041
rect 1666 4833 1700 4849
rect 1780 5025 1814 5041
rect 1780 4833 1814 4849
rect 1876 5025 1910 5041
rect 1876 4833 1910 4849
rect 1990 5025 2024 5041
rect 1990 4833 2024 4849
rect 2086 5025 2120 5041
rect 2086 4833 2120 4849
rect 2200 5025 2234 5041
rect 2200 4833 2234 4849
rect 2296 5025 2330 5041
rect 2296 4833 2330 4849
rect 2410 5025 2444 5041
rect 2410 4833 2444 4849
rect 2506 5025 2540 5041
rect 2506 4833 2540 4849
rect 2620 5025 2654 5041
rect 2620 4833 2654 4849
rect 2716 5025 2750 5041
rect 2716 4833 2750 4849
rect 2830 5025 2864 5041
rect 2830 4833 2864 4849
rect 2926 5025 2960 5041
rect 2926 4833 2960 4849
rect 3040 5025 3074 5041
rect 3040 4833 3074 4849
rect 3136 5025 3170 5041
rect 3136 4833 3170 4849
rect 3250 5025 3284 5041
rect 3250 4833 3284 4849
rect 3346 5025 3380 5041
rect 3346 4833 3380 4849
rect 3460 5025 3494 5041
rect 3460 4833 3494 4849
rect 3556 5025 3590 5041
rect 3556 4833 3590 4849
rect 3670 5025 3704 5041
rect 3670 4833 3704 4849
rect 3766 5025 3800 5041
rect 3766 4833 3800 4849
rect 3880 5025 3914 5041
rect 3880 4833 3914 4849
rect 3976 5025 4010 5041
rect 3976 4833 4010 4849
rect 4090 5025 4124 5041
rect 4090 4833 4124 4849
rect 4186 5025 4220 5041
rect 4186 4833 4220 4849
rect 4300 5025 4334 5041
rect 4300 4833 4334 4849
rect 4396 5025 4430 5041
rect 4396 4833 4430 4849
rect 4510 5025 4544 5041
rect 4510 4833 4544 4849
rect 4606 5025 4640 5041
rect 4606 4833 4640 4849
rect 4720 5025 4754 5041
rect 4720 4833 4754 4849
rect 4816 5025 4850 5041
rect 4816 4833 4850 4849
rect 4930 5025 4964 5041
rect 4930 4833 4964 4849
rect 5026 5025 5060 5041
rect 5026 4833 5060 4849
rect 5140 5025 5174 5041
rect 5140 4833 5174 4849
rect 5236 5025 5270 5041
rect 5236 4833 5270 4849
rect 5350 5025 5384 5041
rect 5350 4833 5384 4849
rect 5446 5025 5480 5041
rect 5446 4833 5480 4849
rect 5560 5025 5594 5041
rect 5560 4833 5594 4849
rect 5656 5025 5690 5041
rect 5656 4833 5690 4849
rect 5770 5025 5804 5041
rect 5770 4833 5804 4849
rect 5866 5025 5900 5041
rect 5866 4833 5900 4849
rect 5980 5025 6014 5075
rect 5980 4833 6014 4849
rect 6076 5025 6110 5075
rect 6076 4833 6110 4849
rect -2710 4765 -2582 4799
rect -2548 4765 -2500 4799
rect -2178 4765 -2162 4799
rect -2128 4765 -2112 4799
rect -1758 4765 -1742 4799
rect -1708 4765 -1692 4799
rect -1338 4765 -1322 4799
rect -1288 4765 -1272 4799
rect -918 4765 -902 4799
rect -868 4765 -852 4799
rect -498 4765 -482 4799
rect -448 4765 -432 4799
rect -78 4765 -62 4799
rect -28 4765 -12 4799
rect 342 4765 358 4799
rect 392 4765 408 4799
rect 762 4765 778 4799
rect 812 4765 828 4799
rect 1182 4765 1198 4799
rect 1232 4765 1248 4799
rect 1602 4765 1618 4799
rect 1652 4765 1668 4799
rect 2022 4765 2038 4799
rect 2072 4765 2088 4799
rect 2442 4765 2458 4799
rect 2492 4765 2508 4799
rect 2862 4765 2878 4799
rect 2912 4765 2928 4799
rect 3282 4765 3298 4799
rect 3332 4765 3348 4799
rect 3702 4765 3718 4799
rect 3752 4765 3768 4799
rect 4122 4765 4138 4799
rect 4172 4765 4188 4799
rect 4542 4765 4558 4799
rect 4592 4765 4608 4799
rect 4962 4765 4978 4799
rect 5012 4765 5028 4799
rect 5382 4765 5398 4799
rect 5432 4765 5448 4799
rect 5802 4765 5818 4799
rect 5852 4765 5868 4799
rect -2744 4697 -2710 4759
rect 7180 7928 7214 7990
rect 6827 7876 6843 7910
rect 7019 7876 7180 7910
rect 7078 7862 7112 7876
rect 6750 7766 6784 7782
rect 6827 7780 6843 7814
rect 7019 7780 7035 7814
rect 7078 7812 7112 7828
rect 6750 7716 6784 7732
rect 6827 7684 6843 7718
rect 7019 7684 7035 7718
rect 7078 7670 7112 7686
rect 6750 7574 6784 7590
rect 6827 7588 6843 7622
rect 7019 7588 7035 7622
rect 7078 7620 7112 7636
rect 6750 7524 6784 7540
rect 6827 7492 6843 7526
rect 7019 7492 7035 7526
rect 7078 7478 7112 7494
rect 6750 7382 6784 7398
rect 6827 7396 6843 7430
rect 7019 7396 7035 7430
rect 7078 7428 7112 7444
rect 6750 7332 6784 7348
rect 6827 7300 6843 7334
rect 7019 7300 7035 7334
rect 7078 7286 7112 7302
rect 6750 7190 6784 7206
rect 6827 7204 6843 7238
rect 7019 7204 7035 7238
rect 7078 7236 7112 7252
rect 6750 7140 6784 7156
rect 6827 7108 6843 7142
rect 7019 7108 7035 7142
rect 7078 7094 7112 7110
rect 6750 6998 6784 7014
rect 6827 7012 6843 7046
rect 7019 7012 7035 7046
rect 7078 7044 7112 7060
rect 6750 6948 6784 6964
rect 6827 6916 6843 6950
rect 7019 6916 7035 6950
rect 7078 6902 7112 6918
rect 6750 6806 6784 6822
rect 6827 6820 6843 6854
rect 7019 6820 7035 6854
rect 7078 6852 7112 6868
rect 6750 6756 6784 6772
rect 6827 6724 6843 6758
rect 7019 6724 7035 6758
rect 7078 6710 7112 6726
rect 6750 6614 6784 6630
rect 6827 6628 6843 6662
rect 7019 6628 7035 6662
rect 7078 6660 7112 6676
rect 6750 6564 6784 6580
rect 6827 6532 6843 6566
rect 7019 6532 7035 6566
rect 7078 6518 7112 6534
rect 6750 6422 6784 6438
rect 6827 6436 6843 6470
rect 7019 6436 7035 6470
rect 7078 6468 7112 6484
rect 6750 6372 6784 6388
rect 6827 6340 6843 6374
rect 7019 6340 7035 6374
rect 7078 6326 7112 6342
rect 6750 6230 6784 6246
rect 6827 6244 6843 6278
rect 7019 6244 7035 6278
rect 7078 6276 7112 6292
rect 6750 6182 6784 6196
rect 6682 6148 6843 6182
rect 7019 6148 7035 6182
rect 6648 6068 6682 6130
rect 7180 6068 7214 6130
rect 6648 6034 6744 6068
rect 7118 6034 7214 6068
rect 6192 4697 6226 4759
rect -2744 4663 -2648 4697
rect 6130 4663 6226 4697
rect 6648 5580 6744 5614
rect 7118 5580 7214 5614
rect 6648 5518 6682 5580
rect -3218 3658 -3184 3720
rect -3750 3657 -3654 3658
rect -3750 3624 -3656 3657
rect -3280 3624 -3184 3658
rect -2744 4242 -2648 4276
rect 6130 4242 6226 4276
rect -2744 4180 -2710 4242
rect 6192 4180 6226 4242
rect -2388 4140 -2372 4174
rect -2338 4140 -2322 4174
rect -1968 4140 -1952 4174
rect -1918 4140 -1902 4174
rect -1548 4140 -1532 4174
rect -1498 4140 -1482 4174
rect -1128 4140 -1112 4174
rect -1078 4140 -1062 4174
rect -708 4140 -692 4174
rect -658 4140 -642 4174
rect -288 4140 -272 4174
rect -238 4140 -222 4174
rect 132 4140 148 4174
rect 182 4140 198 4174
rect 552 4140 568 4174
rect 602 4140 618 4174
rect 972 4140 988 4174
rect 1022 4140 1038 4174
rect 1392 4140 1408 4174
rect 1442 4140 1458 4174
rect 1812 4140 1828 4174
rect 1862 4140 1878 4174
rect 2232 4140 2248 4174
rect 2282 4140 2298 4174
rect 2652 4140 2668 4174
rect 2702 4140 2718 4174
rect 3072 4140 3088 4174
rect 3122 4140 3138 4174
rect 3492 4140 3508 4174
rect 3542 4140 3558 4174
rect 3912 4140 3928 4174
rect 3962 4140 3978 4174
rect 4332 4140 4348 4174
rect 4382 4140 4398 4174
rect 4752 4140 4768 4174
rect 4802 4140 4818 4174
rect 5172 4140 5188 4174
rect 5222 4140 5238 4174
rect 5592 4140 5608 4174
rect 5642 4140 5658 4174
rect 5980 4140 6028 4174
rect 6062 4140 6192 4174
rect -2630 4090 -2596 4106
rect -2630 3864 -2596 3914
rect -2534 4090 -2500 4106
rect -2534 3864 -2500 3914
rect -2420 4090 -2386 4106
rect -2420 3898 -2386 3914
rect -2324 4090 -2290 4106
rect -2324 3898 -2290 3914
rect -2210 4090 -2176 4106
rect -2210 3898 -2176 3914
rect -2114 4090 -2080 4106
rect -2114 3898 -2080 3914
rect -2000 4090 -1966 4106
rect -2000 3898 -1966 3914
rect -1904 4090 -1870 4106
rect -1904 3898 -1870 3914
rect -1790 4090 -1756 4106
rect -1790 3898 -1756 3914
rect -1694 4090 -1660 4106
rect -1694 3898 -1660 3914
rect -1580 4090 -1546 4106
rect -1580 3898 -1546 3914
rect -1484 4090 -1450 4106
rect -1484 3898 -1450 3914
rect -1370 4090 -1336 4106
rect -1370 3898 -1336 3914
rect -1274 4090 -1240 4106
rect -1274 3898 -1240 3914
rect -1160 4090 -1126 4106
rect -1160 3898 -1126 3914
rect -1064 4090 -1030 4106
rect -1064 3898 -1030 3914
rect -950 4090 -916 4106
rect -950 3898 -916 3914
rect -854 4090 -820 4106
rect -854 3898 -820 3914
rect -740 4090 -706 4106
rect -740 3898 -706 3914
rect -644 4090 -610 4106
rect -644 3898 -610 3914
rect -530 4090 -496 4106
rect -530 3898 -496 3914
rect -434 4090 -400 4106
rect -434 3898 -400 3914
rect -320 4090 -286 4106
rect -320 3898 -286 3914
rect -224 4090 -190 4106
rect -224 3898 -190 3914
rect -110 4090 -76 4106
rect -110 3898 -76 3914
rect -14 4090 20 4106
rect -14 3898 20 3914
rect 100 4090 134 4106
rect 100 3898 134 3914
rect 196 4090 230 4106
rect 196 3898 230 3914
rect 310 4090 344 4106
rect 310 3898 344 3914
rect 406 4090 440 4106
rect 406 3898 440 3914
rect 520 4090 554 4106
rect 520 3898 554 3914
rect 616 4090 650 4106
rect 616 3898 650 3914
rect 730 4090 764 4106
rect 730 3898 764 3914
rect 826 4090 860 4106
rect 826 3898 860 3914
rect 940 4090 974 4106
rect 940 3898 974 3914
rect 1036 4090 1070 4106
rect 1036 3898 1070 3914
rect 1150 4090 1184 4106
rect 1150 3898 1184 3914
rect 1246 4090 1280 4106
rect 1246 3898 1280 3914
rect 1360 4090 1394 4106
rect 1360 3898 1394 3914
rect 1456 4090 1490 4106
rect 1456 3898 1490 3914
rect 1570 4090 1604 4106
rect 1570 3898 1604 3914
rect 1666 4090 1700 4106
rect 1666 3898 1700 3914
rect 1780 4090 1814 4106
rect 1780 3898 1814 3914
rect 1876 4090 1910 4106
rect 1876 3898 1910 3914
rect 1990 4090 2024 4106
rect 1990 3898 2024 3914
rect 2086 4090 2120 4106
rect 2086 3898 2120 3914
rect 2200 4090 2234 4106
rect 2200 3898 2234 3914
rect 2296 4090 2330 4106
rect 2296 3898 2330 3914
rect 2410 4090 2444 4106
rect 2410 3898 2444 3914
rect 2506 4090 2540 4106
rect 2506 3898 2540 3914
rect 2620 4090 2654 4106
rect 2620 3898 2654 3914
rect 2716 4090 2750 4106
rect 2716 3898 2750 3914
rect 2830 4090 2864 4106
rect 2830 3898 2864 3914
rect 2926 4090 2960 4106
rect 2926 3898 2960 3914
rect 3040 4090 3074 4106
rect 3040 3898 3074 3914
rect 3136 4090 3170 4106
rect 3136 3898 3170 3914
rect 3250 4090 3284 4106
rect 3250 3898 3284 3914
rect 3346 4090 3380 4106
rect 3346 3898 3380 3914
rect 3460 4090 3494 4106
rect 3460 3898 3494 3914
rect 3556 4090 3590 4106
rect 3556 3898 3590 3914
rect 3670 4090 3704 4106
rect 3670 3898 3704 3914
rect 3766 4090 3800 4106
rect 3766 3898 3800 3914
rect 3880 4090 3914 4106
rect 3880 3898 3914 3914
rect 3976 4090 4010 4106
rect 3976 3898 4010 3914
rect 4090 4090 4124 4106
rect 4090 3898 4124 3914
rect 4186 4090 4220 4106
rect 4186 3898 4220 3914
rect 4300 4090 4334 4106
rect 4300 3898 4334 3914
rect 4396 4090 4430 4106
rect 4396 3898 4430 3914
rect 4510 4090 4544 4106
rect 4510 3898 4544 3914
rect 4606 4090 4640 4106
rect 4606 3898 4640 3914
rect 4720 4090 4754 4106
rect 4720 3898 4754 3914
rect 4816 4090 4850 4106
rect 4816 3898 4850 3914
rect 4930 4090 4964 4106
rect 4930 3898 4964 3914
rect 5026 4090 5060 4106
rect 5026 3898 5060 3914
rect 5140 4090 5174 4106
rect 5140 3898 5174 3914
rect 5236 4090 5270 4106
rect 5236 3898 5270 3914
rect 5350 4090 5384 4106
rect 5350 3898 5384 3914
rect 5446 4090 5480 4106
rect 5446 3898 5480 3914
rect 5560 4090 5594 4106
rect 5560 3898 5594 3914
rect 5656 4090 5690 4106
rect 5656 3898 5690 3914
rect 5770 4090 5804 4106
rect 5770 3898 5804 3914
rect 5866 4090 5900 4106
rect 5866 3898 5900 3914
rect 5980 4090 6014 4140
rect 5980 3898 6014 3914
rect 6076 4090 6110 4140
rect 6076 3898 6110 3914
rect -2710 3830 -2582 3864
rect -2548 3830 -2500 3864
rect -2178 3830 -2162 3864
rect -2128 3830 -2112 3864
rect -1758 3830 -1742 3864
rect -1708 3830 -1692 3864
rect -1338 3830 -1322 3864
rect -1288 3830 -1272 3864
rect -918 3830 -902 3864
rect -868 3830 -852 3864
rect -498 3830 -482 3864
rect -448 3830 -432 3864
rect -78 3830 -62 3864
rect -28 3830 -12 3864
rect 342 3830 358 3864
rect 392 3830 408 3864
rect 762 3830 778 3864
rect 812 3830 828 3864
rect 1182 3830 1198 3864
rect 1232 3830 1248 3864
rect 1602 3830 1618 3864
rect 1652 3830 1668 3864
rect 2022 3830 2038 3864
rect 2072 3830 2088 3864
rect 2442 3830 2458 3864
rect 2492 3830 2508 3864
rect 2862 3830 2878 3864
rect 2912 3830 2928 3864
rect 3282 3830 3298 3864
rect 3332 3830 3348 3864
rect 3702 3830 3718 3864
rect 3752 3830 3768 3864
rect 4122 3830 4138 3864
rect 4172 3830 4188 3864
rect 4542 3830 4558 3864
rect 4592 3830 4608 3864
rect 4962 3830 4978 3864
rect 5012 3830 5028 3864
rect 5382 3830 5398 3864
rect 5432 3830 5448 3864
rect 5802 3830 5818 3864
rect 5852 3830 5868 3864
rect -2388 3700 -2372 3734
rect -2338 3700 -2322 3734
rect -1968 3700 -1952 3734
rect -1918 3700 -1902 3734
rect -1548 3700 -1532 3734
rect -1498 3700 -1482 3734
rect -1128 3700 -1112 3734
rect -1078 3700 -1062 3734
rect -708 3700 -692 3734
rect -658 3700 -642 3734
rect -288 3700 -272 3734
rect -238 3700 -222 3734
rect 132 3700 148 3734
rect 182 3700 198 3734
rect 552 3700 568 3734
rect 602 3700 618 3734
rect 972 3700 988 3734
rect 1022 3700 1038 3734
rect 1392 3700 1408 3734
rect 1442 3700 1458 3734
rect 1812 3700 1828 3734
rect 1862 3700 1878 3734
rect 2232 3700 2248 3734
rect 2282 3700 2298 3734
rect 2652 3700 2668 3734
rect 2702 3700 2718 3734
rect 3072 3700 3088 3734
rect 3122 3700 3138 3734
rect 3492 3700 3508 3734
rect 3542 3700 3558 3734
rect 3912 3700 3928 3734
rect 3962 3700 3978 3734
rect 4332 3700 4348 3734
rect 4382 3700 4398 3734
rect 4752 3700 4768 3734
rect 4802 3700 4818 3734
rect 5172 3700 5188 3734
rect 5222 3700 5238 3734
rect 5592 3700 5608 3734
rect 5642 3700 5658 3734
rect 5980 3700 6028 3734
rect 6062 3700 6192 3734
rect -2630 3650 -2596 3666
rect -2630 3424 -2596 3474
rect -2534 3650 -2500 3666
rect -2534 3424 -2500 3474
rect -2420 3650 -2386 3666
rect -2420 3458 -2386 3474
rect -2324 3650 -2290 3666
rect -2324 3458 -2290 3474
rect -2210 3650 -2176 3666
rect -2210 3458 -2176 3474
rect -2114 3650 -2080 3666
rect -2114 3458 -2080 3474
rect -2000 3650 -1966 3666
rect -2000 3458 -1966 3474
rect -1904 3650 -1870 3666
rect -1904 3458 -1870 3474
rect -1790 3650 -1756 3666
rect -1790 3458 -1756 3474
rect -1694 3650 -1660 3666
rect -1694 3458 -1660 3474
rect -1580 3650 -1546 3666
rect -1580 3458 -1546 3474
rect -1484 3650 -1450 3666
rect -1484 3458 -1450 3474
rect -1370 3650 -1336 3666
rect -1370 3458 -1336 3474
rect -1274 3650 -1240 3666
rect -1274 3458 -1240 3474
rect -1160 3650 -1126 3666
rect -1160 3458 -1126 3474
rect -1064 3650 -1030 3666
rect -1064 3458 -1030 3474
rect -950 3650 -916 3666
rect -950 3458 -916 3474
rect -854 3650 -820 3666
rect -854 3458 -820 3474
rect -740 3650 -706 3666
rect -740 3458 -706 3474
rect -644 3650 -610 3666
rect -644 3458 -610 3474
rect -530 3650 -496 3666
rect -530 3458 -496 3474
rect -434 3650 -400 3666
rect -434 3458 -400 3474
rect -320 3650 -286 3666
rect -320 3458 -286 3474
rect -224 3650 -190 3666
rect -224 3458 -190 3474
rect -110 3650 -76 3666
rect -110 3458 -76 3474
rect -14 3650 20 3666
rect -14 3458 20 3474
rect 100 3650 134 3666
rect 100 3458 134 3474
rect 196 3650 230 3666
rect 196 3458 230 3474
rect 310 3650 344 3666
rect 310 3458 344 3474
rect 406 3650 440 3666
rect 406 3458 440 3474
rect 520 3650 554 3666
rect 520 3458 554 3474
rect 616 3650 650 3666
rect 616 3458 650 3474
rect 730 3650 764 3666
rect 730 3458 764 3474
rect 826 3650 860 3666
rect 826 3458 860 3474
rect 940 3650 974 3666
rect 940 3458 974 3474
rect 1036 3650 1070 3666
rect 1036 3458 1070 3474
rect 1150 3650 1184 3666
rect 1150 3458 1184 3474
rect 1246 3650 1280 3666
rect 1246 3458 1280 3474
rect 1360 3650 1394 3666
rect 1360 3458 1394 3474
rect 1456 3650 1490 3666
rect 1456 3458 1490 3474
rect 1570 3650 1604 3666
rect 1570 3458 1604 3474
rect 1666 3650 1700 3666
rect 1666 3458 1700 3474
rect 1780 3650 1814 3666
rect 1780 3458 1814 3474
rect 1876 3650 1910 3666
rect 1876 3458 1910 3474
rect 1990 3650 2024 3666
rect 1990 3458 2024 3474
rect 2086 3650 2120 3666
rect 2086 3458 2120 3474
rect 2200 3650 2234 3666
rect 2200 3458 2234 3474
rect 2296 3650 2330 3666
rect 2296 3458 2330 3474
rect 2410 3650 2444 3666
rect 2410 3458 2444 3474
rect 2506 3650 2540 3666
rect 2506 3458 2540 3474
rect 2620 3650 2654 3666
rect 2620 3458 2654 3474
rect 2716 3650 2750 3666
rect 2716 3458 2750 3474
rect 2830 3650 2864 3666
rect 2830 3458 2864 3474
rect 2926 3650 2960 3666
rect 2926 3458 2960 3474
rect 3040 3650 3074 3666
rect 3040 3458 3074 3474
rect 3136 3650 3170 3666
rect 3136 3458 3170 3474
rect 3250 3650 3284 3666
rect 3250 3458 3284 3474
rect 3346 3650 3380 3666
rect 3346 3458 3380 3474
rect 3460 3650 3494 3666
rect 3460 3458 3494 3474
rect 3556 3650 3590 3666
rect 3556 3458 3590 3474
rect 3670 3650 3704 3666
rect 3670 3458 3704 3474
rect 3766 3650 3800 3666
rect 3766 3458 3800 3474
rect 3880 3650 3914 3666
rect 3880 3458 3914 3474
rect 3976 3650 4010 3666
rect 3976 3458 4010 3474
rect 4090 3650 4124 3666
rect 4090 3458 4124 3474
rect 4186 3650 4220 3666
rect 4186 3458 4220 3474
rect 4300 3650 4334 3666
rect 4300 3458 4334 3474
rect 4396 3650 4430 3666
rect 4396 3458 4430 3474
rect 4510 3650 4544 3666
rect 4510 3458 4544 3474
rect 4606 3650 4640 3666
rect 4606 3458 4640 3474
rect 4720 3650 4754 3666
rect 4720 3458 4754 3474
rect 4816 3650 4850 3666
rect 4816 3458 4850 3474
rect 4930 3650 4964 3666
rect 4930 3458 4964 3474
rect 5026 3650 5060 3666
rect 5026 3458 5060 3474
rect 5140 3650 5174 3666
rect 5140 3458 5174 3474
rect 5236 3650 5270 3666
rect 5236 3458 5270 3474
rect 5350 3650 5384 3666
rect 5350 3458 5384 3474
rect 5446 3650 5480 3666
rect 5446 3458 5480 3474
rect 5560 3650 5594 3666
rect 5560 3458 5594 3474
rect 5656 3650 5690 3666
rect 5656 3458 5690 3474
rect 5770 3650 5804 3666
rect 5770 3458 5804 3474
rect 5866 3650 5900 3666
rect 5866 3458 5900 3474
rect 5980 3650 6014 3700
rect 5980 3458 6014 3474
rect 6076 3650 6110 3700
rect 6076 3458 6110 3474
rect -2710 3390 -2582 3424
rect -2548 3390 -2500 3424
rect -2178 3390 -2162 3424
rect -2128 3390 -2112 3424
rect -1758 3390 -1742 3424
rect -1708 3390 -1692 3424
rect -1338 3390 -1322 3424
rect -1288 3390 -1272 3424
rect -918 3390 -902 3424
rect -868 3390 -852 3424
rect -498 3390 -482 3424
rect -448 3390 -432 3424
rect -78 3390 -62 3424
rect -28 3390 -12 3424
rect 342 3390 358 3424
rect 392 3390 408 3424
rect 762 3390 778 3424
rect 812 3390 828 3424
rect 1182 3390 1198 3424
rect 1232 3390 1248 3424
rect 1602 3390 1618 3424
rect 1652 3390 1668 3424
rect 2022 3390 2038 3424
rect 2072 3390 2088 3424
rect 2442 3390 2458 3424
rect 2492 3390 2508 3424
rect 2862 3390 2878 3424
rect 2912 3390 2928 3424
rect 3282 3390 3298 3424
rect 3332 3390 3348 3424
rect 3702 3390 3718 3424
rect 3752 3390 3768 3424
rect 4122 3390 4138 3424
rect 4172 3390 4188 3424
rect 4542 3390 4558 3424
rect 4592 3390 4608 3424
rect 4962 3390 4978 3424
rect 5012 3390 5028 3424
rect 5382 3390 5398 3424
rect 5432 3390 5448 3424
rect 5802 3390 5818 3424
rect 5852 3390 5868 3424
rect -2388 3260 -2372 3294
rect -2338 3260 -2322 3294
rect -1968 3260 -1952 3294
rect -1918 3260 -1902 3294
rect -1548 3260 -1532 3294
rect -1498 3260 -1482 3294
rect -1128 3260 -1112 3294
rect -1078 3260 -1062 3294
rect -708 3260 -692 3294
rect -658 3260 -642 3294
rect -288 3260 -272 3294
rect -238 3260 -222 3294
rect 132 3260 148 3294
rect 182 3260 198 3294
rect 552 3260 568 3294
rect 602 3260 618 3294
rect 972 3260 988 3294
rect 1022 3260 1038 3294
rect 1392 3260 1408 3294
rect 1442 3260 1458 3294
rect 1812 3260 1828 3294
rect 1862 3260 1878 3294
rect 2232 3260 2248 3294
rect 2282 3260 2298 3294
rect 2652 3260 2668 3294
rect 2702 3260 2718 3294
rect 3072 3260 3088 3294
rect 3122 3260 3138 3294
rect 3492 3260 3508 3294
rect 3542 3260 3558 3294
rect 3912 3260 3928 3294
rect 3962 3260 3978 3294
rect 4332 3260 4348 3294
rect 4382 3260 4398 3294
rect 4752 3260 4768 3294
rect 4802 3260 4818 3294
rect 5172 3260 5188 3294
rect 5222 3260 5238 3294
rect 5592 3260 5608 3294
rect 5642 3260 5658 3294
rect 5980 3260 6028 3294
rect 6062 3260 6192 3294
rect -2630 3210 -2596 3226
rect -2630 2984 -2596 3034
rect -2534 3210 -2500 3226
rect -2534 2984 -2500 3034
rect -2420 3210 -2386 3226
rect -2420 3018 -2386 3034
rect -2324 3210 -2290 3226
rect -2324 3018 -2290 3034
rect -2210 3210 -2176 3226
rect -2210 3018 -2176 3034
rect -2114 3210 -2080 3226
rect -2114 3018 -2080 3034
rect -2000 3210 -1966 3226
rect -2000 3018 -1966 3034
rect -1904 3210 -1870 3226
rect -1904 3018 -1870 3034
rect -1790 3210 -1756 3226
rect -1790 3018 -1756 3034
rect -1694 3210 -1660 3226
rect -1694 3018 -1660 3034
rect -1580 3210 -1546 3226
rect -1580 3018 -1546 3034
rect -1484 3210 -1450 3226
rect -1484 3018 -1450 3034
rect -1370 3210 -1336 3226
rect -1370 3018 -1336 3034
rect -1274 3210 -1240 3226
rect -1274 3018 -1240 3034
rect -1160 3210 -1126 3226
rect -1160 3018 -1126 3034
rect -1064 3210 -1030 3226
rect -1064 3018 -1030 3034
rect -950 3210 -916 3226
rect -950 3018 -916 3034
rect -854 3210 -820 3226
rect -854 3018 -820 3034
rect -740 3210 -706 3226
rect -740 3018 -706 3034
rect -644 3210 -610 3226
rect -644 3018 -610 3034
rect -530 3210 -496 3226
rect -530 3018 -496 3034
rect -434 3210 -400 3226
rect -434 3018 -400 3034
rect -320 3210 -286 3226
rect -320 3018 -286 3034
rect -224 3210 -190 3226
rect -224 3018 -190 3034
rect -110 3210 -76 3226
rect -110 3018 -76 3034
rect -14 3210 20 3226
rect -14 3018 20 3034
rect 100 3210 134 3226
rect 100 3018 134 3034
rect 196 3210 230 3226
rect 196 3018 230 3034
rect 310 3210 344 3226
rect 310 3018 344 3034
rect 406 3210 440 3226
rect 406 3018 440 3034
rect 520 3210 554 3226
rect 520 3018 554 3034
rect 616 3210 650 3226
rect 616 3018 650 3034
rect 730 3210 764 3226
rect 730 3018 764 3034
rect 826 3210 860 3226
rect 826 3018 860 3034
rect 940 3210 974 3226
rect 940 3018 974 3034
rect 1036 3210 1070 3226
rect 1036 3018 1070 3034
rect 1150 3210 1184 3226
rect 1150 3018 1184 3034
rect 1246 3210 1280 3226
rect 1246 3018 1280 3034
rect 1360 3210 1394 3226
rect 1360 3018 1394 3034
rect 1456 3210 1490 3226
rect 1456 3018 1490 3034
rect 1570 3210 1604 3226
rect 1570 3018 1604 3034
rect 1666 3210 1700 3226
rect 1666 3018 1700 3034
rect 1780 3210 1814 3226
rect 1780 3018 1814 3034
rect 1876 3210 1910 3226
rect 1876 3018 1910 3034
rect 1990 3210 2024 3226
rect 1990 3018 2024 3034
rect 2086 3210 2120 3226
rect 2086 3018 2120 3034
rect 2200 3210 2234 3226
rect 2200 3018 2234 3034
rect 2296 3210 2330 3226
rect 2296 3018 2330 3034
rect 2410 3210 2444 3226
rect 2410 3018 2444 3034
rect 2506 3210 2540 3226
rect 2506 3018 2540 3034
rect 2620 3210 2654 3226
rect 2620 3018 2654 3034
rect 2716 3210 2750 3226
rect 2716 3018 2750 3034
rect 2830 3210 2864 3226
rect 2830 3018 2864 3034
rect 2926 3210 2960 3226
rect 2926 3018 2960 3034
rect 3040 3210 3074 3226
rect 3040 3018 3074 3034
rect 3136 3210 3170 3226
rect 3136 3018 3170 3034
rect 3250 3210 3284 3226
rect 3250 3018 3284 3034
rect 3346 3210 3380 3226
rect 3346 3018 3380 3034
rect 3460 3210 3494 3226
rect 3460 3018 3494 3034
rect 3556 3210 3590 3226
rect 3556 3018 3590 3034
rect 3670 3210 3704 3226
rect 3670 3018 3704 3034
rect 3766 3210 3800 3226
rect 3766 3018 3800 3034
rect 3880 3210 3914 3226
rect 3880 3018 3914 3034
rect 3976 3210 4010 3226
rect 3976 3018 4010 3034
rect 4090 3210 4124 3226
rect 4090 3018 4124 3034
rect 4186 3210 4220 3226
rect 4186 3018 4220 3034
rect 4300 3210 4334 3226
rect 4300 3018 4334 3034
rect 4396 3210 4430 3226
rect 4396 3018 4430 3034
rect 4510 3210 4544 3226
rect 4510 3018 4544 3034
rect 4606 3210 4640 3226
rect 4606 3018 4640 3034
rect 4720 3210 4754 3226
rect 4720 3018 4754 3034
rect 4816 3210 4850 3226
rect 4816 3018 4850 3034
rect 4930 3210 4964 3226
rect 4930 3018 4964 3034
rect 5026 3210 5060 3226
rect 5026 3018 5060 3034
rect 5140 3210 5174 3226
rect 5140 3018 5174 3034
rect 5236 3210 5270 3226
rect 5236 3018 5270 3034
rect 5350 3210 5384 3226
rect 5350 3018 5384 3034
rect 5446 3210 5480 3226
rect 5446 3018 5480 3034
rect 5560 3210 5594 3226
rect 5560 3018 5594 3034
rect 5656 3210 5690 3226
rect 5656 3018 5690 3034
rect 5770 3210 5804 3226
rect 5770 3018 5804 3034
rect 5866 3210 5900 3226
rect 5866 3018 5900 3034
rect 5980 3210 6014 3260
rect 5980 3018 6014 3034
rect 6076 3210 6110 3260
rect 6076 3018 6110 3034
rect -2710 2950 -2582 2984
rect -2548 2950 -2500 2984
rect -2178 2950 -2162 2984
rect -2128 2950 -2112 2984
rect -1758 2950 -1742 2984
rect -1708 2950 -1692 2984
rect -1338 2950 -1322 2984
rect -1288 2950 -1272 2984
rect -918 2950 -902 2984
rect -868 2950 -852 2984
rect -498 2950 -482 2984
rect -448 2950 -432 2984
rect -78 2950 -62 2984
rect -28 2950 -12 2984
rect 342 2950 358 2984
rect 392 2950 408 2984
rect 762 2950 778 2984
rect 812 2950 828 2984
rect 1182 2950 1198 2984
rect 1232 2950 1248 2984
rect 1602 2950 1618 2984
rect 1652 2950 1668 2984
rect 2022 2950 2038 2984
rect 2072 2950 2088 2984
rect 2442 2950 2458 2984
rect 2492 2950 2508 2984
rect 2862 2950 2878 2984
rect 2912 2950 2928 2984
rect 3282 2950 3298 2984
rect 3332 2950 3348 2984
rect 3702 2950 3718 2984
rect 3752 2950 3768 2984
rect 4122 2950 4138 2984
rect 4172 2950 4188 2984
rect 4542 2950 4558 2984
rect 4592 2950 4608 2984
rect 4962 2950 4978 2984
rect 5012 2950 5028 2984
rect 5382 2950 5398 2984
rect 5432 2950 5448 2984
rect 5802 2950 5818 2984
rect 5852 2950 5868 2984
rect -2388 2820 -2372 2854
rect -2338 2820 -2322 2854
rect -1968 2820 -1952 2854
rect -1918 2820 -1902 2854
rect -1548 2820 -1532 2854
rect -1498 2820 -1482 2854
rect -1128 2820 -1112 2854
rect -1078 2820 -1062 2854
rect -708 2820 -692 2854
rect -658 2820 -642 2854
rect -288 2820 -272 2854
rect -238 2820 -222 2854
rect 132 2820 148 2854
rect 182 2820 198 2854
rect 552 2820 568 2854
rect 602 2820 618 2854
rect 972 2820 988 2854
rect 1022 2820 1038 2854
rect 1392 2820 1408 2854
rect 1442 2820 1458 2854
rect 1812 2820 1828 2854
rect 1862 2820 1878 2854
rect 2232 2820 2248 2854
rect 2282 2820 2298 2854
rect 2652 2820 2668 2854
rect 2702 2820 2718 2854
rect 3072 2820 3088 2854
rect 3122 2820 3138 2854
rect 3492 2820 3508 2854
rect 3542 2820 3558 2854
rect 3912 2820 3928 2854
rect 3962 2820 3978 2854
rect 4332 2820 4348 2854
rect 4382 2820 4398 2854
rect 4752 2820 4768 2854
rect 4802 2820 4818 2854
rect 5172 2820 5188 2854
rect 5222 2820 5238 2854
rect 5592 2820 5608 2854
rect 5642 2820 5658 2854
rect 5980 2820 6028 2854
rect 6062 2820 6192 2854
rect -2630 2770 -2596 2786
rect -2630 2544 -2596 2594
rect -2534 2770 -2500 2786
rect -2534 2544 -2500 2594
rect -2420 2770 -2386 2786
rect -2420 2578 -2386 2594
rect -2324 2770 -2290 2786
rect -2324 2578 -2290 2594
rect -2210 2770 -2176 2786
rect -2210 2578 -2176 2594
rect -2114 2770 -2080 2786
rect -2114 2578 -2080 2594
rect -2000 2770 -1966 2786
rect -2000 2578 -1966 2594
rect -1904 2770 -1870 2786
rect -1904 2578 -1870 2594
rect -1790 2770 -1756 2786
rect -1790 2578 -1756 2594
rect -1694 2770 -1660 2786
rect -1694 2578 -1660 2594
rect -1580 2770 -1546 2786
rect -1580 2578 -1546 2594
rect -1484 2770 -1450 2786
rect -1484 2578 -1450 2594
rect -1370 2770 -1336 2786
rect -1370 2578 -1336 2594
rect -1274 2770 -1240 2786
rect -1274 2578 -1240 2594
rect -1160 2770 -1126 2786
rect -1160 2578 -1126 2594
rect -1064 2770 -1030 2786
rect -1064 2578 -1030 2594
rect -950 2770 -916 2786
rect -950 2578 -916 2594
rect -854 2770 -820 2786
rect -854 2578 -820 2594
rect -740 2770 -706 2786
rect -740 2578 -706 2594
rect -644 2770 -610 2786
rect -644 2578 -610 2594
rect -530 2770 -496 2786
rect -530 2578 -496 2594
rect -434 2770 -400 2786
rect -434 2578 -400 2594
rect -320 2770 -286 2786
rect -320 2578 -286 2594
rect -224 2770 -190 2786
rect -224 2578 -190 2594
rect -110 2770 -76 2786
rect -110 2578 -76 2594
rect -14 2770 20 2786
rect -14 2578 20 2594
rect 100 2770 134 2786
rect 100 2578 134 2594
rect 196 2770 230 2786
rect 196 2578 230 2594
rect 310 2770 344 2786
rect 310 2578 344 2594
rect 406 2770 440 2786
rect 406 2578 440 2594
rect 520 2770 554 2786
rect 520 2578 554 2594
rect 616 2770 650 2786
rect 616 2578 650 2594
rect 730 2770 764 2786
rect 730 2578 764 2594
rect 826 2770 860 2786
rect 826 2578 860 2594
rect 940 2770 974 2786
rect 940 2578 974 2594
rect 1036 2770 1070 2786
rect 1036 2578 1070 2594
rect 1150 2770 1184 2786
rect 1150 2578 1184 2594
rect 1246 2770 1280 2786
rect 1246 2578 1280 2594
rect 1360 2770 1394 2786
rect 1360 2578 1394 2594
rect 1456 2770 1490 2786
rect 1456 2578 1490 2594
rect 1570 2770 1604 2786
rect 1570 2578 1604 2594
rect 1666 2770 1700 2786
rect 1666 2578 1700 2594
rect 1780 2770 1814 2786
rect 1780 2578 1814 2594
rect 1876 2770 1910 2786
rect 1876 2578 1910 2594
rect 1990 2770 2024 2786
rect 1990 2578 2024 2594
rect 2086 2770 2120 2786
rect 2086 2578 2120 2594
rect 2200 2770 2234 2786
rect 2200 2578 2234 2594
rect 2296 2770 2330 2786
rect 2296 2578 2330 2594
rect 2410 2770 2444 2786
rect 2410 2578 2444 2594
rect 2506 2770 2540 2786
rect 2506 2578 2540 2594
rect 2620 2770 2654 2786
rect 2620 2578 2654 2594
rect 2716 2770 2750 2786
rect 2716 2578 2750 2594
rect 2830 2770 2864 2786
rect 2830 2578 2864 2594
rect 2926 2770 2960 2786
rect 2926 2578 2960 2594
rect 3040 2770 3074 2786
rect 3040 2578 3074 2594
rect 3136 2770 3170 2786
rect 3136 2578 3170 2594
rect 3250 2770 3284 2786
rect 3250 2578 3284 2594
rect 3346 2770 3380 2786
rect 3346 2578 3380 2594
rect 3460 2770 3494 2786
rect 3460 2578 3494 2594
rect 3556 2770 3590 2786
rect 3556 2578 3590 2594
rect 3670 2770 3704 2786
rect 3670 2578 3704 2594
rect 3766 2770 3800 2786
rect 3766 2578 3800 2594
rect 3880 2770 3914 2786
rect 3880 2578 3914 2594
rect 3976 2770 4010 2786
rect 3976 2578 4010 2594
rect 4090 2770 4124 2786
rect 4090 2578 4124 2594
rect 4186 2770 4220 2786
rect 4186 2578 4220 2594
rect 4300 2770 4334 2786
rect 4300 2578 4334 2594
rect 4396 2770 4430 2786
rect 4396 2578 4430 2594
rect 4510 2770 4544 2786
rect 4510 2578 4544 2594
rect 4606 2770 4640 2786
rect 4606 2578 4640 2594
rect 4720 2770 4754 2786
rect 4720 2578 4754 2594
rect 4816 2770 4850 2786
rect 4816 2578 4850 2594
rect 4930 2770 4964 2786
rect 4930 2578 4964 2594
rect 5026 2770 5060 2786
rect 5026 2578 5060 2594
rect 5140 2770 5174 2786
rect 5140 2578 5174 2594
rect 5236 2770 5270 2786
rect 5236 2578 5270 2594
rect 5350 2770 5384 2786
rect 5350 2578 5384 2594
rect 5446 2770 5480 2786
rect 5446 2578 5480 2594
rect 5560 2770 5594 2786
rect 5560 2578 5594 2594
rect 5656 2770 5690 2786
rect 5656 2578 5690 2594
rect 5770 2770 5804 2786
rect 5770 2578 5804 2594
rect 5866 2770 5900 2786
rect 5866 2578 5900 2594
rect 5980 2770 6014 2820
rect 5980 2578 6014 2594
rect 6076 2770 6110 2820
rect 6076 2578 6110 2594
rect -2710 2510 -2582 2544
rect -2548 2510 -2500 2544
rect -2178 2510 -2162 2544
rect -2128 2510 -2112 2544
rect -1758 2510 -1742 2544
rect -1708 2510 -1692 2544
rect -1338 2510 -1322 2544
rect -1288 2510 -1272 2544
rect -918 2510 -902 2544
rect -868 2510 -852 2544
rect -498 2510 -482 2544
rect -448 2510 -432 2544
rect -78 2510 -62 2544
rect -28 2510 -12 2544
rect 342 2510 358 2544
rect 392 2510 408 2544
rect 762 2510 778 2544
rect 812 2510 828 2544
rect 1182 2510 1198 2544
rect 1232 2510 1248 2544
rect 1602 2510 1618 2544
rect 1652 2510 1668 2544
rect 2022 2510 2038 2544
rect 2072 2510 2088 2544
rect 2442 2510 2458 2544
rect 2492 2510 2508 2544
rect 2862 2510 2878 2544
rect 2912 2510 2928 2544
rect 3282 2510 3298 2544
rect 3332 2510 3348 2544
rect 3702 2510 3718 2544
rect 3752 2510 3768 2544
rect 4122 2510 4138 2544
rect 4172 2510 4188 2544
rect 4542 2510 4558 2544
rect 4592 2510 4608 2544
rect 4962 2510 4978 2544
rect 5012 2510 5028 2544
rect 5382 2510 5398 2544
rect 5432 2510 5448 2544
rect 5802 2510 5818 2544
rect 5852 2510 5868 2544
rect -2388 2380 -2372 2414
rect -2338 2380 -2322 2414
rect -1968 2380 -1952 2414
rect -1918 2380 -1902 2414
rect -1548 2380 -1532 2414
rect -1498 2380 -1482 2414
rect -1128 2380 -1112 2414
rect -1078 2380 -1062 2414
rect -708 2380 -692 2414
rect -658 2380 -642 2414
rect -288 2380 -272 2414
rect -238 2380 -222 2414
rect 132 2380 148 2414
rect 182 2380 198 2414
rect 552 2380 568 2414
rect 602 2380 618 2414
rect 972 2380 988 2414
rect 1022 2380 1038 2414
rect 1392 2380 1408 2414
rect 1442 2380 1458 2414
rect 1812 2380 1828 2414
rect 1862 2380 1878 2414
rect 2232 2380 2248 2414
rect 2282 2380 2298 2414
rect 2652 2380 2668 2414
rect 2702 2380 2718 2414
rect 3072 2380 3088 2414
rect 3122 2380 3138 2414
rect 3492 2380 3508 2414
rect 3542 2380 3558 2414
rect 3912 2380 3928 2414
rect 3962 2380 3978 2414
rect 4332 2380 4348 2414
rect 4382 2380 4398 2414
rect 4752 2380 4768 2414
rect 4802 2380 4818 2414
rect 5172 2380 5188 2414
rect 5222 2380 5238 2414
rect 5592 2380 5608 2414
rect 5642 2380 5658 2414
rect 5980 2380 6028 2414
rect 6062 2380 6192 2414
rect -2630 2330 -2596 2346
rect -2630 2104 -2596 2154
rect -2534 2330 -2500 2346
rect -2534 2104 -2500 2154
rect -2420 2330 -2386 2346
rect -2420 2138 -2386 2154
rect -2324 2330 -2290 2346
rect -2324 2138 -2290 2154
rect -2210 2330 -2176 2346
rect -2210 2138 -2176 2154
rect -2114 2330 -2080 2346
rect -2114 2138 -2080 2154
rect -2000 2330 -1966 2346
rect -2000 2138 -1966 2154
rect -1904 2330 -1870 2346
rect -1904 2138 -1870 2154
rect -1790 2330 -1756 2346
rect -1790 2138 -1756 2154
rect -1694 2330 -1660 2346
rect -1694 2138 -1660 2154
rect -1580 2330 -1546 2346
rect -1580 2138 -1546 2154
rect -1484 2330 -1450 2346
rect -1484 2138 -1450 2154
rect -1370 2330 -1336 2346
rect -1370 2138 -1336 2154
rect -1274 2330 -1240 2346
rect -1274 2138 -1240 2154
rect -1160 2330 -1126 2346
rect -1160 2138 -1126 2154
rect -1064 2330 -1030 2346
rect -1064 2138 -1030 2154
rect -950 2330 -916 2346
rect -950 2138 -916 2154
rect -854 2330 -820 2346
rect -854 2138 -820 2154
rect -740 2330 -706 2346
rect -740 2138 -706 2154
rect -644 2330 -610 2346
rect -644 2138 -610 2154
rect -530 2330 -496 2346
rect -530 2138 -496 2154
rect -434 2330 -400 2346
rect -434 2138 -400 2154
rect -320 2330 -286 2346
rect -320 2138 -286 2154
rect -224 2330 -190 2346
rect -224 2138 -190 2154
rect -110 2330 -76 2346
rect -110 2138 -76 2154
rect -14 2330 20 2346
rect -14 2138 20 2154
rect 100 2330 134 2346
rect 100 2138 134 2154
rect 196 2330 230 2346
rect 196 2138 230 2154
rect 310 2330 344 2346
rect 310 2138 344 2154
rect 406 2330 440 2346
rect 406 2138 440 2154
rect 520 2330 554 2346
rect 520 2138 554 2154
rect 616 2330 650 2346
rect 616 2138 650 2154
rect 730 2330 764 2346
rect 730 2138 764 2154
rect 826 2330 860 2346
rect 826 2138 860 2154
rect 940 2330 974 2346
rect 940 2138 974 2154
rect 1036 2330 1070 2346
rect 1036 2138 1070 2154
rect 1150 2330 1184 2346
rect 1150 2138 1184 2154
rect 1246 2330 1280 2346
rect 1246 2138 1280 2154
rect 1360 2330 1394 2346
rect 1360 2138 1394 2154
rect 1456 2330 1490 2346
rect 1456 2138 1490 2154
rect 1570 2330 1604 2346
rect 1570 2138 1604 2154
rect 1666 2330 1700 2346
rect 1666 2138 1700 2154
rect 1780 2330 1814 2346
rect 1780 2138 1814 2154
rect 1876 2330 1910 2346
rect 1876 2138 1910 2154
rect 1990 2330 2024 2346
rect 1990 2138 2024 2154
rect 2086 2330 2120 2346
rect 2086 2138 2120 2154
rect 2200 2330 2234 2346
rect 2200 2138 2234 2154
rect 2296 2330 2330 2346
rect 2296 2138 2330 2154
rect 2410 2330 2444 2346
rect 2410 2138 2444 2154
rect 2506 2330 2540 2346
rect 2506 2138 2540 2154
rect 2620 2330 2654 2346
rect 2620 2138 2654 2154
rect 2716 2330 2750 2346
rect 2716 2138 2750 2154
rect 2830 2330 2864 2346
rect 2830 2138 2864 2154
rect 2926 2330 2960 2346
rect 2926 2138 2960 2154
rect 3040 2330 3074 2346
rect 3040 2138 3074 2154
rect 3136 2330 3170 2346
rect 3136 2138 3170 2154
rect 3250 2330 3284 2346
rect 3250 2138 3284 2154
rect 3346 2330 3380 2346
rect 3346 2138 3380 2154
rect 3460 2330 3494 2346
rect 3460 2138 3494 2154
rect 3556 2330 3590 2346
rect 3556 2138 3590 2154
rect 3670 2330 3704 2346
rect 3670 2138 3704 2154
rect 3766 2330 3800 2346
rect 3766 2138 3800 2154
rect 3880 2330 3914 2346
rect 3880 2138 3914 2154
rect 3976 2330 4010 2346
rect 3976 2138 4010 2154
rect 4090 2330 4124 2346
rect 4090 2138 4124 2154
rect 4186 2330 4220 2346
rect 4186 2138 4220 2154
rect 4300 2330 4334 2346
rect 4300 2138 4334 2154
rect 4396 2330 4430 2346
rect 4396 2138 4430 2154
rect 4510 2330 4544 2346
rect 4510 2138 4544 2154
rect 4606 2330 4640 2346
rect 4606 2138 4640 2154
rect 4720 2330 4754 2346
rect 4720 2138 4754 2154
rect 4816 2330 4850 2346
rect 4816 2138 4850 2154
rect 4930 2330 4964 2346
rect 4930 2138 4964 2154
rect 5026 2330 5060 2346
rect 5026 2138 5060 2154
rect 5140 2330 5174 2346
rect 5140 2138 5174 2154
rect 5236 2330 5270 2346
rect 5236 2138 5270 2154
rect 5350 2330 5384 2346
rect 5350 2138 5384 2154
rect 5446 2330 5480 2346
rect 5446 2138 5480 2154
rect 5560 2330 5594 2346
rect 5560 2138 5594 2154
rect 5656 2330 5690 2346
rect 5656 2138 5690 2154
rect 5770 2330 5804 2346
rect 5770 2138 5804 2154
rect 5866 2330 5900 2346
rect 5866 2138 5900 2154
rect 5980 2330 6014 2380
rect 5980 2138 6014 2154
rect 6076 2330 6110 2380
rect 6076 2138 6110 2154
rect -2710 2070 -2582 2104
rect -2548 2070 -2500 2104
rect -2178 2070 -2162 2104
rect -2128 2070 -2112 2104
rect -1758 2070 -1742 2104
rect -1708 2070 -1692 2104
rect -1338 2070 -1322 2104
rect -1288 2070 -1272 2104
rect -918 2070 -902 2104
rect -868 2070 -852 2104
rect -498 2070 -482 2104
rect -448 2070 -432 2104
rect -78 2070 -62 2104
rect -28 2070 -12 2104
rect 342 2070 358 2104
rect 392 2070 408 2104
rect 762 2070 778 2104
rect 812 2070 828 2104
rect 1182 2070 1198 2104
rect 1232 2070 1248 2104
rect 1602 2070 1618 2104
rect 1652 2070 1668 2104
rect 2022 2070 2038 2104
rect 2072 2070 2088 2104
rect 2442 2070 2458 2104
rect 2492 2070 2508 2104
rect 2862 2070 2878 2104
rect 2912 2070 2928 2104
rect 3282 2070 3298 2104
rect 3332 2070 3348 2104
rect 3702 2070 3718 2104
rect 3752 2070 3768 2104
rect 4122 2070 4138 2104
rect 4172 2070 4188 2104
rect 4542 2070 4558 2104
rect 4592 2070 4608 2104
rect 4962 2070 4978 2104
rect 5012 2070 5028 2104
rect 5382 2070 5398 2104
rect 5432 2070 5448 2104
rect 5802 2070 5818 2104
rect 5852 2070 5868 2104
rect -2388 1940 -2372 1974
rect -2338 1940 -2322 1974
rect -1968 1940 -1952 1974
rect -1918 1940 -1902 1974
rect -1548 1940 -1532 1974
rect -1498 1940 -1482 1974
rect -1128 1940 -1112 1974
rect -1078 1940 -1062 1974
rect -708 1940 -692 1974
rect -658 1940 -642 1974
rect -288 1940 -272 1974
rect -238 1940 -222 1974
rect 132 1940 148 1974
rect 182 1940 198 1974
rect 552 1940 568 1974
rect 602 1940 618 1974
rect 972 1940 988 1974
rect 1022 1940 1038 1974
rect 1392 1940 1408 1974
rect 1442 1940 1458 1974
rect 1812 1940 1828 1974
rect 1862 1940 1878 1974
rect 2232 1940 2248 1974
rect 2282 1940 2298 1974
rect 2652 1940 2668 1974
rect 2702 1940 2718 1974
rect 3072 1940 3088 1974
rect 3122 1940 3138 1974
rect 3492 1940 3508 1974
rect 3542 1940 3558 1974
rect 3912 1940 3928 1974
rect 3962 1940 3978 1974
rect 4332 1940 4348 1974
rect 4382 1940 4398 1974
rect 4752 1940 4768 1974
rect 4802 1940 4818 1974
rect 5172 1940 5188 1974
rect 5222 1940 5238 1974
rect 5592 1940 5608 1974
rect 5642 1940 5658 1974
rect 5980 1940 6028 1974
rect 6062 1940 6192 1974
rect -2630 1890 -2596 1906
rect -2630 1664 -2596 1714
rect -2534 1890 -2500 1906
rect -2534 1664 -2500 1714
rect -2420 1890 -2386 1906
rect -2420 1698 -2386 1714
rect -2324 1890 -2290 1906
rect -2324 1698 -2290 1714
rect -2210 1890 -2176 1906
rect -2210 1698 -2176 1714
rect -2114 1890 -2080 1906
rect -2114 1698 -2080 1714
rect -2000 1890 -1966 1906
rect -2000 1698 -1966 1714
rect -1904 1890 -1870 1906
rect -1904 1698 -1870 1714
rect -1790 1890 -1756 1906
rect -1790 1698 -1756 1714
rect -1694 1890 -1660 1906
rect -1694 1698 -1660 1714
rect -1580 1890 -1546 1906
rect -1580 1698 -1546 1714
rect -1484 1890 -1450 1906
rect -1484 1698 -1450 1714
rect -1370 1890 -1336 1906
rect -1370 1698 -1336 1714
rect -1274 1890 -1240 1906
rect -1274 1698 -1240 1714
rect -1160 1890 -1126 1906
rect -1160 1698 -1126 1714
rect -1064 1890 -1030 1906
rect -1064 1698 -1030 1714
rect -950 1890 -916 1906
rect -950 1698 -916 1714
rect -854 1890 -820 1906
rect -854 1698 -820 1714
rect -740 1890 -706 1906
rect -740 1698 -706 1714
rect -644 1890 -610 1906
rect -644 1698 -610 1714
rect -530 1890 -496 1906
rect -530 1698 -496 1714
rect -434 1890 -400 1906
rect -434 1698 -400 1714
rect -320 1890 -286 1906
rect -320 1698 -286 1714
rect -224 1890 -190 1906
rect -224 1698 -190 1714
rect -110 1890 -76 1906
rect -110 1698 -76 1714
rect -14 1890 20 1906
rect -14 1698 20 1714
rect 100 1890 134 1906
rect 100 1698 134 1714
rect 196 1890 230 1906
rect 196 1698 230 1714
rect 310 1890 344 1906
rect 310 1698 344 1714
rect 406 1890 440 1906
rect 406 1698 440 1714
rect 520 1890 554 1906
rect 520 1698 554 1714
rect 616 1890 650 1906
rect 616 1698 650 1714
rect 730 1890 764 1906
rect 730 1698 764 1714
rect 826 1890 860 1906
rect 826 1698 860 1714
rect 940 1890 974 1906
rect 940 1698 974 1714
rect 1036 1890 1070 1906
rect 1036 1698 1070 1714
rect 1150 1890 1184 1906
rect 1150 1698 1184 1714
rect 1246 1890 1280 1906
rect 1246 1698 1280 1714
rect 1360 1890 1394 1906
rect 1360 1698 1394 1714
rect 1456 1890 1490 1906
rect 1456 1698 1490 1714
rect 1570 1890 1604 1906
rect 1570 1698 1604 1714
rect 1666 1890 1700 1906
rect 1666 1698 1700 1714
rect 1780 1890 1814 1906
rect 1780 1698 1814 1714
rect 1876 1890 1910 1906
rect 1876 1698 1910 1714
rect 1990 1890 2024 1906
rect 1990 1698 2024 1714
rect 2086 1890 2120 1906
rect 2086 1698 2120 1714
rect 2200 1890 2234 1906
rect 2200 1698 2234 1714
rect 2296 1890 2330 1906
rect 2296 1698 2330 1714
rect 2410 1890 2444 1906
rect 2410 1698 2444 1714
rect 2506 1890 2540 1906
rect 2506 1698 2540 1714
rect 2620 1890 2654 1906
rect 2620 1698 2654 1714
rect 2716 1890 2750 1906
rect 2716 1698 2750 1714
rect 2830 1890 2864 1906
rect 2830 1698 2864 1714
rect 2926 1890 2960 1906
rect 2926 1698 2960 1714
rect 3040 1890 3074 1906
rect 3040 1698 3074 1714
rect 3136 1890 3170 1906
rect 3136 1698 3170 1714
rect 3250 1890 3284 1906
rect 3250 1698 3284 1714
rect 3346 1890 3380 1906
rect 3346 1698 3380 1714
rect 3460 1890 3494 1906
rect 3460 1698 3494 1714
rect 3556 1890 3590 1906
rect 3556 1698 3590 1714
rect 3670 1890 3704 1906
rect 3670 1698 3704 1714
rect 3766 1890 3800 1906
rect 3766 1698 3800 1714
rect 3880 1890 3914 1906
rect 3880 1698 3914 1714
rect 3976 1890 4010 1906
rect 3976 1698 4010 1714
rect 4090 1890 4124 1906
rect 4090 1698 4124 1714
rect 4186 1890 4220 1906
rect 4186 1698 4220 1714
rect 4300 1890 4334 1906
rect 4300 1698 4334 1714
rect 4396 1890 4430 1906
rect 4396 1698 4430 1714
rect 4510 1890 4544 1906
rect 4510 1698 4544 1714
rect 4606 1890 4640 1906
rect 4606 1698 4640 1714
rect 4720 1890 4754 1906
rect 4720 1698 4754 1714
rect 4816 1890 4850 1906
rect 4816 1698 4850 1714
rect 4930 1890 4964 1906
rect 4930 1698 4964 1714
rect 5026 1890 5060 1906
rect 5026 1698 5060 1714
rect 5140 1890 5174 1906
rect 5140 1698 5174 1714
rect 5236 1890 5270 1906
rect 5236 1698 5270 1714
rect 5350 1890 5384 1906
rect 5350 1698 5384 1714
rect 5446 1890 5480 1906
rect 5446 1698 5480 1714
rect 5560 1890 5594 1906
rect 5560 1698 5594 1714
rect 5656 1890 5690 1906
rect 5656 1698 5690 1714
rect 5770 1890 5804 1906
rect 5770 1698 5804 1714
rect 5866 1890 5900 1906
rect 5866 1698 5900 1714
rect 5980 1890 6014 1940
rect 5980 1698 6014 1714
rect 6076 1890 6110 1940
rect 6076 1698 6110 1714
rect -2710 1630 -2582 1664
rect -2548 1630 -2500 1664
rect -2178 1630 -2162 1664
rect -2128 1630 -2112 1664
rect -1758 1630 -1742 1664
rect -1708 1630 -1692 1664
rect -1338 1630 -1322 1664
rect -1288 1630 -1272 1664
rect -918 1630 -902 1664
rect -868 1630 -852 1664
rect -498 1630 -482 1664
rect -448 1630 -432 1664
rect -78 1630 -62 1664
rect -28 1630 -12 1664
rect 342 1630 358 1664
rect 392 1630 408 1664
rect 762 1630 778 1664
rect 812 1630 828 1664
rect 1182 1630 1198 1664
rect 1232 1630 1248 1664
rect 1602 1630 1618 1664
rect 1652 1630 1668 1664
rect 2022 1630 2038 1664
rect 2072 1630 2088 1664
rect 2442 1630 2458 1664
rect 2492 1630 2508 1664
rect 2862 1630 2878 1664
rect 2912 1630 2928 1664
rect 3282 1630 3298 1664
rect 3332 1630 3348 1664
rect 3702 1630 3718 1664
rect 3752 1630 3768 1664
rect 4122 1630 4138 1664
rect 4172 1630 4188 1664
rect 4542 1630 4558 1664
rect 4592 1630 4608 1664
rect 4962 1630 4978 1664
rect 5012 1630 5028 1664
rect 5382 1630 5398 1664
rect 5432 1630 5448 1664
rect 5802 1630 5818 1664
rect 5852 1630 5868 1664
rect -2388 1500 -2372 1534
rect -2338 1500 -2322 1534
rect -1968 1500 -1952 1534
rect -1918 1500 -1902 1534
rect -1548 1500 -1532 1534
rect -1498 1500 -1482 1534
rect -1128 1500 -1112 1534
rect -1078 1500 -1062 1534
rect -708 1500 -692 1534
rect -658 1500 -642 1534
rect -288 1500 -272 1534
rect -238 1500 -222 1534
rect 132 1500 148 1534
rect 182 1500 198 1534
rect 552 1500 568 1534
rect 602 1500 618 1534
rect 972 1500 988 1534
rect 1022 1500 1038 1534
rect 1392 1500 1408 1534
rect 1442 1500 1458 1534
rect 1812 1500 1828 1534
rect 1862 1500 1878 1534
rect 2232 1500 2248 1534
rect 2282 1500 2298 1534
rect 2652 1500 2668 1534
rect 2702 1500 2718 1534
rect 3072 1500 3088 1534
rect 3122 1500 3138 1534
rect 3492 1500 3508 1534
rect 3542 1500 3558 1534
rect 3912 1500 3928 1534
rect 3962 1500 3978 1534
rect 4332 1500 4348 1534
rect 4382 1500 4398 1534
rect 4752 1500 4768 1534
rect 4802 1500 4818 1534
rect 5172 1500 5188 1534
rect 5222 1500 5238 1534
rect 5592 1500 5608 1534
rect 5642 1500 5658 1534
rect 5980 1500 6028 1534
rect 6062 1500 6192 1534
rect -2630 1450 -2596 1466
rect -2630 1224 -2596 1274
rect -2534 1450 -2500 1466
rect -2534 1224 -2500 1274
rect -2420 1450 -2386 1466
rect -2420 1258 -2386 1274
rect -2324 1450 -2290 1466
rect -2324 1258 -2290 1274
rect -2210 1450 -2176 1466
rect -2210 1258 -2176 1274
rect -2114 1450 -2080 1466
rect -2114 1258 -2080 1274
rect -2000 1450 -1966 1466
rect -2000 1258 -1966 1274
rect -1904 1450 -1870 1466
rect -1904 1258 -1870 1274
rect -1790 1450 -1756 1466
rect -1790 1258 -1756 1274
rect -1694 1450 -1660 1466
rect -1694 1258 -1660 1274
rect -1580 1450 -1546 1466
rect -1580 1258 -1546 1274
rect -1484 1450 -1450 1466
rect -1484 1258 -1450 1274
rect -1370 1450 -1336 1466
rect -1370 1258 -1336 1274
rect -1274 1450 -1240 1466
rect -1274 1258 -1240 1274
rect -1160 1450 -1126 1466
rect -1160 1258 -1126 1274
rect -1064 1450 -1030 1466
rect -1064 1258 -1030 1274
rect -950 1450 -916 1466
rect -950 1258 -916 1274
rect -854 1450 -820 1466
rect -854 1258 -820 1274
rect -740 1450 -706 1466
rect -740 1258 -706 1274
rect -644 1450 -610 1466
rect -644 1258 -610 1274
rect -530 1450 -496 1466
rect -530 1258 -496 1274
rect -434 1450 -400 1466
rect -434 1258 -400 1274
rect -320 1450 -286 1466
rect -320 1258 -286 1274
rect -224 1450 -190 1466
rect -224 1258 -190 1274
rect -110 1450 -76 1466
rect -110 1258 -76 1274
rect -14 1450 20 1466
rect -14 1258 20 1274
rect 100 1450 134 1466
rect 100 1258 134 1274
rect 196 1450 230 1466
rect 196 1258 230 1274
rect 310 1450 344 1466
rect 310 1258 344 1274
rect 406 1450 440 1466
rect 406 1258 440 1274
rect 520 1450 554 1466
rect 520 1258 554 1274
rect 616 1450 650 1466
rect 616 1258 650 1274
rect 730 1450 764 1466
rect 730 1258 764 1274
rect 826 1450 860 1466
rect 826 1258 860 1274
rect 940 1450 974 1466
rect 940 1258 974 1274
rect 1036 1450 1070 1466
rect 1036 1258 1070 1274
rect 1150 1450 1184 1466
rect 1150 1258 1184 1274
rect 1246 1450 1280 1466
rect 1246 1258 1280 1274
rect 1360 1450 1394 1466
rect 1360 1258 1394 1274
rect 1456 1450 1490 1466
rect 1456 1258 1490 1274
rect 1570 1450 1604 1466
rect 1570 1258 1604 1274
rect 1666 1450 1700 1466
rect 1666 1258 1700 1274
rect 1780 1450 1814 1466
rect 1780 1258 1814 1274
rect 1876 1450 1910 1466
rect 1876 1258 1910 1274
rect 1990 1450 2024 1466
rect 1990 1258 2024 1274
rect 2086 1450 2120 1466
rect 2086 1258 2120 1274
rect 2200 1450 2234 1466
rect 2200 1258 2234 1274
rect 2296 1450 2330 1466
rect 2296 1258 2330 1274
rect 2410 1450 2444 1466
rect 2410 1258 2444 1274
rect 2506 1450 2540 1466
rect 2506 1258 2540 1274
rect 2620 1450 2654 1466
rect 2620 1258 2654 1274
rect 2716 1450 2750 1466
rect 2716 1258 2750 1274
rect 2830 1450 2864 1466
rect 2830 1258 2864 1274
rect 2926 1450 2960 1466
rect 2926 1258 2960 1274
rect 3040 1450 3074 1466
rect 3040 1258 3074 1274
rect 3136 1450 3170 1466
rect 3136 1258 3170 1274
rect 3250 1450 3284 1466
rect 3250 1258 3284 1274
rect 3346 1450 3380 1466
rect 3346 1258 3380 1274
rect 3460 1450 3494 1466
rect 3460 1258 3494 1274
rect 3556 1450 3590 1466
rect 3556 1258 3590 1274
rect 3670 1450 3704 1466
rect 3670 1258 3704 1274
rect 3766 1450 3800 1466
rect 3766 1258 3800 1274
rect 3880 1450 3914 1466
rect 3880 1258 3914 1274
rect 3976 1450 4010 1466
rect 3976 1258 4010 1274
rect 4090 1450 4124 1466
rect 4090 1258 4124 1274
rect 4186 1450 4220 1466
rect 4186 1258 4220 1274
rect 4300 1450 4334 1466
rect 4300 1258 4334 1274
rect 4396 1450 4430 1466
rect 4396 1258 4430 1274
rect 4510 1450 4544 1466
rect 4510 1258 4544 1274
rect 4606 1450 4640 1466
rect 4606 1258 4640 1274
rect 4720 1450 4754 1466
rect 4720 1258 4754 1274
rect 4816 1450 4850 1466
rect 4816 1258 4850 1274
rect 4930 1450 4964 1466
rect 4930 1258 4964 1274
rect 5026 1450 5060 1466
rect 5026 1258 5060 1274
rect 5140 1450 5174 1466
rect 5140 1258 5174 1274
rect 5236 1450 5270 1466
rect 5236 1258 5270 1274
rect 5350 1450 5384 1466
rect 5350 1258 5384 1274
rect 5446 1450 5480 1466
rect 5446 1258 5480 1274
rect 5560 1450 5594 1466
rect 5560 1258 5594 1274
rect 5656 1450 5690 1466
rect 5656 1258 5690 1274
rect 5770 1450 5804 1466
rect 5770 1258 5804 1274
rect 5866 1450 5900 1466
rect 5866 1258 5900 1274
rect 5980 1450 6014 1500
rect 5980 1258 6014 1274
rect 6076 1450 6110 1500
rect 6076 1258 6110 1274
rect -2710 1190 -2582 1224
rect -2548 1190 -2500 1224
rect -2178 1190 -2162 1224
rect -2128 1190 -2112 1224
rect -1758 1190 -1742 1224
rect -1708 1190 -1692 1224
rect -1338 1190 -1322 1224
rect -1288 1190 -1272 1224
rect -918 1190 -902 1224
rect -868 1190 -852 1224
rect -498 1190 -482 1224
rect -448 1190 -432 1224
rect -78 1190 -62 1224
rect -28 1190 -12 1224
rect 342 1190 358 1224
rect 392 1190 408 1224
rect 762 1190 778 1224
rect 812 1190 828 1224
rect 1182 1190 1198 1224
rect 1232 1190 1248 1224
rect 1602 1190 1618 1224
rect 1652 1190 1668 1224
rect 2022 1190 2038 1224
rect 2072 1190 2088 1224
rect 2442 1190 2458 1224
rect 2492 1190 2508 1224
rect 2862 1190 2878 1224
rect 2912 1190 2928 1224
rect 3282 1190 3298 1224
rect 3332 1190 3348 1224
rect 3702 1190 3718 1224
rect 3752 1190 3768 1224
rect 4122 1190 4138 1224
rect 4172 1190 4188 1224
rect 4542 1190 4558 1224
rect 4592 1190 4608 1224
rect 4962 1190 4978 1224
rect 5012 1190 5028 1224
rect 5382 1190 5398 1224
rect 5432 1190 5448 1224
rect 5802 1190 5818 1224
rect 5852 1190 5868 1224
rect -2388 1060 -2372 1094
rect -2338 1060 -2322 1094
rect -1968 1060 -1952 1094
rect -1918 1060 -1902 1094
rect -1548 1060 -1532 1094
rect -1498 1060 -1482 1094
rect -1128 1060 -1112 1094
rect -1078 1060 -1062 1094
rect -708 1060 -692 1094
rect -658 1060 -642 1094
rect -288 1060 -272 1094
rect -238 1060 -222 1094
rect 132 1060 148 1094
rect 182 1060 198 1094
rect 552 1060 568 1094
rect 602 1060 618 1094
rect 972 1060 988 1094
rect 1022 1060 1038 1094
rect 1392 1060 1408 1094
rect 1442 1060 1458 1094
rect 1812 1060 1828 1094
rect 1862 1060 1878 1094
rect 2232 1060 2248 1094
rect 2282 1060 2298 1094
rect 2652 1060 2668 1094
rect 2702 1060 2718 1094
rect 3072 1060 3088 1094
rect 3122 1060 3138 1094
rect 3492 1060 3508 1094
rect 3542 1060 3558 1094
rect 3912 1060 3928 1094
rect 3962 1060 3978 1094
rect 4332 1060 4348 1094
rect 4382 1060 4398 1094
rect 4752 1060 4768 1094
rect 4802 1060 4818 1094
rect 5172 1060 5188 1094
rect 5222 1060 5238 1094
rect 5592 1060 5608 1094
rect 5642 1060 5658 1094
rect 5980 1060 6028 1094
rect 6062 1093 6110 1094
rect 6062 1060 6192 1093
rect -2630 1010 -2596 1026
rect -2630 784 -2596 834
rect -2534 1010 -2500 1026
rect -2534 784 -2500 834
rect -2420 1010 -2386 1026
rect -2420 818 -2386 834
rect -2324 1010 -2290 1026
rect -2324 818 -2290 834
rect -2210 1010 -2176 1026
rect -2210 818 -2176 834
rect -2114 1010 -2080 1026
rect -2114 818 -2080 834
rect -2000 1010 -1966 1026
rect -2000 818 -1966 834
rect -1904 1010 -1870 1026
rect -1904 818 -1870 834
rect -1790 1010 -1756 1026
rect -1790 818 -1756 834
rect -1694 1010 -1660 1026
rect -1694 818 -1660 834
rect -1580 1010 -1546 1026
rect -1580 818 -1546 834
rect -1484 1010 -1450 1026
rect -1484 818 -1450 834
rect -1370 1010 -1336 1026
rect -1370 818 -1336 834
rect -1274 1010 -1240 1026
rect -1274 818 -1240 834
rect -1160 1010 -1126 1026
rect -1160 818 -1126 834
rect -1064 1010 -1030 1026
rect -1064 818 -1030 834
rect -950 1010 -916 1026
rect -950 818 -916 834
rect -854 1010 -820 1026
rect -854 818 -820 834
rect -740 1010 -706 1026
rect -740 818 -706 834
rect -644 1010 -610 1026
rect -644 818 -610 834
rect -530 1010 -496 1026
rect -530 818 -496 834
rect -434 1010 -400 1026
rect -434 818 -400 834
rect -320 1010 -286 1026
rect -320 818 -286 834
rect -224 1010 -190 1026
rect -224 818 -190 834
rect -110 1010 -76 1026
rect -110 818 -76 834
rect -14 1010 20 1026
rect -14 818 20 834
rect 100 1010 134 1026
rect 100 818 134 834
rect 196 1010 230 1026
rect 196 818 230 834
rect 310 1010 344 1026
rect 310 818 344 834
rect 406 1010 440 1026
rect 406 818 440 834
rect 520 1010 554 1026
rect 520 818 554 834
rect 616 1010 650 1026
rect 616 818 650 834
rect 730 1010 764 1026
rect 730 818 764 834
rect 826 1010 860 1026
rect 826 818 860 834
rect 940 1010 974 1026
rect 940 818 974 834
rect 1036 1010 1070 1026
rect 1036 818 1070 834
rect 1150 1010 1184 1026
rect 1150 818 1184 834
rect 1246 1010 1280 1026
rect 1246 818 1280 834
rect 1360 1010 1394 1026
rect 1360 818 1394 834
rect 1456 1010 1490 1026
rect 1456 818 1490 834
rect 1570 1010 1604 1026
rect 1570 818 1604 834
rect 1666 1010 1700 1026
rect 1666 818 1700 834
rect 1780 1010 1814 1026
rect 1780 818 1814 834
rect 1876 1010 1910 1026
rect 1876 818 1910 834
rect 1990 1010 2024 1026
rect 1990 818 2024 834
rect 2086 1010 2120 1026
rect 2086 818 2120 834
rect 2200 1010 2234 1026
rect 2200 818 2234 834
rect 2296 1010 2330 1026
rect 2296 818 2330 834
rect 2410 1010 2444 1026
rect 2410 818 2444 834
rect 2506 1010 2540 1026
rect 2506 818 2540 834
rect 2620 1010 2654 1026
rect 2620 818 2654 834
rect 2716 1010 2750 1026
rect 2716 818 2750 834
rect 2830 1010 2864 1026
rect 2830 818 2864 834
rect 2926 1010 2960 1026
rect 2926 818 2960 834
rect 3040 1010 3074 1026
rect 3040 818 3074 834
rect 3136 1010 3170 1026
rect 3136 818 3170 834
rect 3250 1010 3284 1026
rect 3250 818 3284 834
rect 3346 1010 3380 1026
rect 3346 818 3380 834
rect 3460 1010 3494 1026
rect 3460 818 3494 834
rect 3556 1010 3590 1026
rect 3556 818 3590 834
rect 3670 1010 3704 1026
rect 3670 818 3704 834
rect 3766 1010 3800 1026
rect 3766 818 3800 834
rect 3880 1010 3914 1026
rect 3880 818 3914 834
rect 3976 1010 4010 1026
rect 3976 818 4010 834
rect 4090 1010 4124 1026
rect 4090 818 4124 834
rect 4186 1010 4220 1026
rect 4186 818 4220 834
rect 4300 1010 4334 1026
rect 4300 818 4334 834
rect 4396 1010 4430 1026
rect 4396 818 4430 834
rect 4510 1010 4544 1026
rect 4510 818 4544 834
rect 4606 1010 4640 1026
rect 4606 818 4640 834
rect 4720 1010 4754 1026
rect 4720 818 4754 834
rect 4816 1010 4850 1026
rect 4816 818 4850 834
rect 4930 1010 4964 1026
rect 4930 818 4964 834
rect 5026 1010 5060 1026
rect 5026 818 5060 834
rect 5140 1010 5174 1026
rect 5140 818 5174 834
rect 5236 1010 5270 1026
rect 5236 818 5270 834
rect 5350 1010 5384 1026
rect 5350 818 5384 834
rect 5446 1010 5480 1026
rect 5446 818 5480 834
rect 5560 1010 5594 1026
rect 5560 818 5594 834
rect 5656 1010 5690 1026
rect 5656 818 5690 834
rect 5770 1010 5804 1026
rect 5770 818 5804 834
rect 5866 1010 5900 1026
rect 5866 818 5900 834
rect 5980 1010 6014 1060
rect 5980 818 6014 834
rect 6076 1059 6192 1060
rect 6076 1010 6110 1059
rect 6076 818 6110 834
rect -2710 750 -2582 784
rect -2548 750 -2500 784
rect -2178 750 -2162 784
rect -2128 750 -2112 784
rect -1758 750 -1742 784
rect -1708 750 -1692 784
rect -1338 750 -1322 784
rect -1288 750 -1272 784
rect -918 750 -902 784
rect -868 750 -852 784
rect -498 750 -482 784
rect -448 750 -432 784
rect -78 750 -62 784
rect -28 750 -12 784
rect 342 750 358 784
rect 392 750 408 784
rect 762 750 778 784
rect 812 750 828 784
rect 1182 750 1198 784
rect 1232 750 1248 784
rect 1602 750 1618 784
rect 1652 750 1668 784
rect 2022 750 2038 784
rect 2072 750 2088 784
rect 2442 750 2458 784
rect 2492 750 2508 784
rect 2862 750 2878 784
rect 2912 750 2928 784
rect 3282 750 3298 784
rect 3332 750 3348 784
rect 3702 750 3718 784
rect 3752 750 3768 784
rect 4122 750 4138 784
rect 4172 750 4188 784
rect 4542 750 4558 784
rect 4592 750 4608 784
rect 4962 750 4978 784
rect 5012 750 5028 784
rect 5382 750 5398 784
rect 5432 750 5448 784
rect 5802 750 5818 784
rect 5852 750 5868 784
rect -2744 682 -2710 745
rect 7180 5518 7214 5580
rect 6827 5466 6843 5500
rect 7019 5466 7180 5500
rect 7078 5452 7112 5466
rect 6750 5356 6784 5372
rect 6827 5370 6843 5404
rect 7019 5370 7035 5404
rect 7078 5402 7112 5418
rect 6750 5306 6784 5322
rect 6827 5274 6843 5308
rect 7019 5274 7035 5308
rect 7078 5260 7112 5276
rect 6750 5164 6784 5180
rect 6827 5178 6843 5212
rect 7019 5178 7035 5212
rect 7078 5210 7112 5226
rect 6750 5114 6784 5130
rect 6827 5082 6843 5116
rect 7019 5082 7035 5116
rect 7078 5068 7112 5084
rect 6750 4972 6784 4988
rect 6827 4986 6843 5020
rect 7019 4986 7035 5020
rect 7078 5018 7112 5034
rect 6750 4922 6784 4938
rect 6827 4890 6843 4924
rect 7019 4890 7035 4924
rect 7078 4876 7112 4892
rect 6750 4780 6784 4796
rect 6827 4794 6843 4828
rect 7019 4794 7035 4828
rect 7078 4826 7112 4842
rect 6750 4730 6784 4746
rect 6827 4698 6843 4732
rect 7019 4698 7035 4732
rect 7078 4684 7112 4700
rect 6750 4588 6784 4604
rect 6827 4602 6843 4636
rect 7019 4602 7035 4636
rect 7078 4634 7112 4650
rect 6750 4538 6784 4554
rect 6827 4506 6843 4540
rect 7019 4506 7035 4540
rect 7078 4492 7112 4508
rect 6750 4396 6784 4412
rect 6827 4410 6843 4444
rect 7019 4410 7035 4444
rect 7078 4442 7112 4458
rect 6750 4346 6784 4362
rect 6827 4314 6843 4348
rect 7019 4314 7035 4348
rect 7078 4300 7112 4316
rect 6750 4204 6784 4220
rect 6827 4218 6843 4252
rect 7019 4218 7035 4252
rect 7078 4250 7112 4266
rect 6750 4154 6784 4170
rect 6827 4122 6843 4156
rect 7019 4122 7035 4156
rect 7078 4108 7112 4124
rect 6750 4012 6784 4028
rect 6827 4026 6843 4060
rect 7019 4026 7035 4060
rect 7078 4058 7112 4074
rect 6750 3962 6784 3978
rect 6827 3930 6843 3964
rect 7019 3930 7035 3964
rect 7078 3916 7112 3932
rect 6750 3820 6784 3836
rect 6827 3834 6843 3868
rect 7019 3834 7035 3868
rect 7078 3866 7112 3882
rect 6750 3772 6784 3786
rect 6682 3738 6843 3772
rect 7019 3738 7035 3772
rect 6648 3658 6682 3720
rect 7180 3658 7214 3720
rect 6648 3624 6744 3658
rect 7118 3624 7214 3658
rect 6192 682 6226 745
rect -2744 648 -2647 682
rect 6129 648 6226 682
rect -24 358 72 392
rect 3406 358 3502 392
rect -24 296 10 358
rect 3468 296 3502 358
rect 266 256 282 290
rect 316 256 332 290
rect 458 256 474 290
rect 508 256 524 290
rect 650 256 666 290
rect 700 256 716 290
rect 842 256 858 290
rect 892 256 908 290
rect 1034 256 1050 290
rect 1084 256 1100 290
rect 1226 256 1242 290
rect 1276 256 1292 290
rect 1418 256 1434 290
rect 1468 256 1484 290
rect 1610 256 1626 290
rect 1660 256 1676 290
rect 1802 256 1818 290
rect 1852 256 1868 290
rect 1994 256 2010 290
rect 2044 256 2060 290
rect 2186 256 2202 290
rect 2236 256 2252 290
rect 2378 256 2394 290
rect 2428 256 2444 290
rect 2570 256 2586 290
rect 2620 256 2636 290
rect 2762 256 2778 290
rect 2812 256 2828 290
rect 2954 256 2970 290
rect 3004 256 3020 290
rect 3146 256 3162 290
rect 3196 256 3212 290
rect -24 -122 10 -60
rect 90 206 124 222
rect 90 -20 124 30
rect 186 206 220 222
rect 186 14 220 30
rect 282 206 316 222
rect 90 -54 138 -20
rect 172 -54 188 -20
rect 90 -122 124 -54
rect 282 -122 316 29
rect 378 206 412 222
rect 378 14 412 30
rect 474 206 508 222
rect 474 -122 508 29
rect 570 206 604 222
rect 570 14 604 30
rect 666 206 700 222
rect 666 -122 700 29
rect 762 206 796 222
rect 762 14 796 30
rect 858 206 892 222
rect 858 -122 892 29
rect 954 206 988 222
rect 954 14 988 30
rect 1050 206 1084 222
rect 1050 -122 1084 29
rect 1146 206 1180 222
rect 1146 14 1180 30
rect 1242 206 1276 222
rect 1242 -122 1276 29
rect 1338 206 1372 222
rect 1338 14 1372 30
rect 1434 206 1468 222
rect 1434 -122 1468 29
rect 1530 206 1564 222
rect 1530 14 1564 30
rect 1626 206 1660 222
rect 1626 -122 1660 29
rect 1722 206 1756 222
rect 1722 14 1756 30
rect 1818 206 1852 222
rect 1818 -122 1852 29
rect 1914 206 1948 222
rect 1914 14 1948 30
rect 2010 206 2044 222
rect 2010 -122 2044 29
rect 2106 206 2140 222
rect 2106 14 2140 30
rect 2202 206 2236 222
rect 2202 -122 2236 29
rect 2298 206 2332 222
rect 2298 14 2332 30
rect 2394 206 2428 222
rect 2394 -122 2428 29
rect 2490 206 2524 222
rect 2490 14 2524 30
rect 2586 206 2620 222
rect 2586 -122 2620 29
rect 2682 206 2716 222
rect 2682 14 2716 30
rect 2778 206 2812 222
rect 2778 -122 2812 29
rect 2874 206 2908 222
rect 2874 14 2908 30
rect 2970 206 3004 222
rect 2970 -122 3004 29
rect 3066 206 3100 222
rect 3066 14 3100 30
rect 3162 206 3196 222
rect 3162 -122 3196 29
rect 3258 206 3292 222
rect 3258 14 3292 30
rect 3354 206 3388 222
rect 3354 -24 3388 30
rect 3290 -58 3306 -24
rect 3340 -58 3388 -24
rect 3354 -122 3388 -58
rect 3468 -122 3502 -60
rect -24 -156 72 -122
rect 3406 -156 3502 -122
<< viali >>
rect 1165 10570 1199 10604
rect 1165 10478 1199 10512
rect 1165 10386 1199 10420
rect 1165 10294 1199 10328
rect 1165 10202 1199 10236
rect 1165 10110 1199 10144
rect 1709 10570 1743 10604
rect 1709 10478 1743 10512
rect 1709 10386 1743 10420
rect 1709 10294 1743 10328
rect 1709 10202 1743 10236
rect 1709 10110 1743 10144
rect 2253 10570 2287 10604
rect 2253 10478 2287 10512
rect 2253 10386 2287 10420
rect 2253 10294 2287 10328
rect 2253 10202 2287 10236
rect 2253 10110 2287 10144
rect 1165 10018 1199 10052
rect 1165 9926 1199 9960
rect 1165 9834 1199 9868
rect 1165 9742 1199 9776
rect 1165 9650 1199 9684
rect 1165 9558 1199 9592
rect 1709 10018 1743 10052
rect 1709 9926 1743 9960
rect 1709 9834 1743 9868
rect 1709 9742 1743 9776
rect 1709 9650 1743 9684
rect 1709 9558 1743 9592
rect 2253 10018 2287 10052
rect 2253 9926 2287 9960
rect 2253 9834 2287 9868
rect 2253 9742 2287 9776
rect 2253 9650 2287 9684
rect 2253 9558 2287 9592
rect 1165 9466 1199 9500
rect 1709 9466 1743 9500
rect 2253 9466 2287 9500
rect 1165 9374 1199 9408
rect 1165 9282 1199 9316
rect 1165 9190 1199 9224
rect 1165 9098 1199 9132
rect 1709 9374 1743 9408
rect 1404 9322 1438 9356
rect 1404 9234 1438 9265
rect 1404 9231 1431 9234
rect 1431 9231 1438 9234
rect 1709 9282 1743 9316
rect 1709 9190 1743 9224
rect 1165 9006 1199 9040
rect 1165 8914 1199 8948
rect 1165 8822 1199 8856
rect 1165 8730 1199 8764
rect 1709 9098 1743 9132
rect 1709 9006 1743 9040
rect 2016 9330 2050 9364
rect 2015 9234 2049 9258
rect 2015 9224 2021 9234
rect 2021 9224 2049 9234
rect 2253 9374 2287 9408
rect 2253 9282 2287 9316
rect 2253 9190 2287 9224
rect 2253 9098 2287 9132
rect 1317 8982 1351 8989
rect 1317 8955 1343 8982
rect 1343 8955 1351 8982
rect 1403 8955 1437 8989
rect 1497 8948 1531 8982
rect 1599 8948 1633 8982
rect 1404 8746 1438 8780
rect 1709 8914 1743 8948
rect 1820 8948 1853 8982
rect 1853 8948 1854 8982
rect 1921 8948 1955 8982
rect 2016 8955 2050 8989
rect 2102 8982 2136 8989
rect 2102 8955 2109 8982
rect 2109 8955 2136 8982
rect 1709 8822 1743 8856
rect 1709 8730 1743 8764
rect 2012 8745 2046 8779
rect 1165 8638 1199 8672
rect 1404 8660 1438 8694
rect 1709 8638 1743 8672
rect 2012 8659 2046 8693
rect 2253 9006 2287 9040
rect 2253 8914 2287 8948
rect 2253 8822 2287 8856
rect 2253 8730 2287 8764
rect 2253 8638 2287 8672
rect 1165 8546 1199 8580
rect 1709 8546 1743 8580
rect 2253 8546 2287 8580
rect 1165 8454 1199 8488
rect 1306 8463 1341 8498
rect 1518 8489 1552 8497
rect 1518 8463 1528 8489
rect 1528 8463 1552 8489
rect 1709 8454 1743 8488
rect 1165 8362 1199 8396
rect 1898 8489 1932 8496
rect 1898 8462 1924 8489
rect 1924 8462 1932 8489
rect 2109 8462 2144 8497
rect 2253 8454 2287 8488
rect 1165 8270 1199 8304
rect 1397 8278 1431 8312
rect 1709 8362 1743 8396
rect 1709 8270 1743 8304
rect 2022 8312 2056 8313
rect 2022 8279 2055 8312
rect 2055 8279 2056 8312
rect 2253 8362 2287 8396
rect 2253 8270 2287 8304
rect -3656 7990 -3282 8023
rect -3656 7989 -3282 7990
rect -3415 7780 -3381 7813
rect -3415 7779 -3381 7780
rect -3322 7732 -3288 7766
rect -3557 7684 -3523 7717
rect -3557 7683 -3523 7684
rect -3650 7636 -3616 7670
rect -3415 7588 -3381 7621
rect -3415 7587 -3381 7588
rect -3322 7540 -3288 7574
rect -3557 7492 -3523 7525
rect -3557 7491 -3523 7492
rect -3650 7444 -3616 7478
rect -3415 7396 -3381 7429
rect -3415 7395 -3381 7396
rect -3322 7348 -3288 7382
rect -3557 7300 -3523 7333
rect -3557 7299 -3523 7300
rect -3650 7252 -3616 7286
rect -3415 7204 -3381 7237
rect -3415 7203 -3381 7204
rect -3322 7156 -3288 7190
rect -3557 7108 -3523 7141
rect -3557 7107 -3523 7108
rect -3650 7060 -3616 7094
rect -3415 7012 -3381 7045
rect -3415 7011 -3381 7012
rect -3322 6964 -3288 6998
rect -3557 6916 -3523 6949
rect -3557 6915 -3523 6916
rect -3650 6868 -3616 6902
rect -3415 6820 -3381 6853
rect -3415 6819 -3381 6820
rect -3322 6772 -3288 6806
rect -3557 6724 -3523 6757
rect -3557 6723 -3523 6724
rect -3650 6676 -3616 6710
rect -3415 6628 -3381 6661
rect -3415 6627 -3381 6628
rect -3322 6580 -3288 6614
rect -3557 6532 -3523 6565
rect -3557 6531 -3523 6532
rect -3650 6484 -3616 6518
rect -3415 6436 -3381 6469
rect -3415 6435 -3381 6436
rect -3322 6388 -3288 6422
rect -3557 6340 -3523 6373
rect -3557 6339 -3523 6340
rect -3650 6292 -3616 6326
rect -3415 6244 -3381 6277
rect -3415 6243 -3381 6244
rect -2662 7989 6114 8023
rect -2386 7887 -2352 7921
rect -1966 7887 -1932 7921
rect -1546 7887 -1512 7921
rect -1126 7887 -1092 7921
rect -706 7887 -672 7921
rect -286 7887 -252 7921
rect 134 7887 168 7921
rect 554 7887 588 7921
rect 974 7887 1008 7921
rect 1394 7887 1428 7921
rect 1814 7887 1848 7921
rect 2234 7887 2268 7921
rect 2654 7887 2688 7921
rect 3074 7887 3108 7921
rect 3494 7887 3528 7921
rect 3914 7887 3948 7921
rect 4334 7887 4368 7921
rect 4754 7887 4788 7921
rect 5174 7887 5208 7921
rect 5594 7887 5628 7921
rect -2434 7794 -2400 7828
rect -2338 7652 -2304 7686
rect -2224 7794 -2190 7828
rect -2128 7652 -2094 7686
rect -2014 7794 -1980 7828
rect -1918 7652 -1884 7686
rect -1804 7794 -1770 7828
rect -1708 7652 -1674 7686
rect -1594 7794 -1560 7828
rect -1498 7652 -1464 7686
rect -1384 7794 -1350 7828
rect -1288 7652 -1254 7686
rect -1174 7794 -1140 7828
rect -1078 7652 -1044 7686
rect -964 7794 -930 7828
rect -868 7652 -834 7686
rect -754 7794 -720 7828
rect -658 7652 -624 7686
rect -544 7794 -510 7828
rect -448 7652 -414 7686
rect -334 7794 -300 7828
rect -238 7652 -204 7686
rect -124 7794 -90 7828
rect -28 7652 6 7686
rect 86 7794 120 7828
rect 182 7652 216 7686
rect 296 7794 330 7828
rect 392 7652 426 7686
rect 506 7794 540 7828
rect 602 7652 636 7686
rect 716 7794 750 7828
rect 812 7652 846 7686
rect 926 7794 960 7828
rect 1022 7652 1056 7686
rect 1136 7794 1170 7828
rect 1232 7652 1266 7686
rect 1346 7794 1380 7828
rect 1442 7652 1476 7686
rect 1556 7794 1590 7828
rect 1652 7652 1686 7686
rect 1766 7794 1800 7828
rect 1862 7652 1896 7686
rect 1976 7794 2010 7828
rect 2072 7652 2106 7686
rect 2186 7794 2220 7828
rect 2282 7652 2316 7686
rect 2396 7794 2430 7828
rect 2492 7652 2526 7686
rect 2606 7794 2640 7828
rect 2702 7652 2736 7686
rect 2816 7794 2850 7828
rect 2912 7652 2946 7686
rect 3026 7794 3060 7828
rect 3122 7652 3156 7686
rect 3236 7794 3270 7828
rect 3332 7652 3366 7686
rect 3446 7794 3480 7828
rect 3542 7652 3576 7686
rect 3656 7794 3690 7828
rect 3752 7652 3786 7686
rect 3866 7794 3900 7828
rect 3962 7652 3996 7686
rect 4076 7794 4110 7828
rect 4172 7652 4206 7686
rect 4286 7794 4320 7828
rect 4382 7652 4416 7686
rect 4496 7794 4530 7828
rect 4592 7652 4626 7686
rect 4706 7794 4740 7828
rect 4802 7652 4836 7686
rect 4916 7794 4950 7828
rect 5012 7652 5046 7686
rect 5126 7794 5160 7828
rect 5222 7652 5256 7686
rect 5336 7794 5370 7828
rect 5432 7652 5466 7686
rect 5546 7794 5580 7828
rect 5642 7652 5676 7686
rect 5756 7794 5790 7828
rect 5852 7652 5886 7686
rect -2176 7559 -2142 7593
rect -1756 7559 -1722 7593
rect -1336 7559 -1302 7593
rect -916 7559 -882 7593
rect -496 7559 -462 7593
rect -76 7559 -42 7593
rect 344 7559 378 7593
rect 764 7559 798 7593
rect 1184 7559 1218 7593
rect 1604 7559 1638 7593
rect 2024 7559 2058 7593
rect 2444 7559 2478 7593
rect 2864 7559 2898 7593
rect 3284 7559 3318 7593
rect 3704 7559 3738 7593
rect 4124 7559 4158 7593
rect 4544 7559 4578 7593
rect 4964 7559 4998 7593
rect 5384 7559 5418 7593
rect 5804 7559 5838 7593
rect -2384 7355 -2350 7389
rect -1964 7355 -1930 7389
rect -1544 7355 -1510 7389
rect -1124 7355 -1090 7389
rect -704 7355 -670 7389
rect -284 7355 -250 7389
rect 136 7355 170 7389
rect 556 7355 590 7389
rect 976 7355 1010 7389
rect 1396 7355 1430 7389
rect 1816 7355 1850 7389
rect 2236 7355 2270 7389
rect 2656 7355 2690 7389
rect 3076 7355 3110 7389
rect 3496 7355 3530 7389
rect 3916 7355 3950 7389
rect 4336 7355 4370 7389
rect 4756 7355 4790 7389
rect 5176 7355 5210 7389
rect 5596 7355 5630 7389
rect -2432 7295 -2398 7296
rect -2432 7262 -2398 7295
rect -2336 7120 -2302 7154
rect -2222 7295 -2188 7296
rect -2222 7262 -2188 7295
rect -2126 7120 -2092 7154
rect -2012 7295 -1978 7296
rect -2012 7262 -1978 7295
rect -1916 7120 -1882 7154
rect -1802 7295 -1768 7296
rect -1802 7262 -1768 7295
rect -1706 7120 -1672 7154
rect -1592 7295 -1558 7296
rect -1592 7262 -1558 7295
rect -1496 7120 -1462 7154
rect -1382 7295 -1348 7296
rect -1382 7262 -1348 7295
rect -1286 7120 -1252 7154
rect -1172 7295 -1138 7296
rect -1172 7262 -1138 7295
rect -1076 7120 -1042 7154
rect -962 7295 -928 7296
rect -962 7262 -928 7295
rect -866 7120 -832 7154
rect -752 7295 -718 7296
rect -752 7262 -718 7295
rect -656 7120 -622 7154
rect -542 7295 -508 7296
rect -542 7262 -508 7295
rect -446 7120 -412 7154
rect -332 7295 -298 7296
rect -332 7262 -298 7295
rect -236 7120 -202 7154
rect -122 7295 -88 7296
rect -122 7262 -88 7295
rect -26 7120 8 7154
rect 88 7295 122 7296
rect 88 7262 122 7295
rect 184 7120 218 7154
rect 298 7295 332 7296
rect 298 7262 332 7295
rect 394 7120 428 7154
rect 508 7295 542 7296
rect 508 7262 542 7295
rect 604 7120 638 7154
rect 718 7295 752 7296
rect 718 7262 752 7295
rect 814 7120 848 7154
rect 928 7295 962 7296
rect 928 7262 962 7295
rect 1024 7120 1058 7154
rect 1138 7295 1172 7296
rect 1138 7262 1172 7295
rect 1234 7120 1268 7154
rect 1348 7295 1382 7296
rect 1348 7262 1382 7295
rect 1444 7120 1478 7154
rect 1558 7295 1592 7296
rect 1558 7262 1592 7295
rect 1654 7120 1688 7154
rect 1768 7295 1802 7296
rect 1768 7262 1802 7295
rect 1864 7120 1898 7154
rect 1978 7295 2012 7296
rect 1978 7262 2012 7295
rect 2074 7120 2108 7154
rect 2188 7295 2222 7296
rect 2188 7262 2222 7295
rect 2284 7120 2318 7154
rect 2398 7295 2432 7296
rect 2398 7262 2432 7295
rect 2494 7120 2528 7154
rect 2608 7295 2642 7296
rect 2608 7262 2642 7295
rect 2704 7120 2738 7154
rect 2818 7295 2852 7296
rect 2818 7262 2852 7295
rect 2914 7120 2948 7154
rect 3028 7295 3062 7296
rect 3028 7262 3062 7295
rect 3124 7120 3158 7154
rect 3238 7295 3272 7296
rect 3238 7262 3272 7295
rect 3334 7120 3368 7154
rect 3448 7295 3482 7296
rect 3448 7262 3482 7295
rect 3544 7120 3578 7154
rect 3658 7295 3692 7296
rect 3658 7262 3692 7295
rect 3754 7120 3788 7154
rect 3868 7295 3902 7296
rect 3868 7262 3902 7295
rect 3964 7120 3998 7154
rect 4078 7295 4112 7296
rect 4078 7262 4112 7295
rect 4174 7120 4208 7154
rect 4288 7295 4322 7296
rect 4288 7262 4322 7295
rect 4384 7120 4418 7154
rect 4498 7295 4532 7296
rect 4498 7262 4532 7295
rect 4594 7120 4628 7154
rect 4708 7295 4742 7296
rect 4708 7262 4742 7295
rect 4804 7120 4838 7154
rect 4918 7295 4952 7296
rect 4918 7262 4952 7295
rect 5014 7120 5048 7154
rect 5128 7295 5162 7296
rect 5128 7262 5162 7295
rect 5224 7120 5258 7154
rect 5338 7295 5372 7296
rect 5338 7262 5372 7295
rect 5434 7120 5468 7154
rect 5548 7295 5582 7296
rect 5548 7262 5582 7295
rect 5644 7120 5678 7154
rect 5758 7295 5792 7296
rect 5758 7262 5792 7295
rect 5854 7120 5888 7154
rect -2174 7026 -2140 7060
rect -1754 7026 -1720 7060
rect -1334 7026 -1300 7060
rect -914 7026 -880 7060
rect -494 7026 -460 7060
rect -74 7026 -40 7060
rect 346 7026 380 7060
rect 766 7026 800 7060
rect 1186 7026 1220 7060
rect 1606 7026 1640 7060
rect 2026 7026 2060 7060
rect 2446 7026 2480 7060
rect 2866 7026 2900 7060
rect 3286 7026 3320 7060
rect 3706 7026 3740 7060
rect 4126 7026 4160 7060
rect 4546 7026 4580 7060
rect 4966 7026 5000 7060
rect 5386 7026 5420 7060
rect 5806 7026 5840 7060
rect 6744 7990 7118 8023
rect 6744 7989 7118 7990
rect -3656 6034 -3282 6067
rect -3656 6033 -3282 6034
rect -3656 5580 -3654 5613
rect -3654 5580 -3282 5613
rect -3656 5579 -3282 5580
rect -3415 5370 -3381 5403
rect -3415 5369 -3381 5370
rect -3320 5322 -3286 5356
rect -3557 5274 -3555 5307
rect -3555 5274 -3523 5307
rect -3557 5273 -3523 5274
rect -3648 5226 -3614 5260
rect -3415 5178 -3381 5211
rect -3415 5177 -3381 5178
rect -3320 5130 -3286 5164
rect -3557 5082 -3555 5115
rect -3555 5082 -3523 5115
rect -3557 5081 -3523 5082
rect -3648 5034 -3614 5068
rect -3415 4986 -3381 5019
rect -3415 4985 -3381 4986
rect -3320 4938 -3286 4972
rect -3557 4890 -3555 4923
rect -3555 4890 -3523 4923
rect -3557 4889 -3523 4890
rect -3648 4842 -3614 4876
rect -3415 4794 -3381 4827
rect -3415 4793 -3381 4794
rect -3320 4746 -3286 4780
rect -3557 4698 -3555 4731
rect -3555 4698 -3523 4731
rect -3557 4697 -3523 4698
rect -3648 4650 -3614 4684
rect -3415 4602 -3381 4635
rect -3415 4601 -3381 4602
rect -3320 4554 -3286 4588
rect -3557 4506 -3555 4539
rect -3555 4506 -3523 4539
rect -3557 4505 -3523 4506
rect -3648 4458 -3614 4492
rect -3415 4410 -3381 4443
rect -3415 4409 -3381 4410
rect -3320 4362 -3286 4396
rect -3557 4314 -3555 4347
rect -3555 4314 -3523 4347
rect -3557 4313 -3523 4314
rect -3648 4266 -3614 4300
rect -3415 4218 -3381 4251
rect -3415 4217 -3381 4218
rect -3320 4170 -3286 4204
rect -3557 4122 -3555 4155
rect -3555 4122 -3523 4155
rect -3557 4121 -3523 4122
rect -3648 4074 -3614 4108
rect -3415 4026 -3381 4059
rect -3415 4025 -3381 4026
rect -3320 3978 -3286 4012
rect -3557 3930 -3555 3963
rect -3555 3930 -3523 3963
rect -3557 3929 -3523 3930
rect -3648 3882 -3614 3916
rect -3415 3834 -3381 3867
rect -3415 3833 -3381 3834
rect -2744 4759 -2710 6435
rect -2372 6395 -2338 6429
rect -1952 6395 -1918 6429
rect -1532 6395 -1498 6429
rect -1112 6395 -1078 6429
rect -692 6395 -658 6429
rect -272 6395 -238 6429
rect 148 6395 182 6429
rect 568 6395 602 6429
rect 988 6395 1022 6429
rect 1408 6395 1442 6429
rect 1828 6395 1862 6429
rect 2248 6395 2282 6429
rect 2668 6395 2702 6429
rect 3088 6395 3122 6429
rect 3508 6395 3542 6429
rect 3928 6395 3962 6429
rect 4348 6395 4382 6429
rect 4768 6395 4802 6429
rect 5188 6395 5222 6429
rect 5608 6395 5642 6429
rect -2420 6311 -2386 6345
rect -2324 6169 -2290 6203
rect -2210 6311 -2176 6345
rect -2114 6169 -2080 6203
rect -2000 6311 -1966 6345
rect -1904 6169 -1870 6203
rect -1790 6311 -1756 6345
rect -1694 6169 -1660 6203
rect -1580 6311 -1546 6345
rect -1484 6169 -1450 6203
rect -1370 6311 -1336 6345
rect -1274 6169 -1240 6203
rect -1160 6311 -1126 6345
rect -1064 6169 -1030 6203
rect -950 6311 -916 6345
rect -854 6169 -820 6203
rect -740 6311 -706 6345
rect -644 6169 -610 6203
rect -530 6311 -496 6345
rect -434 6169 -400 6203
rect -320 6311 -286 6345
rect -224 6169 -190 6203
rect -110 6311 -76 6345
rect -14 6169 20 6203
rect 100 6311 134 6345
rect 196 6169 230 6203
rect 310 6311 344 6345
rect 406 6169 440 6203
rect 520 6311 554 6345
rect 616 6169 650 6203
rect 730 6311 764 6345
rect 826 6169 860 6203
rect 940 6311 974 6345
rect 1036 6169 1070 6203
rect 1150 6311 1184 6345
rect 1246 6169 1280 6203
rect 1360 6311 1394 6345
rect 1456 6169 1490 6203
rect 1570 6311 1604 6345
rect 1666 6169 1700 6203
rect 1780 6311 1814 6345
rect 1876 6169 1910 6203
rect 1990 6311 2024 6345
rect 2086 6169 2120 6203
rect 2200 6311 2234 6345
rect 2296 6169 2330 6203
rect 2410 6311 2444 6345
rect 2506 6169 2540 6203
rect 2620 6311 2654 6345
rect 2716 6169 2750 6203
rect 2830 6311 2864 6345
rect 2926 6169 2960 6203
rect 3040 6311 3074 6345
rect 3136 6169 3170 6203
rect 3250 6311 3284 6345
rect 3346 6169 3380 6203
rect 3460 6311 3494 6345
rect 3556 6169 3590 6203
rect 3670 6311 3704 6345
rect 3766 6169 3800 6203
rect 3880 6311 3914 6345
rect 3976 6169 4010 6203
rect 4090 6311 4124 6345
rect 4186 6169 4220 6203
rect 4300 6311 4334 6345
rect 4396 6169 4430 6203
rect 4510 6311 4544 6345
rect 4606 6169 4640 6203
rect 4720 6311 4754 6345
rect 4816 6169 4850 6203
rect 4930 6311 4964 6345
rect 5026 6169 5060 6203
rect 5140 6311 5174 6345
rect 5236 6169 5270 6203
rect 5350 6311 5384 6345
rect 5446 6169 5480 6203
rect 5560 6311 5594 6345
rect 5656 6169 5690 6203
rect 5770 6311 5804 6345
rect 5866 6169 5900 6203
rect -2162 6085 -2128 6119
rect -1742 6085 -1708 6119
rect -1322 6085 -1288 6119
rect -902 6085 -868 6119
rect -482 6085 -448 6119
rect -62 6085 -28 6119
rect 358 6085 392 6119
rect 778 6085 812 6119
rect 1198 6085 1232 6119
rect 1618 6085 1652 6119
rect 2038 6085 2072 6119
rect 2458 6085 2492 6119
rect 2878 6085 2912 6119
rect 3298 6085 3332 6119
rect 3718 6085 3752 6119
rect 4138 6085 4172 6119
rect 4558 6085 4592 6119
rect 4978 6085 5012 6119
rect 5398 6085 5432 6119
rect 5818 6085 5852 6119
rect -2372 5955 -2338 5989
rect -1952 5955 -1918 5989
rect -1532 5955 -1498 5989
rect -1112 5955 -1078 5989
rect -692 5955 -658 5989
rect -272 5955 -238 5989
rect 148 5955 182 5989
rect 568 5955 602 5989
rect 988 5955 1022 5989
rect 1408 5955 1442 5989
rect 1828 5955 1862 5989
rect 2248 5955 2282 5989
rect 2668 5955 2702 5989
rect 3088 5955 3122 5989
rect 3508 5955 3542 5989
rect 3928 5955 3962 5989
rect 4348 5955 4382 5989
rect 4768 5955 4802 5989
rect 5188 5955 5222 5989
rect 5608 5955 5642 5989
rect -2420 5871 -2386 5905
rect -2324 5729 -2290 5763
rect -2210 5871 -2176 5905
rect -2114 5729 -2080 5763
rect -2000 5871 -1966 5905
rect -1904 5729 -1870 5763
rect -1790 5871 -1756 5905
rect -1694 5729 -1660 5763
rect -1580 5871 -1546 5905
rect -1484 5729 -1450 5763
rect -1370 5871 -1336 5905
rect -1274 5729 -1240 5763
rect -1160 5871 -1126 5905
rect -1064 5729 -1030 5763
rect -950 5871 -916 5905
rect -854 5729 -820 5763
rect -740 5871 -706 5905
rect -644 5729 -610 5763
rect -530 5871 -496 5905
rect -434 5729 -400 5763
rect -320 5871 -286 5905
rect -224 5729 -190 5763
rect -110 5871 -76 5905
rect -14 5729 20 5763
rect 100 5871 134 5905
rect 196 5729 230 5763
rect 310 5871 344 5905
rect 406 5729 440 5763
rect 520 5871 554 5905
rect 616 5729 650 5763
rect 730 5871 764 5905
rect 826 5729 860 5763
rect 940 5871 974 5905
rect 1036 5729 1070 5763
rect 1150 5871 1184 5905
rect 1246 5729 1280 5763
rect 1360 5871 1394 5905
rect 1456 5729 1490 5763
rect 1570 5871 1604 5905
rect 1666 5729 1700 5763
rect 1780 5871 1814 5905
rect 1876 5729 1910 5763
rect 1990 5871 2024 5905
rect 2086 5729 2120 5763
rect 2200 5871 2234 5905
rect 2296 5729 2330 5763
rect 2410 5871 2444 5905
rect 2506 5729 2540 5763
rect 2620 5871 2654 5905
rect 2716 5729 2750 5763
rect 2830 5871 2864 5905
rect 2926 5729 2960 5763
rect 3040 5871 3074 5905
rect 3136 5729 3170 5763
rect 3250 5871 3284 5905
rect 3346 5729 3380 5763
rect 3460 5871 3494 5905
rect 3556 5729 3590 5763
rect 3670 5871 3704 5905
rect 3766 5729 3800 5763
rect 3880 5871 3914 5905
rect 3976 5729 4010 5763
rect 4090 5871 4124 5905
rect 4186 5729 4220 5763
rect 4300 5871 4334 5905
rect 4396 5729 4430 5763
rect 4510 5871 4544 5905
rect 4606 5729 4640 5763
rect 4720 5871 4754 5905
rect 4816 5729 4850 5763
rect 4930 5871 4964 5905
rect 5026 5729 5060 5763
rect 5140 5871 5174 5905
rect 5236 5729 5270 5763
rect 5350 5871 5384 5905
rect 5446 5729 5480 5763
rect 5560 5871 5594 5905
rect 5656 5729 5690 5763
rect 5770 5871 5804 5905
rect 5866 5729 5900 5763
rect -2162 5645 -2128 5679
rect -1742 5645 -1708 5679
rect -1322 5645 -1288 5679
rect -902 5645 -868 5679
rect -482 5645 -448 5679
rect -62 5645 -28 5679
rect 358 5645 392 5679
rect 778 5645 812 5679
rect 1198 5645 1232 5679
rect 1618 5645 1652 5679
rect 2038 5645 2072 5679
rect 2458 5645 2492 5679
rect 2878 5645 2912 5679
rect 3298 5645 3332 5679
rect 3718 5645 3752 5679
rect 4138 5645 4172 5679
rect 4558 5645 4592 5679
rect 4978 5645 5012 5679
rect 5398 5645 5432 5679
rect 5818 5645 5852 5679
rect -2372 5515 -2338 5549
rect -1952 5515 -1918 5549
rect -1532 5515 -1498 5549
rect -1112 5515 -1078 5549
rect -692 5515 -658 5549
rect -272 5515 -238 5549
rect 148 5515 182 5549
rect 568 5515 602 5549
rect 988 5515 1022 5549
rect 1408 5515 1442 5549
rect 1828 5515 1862 5549
rect 2248 5515 2282 5549
rect 2668 5515 2702 5549
rect 3088 5515 3122 5549
rect 3508 5515 3542 5549
rect 3928 5515 3962 5549
rect 4348 5515 4382 5549
rect 4768 5515 4802 5549
rect 5188 5515 5222 5549
rect 5608 5515 5642 5549
rect -2420 5431 -2386 5465
rect -2324 5289 -2290 5323
rect -2210 5431 -2176 5465
rect -2114 5289 -2080 5323
rect -2000 5431 -1966 5465
rect -1904 5289 -1870 5323
rect -1790 5431 -1756 5465
rect -1694 5289 -1660 5323
rect -1580 5431 -1546 5465
rect -1484 5289 -1450 5323
rect -1370 5431 -1336 5465
rect -1274 5289 -1240 5323
rect -1160 5431 -1126 5465
rect -1064 5289 -1030 5323
rect -950 5431 -916 5465
rect -854 5289 -820 5323
rect -740 5431 -706 5465
rect -644 5289 -610 5323
rect -530 5431 -496 5465
rect -434 5289 -400 5323
rect -320 5431 -286 5465
rect -224 5289 -190 5323
rect -110 5431 -76 5465
rect -14 5289 20 5323
rect 100 5431 134 5465
rect 196 5289 230 5323
rect 310 5431 344 5465
rect 406 5289 440 5323
rect 520 5431 554 5465
rect 616 5289 650 5323
rect 730 5431 764 5465
rect 826 5289 860 5323
rect 940 5431 974 5465
rect 1036 5289 1070 5323
rect 1150 5431 1184 5465
rect 1246 5289 1280 5323
rect 1360 5431 1394 5465
rect 1456 5289 1490 5323
rect 1570 5431 1604 5465
rect 1666 5289 1700 5323
rect 1780 5431 1814 5465
rect 1876 5289 1910 5323
rect 1990 5431 2024 5465
rect 2086 5289 2120 5323
rect 2200 5431 2234 5465
rect 2296 5289 2330 5323
rect 2410 5431 2444 5465
rect 2506 5289 2540 5323
rect 2620 5431 2654 5465
rect 2716 5289 2750 5323
rect 2830 5431 2864 5465
rect 2926 5289 2960 5323
rect 3040 5431 3074 5465
rect 3136 5289 3170 5323
rect 3250 5431 3284 5465
rect 3346 5289 3380 5323
rect 3460 5431 3494 5465
rect 3556 5289 3590 5323
rect 3670 5431 3704 5465
rect 3766 5289 3800 5323
rect 3880 5431 3914 5465
rect 3976 5289 4010 5323
rect 4090 5431 4124 5465
rect 4186 5289 4220 5323
rect 4300 5431 4334 5465
rect 4396 5289 4430 5323
rect 4510 5431 4544 5465
rect 4606 5289 4640 5323
rect 4720 5431 4754 5465
rect 4816 5289 4850 5323
rect 4930 5431 4964 5465
rect 5026 5289 5060 5323
rect 5140 5431 5174 5465
rect 5236 5289 5270 5323
rect 5350 5431 5384 5465
rect 5446 5289 5480 5323
rect 5560 5431 5594 5465
rect 5656 5289 5690 5323
rect 5770 5431 5804 5465
rect 5866 5289 5900 5323
rect -2162 5205 -2128 5239
rect -1742 5205 -1708 5239
rect -1322 5205 -1288 5239
rect -902 5205 -868 5239
rect -482 5205 -448 5239
rect -62 5205 -28 5239
rect 358 5205 392 5239
rect 778 5205 812 5239
rect 1198 5205 1232 5239
rect 1618 5205 1652 5239
rect 2038 5205 2072 5239
rect 2458 5205 2492 5239
rect 2878 5205 2912 5239
rect 3298 5205 3332 5239
rect 3718 5205 3752 5239
rect 4138 5205 4172 5239
rect 4558 5205 4592 5239
rect 4978 5205 5012 5239
rect 5398 5205 5432 5239
rect 5818 5205 5852 5239
rect -2372 5075 -2338 5109
rect -1952 5075 -1918 5109
rect -1532 5075 -1498 5109
rect -1112 5075 -1078 5109
rect -692 5075 -658 5109
rect -272 5075 -238 5109
rect 148 5075 182 5109
rect 568 5075 602 5109
rect 988 5075 1022 5109
rect 1408 5075 1442 5109
rect 1828 5075 1862 5109
rect 2248 5075 2282 5109
rect 2668 5075 2702 5109
rect 3088 5075 3122 5109
rect 3508 5075 3542 5109
rect 3928 5075 3962 5109
rect 4348 5075 4382 5109
rect 4768 5075 4802 5109
rect 5188 5075 5222 5109
rect 5608 5075 5642 5109
rect -2420 4991 -2386 5025
rect -2324 4849 -2290 4883
rect -2210 4991 -2176 5025
rect -2114 4849 -2080 4883
rect -2000 4991 -1966 5025
rect -1904 4849 -1870 4883
rect -1790 4991 -1756 5025
rect -1694 4849 -1660 4883
rect -1580 4991 -1546 5025
rect -1484 4849 -1450 4883
rect -1370 4991 -1336 5025
rect -1274 4849 -1240 4883
rect -1160 4991 -1126 5025
rect -1064 4849 -1030 4883
rect -950 4991 -916 5025
rect -854 4849 -820 4883
rect -740 4991 -706 5025
rect -644 4849 -610 4883
rect -530 4991 -496 5025
rect -434 4849 -400 4883
rect -320 4991 -286 5025
rect -224 4849 -190 4883
rect -110 4991 -76 5025
rect -14 4849 20 4883
rect 100 4991 134 5025
rect 196 4849 230 4883
rect 310 4991 344 5025
rect 406 4849 440 4883
rect 520 4991 554 5025
rect 616 4849 650 4883
rect 730 4991 764 5025
rect 826 4849 860 4883
rect 940 4991 974 5025
rect 1036 4849 1070 4883
rect 1150 4991 1184 5025
rect 1246 4849 1280 4883
rect 1360 4991 1394 5025
rect 1456 4849 1490 4883
rect 1570 4991 1604 5025
rect 1666 4849 1700 4883
rect 1780 4991 1814 5025
rect 1876 4849 1910 4883
rect 1990 4991 2024 5025
rect 2086 4849 2120 4883
rect 2200 4991 2234 5025
rect 2296 4849 2330 4883
rect 2410 4991 2444 5025
rect 2506 4849 2540 4883
rect 2620 4991 2654 5025
rect 2716 4849 2750 4883
rect 2830 4991 2864 5025
rect 2926 4849 2960 4883
rect 3040 4991 3074 5025
rect 3136 4849 3170 4883
rect 3250 4991 3284 5025
rect 3346 4849 3380 4883
rect 3460 4991 3494 5025
rect 3556 4849 3590 4883
rect 3670 4991 3704 5025
rect 3766 4849 3800 4883
rect 3880 4991 3914 5025
rect 3976 4849 4010 4883
rect 4090 4991 4124 5025
rect 4186 4849 4220 4883
rect 4300 4991 4334 5025
rect 4396 4849 4430 4883
rect 4510 4991 4544 5025
rect 4606 4849 4640 4883
rect 4720 4991 4754 5025
rect 4816 4849 4850 4883
rect 4930 4991 4964 5025
rect 5026 4849 5060 4883
rect 5140 4991 5174 5025
rect 5236 4849 5270 4883
rect 5350 4991 5384 5025
rect 5446 4849 5480 4883
rect 5560 4991 5594 5025
rect 5656 4849 5690 4883
rect 5770 4991 5804 5025
rect 5866 4849 5900 4883
rect -2162 4765 -2128 4799
rect -1742 4765 -1708 4799
rect -1322 4765 -1288 4799
rect -902 4765 -868 4799
rect -482 4765 -448 4799
rect -62 4765 -28 4799
rect 358 4765 392 4799
rect 778 4765 812 4799
rect 1198 4765 1232 4799
rect 1618 4765 1652 4799
rect 2038 4765 2072 4799
rect 2458 4765 2492 4799
rect 2878 4765 2912 4799
rect 3298 4765 3332 4799
rect 3718 4765 3752 4799
rect 4138 4765 4172 4799
rect 4558 4765 4592 4799
rect 4978 4765 5012 4799
rect 5398 4765 5432 4799
rect 5818 4765 5852 4799
rect 6192 4759 6226 6435
rect 6843 7780 6877 7813
rect 6843 7779 6877 7780
rect 6750 7732 6784 7766
rect 6985 7684 7019 7717
rect 6985 7683 7019 7684
rect 7078 7636 7112 7670
rect 6843 7588 6877 7621
rect 6843 7587 6877 7588
rect 6750 7540 6784 7574
rect 6985 7492 7019 7525
rect 6985 7491 7019 7492
rect 7078 7444 7112 7478
rect 6843 7396 6877 7429
rect 6843 7395 6877 7396
rect 6750 7348 6784 7382
rect 6985 7300 7019 7333
rect 6985 7299 7019 7300
rect 7078 7252 7112 7286
rect 6843 7204 6877 7237
rect 6843 7203 6877 7204
rect 6750 7156 6784 7190
rect 6985 7108 7019 7141
rect 6985 7107 7019 7108
rect 7078 7060 7112 7094
rect 6843 7012 6877 7045
rect 6843 7011 6877 7012
rect 6750 6964 6784 6998
rect 6985 6916 7019 6949
rect 6985 6915 7019 6916
rect 7078 6868 7112 6902
rect 6843 6820 6877 6853
rect 6843 6819 6877 6820
rect 6750 6772 6784 6806
rect 6985 6724 7019 6757
rect 6985 6723 7019 6724
rect 7078 6676 7112 6710
rect 6843 6628 6877 6661
rect 6843 6627 6877 6628
rect 6750 6580 6784 6614
rect 6985 6532 7019 6565
rect 6985 6531 7019 6532
rect 7078 6484 7112 6518
rect 6843 6436 6877 6469
rect 6843 6435 6877 6436
rect 6750 6388 6784 6422
rect 6985 6340 7019 6373
rect 6985 6339 7019 6340
rect 7078 6292 7112 6326
rect 6843 6244 6877 6277
rect 6843 6243 6877 6244
rect 6744 6034 7118 6067
rect 6744 6033 7118 6034
rect 6744 5580 7118 5613
rect 6744 5579 7118 5580
rect -3656 3624 -3654 3657
rect -3654 3624 -3282 3657
rect -3656 3623 -3282 3624
rect -2744 745 -2710 4180
rect -2372 4140 -2338 4174
rect -1952 4140 -1918 4174
rect -1532 4140 -1498 4174
rect -1112 4140 -1078 4174
rect -692 4140 -658 4174
rect -272 4140 -238 4174
rect 148 4140 182 4174
rect 568 4140 602 4174
rect 988 4140 1022 4174
rect 1408 4140 1442 4174
rect 1828 4140 1862 4174
rect 2248 4140 2282 4174
rect 2668 4140 2702 4174
rect 3088 4140 3122 4174
rect 3508 4140 3542 4174
rect 3928 4140 3962 4174
rect 4348 4140 4382 4174
rect 4768 4140 4802 4174
rect 5188 4140 5222 4174
rect 5608 4140 5642 4174
rect -2420 4056 -2386 4090
rect -2324 3914 -2290 3948
rect -2210 4056 -2176 4090
rect -2114 3914 -2080 3948
rect -2000 4056 -1966 4090
rect -1904 3914 -1870 3948
rect -1790 4056 -1756 4090
rect -1694 3914 -1660 3948
rect -1580 4056 -1546 4090
rect -1484 3914 -1450 3948
rect -1370 4056 -1336 4090
rect -1274 3914 -1240 3948
rect -1160 4056 -1126 4090
rect -1064 3914 -1030 3948
rect -950 4056 -916 4090
rect -854 3914 -820 3948
rect -740 4056 -706 4090
rect -644 3914 -610 3948
rect -530 4056 -496 4090
rect -434 3914 -400 3948
rect -320 4056 -286 4090
rect -224 3914 -190 3948
rect -110 4056 -76 4090
rect -14 3914 20 3948
rect 100 4056 134 4090
rect 196 3914 230 3948
rect 310 4056 344 4090
rect 406 3914 440 3948
rect 520 4056 554 4090
rect 616 3914 650 3948
rect 730 4056 764 4090
rect 826 3914 860 3948
rect 940 4056 974 4090
rect 1036 3914 1070 3948
rect 1150 4056 1184 4090
rect 1246 3914 1280 3948
rect 1360 4056 1394 4090
rect 1456 3914 1490 3948
rect 1570 4056 1604 4090
rect 1666 3914 1700 3948
rect 1780 4056 1814 4090
rect 1876 3914 1910 3948
rect 1990 4056 2024 4090
rect 2086 3914 2120 3948
rect 2200 4056 2234 4090
rect 2296 3914 2330 3948
rect 2410 4056 2444 4090
rect 2506 3914 2540 3948
rect 2620 4056 2654 4090
rect 2716 3914 2750 3948
rect 2830 4056 2864 4090
rect 2926 3914 2960 3948
rect 3040 4056 3074 4090
rect 3136 3914 3170 3948
rect 3250 4056 3284 4090
rect 3346 3914 3380 3948
rect 3460 4056 3494 4090
rect 3556 3914 3590 3948
rect 3670 4056 3704 4090
rect 3766 3914 3800 3948
rect 3880 4056 3914 4090
rect 3976 3914 4010 3948
rect 4090 4056 4124 4090
rect 4186 3914 4220 3948
rect 4300 4056 4334 4090
rect 4396 3914 4430 3948
rect 4510 4056 4544 4090
rect 4606 3914 4640 3948
rect 4720 4056 4754 4090
rect 4816 3914 4850 3948
rect 4930 4056 4964 4090
rect 5026 3914 5060 3948
rect 5140 4056 5174 4090
rect 5236 3914 5270 3948
rect 5350 4056 5384 4090
rect 5446 3914 5480 3948
rect 5560 4056 5594 4090
rect 5656 3914 5690 3948
rect 5770 4056 5804 4090
rect 5866 3914 5900 3948
rect -2162 3830 -2128 3864
rect -1742 3830 -1708 3864
rect -1322 3830 -1288 3864
rect -902 3830 -868 3864
rect -482 3830 -448 3864
rect -62 3830 -28 3864
rect 358 3830 392 3864
rect 778 3830 812 3864
rect 1198 3830 1232 3864
rect 1618 3830 1652 3864
rect 2038 3830 2072 3864
rect 2458 3830 2492 3864
rect 2878 3830 2912 3864
rect 3298 3830 3332 3864
rect 3718 3830 3752 3864
rect 4138 3830 4172 3864
rect 4558 3830 4592 3864
rect 4978 3830 5012 3864
rect 5398 3830 5432 3864
rect 5818 3830 5852 3864
rect -2372 3700 -2338 3734
rect -1952 3700 -1918 3734
rect -1532 3700 -1498 3734
rect -1112 3700 -1078 3734
rect -692 3700 -658 3734
rect -272 3700 -238 3734
rect 148 3700 182 3734
rect 568 3700 602 3734
rect 988 3700 1022 3734
rect 1408 3700 1442 3734
rect 1828 3700 1862 3734
rect 2248 3700 2282 3734
rect 2668 3700 2702 3734
rect 3088 3700 3122 3734
rect 3508 3700 3542 3734
rect 3928 3700 3962 3734
rect 4348 3700 4382 3734
rect 4768 3700 4802 3734
rect 5188 3700 5222 3734
rect 5608 3700 5642 3734
rect -2420 3616 -2386 3650
rect -2324 3474 -2290 3508
rect -2210 3616 -2176 3650
rect -2114 3474 -2080 3508
rect -2000 3616 -1966 3650
rect -1904 3474 -1870 3508
rect -1790 3616 -1756 3650
rect -1694 3474 -1660 3508
rect -1580 3616 -1546 3650
rect -1484 3474 -1450 3508
rect -1370 3616 -1336 3650
rect -1274 3474 -1240 3508
rect -1160 3616 -1126 3650
rect -1064 3474 -1030 3508
rect -950 3616 -916 3650
rect -854 3474 -820 3508
rect -740 3616 -706 3650
rect -644 3474 -610 3508
rect -530 3616 -496 3650
rect -434 3474 -400 3508
rect -320 3616 -286 3650
rect -224 3474 -190 3508
rect -110 3616 -76 3650
rect -14 3474 20 3508
rect 100 3616 134 3650
rect 196 3474 230 3508
rect 310 3616 344 3650
rect 406 3474 440 3508
rect 520 3616 554 3650
rect 616 3474 650 3508
rect 730 3616 764 3650
rect 826 3474 860 3508
rect 940 3616 974 3650
rect 1036 3474 1070 3508
rect 1150 3616 1184 3650
rect 1246 3474 1280 3508
rect 1360 3616 1394 3650
rect 1456 3474 1490 3508
rect 1570 3616 1604 3650
rect 1666 3474 1700 3508
rect 1780 3616 1814 3650
rect 1876 3474 1910 3508
rect 1990 3616 2024 3650
rect 2086 3474 2120 3508
rect 2200 3616 2234 3650
rect 2296 3474 2330 3508
rect 2410 3616 2444 3650
rect 2506 3474 2540 3508
rect 2620 3616 2654 3650
rect 2716 3474 2750 3508
rect 2830 3616 2864 3650
rect 2926 3474 2960 3508
rect 3040 3616 3074 3650
rect 3136 3474 3170 3508
rect 3250 3616 3284 3650
rect 3346 3474 3380 3508
rect 3460 3616 3494 3650
rect 3556 3474 3590 3508
rect 3670 3616 3704 3650
rect 3766 3474 3800 3508
rect 3880 3616 3914 3650
rect 3976 3474 4010 3508
rect 4090 3616 4124 3650
rect 4186 3474 4220 3508
rect 4300 3616 4334 3650
rect 4396 3474 4430 3508
rect 4510 3616 4544 3650
rect 4606 3474 4640 3508
rect 4720 3616 4754 3650
rect 4816 3474 4850 3508
rect 4930 3616 4964 3650
rect 5026 3474 5060 3508
rect 5140 3616 5174 3650
rect 5236 3474 5270 3508
rect 5350 3616 5384 3650
rect 5446 3474 5480 3508
rect 5560 3616 5594 3650
rect 5656 3474 5690 3508
rect 5770 3616 5804 3650
rect 5866 3474 5900 3508
rect -2162 3390 -2128 3424
rect -1742 3390 -1708 3424
rect -1322 3390 -1288 3424
rect -902 3390 -868 3424
rect -482 3390 -448 3424
rect -62 3390 -28 3424
rect 358 3390 392 3424
rect 778 3390 812 3424
rect 1198 3390 1232 3424
rect 1618 3390 1652 3424
rect 2038 3390 2072 3424
rect 2458 3390 2492 3424
rect 2878 3390 2912 3424
rect 3298 3390 3332 3424
rect 3718 3390 3752 3424
rect 4138 3390 4172 3424
rect 4558 3390 4592 3424
rect 4978 3390 5012 3424
rect 5398 3390 5432 3424
rect 5818 3390 5852 3424
rect -2372 3260 -2338 3294
rect -1952 3260 -1918 3294
rect -1532 3260 -1498 3294
rect -1112 3260 -1078 3294
rect -692 3260 -658 3294
rect -272 3260 -238 3294
rect 148 3260 182 3294
rect 568 3260 602 3294
rect 988 3260 1022 3294
rect 1408 3260 1442 3294
rect 1828 3260 1862 3294
rect 2248 3260 2282 3294
rect 2668 3260 2702 3294
rect 3088 3260 3122 3294
rect 3508 3260 3542 3294
rect 3928 3260 3962 3294
rect 4348 3260 4382 3294
rect 4768 3260 4802 3294
rect 5188 3260 5222 3294
rect 5608 3260 5642 3294
rect -2420 3176 -2386 3210
rect -2324 3034 -2290 3068
rect -2210 3176 -2176 3210
rect -2114 3034 -2080 3068
rect -2000 3176 -1966 3210
rect -1904 3034 -1870 3068
rect -1790 3176 -1756 3210
rect -1694 3034 -1660 3068
rect -1580 3176 -1546 3210
rect -1484 3034 -1450 3068
rect -1370 3176 -1336 3210
rect -1274 3034 -1240 3068
rect -1160 3176 -1126 3210
rect -1064 3034 -1030 3068
rect -950 3176 -916 3210
rect -854 3034 -820 3068
rect -740 3176 -706 3210
rect -644 3034 -610 3068
rect -530 3176 -496 3210
rect -434 3034 -400 3068
rect -320 3176 -286 3210
rect -224 3034 -190 3068
rect -110 3176 -76 3210
rect -14 3034 20 3068
rect 100 3176 134 3210
rect 196 3034 230 3068
rect 310 3176 344 3210
rect 406 3034 440 3068
rect 520 3176 554 3210
rect 616 3034 650 3068
rect 730 3176 764 3210
rect 826 3034 860 3068
rect 940 3176 974 3210
rect 1036 3034 1070 3068
rect 1150 3176 1184 3210
rect 1246 3034 1280 3068
rect 1360 3176 1394 3210
rect 1456 3034 1490 3068
rect 1570 3176 1604 3210
rect 1666 3034 1700 3068
rect 1780 3176 1814 3210
rect 1876 3034 1910 3068
rect 1990 3176 2024 3210
rect 2086 3034 2120 3068
rect 2200 3176 2234 3210
rect 2296 3034 2330 3068
rect 2410 3176 2444 3210
rect 2506 3034 2540 3068
rect 2620 3176 2654 3210
rect 2716 3034 2750 3068
rect 2830 3176 2864 3210
rect 2926 3034 2960 3068
rect 3040 3176 3074 3210
rect 3136 3034 3170 3068
rect 3250 3176 3284 3210
rect 3346 3034 3380 3068
rect 3460 3176 3494 3210
rect 3556 3034 3590 3068
rect 3670 3176 3704 3210
rect 3766 3034 3800 3068
rect 3880 3176 3914 3210
rect 3976 3034 4010 3068
rect 4090 3176 4124 3210
rect 4186 3034 4220 3068
rect 4300 3176 4334 3210
rect 4396 3034 4430 3068
rect 4510 3176 4544 3210
rect 4606 3034 4640 3068
rect 4720 3176 4754 3210
rect 4816 3034 4850 3068
rect 4930 3176 4964 3210
rect 5026 3034 5060 3068
rect 5140 3176 5174 3210
rect 5236 3034 5270 3068
rect 5350 3176 5384 3210
rect 5446 3034 5480 3068
rect 5560 3176 5594 3210
rect 5656 3034 5690 3068
rect 5770 3176 5804 3210
rect 5866 3034 5900 3068
rect -2162 2950 -2128 2984
rect -1742 2950 -1708 2984
rect -1322 2950 -1288 2984
rect -902 2950 -868 2984
rect -482 2950 -448 2984
rect -62 2950 -28 2984
rect 358 2950 392 2984
rect 778 2950 812 2984
rect 1198 2950 1232 2984
rect 1618 2950 1652 2984
rect 2038 2950 2072 2984
rect 2458 2950 2492 2984
rect 2878 2950 2912 2984
rect 3298 2950 3332 2984
rect 3718 2950 3752 2984
rect 4138 2950 4172 2984
rect 4558 2950 4592 2984
rect 4978 2950 5012 2984
rect 5398 2950 5432 2984
rect 5818 2950 5852 2984
rect -2372 2820 -2338 2854
rect -1952 2820 -1918 2854
rect -1532 2820 -1498 2854
rect -1112 2820 -1078 2854
rect -692 2820 -658 2854
rect -272 2820 -238 2854
rect 148 2820 182 2854
rect 568 2820 602 2854
rect 988 2820 1022 2854
rect 1408 2820 1442 2854
rect 1828 2820 1862 2854
rect 2248 2820 2282 2854
rect 2668 2820 2702 2854
rect 3088 2820 3122 2854
rect 3508 2820 3542 2854
rect 3928 2820 3962 2854
rect 4348 2820 4382 2854
rect 4768 2820 4802 2854
rect 5188 2820 5222 2854
rect 5608 2820 5642 2854
rect -2420 2736 -2386 2770
rect -2324 2594 -2290 2628
rect -2210 2736 -2176 2770
rect -2114 2594 -2080 2628
rect -2000 2736 -1966 2770
rect -1904 2594 -1870 2628
rect -1790 2736 -1756 2770
rect -1694 2594 -1660 2628
rect -1580 2736 -1546 2770
rect -1484 2594 -1450 2628
rect -1370 2736 -1336 2770
rect -1274 2594 -1240 2628
rect -1160 2736 -1126 2770
rect -1064 2594 -1030 2628
rect -950 2736 -916 2770
rect -854 2594 -820 2628
rect -740 2736 -706 2770
rect -644 2594 -610 2628
rect -530 2736 -496 2770
rect -434 2594 -400 2628
rect -320 2736 -286 2770
rect -224 2594 -190 2628
rect -110 2736 -76 2770
rect -14 2594 20 2628
rect 100 2736 134 2770
rect 196 2594 230 2628
rect 310 2736 344 2770
rect 406 2594 440 2628
rect 520 2736 554 2770
rect 616 2594 650 2628
rect 730 2736 764 2770
rect 826 2594 860 2628
rect 940 2736 974 2770
rect 1036 2594 1070 2628
rect 1150 2736 1184 2770
rect 1246 2594 1280 2628
rect 1360 2736 1394 2770
rect 1456 2594 1490 2628
rect 1570 2736 1604 2770
rect 1666 2594 1700 2628
rect 1780 2736 1814 2770
rect 1876 2594 1910 2628
rect 1990 2736 2024 2770
rect 2086 2594 2120 2628
rect 2200 2736 2234 2770
rect 2296 2594 2330 2628
rect 2410 2736 2444 2770
rect 2506 2594 2540 2628
rect 2620 2736 2654 2770
rect 2716 2594 2750 2628
rect 2830 2736 2864 2770
rect 2926 2594 2960 2628
rect 3040 2736 3074 2770
rect 3136 2594 3170 2628
rect 3250 2736 3284 2770
rect 3346 2594 3380 2628
rect 3460 2736 3494 2770
rect 3556 2594 3590 2628
rect 3670 2736 3704 2770
rect 3766 2594 3800 2628
rect 3880 2736 3914 2770
rect 3976 2594 4010 2628
rect 4090 2736 4124 2770
rect 4186 2594 4220 2628
rect 4300 2736 4334 2770
rect 4396 2594 4430 2628
rect 4510 2736 4544 2770
rect 4606 2594 4640 2628
rect 4720 2736 4754 2770
rect 4816 2594 4850 2628
rect 4930 2736 4964 2770
rect 5026 2594 5060 2628
rect 5140 2736 5174 2770
rect 5236 2594 5270 2628
rect 5350 2736 5384 2770
rect 5446 2594 5480 2628
rect 5560 2736 5594 2770
rect 5656 2594 5690 2628
rect 5770 2736 5804 2770
rect 5866 2594 5900 2628
rect -2162 2510 -2128 2544
rect -1742 2510 -1708 2544
rect -1322 2510 -1288 2544
rect -902 2510 -868 2544
rect -482 2510 -448 2544
rect -62 2510 -28 2544
rect 358 2510 392 2544
rect 778 2510 812 2544
rect 1198 2510 1232 2544
rect 1618 2510 1652 2544
rect 2038 2510 2072 2544
rect 2458 2510 2492 2544
rect 2878 2510 2912 2544
rect 3298 2510 3332 2544
rect 3718 2510 3752 2544
rect 4138 2510 4172 2544
rect 4558 2510 4592 2544
rect 4978 2510 5012 2544
rect 5398 2510 5432 2544
rect 5818 2510 5852 2544
rect -2372 2380 -2338 2414
rect -1952 2380 -1918 2414
rect -1532 2380 -1498 2414
rect -1112 2380 -1078 2414
rect -692 2380 -658 2414
rect -272 2380 -238 2414
rect 148 2380 182 2414
rect 568 2380 602 2414
rect 988 2380 1022 2414
rect 1408 2380 1442 2414
rect 1828 2380 1862 2414
rect 2248 2380 2282 2414
rect 2668 2380 2702 2414
rect 3088 2380 3122 2414
rect 3508 2380 3542 2414
rect 3928 2380 3962 2414
rect 4348 2380 4382 2414
rect 4768 2380 4802 2414
rect 5188 2380 5222 2414
rect 5608 2380 5642 2414
rect -2420 2296 -2386 2330
rect -2324 2154 -2290 2188
rect -2210 2296 -2176 2330
rect -2114 2154 -2080 2188
rect -2000 2296 -1966 2330
rect -1904 2154 -1870 2188
rect -1790 2296 -1756 2330
rect -1694 2154 -1660 2188
rect -1580 2296 -1546 2330
rect -1484 2154 -1450 2188
rect -1370 2296 -1336 2330
rect -1274 2154 -1240 2188
rect -1160 2296 -1126 2330
rect -1064 2154 -1030 2188
rect -950 2296 -916 2330
rect -854 2154 -820 2188
rect -740 2296 -706 2330
rect -644 2154 -610 2188
rect -530 2296 -496 2330
rect -434 2154 -400 2188
rect -320 2296 -286 2330
rect -224 2154 -190 2188
rect -110 2296 -76 2330
rect -14 2154 20 2188
rect 100 2296 134 2330
rect 196 2154 230 2188
rect 310 2296 344 2330
rect 406 2154 440 2188
rect 520 2296 554 2330
rect 616 2154 650 2188
rect 730 2296 764 2330
rect 826 2154 860 2188
rect 940 2296 974 2330
rect 1036 2154 1070 2188
rect 1150 2296 1184 2330
rect 1246 2154 1280 2188
rect 1360 2296 1394 2330
rect 1456 2154 1490 2188
rect 1570 2296 1604 2330
rect 1666 2154 1700 2188
rect 1780 2296 1814 2330
rect 1876 2154 1910 2188
rect 1990 2296 2024 2330
rect 2086 2154 2120 2188
rect 2200 2296 2234 2330
rect 2296 2154 2330 2188
rect 2410 2296 2444 2330
rect 2506 2154 2540 2188
rect 2620 2296 2654 2330
rect 2716 2154 2750 2188
rect 2830 2296 2864 2330
rect 2926 2154 2960 2188
rect 3040 2296 3074 2330
rect 3136 2154 3170 2188
rect 3250 2296 3284 2330
rect 3346 2154 3380 2188
rect 3460 2296 3494 2330
rect 3556 2154 3590 2188
rect 3670 2296 3704 2330
rect 3766 2154 3800 2188
rect 3880 2296 3914 2330
rect 3976 2154 4010 2188
rect 4090 2296 4124 2330
rect 4186 2154 4220 2188
rect 4300 2296 4334 2330
rect 4396 2154 4430 2188
rect 4510 2296 4544 2330
rect 4606 2154 4640 2188
rect 4720 2296 4754 2330
rect 4816 2154 4850 2188
rect 4930 2296 4964 2330
rect 5026 2154 5060 2188
rect 5140 2296 5174 2330
rect 5236 2154 5270 2188
rect 5350 2296 5384 2330
rect 5446 2154 5480 2188
rect 5560 2296 5594 2330
rect 5656 2154 5690 2188
rect 5770 2296 5804 2330
rect 5866 2154 5900 2188
rect -2162 2070 -2128 2104
rect -1742 2070 -1708 2104
rect -1322 2070 -1288 2104
rect -902 2070 -868 2104
rect -482 2070 -448 2104
rect -62 2070 -28 2104
rect 358 2070 392 2104
rect 778 2070 812 2104
rect 1198 2070 1232 2104
rect 1618 2070 1652 2104
rect 2038 2070 2072 2104
rect 2458 2070 2492 2104
rect 2878 2070 2912 2104
rect 3298 2070 3332 2104
rect 3718 2070 3752 2104
rect 4138 2070 4172 2104
rect 4558 2070 4592 2104
rect 4978 2070 5012 2104
rect 5398 2070 5432 2104
rect 5818 2070 5852 2104
rect -2372 1940 -2338 1974
rect -1952 1940 -1918 1974
rect -1532 1940 -1498 1974
rect -1112 1940 -1078 1974
rect -692 1940 -658 1974
rect -272 1940 -238 1974
rect 148 1940 182 1974
rect 568 1940 602 1974
rect 988 1940 1022 1974
rect 1408 1940 1442 1974
rect 1828 1940 1862 1974
rect 2248 1940 2282 1974
rect 2668 1940 2702 1974
rect 3088 1940 3122 1974
rect 3508 1940 3542 1974
rect 3928 1940 3962 1974
rect 4348 1940 4382 1974
rect 4768 1940 4802 1974
rect 5188 1940 5222 1974
rect 5608 1940 5642 1974
rect -2420 1856 -2386 1890
rect -2324 1714 -2290 1748
rect -2210 1856 -2176 1890
rect -2114 1714 -2080 1748
rect -2000 1856 -1966 1890
rect -1904 1714 -1870 1748
rect -1790 1856 -1756 1890
rect -1694 1714 -1660 1748
rect -1580 1856 -1546 1890
rect -1484 1714 -1450 1748
rect -1370 1856 -1336 1890
rect -1274 1714 -1240 1748
rect -1160 1856 -1126 1890
rect -1064 1714 -1030 1748
rect -950 1856 -916 1890
rect -854 1714 -820 1748
rect -740 1856 -706 1890
rect -644 1714 -610 1748
rect -530 1856 -496 1890
rect -434 1714 -400 1748
rect -320 1856 -286 1890
rect -224 1714 -190 1748
rect -110 1856 -76 1890
rect -14 1714 20 1748
rect 100 1856 134 1890
rect 196 1714 230 1748
rect 310 1856 344 1890
rect 406 1714 440 1748
rect 520 1856 554 1890
rect 616 1714 650 1748
rect 730 1856 764 1890
rect 826 1714 860 1748
rect 940 1856 974 1890
rect 1036 1714 1070 1748
rect 1150 1856 1184 1890
rect 1246 1714 1280 1748
rect 1360 1856 1394 1890
rect 1456 1714 1490 1748
rect 1570 1856 1604 1890
rect 1666 1714 1700 1748
rect 1780 1856 1814 1890
rect 1876 1714 1910 1748
rect 1990 1856 2024 1890
rect 2086 1714 2120 1748
rect 2200 1856 2234 1890
rect 2296 1714 2330 1748
rect 2410 1856 2444 1890
rect 2506 1714 2540 1748
rect 2620 1856 2654 1890
rect 2716 1714 2750 1748
rect 2830 1856 2864 1890
rect 2926 1714 2960 1748
rect 3040 1856 3074 1890
rect 3136 1714 3170 1748
rect 3250 1856 3284 1890
rect 3346 1714 3380 1748
rect 3460 1856 3494 1890
rect 3556 1714 3590 1748
rect 3670 1856 3704 1890
rect 3766 1714 3800 1748
rect 3880 1856 3914 1890
rect 3976 1714 4010 1748
rect 4090 1856 4124 1890
rect 4186 1714 4220 1748
rect 4300 1856 4334 1890
rect 4396 1714 4430 1748
rect 4510 1856 4544 1890
rect 4606 1714 4640 1748
rect 4720 1856 4754 1890
rect 4816 1714 4850 1748
rect 4930 1856 4964 1890
rect 5026 1714 5060 1748
rect 5140 1856 5174 1890
rect 5236 1714 5270 1748
rect 5350 1856 5384 1890
rect 5446 1714 5480 1748
rect 5560 1856 5594 1890
rect 5656 1714 5690 1748
rect 5770 1856 5804 1890
rect 5866 1714 5900 1748
rect -2162 1630 -2128 1664
rect -1742 1630 -1708 1664
rect -1322 1630 -1288 1664
rect -902 1630 -868 1664
rect -482 1630 -448 1664
rect -62 1630 -28 1664
rect 358 1630 392 1664
rect 778 1630 812 1664
rect 1198 1630 1232 1664
rect 1618 1630 1652 1664
rect 2038 1630 2072 1664
rect 2458 1630 2492 1664
rect 2878 1630 2912 1664
rect 3298 1630 3332 1664
rect 3718 1630 3752 1664
rect 4138 1630 4172 1664
rect 4558 1630 4592 1664
rect 4978 1630 5012 1664
rect 5398 1630 5432 1664
rect 5818 1630 5852 1664
rect -2372 1500 -2338 1534
rect -1952 1500 -1918 1534
rect -1532 1500 -1498 1534
rect -1112 1500 -1078 1534
rect -692 1500 -658 1534
rect -272 1500 -238 1534
rect 148 1500 182 1534
rect 568 1500 602 1534
rect 988 1500 1022 1534
rect 1408 1500 1442 1534
rect 1828 1500 1862 1534
rect 2248 1500 2282 1534
rect 2668 1500 2702 1534
rect 3088 1500 3122 1534
rect 3508 1500 3542 1534
rect 3928 1500 3962 1534
rect 4348 1500 4382 1534
rect 4768 1500 4802 1534
rect 5188 1500 5222 1534
rect 5608 1500 5642 1534
rect -2420 1416 -2386 1450
rect -2324 1274 -2290 1308
rect -2210 1416 -2176 1450
rect -2114 1274 -2080 1308
rect -2000 1416 -1966 1450
rect -1904 1274 -1870 1308
rect -1790 1416 -1756 1450
rect -1694 1274 -1660 1308
rect -1580 1416 -1546 1450
rect -1484 1274 -1450 1308
rect -1370 1416 -1336 1450
rect -1274 1274 -1240 1308
rect -1160 1416 -1126 1450
rect -1064 1274 -1030 1308
rect -950 1416 -916 1450
rect -854 1274 -820 1308
rect -740 1416 -706 1450
rect -644 1274 -610 1308
rect -530 1416 -496 1450
rect -434 1274 -400 1308
rect -320 1416 -286 1450
rect -224 1274 -190 1308
rect -110 1416 -76 1450
rect -14 1274 20 1308
rect 100 1416 134 1450
rect 196 1274 230 1308
rect 310 1416 344 1450
rect 406 1274 440 1308
rect 520 1416 554 1450
rect 616 1274 650 1308
rect 730 1416 764 1450
rect 826 1274 860 1308
rect 940 1416 974 1450
rect 1036 1274 1070 1308
rect 1150 1416 1184 1450
rect 1246 1274 1280 1308
rect 1360 1416 1394 1450
rect 1456 1274 1490 1308
rect 1570 1416 1604 1450
rect 1666 1274 1700 1308
rect 1780 1416 1814 1450
rect 1876 1274 1910 1308
rect 1990 1416 2024 1450
rect 2086 1274 2120 1308
rect 2200 1416 2234 1450
rect 2296 1274 2330 1308
rect 2410 1416 2444 1450
rect 2506 1274 2540 1308
rect 2620 1416 2654 1450
rect 2716 1274 2750 1308
rect 2830 1416 2864 1450
rect 2926 1274 2960 1308
rect 3040 1416 3074 1450
rect 3136 1274 3170 1308
rect 3250 1416 3284 1450
rect 3346 1274 3380 1308
rect 3460 1416 3494 1450
rect 3556 1274 3590 1308
rect 3670 1416 3704 1450
rect 3766 1274 3800 1308
rect 3880 1416 3914 1450
rect 3976 1274 4010 1308
rect 4090 1416 4124 1450
rect 4186 1274 4220 1308
rect 4300 1416 4334 1450
rect 4396 1274 4430 1308
rect 4510 1416 4544 1450
rect 4606 1274 4640 1308
rect 4720 1416 4754 1450
rect 4816 1274 4850 1308
rect 4930 1416 4964 1450
rect 5026 1274 5060 1308
rect 5140 1416 5174 1450
rect 5236 1274 5270 1308
rect 5350 1416 5384 1450
rect 5446 1274 5480 1308
rect 5560 1416 5594 1450
rect 5656 1274 5690 1308
rect 5770 1416 5804 1450
rect 5866 1274 5900 1308
rect -2162 1190 -2128 1224
rect -1742 1190 -1708 1224
rect -1322 1190 -1288 1224
rect -902 1190 -868 1224
rect -482 1190 -448 1224
rect -62 1190 -28 1224
rect 358 1190 392 1224
rect 778 1190 812 1224
rect 1198 1190 1232 1224
rect 1618 1190 1652 1224
rect 2038 1190 2072 1224
rect 2458 1190 2492 1224
rect 2878 1190 2912 1224
rect 3298 1190 3332 1224
rect 3718 1190 3752 1224
rect 4138 1190 4172 1224
rect 4558 1190 4592 1224
rect 4978 1190 5012 1224
rect 5398 1190 5432 1224
rect 5818 1190 5852 1224
rect -2372 1060 -2338 1094
rect -1952 1060 -1918 1094
rect -1532 1060 -1498 1094
rect -1112 1060 -1078 1094
rect -692 1060 -658 1094
rect -272 1060 -238 1094
rect 148 1060 182 1094
rect 568 1060 602 1094
rect 988 1060 1022 1094
rect 1408 1060 1442 1094
rect 1828 1060 1862 1094
rect 2248 1060 2282 1094
rect 2668 1060 2702 1094
rect 3088 1060 3122 1094
rect 3508 1060 3542 1094
rect 3928 1060 3962 1094
rect 4348 1060 4382 1094
rect 4768 1060 4802 1094
rect 5188 1060 5222 1094
rect 5608 1060 5642 1094
rect -2420 976 -2386 1010
rect -2324 834 -2290 868
rect -2210 976 -2176 1010
rect -2114 834 -2080 868
rect -2000 976 -1966 1010
rect -1904 834 -1870 868
rect -1790 976 -1756 1010
rect -1694 834 -1660 868
rect -1580 976 -1546 1010
rect -1484 834 -1450 868
rect -1370 976 -1336 1010
rect -1274 834 -1240 868
rect -1160 976 -1126 1010
rect -1064 834 -1030 868
rect -950 976 -916 1010
rect -854 834 -820 868
rect -740 976 -706 1010
rect -644 834 -610 868
rect -530 976 -496 1010
rect -434 834 -400 868
rect -320 976 -286 1010
rect -224 834 -190 868
rect -110 976 -76 1010
rect -14 834 20 868
rect 100 976 134 1010
rect 196 834 230 868
rect 310 976 344 1010
rect 406 834 440 868
rect 520 976 554 1010
rect 616 834 650 868
rect 730 976 764 1010
rect 826 834 860 868
rect 940 976 974 1010
rect 1036 834 1070 868
rect 1150 976 1184 1010
rect 1246 834 1280 868
rect 1360 976 1394 1010
rect 1456 834 1490 868
rect 1570 976 1604 1010
rect 1666 834 1700 868
rect 1780 976 1814 1010
rect 1876 834 1910 868
rect 1990 976 2024 1010
rect 2086 834 2120 868
rect 2200 976 2234 1010
rect 2296 834 2330 868
rect 2410 976 2444 1010
rect 2506 834 2540 868
rect 2620 976 2654 1010
rect 2716 834 2750 868
rect 2830 976 2864 1010
rect 2926 834 2960 868
rect 3040 976 3074 1010
rect 3136 834 3170 868
rect 3250 976 3284 1010
rect 3346 834 3380 868
rect 3460 976 3494 1010
rect 3556 834 3590 868
rect 3670 976 3704 1010
rect 3766 834 3800 868
rect 3880 976 3914 1010
rect 3976 834 4010 868
rect 4090 976 4124 1010
rect 4186 834 4220 868
rect 4300 976 4334 1010
rect 4396 834 4430 868
rect 4510 976 4544 1010
rect 4606 834 4640 868
rect 4720 976 4754 1010
rect 4816 834 4850 868
rect 4930 976 4964 1010
rect 5026 834 5060 868
rect 5140 976 5174 1010
rect 5236 834 5270 868
rect 5350 976 5384 1010
rect 5446 834 5480 868
rect 5560 976 5594 1010
rect 5656 834 5690 868
rect 5770 976 5804 1010
rect 5866 834 5900 868
rect -2162 750 -2128 784
rect -1742 750 -1708 784
rect -1322 750 -1288 784
rect -902 750 -868 784
rect -482 750 -448 784
rect -62 750 -28 784
rect 358 750 392 784
rect 778 750 812 784
rect 1198 750 1232 784
rect 1618 750 1652 784
rect 2038 750 2072 784
rect 2458 750 2492 784
rect 2878 750 2912 784
rect 3298 750 3332 784
rect 3718 750 3752 784
rect 4138 750 4172 784
rect 4558 750 4592 784
rect 4978 750 5012 784
rect 5398 750 5432 784
rect 5818 750 5852 784
rect 6192 745 6226 4180
rect 6843 5370 6877 5403
rect 6843 5369 6877 5370
rect 6750 5322 6784 5356
rect 6985 5274 7019 5307
rect 6985 5273 7019 5274
rect 7078 5226 7112 5260
rect 6843 5178 6877 5211
rect 6843 5177 6877 5178
rect 6750 5130 6784 5164
rect 6985 5082 7019 5115
rect 6985 5081 7019 5082
rect 7078 5034 7112 5068
rect 6843 4986 6877 5019
rect 6843 4985 6877 4986
rect 6750 4938 6784 4972
rect 6985 4890 7019 4923
rect 6985 4889 7019 4890
rect 7078 4842 7112 4876
rect 6843 4794 6877 4827
rect 6843 4793 6877 4794
rect 6750 4746 6784 4780
rect 6985 4698 7019 4731
rect 6985 4697 7019 4698
rect 7078 4650 7112 4684
rect 6843 4602 6877 4635
rect 6843 4601 6877 4602
rect 6750 4554 6784 4588
rect 6985 4506 7019 4539
rect 6985 4505 7019 4506
rect 7078 4458 7112 4492
rect 6843 4410 6877 4443
rect 6843 4409 6877 4410
rect 6750 4362 6784 4396
rect 6985 4314 7019 4347
rect 6985 4313 7019 4314
rect 7078 4266 7112 4300
rect 6843 4218 6877 4251
rect 6843 4217 6877 4218
rect 6750 4170 6784 4204
rect 6985 4122 7019 4155
rect 6985 4121 7019 4122
rect 7078 4074 7112 4108
rect 6843 4026 6877 4059
rect 6843 4025 6877 4026
rect 6750 3978 6784 4012
rect 6985 3930 7019 3963
rect 6985 3929 7019 3930
rect 7078 3882 7112 3916
rect 6843 3834 6877 3867
rect 6843 3833 6877 3834
rect 6744 3624 7118 3657
rect 6744 3623 7118 3624
rect 282 256 316 290
rect 474 256 508 290
rect 666 256 700 290
rect 858 256 892 290
rect 1050 256 1084 290
rect 1242 256 1276 290
rect 1434 256 1468 290
rect 1626 256 1660 290
rect 1818 256 1852 290
rect 2010 256 2044 290
rect 2202 256 2236 290
rect 2394 256 2428 290
rect 2586 256 2620 290
rect 2778 256 2812 290
rect 2970 256 3004 290
rect 3162 256 3196 290
rect 186 171 220 205
rect 282 30 316 63
rect 282 29 316 30
rect 378 171 412 205
rect 474 30 508 63
rect 474 29 508 30
rect 570 171 604 205
rect 666 30 700 63
rect 666 29 700 30
rect 762 171 796 205
rect 858 30 892 63
rect 858 29 892 30
rect 954 171 988 205
rect 1050 30 1084 63
rect 1050 29 1084 30
rect 1146 171 1180 205
rect 1242 30 1276 63
rect 1242 29 1276 30
rect 1338 171 1372 205
rect 1434 30 1468 63
rect 1434 29 1468 30
rect 1530 171 1564 205
rect 1626 30 1660 63
rect 1626 29 1660 30
rect 1722 171 1756 205
rect 1818 30 1852 63
rect 1818 29 1852 30
rect 1914 171 1948 205
rect 2010 30 2044 63
rect 2010 29 2044 30
rect 2106 171 2140 205
rect 2202 30 2236 63
rect 2202 29 2236 30
rect 2298 171 2332 205
rect 2394 30 2428 63
rect 2394 29 2428 30
rect 2490 171 2524 205
rect 2586 30 2620 63
rect 2586 29 2620 30
rect 2682 171 2716 205
rect 2778 30 2812 63
rect 2778 29 2812 30
rect 2874 171 2908 205
rect 2970 30 3004 63
rect 2970 29 3004 30
rect 3066 171 3100 205
rect 3162 30 3196 63
rect 3162 29 3196 30
rect 3258 171 3292 205
rect 72 -156 3406 -123
rect 72 -157 3406 -156
<< metal1 >>
rect 1134 10604 1230 10729
rect 1134 10570 1165 10604
rect 1199 10570 1230 10604
rect 1134 10512 1230 10570
rect 1134 10478 1165 10512
rect 1199 10478 1230 10512
rect 1134 10420 1230 10478
rect 1134 10386 1165 10420
rect 1199 10386 1230 10420
rect 1134 10328 1230 10386
rect 1134 10294 1165 10328
rect 1199 10294 1230 10328
rect 1134 10236 1230 10294
rect 1134 10202 1165 10236
rect 1199 10202 1230 10236
rect 1134 10144 1230 10202
rect 1134 10110 1165 10144
rect 1199 10110 1230 10144
rect 1134 10052 1230 10110
rect 1134 10018 1165 10052
rect 1199 10018 1230 10052
rect 1134 9960 1230 10018
rect 1134 9926 1165 9960
rect 1199 9926 1230 9960
rect 1134 9868 1230 9926
rect 1134 9834 1165 9868
rect 1199 9834 1230 9868
rect 1134 9790 1230 9834
rect 1134 9738 1156 9790
rect 1208 9738 1230 9790
rect 1134 9684 1230 9738
rect 1134 9650 1165 9684
rect 1199 9650 1230 9684
rect 1134 9649 1230 9650
rect 1134 9597 1156 9649
rect 1208 9597 1230 9649
rect 1134 9592 1230 9597
rect 1134 9558 1165 9592
rect 1199 9558 1230 9592
rect 1134 9508 1230 9558
rect 1134 9456 1156 9508
rect 1208 9456 1230 9508
rect 1134 9408 1230 9456
rect 1134 9374 1165 9408
rect 1199 9374 1230 9408
rect 1134 9367 1230 9374
rect 1134 9315 1156 9367
rect 1208 9315 1230 9367
rect 1134 9282 1165 9315
rect 1199 9282 1230 9315
rect 1134 9226 1230 9282
rect 1134 9174 1156 9226
rect 1208 9174 1230 9226
rect 1134 9132 1230 9174
rect 1134 9098 1165 9132
rect 1199 9098 1230 9132
rect 1134 9040 1230 9098
rect 1134 9006 1165 9040
rect 1199 9006 1230 9040
rect 1134 8948 1230 9006
rect 1317 8995 1351 10729
rect 1678 10604 1774 10729
rect 1678 10570 1709 10604
rect 1743 10570 1774 10604
rect 1678 10512 1774 10570
rect 1678 10478 1709 10512
rect 1743 10478 1774 10512
rect 1678 10420 1774 10478
rect 1678 10386 1709 10420
rect 1743 10386 1774 10420
rect 1678 10328 1774 10386
rect 1678 10294 1709 10328
rect 1743 10294 1774 10328
rect 1678 10236 1774 10294
rect 1678 10202 1709 10236
rect 1743 10202 1774 10236
rect 1678 10144 1774 10202
rect 1678 10110 1709 10144
rect 1743 10110 1774 10144
rect 1678 10052 1774 10110
rect 1678 10018 1709 10052
rect 1743 10018 1774 10052
rect 1678 9960 1774 10018
rect 1678 9926 1709 9960
rect 1743 9926 1774 9960
rect 1678 9868 1774 9926
rect 1678 9834 1709 9868
rect 1743 9834 1774 9868
rect 1678 9776 1774 9834
rect 1678 9742 1709 9776
rect 1743 9742 1774 9776
rect 1678 9684 1774 9742
rect 1678 9650 1709 9684
rect 1743 9650 1774 9684
rect 1678 9592 1774 9650
rect 1678 9558 1709 9592
rect 1743 9558 1774 9592
rect 1678 9500 1774 9558
rect 1678 9466 1709 9500
rect 1743 9466 1774 9500
rect 1678 9408 1774 9466
rect 1678 9374 1709 9408
rect 1743 9374 1774 9408
rect 1397 9362 1449 9374
rect 1392 9356 1450 9362
rect 1392 9322 1404 9356
rect 1438 9322 1450 9356
rect 1392 9316 1450 9322
rect 1397 9271 1449 9316
rect 1392 9265 1450 9271
rect 1566 9268 1576 9320
rect 1628 9268 1638 9320
rect 1678 9316 1774 9374
rect 1993 9320 2003 9372
rect 2055 9320 2065 9372
rect 1678 9282 1709 9316
rect 1743 9282 1774 9316
rect 1392 9231 1404 9265
rect 1438 9231 1450 9265
rect 1392 9225 1450 9231
rect 1397 9154 1449 9225
rect 1387 9102 1397 9154
rect 1449 9102 1459 9154
rect 1305 8989 1363 8995
rect 1391 8989 1449 8995
rect 1576 8991 1628 9268
rect 1678 9224 1774 9282
rect 2003 9268 2055 9320
rect 1678 9190 1709 9224
rect 1743 9190 1774 9224
rect 1993 9216 2003 9268
rect 2055 9216 2065 9268
rect 1678 9132 1774 9190
rect 1678 9098 1709 9132
rect 1743 9098 1774 9132
rect 1813 9102 1823 9154
rect 1875 9102 1885 9154
rect 1678 9040 1774 9098
rect 1678 9006 1709 9040
rect 1743 9006 1774 9040
rect 1305 8955 1317 8989
rect 1351 8955 1403 8989
rect 1437 8955 1449 8989
rect 1305 8949 1363 8955
rect 1391 8949 1449 8955
rect 1134 8914 1165 8948
rect 1199 8914 1230 8948
rect 1477 8939 1487 8991
rect 1539 8939 1576 8991
rect 1628 8988 1638 8991
rect 1628 8982 1645 8988
rect 1633 8948 1645 8982
rect 1628 8942 1645 8948
rect 1678 8948 1774 9006
rect 1823 8991 1875 9102
rect 2102 8995 2136 10729
rect 2222 10604 2318 10729
rect 2222 10570 2253 10604
rect 2287 10570 2318 10604
rect 2222 10512 2318 10570
rect 2222 10478 2253 10512
rect 2287 10478 2318 10512
rect 2222 10420 2318 10478
rect 2222 10386 2253 10420
rect 2287 10386 2318 10420
rect 2222 10328 2318 10386
rect 2222 10294 2253 10328
rect 2287 10294 2318 10328
rect 2222 10236 2318 10294
rect 2222 10202 2253 10236
rect 2287 10202 2318 10236
rect 2222 10144 2318 10202
rect 2222 10110 2253 10144
rect 2287 10110 2318 10144
rect 2222 10052 2318 10110
rect 2222 10018 2253 10052
rect 2287 10018 2318 10052
rect 2222 9960 2318 10018
rect 2222 9926 2253 9960
rect 2287 9926 2318 9960
rect 2222 9868 2318 9926
rect 2222 9834 2253 9868
rect 2287 9834 2318 9868
rect 2222 9792 2318 9834
rect 2222 9740 2244 9792
rect 2296 9740 2318 9792
rect 2222 9684 2318 9740
rect 2222 9651 2253 9684
rect 2287 9651 2318 9684
rect 2222 9599 2244 9651
rect 2296 9599 2318 9651
rect 2222 9592 2318 9599
rect 2222 9558 2253 9592
rect 2287 9558 2318 9592
rect 2222 9510 2318 9558
rect 2222 9458 2244 9510
rect 2296 9458 2318 9510
rect 2222 9408 2318 9458
rect 2222 9374 2253 9408
rect 2287 9374 2318 9408
rect 2222 9369 2318 9374
rect 2222 9317 2244 9369
rect 2296 9317 2318 9369
rect 2222 9316 2318 9317
rect 2222 9282 2253 9316
rect 2287 9282 2318 9316
rect 2222 9228 2318 9282
rect 2222 9176 2244 9228
rect 2296 9176 2318 9228
rect 2222 9132 2318 9176
rect 2222 9098 2253 9132
rect 2287 9098 2318 9132
rect 2222 9040 2318 9098
rect 2222 9006 2253 9040
rect 2287 9006 2318 9040
rect 1813 8988 1823 8991
rect 1628 8939 1638 8942
rect 1134 8856 1230 8914
rect 1134 8822 1165 8856
rect 1199 8822 1230 8856
rect 1134 8764 1230 8822
rect 1678 8914 1709 8948
rect 1743 8914 1774 8948
rect 1808 8982 1823 8988
rect 1808 8948 1820 8982
rect 1808 8942 1823 8948
rect 1813 8939 1823 8942
rect 1875 8939 1912 8991
rect 1964 8939 1974 8991
rect 2004 8989 2148 8995
rect 2004 8955 2016 8989
rect 2050 8955 2102 8989
rect 2136 8955 2148 8989
rect 2004 8949 2148 8955
rect 2222 8948 2318 9006
rect 1678 8856 1774 8914
rect 1678 8822 1709 8856
rect 1743 8822 1774 8856
rect 1134 8730 1165 8764
rect 1199 8730 1230 8764
rect 1392 8780 1450 8786
rect 1392 8746 1404 8780
rect 1438 8746 1450 8780
rect 1392 8740 1450 8746
rect 1678 8764 1774 8822
rect 2222 8914 2253 8948
rect 2287 8914 2318 8948
rect 2222 8856 2318 8914
rect 2222 8822 2253 8856
rect 2287 8822 2318 8856
rect 1134 8672 1230 8730
rect 1403 8700 1438 8740
rect 1678 8730 1709 8764
rect 1743 8730 1774 8764
rect 2000 8779 2058 8785
rect 2000 8745 2012 8779
rect 2046 8745 2058 8779
rect 2000 8739 2058 8745
rect 2222 8764 2318 8822
rect 1134 8638 1165 8672
rect 1199 8638 1230 8672
rect 1392 8694 1450 8700
rect 1392 8660 1404 8694
rect 1438 8660 1450 8694
rect 1392 8654 1450 8660
rect 1678 8672 1774 8730
rect 2012 8699 2047 8739
rect 2222 8730 2253 8764
rect 2287 8730 2318 8764
rect 1134 8580 1230 8638
rect 1134 8546 1165 8580
rect 1199 8546 1230 8580
rect 1134 8488 1230 8546
rect 1403 8505 1438 8654
rect 1678 8638 1709 8672
rect 1743 8638 1774 8672
rect 2000 8693 2058 8699
rect 2000 8659 2012 8693
rect 2046 8659 2058 8693
rect 2000 8653 2058 8659
rect 2222 8672 2318 8730
rect 1678 8580 1774 8638
rect 1678 8546 1709 8580
rect 1743 8546 1774 8580
rect 1134 8454 1165 8488
rect 1199 8454 1230 8488
rect 1294 8498 1564 8505
rect 1294 8463 1306 8498
rect 1341 8497 1564 8498
rect 1341 8470 1518 8497
rect 1341 8463 1353 8470
rect 1294 8457 1353 8463
rect 1506 8463 1518 8470
rect 1552 8463 1564 8497
rect 1506 8457 1564 8463
rect 1678 8488 1774 8546
rect 2012 8504 2047 8653
rect 2222 8638 2253 8672
rect 2287 8638 2318 8672
rect 2222 8580 2318 8638
rect 2222 8546 2253 8580
rect 2287 8546 2318 8580
rect 1134 8396 1230 8454
rect 1134 8362 1165 8396
rect 1199 8362 1230 8396
rect 1134 8304 1230 8362
rect 1678 8454 1709 8488
rect 1743 8454 1774 8488
rect 1886 8497 2156 8504
rect 1886 8496 2109 8497
rect 1886 8462 1898 8496
rect 1932 8469 2109 8496
rect 1932 8462 1944 8469
rect 1886 8456 1944 8462
rect 2097 8462 2109 8469
rect 2144 8462 2156 8497
rect 2097 8456 2156 8462
rect 2222 8488 2318 8546
rect 1678 8396 1774 8454
rect 1678 8362 1709 8396
rect 1743 8362 1774 8396
rect 1134 8270 1165 8304
rect 1199 8270 1230 8304
rect 1379 8270 1389 8322
rect 1441 8270 1451 8322
rect 1678 8304 1774 8362
rect 2222 8454 2253 8488
rect 2287 8454 2318 8488
rect 2222 8396 2318 8454
rect 2222 8362 2253 8396
rect 2287 8362 2318 8396
rect 1678 8270 1709 8304
rect 1743 8270 1774 8304
rect 2003 8271 2013 8323
rect 2065 8271 2075 8323
rect 2222 8304 2318 8362
rect 1134 8241 1230 8270
rect 1678 8131 1774 8270
rect 2222 8270 2253 8304
rect 2287 8270 2318 8304
rect 2222 8241 2318 8270
rect -3788 8041 7250 8131
rect -3788 8023 -1286 8041
rect -1234 8023 287 8041
rect 339 8023 3230 8041
rect 3282 8023 4699 8041
rect 4751 8023 7250 8041
rect -3788 7989 -3656 8023
rect -3282 7989 -2662 8023
rect 6114 7989 6744 8023
rect 7118 7989 7250 8023
rect -3788 7983 7250 7989
rect -3557 7723 -3523 7983
rect -3427 7813 -3369 7819
rect -3427 7779 -3415 7813
rect -3381 7779 -3369 7813
rect -3427 7773 -3369 7779
rect -3322 7778 -3288 7781
rect -3569 7717 -3511 7723
rect -3650 7682 -3616 7685
rect -3569 7683 -3557 7717
rect -3523 7683 -3511 7717
rect -3656 7670 -3610 7682
rect -3569 7677 -3511 7683
rect -3656 7636 -3650 7670
rect -3616 7636 -3610 7670
rect -3656 7624 -3610 7636
rect -3650 7581 -3616 7624
rect -3672 7529 -3662 7581
rect -3610 7529 -3600 7581
rect -3557 7531 -3523 7677
rect -3415 7627 -3381 7773
rect -3328 7766 -3282 7778
rect -3328 7732 -3322 7766
rect -3288 7732 -3282 7766
rect -3328 7720 -3282 7732
rect -3427 7621 -3369 7627
rect -3427 7587 -3415 7621
rect -3381 7587 -3369 7621
rect -3427 7581 -3369 7587
rect -3322 7586 -3288 7720
rect -3328 7581 -3282 7586
rect -3650 7490 -3616 7529
rect -3569 7525 -3511 7531
rect -3569 7491 -3557 7525
rect -3523 7491 -3511 7525
rect -3656 7478 -3610 7490
rect -3569 7485 -3511 7491
rect -3656 7444 -3650 7478
rect -3616 7444 -3610 7478
rect -3656 7432 -3610 7444
rect -3650 7298 -3616 7432
rect -3557 7339 -3523 7485
rect -3415 7435 -3381 7581
rect -3341 7529 -3331 7581
rect -3279 7529 -3269 7581
rect -3328 7528 -3282 7529
rect -3427 7429 -3369 7435
rect -3427 7395 -3415 7429
rect -3381 7395 -3369 7429
rect -3427 7389 -3369 7395
rect -3322 7394 -3288 7528
rect -3569 7333 -3511 7339
rect -3569 7299 -3557 7333
rect -3523 7299 -3511 7333
rect -3656 7286 -3610 7298
rect -3569 7293 -3511 7299
rect -3656 7252 -3650 7286
rect -3616 7252 -3610 7286
rect -3656 7240 -3610 7252
rect -3650 7106 -3616 7240
rect -3557 7147 -3523 7293
rect -3415 7243 -3381 7389
rect -3328 7382 -3282 7394
rect -3328 7348 -3322 7382
rect -3288 7348 -3282 7382
rect -3328 7336 -3282 7348
rect -3427 7237 -3369 7243
rect -3427 7203 -3415 7237
rect -3381 7203 -3369 7237
rect -3427 7197 -3369 7203
rect -3322 7202 -3288 7336
rect -3569 7141 -3511 7147
rect -3569 7107 -3557 7141
rect -3523 7107 -3511 7141
rect -3656 7094 -3610 7106
rect -3569 7101 -3511 7107
rect -3656 7060 -3650 7094
rect -3616 7060 -3610 7094
rect -3656 7048 -3610 7060
rect -3650 6914 -3616 7048
rect -3557 6955 -3523 7101
rect -3415 7051 -3381 7197
rect -3328 7190 -3282 7202
rect -3328 7156 -3322 7190
rect -3288 7156 -3282 7190
rect -3328 7144 -3282 7156
rect -3427 7045 -3369 7051
rect -3427 7011 -3415 7045
rect -3381 7011 -3369 7045
rect -3427 7005 -3369 7011
rect -3322 7010 -3288 7144
rect -3569 6949 -3511 6955
rect -3569 6915 -3557 6949
rect -3523 6915 -3511 6949
rect -3656 6902 -3610 6914
rect -3569 6909 -3511 6915
rect -3656 6868 -3650 6902
rect -3616 6868 -3610 6902
rect -3656 6856 -3610 6868
rect -3650 6722 -3616 6856
rect -3557 6763 -3523 6909
rect -3415 6859 -3381 7005
rect -3328 6998 -3282 7010
rect -3328 6964 -3322 6998
rect -3288 6964 -3282 6998
rect -3328 6952 -3282 6964
rect -3427 6853 -3369 6859
rect -3427 6819 -3415 6853
rect -3381 6819 -3369 6853
rect -3427 6813 -3369 6819
rect -3322 6818 -3288 6952
rect -3569 6757 -3511 6763
rect -3569 6723 -3557 6757
rect -3523 6723 -3511 6757
rect -3656 6710 -3610 6722
rect -3569 6717 -3511 6723
rect -3415 6720 -3381 6813
rect -3328 6806 -3282 6818
rect -3328 6772 -3322 6806
rect -3288 6772 -3282 6806
rect -3328 6760 -3282 6772
rect -3656 6676 -3650 6710
rect -3616 6676 -3610 6710
rect -3656 6664 -3610 6676
rect -3650 6530 -3616 6664
rect -3557 6571 -3523 6717
rect -3433 6668 -3423 6720
rect -3371 6668 -3361 6720
rect -3427 6661 -3369 6668
rect -3427 6627 -3415 6661
rect -3381 6627 -3369 6661
rect -3427 6621 -3369 6627
rect -3322 6626 -3288 6760
rect -3569 6565 -3511 6571
rect -3569 6531 -3557 6565
rect -3523 6531 -3511 6565
rect -3656 6518 -3610 6530
rect -3569 6525 -3511 6531
rect -3656 6484 -3650 6518
rect -3616 6484 -3610 6518
rect -3656 6472 -3610 6484
rect -3650 6431 -3616 6472
rect -3670 6379 -3660 6431
rect -3608 6379 -3598 6431
rect -3557 6379 -3523 6525
rect -3415 6475 -3381 6621
rect -3328 6614 -3282 6626
rect -3328 6580 -3322 6614
rect -3288 6580 -3282 6614
rect -3328 6568 -3282 6580
rect -3427 6469 -3369 6475
rect -3427 6435 -3415 6469
rect -3381 6435 -3369 6469
rect -3427 6429 -3369 6435
rect -3322 6434 -3288 6568
rect -3328 6431 -3282 6434
rect -3650 6338 -3616 6379
rect -3569 6373 -3511 6379
rect -3569 6339 -3557 6373
rect -3523 6339 -3511 6373
rect -3656 6326 -3610 6338
rect -3569 6333 -3511 6339
rect -3656 6292 -3650 6326
rect -3616 6292 -3610 6326
rect -3656 6280 -3610 6292
rect -3650 6275 -3616 6280
rect -3557 6073 -3523 6333
rect -3415 6283 -3381 6429
rect -3341 6379 -3331 6431
rect -3279 6379 -3269 6431
rect -3328 6376 -3282 6379
rect -3322 6371 -3288 6376
rect -3427 6277 -3369 6283
rect -3427 6243 -3415 6277
rect -3381 6243 -3369 6277
rect -3427 6237 -3369 6243
rect -3220 6073 -3150 7983
rect -2398 7921 -2340 7927
rect -1978 7921 -1920 7927
rect -1558 7921 -1500 7927
rect -1138 7921 -1080 7927
rect -718 7921 -660 7927
rect -298 7921 -240 7927
rect 122 7921 180 7927
rect 542 7921 600 7927
rect 962 7921 1020 7927
rect 1382 7921 1440 7927
rect 1802 7921 1860 7927
rect 1960 7921 1970 7930
rect -2446 7887 -2386 7921
rect -2352 7887 -1966 7921
rect -1932 7887 -1546 7921
rect -1512 7887 -1126 7921
rect -1092 7887 -706 7921
rect -672 7887 -286 7921
rect -252 7887 134 7921
rect 168 7887 554 7921
rect 588 7887 974 7921
rect 1008 7887 1394 7921
rect 1428 7887 1814 7921
rect 1848 7887 1970 7921
rect -2398 7881 -2340 7887
rect -1978 7881 -1920 7887
rect -1558 7881 -1500 7887
rect -1138 7881 -1080 7887
rect -718 7881 -660 7887
rect -298 7881 -240 7887
rect 122 7881 180 7887
rect 542 7881 600 7887
rect 962 7881 1020 7887
rect 1382 7881 1440 7887
rect 1802 7881 1860 7887
rect 1960 7878 1970 7887
rect 2022 7921 2032 7930
rect 2222 7921 2280 7927
rect 2642 7921 2700 7927
rect 3062 7921 3120 7927
rect 3482 7921 3540 7927
rect 3902 7921 3960 7927
rect 4322 7921 4380 7927
rect 4742 7921 4800 7927
rect 5162 7921 5220 7927
rect 5582 7921 5640 7927
rect 2022 7887 2234 7921
rect 2268 7887 2654 7921
rect 2688 7887 3074 7921
rect 3108 7887 3494 7921
rect 3528 7887 3914 7921
rect 3948 7887 4334 7921
rect 4368 7887 4754 7921
rect 4788 7887 5174 7921
rect 5208 7887 5594 7921
rect 5628 7887 5898 7921
rect 2022 7878 2032 7887
rect 2222 7881 2280 7887
rect 2642 7881 2700 7887
rect 3062 7881 3120 7887
rect 3482 7881 3540 7887
rect 3902 7881 3960 7887
rect 4322 7881 4380 7887
rect 4742 7881 4800 7887
rect 5162 7881 5220 7887
rect 5582 7881 5640 7887
rect -2446 7828 -2388 7834
rect -2236 7828 -2178 7834
rect -2026 7828 -1968 7834
rect -1816 7828 -1758 7834
rect -1606 7828 -1548 7834
rect -1396 7828 -1338 7834
rect -1186 7828 -1128 7834
rect -976 7828 -918 7834
rect -766 7828 -708 7834
rect -556 7828 -498 7834
rect -346 7828 -288 7834
rect -136 7828 -78 7834
rect 74 7828 132 7834
rect 284 7828 342 7834
rect 494 7828 552 7834
rect 704 7828 762 7834
rect 914 7828 972 7834
rect 1124 7828 1182 7834
rect 1334 7828 1392 7834
rect 1544 7828 1602 7834
rect 1754 7828 1812 7834
rect 1964 7828 2022 7834
rect 2174 7828 2232 7834
rect 2384 7828 2442 7834
rect 2594 7828 2652 7834
rect 2804 7828 2862 7834
rect 3014 7828 3072 7834
rect 3224 7828 3282 7834
rect 3434 7828 3492 7834
rect 3644 7828 3702 7834
rect 3854 7828 3912 7834
rect 4064 7828 4122 7834
rect 4274 7828 4332 7834
rect 4484 7828 4542 7834
rect 4694 7828 4752 7834
rect 4904 7828 4962 7834
rect 5114 7828 5172 7834
rect 5324 7828 5382 7834
rect 5534 7828 5592 7834
rect 5744 7828 5802 7834
rect -2446 7794 -2434 7828
rect -2400 7794 -2224 7828
rect -2190 7794 -2014 7828
rect -1980 7794 -1804 7828
rect -1770 7794 -1594 7828
rect -1560 7794 -1384 7828
rect -1350 7794 -1286 7828
rect -2446 7788 -2388 7794
rect -2236 7788 -2178 7794
rect -2026 7788 -1968 7794
rect -1816 7788 -1758 7794
rect -1606 7788 -1548 7794
rect -1396 7788 -1338 7794
rect -1296 7776 -1286 7794
rect -1234 7794 -1174 7828
rect -1140 7794 -964 7828
rect -930 7794 -754 7828
rect -720 7794 -544 7828
rect -510 7794 -334 7828
rect -300 7794 -124 7828
rect -90 7794 86 7828
rect 120 7794 287 7828
rect 339 7794 506 7828
rect 540 7794 716 7828
rect 750 7794 926 7828
rect 960 7794 1136 7828
rect 1170 7794 1346 7828
rect 1380 7794 1556 7828
rect 1590 7794 1766 7828
rect 1800 7794 1976 7828
rect 2010 7794 2186 7828
rect 2220 7794 2396 7828
rect 2430 7794 2606 7828
rect 2640 7794 2816 7828
rect 2850 7794 3026 7828
rect 3060 7794 3230 7828
rect 3282 7794 3446 7828
rect 3480 7794 3656 7828
rect 3690 7794 3866 7828
rect 3900 7794 4076 7828
rect 4110 7794 4286 7828
rect 4320 7794 4496 7828
rect 4530 7794 4699 7828
rect 4751 7794 4916 7828
rect 4950 7794 5126 7828
rect 5160 7794 5336 7828
rect 5370 7794 5546 7828
rect 5580 7794 5756 7828
rect 5790 7794 5898 7828
rect -1234 7776 -1224 7794
rect -1186 7788 -1128 7794
rect -976 7788 -918 7794
rect -766 7788 -708 7794
rect -556 7788 -498 7794
rect -346 7788 -288 7794
rect -136 7788 -78 7794
rect 74 7788 132 7794
rect 277 7776 287 7794
rect 339 7776 349 7794
rect 494 7788 552 7794
rect 704 7788 762 7794
rect 914 7788 972 7794
rect 1124 7788 1182 7794
rect 1334 7788 1392 7794
rect 1544 7788 1602 7794
rect 1749 7776 1821 7794
rect 1964 7788 2022 7794
rect 2174 7788 2232 7794
rect 2384 7788 2442 7794
rect 2594 7788 2652 7794
rect 2804 7788 2862 7794
rect 3014 7788 3072 7794
rect 3220 7776 3230 7794
rect 3282 7776 3292 7794
rect 3434 7788 3492 7794
rect 3644 7788 3702 7794
rect 3854 7788 3912 7794
rect 4064 7788 4122 7794
rect 4274 7788 4332 7794
rect 4484 7788 4542 7794
rect 4689 7776 4699 7794
rect 4751 7776 4761 7794
rect 4904 7788 4962 7794
rect 5114 7788 5172 7794
rect 5324 7788 5382 7794
rect 5534 7788 5592 7794
rect 5744 7788 5802 7794
rect -2350 7686 -2292 7692
rect -2140 7686 -2082 7692
rect -1930 7686 -1872 7692
rect -1720 7686 -1662 7692
rect -1510 7686 -1452 7692
rect -1300 7686 -1242 7692
rect -1090 7686 -1032 7692
rect -880 7686 -822 7692
rect -670 7686 -612 7692
rect -460 7686 -402 7692
rect -250 7686 -192 7692
rect -40 7686 18 7692
rect 170 7686 228 7692
rect 380 7686 438 7692
rect 590 7686 648 7692
rect 800 7686 858 7692
rect 1010 7686 1068 7692
rect 1220 7686 1278 7692
rect 1430 7686 1488 7692
rect 1640 7686 1698 7692
rect 1850 7686 1908 7692
rect 2060 7686 2118 7692
rect 2270 7686 2328 7692
rect 2391 7686 2401 7704
rect -2446 7652 -2338 7686
rect -2304 7652 -2128 7686
rect -2094 7652 -1918 7686
rect -1884 7652 -1708 7686
rect -1674 7652 -1498 7686
rect -1464 7652 -1288 7686
rect -1254 7652 -1078 7686
rect -1044 7652 -868 7686
rect -834 7652 -658 7686
rect -624 7652 -448 7686
rect -414 7652 -238 7686
rect -204 7652 -28 7686
rect 6 7652 182 7686
rect 216 7652 392 7686
rect 426 7652 602 7686
rect 636 7652 812 7686
rect 846 7652 1022 7686
rect 1056 7652 1232 7686
rect 1266 7652 1442 7686
rect 1476 7652 1652 7686
rect 1686 7652 1862 7686
rect 1896 7652 2072 7686
rect 2106 7652 2282 7686
rect 2316 7652 2401 7686
rect 2453 7692 2463 7704
rect 2453 7686 2538 7692
rect 2690 7686 2748 7692
rect 2900 7686 2958 7692
rect 3110 7686 3168 7692
rect 3320 7686 3378 7692
rect 3530 7686 3588 7692
rect 3740 7686 3798 7692
rect 3861 7686 3871 7704
rect 2453 7652 2492 7686
rect 2526 7652 2702 7686
rect 2736 7652 2912 7686
rect 2946 7652 3122 7686
rect 3156 7652 3332 7686
rect 3366 7652 3542 7686
rect 3576 7652 3752 7686
rect 3786 7652 3871 7686
rect 3923 7692 3933 7704
rect 3923 7686 4008 7692
rect 4160 7686 4218 7692
rect 4370 7686 4428 7692
rect 4580 7686 4638 7692
rect 4790 7686 4848 7692
rect 5000 7686 5058 7692
rect 5210 7686 5268 7692
rect 5330 7686 5340 7704
rect 3923 7652 3962 7686
rect 3996 7652 4172 7686
rect 4206 7652 4382 7686
rect 4416 7652 4592 7686
rect 4626 7652 4802 7686
rect 4836 7652 5012 7686
rect 5046 7652 5222 7686
rect 5256 7652 5340 7686
rect 5392 7692 5402 7704
rect 5392 7686 5478 7692
rect 5630 7686 5688 7692
rect 5840 7686 5898 7692
rect 5392 7652 5432 7686
rect 5466 7652 5642 7686
rect 5676 7652 5852 7686
rect 5886 7652 5898 7686
rect -2350 7646 -2292 7652
rect -2140 7646 -2082 7652
rect -1930 7646 -1872 7652
rect -1720 7646 -1662 7652
rect -1510 7646 -1452 7652
rect -1300 7646 -1242 7652
rect -1090 7646 -1032 7652
rect -880 7646 -822 7652
rect -670 7646 -612 7652
rect -460 7646 -402 7652
rect -250 7646 -192 7652
rect -40 7646 18 7652
rect 170 7646 228 7652
rect 380 7646 438 7652
rect 590 7646 648 7652
rect 800 7646 858 7652
rect 1010 7646 1068 7652
rect 1220 7646 1278 7652
rect 1430 7646 1488 7652
rect 1640 7646 1698 7652
rect 1850 7646 1908 7652
rect 2060 7646 2118 7652
rect 2270 7646 2328 7652
rect 2480 7646 2538 7652
rect 2690 7646 2748 7652
rect 2900 7646 2958 7652
rect 3110 7646 3168 7652
rect 3320 7646 3378 7652
rect 3530 7646 3588 7652
rect 3740 7646 3798 7652
rect 3950 7646 4008 7652
rect 4160 7646 4218 7652
rect 4370 7646 4428 7652
rect 4580 7646 4638 7652
rect 4790 7646 4848 7652
rect 5000 7646 5058 7652
rect 5210 7646 5268 7652
rect 5420 7646 5478 7652
rect 5630 7646 5688 7652
rect 5840 7646 5898 7652
rect -2188 7593 -2130 7599
rect -1768 7593 -1710 7599
rect -1348 7593 -1290 7599
rect -928 7593 -870 7599
rect -508 7593 -450 7599
rect -88 7593 -30 7599
rect 332 7593 390 7599
rect 752 7593 810 7599
rect 1172 7593 1230 7599
rect 1592 7593 1650 7599
rect 1960 7593 1970 7602
rect -2444 7559 -2176 7593
rect -2142 7559 -1756 7593
rect -1722 7559 -1336 7593
rect -1302 7559 -916 7593
rect -882 7559 -496 7593
rect -462 7559 -76 7593
rect -42 7559 344 7593
rect 378 7559 764 7593
rect 798 7559 1184 7593
rect 1218 7559 1604 7593
rect 1638 7559 1970 7593
rect -2188 7553 -2130 7559
rect -1768 7553 -1710 7559
rect -1348 7553 -1290 7559
rect -928 7553 -870 7559
rect -508 7553 -450 7559
rect -88 7553 -30 7559
rect 332 7553 390 7559
rect 752 7553 810 7559
rect 1172 7553 1230 7559
rect 1592 7553 1650 7559
rect 1960 7550 1970 7559
rect 2022 7599 2032 7602
rect 2022 7593 2070 7599
rect 2432 7593 2490 7599
rect 2852 7593 2910 7599
rect 3272 7593 3330 7599
rect 3692 7593 3750 7599
rect 4112 7593 4170 7599
rect 4532 7593 4590 7599
rect 4952 7593 5010 7599
rect 5372 7593 5430 7599
rect 5792 7593 5850 7599
rect 2022 7559 2024 7593
rect 2058 7559 2444 7593
rect 2478 7559 2864 7593
rect 2898 7559 3284 7593
rect 3318 7559 3704 7593
rect 3738 7559 4124 7593
rect 4158 7559 4544 7593
rect 4578 7559 4964 7593
rect 4998 7559 5384 7593
rect 5418 7559 5804 7593
rect 5838 7559 5898 7593
rect 2022 7553 2070 7559
rect 2432 7553 2490 7559
rect 2852 7553 2910 7559
rect 3272 7553 3330 7559
rect 3692 7553 3750 7559
rect 4112 7553 4170 7559
rect 4532 7553 4590 7559
rect 4952 7553 5010 7559
rect 5372 7553 5430 7559
rect 5792 7553 5850 7559
rect 2022 7550 2032 7553
rect 1436 7395 1458 7400
rect -2396 7389 -2338 7395
rect -1976 7389 -1918 7395
rect -1556 7389 -1498 7395
rect -1136 7389 -1078 7395
rect -716 7389 -658 7395
rect -296 7389 -238 7395
rect 124 7389 182 7395
rect 544 7389 602 7395
rect 964 7389 1022 7395
rect 1384 7389 1458 7395
rect -2444 7355 -2384 7389
rect -2350 7355 -1964 7389
rect -1930 7355 -1544 7389
rect -1510 7355 -1124 7389
rect -1090 7355 -704 7389
rect -670 7355 -284 7389
rect -250 7355 136 7389
rect 170 7355 556 7389
rect 590 7355 976 7389
rect 1010 7355 1396 7389
rect 1430 7355 1458 7389
rect -2396 7349 -2338 7355
rect -1976 7349 -1918 7355
rect -1556 7349 -1498 7355
rect -1136 7349 -1078 7355
rect -716 7349 -658 7355
rect -296 7349 -238 7355
rect 124 7349 182 7355
rect 544 7349 602 7355
rect 964 7349 1022 7355
rect 1384 7349 1458 7355
rect 1448 7348 1458 7349
rect 1510 7389 1520 7400
rect 1804 7389 1862 7395
rect 2224 7389 2282 7395
rect 2644 7389 2702 7395
rect 3064 7389 3122 7395
rect 3484 7389 3542 7395
rect 3904 7389 3962 7395
rect 4324 7389 4382 7395
rect 4744 7389 4802 7395
rect 5164 7389 5222 7395
rect 5584 7389 5642 7395
rect 1510 7355 1816 7389
rect 1850 7355 2236 7389
rect 2270 7355 2656 7389
rect 2690 7355 3076 7389
rect 3110 7355 3496 7389
rect 3530 7355 3916 7389
rect 3950 7355 4336 7389
rect 4370 7355 4756 7389
rect 4790 7355 5176 7389
rect 5210 7355 5596 7389
rect 5630 7355 5900 7389
rect 1510 7348 1520 7355
rect 1804 7349 1862 7355
rect 2224 7349 2282 7355
rect 2644 7349 2702 7355
rect 3064 7349 3122 7355
rect 3484 7349 3542 7355
rect 3904 7349 3962 7355
rect 4324 7349 4382 7355
rect 4744 7349 4802 7355
rect 5164 7349 5222 7355
rect 5584 7349 5642 7355
rect -2444 7296 -2386 7302
rect -2234 7296 -2176 7302
rect -2024 7296 -1966 7302
rect -1814 7296 -1756 7302
rect -1604 7296 -1546 7302
rect -1394 7296 -1336 7302
rect -1184 7296 -1126 7302
rect -974 7296 -916 7302
rect -764 7296 -706 7302
rect -554 7296 -496 7302
rect -344 7296 -286 7302
rect -134 7296 -76 7302
rect 76 7296 134 7302
rect 286 7296 344 7302
rect 496 7296 554 7302
rect 706 7296 764 7302
rect 916 7296 974 7302
rect 1126 7296 1184 7302
rect 1336 7296 1394 7302
rect 1546 7296 1604 7302
rect 1756 7296 1814 7302
rect 1966 7296 2024 7302
rect 2176 7296 2234 7302
rect 2386 7296 2444 7302
rect 2596 7296 2654 7302
rect 2806 7296 2864 7302
rect 3016 7296 3074 7302
rect 3226 7296 3284 7302
rect 3436 7296 3494 7302
rect 3646 7296 3704 7302
rect 3856 7296 3914 7302
rect 4066 7296 4124 7302
rect 4276 7296 4334 7302
rect 4486 7296 4544 7302
rect 4696 7296 4754 7302
rect 4906 7296 4964 7302
rect 5116 7296 5174 7302
rect 5326 7296 5384 7302
rect 5536 7296 5594 7302
rect 5746 7296 5804 7302
rect -2444 7262 -2432 7296
rect -2398 7262 -2222 7296
rect -2188 7262 -2012 7296
rect -1978 7262 -1802 7296
rect -1768 7262 -1592 7296
rect -1558 7262 -1382 7296
rect -1348 7262 -1286 7296
rect -2444 7256 -2386 7262
rect -2234 7256 -2176 7262
rect -2024 7256 -1966 7262
rect -1814 7256 -1756 7262
rect -1604 7256 -1546 7262
rect -1394 7256 -1336 7262
rect -1296 7244 -1286 7262
rect -1234 7262 -1172 7296
rect -1138 7262 -962 7296
rect -928 7262 -752 7296
rect -718 7262 -542 7296
rect -508 7262 -332 7296
rect -298 7262 -122 7296
rect -88 7262 88 7296
rect 122 7262 287 7296
rect 339 7262 508 7296
rect 542 7262 718 7296
rect 752 7262 928 7296
rect 962 7262 1138 7296
rect 1172 7262 1348 7296
rect 1382 7262 1558 7296
rect 1592 7262 1768 7296
rect 1802 7262 1978 7296
rect 2012 7262 2188 7296
rect 2222 7262 2398 7296
rect 2432 7262 2608 7296
rect 2642 7262 2818 7296
rect 2852 7262 3028 7296
rect 3062 7262 3230 7296
rect 3282 7262 3448 7296
rect 3482 7262 3658 7296
rect 3692 7262 3868 7296
rect 3902 7262 4078 7296
rect 4112 7262 4288 7296
rect 4322 7262 4498 7296
rect 4532 7262 4699 7296
rect 4751 7262 4918 7296
rect 4952 7262 5128 7296
rect 5162 7262 5338 7296
rect 5372 7262 5548 7296
rect 5582 7262 5758 7296
rect 5792 7262 5900 7296
rect -1234 7244 -1224 7262
rect -1184 7256 -1126 7262
rect -974 7256 -916 7262
rect -764 7256 -706 7262
rect -554 7256 -496 7262
rect -344 7256 -286 7262
rect -134 7256 -76 7262
rect 76 7256 134 7262
rect 277 7244 287 7262
rect 339 7244 349 7262
rect 496 7256 554 7262
rect 706 7256 764 7262
rect 916 7256 974 7262
rect 1126 7256 1184 7262
rect 1336 7256 1394 7262
rect 1546 7256 1604 7262
rect 1749 7244 1821 7262
rect 1966 7256 2024 7262
rect 2176 7256 2234 7262
rect 2386 7256 2444 7262
rect 2596 7256 2654 7262
rect 2806 7256 2864 7262
rect 3016 7256 3074 7262
rect 3220 7244 3230 7262
rect 3282 7244 3292 7262
rect 3436 7256 3494 7262
rect 3646 7256 3704 7262
rect 3856 7256 3914 7262
rect 4066 7256 4124 7262
rect 4276 7256 4334 7262
rect 4486 7256 4544 7262
rect 4689 7244 4699 7262
rect 4751 7244 4761 7262
rect 4906 7256 4964 7262
rect 5116 7256 5174 7262
rect 5326 7256 5384 7262
rect 5536 7256 5594 7262
rect 5746 7256 5804 7262
rect -2348 7154 -2290 7160
rect -2138 7154 -2080 7160
rect -2019 7154 -2009 7172
rect -2444 7120 -2336 7154
rect -2302 7120 -2126 7154
rect -2092 7120 -2009 7154
rect -1957 7160 -1947 7172
rect -1957 7154 -1870 7160
rect -1718 7154 -1660 7160
rect -1508 7154 -1450 7160
rect -1298 7154 -1240 7160
rect -1088 7154 -1030 7160
rect -878 7154 -820 7160
rect -668 7154 -610 7160
rect -549 7154 -539 7172
rect -1957 7120 -1916 7154
rect -1882 7120 -1706 7154
rect -1672 7120 -1496 7154
rect -1462 7120 -1286 7154
rect -1252 7120 -1076 7154
rect -1042 7120 -866 7154
rect -832 7120 -656 7154
rect -622 7120 -539 7154
rect -487 7160 -477 7172
rect -487 7154 -400 7160
rect -248 7154 -190 7160
rect -38 7154 20 7160
rect 172 7154 230 7160
rect 382 7154 440 7160
rect 592 7154 650 7160
rect 802 7154 860 7160
rect 921 7154 931 7172
rect -487 7120 -446 7154
rect -412 7120 -236 7154
rect -202 7120 -26 7154
rect 8 7120 184 7154
rect 218 7120 394 7154
rect 428 7120 604 7154
rect 638 7120 814 7154
rect 848 7120 931 7154
rect 983 7160 993 7172
rect 983 7154 1070 7160
rect 1222 7154 1280 7160
rect 1432 7154 1490 7160
rect 1642 7154 1700 7160
rect 1852 7154 1910 7160
rect 2062 7154 2120 7160
rect 2272 7154 2330 7160
rect 2482 7154 2540 7160
rect 2692 7154 2750 7160
rect 2902 7154 2960 7160
rect 3112 7154 3170 7160
rect 3322 7154 3380 7160
rect 3532 7154 3590 7160
rect 3742 7154 3800 7160
rect 3952 7154 4010 7160
rect 4162 7154 4220 7160
rect 4372 7154 4430 7160
rect 4582 7154 4640 7160
rect 4792 7154 4850 7160
rect 5002 7154 5060 7160
rect 5212 7154 5270 7160
rect 5422 7154 5480 7160
rect 5632 7154 5690 7160
rect 5842 7154 5900 7160
rect 983 7120 1024 7154
rect 1058 7120 1234 7154
rect 1268 7120 1444 7154
rect 1478 7120 1654 7154
rect 1688 7120 1864 7154
rect 1898 7120 2074 7154
rect 2108 7120 2284 7154
rect 2318 7120 2494 7154
rect 2528 7120 2704 7154
rect 2738 7120 2914 7154
rect 2948 7120 3124 7154
rect 3158 7120 3334 7154
rect 3368 7120 3544 7154
rect 3578 7120 3754 7154
rect 3788 7120 3964 7154
rect 3998 7120 4174 7154
rect 4208 7120 4384 7154
rect 4418 7120 4594 7154
rect 4628 7120 4804 7154
rect 4838 7120 5014 7154
rect 5048 7120 5224 7154
rect 5258 7120 5434 7154
rect 5468 7120 5644 7154
rect 5678 7120 5854 7154
rect 5888 7120 5900 7154
rect -2348 7114 -2290 7120
rect -2138 7114 -2080 7120
rect -1928 7114 -1870 7120
rect -1718 7114 -1660 7120
rect -1508 7114 -1450 7120
rect -1298 7114 -1240 7120
rect -1088 7114 -1030 7120
rect -878 7114 -820 7120
rect -668 7114 -610 7120
rect -458 7114 -400 7120
rect -248 7114 -190 7120
rect -38 7114 20 7120
rect 172 7114 230 7120
rect 382 7114 440 7120
rect 592 7114 650 7120
rect 802 7114 860 7120
rect 1012 7114 1070 7120
rect 1222 7114 1280 7120
rect 1432 7114 1490 7120
rect 1642 7114 1700 7120
rect 1852 7114 1910 7120
rect 2062 7114 2120 7120
rect 2272 7114 2330 7120
rect 2482 7114 2540 7120
rect 2692 7114 2750 7120
rect 2902 7114 2960 7120
rect 3112 7114 3170 7120
rect 3322 7114 3380 7120
rect 3532 7114 3590 7120
rect 3742 7114 3800 7120
rect 3952 7114 4010 7120
rect 4162 7114 4220 7120
rect 4372 7114 4430 7120
rect 4582 7114 4640 7120
rect 4792 7114 4850 7120
rect 5002 7114 5060 7120
rect 5212 7114 5270 7120
rect 5422 7114 5480 7120
rect 5632 7114 5690 7120
rect 5842 7114 5900 7120
rect -2186 7061 -2128 7066
rect -1766 7061 -1708 7066
rect -1346 7061 -1288 7066
rect -926 7061 -868 7066
rect -506 7061 -448 7066
rect -86 7061 -28 7066
rect 334 7061 392 7066
rect 754 7061 812 7066
rect 1174 7061 1232 7066
rect 1448 7061 1458 7070
rect -2432 7060 1458 7061
rect -2432 7027 -2174 7060
rect -2186 7026 -2174 7027
rect -2140 7027 -1754 7060
rect -2140 7026 -2128 7027
rect -2186 7020 -2128 7026
rect -1766 7026 -1754 7027
rect -1720 7027 -1334 7060
rect -1720 7026 -1708 7027
rect -1766 7020 -1708 7026
rect -1346 7026 -1334 7027
rect -1300 7027 -914 7060
rect -1300 7026 -1288 7027
rect -1346 7020 -1288 7026
rect -926 7026 -914 7027
rect -880 7027 -494 7060
rect -880 7026 -868 7027
rect -926 7020 -868 7026
rect -506 7026 -494 7027
rect -460 7027 -74 7060
rect -460 7026 -448 7027
rect -506 7020 -448 7026
rect -86 7026 -74 7027
rect -40 7027 346 7060
rect -40 7026 -28 7027
rect -86 7020 -28 7026
rect 334 7026 346 7027
rect 380 7027 766 7060
rect 380 7026 392 7027
rect 334 7020 392 7026
rect 754 7026 766 7027
rect 800 7027 1186 7060
rect 800 7026 812 7027
rect 754 7020 812 7026
rect 1174 7026 1186 7027
rect 1220 7027 1458 7060
rect 1220 7026 1232 7027
rect 1174 7020 1232 7026
rect 1448 7018 1458 7027
rect 1510 7061 1520 7070
rect 1594 7061 1652 7066
rect 2014 7061 2072 7066
rect 2434 7061 2492 7066
rect 2854 7061 2912 7066
rect 3274 7061 3332 7066
rect 3694 7061 3752 7066
rect 4114 7061 4172 7066
rect 4534 7061 4592 7066
rect 4954 7061 5012 7066
rect 5374 7061 5432 7066
rect 5794 7061 5852 7066
rect 1510 7060 5912 7061
rect 1510 7027 1606 7060
rect 1510 7018 1520 7027
rect 1594 7026 1606 7027
rect 1640 7027 2026 7060
rect 1640 7026 1652 7027
rect 1594 7020 1652 7026
rect 2014 7026 2026 7027
rect 2060 7027 2446 7060
rect 2060 7026 2072 7027
rect 2014 7020 2072 7026
rect 2434 7026 2446 7027
rect 2480 7027 2866 7060
rect 2480 7026 2492 7027
rect 2434 7020 2492 7026
rect 2854 7026 2866 7027
rect 2900 7027 3286 7060
rect 2900 7026 2912 7027
rect 2854 7020 2912 7026
rect 3274 7026 3286 7027
rect 3320 7027 3706 7060
rect 3320 7026 3332 7027
rect 3274 7020 3332 7026
rect 3694 7026 3706 7027
rect 3740 7027 4126 7060
rect 3740 7026 3752 7027
rect 3694 7020 3752 7026
rect 4114 7026 4126 7027
rect 4160 7027 4546 7060
rect 4160 7026 4172 7027
rect 4114 7020 4172 7026
rect 4534 7026 4546 7027
rect 4580 7027 4966 7060
rect 4580 7026 4592 7027
rect 4534 7020 4592 7026
rect 4954 7026 4966 7027
rect 5000 7027 5386 7060
rect 5000 7026 5012 7027
rect 4954 7020 5012 7026
rect 5374 7026 5386 7027
rect 5420 7027 5806 7060
rect 5420 7026 5432 7027
rect 5374 7020 5432 7026
rect 5794 7026 5806 7027
rect 5840 7027 5912 7060
rect 5840 7026 5852 7027
rect 5794 7020 5852 7026
rect 921 6793 931 6845
rect 983 6793 1970 6845
rect 2022 6793 2032 6845
rect -3082 6668 -3072 6720
rect -3020 6668 -2009 6720
rect -1957 6668 -1379 6720
rect -1327 6668 -539 6720
rect -487 6668 301 6720
rect 353 6668 931 6720
rect 983 6668 994 6720
rect 2390 6668 2401 6720
rect 2453 6668 3031 6720
rect 3083 6668 3871 6720
rect 3923 6668 4711 6720
rect 4763 6668 5340 6720
rect 5392 6668 6482 6720
rect 6534 6668 6544 6720
rect 1448 6536 1458 6588
rect 1510 6536 2401 6588
rect 2453 6536 2463 6588
rect -3668 6067 -3150 6073
rect -3668 6033 -3656 6067
rect -3282 6033 -3150 6067
rect -3668 6027 -3150 6033
rect -3220 5619 -3150 6027
rect -3668 5613 -3150 5619
rect -3668 5579 -3656 5613
rect -3282 5579 -3150 5613
rect -3668 5573 -3150 5579
rect -3557 5313 -3523 5573
rect -3427 5403 -3369 5409
rect -3427 5369 -3415 5403
rect -3381 5369 -3369 5403
rect -3427 5363 -3369 5369
rect -3322 5368 -3288 5371
rect -3569 5307 -3511 5313
rect -3650 5272 -3616 5275
rect -3569 5273 -3557 5307
rect -3523 5273 -3511 5307
rect -3654 5260 -3608 5272
rect -3569 5267 -3511 5273
rect -3654 5226 -3648 5260
rect -3614 5226 -3608 5260
rect -3654 5214 -3608 5226
rect -3650 5173 -3616 5214
rect -3670 5121 -3660 5173
rect -3608 5121 -3598 5173
rect -3557 5121 -3523 5267
rect -3415 5217 -3381 5363
rect -3326 5356 -3280 5368
rect -3326 5322 -3320 5356
rect -3286 5322 -3280 5356
rect -3326 5310 -3280 5322
rect -3427 5211 -3369 5217
rect -3427 5177 -3415 5211
rect -3381 5177 -3369 5211
rect -3427 5171 -3369 5177
rect -3322 5176 -3288 5310
rect -3326 5173 -3280 5176
rect -3650 5080 -3616 5121
rect -3569 5115 -3511 5121
rect -3569 5081 -3557 5115
rect -3523 5081 -3511 5115
rect -3654 5068 -3608 5080
rect -3569 5075 -3511 5081
rect -3654 5034 -3648 5068
rect -3614 5034 -3608 5068
rect -3654 5022 -3608 5034
rect -3650 4888 -3616 5022
rect -3557 4929 -3523 5075
rect -3415 5025 -3381 5171
rect -3339 5121 -3329 5173
rect -3277 5121 -3267 5173
rect -3326 5118 -3280 5121
rect -3427 5019 -3369 5025
rect -3427 4985 -3415 5019
rect -3381 4985 -3369 5019
rect -3427 4979 -3369 4985
rect -3322 4984 -3288 5118
rect -3569 4923 -3511 4929
rect -3569 4889 -3557 4923
rect -3523 4889 -3511 4923
rect -3654 4876 -3608 4888
rect -3569 4883 -3511 4889
rect -3654 4842 -3648 4876
rect -3614 4842 -3608 4876
rect -3654 4830 -3608 4842
rect -3650 4696 -3616 4830
rect -3557 4737 -3523 4883
rect -3415 4833 -3381 4979
rect -3326 4972 -3280 4984
rect -3326 4938 -3320 4972
rect -3286 4938 -3280 4972
rect -3326 4926 -3280 4938
rect -3427 4827 -3369 4833
rect -3427 4793 -3415 4827
rect -3381 4793 -3369 4827
rect -3427 4787 -3369 4793
rect -3322 4792 -3288 4926
rect -3569 4731 -3511 4737
rect -3569 4697 -3557 4731
rect -3523 4697 -3511 4731
rect -3654 4684 -3608 4696
rect -3569 4691 -3511 4697
rect -3654 4650 -3648 4684
rect -3614 4650 -3608 4684
rect -3654 4638 -3608 4650
rect -3650 4504 -3616 4638
rect -3557 4545 -3523 4691
rect -3415 4641 -3381 4787
rect -3326 4780 -3280 4792
rect -3326 4746 -3320 4780
rect -3286 4746 -3280 4780
rect -3326 4734 -3280 4746
rect -3427 4635 -3369 4641
rect -3427 4601 -3415 4635
rect -3381 4601 -3369 4635
rect -3427 4595 -3369 4601
rect -3322 4600 -3288 4734
rect -3569 4539 -3511 4545
rect -3569 4505 -3557 4539
rect -3523 4505 -3511 4539
rect -3654 4492 -3608 4504
rect -3569 4499 -3511 4505
rect -3654 4458 -3648 4492
rect -3614 4458 -3608 4492
rect -3654 4446 -3608 4458
rect -3650 4312 -3616 4446
rect -3557 4353 -3523 4499
rect -3415 4497 -3381 4595
rect -3326 4588 -3280 4600
rect -3326 4554 -3320 4588
rect -3286 4554 -3280 4588
rect -3326 4542 -3280 4554
rect -3435 4445 -3425 4497
rect -3373 4445 -3363 4497
rect -3427 4443 -3369 4445
rect -3427 4409 -3415 4443
rect -3381 4409 -3369 4443
rect -3427 4403 -3369 4409
rect -3322 4408 -3288 4542
rect -3569 4347 -3511 4353
rect -3569 4313 -3557 4347
rect -3523 4313 -3511 4347
rect -3654 4300 -3608 4312
rect -3569 4307 -3511 4313
rect -3654 4266 -3648 4300
rect -3614 4266 -3608 4300
rect -3654 4254 -3608 4266
rect -3650 4120 -3616 4254
rect -3557 4161 -3523 4307
rect -3415 4257 -3381 4403
rect -3326 4396 -3280 4408
rect -3326 4362 -3320 4396
rect -3286 4362 -3280 4396
rect -3326 4350 -3280 4362
rect -3427 4251 -3369 4257
rect -3427 4217 -3415 4251
rect -3381 4217 -3369 4251
rect -3427 4211 -3369 4217
rect -3322 4216 -3288 4350
rect -3569 4155 -3511 4161
rect -3569 4121 -3557 4155
rect -3523 4121 -3511 4155
rect -3654 4108 -3608 4120
rect -3569 4115 -3511 4121
rect -3654 4074 -3648 4108
rect -3614 4074 -3608 4108
rect -3654 4062 -3608 4074
rect -3650 4021 -3616 4062
rect -3670 3969 -3660 4021
rect -3608 3969 -3598 4021
rect -3557 3969 -3523 4115
rect -3415 4065 -3381 4211
rect -3326 4204 -3280 4216
rect -3326 4170 -3320 4204
rect -3286 4170 -3280 4204
rect -3326 4158 -3280 4170
rect -3427 4059 -3369 4065
rect -3427 4025 -3415 4059
rect -3381 4025 -3369 4059
rect -3427 4019 -3369 4025
rect -3322 4024 -3288 4158
rect -3326 4021 -3280 4024
rect -3650 3928 -3616 3969
rect -3569 3963 -3511 3969
rect -3569 3929 -3557 3963
rect -3523 3929 -3511 3963
rect -3654 3916 -3608 3928
rect -3569 3923 -3511 3929
rect -3654 3882 -3648 3916
rect -3614 3882 -3608 3916
rect -3654 3870 -3608 3882
rect -3415 3873 -3381 4019
rect -3341 3969 -3331 4021
rect -3279 3969 -3269 4021
rect -3326 3966 -3280 3969
rect -3322 3961 -3288 3966
rect -3650 3865 -3616 3870
rect -3427 3867 -3369 3873
rect -3427 3833 -3415 3867
rect -3381 3833 -3369 3867
rect -3427 3827 -3369 3833
rect -3220 3663 -3150 5573
rect -2845 6435 -2704 6447
rect -2845 6412 -2744 6435
rect -2845 6360 -2798 6412
rect -2746 6360 -2744 6412
rect -2845 6271 -2744 6360
rect -2845 6219 -2798 6271
rect -2746 6219 -2744 6271
rect -2845 6130 -2744 6219
rect -2845 6078 -2798 6130
rect -2746 6078 -2744 6130
rect -2845 5989 -2744 6078
rect -2845 5937 -2798 5989
rect -2746 5937 -2744 5989
rect -2845 5848 -2744 5937
rect -2845 5796 -2798 5848
rect -2746 5796 -2744 5848
rect -2845 5707 -2744 5796
rect -2845 5655 -2798 5707
rect -2746 5655 -2744 5707
rect -2845 5566 -2744 5655
rect -2845 5514 -2798 5566
rect -2746 5514 -2744 5566
rect -2845 5425 -2744 5514
rect -2845 5373 -2798 5425
rect -2746 5373 -2744 5425
rect -2845 5284 -2744 5373
rect -2845 5232 -2798 5284
rect -2746 5232 -2744 5284
rect -2845 5143 -2744 5232
rect -2845 5091 -2798 5143
rect -2746 5091 -2744 5143
rect -2845 5002 -2744 5091
rect -2845 4950 -2798 5002
rect -2746 4950 -2744 5002
rect -2845 4861 -2744 4950
rect -2845 4809 -2798 4861
rect -2746 4809 -2744 4861
rect -2845 4759 -2744 4809
rect -2710 4759 -2704 6435
rect -2384 6429 -2326 6435
rect -1964 6429 -1906 6435
rect -1544 6429 -1486 6435
rect -1124 6429 -1066 6435
rect -704 6429 -646 6435
rect -284 6429 -226 6435
rect 136 6429 194 6435
rect 556 6429 614 6435
rect 976 6429 1034 6435
rect 1396 6429 1454 6435
rect 1816 6429 1874 6435
rect 1960 6429 1970 6438
rect -2432 6395 -2372 6429
rect -2338 6395 -1952 6429
rect -1918 6395 -1532 6429
rect -1498 6395 -1112 6429
rect -1078 6395 -692 6429
rect -658 6395 -272 6429
rect -238 6395 148 6429
rect 182 6395 568 6429
rect 602 6395 988 6429
rect 1022 6395 1408 6429
rect 1442 6395 1828 6429
rect 1862 6395 1970 6429
rect -2384 6389 -2326 6395
rect -1964 6389 -1906 6395
rect -1544 6389 -1486 6395
rect -1124 6389 -1066 6395
rect -704 6389 -646 6395
rect -284 6389 -226 6395
rect 136 6389 194 6395
rect 556 6389 614 6395
rect 976 6389 1034 6395
rect 1396 6389 1454 6395
rect 1816 6389 1874 6395
rect 1960 6386 1970 6395
rect 2022 6429 2032 6438
rect 6186 6435 6322 6447
rect 2236 6429 2294 6435
rect 2656 6429 2714 6435
rect 3076 6429 3134 6435
rect 3496 6429 3554 6435
rect 3916 6429 3974 6435
rect 4336 6429 4394 6435
rect 4756 6429 4814 6435
rect 5176 6429 5234 6435
rect 5596 6429 5654 6435
rect 2022 6395 2248 6429
rect 2282 6395 2668 6429
rect 2702 6395 3088 6429
rect 3122 6395 3508 6429
rect 3542 6395 3928 6429
rect 3962 6395 4348 6429
rect 4382 6395 4768 6429
rect 4802 6395 5188 6429
rect 5222 6395 5608 6429
rect 5642 6395 5900 6429
rect 2022 6386 2032 6395
rect 2236 6389 2294 6395
rect 2656 6389 2714 6395
rect 3076 6389 3134 6395
rect 3496 6389 3554 6395
rect 3916 6389 3974 6395
rect 4336 6389 4394 6395
rect 4756 6389 4814 6395
rect 5176 6389 5234 6395
rect 5596 6389 5654 6395
rect -2432 6345 -2374 6351
rect -2222 6345 -2164 6351
rect -2012 6345 -1954 6351
rect -1802 6345 -1744 6351
rect -1592 6345 -1534 6351
rect -1382 6345 -1324 6351
rect -1172 6345 -1114 6351
rect -962 6345 -904 6351
rect -752 6345 -694 6351
rect -542 6345 -484 6351
rect -332 6345 -274 6351
rect -122 6345 -64 6351
rect 88 6345 146 6351
rect 298 6345 356 6351
rect 508 6345 566 6351
rect 718 6345 776 6351
rect 928 6345 986 6351
rect 1138 6345 1196 6351
rect 1348 6345 1406 6351
rect 1558 6345 1616 6351
rect 1768 6345 1826 6351
rect 1978 6345 2036 6351
rect 2188 6345 2246 6351
rect 2398 6345 2456 6351
rect 2608 6345 2666 6351
rect 2818 6345 2876 6351
rect 3028 6345 3086 6351
rect 3238 6345 3296 6351
rect 3448 6345 3506 6351
rect 3658 6345 3716 6351
rect 3868 6345 3926 6351
rect 4078 6345 4136 6351
rect 4288 6345 4346 6351
rect 4498 6345 4556 6351
rect 4708 6345 4766 6351
rect 4918 6345 4976 6351
rect 5128 6345 5186 6351
rect 5338 6345 5396 6351
rect 5548 6345 5606 6351
rect 5758 6345 5816 6351
rect -2432 6311 -2420 6345
rect -2386 6311 -2210 6345
rect -2176 6311 -2000 6345
rect -1966 6311 -1790 6345
rect -1756 6311 -1580 6345
rect -1546 6311 -1370 6345
rect -1336 6311 -1160 6345
rect -1126 6311 -950 6345
rect -916 6311 -740 6345
rect -706 6311 -530 6345
rect -496 6311 -320 6345
rect -286 6311 -110 6345
rect -76 6311 100 6345
rect 134 6311 310 6345
rect 344 6311 520 6345
rect 554 6311 730 6345
rect 764 6311 940 6345
rect 974 6311 1150 6345
rect 1184 6311 1360 6345
rect 1394 6311 1570 6345
rect 1604 6311 1780 6345
rect 1814 6311 1990 6345
rect 2024 6311 2200 6345
rect 2234 6311 2410 6345
rect 2444 6311 2620 6345
rect 2654 6311 2830 6345
rect 2864 6311 3031 6345
rect 3083 6311 3250 6345
rect 3284 6311 3460 6345
rect 3494 6311 3670 6345
rect 3704 6311 3880 6345
rect 3914 6311 4090 6345
rect 4124 6311 4300 6345
rect 4334 6311 4510 6345
rect 4544 6311 4711 6345
rect 4763 6311 4930 6345
rect 4964 6311 5140 6345
rect 5174 6311 5350 6345
rect 5384 6311 5560 6345
rect 5594 6311 5770 6345
rect 5804 6311 5912 6345
rect -2432 6305 -2374 6311
rect -2222 6305 -2164 6311
rect -2012 6305 -1954 6311
rect -1802 6305 -1744 6311
rect -1592 6305 -1534 6311
rect -1382 6305 -1324 6311
rect -1172 6305 -1114 6311
rect -962 6305 -904 6311
rect -752 6305 -694 6311
rect -542 6305 -484 6311
rect -332 6305 -274 6311
rect -122 6305 -64 6311
rect 88 6305 146 6311
rect 298 6305 356 6311
rect 508 6305 566 6311
rect 718 6305 776 6311
rect 928 6305 986 6311
rect 1138 6305 1196 6311
rect 1348 6305 1406 6311
rect 1558 6305 1616 6311
rect 1768 6305 1826 6311
rect 1978 6305 2036 6311
rect 2188 6305 2246 6311
rect 2398 6305 2456 6311
rect 2608 6305 2666 6311
rect 2818 6305 2876 6311
rect 3021 6293 3031 6311
rect 3083 6293 3093 6311
rect 3238 6305 3296 6311
rect 3448 6305 3506 6311
rect 3658 6305 3716 6311
rect 3868 6305 3926 6311
rect 4078 6305 4136 6311
rect 4288 6305 4346 6311
rect 4498 6305 4556 6311
rect 4701 6293 4711 6311
rect 4763 6293 4773 6311
rect 4918 6305 4976 6311
rect 5128 6305 5186 6311
rect 5338 6305 5396 6311
rect 5548 6305 5606 6311
rect 5758 6305 5816 6311
rect -2336 6203 -2278 6209
rect -2126 6203 -2068 6209
rect -1916 6203 -1858 6209
rect -1706 6203 -1648 6209
rect -1496 6203 -1438 6209
rect -1286 6203 -1228 6209
rect -1076 6203 -1018 6209
rect -866 6203 -808 6209
rect -656 6203 -598 6209
rect -446 6203 -388 6209
rect -236 6203 -178 6209
rect -26 6203 32 6209
rect 184 6203 242 6209
rect 394 6203 452 6209
rect 604 6203 662 6209
rect 814 6203 872 6209
rect 1024 6203 1082 6209
rect 1234 6203 1292 6209
rect 1444 6203 1502 6209
rect 1654 6203 1712 6209
rect 1864 6203 1922 6209
rect 2074 6203 2132 6209
rect 2284 6203 2342 6209
rect 2391 6203 2401 6221
rect -2432 6169 -2324 6203
rect -2290 6169 -2114 6203
rect -2080 6169 -1904 6203
rect -1870 6169 -1694 6203
rect -1660 6169 -1484 6203
rect -1450 6169 -1274 6203
rect -1240 6169 -1064 6203
rect -1030 6169 -854 6203
rect -820 6169 -644 6203
rect -610 6169 -434 6203
rect -400 6169 -224 6203
rect -190 6169 -14 6203
rect 20 6169 196 6203
rect 230 6169 406 6203
rect 440 6169 616 6203
rect 650 6169 826 6203
rect 860 6169 1036 6203
rect 1070 6169 1246 6203
rect 1280 6169 1456 6203
rect 1490 6169 1666 6203
rect 1700 6169 1876 6203
rect 1910 6169 2086 6203
rect 2120 6169 2296 6203
rect 2330 6169 2401 6203
rect 2453 6203 2463 6221
rect 2494 6203 2552 6209
rect 2704 6203 2762 6209
rect 2914 6203 2972 6209
rect 3124 6203 3182 6209
rect 3334 6203 3392 6209
rect 3544 6203 3602 6209
rect 3754 6203 3812 6209
rect 3861 6203 3871 6221
rect 2453 6169 2506 6203
rect 2540 6169 2716 6203
rect 2750 6169 2926 6203
rect 2960 6169 3136 6203
rect 3170 6169 3346 6203
rect 3380 6169 3556 6203
rect 3590 6169 3766 6203
rect 3800 6169 3871 6203
rect 3923 6203 3933 6221
rect 3964 6203 4022 6209
rect 4174 6203 4232 6209
rect 4384 6203 4442 6209
rect 4594 6203 4652 6209
rect 4804 6203 4862 6209
rect 5014 6203 5072 6209
rect 5224 6203 5282 6209
rect 5330 6203 5340 6221
rect 3923 6169 3976 6203
rect 4010 6169 4186 6203
rect 4220 6169 4396 6203
rect 4430 6169 4606 6203
rect 4640 6169 4816 6203
rect 4850 6169 5026 6203
rect 5060 6169 5236 6203
rect 5270 6169 5340 6203
rect 5392 6203 5402 6221
rect 5434 6203 5492 6209
rect 5644 6203 5702 6209
rect 5854 6203 5912 6209
rect 5392 6169 5446 6203
rect 5480 6169 5656 6203
rect 5690 6169 5866 6203
rect 5900 6169 5912 6203
rect -2336 6163 -2278 6169
rect -2126 6163 -2068 6169
rect -1916 6163 -1858 6169
rect -1706 6163 -1648 6169
rect -1496 6163 -1438 6169
rect -1286 6163 -1228 6169
rect -1076 6163 -1018 6169
rect -866 6163 -808 6169
rect -656 6163 -598 6169
rect -446 6163 -388 6169
rect -236 6163 -178 6169
rect -26 6163 32 6169
rect 184 6163 242 6169
rect 394 6163 452 6169
rect 604 6163 662 6169
rect 814 6163 872 6169
rect 1024 6163 1082 6169
rect 1234 6163 1292 6169
rect 1444 6163 1502 6169
rect 1654 6163 1712 6169
rect 1864 6163 1922 6169
rect 2074 6163 2132 6169
rect 2284 6163 2342 6169
rect 2494 6163 2552 6169
rect 2704 6163 2762 6169
rect 2914 6163 2972 6169
rect 3124 6163 3182 6169
rect 3334 6163 3392 6169
rect 3544 6163 3602 6169
rect 3754 6163 3812 6169
rect 3964 6163 4022 6169
rect 4174 6163 4232 6169
rect 4384 6163 4442 6169
rect 4594 6163 4652 6169
rect 4804 6163 4862 6169
rect 5014 6163 5072 6169
rect 5224 6163 5282 6169
rect 5434 6163 5492 6169
rect 5644 6163 5702 6169
rect 5854 6163 5912 6169
rect -2174 6119 -2116 6125
rect -1754 6119 -1696 6125
rect -1334 6119 -1276 6125
rect -914 6119 -856 6125
rect -494 6119 -436 6125
rect -74 6119 -16 6125
rect 346 6119 404 6125
rect 766 6119 824 6125
rect 1186 6119 1244 6125
rect 1606 6119 1664 6125
rect 1960 6119 1970 6128
rect -2432 6085 -2162 6119
rect -2128 6085 -1742 6119
rect -1708 6085 -1322 6119
rect -1288 6085 -902 6119
rect -868 6085 -482 6119
rect -448 6085 -62 6119
rect -28 6085 358 6119
rect 392 6085 778 6119
rect 812 6085 1198 6119
rect 1232 6085 1618 6119
rect 1652 6085 1970 6119
rect -2174 6079 -2116 6085
rect -1754 6079 -1696 6085
rect -1334 6079 -1276 6085
rect -914 6079 -856 6085
rect -494 6079 -436 6085
rect -74 6079 -16 6085
rect 346 6079 404 6085
rect 766 6079 824 6085
rect 1186 6079 1244 6085
rect 1606 6079 1664 6085
rect 1960 6076 1970 6085
rect 2022 6125 2032 6128
rect 2022 6119 2084 6125
rect 2446 6119 2504 6125
rect 2866 6119 2924 6125
rect 3286 6119 3344 6125
rect 3706 6119 3764 6125
rect 4126 6119 4184 6125
rect 4546 6119 4604 6125
rect 4966 6119 5024 6125
rect 5386 6119 5444 6125
rect 5806 6119 5864 6125
rect 2022 6085 2038 6119
rect 2072 6085 2458 6119
rect 2492 6085 2878 6119
rect 2912 6085 3298 6119
rect 3332 6085 3718 6119
rect 3752 6085 4138 6119
rect 4172 6085 4558 6119
rect 4592 6085 4978 6119
rect 5012 6085 5398 6119
rect 5432 6085 5818 6119
rect 5852 6085 5900 6119
rect 2022 6079 2084 6085
rect 2446 6079 2504 6085
rect 2866 6079 2924 6085
rect 3286 6079 3344 6085
rect 3706 6079 3764 6085
rect 4126 6079 4184 6085
rect 4546 6079 4604 6085
rect 4966 6079 5024 6085
rect 5386 6079 5444 6085
rect 5806 6079 5864 6085
rect 2022 6076 2032 6079
rect 1448 5995 1458 5998
rect -2384 5989 -2326 5995
rect -1964 5989 -1906 5995
rect -1544 5989 -1486 5995
rect -1124 5989 -1066 5995
rect -704 5989 -646 5995
rect -284 5989 -226 5995
rect 136 5989 194 5995
rect 556 5989 614 5995
rect 976 5989 1034 5995
rect 1396 5989 1458 5995
rect -2432 5955 -2372 5989
rect -2338 5955 -1952 5989
rect -1918 5955 -1532 5989
rect -1498 5955 -1112 5989
rect -1078 5955 -692 5989
rect -658 5955 -272 5989
rect -238 5955 148 5989
rect 182 5955 568 5989
rect 602 5955 988 5989
rect 1022 5955 1408 5989
rect 1442 5955 1458 5989
rect -2384 5949 -2326 5955
rect -1964 5949 -1906 5955
rect -1544 5949 -1486 5955
rect -1124 5949 -1066 5955
rect -704 5949 -646 5955
rect -284 5949 -226 5955
rect 136 5949 194 5955
rect 556 5949 614 5955
rect 976 5949 1034 5955
rect 1396 5949 1458 5955
rect 1448 5946 1458 5949
rect 1510 5989 1520 5998
rect 1816 5989 1874 5995
rect 2236 5989 2294 5995
rect 2656 5989 2714 5995
rect 3076 5989 3134 5995
rect 3496 5989 3554 5995
rect 3916 5989 3974 5995
rect 4336 5989 4394 5995
rect 4756 5989 4814 5995
rect 5176 5989 5234 5995
rect 5596 5989 5654 5995
rect 1510 5955 1828 5989
rect 1862 5955 2248 5989
rect 2282 5955 2668 5989
rect 2702 5955 3088 5989
rect 3122 5955 3508 5989
rect 3542 5955 3928 5989
rect 3962 5955 4348 5989
rect 4382 5955 4768 5989
rect 4802 5955 5188 5989
rect 5222 5955 5608 5989
rect 5642 5955 5900 5989
rect 1510 5946 1520 5955
rect 1816 5949 1874 5955
rect 2236 5949 2294 5955
rect 2656 5949 2714 5955
rect 3076 5949 3134 5955
rect 3496 5949 3554 5955
rect 3916 5949 3974 5955
rect 4336 5949 4394 5955
rect 4756 5949 4814 5955
rect 5176 5949 5234 5955
rect 5596 5949 5654 5955
rect -2432 5905 -2374 5911
rect -2222 5905 -2164 5911
rect -2012 5905 -1954 5911
rect -1802 5905 -1744 5911
rect -1592 5905 -1534 5911
rect -1382 5905 -1324 5911
rect -1172 5905 -1114 5911
rect -962 5905 -904 5911
rect -752 5905 -694 5911
rect -542 5905 -484 5911
rect -332 5905 -274 5911
rect -122 5905 -64 5911
rect 88 5905 146 5911
rect 298 5905 356 5911
rect 508 5905 566 5911
rect 718 5905 776 5911
rect 928 5905 986 5911
rect 1138 5905 1196 5911
rect 1348 5905 1406 5911
rect 1558 5905 1616 5911
rect 1768 5905 1826 5911
rect 1978 5905 2036 5911
rect 2188 5905 2246 5911
rect 2398 5905 2456 5911
rect 2608 5905 2666 5911
rect 2818 5905 2876 5911
rect 3028 5905 3086 5911
rect 3238 5905 3296 5911
rect 3448 5905 3506 5911
rect 3658 5905 3716 5911
rect 3868 5905 3926 5911
rect 4078 5905 4136 5911
rect 4288 5905 4346 5911
rect 4498 5905 4556 5911
rect 4708 5905 4766 5911
rect 4918 5905 4976 5911
rect 5128 5905 5186 5911
rect 5338 5905 5396 5911
rect 5548 5905 5606 5911
rect 5758 5905 5816 5911
rect -2432 5871 -2420 5905
rect -2386 5871 -2210 5905
rect -2176 5871 -2000 5905
rect -1966 5871 -1790 5905
rect -1756 5871 -1580 5905
rect -1546 5871 -1379 5905
rect -1327 5871 -1160 5905
rect -1126 5871 -950 5905
rect -916 5871 -740 5905
rect -706 5871 -530 5905
rect -496 5871 -320 5905
rect -286 5871 -110 5905
rect -76 5871 100 5905
rect 134 5871 301 5905
rect 353 5871 520 5905
rect 554 5871 730 5905
rect 764 5871 940 5905
rect 974 5871 1150 5905
rect 1184 5871 1360 5905
rect 1394 5871 1570 5905
rect 1604 5871 1780 5905
rect 1814 5871 1990 5905
rect 2024 5871 2200 5905
rect 2234 5871 2410 5905
rect 2444 5871 2620 5905
rect 2654 5871 2830 5905
rect 2864 5871 3040 5905
rect 3074 5871 3250 5905
rect 3284 5871 3460 5905
rect 3494 5871 3670 5905
rect 3704 5871 3880 5905
rect 3914 5871 4090 5905
rect 4124 5871 4300 5905
rect 4334 5871 4510 5905
rect 4544 5871 4720 5905
rect 4754 5871 4930 5905
rect 4964 5871 5140 5905
rect 5174 5871 5350 5905
rect 5384 5871 5560 5905
rect 5594 5871 5770 5905
rect 5804 5871 5912 5905
rect -2432 5865 -2374 5871
rect -2222 5865 -2164 5871
rect -2012 5865 -1954 5871
rect -1802 5865 -1744 5871
rect -1592 5865 -1534 5871
rect -1389 5853 -1379 5871
rect -1327 5853 -1317 5871
rect -1172 5865 -1114 5871
rect -962 5865 -904 5871
rect -752 5865 -694 5871
rect -542 5865 -484 5871
rect -332 5865 -274 5871
rect -122 5865 -64 5871
rect 88 5865 146 5871
rect 291 5853 301 5871
rect 353 5853 363 5871
rect 508 5865 566 5871
rect 718 5865 776 5871
rect 928 5865 986 5871
rect 1138 5865 1196 5871
rect 1348 5865 1406 5871
rect 1558 5865 1616 5871
rect 1768 5865 1826 5871
rect 1978 5865 2036 5871
rect 2188 5865 2246 5871
rect 2398 5865 2456 5871
rect 2608 5865 2666 5871
rect 2818 5865 2876 5871
rect 3028 5865 3086 5871
rect 3238 5865 3296 5871
rect 3448 5865 3506 5871
rect 3658 5865 3716 5871
rect 3868 5865 3926 5871
rect 4078 5865 4136 5871
rect 4288 5865 4346 5871
rect 4498 5865 4556 5871
rect 4708 5865 4766 5871
rect 4918 5865 4976 5871
rect 5128 5865 5186 5871
rect 5338 5865 5396 5871
rect 5548 5865 5606 5871
rect 5758 5865 5816 5871
rect -2336 5763 -2278 5769
rect -2126 5763 -2068 5769
rect -2019 5763 -2009 5781
rect -2432 5729 -2324 5763
rect -2290 5729 -2114 5763
rect -2080 5729 -2009 5763
rect -1957 5763 -1947 5781
rect -1916 5763 -1858 5769
rect -1706 5763 -1648 5769
rect -1496 5763 -1438 5769
rect -1286 5763 -1228 5769
rect -1076 5763 -1018 5769
rect -866 5763 -808 5769
rect -656 5763 -598 5769
rect -549 5763 -539 5781
rect -1957 5729 -1904 5763
rect -1870 5729 -1694 5763
rect -1660 5729 -1484 5763
rect -1450 5729 -1274 5763
rect -1240 5729 -1064 5763
rect -1030 5729 -854 5763
rect -820 5729 -644 5763
rect -610 5729 -539 5763
rect -487 5763 -477 5781
rect -446 5763 -388 5769
rect -236 5763 -178 5769
rect -26 5763 32 5769
rect 184 5763 242 5769
rect 394 5763 452 5769
rect 604 5763 662 5769
rect 814 5763 872 5769
rect 921 5763 931 5781
rect -487 5729 -434 5763
rect -400 5729 -224 5763
rect -190 5729 -14 5763
rect 20 5729 196 5763
rect 230 5729 406 5763
rect 440 5729 616 5763
rect 650 5729 826 5763
rect 860 5729 931 5763
rect 983 5763 993 5781
rect 1024 5763 1082 5769
rect 1234 5763 1292 5769
rect 1444 5763 1502 5769
rect 1654 5763 1712 5769
rect 1864 5763 1922 5769
rect 2074 5763 2132 5769
rect 2284 5763 2342 5769
rect 2494 5763 2552 5769
rect 2704 5763 2762 5769
rect 2914 5763 2972 5769
rect 3124 5763 3182 5769
rect 3334 5763 3392 5769
rect 3544 5763 3602 5769
rect 3754 5763 3812 5769
rect 3964 5763 4022 5769
rect 4174 5763 4232 5769
rect 4384 5763 4442 5769
rect 4594 5763 4652 5769
rect 4804 5763 4862 5769
rect 5014 5763 5072 5769
rect 5224 5763 5282 5769
rect 5434 5763 5492 5769
rect 5644 5763 5702 5769
rect 5854 5763 5912 5769
rect 983 5729 1036 5763
rect 1070 5729 1246 5763
rect 1280 5729 1456 5763
rect 1490 5729 1666 5763
rect 1700 5729 1876 5763
rect 1910 5729 2086 5763
rect 2120 5729 2296 5763
rect 2330 5729 2506 5763
rect 2540 5729 2716 5763
rect 2750 5729 2926 5763
rect 2960 5729 3136 5763
rect 3170 5729 3346 5763
rect 3380 5729 3556 5763
rect 3590 5729 3766 5763
rect 3800 5729 3976 5763
rect 4010 5729 4186 5763
rect 4220 5729 4396 5763
rect 4430 5729 4606 5763
rect 4640 5729 4816 5763
rect 4850 5729 5026 5763
rect 5060 5729 5236 5763
rect 5270 5729 5446 5763
rect 5480 5729 5656 5763
rect 5690 5729 5866 5763
rect 5900 5729 5912 5763
rect -2336 5723 -2278 5729
rect -2126 5723 -2068 5729
rect -1916 5723 -1858 5729
rect -1706 5723 -1648 5729
rect -1496 5723 -1438 5729
rect -1286 5723 -1228 5729
rect -1076 5723 -1018 5729
rect -866 5723 -808 5729
rect -656 5723 -598 5729
rect -446 5723 -388 5729
rect -236 5723 -178 5729
rect -26 5723 32 5729
rect 184 5723 242 5729
rect 394 5723 452 5729
rect 604 5723 662 5729
rect 814 5723 872 5729
rect 1024 5723 1082 5729
rect 1234 5723 1292 5729
rect 1444 5723 1502 5729
rect 1654 5723 1712 5729
rect 1864 5723 1922 5729
rect 2074 5723 2132 5729
rect 2284 5723 2342 5729
rect 2494 5723 2552 5729
rect 2704 5723 2762 5729
rect 2914 5723 2972 5729
rect 3124 5723 3182 5729
rect 3334 5723 3392 5729
rect 3544 5723 3602 5729
rect 3754 5723 3812 5729
rect 3964 5723 4022 5729
rect 4174 5723 4232 5729
rect 4384 5723 4442 5729
rect 4594 5723 4652 5729
rect 4804 5723 4862 5729
rect 5014 5723 5072 5729
rect 5224 5723 5282 5729
rect 5434 5723 5492 5729
rect 5644 5723 5702 5729
rect 5854 5723 5912 5729
rect -2174 5679 -2116 5685
rect -1754 5679 -1696 5685
rect -1334 5679 -1276 5685
rect -914 5679 -856 5685
rect -494 5679 -436 5685
rect -74 5679 -16 5685
rect 346 5679 404 5685
rect 766 5679 824 5685
rect 1186 5679 1244 5685
rect 1448 5679 1458 5686
rect -2432 5645 -2162 5679
rect -2128 5645 -1742 5679
rect -1708 5645 -1322 5679
rect -1288 5645 -902 5679
rect -868 5645 -482 5679
rect -448 5645 -62 5679
rect -28 5645 358 5679
rect 392 5645 778 5679
rect 812 5645 1198 5679
rect 1232 5645 1458 5679
rect -2174 5639 -2116 5645
rect -1754 5639 -1696 5645
rect -1334 5639 -1276 5645
rect -914 5639 -856 5645
rect -494 5639 -436 5645
rect -74 5639 -16 5645
rect 346 5639 404 5645
rect 766 5639 824 5645
rect 1186 5639 1244 5645
rect 1448 5634 1458 5645
rect 1510 5679 1520 5686
rect 1606 5679 1664 5685
rect 2026 5679 2084 5685
rect 2446 5679 2504 5685
rect 2866 5679 2924 5685
rect 3286 5679 3344 5685
rect 3706 5679 3764 5685
rect 4126 5679 4184 5685
rect 4546 5679 4604 5685
rect 4966 5679 5024 5685
rect 5386 5679 5444 5685
rect 5806 5679 5864 5685
rect 1510 5645 1618 5679
rect 1652 5645 2038 5679
rect 2072 5645 2458 5679
rect 2492 5645 2878 5679
rect 2912 5645 3298 5679
rect 3332 5645 3718 5679
rect 3752 5645 4138 5679
rect 4172 5645 4558 5679
rect 4592 5645 4978 5679
rect 5012 5645 5398 5679
rect 5432 5645 5818 5679
rect 5852 5645 5900 5679
rect 1510 5634 1520 5645
rect 1606 5639 1664 5645
rect 2026 5639 2084 5645
rect 2446 5639 2504 5645
rect 2866 5639 2924 5645
rect 3286 5639 3344 5645
rect 3706 5639 3764 5645
rect 4126 5639 4184 5645
rect 4546 5639 4604 5645
rect 4966 5639 5024 5645
rect 5386 5639 5444 5645
rect 5806 5639 5864 5645
rect 1448 5555 1458 5558
rect -2384 5549 -2326 5555
rect -1964 5549 -1906 5555
rect -1544 5549 -1486 5555
rect -1124 5549 -1066 5555
rect -704 5549 -646 5555
rect -284 5549 -226 5555
rect 136 5549 194 5555
rect 556 5549 614 5555
rect 976 5549 1034 5555
rect 1396 5549 1458 5555
rect -2432 5515 -2372 5549
rect -2338 5515 -1952 5549
rect -1918 5515 -1532 5549
rect -1498 5515 -1112 5549
rect -1078 5515 -692 5549
rect -658 5515 -272 5549
rect -238 5515 148 5549
rect 182 5515 568 5549
rect 602 5515 988 5549
rect 1022 5515 1408 5549
rect 1442 5515 1458 5549
rect -2384 5509 -2326 5515
rect -1964 5509 -1906 5515
rect -1544 5509 -1486 5515
rect -1124 5509 -1066 5515
rect -704 5509 -646 5515
rect -284 5509 -226 5515
rect 136 5509 194 5515
rect 556 5509 614 5515
rect 976 5509 1034 5515
rect 1396 5509 1458 5515
rect 1448 5506 1458 5509
rect 1510 5549 1520 5558
rect 1816 5549 1874 5555
rect 2236 5549 2294 5555
rect 2656 5549 2714 5555
rect 3076 5549 3134 5555
rect 3496 5549 3554 5555
rect 3916 5549 3974 5555
rect 4336 5549 4394 5555
rect 4756 5549 4814 5555
rect 5176 5549 5234 5555
rect 5596 5549 5654 5555
rect 1510 5515 1828 5549
rect 1862 5515 2248 5549
rect 2282 5515 2668 5549
rect 2702 5515 3088 5549
rect 3122 5515 3508 5549
rect 3542 5515 3928 5549
rect 3962 5515 4348 5549
rect 4382 5515 4768 5549
rect 4802 5515 5188 5549
rect 5222 5515 5608 5549
rect 5642 5515 5900 5549
rect 1510 5506 1520 5515
rect 1816 5509 1874 5515
rect 2236 5509 2294 5515
rect 2656 5509 2714 5515
rect 3076 5509 3134 5515
rect 3496 5509 3554 5515
rect 3916 5509 3974 5515
rect 4336 5509 4394 5515
rect 4756 5509 4814 5515
rect 5176 5509 5234 5515
rect 5596 5509 5654 5515
rect -2432 5465 -2374 5471
rect -2222 5465 -2164 5471
rect -2012 5465 -1954 5471
rect -1802 5465 -1744 5471
rect -1592 5465 -1534 5471
rect -1382 5465 -1324 5471
rect -1172 5465 -1114 5471
rect -962 5465 -904 5471
rect -752 5465 -694 5471
rect -542 5465 -484 5471
rect -332 5465 -274 5471
rect -122 5465 -64 5471
rect 88 5465 146 5471
rect 298 5465 356 5471
rect 508 5465 566 5471
rect 718 5465 776 5471
rect 928 5465 986 5471
rect 1138 5465 1196 5471
rect 1348 5465 1406 5471
rect 1558 5465 1616 5471
rect 1768 5465 1826 5471
rect 1978 5465 2036 5471
rect 2188 5465 2246 5471
rect 2398 5465 2456 5471
rect 2608 5465 2666 5471
rect 2818 5465 2876 5471
rect 3028 5465 3086 5471
rect 3238 5465 3296 5471
rect 3448 5465 3506 5471
rect 3658 5465 3716 5471
rect 3868 5465 3926 5471
rect 4078 5465 4136 5471
rect 4288 5465 4346 5471
rect 4498 5465 4556 5471
rect 4708 5465 4766 5471
rect 4918 5465 4976 5471
rect 5128 5465 5186 5471
rect 5338 5465 5396 5471
rect 5548 5465 5606 5471
rect 5758 5465 5816 5471
rect -2432 5431 -2420 5465
rect -2386 5431 -2210 5465
rect -2176 5431 -2000 5465
rect -1966 5431 -1790 5465
rect -1756 5431 -1580 5465
rect -1546 5431 -1379 5465
rect -1327 5431 -1160 5465
rect -1126 5431 -950 5465
rect -916 5431 -740 5465
rect -706 5431 -530 5465
rect -496 5431 -320 5465
rect -286 5431 -110 5465
rect -76 5431 100 5465
rect 134 5431 301 5465
rect 353 5431 520 5465
rect 554 5431 730 5465
rect 764 5431 940 5465
rect 974 5431 1150 5465
rect 1184 5431 1360 5465
rect 1394 5431 1570 5465
rect 1604 5431 1780 5465
rect 1814 5431 1990 5465
rect 2024 5431 2200 5465
rect 2234 5431 2410 5465
rect 2444 5431 2620 5465
rect 2654 5431 2830 5465
rect 2864 5431 3040 5465
rect 3074 5431 3250 5465
rect 3284 5431 3460 5465
rect 3494 5431 3670 5465
rect 3704 5431 3880 5465
rect 3914 5431 4090 5465
rect 4124 5431 4300 5465
rect 4334 5431 4510 5465
rect 4544 5431 4720 5465
rect 4754 5431 4930 5465
rect 4964 5431 5140 5465
rect 5174 5431 5350 5465
rect 5384 5431 5560 5465
rect 5594 5431 5770 5465
rect 5804 5431 5912 5465
rect -2432 5425 -2374 5431
rect -2222 5425 -2164 5431
rect -2012 5425 -1954 5431
rect -1802 5425 -1744 5431
rect -1592 5425 -1534 5431
rect -1389 5413 -1379 5431
rect -1327 5413 -1317 5431
rect -1172 5425 -1114 5431
rect -962 5425 -904 5431
rect -752 5425 -694 5431
rect -542 5425 -484 5431
rect -332 5425 -274 5431
rect -122 5425 -64 5431
rect 88 5425 146 5431
rect 291 5413 301 5431
rect 353 5413 363 5431
rect 508 5425 566 5431
rect 718 5425 776 5431
rect 928 5425 986 5431
rect 1138 5425 1196 5431
rect 1348 5425 1406 5431
rect 1558 5425 1616 5431
rect 1768 5425 1826 5431
rect 1978 5425 2036 5431
rect 2188 5425 2246 5431
rect 2398 5425 2456 5431
rect 2608 5425 2666 5431
rect 2818 5425 2876 5431
rect 3028 5425 3086 5431
rect 3238 5425 3296 5431
rect 3448 5425 3506 5431
rect 3658 5425 3716 5431
rect 3868 5425 3926 5431
rect 4078 5425 4136 5431
rect 4288 5425 4346 5431
rect 4498 5425 4556 5431
rect 4708 5425 4766 5431
rect 4918 5425 4976 5431
rect 5128 5425 5186 5431
rect 5338 5425 5396 5431
rect 5548 5425 5606 5431
rect 5758 5425 5816 5431
rect -2336 5323 -2278 5329
rect -2126 5323 -2068 5329
rect -2019 5323 -2009 5341
rect -2432 5289 -2324 5323
rect -2290 5289 -2114 5323
rect -2080 5289 -2009 5323
rect -1957 5323 -1947 5341
rect -1916 5323 -1858 5329
rect -1706 5323 -1648 5329
rect -1496 5323 -1438 5329
rect -1286 5323 -1228 5329
rect -1076 5323 -1018 5329
rect -866 5323 -808 5329
rect -656 5323 -598 5329
rect -549 5323 -539 5341
rect -1957 5289 -1904 5323
rect -1870 5289 -1694 5323
rect -1660 5289 -1484 5323
rect -1450 5289 -1274 5323
rect -1240 5289 -1064 5323
rect -1030 5289 -854 5323
rect -820 5289 -644 5323
rect -610 5289 -539 5323
rect -487 5323 -477 5341
rect -446 5323 -388 5329
rect -236 5323 -178 5329
rect -26 5323 32 5329
rect 184 5323 242 5329
rect 394 5323 452 5329
rect 604 5323 662 5329
rect 814 5323 872 5329
rect 921 5323 931 5341
rect -487 5289 -434 5323
rect -400 5289 -224 5323
rect -190 5289 -14 5323
rect 20 5289 196 5323
rect 230 5289 406 5323
rect 440 5289 616 5323
rect 650 5289 826 5323
rect 860 5289 931 5323
rect 983 5323 993 5341
rect 1024 5323 1082 5329
rect 1234 5323 1292 5329
rect 1444 5323 1502 5329
rect 1654 5323 1712 5329
rect 1864 5323 1922 5329
rect 2074 5323 2132 5329
rect 2284 5323 2342 5329
rect 2494 5323 2552 5329
rect 2704 5323 2762 5329
rect 2914 5323 2972 5329
rect 3124 5323 3182 5329
rect 3334 5323 3392 5329
rect 3544 5323 3602 5329
rect 3754 5323 3812 5329
rect 3964 5323 4022 5329
rect 4174 5323 4232 5329
rect 4384 5323 4442 5329
rect 4594 5323 4652 5329
rect 4804 5323 4862 5329
rect 5014 5323 5072 5329
rect 5224 5323 5282 5329
rect 5434 5323 5492 5329
rect 5644 5323 5702 5329
rect 5854 5323 5912 5329
rect 983 5289 1036 5323
rect 1070 5289 1246 5323
rect 1280 5289 1456 5323
rect 1490 5289 1666 5323
rect 1700 5289 1876 5323
rect 1910 5289 2086 5323
rect 2120 5289 2296 5323
rect 2330 5289 2506 5323
rect 2540 5289 2716 5323
rect 2750 5289 2926 5323
rect 2960 5289 3136 5323
rect 3170 5289 3346 5323
rect 3380 5289 3556 5323
rect 3590 5289 3766 5323
rect 3800 5289 3976 5323
rect 4010 5289 4186 5323
rect 4220 5289 4396 5323
rect 4430 5289 4606 5323
rect 4640 5289 4816 5323
rect 4850 5289 5026 5323
rect 5060 5289 5236 5323
rect 5270 5289 5446 5323
rect 5480 5289 5656 5323
rect 5690 5289 5866 5323
rect 5900 5289 5912 5323
rect -2336 5283 -2278 5289
rect -2126 5283 -2068 5289
rect -1916 5283 -1858 5289
rect -1706 5283 -1648 5289
rect -1496 5283 -1438 5289
rect -1286 5283 -1228 5289
rect -1076 5283 -1018 5289
rect -866 5283 -808 5289
rect -656 5283 -598 5289
rect -446 5283 -388 5289
rect -236 5283 -178 5289
rect -26 5283 32 5289
rect 184 5283 242 5289
rect 394 5283 452 5289
rect 604 5283 662 5289
rect 814 5283 872 5289
rect 1024 5283 1082 5289
rect 1234 5283 1292 5289
rect 1444 5283 1502 5289
rect 1654 5283 1712 5289
rect 1864 5283 1922 5289
rect 2074 5283 2132 5289
rect 2284 5283 2342 5289
rect 2494 5283 2552 5289
rect 2704 5283 2762 5289
rect 2914 5283 2972 5289
rect 3124 5283 3182 5289
rect 3334 5283 3392 5289
rect 3544 5283 3602 5289
rect 3754 5283 3812 5289
rect 3964 5283 4022 5289
rect 4174 5283 4232 5289
rect 4384 5283 4442 5289
rect 4594 5283 4652 5289
rect 4804 5283 4862 5289
rect 5014 5283 5072 5289
rect 5224 5283 5282 5289
rect 5434 5283 5492 5289
rect 5644 5283 5702 5289
rect 5854 5283 5912 5289
rect -2174 5239 -2116 5245
rect -1754 5239 -1696 5245
rect -1334 5239 -1276 5245
rect -914 5239 -856 5245
rect -494 5239 -436 5245
rect -74 5239 -16 5245
rect 346 5239 404 5245
rect 766 5239 824 5245
rect 1186 5239 1244 5245
rect 1448 5239 1458 5245
rect -2432 5205 -2162 5239
rect -2128 5205 -1742 5239
rect -1708 5205 -1322 5239
rect -1288 5205 -902 5239
rect -868 5205 -482 5239
rect -448 5205 -62 5239
rect -28 5205 358 5239
rect 392 5205 778 5239
rect 812 5205 1198 5239
rect 1232 5205 1458 5239
rect -2174 5199 -2116 5205
rect -1754 5199 -1696 5205
rect -1334 5199 -1276 5205
rect -914 5199 -856 5205
rect -494 5199 -436 5205
rect -74 5199 -16 5205
rect 346 5199 404 5205
rect 766 5199 824 5205
rect 1186 5199 1244 5205
rect 1448 5193 1458 5205
rect 1510 5239 1520 5245
rect 1606 5239 1664 5245
rect 2026 5239 2084 5245
rect 2446 5239 2504 5245
rect 2866 5239 2924 5245
rect 3286 5239 3344 5245
rect 3706 5239 3764 5245
rect 4126 5239 4184 5245
rect 4546 5239 4604 5245
rect 4966 5239 5024 5245
rect 5386 5239 5444 5245
rect 5806 5239 5864 5245
rect 1510 5205 1618 5239
rect 1652 5205 2038 5239
rect 2072 5205 2458 5239
rect 2492 5205 2878 5239
rect 2912 5205 3298 5239
rect 3332 5205 3718 5239
rect 3752 5205 4138 5239
rect 4172 5205 4558 5239
rect 4592 5205 4978 5239
rect 5012 5205 5398 5239
rect 5432 5205 5818 5239
rect 5852 5205 5900 5239
rect 1510 5193 1520 5205
rect 1606 5199 1664 5205
rect 2026 5199 2084 5205
rect 2446 5199 2504 5205
rect 2866 5199 2924 5205
rect 3286 5199 3344 5205
rect 3706 5199 3764 5205
rect 4126 5199 4184 5205
rect 4546 5199 4604 5205
rect 4966 5199 5024 5205
rect 5386 5199 5444 5205
rect 5806 5199 5864 5205
rect -2384 5109 -2326 5115
rect -1964 5109 -1906 5115
rect -1544 5109 -1486 5115
rect -1124 5109 -1066 5115
rect -704 5109 -646 5115
rect -284 5109 -226 5115
rect 136 5109 194 5115
rect 556 5109 614 5115
rect 976 5109 1034 5115
rect 1396 5109 1454 5115
rect 1816 5109 1874 5115
rect 1960 5109 1970 5119
rect -2432 5075 -2372 5109
rect -2338 5075 -1952 5109
rect -1918 5075 -1532 5109
rect -1498 5075 -1112 5109
rect -1078 5075 -692 5109
rect -658 5075 -272 5109
rect -238 5075 148 5109
rect 182 5075 568 5109
rect 602 5075 988 5109
rect 1022 5075 1408 5109
rect 1442 5075 1828 5109
rect 1862 5075 1970 5109
rect -2384 5069 -2326 5075
rect -1964 5069 -1906 5075
rect -1544 5069 -1486 5075
rect -1124 5069 -1066 5075
rect -704 5069 -646 5075
rect -284 5069 -226 5075
rect 136 5069 194 5075
rect 556 5069 614 5075
rect 976 5069 1034 5075
rect 1396 5069 1454 5075
rect 1816 5069 1874 5075
rect 1960 5067 1970 5075
rect 2022 5109 2032 5119
rect 2236 5109 2294 5115
rect 2656 5109 2714 5115
rect 3076 5109 3134 5115
rect 3496 5109 3554 5115
rect 3916 5109 3974 5115
rect 4336 5109 4394 5115
rect 4756 5109 4814 5115
rect 5176 5109 5234 5115
rect 5596 5109 5654 5115
rect 2022 5075 2248 5109
rect 2282 5075 2668 5109
rect 2702 5075 3088 5109
rect 3122 5075 3508 5109
rect 3542 5075 3928 5109
rect 3962 5075 4348 5109
rect 4382 5075 4768 5109
rect 4802 5075 5188 5109
rect 5222 5075 5608 5109
rect 5642 5075 5900 5109
rect 2022 5067 2032 5075
rect 2236 5069 2294 5075
rect 2656 5069 2714 5075
rect 3076 5069 3134 5075
rect 3496 5069 3554 5075
rect 3916 5069 3974 5075
rect 4336 5069 4394 5075
rect 4756 5069 4814 5075
rect 5176 5069 5234 5075
rect 5596 5069 5654 5075
rect -2432 5025 -2374 5031
rect -2222 5025 -2164 5031
rect -2012 5025 -1954 5031
rect -1802 5025 -1744 5031
rect -1592 5025 -1534 5031
rect -1382 5025 -1324 5031
rect -1172 5025 -1114 5031
rect -962 5025 -904 5031
rect -752 5025 -694 5031
rect -542 5025 -484 5031
rect -332 5025 -274 5031
rect -122 5025 -64 5031
rect 88 5025 146 5031
rect 298 5025 356 5031
rect 508 5025 566 5031
rect 718 5025 776 5031
rect 928 5025 986 5031
rect 1138 5025 1196 5031
rect 1348 5025 1406 5031
rect 1558 5025 1616 5031
rect 1768 5025 1826 5031
rect 1978 5025 2036 5031
rect 2188 5025 2246 5031
rect 2398 5025 2456 5031
rect 2608 5025 2666 5031
rect 2818 5025 2876 5031
rect 3028 5025 3086 5031
rect 3238 5025 3296 5031
rect 3448 5025 3506 5031
rect 3658 5025 3716 5031
rect 3868 5025 3926 5031
rect 4078 5025 4136 5031
rect 4288 5025 4346 5031
rect 4498 5025 4556 5031
rect 4708 5025 4766 5031
rect 4918 5025 4976 5031
rect 5128 5025 5186 5031
rect 5338 5025 5396 5031
rect 5548 5025 5606 5031
rect 5758 5025 5816 5031
rect -2432 4991 -2420 5025
rect -2386 4991 -2210 5025
rect -2176 4991 -2000 5025
rect -1966 4991 -1790 5025
rect -1756 4991 -1580 5025
rect -1546 4991 -1370 5025
rect -1336 4991 -1160 5025
rect -1126 4991 -950 5025
rect -916 4991 -740 5025
rect -706 4991 -530 5025
rect -496 4991 -320 5025
rect -286 4991 -110 5025
rect -76 4991 100 5025
rect 134 4991 310 5025
rect 344 4991 520 5025
rect 554 4991 730 5025
rect 764 4991 940 5025
rect 974 4991 1150 5025
rect 1184 4991 1360 5025
rect 1394 4991 1570 5025
rect 1604 4991 1780 5025
rect 1814 4991 1990 5025
rect 2024 4991 2200 5025
rect 2234 4991 2410 5025
rect 2444 4991 2620 5025
rect 2654 4991 2830 5025
rect 2864 4991 3031 5025
rect 3083 4991 3250 5025
rect 3284 4991 3460 5025
rect 3494 4991 3670 5025
rect 3704 4991 3880 5025
rect 3914 4991 4090 5025
rect 4124 4991 4300 5025
rect 4334 4991 4510 5025
rect 4544 4991 4711 5025
rect 4763 4991 4930 5025
rect 4964 4991 5140 5025
rect 5174 4991 5350 5025
rect 5384 4991 5560 5025
rect 5594 4991 5770 5025
rect 5804 4991 5912 5025
rect -2432 4985 -2374 4991
rect -2222 4985 -2164 4991
rect -2012 4985 -1954 4991
rect -1802 4985 -1744 4991
rect -1592 4985 -1534 4991
rect -1382 4985 -1324 4991
rect -1172 4985 -1114 4991
rect -962 4985 -904 4991
rect -752 4985 -694 4991
rect -542 4985 -484 4991
rect -332 4985 -274 4991
rect -122 4985 -64 4991
rect 88 4985 146 4991
rect 298 4985 356 4991
rect 508 4985 566 4991
rect 718 4985 776 4991
rect 928 4985 986 4991
rect 1138 4985 1196 4991
rect 1348 4985 1406 4991
rect 1558 4985 1616 4991
rect 1768 4985 1826 4991
rect 1978 4985 2036 4991
rect 2188 4985 2246 4991
rect 2398 4985 2456 4991
rect 2608 4985 2666 4991
rect 2818 4985 2876 4991
rect 3021 4973 3031 4991
rect 3083 4973 3093 4991
rect 3238 4985 3296 4991
rect 3448 4985 3506 4991
rect 3658 4985 3716 4991
rect 3868 4985 3926 4991
rect 4078 4985 4136 4991
rect 4288 4985 4346 4991
rect 4498 4985 4556 4991
rect 4701 4973 4711 4991
rect 4763 4973 4773 4991
rect 4918 4985 4976 4991
rect 5128 4985 5186 4991
rect 5338 4985 5396 4991
rect 5548 4985 5606 4991
rect 5758 4985 5816 4991
rect -2336 4883 -2278 4889
rect -2126 4883 -2068 4889
rect -1916 4883 -1858 4889
rect -1706 4883 -1648 4889
rect -1496 4883 -1438 4889
rect -1286 4883 -1228 4889
rect -1076 4883 -1018 4889
rect -866 4883 -808 4889
rect -656 4883 -598 4889
rect -446 4883 -388 4889
rect -236 4883 -178 4889
rect -26 4883 32 4889
rect 184 4883 242 4889
rect 394 4883 452 4889
rect 604 4883 662 4889
rect 814 4883 872 4889
rect 1024 4883 1082 4889
rect 1234 4883 1292 4889
rect 1444 4883 1502 4889
rect 1654 4883 1712 4889
rect 1864 4883 1922 4889
rect 2074 4883 2132 4889
rect 2284 4883 2342 4889
rect 2391 4883 2401 4901
rect -2432 4849 -2324 4883
rect -2290 4849 -2114 4883
rect -2080 4849 -1904 4883
rect -1870 4849 -1694 4883
rect -1660 4849 -1484 4883
rect -1450 4849 -1274 4883
rect -1240 4849 -1064 4883
rect -1030 4849 -854 4883
rect -820 4849 -644 4883
rect -610 4849 -434 4883
rect -400 4849 -224 4883
rect -190 4849 -14 4883
rect 20 4849 196 4883
rect 230 4849 406 4883
rect 440 4849 616 4883
rect 650 4849 826 4883
rect 860 4849 1036 4883
rect 1070 4849 1246 4883
rect 1280 4849 1456 4883
rect 1490 4849 1666 4883
rect 1700 4849 1876 4883
rect 1910 4849 2086 4883
rect 2120 4849 2296 4883
rect 2330 4849 2401 4883
rect 2453 4883 2463 4901
rect 2494 4883 2552 4889
rect 2704 4883 2762 4889
rect 2914 4883 2972 4889
rect 3124 4883 3182 4889
rect 3334 4883 3392 4889
rect 3544 4883 3602 4889
rect 3754 4883 3812 4889
rect 3861 4883 3871 4901
rect 2453 4849 2506 4883
rect 2540 4849 2716 4883
rect 2750 4849 2926 4883
rect 2960 4849 3136 4883
rect 3170 4849 3346 4883
rect 3380 4849 3556 4883
rect 3590 4849 3766 4883
rect 3800 4849 3871 4883
rect 3923 4883 3933 4901
rect 3964 4883 4022 4889
rect 4174 4883 4232 4889
rect 4384 4883 4442 4889
rect 4594 4883 4652 4889
rect 4804 4883 4862 4889
rect 5014 4883 5072 4889
rect 5224 4883 5282 4889
rect 5330 4883 5340 4901
rect 3923 4849 3976 4883
rect 4010 4849 4186 4883
rect 4220 4849 4396 4883
rect 4430 4849 4606 4883
rect 4640 4849 4816 4883
rect 4850 4849 5026 4883
rect 5060 4849 5236 4883
rect 5270 4849 5340 4883
rect 5392 4883 5402 4901
rect 5434 4883 5492 4889
rect 5644 4883 5702 4889
rect 5854 4883 5912 4889
rect 5392 4849 5446 4883
rect 5480 4849 5656 4883
rect 5690 4849 5866 4883
rect 5900 4849 5912 4883
rect -2336 4843 -2278 4849
rect -2126 4843 -2068 4849
rect -1916 4843 -1858 4849
rect -1706 4843 -1648 4849
rect -1496 4843 -1438 4849
rect -1286 4843 -1228 4849
rect -1076 4843 -1018 4849
rect -866 4843 -808 4849
rect -656 4843 -598 4849
rect -446 4843 -388 4849
rect -236 4843 -178 4849
rect -26 4843 32 4849
rect 184 4843 242 4849
rect 394 4843 452 4849
rect 604 4843 662 4849
rect 814 4843 872 4849
rect 1024 4843 1082 4849
rect 1234 4843 1292 4849
rect 1444 4843 1502 4849
rect 1654 4843 1712 4849
rect 1864 4843 1922 4849
rect 2074 4843 2132 4849
rect 2284 4843 2342 4849
rect 2494 4843 2552 4849
rect 2704 4843 2762 4849
rect 2914 4843 2972 4849
rect 3124 4843 3182 4849
rect 3334 4843 3392 4849
rect 3544 4843 3602 4849
rect 3754 4843 3812 4849
rect 3964 4843 4022 4849
rect 4174 4843 4232 4849
rect 4384 4843 4442 4849
rect 4594 4843 4652 4849
rect 4804 4843 4862 4849
rect 5014 4843 5072 4849
rect 5224 4843 5282 4849
rect 5434 4843 5492 4849
rect 5644 4843 5702 4849
rect 5854 4843 5912 4849
rect -2174 4799 -2116 4805
rect -1754 4799 -1696 4805
rect -1334 4799 -1276 4805
rect -914 4799 -856 4805
rect -494 4799 -436 4805
rect -74 4799 -16 4805
rect 346 4799 404 4805
rect 766 4799 824 4805
rect 1186 4799 1244 4805
rect 1606 4799 1664 4805
rect 1960 4799 1970 4808
rect -2432 4765 -2162 4799
rect -2128 4765 -1742 4799
rect -1708 4765 -1322 4799
rect -1288 4765 -902 4799
rect -868 4765 -482 4799
rect -448 4765 -62 4799
rect -28 4765 358 4799
rect 392 4765 778 4799
rect 812 4765 1198 4799
rect 1232 4765 1618 4799
rect 1652 4765 1970 4799
rect -2174 4759 -2116 4765
rect -1754 4759 -1696 4765
rect -1334 4759 -1276 4765
rect -914 4759 -856 4765
rect -494 4759 -436 4765
rect -74 4759 -16 4765
rect 346 4759 404 4765
rect 766 4759 824 4765
rect 1186 4759 1244 4765
rect 1606 4759 1664 4765
rect -2845 4747 -2704 4759
rect 1960 4756 1970 4765
rect 2022 4805 2032 4808
rect 2022 4799 2084 4805
rect 2446 4799 2504 4805
rect 2866 4799 2924 4805
rect 3286 4799 3344 4805
rect 3706 4799 3764 4805
rect 4126 4799 4184 4805
rect 4546 4799 4604 4805
rect 4966 4799 5024 4805
rect 5386 4799 5444 4805
rect 5806 4799 5864 4805
rect 2022 4765 2038 4799
rect 2072 4765 2458 4799
rect 2492 4765 2878 4799
rect 2912 4765 3298 4799
rect 3332 4765 3718 4799
rect 3752 4765 4138 4799
rect 4172 4765 4558 4799
rect 4592 4765 4978 4799
rect 5012 4765 5398 4799
rect 5432 4765 5818 4799
rect 5852 4765 5900 4799
rect 2022 4759 2084 4765
rect 2446 4759 2504 4765
rect 2866 4759 2924 4765
rect 3286 4759 3344 4765
rect 3706 4759 3764 4765
rect 4126 4759 4184 4765
rect 4546 4759 4604 4765
rect 4966 4759 5024 4765
rect 5386 4759 5444 4765
rect 5806 4759 5864 4765
rect 6186 4759 6192 6435
rect 6226 6412 6322 6435
rect 6226 6360 6229 6412
rect 6281 6360 6322 6412
rect 6226 6271 6322 6360
rect 6226 6219 6229 6271
rect 6281 6219 6322 6271
rect 6226 6130 6322 6219
rect 6226 6078 6229 6130
rect 6281 6078 6322 6130
rect 6226 5989 6322 6078
rect 6226 5937 6229 5989
rect 6281 5937 6322 5989
rect 6226 5848 6322 5937
rect 6226 5796 6229 5848
rect 6281 5796 6322 5848
rect 6226 5707 6322 5796
rect 6226 5655 6229 5707
rect 6281 5655 6322 5707
rect 6226 5566 6322 5655
rect 6226 5514 6229 5566
rect 6281 5514 6322 5566
rect 6226 5425 6322 5514
rect 6226 5373 6229 5425
rect 6281 5373 6322 5425
rect 6226 5284 6322 5373
rect 6226 5232 6229 5284
rect 6281 5232 6322 5284
rect 6226 5143 6322 5232
rect 6226 5091 6229 5143
rect 6281 5091 6322 5143
rect 6226 5002 6322 5091
rect 6226 4950 6229 5002
rect 6281 4950 6322 5002
rect 6226 4861 6322 4950
rect 6226 4809 6229 4861
rect 6281 4809 6322 4861
rect 6226 4759 6322 4809
rect 2022 4756 2032 4759
rect 6186 4747 6322 4759
rect 6612 6073 6682 7983
rect 6831 7813 6889 7819
rect 6750 7778 6784 7781
rect 6831 7779 6843 7813
rect 6877 7779 6889 7813
rect 6744 7766 6790 7778
rect 6831 7773 6889 7779
rect 6744 7732 6750 7766
rect 6784 7732 6790 7766
rect 6744 7720 6790 7732
rect 6750 7586 6784 7720
rect 6843 7627 6877 7773
rect 6985 7723 7019 7983
rect 6973 7717 7031 7723
rect 6973 7683 6985 7717
rect 7019 7683 7031 7717
rect 6973 7677 7031 7683
rect 7078 7682 7112 7685
rect 6831 7621 6889 7627
rect 6831 7587 6843 7621
rect 6877 7587 6889 7621
rect 6744 7581 6790 7586
rect 6831 7581 6889 7587
rect 6731 7529 6741 7581
rect 6793 7529 6803 7581
rect 6744 7528 6790 7529
rect 6750 7394 6784 7528
rect 6843 7435 6877 7581
rect 6985 7531 7019 7677
rect 7072 7670 7118 7682
rect 7072 7636 7078 7670
rect 7112 7636 7118 7670
rect 7072 7624 7118 7636
rect 7078 7581 7112 7624
rect 6973 7525 7031 7531
rect 7062 7529 7072 7581
rect 7124 7529 7134 7581
rect 6973 7491 6985 7525
rect 7019 7491 7031 7525
rect 6973 7485 7031 7491
rect 7078 7490 7112 7529
rect 6831 7429 6889 7435
rect 6831 7395 6843 7429
rect 6877 7395 6889 7429
rect 6744 7382 6790 7394
rect 6831 7389 6889 7395
rect 6744 7348 6750 7382
rect 6784 7348 6790 7382
rect 6744 7336 6790 7348
rect 6750 7202 6784 7336
rect 6843 7243 6877 7389
rect 6985 7339 7019 7485
rect 7072 7478 7118 7490
rect 7072 7444 7078 7478
rect 7112 7444 7118 7478
rect 7072 7432 7118 7444
rect 6973 7333 7031 7339
rect 6973 7299 6985 7333
rect 7019 7299 7031 7333
rect 6973 7293 7031 7299
rect 7078 7298 7112 7432
rect 6831 7237 6889 7243
rect 6831 7203 6843 7237
rect 6877 7203 6889 7237
rect 6744 7190 6790 7202
rect 6831 7197 6889 7203
rect 6744 7156 6750 7190
rect 6784 7156 6790 7190
rect 6744 7144 6790 7156
rect 6750 7010 6784 7144
rect 6843 7051 6877 7197
rect 6985 7147 7019 7293
rect 7072 7286 7118 7298
rect 7072 7252 7078 7286
rect 7112 7252 7118 7286
rect 7072 7240 7118 7252
rect 6973 7141 7031 7147
rect 6973 7107 6985 7141
rect 7019 7107 7031 7141
rect 6973 7101 7031 7107
rect 7078 7106 7112 7240
rect 6831 7045 6889 7051
rect 6831 7011 6843 7045
rect 6877 7011 6889 7045
rect 6744 6998 6790 7010
rect 6831 7005 6889 7011
rect 6744 6964 6750 6998
rect 6784 6964 6790 6998
rect 6744 6952 6790 6964
rect 6750 6818 6784 6952
rect 6843 6859 6877 7005
rect 6985 6955 7019 7101
rect 7072 7094 7118 7106
rect 7072 7060 7078 7094
rect 7112 7060 7118 7094
rect 7072 7048 7118 7060
rect 6973 6949 7031 6955
rect 6973 6915 6985 6949
rect 7019 6915 7031 6949
rect 6973 6909 7031 6915
rect 7078 6914 7112 7048
rect 6831 6853 6889 6859
rect 6831 6819 6843 6853
rect 6877 6819 6889 6853
rect 6744 6806 6790 6818
rect 6831 6813 6889 6819
rect 6744 6772 6750 6806
rect 6784 6772 6790 6806
rect 6744 6760 6790 6772
rect 6750 6626 6784 6760
rect 6843 6720 6877 6813
rect 6985 6763 7019 6909
rect 7072 6902 7118 6914
rect 7072 6868 7078 6902
rect 7112 6868 7118 6902
rect 7072 6856 7118 6868
rect 6973 6757 7031 6763
rect 6973 6723 6985 6757
rect 7019 6723 7031 6757
rect 6823 6668 6833 6720
rect 6885 6668 6895 6720
rect 6973 6717 7031 6723
rect 7078 6722 7112 6856
rect 6831 6661 6889 6668
rect 6831 6627 6843 6661
rect 6877 6627 6889 6661
rect 6744 6614 6790 6626
rect 6831 6621 6889 6627
rect 6744 6580 6750 6614
rect 6784 6580 6790 6614
rect 6744 6568 6790 6580
rect 6750 6434 6784 6568
rect 6843 6475 6877 6621
rect 6985 6571 7019 6717
rect 7072 6710 7118 6722
rect 7072 6676 7078 6710
rect 7112 6676 7118 6710
rect 7072 6664 7118 6676
rect 6973 6565 7031 6571
rect 6973 6531 6985 6565
rect 7019 6531 7031 6565
rect 6973 6525 7031 6531
rect 7078 6530 7112 6664
rect 6831 6469 6889 6475
rect 6831 6435 6843 6469
rect 6877 6435 6889 6469
rect 6744 6431 6790 6434
rect 6731 6379 6741 6431
rect 6793 6379 6803 6431
rect 6831 6429 6889 6435
rect 6744 6376 6790 6379
rect 6750 6371 6784 6376
rect 6843 6283 6877 6429
rect 6985 6379 7019 6525
rect 7072 6518 7118 6530
rect 7072 6484 7078 6518
rect 7112 6484 7118 6518
rect 7072 6472 7118 6484
rect 7078 6431 7112 6472
rect 7060 6379 7070 6431
rect 7122 6379 7132 6431
rect 6973 6373 7031 6379
rect 6973 6339 6985 6373
rect 7019 6339 7031 6373
rect 6973 6333 7031 6339
rect 7078 6338 7112 6379
rect 6831 6277 6889 6283
rect 6831 6243 6843 6277
rect 6877 6243 6889 6277
rect 6831 6237 6889 6243
rect 6985 6073 7019 6333
rect 7072 6326 7118 6338
rect 7072 6292 7078 6326
rect 7112 6292 7118 6326
rect 7072 6280 7118 6292
rect 7078 6275 7112 6280
rect 6612 6067 7130 6073
rect 6612 6033 6744 6067
rect 7118 6033 7130 6067
rect 6612 6027 7130 6033
rect 6612 5619 6682 6027
rect 6612 5613 7130 5619
rect 6612 5579 6744 5613
rect 7118 5579 7130 5613
rect 6612 5573 7130 5579
rect -3082 4445 -3072 4497
rect -3020 4445 -2009 4497
rect -1957 4445 -539 4497
rect -487 4445 931 4497
rect 983 4445 999 4497
rect 2391 4445 2401 4497
rect 2453 4445 3871 4497
rect 3923 4445 5340 4497
rect 5392 4445 6482 4497
rect 6534 4445 6544 4497
rect -3668 3657 -3150 3663
rect -3668 3623 -3656 3657
rect -3282 3623 -3150 3657
rect -3668 3617 -3150 3623
rect -3220 3587 -3150 3617
rect -2845 4180 -2704 4192
rect -2845 4144 -2744 4180
rect -2845 4092 -2798 4144
rect -2746 4092 -2744 4144
rect -2845 4003 -2744 4092
rect -2845 3951 -2798 4003
rect -2746 3951 -2744 4003
rect -2845 3862 -2744 3951
rect -2845 3810 -2798 3862
rect -2746 3810 -2744 3862
rect -2845 3721 -2744 3810
rect -2845 3669 -2798 3721
rect -2746 3669 -2744 3721
rect -2845 3580 -2744 3669
rect -2845 3528 -2798 3580
rect -2746 3528 -2744 3580
rect -2845 3439 -2744 3528
rect -2845 3387 -2798 3439
rect -2746 3387 -2744 3439
rect -2845 3298 -2744 3387
rect -2845 3246 -2798 3298
rect -2746 3246 -2744 3298
rect -2845 3157 -2744 3246
rect -2845 3105 -2798 3157
rect -2746 3105 -2744 3157
rect -2845 3016 -2744 3105
rect -2845 2964 -2798 3016
rect -2746 2964 -2744 3016
rect -2845 2875 -2744 2964
rect -2845 2823 -2798 2875
rect -2746 2823 -2744 2875
rect -2845 2734 -2744 2823
rect -2845 2682 -2798 2734
rect -2746 2682 -2744 2734
rect -2845 1549 -2744 2682
rect -2845 1497 -2798 1549
rect -2746 1497 -2744 1549
rect -2845 1408 -2744 1497
rect -2845 1356 -2798 1408
rect -2746 1356 -2744 1408
rect -2845 1267 -2744 1356
rect -2845 1215 -2798 1267
rect -2746 1215 -2744 1267
rect -2845 1126 -2744 1215
rect -2845 1074 -2798 1126
rect -2746 1074 -2744 1126
rect -2845 985 -2744 1074
rect -2845 933 -2798 985
rect -2746 933 -2744 985
rect -2845 844 -2744 933
rect -2845 792 -2798 844
rect -2746 792 -2744 844
rect -2845 745 -2744 792
rect -2710 745 -2704 4180
rect -2598 4131 -2588 4183
rect -2536 4174 -2526 4183
rect -2391 4174 -2319 4183
rect -1964 4174 -1906 4180
rect -1551 4174 -1479 4183
rect -1124 4174 -1066 4180
rect -711 4174 -639 4183
rect -284 4174 -226 4180
rect 129 4174 201 4183
rect 556 4174 614 4180
rect 969 4174 1041 4183
rect 6186 4180 6322 4192
rect 1396 4174 1454 4180
rect 1816 4174 1874 4180
rect 2236 4174 2294 4180
rect 2656 4174 2714 4180
rect 3076 4174 3134 4180
rect 3496 4174 3554 4180
rect 3916 4174 3974 4180
rect 4336 4174 4394 4180
rect 4756 4174 4814 4180
rect 5176 4174 5234 4180
rect 5596 4174 5654 4180
rect -2536 4140 -2372 4174
rect -2338 4140 -1952 4174
rect -1918 4140 -1532 4174
rect -1498 4140 -1112 4174
rect -1078 4140 -692 4174
rect -658 4140 -272 4174
rect -238 4140 148 4174
rect 182 4140 568 4174
rect 602 4140 988 4174
rect 1022 4140 1408 4174
rect 1442 4140 1828 4174
rect 1862 4140 2248 4174
rect 2282 4140 2668 4174
rect 2702 4140 3088 4174
rect 3122 4140 3508 4174
rect 3542 4140 3928 4174
rect 3962 4140 4348 4174
rect 4382 4140 4768 4174
rect 4802 4140 5188 4174
rect 5222 4140 5608 4174
rect 5642 4140 5912 4174
rect -2536 4131 -2526 4140
rect -2391 4131 -2319 4140
rect -1964 4134 -1906 4140
rect -1551 4131 -1479 4140
rect -1124 4134 -1066 4140
rect -711 4131 -639 4140
rect -284 4134 -226 4140
rect 129 4131 201 4140
rect 556 4134 614 4140
rect 969 4131 1041 4140
rect 1396 4134 1454 4140
rect 1816 4134 1874 4140
rect 2236 4134 2294 4140
rect 2656 4134 2714 4140
rect 3076 4134 3134 4140
rect 3496 4134 3554 4140
rect 3916 4134 3974 4140
rect 4336 4134 4394 4140
rect 4756 4134 4814 4140
rect 5176 4134 5234 4140
rect 5596 4134 5654 4140
rect -2432 4090 -2374 4096
rect -2229 4090 -2157 4096
rect -2012 4090 -1954 4096
rect -1802 4090 -1744 4096
rect -1592 4090 -1534 4096
rect -1382 4090 -1324 4096
rect -1172 4090 -1114 4096
rect -962 4090 -904 4096
rect -752 4090 -694 4096
rect -549 4090 -539 4096
rect -487 4090 -477 4096
rect -332 4090 -274 4096
rect -122 4090 -64 4096
rect 88 4090 146 4096
rect 298 4090 356 4096
rect 508 4090 566 4096
rect 718 4090 776 4096
rect 928 4090 986 4096
rect 1138 4090 1196 4096
rect 1348 4090 1406 4096
rect 1558 4090 1616 4096
rect 1768 4090 1826 4096
rect 1978 4090 2036 4096
rect 2188 4090 2246 4096
rect 2398 4090 2456 4096
rect 2608 4090 2666 4096
rect 2818 4090 2876 4096
rect 3028 4090 3086 4096
rect 3238 4090 3296 4096
rect 3448 4090 3506 4096
rect 3658 4090 3716 4096
rect 3868 4090 3926 4096
rect 4078 4090 4136 4096
rect 4288 4090 4346 4096
rect 4498 4090 4556 4096
rect 4708 4090 4766 4096
rect 4918 4090 4976 4096
rect 5128 4090 5186 4096
rect 5338 4090 5396 4096
rect 5548 4090 5606 4096
rect 5758 4090 5816 4096
rect -2432 4056 -2420 4090
rect -2386 4056 -2210 4090
rect -2176 4056 -2009 4090
rect -1957 4056 -1790 4090
rect -1756 4056 -1580 4090
rect -1546 4056 -1370 4090
rect -1336 4056 -1160 4090
rect -1126 4056 -950 4090
rect -916 4056 -740 4090
rect -706 4056 -539 4090
rect -487 4056 -320 4090
rect -286 4056 -110 4090
rect -76 4056 100 4090
rect 134 4056 310 4090
rect 344 4056 520 4090
rect 554 4056 730 4090
rect 764 4056 931 4090
rect 983 4056 1150 4090
rect 1184 4056 1360 4090
rect 1394 4056 1570 4090
rect 1604 4056 1780 4090
rect 1814 4056 1990 4090
rect 2024 4056 2200 4090
rect 2234 4056 2410 4090
rect 2444 4056 2620 4090
rect 2654 4056 2830 4090
rect 2864 4056 3040 4090
rect 3074 4056 3250 4090
rect 3284 4056 3460 4090
rect 3494 4056 3670 4090
rect 3704 4056 3880 4090
rect 3914 4056 4090 4090
rect 4124 4056 4300 4090
rect 4334 4056 4510 4090
rect 4544 4056 4720 4090
rect 4754 4056 4930 4090
rect 4964 4056 5140 4090
rect 5174 4056 5350 4090
rect 5384 4056 5560 4090
rect 5594 4056 5770 4090
rect 5804 4056 5912 4090
rect -2432 4050 -2374 4056
rect -2229 4044 -2157 4056
rect -2019 4038 -2009 4056
rect -1957 4038 -1947 4056
rect -1802 4050 -1744 4056
rect -1592 4050 -1534 4056
rect -1382 4050 -1324 4056
rect -1172 4050 -1114 4056
rect -962 4050 -904 4056
rect -752 4050 -694 4056
rect -549 4044 -539 4056
rect -487 4044 -477 4056
rect -332 4050 -274 4056
rect -122 4050 -64 4056
rect 88 4050 146 4056
rect 298 4050 356 4056
rect 508 4050 566 4056
rect 718 4050 776 4056
rect 921 4038 931 4056
rect 983 4038 993 4056
rect 1138 4050 1196 4056
rect 1348 4050 1406 4056
rect 1558 4050 1616 4056
rect 1768 4050 1826 4056
rect 1978 4050 2036 4056
rect 2188 4050 2246 4056
rect 2398 4050 2456 4056
rect 2608 4050 2666 4056
rect 2818 4050 2876 4056
rect 3028 4050 3086 4056
rect 3238 4050 3296 4056
rect 3448 4050 3506 4056
rect 3658 4050 3716 4056
rect 3868 4050 3926 4056
rect 4078 4050 4136 4056
rect 4288 4050 4346 4056
rect 4498 4050 4556 4056
rect 4708 4050 4766 4056
rect 4918 4050 4976 4056
rect 5128 4050 5186 4056
rect 5338 4050 5396 4056
rect 5548 4050 5606 4056
rect 5758 4050 5816 4056
rect -2336 3948 -2278 3954
rect -2126 3948 -2068 3954
rect -1916 3948 -1858 3954
rect -1706 3948 -1648 3954
rect -1496 3948 -1438 3954
rect -1293 3948 -1283 3960
rect -1231 3948 -1221 3960
rect -1076 3948 -1018 3954
rect -866 3948 -808 3954
rect -656 3948 -598 3954
rect -446 3948 -388 3954
rect -236 3948 -178 3954
rect -26 3948 32 3954
rect 184 3948 242 3954
rect 292 3948 302 3960
rect -2432 3914 -2324 3948
rect -2290 3914 -2114 3948
rect -2080 3914 -1904 3948
rect -1870 3914 -1694 3948
rect -1660 3914 -1484 3948
rect -1450 3914 -1283 3948
rect -1231 3914 -1064 3948
rect -1030 3914 -854 3948
rect -820 3914 -644 3948
rect -610 3914 -434 3948
rect -400 3914 -224 3948
rect -190 3914 -14 3948
rect 20 3914 196 3948
rect 230 3914 302 3948
rect -2336 3908 -2278 3914
rect -2126 3908 -2068 3914
rect -1916 3908 -1858 3914
rect -1706 3908 -1648 3914
rect -1496 3908 -1438 3914
rect -1293 3908 -1283 3914
rect -1231 3908 -1221 3914
rect -1076 3908 -1018 3914
rect -866 3908 -808 3914
rect -656 3908 -598 3914
rect -446 3908 -388 3914
rect -236 3908 -178 3914
rect -26 3908 32 3914
rect 184 3908 242 3914
rect 292 3908 302 3914
rect 354 3948 364 3960
rect 394 3948 452 3954
rect 604 3948 662 3954
rect 814 3948 872 3954
rect 1024 3948 1082 3954
rect 1234 3948 1292 3954
rect 1444 3948 1502 3954
rect 1647 3948 1657 3960
rect 1709 3948 1719 3960
rect 1864 3948 1922 3954
rect 2074 3948 2132 3954
rect 2284 3948 2342 3954
rect 2494 3948 2552 3954
rect 2704 3948 2762 3954
rect 2907 3948 2917 3960
rect 2969 3948 2979 3960
rect 3124 3948 3182 3954
rect 3334 3948 3392 3954
rect 3544 3948 3602 3954
rect 3754 3948 3812 3954
rect 3964 3948 4022 3954
rect 4174 3948 4232 3954
rect 4384 3948 4442 3954
rect 4594 3948 4652 3954
rect 4804 3948 4862 3954
rect 4911 3948 4921 3960
rect 354 3914 406 3948
rect 440 3914 616 3948
rect 650 3914 826 3948
rect 860 3914 1036 3948
rect 1070 3914 1246 3948
rect 1280 3914 1456 3948
rect 1490 3914 1657 3948
rect 1709 3914 1876 3948
rect 1910 3914 2086 3948
rect 2120 3914 2296 3948
rect 2330 3914 2506 3948
rect 2540 3914 2716 3948
rect 2750 3914 2917 3948
rect 2969 3914 3136 3948
rect 3170 3914 3346 3948
rect 3380 3914 3556 3948
rect 3590 3914 3766 3948
rect 3800 3914 3976 3948
rect 4010 3914 4186 3948
rect 4220 3914 4396 3948
rect 4430 3914 4606 3948
rect 4640 3914 4816 3948
rect 4850 3914 4921 3948
rect 354 3908 364 3914
rect 394 3908 452 3914
rect 604 3908 662 3914
rect 814 3908 872 3914
rect 1024 3908 1082 3914
rect 1234 3908 1292 3914
rect 1444 3908 1502 3914
rect 1647 3908 1657 3914
rect 1709 3908 1719 3914
rect 1864 3908 1922 3914
rect 2074 3908 2132 3914
rect 2284 3908 2342 3914
rect 2494 3908 2552 3914
rect 2704 3908 2762 3914
rect 2907 3908 2917 3914
rect 2969 3908 2979 3914
rect 3124 3908 3182 3914
rect 3334 3908 3392 3914
rect 3544 3908 3602 3914
rect 3754 3908 3812 3914
rect 3964 3908 4022 3914
rect 4174 3908 4232 3914
rect 4384 3908 4442 3914
rect 4594 3908 4652 3914
rect 4804 3908 4862 3914
rect 4911 3908 4921 3914
rect 4973 3948 4983 3960
rect 5014 3948 5072 3954
rect 5224 3948 5282 3954
rect 5434 3948 5492 3954
rect 5644 3948 5702 3954
rect 5854 3948 5912 3954
rect 4973 3914 5026 3948
rect 5060 3914 5236 3948
rect 5270 3914 5446 3948
rect 5480 3914 5656 3948
rect 5690 3914 5866 3948
rect 5900 3914 5912 3948
rect 4973 3908 4983 3914
rect 5014 3908 5072 3914
rect 5224 3908 5282 3914
rect 5434 3908 5492 3914
rect 5644 3908 5702 3914
rect 5854 3908 5912 3914
rect -2598 3821 -2588 3873
rect -2536 3864 -2526 3873
rect -2181 3864 -2109 3873
rect -1754 3864 -1696 3870
rect -1341 3864 -1269 3873
rect -914 3864 -856 3870
rect -501 3864 -429 3873
rect -74 3864 -16 3870
rect 339 3864 411 3873
rect 766 3864 824 3870
rect 1179 3864 1251 3873
rect 1606 3864 1664 3870
rect 2026 3864 2084 3870
rect 2446 3864 2504 3870
rect 2866 3864 2924 3870
rect 3286 3864 3344 3870
rect 3706 3864 3764 3870
rect 4126 3864 4184 3870
rect 4546 3864 4604 3870
rect 4966 3864 5024 3870
rect 5386 3864 5444 3870
rect 5806 3864 5864 3870
rect -2536 3830 -2162 3864
rect -2128 3830 -1742 3864
rect -1708 3830 -1322 3864
rect -1288 3830 -902 3864
rect -868 3830 -482 3864
rect -448 3830 -62 3864
rect -28 3830 358 3864
rect 392 3830 778 3864
rect 812 3830 1198 3864
rect 1232 3830 1618 3864
rect 1652 3830 2038 3864
rect 2072 3830 2458 3864
rect 2492 3830 2878 3864
rect 2912 3830 3298 3864
rect 3332 3830 3718 3864
rect 3752 3830 4138 3864
rect 4172 3830 4558 3864
rect 4592 3830 4978 3864
rect 5012 3830 5398 3864
rect 5432 3830 5818 3864
rect 5852 3830 5912 3864
rect -2536 3821 -2526 3830
rect -2181 3821 -2109 3830
rect -1754 3824 -1696 3830
rect -1341 3821 -1269 3830
rect -914 3824 -856 3830
rect -501 3821 -429 3830
rect -74 3824 -16 3830
rect 339 3821 411 3830
rect 766 3824 824 3830
rect 1179 3821 1251 3830
rect 1606 3824 1664 3830
rect 2026 3824 2084 3830
rect 2446 3824 2504 3830
rect 2866 3824 2924 3830
rect 3286 3824 3344 3830
rect 3706 3824 3764 3830
rect 4126 3824 4184 3830
rect 4546 3824 4604 3830
rect 4966 3824 5024 3830
rect 5386 3824 5444 3830
rect 5806 3824 5864 3830
rect -2384 3734 -2326 3740
rect -1971 3734 -1899 3743
rect -1544 3734 -1486 3740
rect -1124 3734 -1066 3740
rect -704 3734 -646 3740
rect -291 3734 -219 3743
rect 136 3734 194 3740
rect 556 3734 614 3740
rect 976 3734 1034 3740
rect 1389 3734 1461 3743
rect 1816 3734 1874 3740
rect 2236 3734 2294 3740
rect 2656 3734 2714 3740
rect 3076 3734 3134 3740
rect 3496 3734 3554 3740
rect 3916 3734 3974 3740
rect 4336 3734 4394 3740
rect 4756 3734 4814 3740
rect 5176 3734 5234 3740
rect 5596 3734 5654 3740
rect 6010 3734 6020 3743
rect -2432 3700 -2372 3734
rect -2338 3700 -1952 3734
rect -1918 3700 -1532 3734
rect -1498 3700 -1112 3734
rect -1078 3700 -692 3734
rect -658 3700 -272 3734
rect -238 3700 148 3734
rect 182 3700 568 3734
rect 602 3700 988 3734
rect 1022 3700 1408 3734
rect 1442 3700 1828 3734
rect 1862 3700 2248 3734
rect 2282 3700 2668 3734
rect 2702 3700 3088 3734
rect 3122 3700 3508 3734
rect 3542 3700 3928 3734
rect 3962 3700 4348 3734
rect 4382 3700 4768 3734
rect 4802 3700 5188 3734
rect 5222 3700 5608 3734
rect 5642 3700 6020 3734
rect -2384 3694 -2326 3700
rect -1971 3691 -1899 3700
rect -1544 3694 -1486 3700
rect -1124 3694 -1066 3700
rect -704 3694 -646 3700
rect -291 3691 -219 3700
rect 136 3694 194 3700
rect 556 3694 614 3700
rect 976 3694 1034 3700
rect 1389 3691 1461 3700
rect 1816 3694 1874 3700
rect 2236 3694 2294 3700
rect 2656 3694 2714 3700
rect 3076 3694 3134 3700
rect 3496 3694 3554 3700
rect 3916 3694 3974 3700
rect 4336 3694 4394 3700
rect 4756 3694 4814 3700
rect 5176 3694 5234 3700
rect 5596 3694 5654 3700
rect 6010 3691 6020 3700
rect 6072 3691 6082 3743
rect -2432 3650 -2374 3656
rect -2222 3650 -2164 3656
rect -2012 3650 -1954 3656
rect -1802 3650 -1744 3656
rect -1592 3650 -1534 3656
rect -1382 3650 -1324 3656
rect -1172 3650 -1114 3656
rect -962 3650 -904 3656
rect -752 3650 -694 3656
rect -542 3650 -484 3656
rect -332 3650 -274 3656
rect -122 3650 -64 3656
rect 88 3650 146 3656
rect 298 3650 356 3656
rect 508 3650 566 3656
rect 718 3650 776 3656
rect 928 3650 986 3656
rect 1138 3650 1196 3656
rect 1348 3650 1406 3656
rect 1558 3650 1616 3656
rect 1768 3650 1826 3656
rect 1978 3650 2036 3656
rect 2188 3650 2246 3656
rect 2398 3650 2456 3656
rect 2608 3650 2666 3656
rect 2818 3650 2876 3656
rect 3028 3650 3086 3656
rect 3238 3650 3296 3656
rect 3448 3650 3506 3656
rect 3658 3650 3716 3656
rect 3868 3650 3926 3656
rect 4078 3650 4136 3656
rect 4288 3650 4346 3656
rect 4498 3650 4556 3656
rect 4708 3650 4766 3656
rect 4918 3650 4976 3656
rect 5128 3650 5186 3656
rect 5338 3650 5396 3656
rect 5548 3650 5606 3656
rect 5758 3650 5816 3656
rect -2432 3616 -2420 3650
rect -2386 3616 -2210 3650
rect -2176 3616 -2000 3650
rect -1966 3616 -1790 3650
rect -1756 3616 -1580 3650
rect -1546 3616 -1370 3650
rect -1336 3616 -1160 3650
rect -1126 3616 -950 3650
rect -916 3616 -740 3650
rect -706 3616 -530 3650
rect -496 3616 -320 3650
rect -286 3616 -110 3650
rect -76 3616 100 3650
rect 134 3616 310 3650
rect 344 3616 520 3650
rect 554 3616 730 3650
rect 764 3616 940 3650
rect 974 3616 1150 3650
rect 1184 3616 1360 3650
rect 1394 3616 1570 3650
rect 1604 3616 1780 3650
rect 1814 3616 1990 3650
rect 2024 3616 2200 3650
rect 2234 3616 2401 3650
rect 2453 3616 2620 3650
rect 2654 3616 2830 3650
rect 2864 3616 3040 3650
rect 3074 3616 3250 3650
rect 3284 3616 3460 3650
rect 3494 3616 3670 3650
rect 3704 3616 3871 3650
rect 3923 3616 4090 3650
rect 4124 3616 4300 3650
rect 4334 3616 4510 3650
rect 4544 3616 4720 3650
rect 4754 3616 4930 3650
rect 4964 3616 5140 3650
rect 5174 3616 5340 3650
rect 5392 3616 5560 3650
rect 5594 3616 5770 3650
rect 5804 3616 5912 3650
rect -2432 3610 -2374 3616
rect -2222 3610 -2164 3616
rect -2012 3610 -1954 3616
rect -1802 3610 -1744 3616
rect -1592 3610 -1534 3616
rect -1382 3610 -1324 3616
rect -1172 3610 -1114 3616
rect -962 3610 -904 3616
rect -752 3610 -694 3616
rect -542 3610 -484 3616
rect -332 3610 -274 3616
rect -122 3610 -64 3616
rect 88 3610 146 3616
rect 298 3610 356 3616
rect 508 3610 566 3616
rect 718 3610 776 3616
rect 928 3610 986 3616
rect 1138 3610 1196 3616
rect 1348 3610 1406 3616
rect 1558 3610 1616 3616
rect 1768 3610 1826 3616
rect 1978 3610 2036 3616
rect 2188 3610 2246 3616
rect 2391 3598 2401 3616
rect 2453 3598 2463 3616
rect 2608 3610 2666 3616
rect 2818 3610 2876 3616
rect 3028 3610 3086 3616
rect 3238 3610 3296 3616
rect 3448 3610 3506 3616
rect 3658 3610 3716 3616
rect 3861 3598 3871 3616
rect 3923 3598 3933 3616
rect 4078 3610 4136 3616
rect 4288 3610 4346 3616
rect 4498 3610 4556 3616
rect 4708 3610 4766 3616
rect 4918 3610 4976 3616
rect 5128 3610 5186 3616
rect 5330 3598 5340 3616
rect 5392 3598 5402 3616
rect 5548 3610 5606 3616
rect 5758 3610 5816 3616
rect -2336 3508 -2278 3514
rect -2126 3508 -2068 3514
rect -1916 3508 -1858 3514
rect -1706 3508 -1648 3514
rect -1496 3508 -1438 3514
rect -1293 3508 -1283 3520
rect -1231 3508 -1221 3520
rect -1076 3508 -1018 3514
rect -866 3508 -808 3514
rect -656 3508 -598 3514
rect -446 3508 -388 3514
rect -236 3508 -178 3514
rect -26 3508 32 3514
rect 184 3508 242 3514
rect 292 3508 302 3520
rect -2432 3474 -2324 3508
rect -2290 3474 -2114 3508
rect -2080 3474 -1904 3508
rect -1870 3474 -1694 3508
rect -1660 3474 -1484 3508
rect -1450 3474 -1283 3508
rect -1231 3474 -1064 3508
rect -1030 3474 -854 3508
rect -820 3474 -644 3508
rect -610 3474 -434 3508
rect -400 3474 -224 3508
rect -190 3474 -14 3508
rect 20 3474 196 3508
rect 230 3474 302 3508
rect -2336 3468 -2278 3474
rect -2126 3468 -2068 3474
rect -1916 3468 -1858 3474
rect -1706 3468 -1648 3474
rect -1496 3468 -1438 3474
rect -1293 3468 -1283 3474
rect -1231 3468 -1221 3474
rect -1076 3468 -1018 3474
rect -866 3468 -808 3474
rect -656 3468 -598 3474
rect -446 3468 -388 3474
rect -236 3468 -178 3474
rect -26 3468 32 3474
rect 184 3468 242 3474
rect 292 3468 302 3474
rect 354 3508 364 3520
rect 394 3508 452 3514
rect 604 3508 662 3514
rect 814 3508 872 3514
rect 1024 3508 1082 3514
rect 1234 3508 1292 3514
rect 1444 3508 1502 3514
rect 1647 3508 1657 3520
rect 1709 3508 1719 3520
rect 1864 3508 1922 3514
rect 2074 3508 2132 3514
rect 2284 3508 2342 3514
rect 2494 3508 2552 3514
rect 2704 3508 2762 3514
rect 2907 3508 2917 3520
rect 2969 3508 2979 3520
rect 3124 3508 3182 3514
rect 3334 3508 3392 3514
rect 3544 3508 3602 3514
rect 3754 3508 3812 3514
rect 3964 3508 4022 3514
rect 4174 3508 4232 3514
rect 4384 3508 4442 3514
rect 4594 3508 4652 3514
rect 4804 3508 4862 3514
rect 4911 3508 4921 3520
rect 354 3474 406 3508
rect 440 3474 616 3508
rect 650 3474 826 3508
rect 860 3474 1036 3508
rect 1070 3474 1246 3508
rect 1280 3474 1456 3508
rect 1490 3474 1657 3508
rect 1709 3474 1876 3508
rect 1910 3474 2086 3508
rect 2120 3474 2296 3508
rect 2330 3474 2506 3508
rect 2540 3474 2716 3508
rect 2750 3474 2917 3508
rect 2969 3474 3136 3508
rect 3170 3474 3346 3508
rect 3380 3474 3556 3508
rect 3590 3474 3766 3508
rect 3800 3474 3976 3508
rect 4010 3474 4186 3508
rect 4220 3474 4396 3508
rect 4430 3474 4606 3508
rect 4640 3474 4816 3508
rect 4850 3474 4921 3508
rect 354 3468 364 3474
rect 394 3468 452 3474
rect 604 3468 662 3474
rect 814 3468 872 3474
rect 1024 3468 1082 3474
rect 1234 3468 1292 3474
rect 1444 3468 1502 3474
rect 1647 3468 1657 3474
rect 1709 3468 1719 3474
rect 1864 3468 1922 3474
rect 2074 3468 2132 3474
rect 2284 3468 2342 3474
rect 2494 3468 2552 3474
rect 2704 3468 2762 3474
rect 2907 3468 2917 3474
rect 2969 3468 2979 3474
rect 3124 3468 3182 3474
rect 3334 3468 3392 3474
rect 3544 3468 3602 3474
rect 3754 3468 3812 3474
rect 3964 3468 4022 3474
rect 4174 3468 4232 3474
rect 4384 3468 4442 3474
rect 4594 3468 4652 3474
rect 4804 3468 4862 3474
rect 4911 3468 4921 3474
rect 4973 3508 4983 3520
rect 5014 3508 5072 3514
rect 5224 3508 5282 3514
rect 5434 3508 5492 3514
rect 5644 3508 5702 3514
rect 5854 3508 5912 3514
rect 4973 3474 5026 3508
rect 5060 3474 5236 3508
rect 5270 3474 5446 3508
rect 5480 3474 5656 3508
rect 5690 3474 5866 3508
rect 5900 3474 5912 3508
rect 4973 3468 4983 3474
rect 5014 3468 5072 3474
rect 5224 3468 5282 3474
rect 5434 3468 5492 3474
rect 5644 3468 5702 3474
rect 5854 3468 5912 3474
rect -2174 3424 -2116 3430
rect -1761 3424 -1689 3433
rect -1334 3424 -1276 3430
rect -914 3424 -856 3430
rect -494 3424 -436 3430
rect -81 3424 -9 3433
rect 346 3424 404 3430
rect 766 3424 824 3430
rect 1186 3424 1244 3430
rect 1599 3424 1671 3433
rect 2026 3424 2084 3430
rect 2446 3424 2504 3430
rect 2866 3424 2924 3430
rect 3286 3424 3344 3430
rect 3706 3424 3764 3430
rect 4126 3424 4184 3430
rect 4546 3424 4604 3430
rect 4966 3424 5024 3430
rect 5386 3424 5444 3430
rect 5806 3424 5864 3430
rect 6010 3424 6020 3433
rect -2432 3390 -2162 3424
rect -2128 3390 -1742 3424
rect -1708 3390 -1322 3424
rect -1288 3390 -902 3424
rect -868 3390 -482 3424
rect -448 3390 -62 3424
rect -28 3390 358 3424
rect 392 3390 778 3424
rect 812 3390 1198 3424
rect 1232 3390 1618 3424
rect 1652 3390 2038 3424
rect 2072 3390 2458 3424
rect 2492 3390 2878 3424
rect 2912 3390 3298 3424
rect 3332 3390 3718 3424
rect 3752 3390 4138 3424
rect 4172 3390 4558 3424
rect 4592 3390 4978 3424
rect 5012 3390 5398 3424
rect 5432 3390 5818 3424
rect 5852 3390 6020 3424
rect -2174 3384 -2116 3390
rect -1761 3381 -1689 3390
rect -1334 3384 -1276 3390
rect -914 3384 -856 3390
rect -494 3384 -436 3390
rect -81 3381 -9 3390
rect 346 3384 404 3390
rect 766 3384 824 3390
rect 1186 3384 1244 3390
rect 1599 3381 1671 3390
rect 2026 3384 2084 3390
rect 2446 3384 2504 3390
rect 2866 3384 2924 3390
rect 3286 3384 3344 3390
rect 3706 3384 3764 3390
rect 4126 3384 4184 3390
rect 4546 3384 4604 3390
rect 4966 3384 5024 3390
rect 5386 3384 5444 3390
rect 5806 3384 5864 3390
rect 6010 3381 6020 3390
rect 6072 3381 6082 3433
rect -2391 3294 -2319 3303
rect -1964 3294 -1906 3300
rect -1551 3294 -1479 3303
rect -1124 3294 -1066 3300
rect -711 3294 -639 3303
rect -284 3294 -226 3300
rect 129 3294 201 3303
rect 556 3294 614 3300
rect 969 3294 1041 3303
rect 1396 3294 1454 3300
rect 1816 3294 1874 3300
rect 2236 3294 2294 3300
rect 2656 3294 2714 3300
rect 3076 3294 3134 3300
rect 3496 3294 3554 3300
rect 3916 3294 3974 3300
rect 4336 3294 4394 3300
rect 4756 3294 4814 3300
rect 5176 3294 5234 3300
rect 5596 3294 5654 3300
rect 6010 3294 6020 3305
rect -2432 3260 -2372 3294
rect -2338 3260 -1952 3294
rect -1918 3260 -1532 3294
rect -1498 3260 -1112 3294
rect -1078 3260 -692 3294
rect -658 3260 -272 3294
rect -238 3260 148 3294
rect 182 3260 568 3294
rect 602 3260 988 3294
rect 1022 3260 1408 3294
rect 1442 3260 1828 3294
rect 1862 3260 2248 3294
rect 2282 3260 2668 3294
rect 2702 3260 3088 3294
rect 3122 3260 3508 3294
rect 3542 3260 3928 3294
rect 3962 3260 4348 3294
rect 4382 3260 4768 3294
rect 4802 3260 5188 3294
rect 5222 3260 5608 3294
rect 5642 3260 6020 3294
rect -2391 3251 -2319 3260
rect -1964 3254 -1906 3260
rect -1551 3251 -1479 3260
rect -1124 3254 -1066 3260
rect -711 3251 -639 3260
rect -284 3254 -226 3260
rect 129 3251 201 3260
rect 556 3254 614 3260
rect 969 3251 1041 3260
rect 1396 3254 1454 3260
rect 1816 3254 1874 3260
rect 2236 3254 2294 3260
rect 2656 3254 2714 3260
rect 3076 3254 3134 3260
rect 3496 3254 3554 3260
rect 3916 3254 3974 3260
rect 4336 3254 4394 3260
rect 4756 3254 4814 3260
rect 5176 3254 5234 3260
rect 5596 3254 5654 3260
rect 6010 3253 6020 3260
rect 6072 3253 6082 3305
rect -2432 3210 -2374 3216
rect -2222 3210 -2164 3216
rect -2012 3210 -1954 3216
rect -1802 3210 -1744 3216
rect -1592 3210 -1534 3216
rect -1382 3210 -1324 3216
rect -1172 3210 -1114 3216
rect -962 3210 -904 3216
rect -752 3210 -694 3216
rect -542 3210 -484 3216
rect -332 3210 -274 3216
rect -122 3210 -64 3216
rect 88 3210 146 3216
rect 298 3210 356 3216
rect 508 3210 566 3216
rect 718 3210 776 3216
rect 928 3210 986 3216
rect 1138 3210 1196 3216
rect 1348 3210 1406 3216
rect 1558 3210 1616 3216
rect 1768 3210 1826 3216
rect 1978 3210 2036 3216
rect 2188 3210 2246 3216
rect 2398 3210 2456 3216
rect 2608 3210 2666 3216
rect 2818 3210 2876 3216
rect 3028 3210 3086 3216
rect 3238 3210 3296 3216
rect 3448 3210 3506 3216
rect 3658 3210 3716 3216
rect 3868 3210 3926 3216
rect 4078 3210 4136 3216
rect 4288 3210 4346 3216
rect 4498 3210 4556 3216
rect 4708 3210 4766 3216
rect 4918 3210 4976 3216
rect 5128 3210 5186 3216
rect 5338 3210 5396 3216
rect 5548 3210 5606 3216
rect 5758 3210 5816 3216
rect -2432 3176 -2420 3210
rect -2386 3176 -2210 3210
rect -2176 3176 -2000 3210
rect -1966 3176 -1790 3210
rect -1756 3176 -1580 3210
rect -1546 3176 -1370 3210
rect -1336 3176 -1160 3210
rect -1126 3176 -950 3210
rect -916 3176 -740 3210
rect -706 3176 -530 3210
rect -496 3176 -320 3210
rect -286 3176 -110 3210
rect -76 3176 100 3210
rect 134 3176 310 3210
rect 344 3176 520 3210
rect 554 3176 730 3210
rect 764 3176 940 3210
rect 974 3176 1150 3210
rect 1184 3176 1360 3210
rect 1394 3176 1570 3210
rect 1604 3176 1780 3210
rect 1814 3176 1990 3210
rect 2024 3176 2200 3210
rect 2234 3176 2401 3210
rect 2453 3176 2620 3210
rect 2654 3176 2830 3210
rect 2864 3176 3040 3210
rect 3074 3176 3250 3210
rect 3284 3176 3460 3210
rect 3494 3176 3670 3210
rect 3704 3176 3871 3210
rect 3923 3176 4090 3210
rect 4124 3176 4300 3210
rect 4334 3176 4510 3210
rect 4544 3176 4720 3210
rect 4754 3176 4930 3210
rect 4964 3176 5140 3210
rect 5174 3176 5340 3210
rect 5392 3176 5560 3210
rect 5594 3176 5770 3210
rect 5804 3176 5912 3210
rect -2432 3170 -2374 3176
rect -2222 3170 -2164 3176
rect -2012 3170 -1954 3176
rect -1802 3170 -1744 3176
rect -1592 3170 -1534 3176
rect -1382 3170 -1324 3176
rect -1172 3170 -1114 3176
rect -962 3170 -904 3176
rect -752 3170 -694 3176
rect -542 3170 -484 3176
rect -332 3170 -274 3176
rect -122 3170 -64 3176
rect 88 3170 146 3176
rect 298 3170 356 3176
rect 508 3170 566 3176
rect 718 3170 776 3176
rect 928 3170 986 3176
rect 1138 3170 1196 3176
rect 1348 3170 1406 3176
rect 1558 3170 1616 3176
rect 1768 3170 1826 3176
rect 1978 3170 2036 3176
rect 2188 3170 2246 3176
rect 2391 3158 2401 3176
rect 2453 3158 2463 3176
rect 2608 3170 2666 3176
rect 2818 3170 2876 3176
rect 3028 3170 3086 3176
rect 3238 3170 3296 3176
rect 3448 3170 3506 3176
rect 3658 3170 3716 3176
rect 3861 3158 3871 3176
rect 3923 3158 3933 3176
rect 4078 3170 4136 3176
rect 4288 3170 4346 3176
rect 4498 3170 4556 3176
rect 4708 3170 4766 3176
rect 4918 3170 4976 3176
rect 5128 3170 5186 3176
rect 5330 3158 5340 3176
rect 5392 3158 5402 3176
rect 5548 3170 5606 3176
rect 5758 3170 5816 3176
rect -2336 3068 -2278 3074
rect -2126 3068 -2068 3074
rect -1916 3068 -1858 3074
rect -1706 3068 -1648 3074
rect -1496 3068 -1438 3074
rect -1293 3068 -1283 3080
rect -1231 3068 -1221 3080
rect -1076 3068 -1018 3074
rect -866 3068 -808 3074
rect -656 3068 -598 3074
rect -446 3068 -388 3074
rect -236 3068 -178 3074
rect -26 3068 32 3074
rect 184 3068 242 3074
rect 292 3068 302 3080
rect -2432 3034 -2324 3068
rect -2290 3034 -2114 3068
rect -2080 3034 -1904 3068
rect -1870 3034 -1694 3068
rect -1660 3034 -1484 3068
rect -1450 3034 -1283 3068
rect -1231 3034 -1064 3068
rect -1030 3034 -854 3068
rect -820 3034 -644 3068
rect -610 3034 -434 3068
rect -400 3034 -224 3068
rect -190 3034 -14 3068
rect 20 3034 196 3068
rect 230 3034 302 3068
rect -2336 3028 -2278 3034
rect -2126 3028 -2068 3034
rect -1916 3028 -1858 3034
rect -1706 3028 -1648 3034
rect -1496 3028 -1438 3034
rect -1293 3028 -1283 3034
rect -1231 3028 -1221 3034
rect -1076 3028 -1018 3034
rect -866 3028 -808 3034
rect -656 3028 -598 3034
rect -446 3028 -388 3034
rect -236 3028 -178 3034
rect -26 3028 32 3034
rect 184 3028 242 3034
rect 292 3028 302 3034
rect 354 3068 364 3080
rect 394 3068 452 3074
rect 604 3068 662 3074
rect 814 3068 872 3074
rect 1024 3068 1082 3074
rect 1234 3068 1292 3074
rect 1444 3068 1502 3074
rect 1647 3068 1657 3080
rect 1709 3068 1719 3080
rect 1864 3068 1922 3074
rect 2074 3068 2132 3074
rect 2284 3068 2342 3074
rect 2494 3068 2552 3074
rect 2704 3068 2762 3074
rect 2907 3068 2917 3080
rect 2969 3068 2979 3080
rect 3124 3068 3182 3074
rect 3334 3068 3392 3074
rect 3544 3068 3602 3074
rect 3754 3068 3812 3074
rect 3964 3068 4022 3074
rect 4174 3068 4232 3074
rect 4384 3068 4442 3074
rect 4594 3068 4652 3074
rect 4804 3068 4862 3074
rect 4911 3068 4921 3080
rect 354 3034 406 3068
rect 440 3034 616 3068
rect 650 3034 826 3068
rect 860 3034 1036 3068
rect 1070 3034 1246 3068
rect 1280 3034 1456 3068
rect 1490 3034 1657 3068
rect 1709 3034 1876 3068
rect 1910 3034 2086 3068
rect 2120 3034 2296 3068
rect 2330 3034 2506 3068
rect 2540 3034 2716 3068
rect 2750 3034 2917 3068
rect 2969 3034 3136 3068
rect 3170 3034 3346 3068
rect 3380 3034 3556 3068
rect 3590 3034 3766 3068
rect 3800 3034 3976 3068
rect 4010 3034 4186 3068
rect 4220 3034 4396 3068
rect 4430 3034 4606 3068
rect 4640 3034 4816 3068
rect 4850 3034 4921 3068
rect 354 3028 364 3034
rect 394 3028 452 3034
rect 604 3028 662 3034
rect 814 3028 872 3034
rect 1024 3028 1082 3034
rect 1234 3028 1292 3034
rect 1444 3028 1502 3034
rect 1647 3028 1657 3034
rect 1709 3028 1719 3034
rect 1864 3028 1922 3034
rect 2074 3028 2132 3034
rect 2284 3028 2342 3034
rect 2494 3028 2552 3034
rect 2704 3028 2762 3034
rect 2907 3028 2917 3034
rect 2969 3028 2979 3034
rect 3124 3028 3182 3034
rect 3334 3028 3392 3034
rect 3544 3028 3602 3034
rect 3754 3028 3812 3034
rect 3964 3028 4022 3034
rect 4174 3028 4232 3034
rect 4384 3028 4442 3034
rect 4594 3028 4652 3034
rect 4804 3028 4862 3034
rect 4911 3028 4921 3034
rect 4973 3068 4983 3080
rect 5014 3068 5072 3074
rect 5224 3068 5282 3074
rect 5434 3068 5492 3074
rect 5644 3068 5702 3074
rect 5854 3068 5912 3074
rect 4973 3034 5026 3068
rect 5060 3034 5236 3068
rect 5270 3034 5446 3068
rect 5480 3034 5656 3068
rect 5690 3034 5866 3068
rect 5900 3034 5912 3068
rect 4973 3028 4983 3034
rect 5014 3028 5072 3034
rect 5224 3028 5282 3034
rect 5434 3028 5492 3034
rect 5644 3028 5702 3034
rect 5854 3028 5912 3034
rect -2181 2984 -2109 2993
rect -1754 2984 -1696 2990
rect -1341 2984 -1269 2993
rect -914 2984 -856 2990
rect -501 2984 -429 2993
rect -74 2984 -16 2990
rect 339 2984 411 2993
rect 766 2984 824 2990
rect 1179 2984 1251 2993
rect 1606 2984 1664 2990
rect 2026 2984 2084 2990
rect 2446 2984 2504 2990
rect 2866 2984 2924 2990
rect 3286 2984 3344 2990
rect 3706 2984 3764 2990
rect 4126 2984 4184 2990
rect 4546 2984 4604 2990
rect 4966 2984 5024 2990
rect 5386 2984 5444 2990
rect 5806 2984 5864 2990
rect 6010 2984 6020 2991
rect -2432 2950 -2162 2984
rect -2128 2950 -1742 2984
rect -1708 2950 -1322 2984
rect -1288 2950 -902 2984
rect -868 2950 -482 2984
rect -448 2950 -62 2984
rect -28 2950 358 2984
rect 392 2950 778 2984
rect 812 2950 1198 2984
rect 1232 2950 1618 2984
rect 1652 2950 2038 2984
rect 2072 2950 2458 2984
rect 2492 2950 2878 2984
rect 2912 2950 3298 2984
rect 3332 2950 3718 2984
rect 3752 2950 4138 2984
rect 4172 2950 4558 2984
rect 4592 2950 4978 2984
rect 5012 2950 5398 2984
rect 5432 2950 5818 2984
rect 5852 2950 6020 2984
rect -2181 2941 -2109 2950
rect -1754 2944 -1696 2950
rect -1341 2941 -1269 2950
rect -914 2944 -856 2950
rect -501 2941 -429 2950
rect -74 2944 -16 2950
rect 339 2941 411 2950
rect 766 2944 824 2950
rect 1179 2941 1251 2950
rect 1606 2944 1664 2950
rect 2026 2944 2084 2950
rect 2446 2944 2504 2950
rect 2866 2944 2924 2950
rect 3286 2944 3344 2950
rect 3706 2944 3764 2950
rect 4126 2944 4184 2950
rect 4546 2944 4604 2950
rect 4966 2944 5024 2950
rect 5386 2944 5444 2950
rect 5806 2944 5864 2950
rect 6010 2939 6020 2950
rect 6072 2939 6082 2991
rect -2598 2811 -2588 2863
rect -2536 2854 -2526 2863
rect -2384 2854 -2326 2860
rect -1971 2854 -1899 2863
rect -1544 2854 -1486 2860
rect -1124 2854 -1066 2860
rect -704 2854 -646 2860
rect -291 2854 -219 2863
rect 136 2854 194 2860
rect 556 2854 614 2860
rect 976 2854 1034 2860
rect 1389 2854 1461 2863
rect 1816 2854 1874 2860
rect 2236 2854 2294 2860
rect 2656 2854 2714 2860
rect 3076 2854 3134 2860
rect 3496 2854 3554 2860
rect 3916 2854 3974 2860
rect 4336 2854 4394 2860
rect 4756 2854 4814 2860
rect 5176 2854 5234 2860
rect 5596 2854 5654 2860
rect -2536 2820 -2372 2854
rect -2338 2820 -1952 2854
rect -1918 2820 -1532 2854
rect -1498 2820 -1112 2854
rect -1078 2820 -692 2854
rect -658 2820 -272 2854
rect -238 2820 148 2854
rect 182 2820 568 2854
rect 602 2820 988 2854
rect 1022 2820 1408 2854
rect 1442 2820 1828 2854
rect 1862 2820 2248 2854
rect 2282 2820 2668 2854
rect 2702 2820 3088 2854
rect 3122 2820 3508 2854
rect 3542 2820 3928 2854
rect 3962 2820 4348 2854
rect 4382 2820 4768 2854
rect 4802 2820 5188 2854
rect 5222 2820 5608 2854
rect 5642 2820 5912 2854
rect -2536 2811 -2526 2820
rect -2384 2814 -2326 2820
rect -1971 2811 -1899 2820
rect -1544 2814 -1486 2820
rect -1124 2814 -1066 2820
rect -704 2814 -646 2820
rect -291 2811 -219 2820
rect 136 2814 194 2820
rect 556 2814 614 2820
rect 976 2814 1034 2820
rect 1389 2811 1461 2820
rect 1816 2814 1874 2820
rect 2236 2814 2294 2820
rect 2656 2814 2714 2820
rect 3076 2814 3134 2820
rect 3496 2814 3554 2820
rect 3916 2814 3974 2820
rect 4336 2814 4394 2820
rect 4756 2814 4814 2820
rect 5176 2814 5234 2820
rect 5596 2814 5654 2820
rect -2432 2770 -2374 2776
rect -2229 2770 -2157 2776
rect -2012 2770 -1954 2776
rect -1802 2770 -1744 2776
rect -1592 2770 -1534 2776
rect -1382 2770 -1324 2776
rect -1172 2770 -1114 2776
rect -962 2770 -904 2776
rect -752 2770 -694 2776
rect -549 2770 -539 2776
rect -487 2770 -477 2776
rect -332 2770 -274 2776
rect -122 2770 -64 2776
rect 88 2770 146 2776
rect 298 2770 356 2776
rect 508 2770 566 2776
rect 718 2770 776 2776
rect 928 2770 986 2776
rect 1138 2770 1196 2776
rect 1348 2770 1406 2776
rect 1558 2770 1616 2776
rect 1768 2770 1826 2776
rect 1978 2770 2036 2776
rect 2188 2770 2246 2776
rect 2398 2770 2456 2776
rect 2608 2770 2666 2776
rect 2818 2770 2876 2776
rect 3028 2770 3086 2776
rect 3238 2770 3296 2776
rect 3448 2770 3506 2776
rect 3658 2770 3716 2776
rect 3868 2770 3926 2776
rect 4078 2770 4136 2776
rect 4288 2770 4346 2776
rect 4498 2770 4556 2776
rect 4708 2770 4766 2776
rect 4918 2770 4976 2776
rect 5128 2770 5186 2776
rect 5338 2770 5396 2776
rect 5548 2770 5606 2776
rect 5758 2770 5816 2776
rect -2432 2736 -2420 2770
rect -2386 2736 -2210 2770
rect -2176 2736 -2009 2770
rect -1957 2736 -1790 2770
rect -1756 2736 -1580 2770
rect -1546 2736 -1370 2770
rect -1336 2736 -1160 2770
rect -1126 2736 -950 2770
rect -916 2736 -740 2770
rect -706 2736 -539 2770
rect -487 2736 -320 2770
rect -286 2736 -110 2770
rect -76 2736 100 2770
rect 134 2736 310 2770
rect 344 2736 520 2770
rect 554 2736 730 2770
rect 764 2736 931 2770
rect 983 2736 1150 2770
rect 1184 2736 1360 2770
rect 1394 2736 1570 2770
rect 1604 2736 1780 2770
rect 1814 2736 1990 2770
rect 2024 2736 2200 2770
rect 2234 2736 2410 2770
rect 2444 2736 2620 2770
rect 2654 2736 2830 2770
rect 2864 2736 3040 2770
rect 3074 2736 3250 2770
rect 3284 2736 3460 2770
rect 3494 2736 3670 2770
rect 3704 2736 3880 2770
rect 3914 2736 4090 2770
rect 4124 2736 4300 2770
rect 4334 2736 4510 2770
rect 4544 2736 4720 2770
rect 4754 2736 4930 2770
rect 4964 2736 5140 2770
rect 5174 2736 5350 2770
rect 5384 2736 5560 2770
rect 5594 2736 5770 2770
rect 5804 2736 5912 2770
rect -2432 2730 -2374 2736
rect -2229 2724 -2157 2736
rect -2019 2718 -2009 2736
rect -1957 2718 -1947 2736
rect -1802 2730 -1744 2736
rect -1592 2730 -1534 2736
rect -1382 2730 -1324 2736
rect -1172 2730 -1114 2736
rect -962 2730 -904 2736
rect -752 2730 -694 2736
rect -549 2724 -539 2736
rect -487 2724 -477 2736
rect -332 2730 -274 2736
rect -122 2730 -64 2736
rect 88 2730 146 2736
rect 298 2730 356 2736
rect 508 2730 566 2736
rect 718 2730 776 2736
rect 921 2718 931 2736
rect 983 2718 993 2736
rect 1138 2730 1196 2736
rect 1348 2730 1406 2736
rect 1558 2730 1616 2736
rect 1768 2730 1826 2736
rect 1978 2730 2036 2736
rect 2188 2730 2246 2736
rect 2398 2730 2456 2736
rect 2608 2730 2666 2736
rect 2818 2730 2876 2736
rect 3028 2730 3086 2736
rect 3238 2730 3296 2736
rect 3448 2730 3506 2736
rect 3658 2730 3716 2736
rect 3868 2730 3926 2736
rect 4078 2730 4136 2736
rect 4288 2730 4346 2736
rect 4498 2730 4556 2736
rect 4708 2730 4766 2736
rect 4918 2730 4976 2736
rect 5128 2730 5186 2736
rect 5338 2730 5396 2736
rect 5548 2730 5606 2736
rect 5758 2730 5816 2736
rect -2336 2628 -2278 2634
rect -2126 2628 -2068 2634
rect -1916 2628 -1858 2634
rect -1706 2628 -1648 2634
rect -1496 2628 -1438 2634
rect -1293 2628 -1283 2640
rect -1231 2628 -1221 2640
rect -1076 2628 -1018 2634
rect -866 2628 -808 2634
rect -656 2628 -598 2634
rect -446 2628 -388 2634
rect -236 2628 -178 2634
rect -26 2628 32 2634
rect 184 2628 242 2634
rect 292 2628 302 2640
rect -2432 2594 -2324 2628
rect -2290 2594 -2114 2628
rect -2080 2594 -1904 2628
rect -1870 2594 -1694 2628
rect -1660 2594 -1484 2628
rect -1450 2594 -1283 2628
rect -1231 2594 -1064 2628
rect -1030 2594 -854 2628
rect -820 2594 -644 2628
rect -610 2594 -434 2628
rect -400 2594 -224 2628
rect -190 2594 -14 2628
rect 20 2594 196 2628
rect 230 2594 302 2628
rect -2336 2588 -2278 2594
rect -2126 2588 -2068 2594
rect -1916 2588 -1858 2594
rect -1706 2588 -1648 2594
rect -1496 2588 -1438 2594
rect -1293 2588 -1283 2594
rect -1231 2588 -1221 2594
rect -1076 2588 -1018 2594
rect -866 2588 -808 2594
rect -656 2588 -598 2594
rect -446 2588 -388 2594
rect -236 2588 -178 2594
rect -26 2588 32 2594
rect 184 2588 242 2594
rect 292 2588 302 2594
rect 354 2628 364 2640
rect 394 2628 452 2634
rect 604 2628 662 2634
rect 814 2628 872 2634
rect 1024 2628 1082 2634
rect 1234 2628 1292 2634
rect 1444 2628 1502 2634
rect 1647 2628 1657 2640
rect 1709 2628 1719 2640
rect 1864 2628 1922 2634
rect 2074 2628 2132 2634
rect 2284 2628 2342 2634
rect 2494 2628 2552 2634
rect 2704 2628 2762 2634
rect 2907 2628 2917 2640
rect 2969 2628 2979 2640
rect 3124 2628 3182 2634
rect 3334 2628 3392 2634
rect 3544 2628 3602 2634
rect 3754 2628 3812 2634
rect 3964 2628 4022 2634
rect 4174 2628 4232 2634
rect 4384 2628 4442 2634
rect 4594 2628 4652 2634
rect 4804 2628 4862 2634
rect 4911 2628 4921 2640
rect 354 2594 406 2628
rect 440 2594 616 2628
rect 650 2594 826 2628
rect 860 2594 1036 2628
rect 1070 2594 1246 2628
rect 1280 2594 1456 2628
rect 1490 2594 1657 2628
rect 1709 2594 1876 2628
rect 1910 2594 2086 2628
rect 2120 2594 2296 2628
rect 2330 2594 2506 2628
rect 2540 2594 2716 2628
rect 2750 2594 2917 2628
rect 2969 2594 3136 2628
rect 3170 2594 3346 2628
rect 3380 2594 3556 2628
rect 3590 2594 3766 2628
rect 3800 2594 3976 2628
rect 4010 2594 4186 2628
rect 4220 2594 4396 2628
rect 4430 2594 4606 2628
rect 4640 2594 4816 2628
rect 4850 2594 4921 2628
rect 354 2588 364 2594
rect 394 2588 452 2594
rect 604 2588 662 2594
rect 814 2588 872 2594
rect 1024 2588 1082 2594
rect 1234 2588 1292 2594
rect 1444 2588 1502 2594
rect 1647 2588 1657 2594
rect 1709 2588 1719 2594
rect 1864 2588 1922 2594
rect 2074 2588 2132 2594
rect 2284 2588 2342 2594
rect 2494 2588 2552 2594
rect 2704 2588 2762 2594
rect 2907 2588 2917 2594
rect 2969 2588 2979 2594
rect 3124 2588 3182 2594
rect 3334 2588 3392 2594
rect 3544 2588 3602 2594
rect 3754 2588 3812 2594
rect 3964 2588 4022 2594
rect 4174 2588 4232 2594
rect 4384 2588 4442 2594
rect 4594 2588 4652 2594
rect 4804 2588 4862 2594
rect 4911 2588 4921 2594
rect 4973 2628 4983 2640
rect 5014 2628 5072 2634
rect 5224 2628 5282 2634
rect 5434 2628 5492 2634
rect 5644 2628 5702 2634
rect 5854 2628 5912 2634
rect 4973 2594 5026 2628
rect 5060 2594 5236 2628
rect 5270 2594 5446 2628
rect 5480 2594 5656 2628
rect 5690 2594 5866 2628
rect 5900 2594 5912 2628
rect 4973 2588 4983 2594
rect 5014 2588 5072 2594
rect 5224 2588 5282 2594
rect 5434 2588 5492 2594
rect 5644 2588 5702 2594
rect 5854 2588 5912 2594
rect -2598 2501 -2588 2553
rect -2536 2544 -2526 2553
rect -2174 2544 -2116 2550
rect -1761 2544 -1689 2553
rect -1334 2544 -1276 2550
rect -914 2544 -856 2550
rect -494 2544 -436 2550
rect -81 2544 -9 2553
rect 346 2544 404 2550
rect 766 2544 824 2550
rect 1186 2544 1244 2550
rect 1599 2544 1671 2553
rect 2026 2544 2084 2550
rect 2446 2544 2504 2550
rect 2866 2544 2924 2550
rect 3286 2544 3344 2550
rect 3706 2544 3764 2550
rect 4126 2544 4184 2550
rect 4546 2544 4604 2550
rect 4966 2544 5024 2550
rect 5386 2544 5444 2550
rect 5806 2544 5864 2550
rect -2536 2510 -2162 2544
rect -2128 2510 -1742 2544
rect -1708 2510 -1322 2544
rect -1288 2510 -902 2544
rect -868 2510 -482 2544
rect -448 2510 -62 2544
rect -28 2510 358 2544
rect 392 2510 778 2544
rect 812 2510 1198 2544
rect 1232 2510 1618 2544
rect 1652 2510 2038 2544
rect 2072 2510 2458 2544
rect 2492 2510 2878 2544
rect 2912 2510 3298 2544
rect 3332 2510 3718 2544
rect 3752 2510 4138 2544
rect 4172 2510 4558 2544
rect 4592 2510 4978 2544
rect 5012 2510 5398 2544
rect 5432 2510 5818 2544
rect 5852 2510 5912 2544
rect -2536 2501 -2526 2510
rect -2174 2504 -2116 2510
rect -1761 2501 -1689 2510
rect -1334 2504 -1276 2510
rect -914 2504 -856 2510
rect -494 2504 -436 2510
rect -81 2501 -9 2510
rect 346 2504 404 2510
rect 766 2504 824 2510
rect 1186 2504 1244 2510
rect 1599 2501 1671 2510
rect 2026 2504 2084 2510
rect 2446 2504 2504 2510
rect 2866 2504 2924 2510
rect 3286 2504 3344 2510
rect 3706 2504 3764 2510
rect 4126 2504 4184 2510
rect 4546 2504 4604 2510
rect 4966 2504 5024 2510
rect 5386 2504 5444 2510
rect 5806 2504 5864 2510
rect -2598 2424 -2546 2501
rect -2598 2372 -2588 2424
rect -2536 2414 -2526 2424
rect -2391 2414 -2319 2423
rect -1964 2414 -1906 2420
rect -1551 2414 -1479 2423
rect -1124 2414 -1066 2420
rect -711 2414 -639 2423
rect -284 2414 -226 2420
rect 129 2414 201 2423
rect 556 2414 614 2420
rect 969 2414 1041 2423
rect 1396 2414 1454 2420
rect 1816 2414 1874 2420
rect 2236 2414 2294 2420
rect 2656 2414 2714 2420
rect 3076 2414 3134 2420
rect 3496 2414 3554 2420
rect 3916 2414 3974 2420
rect 4336 2414 4394 2420
rect 4756 2414 4814 2420
rect 5176 2414 5234 2420
rect 5596 2414 5654 2420
rect -2536 2380 -2372 2414
rect -2338 2380 -1952 2414
rect -1918 2380 -1532 2414
rect -1498 2380 -1112 2414
rect -1078 2380 -692 2414
rect -658 2380 -272 2414
rect -238 2380 148 2414
rect 182 2380 568 2414
rect 602 2380 988 2414
rect 1022 2380 1408 2414
rect 1442 2380 1828 2414
rect 1862 2380 2248 2414
rect 2282 2380 2668 2414
rect 2702 2380 3088 2414
rect 3122 2380 3508 2414
rect 3542 2380 3928 2414
rect 3962 2380 4348 2414
rect 4382 2380 4768 2414
rect 4802 2380 5188 2414
rect 5222 2380 5608 2414
rect 5642 2380 5912 2414
rect -2536 2372 -2526 2380
rect -2391 2371 -2319 2380
rect -1964 2374 -1906 2380
rect -1551 2371 -1479 2380
rect -1124 2374 -1066 2380
rect -711 2371 -639 2380
rect -284 2374 -226 2380
rect 129 2371 201 2380
rect 556 2374 614 2380
rect 969 2371 1041 2380
rect 1396 2374 1454 2380
rect 1816 2374 1874 2380
rect 2236 2374 2294 2380
rect 2656 2374 2714 2380
rect 3076 2374 3134 2380
rect 3496 2374 3554 2380
rect 3916 2374 3974 2380
rect 4336 2374 4394 2380
rect 4756 2374 4814 2380
rect 5176 2374 5234 2380
rect 5596 2374 5654 2380
rect -2432 2330 -2374 2336
rect -2229 2330 -2157 2336
rect -2012 2330 -1954 2336
rect -1802 2330 -1744 2336
rect -1592 2330 -1534 2336
rect -1382 2330 -1324 2336
rect -1172 2330 -1114 2336
rect -962 2330 -904 2336
rect -752 2330 -694 2336
rect -549 2330 -539 2336
rect -487 2330 -477 2336
rect -332 2330 -274 2336
rect -122 2330 -64 2336
rect 88 2330 146 2336
rect 298 2330 356 2336
rect 508 2330 566 2336
rect 718 2330 776 2336
rect 928 2330 986 2336
rect 1138 2330 1196 2336
rect 1348 2330 1406 2336
rect 1558 2330 1616 2336
rect 1768 2330 1826 2336
rect 1978 2330 2036 2336
rect 2188 2330 2246 2336
rect 2398 2330 2456 2336
rect 2608 2330 2666 2336
rect 2818 2330 2876 2336
rect 3028 2330 3086 2336
rect 3238 2330 3296 2336
rect 3448 2330 3506 2336
rect 3658 2330 3716 2336
rect 3868 2330 3926 2336
rect 4078 2330 4136 2336
rect 4288 2330 4346 2336
rect 4498 2330 4556 2336
rect 4708 2330 4766 2336
rect 4918 2330 4976 2336
rect 5128 2330 5186 2336
rect 5338 2330 5396 2336
rect 5548 2330 5606 2336
rect 5758 2330 5816 2336
rect -2432 2296 -2420 2330
rect -2386 2296 -2210 2330
rect -2176 2296 -2009 2330
rect -1957 2296 -1790 2330
rect -1756 2296 -1580 2330
rect -1546 2296 -1370 2330
rect -1336 2296 -1160 2330
rect -1126 2296 -950 2330
rect -916 2296 -740 2330
rect -706 2296 -539 2330
rect -487 2296 -320 2330
rect -286 2296 -110 2330
rect -76 2296 100 2330
rect 134 2296 310 2330
rect 344 2296 520 2330
rect 554 2296 730 2330
rect 764 2296 931 2330
rect 983 2296 1150 2330
rect 1184 2296 1360 2330
rect 1394 2296 1570 2330
rect 1604 2296 1780 2330
rect 1814 2296 1990 2330
rect 2024 2296 2200 2330
rect 2234 2296 2410 2330
rect 2444 2296 2620 2330
rect 2654 2296 2830 2330
rect 2864 2296 3040 2330
rect 3074 2296 3250 2330
rect 3284 2296 3460 2330
rect 3494 2296 3670 2330
rect 3704 2296 3880 2330
rect 3914 2296 4090 2330
rect 4124 2296 4300 2330
rect 4334 2296 4510 2330
rect 4544 2296 4720 2330
rect 4754 2296 4930 2330
rect 4964 2296 5140 2330
rect 5174 2296 5350 2330
rect 5384 2296 5560 2330
rect 5594 2296 5770 2330
rect 5804 2296 5912 2330
rect -2432 2290 -2374 2296
rect -2229 2284 -2157 2296
rect -2019 2278 -2009 2296
rect -1957 2278 -1947 2296
rect -1802 2290 -1744 2296
rect -1592 2290 -1534 2296
rect -1382 2290 -1324 2296
rect -1172 2290 -1114 2296
rect -962 2290 -904 2296
rect -752 2290 -694 2296
rect -549 2284 -539 2296
rect -487 2284 -477 2296
rect -332 2290 -274 2296
rect -122 2290 -64 2296
rect 88 2290 146 2296
rect 298 2290 356 2296
rect 508 2290 566 2296
rect 718 2290 776 2296
rect 921 2278 931 2296
rect 983 2278 993 2296
rect 1138 2290 1196 2296
rect 1348 2290 1406 2296
rect 1558 2290 1616 2296
rect 1768 2290 1826 2296
rect 1978 2290 2036 2296
rect 2188 2290 2246 2296
rect 2398 2290 2456 2296
rect 2608 2290 2666 2296
rect 2818 2290 2876 2296
rect 3028 2290 3086 2296
rect 3238 2290 3296 2296
rect 3448 2290 3506 2296
rect 3658 2290 3716 2296
rect 3868 2290 3926 2296
rect 4078 2290 4136 2296
rect 4288 2290 4346 2296
rect 4498 2290 4556 2296
rect 4708 2290 4766 2296
rect 4918 2290 4976 2296
rect 5128 2290 5186 2296
rect 5338 2290 5396 2296
rect 5548 2290 5606 2296
rect 5758 2290 5816 2296
rect -2336 2188 -2278 2194
rect -2126 2188 -2068 2194
rect -1916 2188 -1858 2194
rect -1706 2188 -1648 2194
rect -1496 2188 -1438 2194
rect -1293 2188 -1283 2200
rect -1231 2188 -1221 2200
rect -1076 2188 -1018 2194
rect -866 2188 -808 2194
rect -656 2188 -598 2194
rect -446 2188 -388 2194
rect -236 2188 -178 2194
rect -26 2188 32 2194
rect 184 2188 242 2194
rect 292 2188 302 2200
rect -2432 2154 -2324 2188
rect -2290 2154 -2114 2188
rect -2080 2154 -1904 2188
rect -1870 2154 -1694 2188
rect -1660 2154 -1484 2188
rect -1450 2154 -1283 2188
rect -1231 2154 -1064 2188
rect -1030 2154 -854 2188
rect -820 2154 -644 2188
rect -610 2154 -434 2188
rect -400 2154 -224 2188
rect -190 2154 -14 2188
rect 20 2154 196 2188
rect 230 2154 302 2188
rect -2336 2148 -2278 2154
rect -2126 2148 -2068 2154
rect -1916 2148 -1858 2154
rect -1706 2148 -1648 2154
rect -1496 2148 -1438 2154
rect -1293 2148 -1283 2154
rect -1231 2148 -1221 2154
rect -1076 2148 -1018 2154
rect -866 2148 -808 2154
rect -656 2148 -598 2154
rect -446 2148 -388 2154
rect -236 2148 -178 2154
rect -26 2148 32 2154
rect 184 2148 242 2154
rect 292 2148 302 2154
rect 354 2188 364 2200
rect 394 2188 452 2194
rect 604 2188 662 2194
rect 814 2188 872 2194
rect 1024 2188 1082 2194
rect 1234 2188 1292 2194
rect 1444 2188 1502 2194
rect 1647 2188 1657 2200
rect 1709 2188 1719 2200
rect 1864 2188 1922 2194
rect 2074 2188 2132 2194
rect 2284 2188 2342 2194
rect 2494 2188 2552 2194
rect 2704 2188 2762 2194
rect 2907 2188 2917 2200
rect 2969 2188 2979 2200
rect 3124 2188 3182 2194
rect 3334 2188 3392 2194
rect 3544 2188 3602 2194
rect 3754 2188 3812 2194
rect 3964 2188 4022 2194
rect 4174 2188 4232 2194
rect 4384 2188 4442 2194
rect 4594 2188 4652 2194
rect 4804 2188 4862 2194
rect 4911 2188 4921 2200
rect 354 2154 406 2188
rect 440 2154 616 2188
rect 650 2154 826 2188
rect 860 2154 1036 2188
rect 1070 2154 1246 2188
rect 1280 2154 1456 2188
rect 1490 2154 1657 2188
rect 1709 2154 1876 2188
rect 1910 2154 2086 2188
rect 2120 2154 2296 2188
rect 2330 2154 2506 2188
rect 2540 2154 2716 2188
rect 2750 2154 2917 2188
rect 2969 2154 3136 2188
rect 3170 2154 3346 2188
rect 3380 2154 3556 2188
rect 3590 2154 3766 2188
rect 3800 2154 3976 2188
rect 4010 2154 4186 2188
rect 4220 2154 4396 2188
rect 4430 2154 4606 2188
rect 4640 2154 4816 2188
rect 4850 2154 4921 2188
rect 354 2148 364 2154
rect 394 2148 452 2154
rect 604 2148 662 2154
rect 814 2148 872 2154
rect 1024 2148 1082 2154
rect 1234 2148 1292 2154
rect 1444 2148 1502 2154
rect 1647 2148 1657 2154
rect 1709 2148 1719 2154
rect 1864 2148 1922 2154
rect 2074 2148 2132 2154
rect 2284 2148 2342 2154
rect 2494 2148 2552 2154
rect 2704 2148 2762 2154
rect 2907 2148 2917 2154
rect 2969 2148 2979 2154
rect 3124 2148 3182 2154
rect 3334 2148 3392 2154
rect 3544 2148 3602 2154
rect 3754 2148 3812 2154
rect 3964 2148 4022 2154
rect 4174 2148 4232 2154
rect 4384 2148 4442 2154
rect 4594 2148 4652 2154
rect 4804 2148 4862 2154
rect 4911 2148 4921 2154
rect 4973 2188 4983 2200
rect 5014 2188 5072 2194
rect 5224 2188 5282 2194
rect 5434 2188 5492 2194
rect 5644 2188 5702 2194
rect 5854 2188 5912 2194
rect 4973 2154 5026 2188
rect 5060 2154 5236 2188
rect 5270 2154 5446 2188
rect 5480 2154 5656 2188
rect 5690 2154 5866 2188
rect 5900 2154 5912 2188
rect 4973 2148 4983 2154
rect 5014 2148 5072 2154
rect 5224 2148 5282 2154
rect 5434 2148 5492 2154
rect 5644 2148 5702 2154
rect 5854 2148 5912 2154
rect -2598 2061 -2588 2113
rect -2536 2104 -2526 2113
rect -2181 2104 -2109 2113
rect -1754 2104 -1696 2110
rect -1341 2104 -1269 2113
rect -914 2104 -856 2110
rect -501 2104 -429 2113
rect -74 2104 -16 2110
rect 339 2104 411 2113
rect 766 2104 824 2110
rect 1179 2104 1251 2113
rect 1606 2104 1664 2110
rect 2026 2104 2084 2110
rect 2446 2104 2504 2110
rect 2866 2104 2924 2110
rect 3286 2104 3344 2110
rect 3706 2104 3764 2110
rect 4126 2104 4184 2110
rect 4546 2104 4604 2110
rect 4966 2104 5024 2110
rect 5386 2104 5444 2110
rect 5806 2104 5864 2110
rect -2536 2070 -2162 2104
rect -2128 2070 -1742 2104
rect -1708 2070 -1322 2104
rect -1288 2070 -902 2104
rect -868 2070 -482 2104
rect -448 2070 -62 2104
rect -28 2070 358 2104
rect 392 2070 778 2104
rect 812 2070 1198 2104
rect 1232 2070 1618 2104
rect 1652 2070 2038 2104
rect 2072 2070 2458 2104
rect 2492 2070 2878 2104
rect 2912 2070 3298 2104
rect 3332 2070 3718 2104
rect 3752 2070 4138 2104
rect 4172 2070 4558 2104
rect 4592 2070 4978 2104
rect 5012 2070 5398 2104
rect 5432 2070 5818 2104
rect 5852 2070 5912 2104
rect -2536 2061 -2526 2070
rect -2181 2061 -2109 2070
rect -1754 2064 -1696 2070
rect -1341 2061 -1269 2070
rect -914 2064 -856 2070
rect -501 2061 -429 2070
rect -74 2064 -16 2070
rect 339 2061 411 2070
rect 766 2064 824 2070
rect 1179 2061 1251 2070
rect 1606 2064 1664 2070
rect 2026 2064 2084 2070
rect 2446 2064 2504 2070
rect 2866 2064 2924 2070
rect 3286 2064 3344 2070
rect 3706 2064 3764 2070
rect 4126 2064 4184 2070
rect 4546 2064 4604 2070
rect 4966 2064 5024 2070
rect 5386 2064 5444 2070
rect 5806 2064 5864 2070
rect -2384 1974 -2326 1980
rect -1971 1974 -1899 1983
rect -1544 1974 -1486 1980
rect -1124 1974 -1066 1980
rect -704 1974 -646 1980
rect -291 1974 -219 1983
rect 136 1974 194 1980
rect 556 1974 614 1980
rect 976 1974 1034 1980
rect 1389 1974 1461 1983
rect 1816 1974 1874 1980
rect 2236 1974 2294 1980
rect 2656 1974 2714 1980
rect 3076 1974 3134 1980
rect 3496 1974 3554 1980
rect 3916 1974 3974 1980
rect 4336 1974 4394 1980
rect 4756 1974 4814 1980
rect 5176 1974 5234 1980
rect 5596 1974 5654 1980
rect 6010 1974 6020 1985
rect -2432 1940 -2372 1974
rect -2338 1940 -1952 1974
rect -1918 1940 -1532 1974
rect -1498 1940 -1112 1974
rect -1078 1940 -692 1974
rect -658 1940 -272 1974
rect -238 1940 148 1974
rect 182 1940 568 1974
rect 602 1940 988 1974
rect 1022 1940 1408 1974
rect 1442 1940 1828 1974
rect 1862 1940 2248 1974
rect 2282 1940 2668 1974
rect 2702 1940 3088 1974
rect 3122 1940 3508 1974
rect 3542 1940 3928 1974
rect 3962 1940 4348 1974
rect 4382 1940 4768 1974
rect 4802 1940 5188 1974
rect 5222 1940 5608 1974
rect 5642 1940 6020 1974
rect -2384 1934 -2326 1940
rect -1971 1931 -1899 1940
rect -1544 1934 -1486 1940
rect -1124 1934 -1066 1940
rect -704 1934 -646 1940
rect -291 1931 -219 1940
rect 136 1934 194 1940
rect 556 1934 614 1940
rect 976 1934 1034 1940
rect 1389 1931 1461 1940
rect 1816 1934 1874 1940
rect 2236 1934 2294 1940
rect 2656 1934 2714 1940
rect 3076 1934 3134 1940
rect 3496 1934 3554 1940
rect 3916 1934 3974 1940
rect 4336 1934 4394 1940
rect 4756 1934 4814 1940
rect 5176 1934 5234 1940
rect 5596 1934 5654 1940
rect 6010 1933 6020 1940
rect 6072 1974 6082 1985
rect 6072 1940 6088 1974
rect 6072 1933 6082 1940
rect -2432 1890 -2374 1896
rect -2222 1890 -2164 1896
rect -2012 1890 -1954 1896
rect -1802 1890 -1744 1896
rect -1592 1890 -1534 1896
rect -1382 1890 -1324 1896
rect -1172 1890 -1114 1896
rect -962 1890 -904 1896
rect -752 1890 -694 1896
rect -542 1890 -484 1896
rect -332 1890 -274 1896
rect -122 1890 -64 1896
rect 88 1890 146 1896
rect 298 1890 356 1896
rect 508 1890 566 1896
rect 718 1890 776 1896
rect 928 1890 986 1896
rect 1138 1890 1196 1896
rect 1348 1890 1406 1896
rect 1558 1890 1616 1896
rect 1768 1890 1826 1896
rect 1978 1890 2036 1896
rect 2188 1890 2246 1896
rect 2398 1890 2456 1896
rect 2608 1890 2666 1896
rect 2818 1890 2876 1896
rect 3028 1890 3086 1896
rect 3238 1890 3296 1896
rect 3448 1890 3506 1896
rect 3658 1890 3716 1896
rect 3868 1890 3926 1896
rect 4078 1890 4136 1896
rect 4288 1890 4346 1896
rect 4498 1890 4556 1896
rect 4708 1890 4766 1896
rect 4918 1890 4976 1896
rect 5128 1890 5186 1896
rect 5338 1890 5396 1896
rect 5548 1890 5606 1896
rect 5758 1890 5816 1896
rect -2432 1856 -2420 1890
rect -2386 1856 -2210 1890
rect -2176 1856 -2000 1890
rect -1966 1856 -1790 1890
rect -1756 1856 -1580 1890
rect -1546 1856 -1370 1890
rect -1336 1856 -1160 1890
rect -1126 1856 -950 1890
rect -916 1856 -740 1890
rect -706 1856 -530 1890
rect -496 1856 -320 1890
rect -286 1856 -110 1890
rect -76 1856 100 1890
rect 134 1856 310 1890
rect 344 1856 520 1890
rect 554 1856 730 1890
rect 764 1856 940 1890
rect 974 1856 1150 1890
rect 1184 1856 1360 1890
rect 1394 1856 1570 1890
rect 1604 1856 1780 1890
rect 1814 1856 1990 1890
rect 2024 1856 2200 1890
rect 2234 1856 2401 1890
rect 2453 1856 2620 1890
rect 2654 1856 2830 1890
rect 2864 1856 3040 1890
rect 3074 1856 3250 1890
rect 3284 1856 3460 1890
rect 3494 1856 3670 1890
rect 3704 1856 3871 1890
rect 3923 1856 4090 1890
rect 4124 1856 4300 1890
rect 4334 1856 4510 1890
rect 4544 1856 4720 1890
rect 4754 1856 4930 1890
rect 4964 1856 5140 1890
rect 5174 1856 5340 1890
rect 5392 1856 5560 1890
rect 5594 1856 5770 1890
rect 5804 1856 5912 1890
rect -2432 1850 -2374 1856
rect -2222 1850 -2164 1856
rect -2012 1850 -1954 1856
rect -1802 1850 -1744 1856
rect -1592 1850 -1534 1856
rect -1382 1850 -1324 1856
rect -1172 1850 -1114 1856
rect -962 1850 -904 1856
rect -752 1850 -694 1856
rect -542 1850 -484 1856
rect -332 1850 -274 1856
rect -122 1850 -64 1856
rect 88 1850 146 1856
rect 298 1850 356 1856
rect 508 1850 566 1856
rect 718 1850 776 1856
rect 928 1850 986 1856
rect 1138 1850 1196 1856
rect 1348 1850 1406 1856
rect 1558 1850 1616 1856
rect 1768 1850 1826 1856
rect 1978 1850 2036 1856
rect 2188 1850 2246 1856
rect 2391 1838 2401 1856
rect 2453 1838 2463 1856
rect 2608 1850 2666 1856
rect 2818 1850 2876 1856
rect 3028 1850 3086 1856
rect 3238 1850 3296 1856
rect 3448 1850 3506 1856
rect 3658 1850 3716 1856
rect 3861 1838 3871 1856
rect 3923 1838 3933 1856
rect 4078 1850 4136 1856
rect 4288 1850 4346 1856
rect 4498 1850 4556 1856
rect 4708 1850 4766 1856
rect 4918 1850 4976 1856
rect 5128 1850 5186 1856
rect 5330 1838 5340 1856
rect 5392 1838 5402 1856
rect 5548 1850 5606 1856
rect 5758 1850 5816 1856
rect -2336 1748 -2278 1754
rect -2126 1748 -2068 1754
rect -1916 1748 -1858 1754
rect -1706 1748 -1648 1754
rect -1496 1748 -1438 1754
rect -1293 1748 -1283 1760
rect -1231 1748 -1221 1760
rect -1076 1748 -1018 1754
rect -866 1748 -808 1754
rect -656 1748 -598 1754
rect -446 1748 -388 1754
rect -236 1748 -178 1754
rect -26 1748 32 1754
rect 184 1748 242 1754
rect 292 1748 302 1760
rect -2432 1714 -2324 1748
rect -2290 1714 -2114 1748
rect -2080 1714 -1904 1748
rect -1870 1714 -1694 1748
rect -1660 1714 -1484 1748
rect -1450 1714 -1283 1748
rect -1231 1714 -1064 1748
rect -1030 1714 -854 1748
rect -820 1714 -644 1748
rect -610 1714 -434 1748
rect -400 1714 -224 1748
rect -190 1714 -14 1748
rect 20 1714 196 1748
rect 230 1714 302 1748
rect -2336 1708 -2278 1714
rect -2126 1708 -2068 1714
rect -1916 1708 -1858 1714
rect -1706 1708 -1648 1714
rect -1496 1708 -1438 1714
rect -1293 1708 -1283 1714
rect -1231 1708 -1221 1714
rect -1076 1708 -1018 1714
rect -866 1708 -808 1714
rect -656 1708 -598 1714
rect -446 1708 -388 1714
rect -236 1708 -178 1714
rect -26 1708 32 1714
rect 184 1708 242 1714
rect 292 1708 302 1714
rect 354 1748 364 1760
rect 394 1748 452 1754
rect 604 1748 662 1754
rect 814 1748 872 1754
rect 1024 1748 1082 1754
rect 1234 1748 1292 1754
rect 1444 1748 1502 1754
rect 1647 1748 1657 1760
rect 1709 1748 1719 1760
rect 1864 1748 1922 1754
rect 2074 1748 2132 1754
rect 2284 1748 2342 1754
rect 2494 1748 2552 1754
rect 2704 1748 2762 1754
rect 2907 1748 2917 1760
rect 2969 1748 2979 1760
rect 3124 1748 3182 1754
rect 3334 1748 3392 1754
rect 3544 1748 3602 1754
rect 3754 1748 3812 1754
rect 3964 1748 4022 1754
rect 4174 1748 4232 1754
rect 4384 1748 4442 1754
rect 4594 1748 4652 1754
rect 4804 1748 4862 1754
rect 4911 1748 4921 1760
rect 354 1714 406 1748
rect 440 1714 616 1748
rect 650 1714 826 1748
rect 860 1714 1036 1748
rect 1070 1714 1246 1748
rect 1280 1714 1456 1748
rect 1490 1714 1657 1748
rect 1709 1714 1876 1748
rect 1910 1714 2086 1748
rect 2120 1714 2296 1748
rect 2330 1714 2506 1748
rect 2540 1714 2716 1748
rect 2750 1714 2917 1748
rect 2969 1714 3136 1748
rect 3170 1714 3346 1748
rect 3380 1714 3556 1748
rect 3590 1714 3766 1748
rect 3800 1714 3976 1748
rect 4010 1714 4186 1748
rect 4220 1714 4396 1748
rect 4430 1714 4606 1748
rect 4640 1714 4816 1748
rect 4850 1714 4921 1748
rect 354 1708 364 1714
rect 394 1708 452 1714
rect 604 1708 662 1714
rect 814 1708 872 1714
rect 1024 1708 1082 1714
rect 1234 1708 1292 1714
rect 1444 1708 1502 1714
rect 1647 1708 1657 1714
rect 1709 1708 1719 1714
rect 1864 1708 1922 1714
rect 2074 1708 2132 1714
rect 2284 1708 2342 1714
rect 2494 1708 2552 1714
rect 2704 1708 2762 1714
rect 2907 1708 2917 1714
rect 2969 1708 2979 1714
rect 3124 1708 3182 1714
rect 3334 1708 3392 1714
rect 3544 1708 3602 1714
rect 3754 1708 3812 1714
rect 3964 1708 4022 1714
rect 4174 1708 4232 1714
rect 4384 1708 4442 1714
rect 4594 1708 4652 1714
rect 4804 1708 4862 1714
rect 4911 1708 4921 1714
rect 4973 1748 4983 1760
rect 5014 1748 5072 1754
rect 5224 1748 5282 1754
rect 5434 1748 5492 1754
rect 5644 1748 5702 1754
rect 5854 1748 5912 1754
rect 4973 1714 5026 1748
rect 5060 1714 5236 1748
rect 5270 1714 5446 1748
rect 5480 1714 5656 1748
rect 5690 1714 5866 1748
rect 5900 1714 5912 1748
rect 4973 1708 4983 1714
rect 5014 1708 5072 1714
rect 5224 1708 5282 1714
rect 5434 1708 5492 1714
rect 5644 1708 5702 1714
rect 5854 1708 5912 1714
rect -2174 1664 -2116 1670
rect -1761 1664 -1689 1673
rect -1334 1664 -1276 1670
rect -914 1664 -856 1670
rect -494 1664 -436 1670
rect -81 1664 -9 1673
rect 346 1664 404 1670
rect 766 1664 824 1670
rect 1186 1664 1244 1670
rect 1599 1664 1671 1673
rect 2026 1664 2084 1670
rect 2446 1664 2504 1670
rect 2866 1664 2924 1670
rect 3286 1664 3344 1670
rect 3706 1664 3764 1670
rect 4126 1664 4184 1670
rect 4546 1664 4604 1670
rect 4966 1664 5024 1670
rect 5386 1664 5444 1670
rect 5806 1664 5864 1670
rect 6010 1664 6020 1671
rect -2432 1630 -2162 1664
rect -2128 1630 -1742 1664
rect -1708 1630 -1322 1664
rect -1288 1630 -902 1664
rect -868 1630 -482 1664
rect -448 1630 -62 1664
rect -28 1630 358 1664
rect 392 1630 778 1664
rect 812 1630 1198 1664
rect 1232 1630 1618 1664
rect 1652 1630 2038 1664
rect 2072 1630 2458 1664
rect 2492 1630 2878 1664
rect 2912 1630 3298 1664
rect 3332 1630 3718 1664
rect 3752 1630 4138 1664
rect 4172 1630 4558 1664
rect 4592 1630 4978 1664
rect 5012 1630 5398 1664
rect 5432 1630 5818 1664
rect 5852 1630 6020 1664
rect -2174 1624 -2116 1630
rect -1761 1621 -1689 1630
rect -1334 1624 -1276 1630
rect -914 1624 -856 1630
rect -494 1624 -436 1630
rect -81 1621 -9 1630
rect 346 1624 404 1630
rect 766 1624 824 1630
rect 1186 1624 1244 1630
rect 1599 1621 1671 1630
rect 2026 1624 2084 1630
rect 2446 1624 2504 1630
rect 2866 1624 2924 1630
rect 3286 1624 3344 1630
rect 3706 1624 3764 1630
rect 4126 1624 4184 1630
rect 4546 1624 4604 1630
rect 4966 1624 5024 1630
rect 5386 1624 5444 1630
rect 5806 1624 5864 1630
rect 6010 1619 6020 1630
rect 6072 1664 6082 1671
rect 6072 1630 6083 1664
rect 6072 1619 6082 1630
rect -2391 1534 -2319 1543
rect -1964 1534 -1906 1540
rect -1551 1534 -1479 1543
rect -1124 1534 -1066 1540
rect -711 1534 -639 1543
rect -284 1534 -226 1540
rect 129 1534 201 1543
rect 556 1534 614 1540
rect 969 1534 1041 1543
rect 1396 1534 1454 1540
rect 1816 1534 1874 1540
rect 2236 1534 2294 1540
rect 2656 1534 2714 1540
rect 3076 1534 3134 1540
rect 3496 1534 3554 1540
rect 3916 1534 3974 1540
rect 4336 1534 4394 1540
rect 4756 1534 4814 1540
rect 5176 1534 5234 1540
rect 5596 1534 5654 1540
rect 6010 1534 6020 1544
rect -2432 1500 -2372 1534
rect -2338 1500 -1952 1534
rect -1918 1500 -1532 1534
rect -1498 1500 -1112 1534
rect -1078 1500 -692 1534
rect -658 1500 -272 1534
rect -238 1500 148 1534
rect 182 1500 568 1534
rect 602 1500 988 1534
rect 1022 1500 1408 1534
rect 1442 1500 1828 1534
rect 1862 1500 2248 1534
rect 2282 1500 2668 1534
rect 2702 1500 3088 1534
rect 3122 1500 3508 1534
rect 3542 1500 3928 1534
rect 3962 1500 4348 1534
rect 4382 1500 4768 1534
rect 4802 1500 5188 1534
rect 5222 1500 5608 1534
rect 5642 1500 6020 1534
rect -2391 1491 -2319 1500
rect -1964 1494 -1906 1500
rect -1551 1491 -1479 1500
rect -1124 1494 -1066 1500
rect -711 1491 -639 1500
rect -284 1494 -226 1500
rect 129 1491 201 1500
rect 556 1494 614 1500
rect 969 1491 1041 1500
rect 1396 1494 1454 1500
rect 1816 1494 1874 1500
rect 2236 1494 2294 1500
rect 2656 1494 2714 1500
rect 3076 1494 3134 1500
rect 3496 1494 3554 1500
rect 3916 1494 3974 1500
rect 4336 1494 4394 1500
rect 4756 1494 4814 1500
rect 5176 1494 5234 1500
rect 5596 1494 5654 1500
rect 6010 1492 6020 1500
rect 6072 1492 6082 1544
rect -2432 1450 -2374 1456
rect -2222 1450 -2164 1456
rect -2012 1450 -1954 1456
rect -1802 1450 -1744 1456
rect -1592 1450 -1534 1456
rect -1382 1450 -1324 1456
rect -1172 1450 -1114 1456
rect -962 1450 -904 1456
rect -752 1450 -694 1456
rect -542 1450 -484 1456
rect -332 1450 -274 1456
rect -122 1450 -64 1456
rect 88 1450 146 1456
rect 298 1450 356 1456
rect 508 1450 566 1456
rect 718 1450 776 1456
rect 928 1450 986 1456
rect 1138 1450 1196 1456
rect 1348 1450 1406 1456
rect 1558 1450 1616 1456
rect 1768 1450 1826 1456
rect 1978 1450 2036 1456
rect 2188 1450 2246 1456
rect 2398 1450 2456 1456
rect 2608 1450 2666 1456
rect 2818 1450 2876 1456
rect 3028 1450 3086 1456
rect 3238 1450 3296 1456
rect 3448 1450 3506 1456
rect 3658 1450 3716 1456
rect 3868 1450 3926 1456
rect 4078 1450 4136 1456
rect 4288 1450 4346 1456
rect 4498 1450 4556 1456
rect 4708 1450 4766 1456
rect 4918 1450 4976 1456
rect 5128 1450 5186 1456
rect 5338 1450 5396 1456
rect 5548 1450 5606 1456
rect 5758 1450 5816 1456
rect -2432 1416 -2420 1450
rect -2386 1416 -2210 1450
rect -2176 1416 -2000 1450
rect -1966 1416 -1790 1450
rect -1756 1416 -1580 1450
rect -1546 1416 -1370 1450
rect -1336 1416 -1160 1450
rect -1126 1416 -950 1450
rect -916 1416 -740 1450
rect -706 1416 -530 1450
rect -496 1416 -320 1450
rect -286 1416 -110 1450
rect -76 1416 100 1450
rect 134 1416 310 1450
rect 344 1416 520 1450
rect 554 1416 730 1450
rect 764 1416 940 1450
rect 974 1416 1150 1450
rect 1184 1416 1360 1450
rect 1394 1416 1570 1450
rect 1604 1416 1780 1450
rect 1814 1416 1990 1450
rect 2024 1416 2200 1450
rect 2234 1416 2401 1450
rect 2453 1416 2620 1450
rect 2654 1416 2830 1450
rect 2864 1416 3040 1450
rect 3074 1416 3250 1450
rect 3284 1416 3460 1450
rect 3494 1416 3670 1450
rect 3704 1416 3871 1450
rect 3923 1416 4090 1450
rect 4124 1416 4300 1450
rect 4334 1416 4510 1450
rect 4544 1416 4720 1450
rect 4754 1416 4930 1450
rect 4964 1416 5140 1450
rect 5174 1416 5340 1450
rect 5392 1416 5560 1450
rect 5594 1416 5770 1450
rect 5804 1416 5912 1450
rect -2432 1410 -2374 1416
rect -2222 1410 -2164 1416
rect -2012 1410 -1954 1416
rect -1802 1410 -1744 1416
rect -1592 1410 -1534 1416
rect -1382 1410 -1324 1416
rect -1172 1410 -1114 1416
rect -962 1410 -904 1416
rect -752 1410 -694 1416
rect -542 1410 -484 1416
rect -332 1410 -274 1416
rect -122 1410 -64 1416
rect 88 1410 146 1416
rect 298 1410 356 1416
rect 508 1410 566 1416
rect 718 1410 776 1416
rect 928 1410 986 1416
rect 1138 1410 1196 1416
rect 1348 1410 1406 1416
rect 1558 1410 1616 1416
rect 1768 1410 1826 1416
rect 1978 1410 2036 1416
rect 2188 1410 2246 1416
rect 2391 1398 2401 1416
rect 2453 1398 2463 1416
rect 2608 1410 2666 1416
rect 2818 1410 2876 1416
rect 3028 1410 3086 1416
rect 3238 1410 3296 1416
rect 3448 1410 3506 1416
rect 3658 1410 3716 1416
rect 3861 1398 3871 1416
rect 3923 1398 3933 1416
rect 4078 1410 4136 1416
rect 4288 1410 4346 1416
rect 4498 1410 4556 1416
rect 4708 1410 4766 1416
rect 4918 1410 4976 1416
rect 5128 1410 5186 1416
rect 5330 1398 5340 1416
rect 5392 1398 5402 1416
rect 5548 1410 5606 1416
rect 5758 1410 5816 1416
rect -2336 1308 -2278 1314
rect -2126 1308 -2068 1314
rect -1916 1308 -1858 1314
rect -1706 1308 -1648 1314
rect -1496 1308 -1438 1314
rect -1293 1308 -1283 1320
rect -1231 1308 -1221 1320
rect -1076 1308 -1018 1314
rect -866 1308 -808 1314
rect -656 1308 -598 1314
rect -446 1308 -388 1314
rect -236 1308 -178 1314
rect -26 1308 32 1314
rect 184 1308 242 1314
rect 292 1308 302 1320
rect -2432 1274 -2324 1308
rect -2290 1274 -2114 1308
rect -2080 1274 -1904 1308
rect -1870 1274 -1694 1308
rect -1660 1274 -1484 1308
rect -1450 1274 -1283 1308
rect -1231 1274 -1064 1308
rect -1030 1274 -854 1308
rect -820 1274 -644 1308
rect -610 1274 -434 1308
rect -400 1274 -224 1308
rect -190 1274 -14 1308
rect 20 1274 196 1308
rect 230 1274 302 1308
rect -2336 1268 -2278 1274
rect -2126 1268 -2068 1274
rect -1916 1268 -1858 1274
rect -1706 1268 -1648 1274
rect -1496 1268 -1438 1274
rect -1293 1268 -1283 1274
rect -1231 1268 -1221 1274
rect -1076 1268 -1018 1274
rect -866 1268 -808 1274
rect -656 1268 -598 1274
rect -446 1268 -388 1274
rect -236 1268 -178 1274
rect -26 1268 32 1274
rect 184 1268 242 1274
rect 292 1268 302 1274
rect 354 1308 364 1320
rect 394 1308 452 1314
rect 604 1308 662 1314
rect 814 1308 872 1314
rect 1024 1308 1082 1314
rect 1234 1308 1292 1314
rect 1444 1308 1502 1314
rect 1647 1308 1657 1320
rect 1709 1308 1719 1320
rect 1864 1308 1922 1314
rect 2074 1308 2132 1314
rect 2284 1308 2342 1314
rect 2494 1308 2552 1314
rect 2704 1308 2762 1314
rect 2907 1308 2917 1320
rect 2969 1308 2979 1320
rect 3124 1308 3182 1314
rect 3334 1308 3392 1314
rect 3544 1308 3602 1314
rect 3754 1308 3812 1314
rect 3964 1308 4022 1314
rect 4174 1308 4232 1314
rect 4384 1308 4442 1314
rect 4594 1308 4652 1314
rect 4804 1308 4862 1314
rect 4911 1308 4921 1320
rect 354 1274 406 1308
rect 440 1274 616 1308
rect 650 1274 826 1308
rect 860 1274 1036 1308
rect 1070 1274 1246 1308
rect 1280 1274 1456 1308
rect 1490 1274 1657 1308
rect 1709 1274 1876 1308
rect 1910 1274 2086 1308
rect 2120 1274 2296 1308
rect 2330 1274 2506 1308
rect 2540 1274 2716 1308
rect 2750 1274 2917 1308
rect 2969 1274 3136 1308
rect 3170 1274 3346 1308
rect 3380 1274 3556 1308
rect 3590 1274 3766 1308
rect 3800 1274 3976 1308
rect 4010 1274 4186 1308
rect 4220 1274 4396 1308
rect 4430 1274 4606 1308
rect 4640 1274 4816 1308
rect 4850 1274 4921 1308
rect 354 1268 364 1274
rect 394 1268 452 1274
rect 604 1268 662 1274
rect 814 1268 872 1274
rect 1024 1268 1082 1274
rect 1234 1268 1292 1274
rect 1444 1268 1502 1274
rect 1647 1268 1657 1274
rect 1709 1268 1719 1274
rect 1864 1268 1922 1274
rect 2074 1268 2132 1274
rect 2284 1268 2342 1274
rect 2494 1268 2552 1274
rect 2704 1268 2762 1274
rect 2907 1268 2917 1274
rect 2969 1268 2979 1274
rect 3124 1268 3182 1274
rect 3334 1268 3392 1274
rect 3544 1268 3602 1274
rect 3754 1268 3812 1274
rect 3964 1268 4022 1274
rect 4174 1268 4232 1274
rect 4384 1268 4442 1274
rect 4594 1268 4652 1274
rect 4804 1268 4862 1274
rect 4911 1268 4921 1274
rect 4973 1308 4983 1320
rect 5014 1308 5072 1314
rect 5224 1308 5282 1314
rect 5434 1308 5492 1314
rect 5644 1308 5702 1314
rect 5854 1308 5912 1314
rect 4973 1274 5026 1308
rect 5060 1274 5236 1308
rect 5270 1274 5446 1308
rect 5480 1274 5656 1308
rect 5690 1274 5866 1308
rect 5900 1274 5912 1308
rect 4973 1268 4983 1274
rect 5014 1268 5072 1274
rect 5224 1268 5282 1274
rect 5434 1268 5492 1274
rect 5644 1268 5702 1274
rect 5854 1268 5912 1274
rect -2181 1224 -2109 1233
rect -1754 1224 -1696 1230
rect -1341 1224 -1269 1233
rect -914 1224 -856 1230
rect -501 1224 -429 1233
rect -74 1224 -16 1230
rect 339 1224 411 1233
rect 766 1224 824 1230
rect 1179 1224 1251 1233
rect 1606 1224 1664 1230
rect 2026 1224 2084 1230
rect 2446 1224 2504 1230
rect 2866 1224 2924 1230
rect 3286 1224 3344 1230
rect 3706 1224 3764 1230
rect 4126 1224 4184 1230
rect 4546 1224 4604 1230
rect 4966 1224 5024 1230
rect 5386 1224 5444 1230
rect 5806 1224 5864 1230
rect 6010 1224 6020 1233
rect -2432 1190 -2162 1224
rect -2128 1190 -1742 1224
rect -1708 1190 -1322 1224
rect -1288 1190 -902 1224
rect -868 1190 -482 1224
rect -448 1190 -62 1224
rect -28 1190 358 1224
rect 392 1190 778 1224
rect 812 1190 1198 1224
rect 1232 1190 1618 1224
rect 1652 1190 2038 1224
rect 2072 1190 2458 1224
rect 2492 1190 2878 1224
rect 2912 1190 3298 1224
rect 3332 1190 3718 1224
rect 3752 1190 4138 1224
rect 4172 1190 4558 1224
rect 4592 1190 4978 1224
rect 5012 1190 5398 1224
rect 5432 1190 5818 1224
rect 5852 1190 6020 1224
rect -2181 1181 -2109 1190
rect -1754 1184 -1696 1190
rect -1341 1181 -1269 1190
rect -914 1184 -856 1190
rect -501 1181 -429 1190
rect -74 1184 -16 1190
rect 339 1181 411 1190
rect 766 1184 824 1190
rect 1179 1181 1251 1190
rect 1606 1184 1664 1190
rect 2026 1184 2084 1190
rect 2446 1184 2504 1190
rect 2866 1184 2924 1190
rect 3286 1184 3344 1190
rect 3706 1184 3764 1190
rect 4126 1184 4184 1190
rect 4546 1184 4604 1190
rect 4966 1184 5024 1190
rect 5386 1184 5444 1190
rect 5806 1184 5864 1190
rect 6010 1181 6020 1190
rect 6072 1181 6082 1233
rect -2598 1051 -2588 1103
rect -2536 1094 -2526 1103
rect -2384 1094 -2326 1100
rect -1971 1094 -1899 1103
rect -1544 1094 -1486 1100
rect -1124 1094 -1066 1100
rect -704 1094 -646 1100
rect -291 1094 -219 1103
rect 136 1094 194 1100
rect 556 1094 614 1100
rect 976 1094 1034 1100
rect 1389 1094 1461 1103
rect 1816 1094 1874 1100
rect 2236 1094 2294 1100
rect 2656 1094 2714 1100
rect 3076 1094 3134 1100
rect 3496 1094 3554 1100
rect 3916 1094 3974 1100
rect 4336 1094 4394 1100
rect 4756 1094 4814 1100
rect 5176 1094 5234 1100
rect 5596 1094 5654 1100
rect -2536 1060 -2372 1094
rect -2338 1060 -1952 1094
rect -1918 1060 -1532 1094
rect -1498 1060 -1112 1094
rect -1078 1060 -692 1094
rect -658 1060 -272 1094
rect -238 1060 148 1094
rect 182 1060 568 1094
rect 602 1060 988 1094
rect 1022 1060 1408 1094
rect 1442 1060 1828 1094
rect 1862 1060 2248 1094
rect 2282 1060 2668 1094
rect 2702 1060 3088 1094
rect 3122 1060 3508 1094
rect 3542 1060 3928 1094
rect 3962 1060 4348 1094
rect 4382 1060 4768 1094
rect 4802 1060 5188 1094
rect 5222 1060 5608 1094
rect 5642 1060 5912 1094
rect -2536 1051 -2526 1060
rect -2384 1054 -2326 1060
rect -1971 1051 -1899 1060
rect -1544 1054 -1486 1060
rect -1124 1054 -1066 1060
rect -704 1054 -646 1060
rect -291 1051 -219 1060
rect 136 1054 194 1060
rect 556 1054 614 1060
rect 976 1054 1034 1060
rect 1389 1051 1461 1060
rect 1816 1054 1874 1060
rect 2236 1054 2294 1060
rect 2656 1054 2714 1060
rect 3076 1054 3134 1060
rect 3496 1054 3554 1060
rect 3916 1054 3974 1060
rect 4336 1054 4394 1060
rect 4756 1054 4814 1060
rect 5176 1054 5234 1060
rect 5596 1054 5654 1060
rect -2432 1010 -2374 1016
rect -2229 1010 -2157 1016
rect -2012 1010 -1954 1016
rect -1802 1010 -1744 1016
rect -1592 1010 -1534 1016
rect -1382 1010 -1324 1016
rect -1172 1010 -1114 1016
rect -962 1010 -904 1016
rect -752 1010 -694 1016
rect -549 1010 -539 1016
rect -487 1010 -477 1016
rect -332 1010 -274 1016
rect -122 1010 -64 1016
rect 88 1010 146 1016
rect 298 1010 356 1016
rect 508 1010 566 1016
rect 718 1010 776 1016
rect 928 1010 986 1016
rect 1138 1010 1196 1016
rect 1348 1010 1406 1016
rect 1558 1010 1616 1016
rect 1768 1010 1826 1016
rect 1978 1010 2036 1016
rect 2188 1010 2246 1016
rect 2398 1010 2456 1016
rect 2608 1010 2666 1016
rect 2818 1010 2876 1016
rect 3028 1010 3086 1016
rect 3238 1010 3296 1016
rect 3448 1010 3506 1016
rect 3658 1010 3716 1016
rect 3868 1010 3926 1016
rect 4078 1010 4136 1016
rect 4288 1010 4346 1016
rect 4498 1010 4556 1016
rect 4708 1010 4766 1016
rect 4918 1010 4976 1016
rect 5128 1010 5186 1016
rect 5338 1010 5396 1016
rect 5548 1010 5606 1016
rect 5758 1010 5816 1016
rect -2432 976 -2420 1010
rect -2386 976 -2210 1010
rect -2176 976 -2009 1010
rect -1957 976 -1790 1010
rect -1756 976 -1580 1010
rect -1546 976 -1370 1010
rect -1336 976 -1160 1010
rect -1126 976 -950 1010
rect -916 976 -740 1010
rect -706 976 -539 1010
rect -487 976 -320 1010
rect -286 976 -110 1010
rect -76 976 100 1010
rect 134 976 310 1010
rect 344 976 520 1010
rect 554 976 730 1010
rect 764 976 931 1010
rect 983 976 1150 1010
rect 1184 976 1360 1010
rect 1394 976 1570 1010
rect 1604 976 1780 1010
rect 1814 976 1990 1010
rect 2024 976 2200 1010
rect 2234 976 2410 1010
rect 2444 976 2620 1010
rect 2654 976 2830 1010
rect 2864 976 3040 1010
rect 3074 976 3250 1010
rect 3284 976 3460 1010
rect 3494 976 3670 1010
rect 3704 976 3880 1010
rect 3914 976 4090 1010
rect 4124 976 4300 1010
rect 4334 976 4510 1010
rect 4544 976 4720 1010
rect 4754 976 4930 1010
rect 4964 976 5140 1010
rect 5174 976 5350 1010
rect 5384 976 5560 1010
rect 5594 976 5770 1010
rect 5804 976 5912 1010
rect -2432 970 -2374 976
rect -2229 964 -2157 976
rect -2019 958 -2009 976
rect -1957 958 -1947 976
rect -1802 970 -1744 976
rect -1592 970 -1534 976
rect -1382 970 -1324 976
rect -1172 970 -1114 976
rect -962 970 -904 976
rect -752 970 -694 976
rect -549 964 -539 976
rect -487 964 -477 976
rect -332 970 -274 976
rect -122 970 -64 976
rect 88 970 146 976
rect 298 970 356 976
rect 508 970 566 976
rect 718 970 776 976
rect 921 958 931 976
rect 983 958 993 976
rect 1138 970 1196 976
rect 1348 970 1406 976
rect 1558 970 1616 976
rect 1768 970 1826 976
rect 1978 970 2036 976
rect 2188 970 2246 976
rect 2398 970 2456 976
rect 2608 970 2666 976
rect 2818 970 2876 976
rect 3028 970 3086 976
rect 3238 970 3296 976
rect 3448 970 3506 976
rect 3658 970 3716 976
rect 3868 970 3926 976
rect 4078 970 4136 976
rect 4288 970 4346 976
rect 4498 970 4556 976
rect 4708 970 4766 976
rect 4918 970 4976 976
rect 5128 970 5186 976
rect 5338 970 5396 976
rect 5548 970 5606 976
rect 5758 970 5816 976
rect -2336 868 -2278 874
rect -2126 868 -2068 874
rect -1916 868 -1858 874
rect -1706 868 -1648 874
rect -1496 868 -1438 874
rect -1293 868 -1283 880
rect -1231 868 -1221 880
rect -1076 868 -1018 874
rect -866 868 -808 874
rect -656 868 -598 874
rect -446 868 -388 874
rect -236 868 -178 874
rect -26 868 32 874
rect 184 868 242 874
rect 292 868 302 880
rect -2432 834 -2324 868
rect -2290 834 -2114 868
rect -2080 834 -1904 868
rect -1870 834 -1694 868
rect -1660 834 -1484 868
rect -1450 834 -1283 868
rect -1231 834 -1064 868
rect -1030 834 -854 868
rect -820 834 -644 868
rect -610 834 -434 868
rect -400 834 -224 868
rect -190 834 -14 868
rect 20 834 196 868
rect 230 834 302 868
rect -2336 828 -2278 834
rect -2126 828 -2068 834
rect -1916 828 -1858 834
rect -1706 828 -1648 834
rect -1496 828 -1438 834
rect -1293 828 -1283 834
rect -1231 828 -1221 834
rect -1076 828 -1018 834
rect -866 828 -808 834
rect -656 828 -598 834
rect -446 828 -388 834
rect -236 828 -178 834
rect -26 828 32 834
rect 184 828 242 834
rect 292 828 302 834
rect 354 868 364 880
rect 394 868 452 874
rect 604 868 662 874
rect 814 868 872 874
rect 1024 868 1082 874
rect 1234 868 1292 874
rect 1444 868 1502 874
rect 1647 868 1657 880
rect 1709 868 1719 880
rect 1864 868 1922 874
rect 2074 868 2132 874
rect 2284 868 2342 874
rect 2494 868 2552 874
rect 2704 868 2762 874
rect 2907 868 2917 880
rect 2969 868 2979 880
rect 3124 868 3182 874
rect 3334 868 3392 874
rect 3544 868 3602 874
rect 3754 868 3812 874
rect 3964 868 4022 874
rect 4174 868 4232 874
rect 4384 868 4442 874
rect 4594 868 4652 874
rect 4804 868 4862 874
rect 4911 868 4921 880
rect 354 834 406 868
rect 440 834 616 868
rect 650 834 826 868
rect 860 834 1036 868
rect 1070 834 1246 868
rect 1280 834 1456 868
rect 1490 834 1657 868
rect 1709 834 1876 868
rect 1910 834 2086 868
rect 2120 834 2296 868
rect 2330 834 2506 868
rect 2540 834 2716 868
rect 2750 834 2917 868
rect 2969 834 3136 868
rect 3170 834 3346 868
rect 3380 834 3556 868
rect 3590 834 3766 868
rect 3800 834 3976 868
rect 4010 834 4186 868
rect 4220 834 4396 868
rect 4430 834 4606 868
rect 4640 834 4816 868
rect 4850 834 4921 868
rect 354 828 364 834
rect 394 828 452 834
rect 604 828 662 834
rect 814 828 872 834
rect 1024 828 1082 834
rect 1234 828 1292 834
rect 1444 828 1502 834
rect 1647 828 1657 834
rect 1709 828 1719 834
rect 1864 828 1922 834
rect 2074 828 2132 834
rect 2284 828 2342 834
rect 2494 828 2552 834
rect 2704 828 2762 834
rect 2907 828 2917 834
rect 2969 828 2979 834
rect 3124 828 3182 834
rect 3334 828 3392 834
rect 3544 828 3602 834
rect 3754 828 3812 834
rect 3964 828 4022 834
rect 4174 828 4232 834
rect 4384 828 4442 834
rect 4594 828 4652 834
rect 4804 828 4862 834
rect 4911 828 4921 834
rect 4973 868 4983 880
rect 5014 868 5072 874
rect 5224 868 5282 874
rect 5434 868 5492 874
rect 5644 868 5702 874
rect 5854 868 5912 874
rect 4973 834 5026 868
rect 5060 834 5236 868
rect 5270 834 5446 868
rect 5480 834 5656 868
rect 5690 834 5866 868
rect 5900 834 5912 868
rect 4973 828 4983 834
rect 5014 828 5072 834
rect 5224 828 5282 834
rect 5434 828 5492 834
rect 5644 828 5702 834
rect 5854 828 5912 834
rect -2845 733 -2704 745
rect -2598 741 -2588 793
rect -2536 784 -2526 793
rect -2174 784 -2116 790
rect -1761 784 -1689 793
rect -1334 784 -1276 790
rect -914 784 -856 790
rect -494 784 -436 790
rect -81 784 -9 793
rect 346 784 404 790
rect 766 784 824 790
rect 1186 784 1244 790
rect 1599 784 1671 793
rect 2026 784 2084 790
rect 2446 784 2504 790
rect 2866 784 2924 790
rect 3286 784 3344 790
rect 3706 784 3764 790
rect 4126 784 4184 790
rect 4546 784 4604 790
rect 4966 784 5024 790
rect 5386 784 5444 790
rect 5806 784 5864 790
rect -2536 750 -2162 784
rect -2128 750 -1742 784
rect -1708 750 -1322 784
rect -1288 750 -902 784
rect -868 750 -482 784
rect -448 750 -62 784
rect -28 750 358 784
rect 392 750 778 784
rect 812 750 1198 784
rect 1232 750 1618 784
rect 1652 750 2038 784
rect 2072 750 2458 784
rect 2492 750 2878 784
rect 2912 750 3298 784
rect 3332 750 3718 784
rect 3752 750 4138 784
rect 4172 750 4558 784
rect 4592 750 4978 784
rect 5012 750 5398 784
rect 5432 750 5818 784
rect 5852 750 5912 784
rect -2536 741 -2526 750
rect -2174 744 -2116 750
rect -1761 741 -1689 750
rect -1334 744 -1276 750
rect -914 744 -856 750
rect -494 744 -436 750
rect -81 741 -9 750
rect 346 744 404 750
rect 766 744 824 750
rect 1186 744 1244 750
rect 1599 741 1671 750
rect 2026 744 2084 750
rect 2446 744 2504 750
rect 2866 744 2924 750
rect 3286 744 3344 750
rect 3706 744 3764 750
rect 4126 744 4184 750
rect 4546 744 4604 750
rect 4966 744 5024 750
rect 5386 744 5444 750
rect 5806 744 5864 750
rect 6186 745 6192 4180
rect 6226 4144 6322 4180
rect 6226 4092 6229 4144
rect 6281 4092 6322 4144
rect 6226 4003 6322 4092
rect 6226 3951 6229 4003
rect 6281 3951 6322 4003
rect 6226 3862 6322 3951
rect 6226 3810 6229 3862
rect 6281 3810 6322 3862
rect 6226 3721 6322 3810
rect 6226 3669 6229 3721
rect 6281 3669 6322 3721
rect 6226 3580 6322 3669
rect 6612 3663 6682 5573
rect 6831 5403 6889 5409
rect 6750 5368 6784 5371
rect 6831 5369 6843 5403
rect 6877 5369 6889 5403
rect 6744 5356 6790 5368
rect 6831 5363 6889 5369
rect 6744 5322 6750 5356
rect 6784 5322 6790 5356
rect 6744 5310 6790 5322
rect 6750 5176 6784 5310
rect 6843 5217 6877 5363
rect 6985 5313 7019 5573
rect 6973 5307 7031 5313
rect 6973 5273 6985 5307
rect 7019 5273 7031 5307
rect 6973 5267 7031 5273
rect 7078 5272 7112 5275
rect 6831 5211 6889 5217
rect 6831 5177 6843 5211
rect 6877 5177 6889 5211
rect 6744 5173 6790 5176
rect 6729 5121 6739 5173
rect 6791 5121 6801 5173
rect 6831 5171 6889 5177
rect 6744 5118 6790 5121
rect 6750 4984 6784 5118
rect 6843 5025 6877 5171
rect 6985 5121 7019 5267
rect 7072 5260 7118 5272
rect 7072 5226 7078 5260
rect 7112 5226 7118 5260
rect 7072 5214 7118 5226
rect 7078 5173 7112 5214
rect 7060 5121 7070 5173
rect 7122 5121 7132 5173
rect 6973 5115 7031 5121
rect 6973 5081 6985 5115
rect 7019 5081 7031 5115
rect 6973 5075 7031 5081
rect 7078 5080 7112 5121
rect 6831 5019 6889 5025
rect 6831 4985 6843 5019
rect 6877 4985 6889 5019
rect 6744 4972 6790 4984
rect 6831 4979 6889 4985
rect 6744 4938 6750 4972
rect 6784 4938 6790 4972
rect 6744 4926 6790 4938
rect 6750 4792 6784 4926
rect 6843 4833 6877 4979
rect 6985 4929 7019 5075
rect 7072 5068 7118 5080
rect 7072 5034 7078 5068
rect 7112 5034 7118 5068
rect 7072 5022 7118 5034
rect 6973 4923 7031 4929
rect 6973 4889 6985 4923
rect 7019 4889 7031 4923
rect 6973 4883 7031 4889
rect 7078 4888 7112 5022
rect 6831 4827 6889 4833
rect 6831 4793 6843 4827
rect 6877 4793 6889 4827
rect 6744 4780 6790 4792
rect 6831 4787 6889 4793
rect 6744 4746 6750 4780
rect 6784 4746 6790 4780
rect 6744 4734 6790 4746
rect 6750 4600 6784 4734
rect 6843 4641 6877 4787
rect 6985 4737 7019 4883
rect 7072 4876 7118 4888
rect 7072 4842 7078 4876
rect 7112 4842 7118 4876
rect 7072 4830 7118 4842
rect 6973 4731 7031 4737
rect 6973 4697 6985 4731
rect 7019 4697 7031 4731
rect 6973 4691 7031 4697
rect 7078 4696 7112 4830
rect 6831 4635 6889 4641
rect 6831 4601 6843 4635
rect 6877 4601 6889 4635
rect 6744 4588 6790 4600
rect 6831 4595 6889 4601
rect 6744 4554 6750 4588
rect 6784 4554 6790 4588
rect 6744 4542 6790 4554
rect 6750 4408 6784 4542
rect 6843 4497 6877 4595
rect 6985 4545 7019 4691
rect 7072 4684 7118 4696
rect 7072 4650 7078 4684
rect 7112 4650 7118 4684
rect 7072 4638 7118 4650
rect 6973 4539 7031 4545
rect 6973 4505 6985 4539
rect 7019 4505 7031 4539
rect 6973 4499 7031 4505
rect 7078 4504 7112 4638
rect 6825 4445 6835 4497
rect 6887 4445 6897 4497
rect 6831 4443 6889 4445
rect 6831 4409 6843 4443
rect 6877 4409 6889 4443
rect 6744 4396 6790 4408
rect 6831 4403 6889 4409
rect 6744 4362 6750 4396
rect 6784 4362 6790 4396
rect 6744 4350 6790 4362
rect 6750 4216 6784 4350
rect 6843 4257 6877 4403
rect 6985 4353 7019 4499
rect 7072 4492 7118 4504
rect 7072 4458 7078 4492
rect 7112 4458 7118 4492
rect 7072 4446 7118 4458
rect 6973 4347 7031 4353
rect 6973 4313 6985 4347
rect 7019 4313 7031 4347
rect 6973 4307 7031 4313
rect 7078 4312 7112 4446
rect 6831 4251 6889 4257
rect 6831 4217 6843 4251
rect 6877 4217 6889 4251
rect 6744 4204 6790 4216
rect 6831 4211 6889 4217
rect 6744 4170 6750 4204
rect 6784 4170 6790 4204
rect 6744 4158 6790 4170
rect 6750 4024 6784 4158
rect 6843 4065 6877 4211
rect 6985 4161 7019 4307
rect 7072 4300 7118 4312
rect 7072 4266 7078 4300
rect 7112 4266 7118 4300
rect 7072 4254 7118 4266
rect 6973 4155 7031 4161
rect 6973 4121 6985 4155
rect 7019 4121 7031 4155
rect 6973 4115 7031 4121
rect 7078 4120 7112 4254
rect 6831 4059 6889 4065
rect 6831 4025 6843 4059
rect 6877 4025 6889 4059
rect 6744 4021 6790 4024
rect 6731 3969 6741 4021
rect 6793 3969 6803 4021
rect 6831 4019 6889 4025
rect 6744 3966 6790 3969
rect 6750 3961 6784 3966
rect 6843 3873 6877 4019
rect 6985 3969 7019 4115
rect 7072 4108 7118 4120
rect 7072 4074 7078 4108
rect 7112 4074 7118 4108
rect 7072 4062 7118 4074
rect 7078 4021 7112 4062
rect 7060 3969 7070 4021
rect 7122 3969 7132 4021
rect 6973 3963 7031 3969
rect 6973 3929 6985 3963
rect 7019 3929 7031 3963
rect 6973 3923 7031 3929
rect 7078 3928 7112 3969
rect 7072 3916 7118 3928
rect 7072 3882 7078 3916
rect 7112 3882 7118 3916
rect 6831 3867 6889 3873
rect 7072 3870 7118 3882
rect 6831 3833 6843 3867
rect 6877 3833 6889 3867
rect 7078 3865 7112 3870
rect 6831 3827 6889 3833
rect 6612 3657 7130 3663
rect 6612 3623 6744 3657
rect 7118 3623 7130 3657
rect 6612 3617 7130 3623
rect 6612 3587 6682 3617
rect 6226 3528 6229 3580
rect 6281 3528 6322 3580
rect 6226 3439 6322 3528
rect 6226 3387 6229 3439
rect 6281 3387 6322 3439
rect 6226 3298 6322 3387
rect 6226 3246 6229 3298
rect 6281 3246 6322 3298
rect 6226 3157 6322 3246
rect 6226 3105 6229 3157
rect 6281 3105 6322 3157
rect 6226 3016 6322 3105
rect 6226 2964 6229 3016
rect 6281 2964 6322 3016
rect 6226 2875 6322 2964
rect 6226 2823 6229 2875
rect 6281 2823 6322 2875
rect 6226 2734 6322 2823
rect 6226 2682 6229 2734
rect 6281 2682 6322 2734
rect 6226 1549 6322 2682
rect 6226 1497 6229 1549
rect 6281 1497 6322 1549
rect 6226 1408 6322 1497
rect 6226 1356 6229 1408
rect 6281 1356 6322 1408
rect 6226 1267 6322 1356
rect 6226 1215 6229 1267
rect 6281 1215 6322 1267
rect 6226 1126 6322 1215
rect 6226 1074 6229 1126
rect 6281 1074 6322 1126
rect 6226 985 6322 1074
rect 6226 933 6229 985
rect 6281 933 6322 985
rect 6226 844 6322 933
rect 6226 792 6229 844
rect 6281 792 6322 844
rect 6226 745 6322 792
rect 6186 733 6322 745
rect -1297 463 -1283 567
rect -1231 463 302 567
rect 354 463 1657 567
rect 1709 463 2917 567
rect 2969 463 4921 567
rect 4973 463 4983 567
rect -1297 462 4983 463
rect 270 290 328 296
rect 270 289 282 290
rect 218 256 282 289
rect 316 289 328 290
rect 462 290 520 296
rect 462 289 474 290
rect 316 256 474 289
rect 508 289 520 290
rect 654 290 712 296
rect 654 289 666 290
rect 508 256 666 289
rect 700 289 712 290
rect 846 290 904 296
rect 846 289 858 290
rect 700 256 858 289
rect 892 289 904 290
rect 1032 289 1042 303
rect 892 256 1042 289
rect 1094 289 1104 303
rect 1230 290 1288 296
rect 1230 289 1242 290
rect 1094 256 1242 289
rect 1276 289 1288 290
rect 1422 290 1480 296
rect 1422 289 1434 290
rect 1276 256 1434 289
rect 1468 289 1480 290
rect 1614 290 1672 296
rect 1614 289 1626 290
rect 1468 256 1626 289
rect 1660 289 1672 290
rect 1806 290 1864 296
rect 1806 289 1818 290
rect 1660 256 1818 289
rect 1852 289 1864 290
rect 1998 290 2056 296
rect 1998 289 2010 290
rect 1852 256 2010 289
rect 2044 289 2056 290
rect 2190 290 2248 296
rect 2190 289 2202 290
rect 2044 256 2202 289
rect 2236 289 2248 290
rect 2375 289 2385 303
rect 2236 256 2385 289
rect 2437 289 2447 303
rect 2574 290 2632 296
rect 2574 289 2586 290
rect 2437 256 2586 289
rect 2620 289 2632 290
rect 2766 290 2824 296
rect 2766 289 2778 290
rect 2620 256 2778 289
rect 2812 289 2824 290
rect 2958 290 3016 296
rect 2958 289 2970 290
rect 2812 256 2970 289
rect 3004 289 3016 290
rect 3150 290 3208 296
rect 3150 289 3162 290
rect 3004 256 3162 289
rect 3196 256 3208 290
rect 218 255 1042 256
rect 270 250 328 255
rect 462 250 520 255
rect 654 250 712 255
rect 846 250 904 255
rect 1032 251 1042 255
rect 1094 255 2385 256
rect 1094 251 1104 255
rect 1038 250 1096 251
rect 1230 250 1288 255
rect 1422 250 1480 255
rect 1614 250 1672 255
rect 1806 250 1864 255
rect 1998 250 2056 255
rect 2190 250 2248 255
rect 2375 251 2385 255
rect 2437 255 3208 256
rect 2437 251 2447 255
rect 2382 250 2440 251
rect 2574 250 2632 255
rect 2766 250 2824 255
rect 2958 250 3016 255
rect 3150 250 3208 255
rect 174 205 232 211
rect 292 205 302 211
rect 174 171 186 205
rect 220 171 302 205
rect 174 165 232 171
rect 292 159 302 171
rect 354 205 424 211
rect 558 205 616 211
rect 750 205 808 211
rect 942 205 1000 211
rect 1134 205 1192 211
rect 1326 205 1384 211
rect 1518 205 1576 211
rect 1647 205 1657 211
rect 354 171 378 205
rect 412 171 570 205
rect 604 171 762 205
rect 796 171 954 205
rect 988 171 1146 205
rect 1180 171 1338 205
rect 1372 171 1530 205
rect 1564 171 1657 205
rect 354 165 424 171
rect 558 165 616 171
rect 750 165 808 171
rect 942 165 1000 171
rect 1134 165 1192 171
rect 1326 165 1384 171
rect 1518 165 1576 171
rect 354 159 364 165
rect 1647 159 1657 171
rect 1709 205 1768 211
rect 1902 205 1960 211
rect 2094 205 2152 211
rect 2286 205 2344 211
rect 2478 205 2536 211
rect 2670 205 2728 211
rect 2862 205 2917 211
rect 1709 171 1722 205
rect 1756 171 1914 205
rect 1948 171 2106 205
rect 2140 171 2298 205
rect 2332 171 2490 205
rect 2524 171 2682 205
rect 2716 171 2874 205
rect 2908 171 2917 205
rect 1709 165 1768 171
rect 1902 165 1960 171
rect 2094 165 2152 171
rect 2286 165 2344 171
rect 2478 165 2536 171
rect 2670 165 2728 171
rect 2862 165 2917 171
rect 1709 159 1719 165
rect 2907 159 2917 165
rect 2969 205 2979 211
rect 3054 205 3112 211
rect 3246 205 3304 211
rect 2969 171 3066 205
rect 3100 171 3258 205
rect 3292 171 3304 205
rect 2969 159 2979 171
rect 3054 165 3112 171
rect 3246 165 3304 171
rect 270 63 328 69
rect 462 63 520 69
rect 654 63 712 69
rect 846 63 904 69
rect 1038 63 1096 69
rect 1230 63 1288 69
rect 1422 63 1480 69
rect 1614 63 1672 69
rect 1806 63 1864 69
rect 1998 63 2056 69
rect 2190 63 2248 69
rect 2382 63 2440 69
rect 2574 63 2632 69
rect 2766 63 2824 69
rect 2958 63 3016 69
rect 3150 63 3208 69
rect 270 29 282 63
rect 316 29 474 63
rect 508 29 666 63
rect 700 29 858 63
rect 892 29 1050 63
rect 1084 29 1242 63
rect 1276 29 1434 63
rect 1468 29 1626 63
rect 1660 29 1818 63
rect 1852 29 2010 63
rect 2044 29 2202 63
rect 2236 29 2394 63
rect 2428 29 2586 63
rect 2620 29 2778 63
rect 2812 29 2970 63
rect 3004 29 3162 63
rect 3196 29 3208 63
rect 270 23 328 29
rect 462 23 520 29
rect 654 23 712 29
rect 846 23 904 29
rect 1038 23 1096 29
rect 1230 23 1288 29
rect 1422 23 1480 29
rect 1614 23 1672 29
rect 1806 23 1864 29
rect 1998 23 2056 29
rect 2190 23 2248 29
rect 2382 23 2440 29
rect 2574 23 2632 29
rect 2766 23 2824 29
rect 2958 23 3016 29
rect 3150 23 3208 29
rect -3246 -114 6607 -82
rect -3246 -115 5523 -114
rect -3246 -167 -2798 -115
rect -2746 -167 -2657 -115
rect -2605 -167 -2516 -115
rect -2464 -167 -2375 -115
rect -2323 -167 -2234 -115
rect -2182 -167 -2093 -115
rect -2041 -123 5523 -115
rect -2041 -157 72 -123
rect 3406 -157 5523 -123
rect -2041 -166 5523 -157
rect 5575 -166 5664 -114
rect 5716 -166 5805 -114
rect 5857 -166 5946 -114
rect 5998 -166 6087 -114
rect 6139 -166 6228 -114
rect 6280 -166 6607 -114
rect -2041 -167 6607 -166
rect -3246 -193 6607 -167
<< via1 >>
rect 1156 9776 1208 9790
rect 1156 9742 1165 9776
rect 1165 9742 1199 9776
rect 1199 9742 1208 9776
rect 1156 9738 1208 9742
rect 1156 9597 1208 9649
rect 1156 9500 1208 9508
rect 1156 9466 1165 9500
rect 1165 9466 1199 9500
rect 1199 9466 1208 9500
rect 1156 9456 1208 9466
rect 1156 9316 1208 9367
rect 1156 9315 1165 9316
rect 1165 9315 1199 9316
rect 1199 9315 1208 9316
rect 1156 9224 1208 9226
rect 1156 9190 1165 9224
rect 1165 9190 1199 9224
rect 1199 9190 1208 9224
rect 1156 9174 1208 9190
rect 1576 9268 1628 9320
rect 2003 9364 2055 9372
rect 2003 9330 2016 9364
rect 2016 9330 2050 9364
rect 2050 9330 2055 9364
rect 2003 9320 2055 9330
rect 1397 9102 1449 9154
rect 2003 9258 2055 9268
rect 2003 9224 2015 9258
rect 2015 9224 2049 9258
rect 2049 9224 2055 9258
rect 2003 9216 2055 9224
rect 1823 9102 1875 9154
rect 1487 8982 1539 8991
rect 1487 8948 1497 8982
rect 1497 8948 1531 8982
rect 1531 8948 1539 8982
rect 1487 8939 1539 8948
rect 1576 8982 1628 8991
rect 1576 8948 1599 8982
rect 1599 8948 1628 8982
rect 1576 8939 1628 8948
rect 2244 9776 2296 9792
rect 2244 9742 2253 9776
rect 2253 9742 2287 9776
rect 2287 9742 2296 9776
rect 2244 9740 2296 9742
rect 2244 9650 2253 9651
rect 2253 9650 2287 9651
rect 2287 9650 2296 9651
rect 2244 9599 2296 9650
rect 2244 9500 2296 9510
rect 2244 9466 2253 9500
rect 2253 9466 2287 9500
rect 2287 9466 2296 9500
rect 2244 9458 2296 9466
rect 2244 9317 2296 9369
rect 2244 9224 2296 9228
rect 2244 9190 2253 9224
rect 2253 9190 2287 9224
rect 2287 9190 2296 9224
rect 2244 9176 2296 9190
rect 1823 8982 1875 8991
rect 1823 8948 1854 8982
rect 1854 8948 1875 8982
rect 1823 8939 1875 8948
rect 1912 8982 1964 8991
rect 1912 8948 1921 8982
rect 1921 8948 1955 8982
rect 1955 8948 1964 8982
rect 1912 8939 1964 8948
rect 1389 8312 1441 8322
rect 1389 8278 1397 8312
rect 1397 8278 1431 8312
rect 1431 8278 1441 8312
rect 1389 8270 1441 8278
rect 2013 8313 2065 8323
rect 2013 8279 2022 8313
rect 2022 8279 2056 8313
rect 2056 8279 2065 8313
rect 2013 8271 2065 8279
rect -1286 8023 -1234 8041
rect 287 8023 339 8041
rect 3230 8023 3282 8041
rect 4699 8023 4751 8041
rect -1286 7989 -1234 8023
rect 287 7989 339 8023
rect 3230 7989 3282 8023
rect 4699 7989 4751 8023
rect -3662 7529 -3610 7581
rect -3331 7574 -3279 7581
rect -3331 7540 -3322 7574
rect -3322 7540 -3288 7574
rect -3288 7540 -3279 7574
rect -3331 7529 -3279 7540
rect -3423 6668 -3371 6720
rect -3660 6379 -3608 6431
rect -3331 6422 -3279 6431
rect -3331 6388 -3322 6422
rect -3322 6388 -3288 6422
rect -3288 6388 -3279 6422
rect -3331 6379 -3279 6388
rect 1970 7878 2022 7930
rect -1286 7776 -1234 7828
rect 287 7794 296 7828
rect 296 7794 330 7828
rect 330 7794 339 7828
rect 3230 7794 3236 7828
rect 3236 7794 3270 7828
rect 3270 7794 3282 7828
rect 4699 7794 4706 7828
rect 4706 7794 4740 7828
rect 4740 7794 4751 7828
rect 287 7776 339 7794
rect 3230 7776 3282 7794
rect 4699 7776 4751 7794
rect 2401 7652 2453 7704
rect 3871 7652 3923 7704
rect 5340 7652 5392 7704
rect 1970 7550 2022 7602
rect 1458 7348 1510 7400
rect -1286 7244 -1234 7296
rect 287 7262 298 7296
rect 298 7262 332 7296
rect 332 7262 339 7296
rect 3230 7262 3238 7296
rect 3238 7262 3272 7296
rect 3272 7262 3282 7296
rect 4699 7262 4708 7296
rect 4708 7262 4742 7296
rect 4742 7262 4751 7296
rect 287 7244 339 7262
rect 3230 7244 3282 7262
rect 4699 7244 4751 7262
rect -2009 7120 -1957 7172
rect -539 7120 -487 7172
rect 931 7120 983 7172
rect 1458 7018 1510 7070
rect 931 6793 983 6845
rect 1970 6793 2022 6845
rect -3072 6668 -3020 6720
rect -2009 6668 -1957 6720
rect -1379 6668 -1327 6720
rect -539 6668 -487 6720
rect 301 6668 353 6720
rect 931 6668 983 6720
rect 2401 6668 2453 6720
rect 3031 6668 3083 6720
rect 3871 6668 3923 6720
rect 4711 6668 4763 6720
rect 5340 6668 5392 6720
rect 6482 6668 6534 6720
rect 1458 6536 1510 6588
rect 2401 6536 2453 6588
rect -3660 5121 -3608 5173
rect -3329 5164 -3277 5173
rect -3329 5130 -3320 5164
rect -3320 5130 -3286 5164
rect -3286 5130 -3277 5164
rect -3329 5121 -3277 5130
rect -3425 4445 -3373 4497
rect -3660 3969 -3608 4021
rect -3331 4012 -3279 4021
rect -3331 3978 -3320 4012
rect -3320 3978 -3286 4012
rect -3286 3978 -3279 4012
rect -3331 3969 -3279 3978
rect -2798 6360 -2746 6412
rect -2798 6219 -2746 6271
rect -2798 6078 -2746 6130
rect -2798 5937 -2746 5989
rect -2798 5796 -2746 5848
rect -2798 5655 -2746 5707
rect -2798 5514 -2746 5566
rect -2798 5373 -2746 5425
rect -2798 5232 -2746 5284
rect -2798 5091 -2746 5143
rect -2798 4950 -2746 5002
rect -2798 4809 -2746 4861
rect 1970 6386 2022 6438
rect 3031 6311 3040 6345
rect 3040 6311 3074 6345
rect 3074 6311 3083 6345
rect 4711 6311 4720 6345
rect 4720 6311 4754 6345
rect 4754 6311 4763 6345
rect 3031 6293 3083 6311
rect 4711 6293 4763 6311
rect 2401 6169 2453 6221
rect 3871 6169 3923 6221
rect 5340 6169 5392 6221
rect 1970 6076 2022 6128
rect 1458 5946 1510 5998
rect -1379 5871 -1370 5905
rect -1370 5871 -1336 5905
rect -1336 5871 -1327 5905
rect 301 5871 310 5905
rect 310 5871 344 5905
rect 344 5871 353 5905
rect -1379 5853 -1327 5871
rect 301 5853 353 5871
rect -2009 5729 -1957 5781
rect -539 5729 -487 5781
rect 931 5729 983 5781
rect 1458 5634 1510 5686
rect 1458 5506 1510 5558
rect -1379 5431 -1370 5465
rect -1370 5431 -1336 5465
rect -1336 5431 -1327 5465
rect 301 5431 310 5465
rect 310 5431 344 5465
rect 344 5431 353 5465
rect -1379 5413 -1327 5431
rect 301 5413 353 5431
rect -2009 5289 -1957 5341
rect -539 5289 -487 5341
rect 931 5289 983 5341
rect 1458 5193 1510 5245
rect 1970 5067 2022 5119
rect 3031 4991 3040 5025
rect 3040 4991 3074 5025
rect 3074 4991 3083 5025
rect 4711 4991 4720 5025
rect 4720 4991 4754 5025
rect 4754 4991 4763 5025
rect 3031 4973 3083 4991
rect 4711 4973 4763 4991
rect 2401 4849 2453 4901
rect 3871 4849 3923 4901
rect 5340 4849 5392 4901
rect 1970 4756 2022 4808
rect 6229 6360 6281 6412
rect 6229 6219 6281 6271
rect 6229 6078 6281 6130
rect 6229 5937 6281 5989
rect 6229 5796 6281 5848
rect 6229 5655 6281 5707
rect 6229 5514 6281 5566
rect 6229 5373 6281 5425
rect 6229 5232 6281 5284
rect 6229 5091 6281 5143
rect 6229 4950 6281 5002
rect 6229 4809 6281 4861
rect 6741 7574 6793 7581
rect 6741 7540 6750 7574
rect 6750 7540 6784 7574
rect 6784 7540 6793 7574
rect 6741 7529 6793 7540
rect 7072 7529 7124 7581
rect 6833 6668 6885 6720
rect 6741 6422 6793 6431
rect 6741 6388 6750 6422
rect 6750 6388 6784 6422
rect 6784 6388 6793 6422
rect 6741 6379 6793 6388
rect 7070 6379 7122 6431
rect -3072 4445 -3020 4497
rect -2009 4445 -1957 4497
rect -539 4445 -487 4497
rect 931 4445 983 4497
rect 2401 4445 2453 4497
rect 3871 4445 3923 4497
rect 5340 4445 5392 4497
rect 6482 4445 6534 4497
rect -2798 4092 -2746 4144
rect -2798 3951 -2746 4003
rect -2798 3810 -2746 3862
rect -2798 3669 -2746 3721
rect -2798 3528 -2746 3580
rect -2798 3387 -2746 3439
rect -2798 3246 -2746 3298
rect -2798 3105 -2746 3157
rect -2798 2964 -2746 3016
rect -2798 2823 -2746 2875
rect -2798 2682 -2746 2734
rect -2798 1497 -2746 1549
rect -2798 1356 -2746 1408
rect -2798 1215 -2746 1267
rect -2798 1074 -2746 1126
rect -2798 933 -2746 985
rect -2798 792 -2746 844
rect -2588 4131 -2536 4183
rect -539 4090 -487 4096
rect -2009 4056 -2000 4090
rect -2000 4056 -1966 4090
rect -1966 4056 -1957 4090
rect -539 4056 -530 4090
rect -530 4056 -496 4090
rect -496 4056 -487 4090
rect 931 4056 940 4090
rect 940 4056 974 4090
rect 974 4056 983 4090
rect -2009 4038 -1957 4056
rect -539 4044 -487 4056
rect 931 4038 983 4056
rect -1283 3948 -1231 3960
rect -1283 3914 -1274 3948
rect -1274 3914 -1240 3948
rect -1240 3914 -1231 3948
rect -1283 3908 -1231 3914
rect 302 3908 354 3960
rect 1657 3948 1709 3960
rect 2917 3948 2969 3960
rect 1657 3914 1666 3948
rect 1666 3914 1700 3948
rect 1700 3914 1709 3948
rect 2917 3914 2926 3948
rect 2926 3914 2960 3948
rect 2960 3914 2969 3948
rect 1657 3908 1709 3914
rect 2917 3908 2969 3914
rect 4921 3908 4973 3960
rect -2588 3821 -2536 3873
rect 6020 3691 6072 3743
rect 2401 3616 2410 3650
rect 2410 3616 2444 3650
rect 2444 3616 2453 3650
rect 3871 3616 3880 3650
rect 3880 3616 3914 3650
rect 3914 3616 3923 3650
rect 5340 3616 5350 3650
rect 5350 3616 5384 3650
rect 5384 3616 5392 3650
rect 2401 3598 2453 3616
rect 3871 3598 3923 3616
rect 5340 3598 5392 3616
rect -1283 3508 -1231 3520
rect -1283 3474 -1274 3508
rect -1274 3474 -1240 3508
rect -1240 3474 -1231 3508
rect -1283 3468 -1231 3474
rect 302 3468 354 3520
rect 1657 3508 1709 3520
rect 2917 3508 2969 3520
rect 1657 3474 1666 3508
rect 1666 3474 1700 3508
rect 1700 3474 1709 3508
rect 2917 3474 2926 3508
rect 2926 3474 2960 3508
rect 2960 3474 2969 3508
rect 1657 3468 1709 3474
rect 2917 3468 2969 3474
rect 4921 3468 4973 3520
rect 6020 3381 6072 3433
rect 6020 3253 6072 3305
rect 2401 3176 2410 3210
rect 2410 3176 2444 3210
rect 2444 3176 2453 3210
rect 3871 3176 3880 3210
rect 3880 3176 3914 3210
rect 3914 3176 3923 3210
rect 5340 3176 5350 3210
rect 5350 3176 5384 3210
rect 5384 3176 5392 3210
rect 2401 3158 2453 3176
rect 3871 3158 3923 3176
rect 5340 3158 5392 3176
rect -1283 3068 -1231 3080
rect -1283 3034 -1274 3068
rect -1274 3034 -1240 3068
rect -1240 3034 -1231 3068
rect -1283 3028 -1231 3034
rect 302 3028 354 3080
rect 1657 3068 1709 3080
rect 2917 3068 2969 3080
rect 1657 3034 1666 3068
rect 1666 3034 1700 3068
rect 1700 3034 1709 3068
rect 2917 3034 2926 3068
rect 2926 3034 2960 3068
rect 2960 3034 2969 3068
rect 1657 3028 1709 3034
rect 2917 3028 2969 3034
rect 4921 3028 4973 3080
rect 6020 2939 6072 2991
rect -2588 2811 -2536 2863
rect -539 2770 -487 2776
rect -2009 2736 -2000 2770
rect -2000 2736 -1966 2770
rect -1966 2736 -1957 2770
rect -539 2736 -530 2770
rect -530 2736 -496 2770
rect -496 2736 -487 2770
rect 931 2736 940 2770
rect 940 2736 974 2770
rect 974 2736 983 2770
rect -2009 2718 -1957 2736
rect -539 2724 -487 2736
rect 931 2718 983 2736
rect -1283 2628 -1231 2640
rect -1283 2594 -1274 2628
rect -1274 2594 -1240 2628
rect -1240 2594 -1231 2628
rect -1283 2588 -1231 2594
rect 302 2588 354 2640
rect 1657 2628 1709 2640
rect 2917 2628 2969 2640
rect 1657 2594 1666 2628
rect 1666 2594 1700 2628
rect 1700 2594 1709 2628
rect 2917 2594 2926 2628
rect 2926 2594 2960 2628
rect 2960 2594 2969 2628
rect 1657 2588 1709 2594
rect 2917 2588 2969 2594
rect 4921 2588 4973 2640
rect -2588 2501 -2536 2553
rect -2588 2372 -2536 2424
rect -539 2330 -487 2336
rect -2009 2296 -2000 2330
rect -2000 2296 -1966 2330
rect -1966 2296 -1957 2330
rect -539 2296 -530 2330
rect -530 2296 -496 2330
rect -496 2296 -487 2330
rect 931 2296 940 2330
rect 940 2296 974 2330
rect 974 2296 983 2330
rect -2009 2278 -1957 2296
rect -539 2284 -487 2296
rect 931 2278 983 2296
rect -1283 2188 -1231 2200
rect -1283 2154 -1274 2188
rect -1274 2154 -1240 2188
rect -1240 2154 -1231 2188
rect -1283 2148 -1231 2154
rect 302 2148 354 2200
rect 1657 2188 1709 2200
rect 2917 2188 2969 2200
rect 1657 2154 1666 2188
rect 1666 2154 1700 2188
rect 1700 2154 1709 2188
rect 2917 2154 2926 2188
rect 2926 2154 2960 2188
rect 2960 2154 2969 2188
rect 1657 2148 1709 2154
rect 2917 2148 2969 2154
rect 4921 2148 4973 2200
rect -2588 2061 -2536 2113
rect 6020 1933 6072 1985
rect 2401 1856 2410 1890
rect 2410 1856 2444 1890
rect 2444 1856 2453 1890
rect 3871 1856 3880 1890
rect 3880 1856 3914 1890
rect 3914 1856 3923 1890
rect 5340 1856 5350 1890
rect 5350 1856 5384 1890
rect 5384 1856 5392 1890
rect 2401 1838 2453 1856
rect 3871 1838 3923 1856
rect 5340 1838 5392 1856
rect -1283 1748 -1231 1760
rect -1283 1714 -1274 1748
rect -1274 1714 -1240 1748
rect -1240 1714 -1231 1748
rect -1283 1708 -1231 1714
rect 302 1708 354 1760
rect 1657 1748 1709 1760
rect 2917 1748 2969 1760
rect 1657 1714 1666 1748
rect 1666 1714 1700 1748
rect 1700 1714 1709 1748
rect 2917 1714 2926 1748
rect 2926 1714 2960 1748
rect 2960 1714 2969 1748
rect 1657 1708 1709 1714
rect 2917 1708 2969 1714
rect 4921 1708 4973 1760
rect 6020 1619 6072 1671
rect 6020 1492 6072 1544
rect 2401 1416 2410 1450
rect 2410 1416 2444 1450
rect 2444 1416 2453 1450
rect 3871 1416 3880 1450
rect 3880 1416 3914 1450
rect 3914 1416 3923 1450
rect 5340 1416 5350 1450
rect 5350 1416 5384 1450
rect 5384 1416 5392 1450
rect 2401 1398 2453 1416
rect 3871 1398 3923 1416
rect 5340 1398 5392 1416
rect -1283 1308 -1231 1320
rect -1283 1274 -1274 1308
rect -1274 1274 -1240 1308
rect -1240 1274 -1231 1308
rect -1283 1268 -1231 1274
rect 302 1268 354 1320
rect 1657 1308 1709 1320
rect 2917 1308 2969 1320
rect 1657 1274 1666 1308
rect 1666 1274 1700 1308
rect 1700 1274 1709 1308
rect 2917 1274 2926 1308
rect 2926 1274 2960 1308
rect 2960 1274 2969 1308
rect 1657 1268 1709 1274
rect 2917 1268 2969 1274
rect 4921 1268 4973 1320
rect 6020 1181 6072 1233
rect -2588 1051 -2536 1103
rect -539 1010 -487 1016
rect -2009 976 -2000 1010
rect -2000 976 -1966 1010
rect -1966 976 -1957 1010
rect -539 976 -530 1010
rect -530 976 -496 1010
rect -496 976 -487 1010
rect 931 976 940 1010
rect 940 976 974 1010
rect 974 976 983 1010
rect -2009 958 -1957 976
rect -539 964 -487 976
rect 931 958 983 976
rect -1283 868 -1231 880
rect -1283 834 -1274 868
rect -1274 834 -1240 868
rect -1240 834 -1231 868
rect -1283 828 -1231 834
rect 302 828 354 880
rect 1657 868 1709 880
rect 2917 868 2969 880
rect 1657 834 1666 868
rect 1666 834 1700 868
rect 1700 834 1709 868
rect 2917 834 2926 868
rect 2926 834 2960 868
rect 2960 834 2969 868
rect 1657 828 1709 834
rect 2917 828 2969 834
rect 4921 828 4973 880
rect -2588 741 -2536 793
rect 6229 4092 6281 4144
rect 6229 3951 6281 4003
rect 6229 3810 6281 3862
rect 6229 3669 6281 3721
rect 6739 5164 6791 5173
rect 6739 5130 6750 5164
rect 6750 5130 6784 5164
rect 6784 5130 6791 5164
rect 6739 5121 6791 5130
rect 7070 5121 7122 5173
rect 6835 4445 6887 4497
rect 6741 4012 6793 4021
rect 6741 3978 6750 4012
rect 6750 3978 6784 4012
rect 6784 3978 6793 4012
rect 6741 3969 6793 3978
rect 7070 3969 7122 4021
rect 6229 3528 6281 3580
rect 6229 3387 6281 3439
rect 6229 3246 6281 3298
rect 6229 3105 6281 3157
rect 6229 2964 6281 3016
rect 6229 2823 6281 2875
rect 6229 2682 6281 2734
rect 6229 1497 6281 1549
rect 6229 1356 6281 1408
rect 6229 1215 6281 1267
rect 6229 1074 6281 1126
rect 6229 933 6281 985
rect 6229 792 6281 844
rect -1283 463 -1231 567
rect 302 463 354 567
rect 1657 463 1709 567
rect 2917 463 2969 567
rect 4921 463 4973 567
rect 1042 290 1094 303
rect 1042 256 1050 290
rect 1050 256 1084 290
rect 1084 256 1094 290
rect 2385 290 2437 303
rect 2385 256 2394 290
rect 2394 256 2428 290
rect 2428 256 2437 290
rect 1042 251 1094 256
rect 2385 251 2437 256
rect 302 159 354 211
rect 1657 159 1709 211
rect 2917 159 2969 211
rect -2798 -167 -2746 -115
rect -2657 -167 -2605 -115
rect -2516 -167 -2464 -115
rect -2375 -167 -2323 -115
rect -2234 -167 -2182 -115
rect -2093 -167 -2041 -115
rect 5523 -166 5575 -114
rect 5664 -166 5716 -114
rect 5805 -166 5857 -114
rect 5946 -166 5998 -114
rect 6087 -166 6139 -114
rect 6228 -166 6280 -114
<< metal2 >>
rect 1134 9790 1230 9800
rect 1134 9738 1156 9790
rect 1208 9738 1230 9790
rect 1134 9649 1230 9738
rect 1134 9597 1156 9649
rect 1208 9597 1230 9649
rect 1134 9553 1230 9597
rect -2845 9508 1230 9553
rect -2845 9456 1156 9508
rect 1208 9456 1230 9508
rect -2845 9412 1230 9456
rect -3662 7581 -3610 7591
rect -3331 7581 -3279 7591
rect -3610 7529 -3331 7581
rect -3662 7519 -3608 7529
rect -3331 7519 -3279 7529
rect -3660 6431 -3608 7519
rect -3423 6720 -3371 6730
rect -3072 6720 -3020 6730
rect -3427 6668 -3423 6720
rect -3371 6668 -3072 6720
rect -3020 6668 -3010 6720
rect -3423 6658 -3371 6668
rect -3072 6658 -3020 6668
rect -3331 6431 -3279 6441
rect -3608 6379 -3331 6431
rect -3660 5871 -3608 6379
rect -3331 6369 -3279 6379
rect -2845 6412 -2704 9412
rect 1134 9367 1230 9412
rect 2222 9792 2318 9802
rect 2222 9740 2244 9792
rect 2296 9740 2318 9792
rect 2222 9651 2318 9740
rect 2222 9599 2244 9651
rect 2296 9599 2318 9651
rect 2222 9552 2318 9599
rect 2222 9510 6322 9552
rect 2222 9458 2244 9510
rect 2296 9458 6322 9510
rect 2222 9416 6322 9458
rect 1134 9315 1156 9367
rect 1208 9315 1230 9367
rect 2003 9372 2055 9382
rect 1134 9226 1230 9315
rect 1576 9320 1628 9330
rect 1628 9268 2055 9320
rect 1576 9258 1628 9268
rect 1134 9174 1156 9226
rect 1208 9174 1230 9226
rect 2003 9206 2055 9216
rect 2222 9369 2318 9416
rect 2222 9317 2244 9369
rect 2296 9317 2318 9369
rect 2222 9228 2318 9317
rect 1134 9164 1230 9174
rect 2222 9176 2244 9228
rect 2296 9176 2318 9228
rect 2222 9166 2318 9176
rect 1397 9154 1449 9164
rect 1823 9154 1875 9164
rect 1449 9102 1823 9154
rect 1397 9092 1449 9102
rect 1823 9092 1875 9102
rect 1487 8991 1628 9001
rect 1539 8939 1576 8991
rect 1487 8929 1539 8939
rect 1576 8929 1628 8939
rect 1823 8991 1875 9001
rect 1912 8991 1964 9001
rect 1875 8939 1912 8991
rect 1823 8929 1875 8939
rect 1912 8929 1964 8939
rect 1389 8322 1441 8332
rect 2013 8323 2065 8333
rect 1379 8270 1389 8322
rect 1441 8270 1510 8322
rect 1389 8260 1510 8270
rect -1286 8041 -1234 8051
rect -1286 7828 -1234 7989
rect -1286 7296 -1234 7776
rect -1286 7234 -1234 7244
rect 287 8041 339 8051
rect 287 7828 339 7989
rect 287 7296 339 7776
rect 287 7234 339 7244
rect 1458 7400 1510 8260
rect -2009 7172 -1957 7182
rect -2009 6720 -1957 7120
rect -539 7172 -487 7182
rect -2009 6652 -1957 6668
rect -1379 6720 -1327 6727
rect -2845 6360 -2798 6412
rect -2746 6360 -2704 6412
rect -2845 6271 -2704 6360
rect -2845 6219 -2798 6271
rect -2746 6219 -2704 6271
rect -2845 6130 -2704 6219
rect -2845 6078 -2798 6130
rect -2746 6078 -2704 6130
rect -2845 5989 -2704 6078
rect -2845 5937 -2798 5989
rect -2746 5937 -2704 5989
rect -3667 5861 -3603 5871
rect -3667 5787 -3603 5797
rect -2845 5848 -2704 5937
rect -2845 5796 -2798 5848
rect -2746 5796 -2704 5848
rect -1379 5905 -1327 6668
rect -539 6720 -487 7120
rect 931 7172 983 7182
rect 931 6845 983 7120
rect -539 6652 -487 6668
rect 301 6720 353 6730
rect -3660 5173 -3608 5787
rect -2845 5707 -2704 5796
rect -2845 5655 -2798 5707
rect -2746 5655 -2704 5707
rect -2845 5566 -2704 5655
rect -2845 5514 -2798 5566
rect -2746 5514 -2704 5566
rect -2845 5425 -2704 5514
rect -2845 5373 -2798 5425
rect -2746 5373 -2704 5425
rect -2845 5284 -2704 5373
rect -2845 5232 -2798 5284
rect -2746 5232 -2704 5284
rect -3329 5173 -3277 5183
rect -3608 5121 -3329 5173
rect -3660 4021 -3608 5121
rect -3329 5111 -3277 5121
rect -2845 5143 -2704 5232
rect -2845 5091 -2798 5143
rect -2746 5091 -2704 5143
rect -2845 5002 -2704 5091
rect -2845 4950 -2798 5002
rect -2746 4950 -2704 5002
rect -2845 4861 -2704 4950
rect -2845 4809 -2798 4861
rect -2746 4809 -2704 4861
rect -3425 4497 -3373 4507
rect -3072 4497 -3020 4507
rect -3427 4445 -3425 4497
rect -3373 4445 -3072 4497
rect -3020 4445 -3010 4497
rect -3425 4435 -3373 4445
rect -3072 4435 -3020 4445
rect -2845 4144 -2704 4809
rect -2009 5781 -1957 5796
rect -2009 5341 -1957 5729
rect -1379 5465 -1327 5853
rect 301 5905 353 6668
rect 931 6720 983 6793
rect 931 6652 983 6668
rect 1458 7070 1510 7348
rect -1379 5403 -1327 5413
rect -539 5781 -487 5791
rect -2009 4497 -1957 5289
rect -2845 4092 -2798 4144
rect -2746 4092 -2704 4144
rect -3331 4021 -3279 4031
rect -3608 3969 -3331 4021
rect -3660 3959 -3608 3969
rect -3331 3959 -3279 3969
rect -2845 4003 -2704 4092
rect -2845 3951 -2798 4003
rect -2746 3951 -2704 4003
rect -2845 3862 -2704 3951
rect -2845 3810 -2798 3862
rect -2746 3810 -2704 3862
rect -2845 3721 -2704 3810
rect -2845 3669 -2798 3721
rect -2746 3669 -2704 3721
rect -2845 3580 -2704 3669
rect -2845 3528 -2798 3580
rect -2746 3528 -2704 3580
rect -2845 3439 -2704 3528
rect -2845 3387 -2798 3439
rect -2746 3387 -2704 3439
rect -2845 3298 -2704 3387
rect -2845 3246 -2798 3298
rect -2746 3246 -2704 3298
rect -2845 3157 -2704 3246
rect -2845 3105 -2798 3157
rect -2746 3105 -2704 3157
rect -2845 3016 -2704 3105
rect -2845 2964 -2798 3016
rect -2746 2964 -2704 3016
rect -2845 2875 -2704 2964
rect -2845 2823 -2798 2875
rect -2746 2823 -2704 2875
rect -2845 2734 -2704 2823
rect -2845 2682 -2798 2734
rect -2746 2682 -2704 2734
rect -2845 2672 -2704 2682
rect -2588 4183 -2536 4193
rect -2588 3873 -2536 4131
rect -2588 2863 -2536 3821
rect -2588 2553 -2536 2811
rect -2588 2424 -2536 2501
rect -2588 2113 -2536 2372
rect -2845 1549 -2704 1559
rect -2845 1497 -2798 1549
rect -2746 1497 -2704 1549
rect -2845 1408 -2704 1497
rect -2845 1356 -2798 1408
rect -2746 1356 -2704 1408
rect -2845 1267 -2704 1356
rect -2845 1215 -2798 1267
rect -2746 1215 -2704 1267
rect -2845 1126 -2704 1215
rect -2845 1074 -2798 1126
rect -2746 1074 -2704 1126
rect -2845 985 -2704 1074
rect -2845 933 -2798 985
rect -2746 933 -2704 985
rect -2845 844 -2704 933
rect -2845 792 -2798 844
rect -2746 792 -2704 844
rect -2845 -52 -2704 792
rect -2588 1103 -2536 2061
rect -2588 793 -2536 1051
rect -2009 4090 -1957 4445
rect -2009 2770 -1957 4038
rect -539 5341 -487 5729
rect 301 5465 353 5853
rect 1458 6588 1510 7018
rect 1458 5998 1510 6536
rect 301 5403 353 5413
rect 931 5781 983 5794
rect -539 4497 -487 5289
rect -539 4096 -487 4445
rect -2009 2330 -1957 2718
rect -2009 1010 -1957 2278
rect -2009 948 -1957 958
rect -1283 3960 -1231 3970
rect -1283 3520 -1231 3908
rect -1283 3080 -1231 3468
rect -1283 2640 -1231 3028
rect -1283 2200 -1231 2588
rect -1283 1760 -1231 2148
rect -1283 1320 -1231 1708
rect -2588 731 -2536 741
rect -1283 880 -1231 1268
rect -539 2776 -487 4044
rect 931 5341 983 5729
rect 931 4497 983 5289
rect 1458 5686 1510 5946
rect 1458 5558 1510 5634
rect 1458 5245 1510 5506
rect 1458 5183 1510 5193
rect 1970 8271 2013 8323
rect 2065 8271 2071 8323
rect 1970 8261 2065 8271
rect 1970 7930 2022 8261
rect 1970 7602 2022 7878
rect 3230 8041 3282 8051
rect 3230 7828 3282 7989
rect 1970 6845 2022 7550
rect 1970 6438 2022 6793
rect 2401 7704 2453 7711
rect 2401 6720 2453 7652
rect 3230 7296 3282 7776
rect 4699 8041 4751 8051
rect 4699 7828 4751 7989
rect 3230 7234 3282 7244
rect 3871 7704 3923 7714
rect 2401 6588 2453 6668
rect 2401 6526 2453 6536
rect 3031 6720 3083 6730
rect 1970 6128 2022 6386
rect 3031 6345 3083 6668
rect 3871 6720 3923 7652
rect 4699 7296 4751 7776
rect 4699 7234 4751 7244
rect 5340 7704 5392 7714
rect 3871 6657 3923 6668
rect 4711 6720 4763 6730
rect 1970 5119 2022 6076
rect 1970 4808 2022 5067
rect 1970 4746 2022 4756
rect 2401 6221 2453 6240
rect 2401 4901 2453 6169
rect 3031 5025 3083 6293
rect 4711 6345 4763 6668
rect 5340 6720 5392 7652
rect 5340 6657 5392 6668
rect 3031 4963 3083 4973
rect 3871 6221 3923 6236
rect 931 4090 983 4445
rect -539 2336 -487 2724
rect -539 1016 -487 2284
rect -539 954 -487 964
rect 302 3960 354 3970
rect 302 3520 354 3908
rect 302 3080 354 3468
rect 302 2640 354 3028
rect 302 2200 354 2588
rect 302 1760 354 2148
rect 302 1320 354 1708
rect -1283 567 -1231 828
rect -1283 457 -1231 463
rect 302 880 354 1268
rect 931 2770 983 4038
rect 2401 4497 2453 4849
rect 931 2330 983 2718
rect 931 1010 983 2278
rect 931 948 983 958
rect 1657 3960 1709 3975
rect 1657 3520 1709 3908
rect 1657 3080 1709 3468
rect 1657 2640 1709 3028
rect 1657 2200 1709 2588
rect 1657 1760 1709 2148
rect 1657 1320 1709 1708
rect 2401 3650 2453 4445
rect 3871 4901 3923 6169
rect 4711 5025 4763 6293
rect 6186 6412 6322 9416
rect 6741 7581 6793 7591
rect 7072 7581 7124 7591
rect 6793 7529 7072 7581
rect 6741 7519 6793 7529
rect 7070 7519 7124 7529
rect 6482 6720 6534 6730
rect 6833 6720 6885 6730
rect 6462 6668 6482 6720
rect 6534 6668 6833 6720
rect 6885 6668 6889 6720
rect 6482 6658 6534 6668
rect 6833 6658 6885 6668
rect 6186 6360 6229 6412
rect 6281 6360 6322 6412
rect 6741 6431 6793 6441
rect 7070 6431 7122 7519
rect 6793 6379 7070 6431
rect 6741 6369 6793 6379
rect 6186 6271 6322 6360
rect 4711 4963 4763 4973
rect 5340 6221 5392 6237
rect 3871 4497 3923 4849
rect 2401 3210 2453 3598
rect 2401 1890 2453 3158
rect 2401 1450 2453 1838
rect 2401 1388 2453 1398
rect 2917 3960 2969 3974
rect 2917 3520 2969 3908
rect 2917 3080 2969 3468
rect 2917 2640 2969 3028
rect 2917 2200 2969 2588
rect 2917 1760 2969 2148
rect 302 567 354 828
rect 302 211 354 463
rect 1657 880 1709 1268
rect 1657 567 1709 828
rect 1036 313 1100 323
rect 1036 239 1100 249
rect 302 149 354 159
rect 1657 211 1709 463
rect 2917 1320 2969 1708
rect 3871 3650 3923 4445
rect 5340 4901 5392 6169
rect 5340 4497 5392 4849
rect 3871 3210 3923 3598
rect 3871 1890 3923 3158
rect 3871 1450 3923 1838
rect 3871 1388 3923 1398
rect 4921 3960 4973 3970
rect 4921 3520 4973 3908
rect 4921 3080 4973 3468
rect 4921 2640 4973 3028
rect 4921 2200 4973 2588
rect 4921 1760 4973 2148
rect 2917 880 2969 1268
rect 2917 567 2969 828
rect 2380 313 2444 323
rect 2380 239 2444 249
rect 1657 149 1709 159
rect 2917 211 2969 463
rect 4921 1320 4973 1708
rect 5340 3650 5392 4445
rect 6186 6219 6229 6271
rect 6281 6219 6322 6271
rect 6186 6130 6322 6219
rect 6186 6078 6229 6130
rect 6281 6078 6322 6130
rect 6186 5989 6322 6078
rect 6186 5937 6229 5989
rect 6281 5937 6322 5989
rect 6186 5848 6322 5937
rect 7070 5871 7122 6379
rect 6186 5796 6229 5848
rect 6281 5796 6322 5848
rect 6186 5707 6322 5796
rect 7064 5861 7128 5871
rect 7064 5787 7128 5797
rect 6186 5655 6229 5707
rect 6281 5655 6322 5707
rect 6186 5566 6322 5655
rect 6186 5514 6229 5566
rect 6281 5514 6322 5566
rect 6186 5425 6322 5514
rect 6186 5373 6229 5425
rect 6281 5373 6322 5425
rect 6186 5284 6322 5373
rect 6186 5232 6229 5284
rect 6281 5232 6322 5284
rect 6186 5143 6322 5232
rect 6186 5091 6229 5143
rect 6281 5091 6322 5143
rect 6739 5173 6791 5183
rect 7070 5173 7122 5787
rect 6791 5121 7070 5173
rect 6739 5111 6791 5121
rect 6186 5002 6322 5091
rect 6186 4950 6229 5002
rect 6281 4950 6322 5002
rect 6186 4861 6322 4950
rect 6186 4809 6229 4861
rect 6281 4809 6322 4861
rect 6186 4144 6322 4809
rect 6482 4497 6534 4507
rect 6835 4497 6887 4507
rect 6462 4445 6482 4497
rect 6534 4445 6835 4497
rect 6887 4445 6889 4497
rect 6482 4435 6534 4445
rect 6835 4435 6887 4445
rect 6186 4092 6229 4144
rect 6281 4092 6322 4144
rect 6186 4003 6322 4092
rect 6186 3951 6229 4003
rect 6281 3951 6322 4003
rect 6741 4021 6793 4031
rect 7070 4021 7122 5121
rect 6793 3969 7070 4021
rect 6741 3959 6793 3969
rect 7070 3959 7122 3969
rect 6186 3862 6322 3951
rect 6186 3810 6229 3862
rect 6281 3810 6322 3862
rect 5340 3210 5392 3598
rect 5340 1890 5392 3158
rect 5340 1450 5392 1838
rect 5340 1388 5392 1398
rect 6020 3743 6072 3753
rect 6020 3433 6072 3691
rect 6020 3305 6072 3381
rect 6020 2991 6072 3253
rect 6020 1985 6072 2939
rect 6186 3721 6322 3810
rect 6186 3669 6229 3721
rect 6281 3669 6322 3721
rect 6186 3580 6322 3669
rect 6186 3528 6229 3580
rect 6281 3528 6322 3580
rect 6186 3439 6322 3528
rect 6186 3387 6229 3439
rect 6281 3387 6322 3439
rect 6186 3298 6322 3387
rect 6186 3246 6229 3298
rect 6281 3246 6322 3298
rect 6186 3157 6322 3246
rect 6186 3105 6229 3157
rect 6281 3105 6322 3157
rect 6186 3016 6322 3105
rect 6186 2964 6229 3016
rect 6281 2964 6322 3016
rect 6186 2875 6322 2964
rect 6186 2823 6229 2875
rect 6281 2823 6322 2875
rect 6186 2734 6322 2823
rect 6186 2682 6229 2734
rect 6281 2682 6322 2734
rect 6186 2672 6322 2682
rect 6020 1671 6072 1933
rect 6020 1544 6072 1619
rect 4921 880 4973 1268
rect 6020 1233 6072 1492
rect 6020 1168 6072 1181
rect 6186 1549 6322 1559
rect 6186 1497 6229 1549
rect 6281 1497 6322 1549
rect 6186 1408 6322 1497
rect 6186 1356 6229 1408
rect 6281 1356 6322 1408
rect 6186 1267 6322 1356
rect 6186 1215 6229 1267
rect 6281 1215 6322 1267
rect 4921 567 4973 828
rect 4921 453 4973 463
rect 6186 1126 6322 1215
rect 6186 1074 6229 1126
rect 6281 1074 6322 1126
rect 6186 985 6322 1074
rect 6186 933 6229 985
rect 6281 933 6322 985
rect 6186 844 6322 933
rect 6186 792 6229 844
rect 6281 792 6322 844
rect 2917 149 2969 159
rect -2845 -115 -2004 -52
rect 6186 -57 6322 792
rect -2845 -167 -2798 -115
rect -2746 -167 -2657 -115
rect -2605 -167 -2516 -115
rect -2464 -167 -2375 -115
rect -2323 -167 -2234 -115
rect -2182 -167 -2093 -115
rect -2041 -167 -2004 -115
rect -2845 -193 -2004 -167
rect 5496 -114 6322 -57
rect 5496 -166 5523 -114
rect 5575 -166 5664 -114
rect 5716 -166 5805 -114
rect 5857 -166 5946 -114
rect 5998 -166 6087 -114
rect 6139 -166 6228 -114
rect 6280 -166 6322 -114
rect 5496 -193 6322 -166
<< via2 >>
rect -3667 5797 -3603 5861
rect 1036 303 1100 313
rect 1036 251 1042 303
rect 1042 251 1094 303
rect 1094 251 1100 303
rect 1036 249 1100 251
rect 2380 303 2444 313
rect 2380 251 2385 303
rect 2385 251 2437 303
rect 2437 251 2444 303
rect 2380 249 2444 251
rect 7064 5797 7128 5861
<< metal3 >>
rect -3677 5861 -3593 5866
rect 7054 5861 7138 5866
rect -3677 5797 -3667 5861
rect -3603 5797 7064 5861
rect 7128 5797 7138 5861
rect -3677 5792 -3593 5797
rect 1698 492 1762 5797
rect 7054 5792 7138 5797
rect 1036 428 2444 492
rect 1036 318 1100 428
rect 2380 318 2444 428
rect 1026 313 1110 318
rect 1026 249 1036 313
rect 1100 249 1110 313
rect 1026 244 1110 249
rect 2370 313 2454 318
rect 2370 249 2380 313
rect 2444 249 2454 313
rect 2370 244 2454 249
rect 2380 242 2444 244
<< labels >>
flabel metal1 1334 10724 1334 10724 5 FreeSans 400 0 0 0 outn
port 5 s
flabel metal1 2119 10721 2119 10721 1 FreeSans 400 0 0 0 outp
port 4 n
flabel metal3 1730 4459 1730 4459 1 FreeSans 400 0 0 0 clk
port 1 n
flabel metal1 -3776 8059 -3776 8059 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 -3228 -136 -3228 -136 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
flabel metal2 6063 2476 6063 2476 1 FreeSans 400 0 0 0 in
port 3 n
flabel metal2 -2580 2466 -2580 2466 1 FreeSans 400 0 0 0 ip
port 2 n
flabel metal1 1709 8270 1743 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VPWR
flabel metal1 2253 8270 2287 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VGND
flabel locali 1709 8270 1743 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VPWR
flabel locali 2253 8270 2287 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VGND
flabel locali 2151 8453 2185 8487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/X
flabel locali 1879 8453 1913 8487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/X
flabel locali 1811 8453 1845 8487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/X
flabel locali 2015 8270 2049 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/A
flabel nwell 1709 8270 1743 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VPB
flabel pwell 2253 8270 2287 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_0/VNB
rlabel comment 2270 8241 2270 8241 2 sky130_fd_sc_hd__buf_2_0/buf_2
rlabel metal1 2222 8241 2318 8609 7 sky130_fd_sc_hd__buf_2_0/VGND
rlabel metal1 1678 8241 1774 8609 7 sky130_fd_sc_hd__buf_2_0/VPWR
flabel metal1 1709 8270 1743 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VPWR
flabel metal1 1165 8270 1199 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VGND
flabel locali 1709 8270 1743 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VPWR
flabel locali 1165 8270 1199 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VGND
flabel locali 1267 8453 1301 8487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/X
flabel locali 1539 8453 1573 8487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/X
flabel locali 1607 8453 1641 8487 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/X
flabel locali 1403 8270 1437 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/A
flabel nwell 1709 8270 1743 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VPB
flabel pwell 1165 8270 1199 8304 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__buf_2_1/VNB
rlabel comment 1182 8241 1182 8241 8 sky130_fd_sc_hd__buf_2_1/buf_2
rlabel metal1 1134 8241 1230 8609 3 sky130_fd_sc_hd__buf_2_1/VGND
rlabel metal1 1678 8241 1774 8609 3 sky130_fd_sc_hd__buf_2_1/VPWR
flabel metal1 1165 10570 1199 10604 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VGND
flabel metal1 1709 10570 1743 10604 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VPWR
flabel nwell 1709 10570 1743 10604 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VPB
flabel pwell 1165 10570 1199 10604 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_0/VNB
rlabel comment 1182 10633 1182 10633 6 sky130_fd_sc_hd__decap_12_0/decap_12
rlabel metal1 1134 9529 1230 10633 3 sky130_fd_sc_hd__decap_12_0/VGND
rlabel metal1 1678 9529 1774 10633 3 sky130_fd_sc_hd__decap_12_0/VPWR
flabel metal1 2253 9558 2287 9592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VGND
flabel metal1 1709 9558 1743 9592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VPWR
flabel nwell 1709 9558 1743 9592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VPB
flabel pwell 2253 9558 2287 9592 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__decap_12_1/VNB
rlabel comment 2270 9529 2270 9529 2 sky130_fd_sc_hd__decap_12_1/decap_12
rlabel metal1 2222 9529 2318 10633 7 sky130_fd_sc_hd__decap_12_1/VGND
rlabel metal1 1678 9529 1774 10633 7 sky130_fd_sc_hd__decap_12_1/VPWR
flabel locali 1403 9005 1437 9039 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/Y
flabel locali 1471 9005 1505 9039 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/Y
flabel locali 1403 8729 1437 8763 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/A
flabel locali 1403 8821 1437 8855 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/A
flabel locali 1403 9097 1437 9131 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 1403 9189 1437 9223 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 1403 9373 1437 9407 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel locali 1403 9281 1437 9315 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_0/B
flabel nwell 1709 9373 1743 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VPB
flabel pwell 1165 9373 1199 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VNB
flabel metal1 1165 9373 1199 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VGND
flabel metal1 1709 9373 1743 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_0/VPWR
rlabel comment 1182 9437 1182 9437 6 sky130_fd_sc_hd__nand2_4_0/nand2_4
rlabel metal1 1134 8609 1230 9437 3 sky130_fd_sc_hd__nand2_4_0/VGND
rlabel metal1 1678 8609 1774 9437 3 sky130_fd_sc_hd__nand2_4_0/VPWR
flabel locali 2015 9005 2049 9039 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/Y
flabel locali 1947 9005 1981 9039 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/Y
flabel locali 2015 8729 2049 8763 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/A
flabel locali 2015 8821 2049 8855 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/A
flabel locali 2015 9097 2049 9131 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 2015 9189 2049 9223 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 2015 9373 2049 9407 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel locali 2015 9281 2049 9315 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_4_1/B
flabel nwell 1709 9373 1743 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VPB
flabel pwell 2253 9373 2287 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VNB
flabel metal1 2253 9373 2287 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VGND
flabel metal1 1709 9373 1743 9407 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_4_1/VPWR
rlabel comment 2270 9437 2270 9437 4 sky130_fd_sc_hd__nand2_4_1/nand2_4
rlabel metal1 2222 8609 2318 9437 7 sky130_fd_sc_hd__nand2_4_1/VGND
rlabel metal1 1678 8609 1774 9437 7 sky130_fd_sc_hd__nand2_4_1/VPWR
flabel metal1 1706 9454 1735 9507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 1164 9457 1202 9508 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment 1182 9529 1182 9529 6 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
rlabel metal1 1134 9437 1230 9529 3 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel metal1 1678 9437 1774 9529 3 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 1717 9459 1746 9512 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 2250 9458 2288 9509 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment 2270 9437 2270 9437 2 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
rlabel metal1 2222 9437 2318 9529 7 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel metal1 1678 9437 1774 9529 7 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
<< end >>
