magic
tech sky130A
magscale 1 2
timestamp 1653460579
<< nwell >>
rect -2098 7664 -804 8314
rect 6902 7664 8196 8314
rect -2098 5864 -804 6514
rect 6902 5864 8196 6514
rect -2098 4064 -804 4714
rect 6902 4064 8196 4714
rect -2098 2264 -804 2914
rect 6902 2264 8196 2914
rect -2098 464 -804 1114
rect 6902 464 8196 1114
rect -2098 -1336 -804 -686
rect 6902 -1336 8196 -686
<< pwell >>
rect -2098 7200 -804 7664
rect 6902 7200 8196 7664
rect -2098 5400 -804 5864
rect 6902 5400 8196 5864
rect -2098 3600 -804 4064
rect 6902 3600 8196 4064
rect -2098 1800 -804 2264
rect 6902 1800 8196 2264
rect -2098 0 -804 464
rect 6902 0 8196 464
rect -2098 -1800 -804 -1336
rect 6902 -1800 8196 -1336
<< nmos >>
rect -1898 7410 -1868 7516
rect -1802 7410 -1772 7516
rect -1706 7410 -1676 7516
rect -1610 7410 -1580 7516
rect -1514 7410 -1484 7516
rect -1418 7410 -1388 7516
rect -1322 7410 -1292 7516
rect -1226 7410 -1196 7516
rect -1130 7410 -1100 7516
rect -1034 7410 -1004 7516
rect 7102 7410 7132 7516
rect 7198 7410 7228 7516
rect 7294 7410 7324 7516
rect 7390 7410 7420 7516
rect 7486 7410 7516 7516
rect 7582 7410 7612 7516
rect 7678 7410 7708 7516
rect 7774 7410 7804 7516
rect 7870 7410 7900 7516
rect 7966 7410 7996 7516
rect -1898 5610 -1868 5716
rect -1802 5610 -1772 5716
rect -1706 5610 -1676 5716
rect -1610 5610 -1580 5716
rect -1514 5610 -1484 5716
rect -1418 5610 -1388 5716
rect -1322 5610 -1292 5716
rect -1226 5610 -1196 5716
rect -1130 5610 -1100 5716
rect -1034 5610 -1004 5716
rect 7102 5610 7132 5716
rect 7198 5610 7228 5716
rect 7294 5610 7324 5716
rect 7390 5610 7420 5716
rect 7486 5610 7516 5716
rect 7582 5610 7612 5716
rect 7678 5610 7708 5716
rect 7774 5610 7804 5716
rect 7870 5610 7900 5716
rect 7966 5610 7996 5716
rect -1898 3810 -1868 3916
rect -1802 3810 -1772 3916
rect -1706 3810 -1676 3916
rect -1610 3810 -1580 3916
rect -1514 3810 -1484 3916
rect -1418 3810 -1388 3916
rect -1322 3810 -1292 3916
rect -1226 3810 -1196 3916
rect -1130 3810 -1100 3916
rect -1034 3810 -1004 3916
rect 7102 3810 7132 3916
rect 7198 3810 7228 3916
rect 7294 3810 7324 3916
rect 7390 3810 7420 3916
rect 7486 3810 7516 3916
rect 7582 3810 7612 3916
rect 7678 3810 7708 3916
rect 7774 3810 7804 3916
rect 7870 3810 7900 3916
rect 7966 3810 7996 3916
rect -1898 2010 -1868 2116
rect -1802 2010 -1772 2116
rect -1706 2010 -1676 2116
rect -1610 2010 -1580 2116
rect -1514 2010 -1484 2116
rect -1418 2010 -1388 2116
rect -1322 2010 -1292 2116
rect -1226 2010 -1196 2116
rect -1130 2010 -1100 2116
rect -1034 2010 -1004 2116
rect 7102 2010 7132 2116
rect 7198 2010 7228 2116
rect 7294 2010 7324 2116
rect 7390 2010 7420 2116
rect 7486 2010 7516 2116
rect 7582 2010 7612 2116
rect 7678 2010 7708 2116
rect 7774 2010 7804 2116
rect 7870 2010 7900 2116
rect 7966 2010 7996 2116
rect -1898 210 -1868 316
rect -1802 210 -1772 316
rect -1706 210 -1676 316
rect -1610 210 -1580 316
rect -1514 210 -1484 316
rect -1418 210 -1388 316
rect -1322 210 -1292 316
rect -1226 210 -1196 316
rect -1130 210 -1100 316
rect -1034 210 -1004 316
rect 7102 210 7132 316
rect 7198 210 7228 316
rect 7294 210 7324 316
rect 7390 210 7420 316
rect 7486 210 7516 316
rect 7582 210 7612 316
rect 7678 210 7708 316
rect 7774 210 7804 316
rect 7870 210 7900 316
rect 7966 210 7996 316
rect -1898 -1590 -1868 -1484
rect -1802 -1590 -1772 -1484
rect -1706 -1590 -1676 -1484
rect -1610 -1590 -1580 -1484
rect -1514 -1590 -1484 -1484
rect -1418 -1590 -1388 -1484
rect -1322 -1590 -1292 -1484
rect -1226 -1590 -1196 -1484
rect -1130 -1590 -1100 -1484
rect -1034 -1590 -1004 -1484
rect 7102 -1590 7132 -1484
rect 7198 -1590 7228 -1484
rect 7294 -1590 7324 -1484
rect 7390 -1590 7420 -1484
rect 7486 -1590 7516 -1484
rect 7582 -1590 7612 -1484
rect 7678 -1590 7708 -1484
rect 7774 -1590 7804 -1484
rect 7870 -1590 7900 -1484
rect 7966 -1590 7996 -1484
<< pmos >>
rect -1898 7821 -1868 8095
rect -1802 7821 -1772 8095
rect -1706 7821 -1676 8095
rect -1610 7821 -1580 8095
rect -1514 7821 -1484 8095
rect -1418 7821 -1388 8095
rect -1322 7821 -1292 8095
rect -1226 7821 -1196 8095
rect -1130 7821 -1100 8095
rect -1034 7821 -1004 8095
rect 7102 7821 7132 8095
rect 7198 7821 7228 8095
rect 7294 7821 7324 8095
rect 7390 7821 7420 8095
rect 7486 7821 7516 8095
rect 7582 7821 7612 8095
rect 7678 7821 7708 8095
rect 7774 7821 7804 8095
rect 7870 7821 7900 8095
rect 7966 7821 7996 8095
rect -1898 6021 -1868 6295
rect -1802 6021 -1772 6295
rect -1706 6021 -1676 6295
rect -1610 6021 -1580 6295
rect -1514 6021 -1484 6295
rect -1418 6021 -1388 6295
rect -1322 6021 -1292 6295
rect -1226 6021 -1196 6295
rect -1130 6021 -1100 6295
rect -1034 6021 -1004 6295
rect 7102 6021 7132 6295
rect 7198 6021 7228 6295
rect 7294 6021 7324 6295
rect 7390 6021 7420 6295
rect 7486 6021 7516 6295
rect 7582 6021 7612 6295
rect 7678 6021 7708 6295
rect 7774 6021 7804 6295
rect 7870 6021 7900 6295
rect 7966 6021 7996 6295
rect -1898 4221 -1868 4495
rect -1802 4221 -1772 4495
rect -1706 4221 -1676 4495
rect -1610 4221 -1580 4495
rect -1514 4221 -1484 4495
rect -1418 4221 -1388 4495
rect -1322 4221 -1292 4495
rect -1226 4221 -1196 4495
rect -1130 4221 -1100 4495
rect -1034 4221 -1004 4495
rect 7102 4221 7132 4495
rect 7198 4221 7228 4495
rect 7294 4221 7324 4495
rect 7390 4221 7420 4495
rect 7486 4221 7516 4495
rect 7582 4221 7612 4495
rect 7678 4221 7708 4495
rect 7774 4221 7804 4495
rect 7870 4221 7900 4495
rect 7966 4221 7996 4495
rect -1898 2421 -1868 2695
rect -1802 2421 -1772 2695
rect -1706 2421 -1676 2695
rect -1610 2421 -1580 2695
rect -1514 2421 -1484 2695
rect -1418 2421 -1388 2695
rect -1322 2421 -1292 2695
rect -1226 2421 -1196 2695
rect -1130 2421 -1100 2695
rect -1034 2421 -1004 2695
rect 7102 2421 7132 2695
rect 7198 2421 7228 2695
rect 7294 2421 7324 2695
rect 7390 2421 7420 2695
rect 7486 2421 7516 2695
rect 7582 2421 7612 2695
rect 7678 2421 7708 2695
rect 7774 2421 7804 2695
rect 7870 2421 7900 2695
rect 7966 2421 7996 2695
rect -1898 621 -1868 895
rect -1802 621 -1772 895
rect -1706 621 -1676 895
rect -1610 621 -1580 895
rect -1514 621 -1484 895
rect -1418 621 -1388 895
rect -1322 621 -1292 895
rect -1226 621 -1196 895
rect -1130 621 -1100 895
rect -1034 621 -1004 895
rect 7102 621 7132 895
rect 7198 621 7228 895
rect 7294 621 7324 895
rect 7390 621 7420 895
rect 7486 621 7516 895
rect 7582 621 7612 895
rect 7678 621 7708 895
rect 7774 621 7804 895
rect 7870 621 7900 895
rect 7966 621 7996 895
rect -1898 -1179 -1868 -905
rect -1802 -1179 -1772 -905
rect -1706 -1179 -1676 -905
rect -1610 -1179 -1580 -905
rect -1514 -1179 -1484 -905
rect -1418 -1179 -1388 -905
rect -1322 -1179 -1292 -905
rect -1226 -1179 -1196 -905
rect -1130 -1179 -1100 -905
rect -1034 -1179 -1004 -905
rect 7102 -1179 7132 -905
rect 7198 -1179 7228 -905
rect 7294 -1179 7324 -905
rect 7390 -1179 7420 -905
rect 7486 -1179 7516 -905
rect 7582 -1179 7612 -905
rect 7678 -1179 7708 -905
rect 7774 -1179 7804 -905
rect 7870 -1179 7900 -905
rect 7966 -1179 7996 -905
<< ndiff >>
rect -1960 7504 -1898 7516
rect -1960 7422 -1948 7504
rect -1914 7422 -1898 7504
rect -1960 7410 -1898 7422
rect -1868 7504 -1802 7516
rect -1868 7422 -1852 7504
rect -1818 7422 -1802 7504
rect -1868 7410 -1802 7422
rect -1772 7504 -1706 7516
rect -1772 7422 -1756 7504
rect -1722 7422 -1706 7504
rect -1772 7410 -1706 7422
rect -1676 7504 -1610 7516
rect -1676 7422 -1660 7504
rect -1626 7422 -1610 7504
rect -1676 7410 -1610 7422
rect -1580 7504 -1514 7516
rect -1580 7422 -1564 7504
rect -1530 7422 -1514 7504
rect -1580 7410 -1514 7422
rect -1484 7504 -1418 7516
rect -1484 7422 -1468 7504
rect -1434 7422 -1418 7504
rect -1484 7410 -1418 7422
rect -1388 7504 -1322 7516
rect -1388 7422 -1372 7504
rect -1338 7422 -1322 7504
rect -1388 7410 -1322 7422
rect -1292 7504 -1226 7516
rect -1292 7422 -1276 7504
rect -1242 7422 -1226 7504
rect -1292 7410 -1226 7422
rect -1196 7504 -1130 7516
rect -1196 7422 -1180 7504
rect -1146 7422 -1130 7504
rect -1196 7410 -1130 7422
rect -1100 7504 -1034 7516
rect -1100 7422 -1084 7504
rect -1050 7422 -1034 7504
rect -1100 7410 -1034 7422
rect -1004 7504 -942 7516
rect -1004 7422 -988 7504
rect -954 7422 -942 7504
rect -1004 7410 -942 7422
rect 7040 7504 7102 7516
rect 7040 7422 7052 7504
rect 7086 7422 7102 7504
rect 7040 7410 7102 7422
rect 7132 7504 7198 7516
rect 7132 7422 7148 7504
rect 7182 7422 7198 7504
rect 7132 7410 7198 7422
rect 7228 7504 7294 7516
rect 7228 7422 7244 7504
rect 7278 7422 7294 7504
rect 7228 7410 7294 7422
rect 7324 7504 7390 7516
rect 7324 7422 7340 7504
rect 7374 7422 7390 7504
rect 7324 7410 7390 7422
rect 7420 7504 7486 7516
rect 7420 7422 7436 7504
rect 7470 7422 7486 7504
rect 7420 7410 7486 7422
rect 7516 7504 7582 7516
rect 7516 7422 7532 7504
rect 7566 7422 7582 7504
rect 7516 7410 7582 7422
rect 7612 7504 7678 7516
rect 7612 7422 7628 7504
rect 7662 7422 7678 7504
rect 7612 7410 7678 7422
rect 7708 7504 7774 7516
rect 7708 7422 7724 7504
rect 7758 7422 7774 7504
rect 7708 7410 7774 7422
rect 7804 7504 7870 7516
rect 7804 7422 7820 7504
rect 7854 7422 7870 7504
rect 7804 7410 7870 7422
rect 7900 7504 7966 7516
rect 7900 7422 7916 7504
rect 7950 7422 7966 7504
rect 7900 7410 7966 7422
rect 7996 7504 8058 7516
rect 7996 7422 8012 7504
rect 8046 7422 8058 7504
rect 7996 7410 8058 7422
rect -1960 5704 -1898 5716
rect -1960 5622 -1948 5704
rect -1914 5622 -1898 5704
rect -1960 5610 -1898 5622
rect -1868 5704 -1802 5716
rect -1868 5622 -1852 5704
rect -1818 5622 -1802 5704
rect -1868 5610 -1802 5622
rect -1772 5704 -1706 5716
rect -1772 5622 -1756 5704
rect -1722 5622 -1706 5704
rect -1772 5610 -1706 5622
rect -1676 5704 -1610 5716
rect -1676 5622 -1660 5704
rect -1626 5622 -1610 5704
rect -1676 5610 -1610 5622
rect -1580 5704 -1514 5716
rect -1580 5622 -1564 5704
rect -1530 5622 -1514 5704
rect -1580 5610 -1514 5622
rect -1484 5704 -1418 5716
rect -1484 5622 -1468 5704
rect -1434 5622 -1418 5704
rect -1484 5610 -1418 5622
rect -1388 5704 -1322 5716
rect -1388 5622 -1372 5704
rect -1338 5622 -1322 5704
rect -1388 5610 -1322 5622
rect -1292 5704 -1226 5716
rect -1292 5622 -1276 5704
rect -1242 5622 -1226 5704
rect -1292 5610 -1226 5622
rect -1196 5704 -1130 5716
rect -1196 5622 -1180 5704
rect -1146 5622 -1130 5704
rect -1196 5610 -1130 5622
rect -1100 5704 -1034 5716
rect -1100 5622 -1084 5704
rect -1050 5622 -1034 5704
rect -1100 5610 -1034 5622
rect -1004 5704 -942 5716
rect -1004 5622 -988 5704
rect -954 5622 -942 5704
rect -1004 5610 -942 5622
rect 7040 5704 7102 5716
rect 7040 5622 7052 5704
rect 7086 5622 7102 5704
rect 7040 5610 7102 5622
rect 7132 5704 7198 5716
rect 7132 5622 7148 5704
rect 7182 5622 7198 5704
rect 7132 5610 7198 5622
rect 7228 5704 7294 5716
rect 7228 5622 7244 5704
rect 7278 5622 7294 5704
rect 7228 5610 7294 5622
rect 7324 5704 7390 5716
rect 7324 5622 7340 5704
rect 7374 5622 7390 5704
rect 7324 5610 7390 5622
rect 7420 5704 7486 5716
rect 7420 5622 7436 5704
rect 7470 5622 7486 5704
rect 7420 5610 7486 5622
rect 7516 5704 7582 5716
rect 7516 5622 7532 5704
rect 7566 5622 7582 5704
rect 7516 5610 7582 5622
rect 7612 5704 7678 5716
rect 7612 5622 7628 5704
rect 7662 5622 7678 5704
rect 7612 5610 7678 5622
rect 7708 5704 7774 5716
rect 7708 5622 7724 5704
rect 7758 5622 7774 5704
rect 7708 5610 7774 5622
rect 7804 5704 7870 5716
rect 7804 5622 7820 5704
rect 7854 5622 7870 5704
rect 7804 5610 7870 5622
rect 7900 5704 7966 5716
rect 7900 5622 7916 5704
rect 7950 5622 7966 5704
rect 7900 5610 7966 5622
rect 7996 5704 8058 5716
rect 7996 5622 8012 5704
rect 8046 5622 8058 5704
rect 7996 5610 8058 5622
rect -1960 3904 -1898 3916
rect -1960 3822 -1948 3904
rect -1914 3822 -1898 3904
rect -1960 3810 -1898 3822
rect -1868 3904 -1802 3916
rect -1868 3822 -1852 3904
rect -1818 3822 -1802 3904
rect -1868 3810 -1802 3822
rect -1772 3904 -1706 3916
rect -1772 3822 -1756 3904
rect -1722 3822 -1706 3904
rect -1772 3810 -1706 3822
rect -1676 3904 -1610 3916
rect -1676 3822 -1660 3904
rect -1626 3822 -1610 3904
rect -1676 3810 -1610 3822
rect -1580 3904 -1514 3916
rect -1580 3822 -1564 3904
rect -1530 3822 -1514 3904
rect -1580 3810 -1514 3822
rect -1484 3904 -1418 3916
rect -1484 3822 -1468 3904
rect -1434 3822 -1418 3904
rect -1484 3810 -1418 3822
rect -1388 3904 -1322 3916
rect -1388 3822 -1372 3904
rect -1338 3822 -1322 3904
rect -1388 3810 -1322 3822
rect -1292 3904 -1226 3916
rect -1292 3822 -1276 3904
rect -1242 3822 -1226 3904
rect -1292 3810 -1226 3822
rect -1196 3904 -1130 3916
rect -1196 3822 -1180 3904
rect -1146 3822 -1130 3904
rect -1196 3810 -1130 3822
rect -1100 3904 -1034 3916
rect -1100 3822 -1084 3904
rect -1050 3822 -1034 3904
rect -1100 3810 -1034 3822
rect -1004 3904 -942 3916
rect -1004 3822 -988 3904
rect -954 3822 -942 3904
rect -1004 3810 -942 3822
rect 7040 3904 7102 3916
rect 7040 3822 7052 3904
rect 7086 3822 7102 3904
rect 7040 3810 7102 3822
rect 7132 3904 7198 3916
rect 7132 3822 7148 3904
rect 7182 3822 7198 3904
rect 7132 3810 7198 3822
rect 7228 3904 7294 3916
rect 7228 3822 7244 3904
rect 7278 3822 7294 3904
rect 7228 3810 7294 3822
rect 7324 3904 7390 3916
rect 7324 3822 7340 3904
rect 7374 3822 7390 3904
rect 7324 3810 7390 3822
rect 7420 3904 7486 3916
rect 7420 3822 7436 3904
rect 7470 3822 7486 3904
rect 7420 3810 7486 3822
rect 7516 3904 7582 3916
rect 7516 3822 7532 3904
rect 7566 3822 7582 3904
rect 7516 3810 7582 3822
rect 7612 3904 7678 3916
rect 7612 3822 7628 3904
rect 7662 3822 7678 3904
rect 7612 3810 7678 3822
rect 7708 3904 7774 3916
rect 7708 3822 7724 3904
rect 7758 3822 7774 3904
rect 7708 3810 7774 3822
rect 7804 3904 7870 3916
rect 7804 3822 7820 3904
rect 7854 3822 7870 3904
rect 7804 3810 7870 3822
rect 7900 3904 7966 3916
rect 7900 3822 7916 3904
rect 7950 3822 7966 3904
rect 7900 3810 7966 3822
rect 7996 3904 8058 3916
rect 7996 3822 8012 3904
rect 8046 3822 8058 3904
rect 7996 3810 8058 3822
rect -1960 2104 -1898 2116
rect -1960 2022 -1948 2104
rect -1914 2022 -1898 2104
rect -1960 2010 -1898 2022
rect -1868 2104 -1802 2116
rect -1868 2022 -1852 2104
rect -1818 2022 -1802 2104
rect -1868 2010 -1802 2022
rect -1772 2104 -1706 2116
rect -1772 2022 -1756 2104
rect -1722 2022 -1706 2104
rect -1772 2010 -1706 2022
rect -1676 2104 -1610 2116
rect -1676 2022 -1660 2104
rect -1626 2022 -1610 2104
rect -1676 2010 -1610 2022
rect -1580 2104 -1514 2116
rect -1580 2022 -1564 2104
rect -1530 2022 -1514 2104
rect -1580 2010 -1514 2022
rect -1484 2104 -1418 2116
rect -1484 2022 -1468 2104
rect -1434 2022 -1418 2104
rect -1484 2010 -1418 2022
rect -1388 2104 -1322 2116
rect -1388 2022 -1372 2104
rect -1338 2022 -1322 2104
rect -1388 2010 -1322 2022
rect -1292 2104 -1226 2116
rect -1292 2022 -1276 2104
rect -1242 2022 -1226 2104
rect -1292 2010 -1226 2022
rect -1196 2104 -1130 2116
rect -1196 2022 -1180 2104
rect -1146 2022 -1130 2104
rect -1196 2010 -1130 2022
rect -1100 2104 -1034 2116
rect -1100 2022 -1084 2104
rect -1050 2022 -1034 2104
rect -1100 2010 -1034 2022
rect -1004 2104 -942 2116
rect -1004 2022 -988 2104
rect -954 2022 -942 2104
rect -1004 2010 -942 2022
rect 7040 2104 7102 2116
rect 7040 2022 7052 2104
rect 7086 2022 7102 2104
rect 7040 2010 7102 2022
rect 7132 2104 7198 2116
rect 7132 2022 7148 2104
rect 7182 2022 7198 2104
rect 7132 2010 7198 2022
rect 7228 2104 7294 2116
rect 7228 2022 7244 2104
rect 7278 2022 7294 2104
rect 7228 2010 7294 2022
rect 7324 2104 7390 2116
rect 7324 2022 7340 2104
rect 7374 2022 7390 2104
rect 7324 2010 7390 2022
rect 7420 2104 7486 2116
rect 7420 2022 7436 2104
rect 7470 2022 7486 2104
rect 7420 2010 7486 2022
rect 7516 2104 7582 2116
rect 7516 2022 7532 2104
rect 7566 2022 7582 2104
rect 7516 2010 7582 2022
rect 7612 2104 7678 2116
rect 7612 2022 7628 2104
rect 7662 2022 7678 2104
rect 7612 2010 7678 2022
rect 7708 2104 7774 2116
rect 7708 2022 7724 2104
rect 7758 2022 7774 2104
rect 7708 2010 7774 2022
rect 7804 2104 7870 2116
rect 7804 2022 7820 2104
rect 7854 2022 7870 2104
rect 7804 2010 7870 2022
rect 7900 2104 7966 2116
rect 7900 2022 7916 2104
rect 7950 2022 7966 2104
rect 7900 2010 7966 2022
rect 7996 2104 8058 2116
rect 7996 2022 8012 2104
rect 8046 2022 8058 2104
rect 7996 2010 8058 2022
rect -1960 304 -1898 316
rect -1960 222 -1948 304
rect -1914 222 -1898 304
rect -1960 210 -1898 222
rect -1868 304 -1802 316
rect -1868 222 -1852 304
rect -1818 222 -1802 304
rect -1868 210 -1802 222
rect -1772 304 -1706 316
rect -1772 222 -1756 304
rect -1722 222 -1706 304
rect -1772 210 -1706 222
rect -1676 304 -1610 316
rect -1676 222 -1660 304
rect -1626 222 -1610 304
rect -1676 210 -1610 222
rect -1580 304 -1514 316
rect -1580 222 -1564 304
rect -1530 222 -1514 304
rect -1580 210 -1514 222
rect -1484 304 -1418 316
rect -1484 222 -1468 304
rect -1434 222 -1418 304
rect -1484 210 -1418 222
rect -1388 304 -1322 316
rect -1388 222 -1372 304
rect -1338 222 -1322 304
rect -1388 210 -1322 222
rect -1292 304 -1226 316
rect -1292 222 -1276 304
rect -1242 222 -1226 304
rect -1292 210 -1226 222
rect -1196 304 -1130 316
rect -1196 222 -1180 304
rect -1146 222 -1130 304
rect -1196 210 -1130 222
rect -1100 304 -1034 316
rect -1100 222 -1084 304
rect -1050 222 -1034 304
rect -1100 210 -1034 222
rect -1004 304 -942 316
rect -1004 222 -988 304
rect -954 222 -942 304
rect -1004 210 -942 222
rect 7040 304 7102 316
rect 7040 222 7052 304
rect 7086 222 7102 304
rect 7040 210 7102 222
rect 7132 304 7198 316
rect 7132 222 7148 304
rect 7182 222 7198 304
rect 7132 210 7198 222
rect 7228 304 7294 316
rect 7228 222 7244 304
rect 7278 222 7294 304
rect 7228 210 7294 222
rect 7324 304 7390 316
rect 7324 222 7340 304
rect 7374 222 7390 304
rect 7324 210 7390 222
rect 7420 304 7486 316
rect 7420 222 7436 304
rect 7470 222 7486 304
rect 7420 210 7486 222
rect 7516 304 7582 316
rect 7516 222 7532 304
rect 7566 222 7582 304
rect 7516 210 7582 222
rect 7612 304 7678 316
rect 7612 222 7628 304
rect 7662 222 7678 304
rect 7612 210 7678 222
rect 7708 304 7774 316
rect 7708 222 7724 304
rect 7758 222 7774 304
rect 7708 210 7774 222
rect 7804 304 7870 316
rect 7804 222 7820 304
rect 7854 222 7870 304
rect 7804 210 7870 222
rect 7900 304 7966 316
rect 7900 222 7916 304
rect 7950 222 7966 304
rect 7900 210 7966 222
rect 7996 304 8058 316
rect 7996 222 8012 304
rect 8046 222 8058 304
rect 7996 210 8058 222
rect -1960 -1496 -1898 -1484
rect -1960 -1578 -1948 -1496
rect -1914 -1578 -1898 -1496
rect -1960 -1590 -1898 -1578
rect -1868 -1496 -1802 -1484
rect -1868 -1578 -1852 -1496
rect -1818 -1578 -1802 -1496
rect -1868 -1590 -1802 -1578
rect -1772 -1496 -1706 -1484
rect -1772 -1578 -1756 -1496
rect -1722 -1578 -1706 -1496
rect -1772 -1590 -1706 -1578
rect -1676 -1496 -1610 -1484
rect -1676 -1578 -1660 -1496
rect -1626 -1578 -1610 -1496
rect -1676 -1590 -1610 -1578
rect -1580 -1496 -1514 -1484
rect -1580 -1578 -1564 -1496
rect -1530 -1578 -1514 -1496
rect -1580 -1590 -1514 -1578
rect -1484 -1496 -1418 -1484
rect -1484 -1578 -1468 -1496
rect -1434 -1578 -1418 -1496
rect -1484 -1590 -1418 -1578
rect -1388 -1496 -1322 -1484
rect -1388 -1578 -1372 -1496
rect -1338 -1578 -1322 -1496
rect -1388 -1590 -1322 -1578
rect -1292 -1496 -1226 -1484
rect -1292 -1578 -1276 -1496
rect -1242 -1578 -1226 -1496
rect -1292 -1590 -1226 -1578
rect -1196 -1496 -1130 -1484
rect -1196 -1578 -1180 -1496
rect -1146 -1578 -1130 -1496
rect -1196 -1590 -1130 -1578
rect -1100 -1496 -1034 -1484
rect -1100 -1578 -1084 -1496
rect -1050 -1578 -1034 -1496
rect -1100 -1590 -1034 -1578
rect -1004 -1496 -942 -1484
rect -1004 -1578 -988 -1496
rect -954 -1578 -942 -1496
rect -1004 -1590 -942 -1578
rect 7040 -1496 7102 -1484
rect 7040 -1578 7052 -1496
rect 7086 -1578 7102 -1496
rect 7040 -1590 7102 -1578
rect 7132 -1496 7198 -1484
rect 7132 -1578 7148 -1496
rect 7182 -1578 7198 -1496
rect 7132 -1590 7198 -1578
rect 7228 -1496 7294 -1484
rect 7228 -1578 7244 -1496
rect 7278 -1578 7294 -1496
rect 7228 -1590 7294 -1578
rect 7324 -1496 7390 -1484
rect 7324 -1578 7340 -1496
rect 7374 -1578 7390 -1496
rect 7324 -1590 7390 -1578
rect 7420 -1496 7486 -1484
rect 7420 -1578 7436 -1496
rect 7470 -1578 7486 -1496
rect 7420 -1590 7486 -1578
rect 7516 -1496 7582 -1484
rect 7516 -1578 7532 -1496
rect 7566 -1578 7582 -1496
rect 7516 -1590 7582 -1578
rect 7612 -1496 7678 -1484
rect 7612 -1578 7628 -1496
rect 7662 -1578 7678 -1496
rect 7612 -1590 7678 -1578
rect 7708 -1496 7774 -1484
rect 7708 -1578 7724 -1496
rect 7758 -1578 7774 -1496
rect 7708 -1590 7774 -1578
rect 7804 -1496 7870 -1484
rect 7804 -1578 7820 -1496
rect 7854 -1578 7870 -1496
rect 7804 -1590 7870 -1578
rect 7900 -1496 7966 -1484
rect 7900 -1578 7916 -1496
rect 7950 -1578 7966 -1496
rect 7900 -1590 7966 -1578
rect 7996 -1496 8058 -1484
rect 7996 -1578 8012 -1496
rect 8046 -1578 8058 -1496
rect 7996 -1590 8058 -1578
<< pdiff >>
rect -1960 8083 -1898 8095
rect -1960 7833 -1948 8083
rect -1914 7833 -1898 8083
rect -1960 7821 -1898 7833
rect -1868 8083 -1802 8095
rect -1868 7833 -1852 8083
rect -1818 7833 -1802 8083
rect -1868 7821 -1802 7833
rect -1772 8083 -1706 8095
rect -1772 7833 -1756 8083
rect -1722 7833 -1706 8083
rect -1772 7821 -1706 7833
rect -1676 8083 -1610 8095
rect -1676 7833 -1660 8083
rect -1626 7833 -1610 8083
rect -1676 7821 -1610 7833
rect -1580 8083 -1514 8095
rect -1580 7833 -1564 8083
rect -1530 7833 -1514 8083
rect -1580 7821 -1514 7833
rect -1484 8083 -1418 8095
rect -1484 7833 -1468 8083
rect -1434 7833 -1418 8083
rect -1484 7821 -1418 7833
rect -1388 8083 -1322 8095
rect -1388 7833 -1372 8083
rect -1338 7833 -1322 8083
rect -1388 7821 -1322 7833
rect -1292 8083 -1226 8095
rect -1292 7833 -1276 8083
rect -1242 7833 -1226 8083
rect -1292 7821 -1226 7833
rect -1196 8083 -1130 8095
rect -1196 7833 -1180 8083
rect -1146 7833 -1130 8083
rect -1196 7821 -1130 7833
rect -1100 8083 -1034 8095
rect -1100 7833 -1084 8083
rect -1050 7833 -1034 8083
rect -1100 7821 -1034 7833
rect -1004 8083 -942 8095
rect -1004 7833 -988 8083
rect -954 7833 -942 8083
rect -1004 7821 -942 7833
rect 7040 8083 7102 8095
rect 7040 7833 7052 8083
rect 7086 7833 7102 8083
rect 7040 7821 7102 7833
rect 7132 8083 7198 8095
rect 7132 7833 7148 8083
rect 7182 7833 7198 8083
rect 7132 7821 7198 7833
rect 7228 8083 7294 8095
rect 7228 7833 7244 8083
rect 7278 7833 7294 8083
rect 7228 7821 7294 7833
rect 7324 8083 7390 8095
rect 7324 7833 7340 8083
rect 7374 7833 7390 8083
rect 7324 7821 7390 7833
rect 7420 8083 7486 8095
rect 7420 7833 7436 8083
rect 7470 7833 7486 8083
rect 7420 7821 7486 7833
rect 7516 8083 7582 8095
rect 7516 7833 7532 8083
rect 7566 7833 7582 8083
rect 7516 7821 7582 7833
rect 7612 8083 7678 8095
rect 7612 7833 7628 8083
rect 7662 7833 7678 8083
rect 7612 7821 7678 7833
rect 7708 8083 7774 8095
rect 7708 7833 7724 8083
rect 7758 7833 7774 8083
rect 7708 7821 7774 7833
rect 7804 8083 7870 8095
rect 7804 7833 7820 8083
rect 7854 7833 7870 8083
rect 7804 7821 7870 7833
rect 7900 8083 7966 8095
rect 7900 7833 7916 8083
rect 7950 7833 7966 8083
rect 7900 7821 7966 7833
rect 7996 8083 8058 8095
rect 7996 7833 8012 8083
rect 8046 7833 8058 8083
rect 7996 7821 8058 7833
rect -1960 6283 -1898 6295
rect -1960 6033 -1948 6283
rect -1914 6033 -1898 6283
rect -1960 6021 -1898 6033
rect -1868 6283 -1802 6295
rect -1868 6033 -1852 6283
rect -1818 6033 -1802 6283
rect -1868 6021 -1802 6033
rect -1772 6283 -1706 6295
rect -1772 6033 -1756 6283
rect -1722 6033 -1706 6283
rect -1772 6021 -1706 6033
rect -1676 6283 -1610 6295
rect -1676 6033 -1660 6283
rect -1626 6033 -1610 6283
rect -1676 6021 -1610 6033
rect -1580 6283 -1514 6295
rect -1580 6033 -1564 6283
rect -1530 6033 -1514 6283
rect -1580 6021 -1514 6033
rect -1484 6283 -1418 6295
rect -1484 6033 -1468 6283
rect -1434 6033 -1418 6283
rect -1484 6021 -1418 6033
rect -1388 6283 -1322 6295
rect -1388 6033 -1372 6283
rect -1338 6033 -1322 6283
rect -1388 6021 -1322 6033
rect -1292 6283 -1226 6295
rect -1292 6033 -1276 6283
rect -1242 6033 -1226 6283
rect -1292 6021 -1226 6033
rect -1196 6283 -1130 6295
rect -1196 6033 -1180 6283
rect -1146 6033 -1130 6283
rect -1196 6021 -1130 6033
rect -1100 6283 -1034 6295
rect -1100 6033 -1084 6283
rect -1050 6033 -1034 6283
rect -1100 6021 -1034 6033
rect -1004 6283 -942 6295
rect -1004 6033 -988 6283
rect -954 6033 -942 6283
rect -1004 6021 -942 6033
rect 7040 6283 7102 6295
rect 7040 6033 7052 6283
rect 7086 6033 7102 6283
rect 7040 6021 7102 6033
rect 7132 6283 7198 6295
rect 7132 6033 7148 6283
rect 7182 6033 7198 6283
rect 7132 6021 7198 6033
rect 7228 6283 7294 6295
rect 7228 6033 7244 6283
rect 7278 6033 7294 6283
rect 7228 6021 7294 6033
rect 7324 6283 7390 6295
rect 7324 6033 7340 6283
rect 7374 6033 7390 6283
rect 7324 6021 7390 6033
rect 7420 6283 7486 6295
rect 7420 6033 7436 6283
rect 7470 6033 7486 6283
rect 7420 6021 7486 6033
rect 7516 6283 7582 6295
rect 7516 6033 7532 6283
rect 7566 6033 7582 6283
rect 7516 6021 7582 6033
rect 7612 6283 7678 6295
rect 7612 6033 7628 6283
rect 7662 6033 7678 6283
rect 7612 6021 7678 6033
rect 7708 6283 7774 6295
rect 7708 6033 7724 6283
rect 7758 6033 7774 6283
rect 7708 6021 7774 6033
rect 7804 6283 7870 6295
rect 7804 6033 7820 6283
rect 7854 6033 7870 6283
rect 7804 6021 7870 6033
rect 7900 6283 7966 6295
rect 7900 6033 7916 6283
rect 7950 6033 7966 6283
rect 7900 6021 7966 6033
rect 7996 6283 8058 6295
rect 7996 6033 8012 6283
rect 8046 6033 8058 6283
rect 7996 6021 8058 6033
rect -1960 4483 -1898 4495
rect -1960 4233 -1948 4483
rect -1914 4233 -1898 4483
rect -1960 4221 -1898 4233
rect -1868 4483 -1802 4495
rect -1868 4233 -1852 4483
rect -1818 4233 -1802 4483
rect -1868 4221 -1802 4233
rect -1772 4483 -1706 4495
rect -1772 4233 -1756 4483
rect -1722 4233 -1706 4483
rect -1772 4221 -1706 4233
rect -1676 4483 -1610 4495
rect -1676 4233 -1660 4483
rect -1626 4233 -1610 4483
rect -1676 4221 -1610 4233
rect -1580 4483 -1514 4495
rect -1580 4233 -1564 4483
rect -1530 4233 -1514 4483
rect -1580 4221 -1514 4233
rect -1484 4483 -1418 4495
rect -1484 4233 -1468 4483
rect -1434 4233 -1418 4483
rect -1484 4221 -1418 4233
rect -1388 4483 -1322 4495
rect -1388 4233 -1372 4483
rect -1338 4233 -1322 4483
rect -1388 4221 -1322 4233
rect -1292 4483 -1226 4495
rect -1292 4233 -1276 4483
rect -1242 4233 -1226 4483
rect -1292 4221 -1226 4233
rect -1196 4483 -1130 4495
rect -1196 4233 -1180 4483
rect -1146 4233 -1130 4483
rect -1196 4221 -1130 4233
rect -1100 4483 -1034 4495
rect -1100 4233 -1084 4483
rect -1050 4233 -1034 4483
rect -1100 4221 -1034 4233
rect -1004 4483 -942 4495
rect -1004 4233 -988 4483
rect -954 4233 -942 4483
rect -1004 4221 -942 4233
rect 7040 4483 7102 4495
rect 7040 4233 7052 4483
rect 7086 4233 7102 4483
rect 7040 4221 7102 4233
rect 7132 4483 7198 4495
rect 7132 4233 7148 4483
rect 7182 4233 7198 4483
rect 7132 4221 7198 4233
rect 7228 4483 7294 4495
rect 7228 4233 7244 4483
rect 7278 4233 7294 4483
rect 7228 4221 7294 4233
rect 7324 4483 7390 4495
rect 7324 4233 7340 4483
rect 7374 4233 7390 4483
rect 7324 4221 7390 4233
rect 7420 4483 7486 4495
rect 7420 4233 7436 4483
rect 7470 4233 7486 4483
rect 7420 4221 7486 4233
rect 7516 4483 7582 4495
rect 7516 4233 7532 4483
rect 7566 4233 7582 4483
rect 7516 4221 7582 4233
rect 7612 4483 7678 4495
rect 7612 4233 7628 4483
rect 7662 4233 7678 4483
rect 7612 4221 7678 4233
rect 7708 4483 7774 4495
rect 7708 4233 7724 4483
rect 7758 4233 7774 4483
rect 7708 4221 7774 4233
rect 7804 4483 7870 4495
rect 7804 4233 7820 4483
rect 7854 4233 7870 4483
rect 7804 4221 7870 4233
rect 7900 4483 7966 4495
rect 7900 4233 7916 4483
rect 7950 4233 7966 4483
rect 7900 4221 7966 4233
rect 7996 4483 8058 4495
rect 7996 4233 8012 4483
rect 8046 4233 8058 4483
rect 7996 4221 8058 4233
rect -1960 2683 -1898 2695
rect -1960 2433 -1948 2683
rect -1914 2433 -1898 2683
rect -1960 2421 -1898 2433
rect -1868 2683 -1802 2695
rect -1868 2433 -1852 2683
rect -1818 2433 -1802 2683
rect -1868 2421 -1802 2433
rect -1772 2683 -1706 2695
rect -1772 2433 -1756 2683
rect -1722 2433 -1706 2683
rect -1772 2421 -1706 2433
rect -1676 2683 -1610 2695
rect -1676 2433 -1660 2683
rect -1626 2433 -1610 2683
rect -1676 2421 -1610 2433
rect -1580 2683 -1514 2695
rect -1580 2433 -1564 2683
rect -1530 2433 -1514 2683
rect -1580 2421 -1514 2433
rect -1484 2683 -1418 2695
rect -1484 2433 -1468 2683
rect -1434 2433 -1418 2683
rect -1484 2421 -1418 2433
rect -1388 2683 -1322 2695
rect -1388 2433 -1372 2683
rect -1338 2433 -1322 2683
rect -1388 2421 -1322 2433
rect -1292 2683 -1226 2695
rect -1292 2433 -1276 2683
rect -1242 2433 -1226 2683
rect -1292 2421 -1226 2433
rect -1196 2683 -1130 2695
rect -1196 2433 -1180 2683
rect -1146 2433 -1130 2683
rect -1196 2421 -1130 2433
rect -1100 2683 -1034 2695
rect -1100 2433 -1084 2683
rect -1050 2433 -1034 2683
rect -1100 2421 -1034 2433
rect -1004 2683 -942 2695
rect -1004 2433 -988 2683
rect -954 2433 -942 2683
rect -1004 2421 -942 2433
rect 7040 2683 7102 2695
rect 7040 2433 7052 2683
rect 7086 2433 7102 2683
rect 7040 2421 7102 2433
rect 7132 2683 7198 2695
rect 7132 2433 7148 2683
rect 7182 2433 7198 2683
rect 7132 2421 7198 2433
rect 7228 2683 7294 2695
rect 7228 2433 7244 2683
rect 7278 2433 7294 2683
rect 7228 2421 7294 2433
rect 7324 2683 7390 2695
rect 7324 2433 7340 2683
rect 7374 2433 7390 2683
rect 7324 2421 7390 2433
rect 7420 2683 7486 2695
rect 7420 2433 7436 2683
rect 7470 2433 7486 2683
rect 7420 2421 7486 2433
rect 7516 2683 7582 2695
rect 7516 2433 7532 2683
rect 7566 2433 7582 2683
rect 7516 2421 7582 2433
rect 7612 2683 7678 2695
rect 7612 2433 7628 2683
rect 7662 2433 7678 2683
rect 7612 2421 7678 2433
rect 7708 2683 7774 2695
rect 7708 2433 7724 2683
rect 7758 2433 7774 2683
rect 7708 2421 7774 2433
rect 7804 2683 7870 2695
rect 7804 2433 7820 2683
rect 7854 2433 7870 2683
rect 7804 2421 7870 2433
rect 7900 2683 7966 2695
rect 7900 2433 7916 2683
rect 7950 2433 7966 2683
rect 7900 2421 7966 2433
rect 7996 2683 8058 2695
rect 7996 2433 8012 2683
rect 8046 2433 8058 2683
rect 7996 2421 8058 2433
rect -1960 883 -1898 895
rect -1960 633 -1948 883
rect -1914 633 -1898 883
rect -1960 621 -1898 633
rect -1868 883 -1802 895
rect -1868 633 -1852 883
rect -1818 633 -1802 883
rect -1868 621 -1802 633
rect -1772 883 -1706 895
rect -1772 633 -1756 883
rect -1722 633 -1706 883
rect -1772 621 -1706 633
rect -1676 883 -1610 895
rect -1676 633 -1660 883
rect -1626 633 -1610 883
rect -1676 621 -1610 633
rect -1580 883 -1514 895
rect -1580 633 -1564 883
rect -1530 633 -1514 883
rect -1580 621 -1514 633
rect -1484 883 -1418 895
rect -1484 633 -1468 883
rect -1434 633 -1418 883
rect -1484 621 -1418 633
rect -1388 883 -1322 895
rect -1388 633 -1372 883
rect -1338 633 -1322 883
rect -1388 621 -1322 633
rect -1292 883 -1226 895
rect -1292 633 -1276 883
rect -1242 633 -1226 883
rect -1292 621 -1226 633
rect -1196 883 -1130 895
rect -1196 633 -1180 883
rect -1146 633 -1130 883
rect -1196 621 -1130 633
rect -1100 883 -1034 895
rect -1100 633 -1084 883
rect -1050 633 -1034 883
rect -1100 621 -1034 633
rect -1004 883 -942 895
rect -1004 633 -988 883
rect -954 633 -942 883
rect -1004 621 -942 633
rect 7040 883 7102 895
rect 7040 633 7052 883
rect 7086 633 7102 883
rect 7040 621 7102 633
rect 7132 883 7198 895
rect 7132 633 7148 883
rect 7182 633 7198 883
rect 7132 621 7198 633
rect 7228 883 7294 895
rect 7228 633 7244 883
rect 7278 633 7294 883
rect 7228 621 7294 633
rect 7324 883 7390 895
rect 7324 633 7340 883
rect 7374 633 7390 883
rect 7324 621 7390 633
rect 7420 883 7486 895
rect 7420 633 7436 883
rect 7470 633 7486 883
rect 7420 621 7486 633
rect 7516 883 7582 895
rect 7516 633 7532 883
rect 7566 633 7582 883
rect 7516 621 7582 633
rect 7612 883 7678 895
rect 7612 633 7628 883
rect 7662 633 7678 883
rect 7612 621 7678 633
rect 7708 883 7774 895
rect 7708 633 7724 883
rect 7758 633 7774 883
rect 7708 621 7774 633
rect 7804 883 7870 895
rect 7804 633 7820 883
rect 7854 633 7870 883
rect 7804 621 7870 633
rect 7900 883 7966 895
rect 7900 633 7916 883
rect 7950 633 7966 883
rect 7900 621 7966 633
rect 7996 883 8058 895
rect 7996 633 8012 883
rect 8046 633 8058 883
rect 7996 621 8058 633
rect -1960 -917 -1898 -905
rect -1960 -1167 -1948 -917
rect -1914 -1167 -1898 -917
rect -1960 -1179 -1898 -1167
rect -1868 -917 -1802 -905
rect -1868 -1167 -1852 -917
rect -1818 -1167 -1802 -917
rect -1868 -1179 -1802 -1167
rect -1772 -917 -1706 -905
rect -1772 -1167 -1756 -917
rect -1722 -1167 -1706 -917
rect -1772 -1179 -1706 -1167
rect -1676 -917 -1610 -905
rect -1676 -1167 -1660 -917
rect -1626 -1167 -1610 -917
rect -1676 -1179 -1610 -1167
rect -1580 -917 -1514 -905
rect -1580 -1167 -1564 -917
rect -1530 -1167 -1514 -917
rect -1580 -1179 -1514 -1167
rect -1484 -917 -1418 -905
rect -1484 -1167 -1468 -917
rect -1434 -1167 -1418 -917
rect -1484 -1179 -1418 -1167
rect -1388 -917 -1322 -905
rect -1388 -1167 -1372 -917
rect -1338 -1167 -1322 -917
rect -1388 -1179 -1322 -1167
rect -1292 -917 -1226 -905
rect -1292 -1167 -1276 -917
rect -1242 -1167 -1226 -917
rect -1292 -1179 -1226 -1167
rect -1196 -917 -1130 -905
rect -1196 -1167 -1180 -917
rect -1146 -1167 -1130 -917
rect -1196 -1179 -1130 -1167
rect -1100 -917 -1034 -905
rect -1100 -1167 -1084 -917
rect -1050 -1167 -1034 -917
rect -1100 -1179 -1034 -1167
rect -1004 -917 -942 -905
rect -1004 -1167 -988 -917
rect -954 -1167 -942 -917
rect -1004 -1179 -942 -1167
rect 7040 -917 7102 -905
rect 7040 -1167 7052 -917
rect 7086 -1167 7102 -917
rect 7040 -1179 7102 -1167
rect 7132 -917 7198 -905
rect 7132 -1167 7148 -917
rect 7182 -1167 7198 -917
rect 7132 -1179 7198 -1167
rect 7228 -917 7294 -905
rect 7228 -1167 7244 -917
rect 7278 -1167 7294 -917
rect 7228 -1179 7294 -1167
rect 7324 -917 7390 -905
rect 7324 -1167 7340 -917
rect 7374 -1167 7390 -917
rect 7324 -1179 7390 -1167
rect 7420 -917 7486 -905
rect 7420 -1167 7436 -917
rect 7470 -1167 7486 -917
rect 7420 -1179 7486 -1167
rect 7516 -917 7582 -905
rect 7516 -1167 7532 -917
rect 7566 -1167 7582 -917
rect 7516 -1179 7582 -1167
rect 7612 -917 7678 -905
rect 7612 -1167 7628 -917
rect 7662 -1167 7678 -917
rect 7612 -1179 7678 -1167
rect 7708 -917 7774 -905
rect 7708 -1167 7724 -917
rect 7758 -1167 7774 -917
rect 7708 -1179 7774 -1167
rect 7804 -917 7870 -905
rect 7804 -1167 7820 -917
rect 7854 -1167 7870 -917
rect 7804 -1179 7870 -1167
rect 7900 -917 7966 -905
rect 7900 -1167 7916 -917
rect 7950 -1167 7966 -917
rect 7900 -1179 7966 -1167
rect 7996 -917 8058 -905
rect 7996 -1167 8012 -917
rect 8046 -1167 8058 -917
rect 7996 -1179 8058 -1167
<< ndiffc >>
rect -1948 7422 -1914 7504
rect -1852 7422 -1818 7504
rect -1756 7422 -1722 7504
rect -1660 7422 -1626 7504
rect -1564 7422 -1530 7504
rect -1468 7422 -1434 7504
rect -1372 7422 -1338 7504
rect -1276 7422 -1242 7504
rect -1180 7422 -1146 7504
rect -1084 7422 -1050 7504
rect -988 7422 -954 7504
rect 7052 7422 7086 7504
rect 7148 7422 7182 7504
rect 7244 7422 7278 7504
rect 7340 7422 7374 7504
rect 7436 7422 7470 7504
rect 7532 7422 7566 7504
rect 7628 7422 7662 7504
rect 7724 7422 7758 7504
rect 7820 7422 7854 7504
rect 7916 7422 7950 7504
rect 8012 7422 8046 7504
rect -1948 5622 -1914 5704
rect -1852 5622 -1818 5704
rect -1756 5622 -1722 5704
rect -1660 5622 -1626 5704
rect -1564 5622 -1530 5704
rect -1468 5622 -1434 5704
rect -1372 5622 -1338 5704
rect -1276 5622 -1242 5704
rect -1180 5622 -1146 5704
rect -1084 5622 -1050 5704
rect -988 5622 -954 5704
rect 7052 5622 7086 5704
rect 7148 5622 7182 5704
rect 7244 5622 7278 5704
rect 7340 5622 7374 5704
rect 7436 5622 7470 5704
rect 7532 5622 7566 5704
rect 7628 5622 7662 5704
rect 7724 5622 7758 5704
rect 7820 5622 7854 5704
rect 7916 5622 7950 5704
rect 8012 5622 8046 5704
rect -1948 3822 -1914 3904
rect -1852 3822 -1818 3904
rect -1756 3822 -1722 3904
rect -1660 3822 -1626 3904
rect -1564 3822 -1530 3904
rect -1468 3822 -1434 3904
rect -1372 3822 -1338 3904
rect -1276 3822 -1242 3904
rect -1180 3822 -1146 3904
rect -1084 3822 -1050 3904
rect -988 3822 -954 3904
rect 7052 3822 7086 3904
rect 7148 3822 7182 3904
rect 7244 3822 7278 3904
rect 7340 3822 7374 3904
rect 7436 3822 7470 3904
rect 7532 3822 7566 3904
rect 7628 3822 7662 3904
rect 7724 3822 7758 3904
rect 7820 3822 7854 3904
rect 7916 3822 7950 3904
rect 8012 3822 8046 3904
rect -1948 2022 -1914 2104
rect -1852 2022 -1818 2104
rect -1756 2022 -1722 2104
rect -1660 2022 -1626 2104
rect -1564 2022 -1530 2104
rect -1468 2022 -1434 2104
rect -1372 2022 -1338 2104
rect -1276 2022 -1242 2104
rect -1180 2022 -1146 2104
rect -1084 2022 -1050 2104
rect -988 2022 -954 2104
rect 7052 2022 7086 2104
rect 7148 2022 7182 2104
rect 7244 2022 7278 2104
rect 7340 2022 7374 2104
rect 7436 2022 7470 2104
rect 7532 2022 7566 2104
rect 7628 2022 7662 2104
rect 7724 2022 7758 2104
rect 7820 2022 7854 2104
rect 7916 2022 7950 2104
rect 8012 2022 8046 2104
rect -1948 222 -1914 304
rect -1852 222 -1818 304
rect -1756 222 -1722 304
rect -1660 222 -1626 304
rect -1564 222 -1530 304
rect -1468 222 -1434 304
rect -1372 222 -1338 304
rect -1276 222 -1242 304
rect -1180 222 -1146 304
rect -1084 222 -1050 304
rect -988 222 -954 304
rect 7052 222 7086 304
rect 7148 222 7182 304
rect 7244 222 7278 304
rect 7340 222 7374 304
rect 7436 222 7470 304
rect 7532 222 7566 304
rect 7628 222 7662 304
rect 7724 222 7758 304
rect 7820 222 7854 304
rect 7916 222 7950 304
rect 8012 222 8046 304
rect -1948 -1578 -1914 -1496
rect -1852 -1578 -1818 -1496
rect -1756 -1578 -1722 -1496
rect -1660 -1578 -1626 -1496
rect -1564 -1578 -1530 -1496
rect -1468 -1578 -1434 -1496
rect -1372 -1578 -1338 -1496
rect -1276 -1578 -1242 -1496
rect -1180 -1578 -1146 -1496
rect -1084 -1578 -1050 -1496
rect -988 -1578 -954 -1496
rect 7052 -1578 7086 -1496
rect 7148 -1578 7182 -1496
rect 7244 -1578 7278 -1496
rect 7340 -1578 7374 -1496
rect 7436 -1578 7470 -1496
rect 7532 -1578 7566 -1496
rect 7628 -1578 7662 -1496
rect 7724 -1578 7758 -1496
rect 7820 -1578 7854 -1496
rect 7916 -1578 7950 -1496
rect 8012 -1578 8046 -1496
<< pdiffc >>
rect -1948 7833 -1914 8083
rect -1852 7833 -1818 8083
rect -1756 7833 -1722 8083
rect -1660 7833 -1626 8083
rect -1564 7833 -1530 8083
rect -1468 7833 -1434 8083
rect -1372 7833 -1338 8083
rect -1276 7833 -1242 8083
rect -1180 7833 -1146 8083
rect -1084 7833 -1050 8083
rect -988 7833 -954 8083
rect 7052 7833 7086 8083
rect 7148 7833 7182 8083
rect 7244 7833 7278 8083
rect 7340 7833 7374 8083
rect 7436 7833 7470 8083
rect 7532 7833 7566 8083
rect 7628 7833 7662 8083
rect 7724 7833 7758 8083
rect 7820 7833 7854 8083
rect 7916 7833 7950 8083
rect 8012 7833 8046 8083
rect -1948 6033 -1914 6283
rect -1852 6033 -1818 6283
rect -1756 6033 -1722 6283
rect -1660 6033 -1626 6283
rect -1564 6033 -1530 6283
rect -1468 6033 -1434 6283
rect -1372 6033 -1338 6283
rect -1276 6033 -1242 6283
rect -1180 6033 -1146 6283
rect -1084 6033 -1050 6283
rect -988 6033 -954 6283
rect 7052 6033 7086 6283
rect 7148 6033 7182 6283
rect 7244 6033 7278 6283
rect 7340 6033 7374 6283
rect 7436 6033 7470 6283
rect 7532 6033 7566 6283
rect 7628 6033 7662 6283
rect 7724 6033 7758 6283
rect 7820 6033 7854 6283
rect 7916 6033 7950 6283
rect 8012 6033 8046 6283
rect -1948 4233 -1914 4483
rect -1852 4233 -1818 4483
rect -1756 4233 -1722 4483
rect -1660 4233 -1626 4483
rect -1564 4233 -1530 4483
rect -1468 4233 -1434 4483
rect -1372 4233 -1338 4483
rect -1276 4233 -1242 4483
rect -1180 4233 -1146 4483
rect -1084 4233 -1050 4483
rect -988 4233 -954 4483
rect 7052 4233 7086 4483
rect 7148 4233 7182 4483
rect 7244 4233 7278 4483
rect 7340 4233 7374 4483
rect 7436 4233 7470 4483
rect 7532 4233 7566 4483
rect 7628 4233 7662 4483
rect 7724 4233 7758 4483
rect 7820 4233 7854 4483
rect 7916 4233 7950 4483
rect 8012 4233 8046 4483
rect -1948 2433 -1914 2683
rect -1852 2433 -1818 2683
rect -1756 2433 -1722 2683
rect -1660 2433 -1626 2683
rect -1564 2433 -1530 2683
rect -1468 2433 -1434 2683
rect -1372 2433 -1338 2683
rect -1276 2433 -1242 2683
rect -1180 2433 -1146 2683
rect -1084 2433 -1050 2683
rect -988 2433 -954 2683
rect 7052 2433 7086 2683
rect 7148 2433 7182 2683
rect 7244 2433 7278 2683
rect 7340 2433 7374 2683
rect 7436 2433 7470 2683
rect 7532 2433 7566 2683
rect 7628 2433 7662 2683
rect 7724 2433 7758 2683
rect 7820 2433 7854 2683
rect 7916 2433 7950 2683
rect 8012 2433 8046 2683
rect -1948 633 -1914 883
rect -1852 633 -1818 883
rect -1756 633 -1722 883
rect -1660 633 -1626 883
rect -1564 633 -1530 883
rect -1468 633 -1434 883
rect -1372 633 -1338 883
rect -1276 633 -1242 883
rect -1180 633 -1146 883
rect -1084 633 -1050 883
rect -988 633 -954 883
rect 7052 633 7086 883
rect 7148 633 7182 883
rect 7244 633 7278 883
rect 7340 633 7374 883
rect 7436 633 7470 883
rect 7532 633 7566 883
rect 7628 633 7662 883
rect 7724 633 7758 883
rect 7820 633 7854 883
rect 7916 633 7950 883
rect 8012 633 8046 883
rect -1948 -1167 -1914 -917
rect -1852 -1167 -1818 -917
rect -1756 -1167 -1722 -917
rect -1660 -1167 -1626 -917
rect -1564 -1167 -1530 -917
rect -1468 -1167 -1434 -917
rect -1372 -1167 -1338 -917
rect -1276 -1167 -1242 -917
rect -1180 -1167 -1146 -917
rect -1084 -1167 -1050 -917
rect -988 -1167 -954 -917
rect 7052 -1167 7086 -917
rect 7148 -1167 7182 -917
rect 7244 -1167 7278 -917
rect 7340 -1167 7374 -917
rect 7436 -1167 7470 -917
rect 7532 -1167 7566 -917
rect 7628 -1167 7662 -917
rect 7724 -1167 7758 -917
rect 7820 -1167 7854 -917
rect 7916 -1167 7950 -917
rect 8012 -1167 8046 -917
<< psubdiff >>
rect -2062 7594 -1966 7628
rect -936 7594 -840 7628
rect -2062 7532 -2028 7594
rect -874 7532 -840 7594
rect -2062 7270 -2028 7332
rect -874 7270 -840 7332
rect -2062 7236 -1966 7270
rect -936 7236 -840 7270
rect 6938 7594 7034 7628
rect 8064 7594 8160 7628
rect 6938 7532 6972 7594
rect 8126 7532 8160 7594
rect 6938 7270 6972 7332
rect 8126 7270 8160 7332
rect 6938 7236 7034 7270
rect 8064 7236 8160 7270
rect -2062 5794 -1966 5828
rect -936 5794 -840 5828
rect -2062 5732 -2028 5794
rect -874 5732 -840 5794
rect -2062 5470 -2028 5532
rect -874 5470 -840 5532
rect -2062 5436 -1966 5470
rect -936 5436 -840 5470
rect 6938 5794 7034 5828
rect 8064 5794 8160 5828
rect 6938 5732 6972 5794
rect 8126 5732 8160 5794
rect 6938 5470 6972 5532
rect 8126 5470 8160 5532
rect 6938 5436 7034 5470
rect 8064 5436 8160 5470
rect -2062 3994 -1966 4028
rect -936 3994 -840 4028
rect -2062 3932 -2028 3994
rect -874 3932 -840 3994
rect -2062 3670 -2028 3732
rect -874 3670 -840 3732
rect -2062 3636 -1966 3670
rect -936 3636 -840 3670
rect 6938 3994 7034 4028
rect 8064 3994 8160 4028
rect 6938 3932 6972 3994
rect 8126 3932 8160 3994
rect 6938 3670 6972 3732
rect 8126 3670 8160 3732
rect 6938 3636 7034 3670
rect 8064 3636 8160 3670
rect -2062 2194 -1966 2228
rect -936 2194 -840 2228
rect -2062 2132 -2028 2194
rect -874 2132 -840 2194
rect -2062 1870 -2028 1932
rect -874 1870 -840 1932
rect -2062 1836 -1966 1870
rect -936 1836 -840 1870
rect 6938 2194 7034 2228
rect 8064 2194 8160 2228
rect 6938 2132 6972 2194
rect 8126 2132 8160 2194
rect 6938 1870 6972 1932
rect 8126 1870 8160 1932
rect 6938 1836 7034 1870
rect 8064 1836 8160 1870
rect -2062 394 -1966 428
rect -936 394 -840 428
rect -2062 332 -2028 394
rect -874 332 -840 394
rect -2062 70 -2028 132
rect -874 70 -840 132
rect -2062 36 -1966 70
rect -936 36 -840 70
rect 6938 394 7034 428
rect 8064 394 8160 428
rect 6938 332 6972 394
rect 8126 332 8160 394
rect 6938 70 6972 132
rect 8126 70 8160 132
rect 6938 36 7034 70
rect 8064 36 8160 70
rect -2062 -1406 -1966 -1372
rect -936 -1406 -840 -1372
rect -2062 -1468 -2028 -1406
rect -874 -1468 -840 -1406
rect -2062 -1730 -2028 -1668
rect -874 -1730 -840 -1668
rect -2062 -1764 -1966 -1730
rect -936 -1764 -840 -1730
rect 6938 -1406 7034 -1372
rect 8064 -1406 8160 -1372
rect 6938 -1468 6972 -1406
rect 8126 -1468 8160 -1406
rect 6938 -1730 6972 -1668
rect 8126 -1730 8160 -1668
rect 6938 -1764 7034 -1730
rect 8064 -1764 8160 -1730
<< nsubdiff >>
rect -2062 8244 -1966 8278
rect -936 8244 -840 8278
rect -2062 8182 -2028 8244
rect -874 8182 -840 8244
rect -2062 7734 -2028 7796
rect -874 7734 -840 7796
rect -2062 7700 -1966 7734
rect -936 7700 -840 7734
rect 6938 8244 7034 8278
rect 8064 8244 8160 8278
rect 6938 8182 6972 8244
rect 8126 8182 8160 8244
rect 6938 7734 6972 7796
rect 8126 7734 8160 7796
rect 6938 7700 7034 7734
rect 8064 7700 8160 7734
rect -2062 6444 -1966 6478
rect -936 6444 -840 6478
rect -2062 6382 -2028 6444
rect -874 6382 -840 6444
rect -2062 5934 -2028 5996
rect -874 5934 -840 5996
rect -2062 5900 -1966 5934
rect -936 5900 -840 5934
rect 6938 6444 7034 6478
rect 8064 6444 8160 6478
rect 6938 6382 6972 6444
rect 8126 6382 8160 6444
rect 6938 5934 6972 5996
rect 8126 5934 8160 5996
rect 6938 5900 7034 5934
rect 8064 5900 8160 5934
rect -2062 4644 -1966 4678
rect -936 4644 -840 4678
rect -2062 4582 -2028 4644
rect -874 4582 -840 4644
rect -2062 4134 -2028 4196
rect -874 4134 -840 4196
rect -2062 4100 -1966 4134
rect -936 4100 -840 4134
rect 6938 4644 7034 4678
rect 8064 4644 8160 4678
rect 6938 4582 6972 4644
rect 8126 4582 8160 4644
rect 6938 4134 6972 4196
rect 8126 4134 8160 4196
rect 6938 4100 7034 4134
rect 8064 4100 8160 4134
rect -2062 2844 -1966 2878
rect -936 2844 -840 2878
rect -2062 2782 -2028 2844
rect -874 2782 -840 2844
rect -2062 2334 -2028 2396
rect -874 2334 -840 2396
rect -2062 2300 -1966 2334
rect -936 2300 -840 2334
rect 6938 2844 7034 2878
rect 8064 2844 8160 2878
rect 6938 2782 6972 2844
rect 8126 2782 8160 2844
rect 6938 2334 6972 2396
rect 8126 2334 8160 2396
rect 6938 2300 7034 2334
rect 8064 2300 8160 2334
rect -2062 1044 -1966 1078
rect -936 1044 -840 1078
rect -2062 982 -2028 1044
rect -874 982 -840 1044
rect -2062 534 -2028 596
rect -874 534 -840 596
rect -2062 500 -1966 534
rect -936 500 -840 534
rect 6938 1044 7034 1078
rect 8064 1044 8160 1078
rect 6938 982 6972 1044
rect 8126 982 8160 1044
rect 6938 534 6972 596
rect 8126 534 8160 596
rect 6938 500 7034 534
rect 8064 500 8160 534
rect -2062 -756 -1966 -722
rect -936 -756 -840 -722
rect -2062 -818 -2028 -756
rect -874 -818 -840 -756
rect -2062 -1266 -2028 -1204
rect -874 -1266 -840 -1204
rect -2062 -1300 -1966 -1266
rect -936 -1300 -840 -1266
rect 6938 -756 7034 -722
rect 8064 -756 8160 -722
rect 6938 -818 6972 -756
rect 8126 -818 8160 -756
rect 6938 -1266 6972 -1204
rect 8126 -1266 8160 -1204
rect 6938 -1300 7034 -1266
rect 8064 -1300 8160 -1266
<< psubdiffcont >>
rect -1966 7594 -936 7628
rect -2062 7332 -2028 7532
rect -874 7332 -840 7532
rect -1966 7236 -936 7270
rect 7034 7594 8064 7628
rect 6938 7332 6972 7532
rect 8126 7332 8160 7532
rect 7034 7236 8064 7270
rect -1966 5794 -936 5828
rect -2062 5532 -2028 5732
rect -874 5532 -840 5732
rect -1966 5436 -936 5470
rect 7034 5794 8064 5828
rect 6938 5532 6972 5732
rect 8126 5532 8160 5732
rect 7034 5436 8064 5470
rect -1966 3994 -936 4028
rect -2062 3732 -2028 3932
rect -874 3732 -840 3932
rect -1966 3636 -936 3670
rect 7034 3994 8064 4028
rect 6938 3732 6972 3932
rect 8126 3732 8160 3932
rect 7034 3636 8064 3670
rect -1966 2194 -936 2228
rect -2062 1932 -2028 2132
rect -874 1932 -840 2132
rect -1966 1836 -936 1870
rect 7034 2194 8064 2228
rect 6938 1932 6972 2132
rect 8126 1932 8160 2132
rect 7034 1836 8064 1870
rect -1966 394 -936 428
rect -2062 132 -2028 332
rect -874 132 -840 332
rect -1966 36 -936 70
rect 7034 394 8064 428
rect 6938 132 6972 332
rect 8126 132 8160 332
rect 7034 36 8064 70
rect -1966 -1406 -936 -1372
rect -2062 -1668 -2028 -1468
rect -874 -1668 -840 -1468
rect -1966 -1764 -936 -1730
rect 7034 -1406 8064 -1372
rect 6938 -1668 6972 -1468
rect 8126 -1668 8160 -1468
rect 7034 -1764 8064 -1730
<< nsubdiffcont >>
rect -1966 8244 -936 8278
rect -2062 7796 -2028 8182
rect -874 7796 -840 8182
rect -1966 7700 -936 7734
rect 7034 8244 8064 8278
rect 6938 7796 6972 8182
rect 8126 7796 8160 8182
rect 7034 7700 8064 7734
rect -1966 6444 -936 6478
rect -2062 5996 -2028 6382
rect -874 5996 -840 6382
rect -1966 5900 -936 5934
rect 7034 6444 8064 6478
rect 6938 5996 6972 6382
rect 8126 5996 8160 6382
rect 7034 5900 8064 5934
rect -1966 4644 -936 4678
rect -2062 4196 -2028 4582
rect -874 4196 -840 4582
rect -1966 4100 -936 4134
rect 7034 4644 8064 4678
rect 6938 4196 6972 4582
rect 8126 4196 8160 4582
rect 7034 4100 8064 4134
rect -1966 2844 -936 2878
rect -2062 2396 -2028 2782
rect -874 2396 -840 2782
rect -1966 2300 -936 2334
rect 7034 2844 8064 2878
rect 6938 2396 6972 2782
rect 8126 2396 8160 2782
rect 7034 2300 8064 2334
rect -1966 1044 -936 1078
rect -2062 596 -2028 982
rect -874 596 -840 982
rect -1966 500 -936 534
rect 7034 1044 8064 1078
rect 6938 596 6972 982
rect 8126 596 8160 982
rect 7034 500 8064 534
rect -1966 -756 -936 -722
rect -2062 -1204 -2028 -818
rect -874 -1204 -840 -818
rect -1966 -1300 -936 -1266
rect 7034 -756 8064 -722
rect 6938 -1204 6972 -818
rect 8126 -1204 8160 -818
rect 7034 -1300 8064 -1266
<< poly >>
rect -1964 8176 -938 8192
rect -1964 8142 -1948 8176
rect -1914 8142 -1756 8176
rect -1722 8142 -1564 8176
rect -1530 8142 -1372 8176
rect -1338 8142 -1180 8176
rect -1146 8142 -988 8176
rect -954 8142 -938 8176
rect -1964 8126 -938 8142
rect -1898 8095 -1868 8126
rect -1802 8095 -1772 8126
rect -1706 8095 -1676 8126
rect -1610 8095 -1580 8126
rect -1514 8095 -1484 8126
rect -1418 8095 -1388 8126
rect -1322 8095 -1292 8126
rect -1226 8095 -1196 8126
rect -1130 8095 -1100 8126
rect -1034 8095 -1004 8126
rect -1898 7795 -1868 7821
rect -1802 7795 -1772 7821
rect -1706 7795 -1676 7821
rect -1610 7795 -1580 7821
rect -1514 7795 -1484 7821
rect -1418 7795 -1388 7821
rect -1322 7795 -1292 7821
rect -1226 7795 -1196 7821
rect -1130 7795 -1100 7821
rect -1034 7795 -1004 7821
rect 7036 8176 8062 8192
rect 7036 8142 7052 8176
rect 7086 8142 7244 8176
rect 7278 8142 7436 8176
rect 7470 8142 7628 8176
rect 7662 8142 7820 8176
rect 7854 8142 8012 8176
rect 8046 8142 8062 8176
rect 7036 8126 8062 8142
rect 7102 8095 7132 8126
rect 7198 8095 7228 8126
rect 7294 8095 7324 8126
rect 7390 8095 7420 8126
rect 7486 8095 7516 8126
rect 7582 8095 7612 8126
rect 7678 8095 7708 8126
rect 7774 8095 7804 8126
rect 7870 8095 7900 8126
rect 7966 8095 7996 8126
rect 7102 7795 7132 7821
rect 7198 7795 7228 7821
rect 7294 7795 7324 7821
rect 7390 7795 7420 7821
rect 7486 7795 7516 7821
rect 7582 7795 7612 7821
rect 7678 7795 7708 7821
rect 7774 7795 7804 7821
rect 7870 7795 7900 7821
rect 7966 7795 7996 7821
rect -1898 7516 -1868 7542
rect -1802 7516 -1772 7542
rect -1706 7516 -1676 7542
rect -1610 7516 -1580 7542
rect -1514 7516 -1484 7542
rect -1418 7516 -1388 7542
rect -1322 7516 -1292 7542
rect -1226 7516 -1196 7542
rect -1130 7516 -1100 7542
rect -1034 7516 -1004 7542
rect -1898 7388 -1868 7410
rect -1802 7388 -1772 7410
rect -1706 7388 -1676 7410
rect -1610 7388 -1580 7410
rect -1514 7388 -1484 7410
rect -1418 7388 -1388 7410
rect -1322 7388 -1292 7410
rect -1226 7388 -1196 7410
rect -1130 7388 -1100 7410
rect -1034 7388 -1004 7410
rect -1964 7369 -938 7388
rect -1964 7335 -1948 7369
rect -1914 7335 -1756 7369
rect -1722 7335 -1564 7369
rect -1530 7335 -1372 7369
rect -1338 7335 -1180 7369
rect -1146 7335 -988 7369
rect -954 7335 -938 7369
rect -1964 7322 -938 7335
rect 7102 7516 7132 7542
rect 7198 7516 7228 7542
rect 7294 7516 7324 7542
rect 7390 7516 7420 7542
rect 7486 7516 7516 7542
rect 7582 7516 7612 7542
rect 7678 7516 7708 7542
rect 7774 7516 7804 7542
rect 7870 7516 7900 7542
rect 7966 7516 7996 7542
rect 7102 7388 7132 7410
rect 7198 7388 7228 7410
rect 7294 7388 7324 7410
rect 7390 7388 7420 7410
rect 7486 7388 7516 7410
rect 7582 7388 7612 7410
rect 7678 7388 7708 7410
rect 7774 7388 7804 7410
rect 7870 7388 7900 7410
rect 7966 7388 7996 7410
rect 7036 7369 8062 7388
rect 7036 7335 7052 7369
rect 7086 7335 7244 7369
rect 7278 7335 7436 7369
rect 7470 7335 7628 7369
rect 7662 7335 7820 7369
rect 7854 7335 8012 7369
rect 8046 7335 8062 7369
rect 7036 7322 8062 7335
rect -1964 6376 -938 6392
rect -1964 6342 -1948 6376
rect -1914 6342 -1756 6376
rect -1722 6342 -1564 6376
rect -1530 6342 -1372 6376
rect -1338 6342 -1180 6376
rect -1146 6342 -988 6376
rect -954 6342 -938 6376
rect -1964 6326 -938 6342
rect -1898 6295 -1868 6326
rect -1802 6295 -1772 6326
rect -1706 6295 -1676 6326
rect -1610 6295 -1580 6326
rect -1514 6295 -1484 6326
rect -1418 6295 -1388 6326
rect -1322 6295 -1292 6326
rect -1226 6295 -1196 6326
rect -1130 6295 -1100 6326
rect -1034 6295 -1004 6326
rect -1898 5995 -1868 6021
rect -1802 5995 -1772 6021
rect -1706 5995 -1676 6021
rect -1610 5995 -1580 6021
rect -1514 5995 -1484 6021
rect -1418 5995 -1388 6021
rect -1322 5995 -1292 6021
rect -1226 5995 -1196 6021
rect -1130 5995 -1100 6021
rect -1034 5995 -1004 6021
rect 7036 6376 8062 6392
rect 7036 6342 7052 6376
rect 7086 6342 7244 6376
rect 7278 6342 7436 6376
rect 7470 6342 7628 6376
rect 7662 6342 7820 6376
rect 7854 6342 8012 6376
rect 8046 6342 8062 6376
rect 7036 6326 8062 6342
rect 7102 6295 7132 6326
rect 7198 6295 7228 6326
rect 7294 6295 7324 6326
rect 7390 6295 7420 6326
rect 7486 6295 7516 6326
rect 7582 6295 7612 6326
rect 7678 6295 7708 6326
rect 7774 6295 7804 6326
rect 7870 6295 7900 6326
rect 7966 6295 7996 6326
rect 7102 5995 7132 6021
rect 7198 5995 7228 6021
rect 7294 5995 7324 6021
rect 7390 5995 7420 6021
rect 7486 5995 7516 6021
rect 7582 5995 7612 6021
rect 7678 5995 7708 6021
rect 7774 5995 7804 6021
rect 7870 5995 7900 6021
rect 7966 5995 7996 6021
rect -1898 5716 -1868 5742
rect -1802 5716 -1772 5742
rect -1706 5716 -1676 5742
rect -1610 5716 -1580 5742
rect -1514 5716 -1484 5742
rect -1418 5716 -1388 5742
rect -1322 5716 -1292 5742
rect -1226 5716 -1196 5742
rect -1130 5716 -1100 5742
rect -1034 5716 -1004 5742
rect -1898 5588 -1868 5610
rect -1802 5588 -1772 5610
rect -1706 5588 -1676 5610
rect -1610 5588 -1580 5610
rect -1514 5588 -1484 5610
rect -1418 5588 -1388 5610
rect -1322 5588 -1292 5610
rect -1226 5588 -1196 5610
rect -1130 5588 -1100 5610
rect -1034 5588 -1004 5610
rect -1964 5569 -938 5588
rect -1964 5535 -1948 5569
rect -1914 5535 -1756 5569
rect -1722 5535 -1564 5569
rect -1530 5535 -1372 5569
rect -1338 5535 -1180 5569
rect -1146 5535 -988 5569
rect -954 5535 -938 5569
rect -1964 5522 -938 5535
rect 7102 5716 7132 5742
rect 7198 5716 7228 5742
rect 7294 5716 7324 5742
rect 7390 5716 7420 5742
rect 7486 5716 7516 5742
rect 7582 5716 7612 5742
rect 7678 5716 7708 5742
rect 7774 5716 7804 5742
rect 7870 5716 7900 5742
rect 7966 5716 7996 5742
rect 7102 5588 7132 5610
rect 7198 5588 7228 5610
rect 7294 5588 7324 5610
rect 7390 5588 7420 5610
rect 7486 5588 7516 5610
rect 7582 5588 7612 5610
rect 7678 5588 7708 5610
rect 7774 5588 7804 5610
rect 7870 5588 7900 5610
rect 7966 5588 7996 5610
rect 7036 5569 8062 5588
rect 7036 5535 7052 5569
rect 7086 5535 7244 5569
rect 7278 5535 7436 5569
rect 7470 5535 7628 5569
rect 7662 5535 7820 5569
rect 7854 5535 8012 5569
rect 8046 5535 8062 5569
rect 7036 5522 8062 5535
rect -1964 4576 -938 4592
rect -1964 4542 -1948 4576
rect -1914 4542 -1756 4576
rect -1722 4542 -1564 4576
rect -1530 4542 -1372 4576
rect -1338 4542 -1180 4576
rect -1146 4542 -988 4576
rect -954 4542 -938 4576
rect -1964 4526 -938 4542
rect -1898 4495 -1868 4526
rect -1802 4495 -1772 4526
rect -1706 4495 -1676 4526
rect -1610 4495 -1580 4526
rect -1514 4495 -1484 4526
rect -1418 4495 -1388 4526
rect -1322 4495 -1292 4526
rect -1226 4495 -1196 4526
rect -1130 4495 -1100 4526
rect -1034 4495 -1004 4526
rect -1898 4195 -1868 4221
rect -1802 4195 -1772 4221
rect -1706 4195 -1676 4221
rect -1610 4195 -1580 4221
rect -1514 4195 -1484 4221
rect -1418 4195 -1388 4221
rect -1322 4195 -1292 4221
rect -1226 4195 -1196 4221
rect -1130 4195 -1100 4221
rect -1034 4195 -1004 4221
rect 7036 4576 8062 4592
rect 7036 4542 7052 4576
rect 7086 4542 7244 4576
rect 7278 4542 7436 4576
rect 7470 4542 7628 4576
rect 7662 4542 7820 4576
rect 7854 4542 8012 4576
rect 8046 4542 8062 4576
rect 7036 4526 8062 4542
rect 7102 4495 7132 4526
rect 7198 4495 7228 4526
rect 7294 4495 7324 4526
rect 7390 4495 7420 4526
rect 7486 4495 7516 4526
rect 7582 4495 7612 4526
rect 7678 4495 7708 4526
rect 7774 4495 7804 4526
rect 7870 4495 7900 4526
rect 7966 4495 7996 4526
rect 7102 4195 7132 4221
rect 7198 4195 7228 4221
rect 7294 4195 7324 4221
rect 7390 4195 7420 4221
rect 7486 4195 7516 4221
rect 7582 4195 7612 4221
rect 7678 4195 7708 4221
rect 7774 4195 7804 4221
rect 7870 4195 7900 4221
rect 7966 4195 7996 4221
rect -1898 3916 -1868 3942
rect -1802 3916 -1772 3942
rect -1706 3916 -1676 3942
rect -1610 3916 -1580 3942
rect -1514 3916 -1484 3942
rect -1418 3916 -1388 3942
rect -1322 3916 -1292 3942
rect -1226 3916 -1196 3942
rect -1130 3916 -1100 3942
rect -1034 3916 -1004 3942
rect -1898 3788 -1868 3810
rect -1802 3788 -1772 3810
rect -1706 3788 -1676 3810
rect -1610 3788 -1580 3810
rect -1514 3788 -1484 3810
rect -1418 3788 -1388 3810
rect -1322 3788 -1292 3810
rect -1226 3788 -1196 3810
rect -1130 3788 -1100 3810
rect -1034 3788 -1004 3810
rect -1964 3769 -938 3788
rect -1964 3735 -1948 3769
rect -1914 3735 -1756 3769
rect -1722 3735 -1564 3769
rect -1530 3735 -1372 3769
rect -1338 3735 -1180 3769
rect -1146 3735 -988 3769
rect -954 3735 -938 3769
rect -1964 3722 -938 3735
rect 7102 3916 7132 3942
rect 7198 3916 7228 3942
rect 7294 3916 7324 3942
rect 7390 3916 7420 3942
rect 7486 3916 7516 3942
rect 7582 3916 7612 3942
rect 7678 3916 7708 3942
rect 7774 3916 7804 3942
rect 7870 3916 7900 3942
rect 7966 3916 7996 3942
rect 7102 3788 7132 3810
rect 7198 3788 7228 3810
rect 7294 3788 7324 3810
rect 7390 3788 7420 3810
rect 7486 3788 7516 3810
rect 7582 3788 7612 3810
rect 7678 3788 7708 3810
rect 7774 3788 7804 3810
rect 7870 3788 7900 3810
rect 7966 3788 7996 3810
rect 7036 3769 8062 3788
rect 7036 3735 7052 3769
rect 7086 3735 7244 3769
rect 7278 3735 7436 3769
rect 7470 3735 7628 3769
rect 7662 3735 7820 3769
rect 7854 3735 8012 3769
rect 8046 3735 8062 3769
rect 7036 3722 8062 3735
rect -1964 2776 -938 2792
rect -1964 2742 -1948 2776
rect -1914 2742 -1756 2776
rect -1722 2742 -1564 2776
rect -1530 2742 -1372 2776
rect -1338 2742 -1180 2776
rect -1146 2742 -988 2776
rect -954 2742 -938 2776
rect -1964 2726 -938 2742
rect -1898 2695 -1868 2726
rect -1802 2695 -1772 2726
rect -1706 2695 -1676 2726
rect -1610 2695 -1580 2726
rect -1514 2695 -1484 2726
rect -1418 2695 -1388 2726
rect -1322 2695 -1292 2726
rect -1226 2695 -1196 2726
rect -1130 2695 -1100 2726
rect -1034 2695 -1004 2726
rect -1898 2395 -1868 2421
rect -1802 2395 -1772 2421
rect -1706 2395 -1676 2421
rect -1610 2395 -1580 2421
rect -1514 2395 -1484 2421
rect -1418 2395 -1388 2421
rect -1322 2395 -1292 2421
rect -1226 2395 -1196 2421
rect -1130 2395 -1100 2421
rect -1034 2395 -1004 2421
rect 7036 2776 8062 2792
rect 7036 2742 7052 2776
rect 7086 2742 7244 2776
rect 7278 2742 7436 2776
rect 7470 2742 7628 2776
rect 7662 2742 7820 2776
rect 7854 2742 8012 2776
rect 8046 2742 8062 2776
rect 7036 2726 8062 2742
rect 7102 2695 7132 2726
rect 7198 2695 7228 2726
rect 7294 2695 7324 2726
rect 7390 2695 7420 2726
rect 7486 2695 7516 2726
rect 7582 2695 7612 2726
rect 7678 2695 7708 2726
rect 7774 2695 7804 2726
rect 7870 2695 7900 2726
rect 7966 2695 7996 2726
rect 7102 2395 7132 2421
rect 7198 2395 7228 2421
rect 7294 2395 7324 2421
rect 7390 2395 7420 2421
rect 7486 2395 7516 2421
rect 7582 2395 7612 2421
rect 7678 2395 7708 2421
rect 7774 2395 7804 2421
rect 7870 2395 7900 2421
rect 7966 2395 7996 2421
rect -1898 2116 -1868 2142
rect -1802 2116 -1772 2142
rect -1706 2116 -1676 2142
rect -1610 2116 -1580 2142
rect -1514 2116 -1484 2142
rect -1418 2116 -1388 2142
rect -1322 2116 -1292 2142
rect -1226 2116 -1196 2142
rect -1130 2116 -1100 2142
rect -1034 2116 -1004 2142
rect -1898 1988 -1868 2010
rect -1802 1988 -1772 2010
rect -1706 1988 -1676 2010
rect -1610 1988 -1580 2010
rect -1514 1988 -1484 2010
rect -1418 1988 -1388 2010
rect -1322 1988 -1292 2010
rect -1226 1988 -1196 2010
rect -1130 1988 -1100 2010
rect -1034 1988 -1004 2010
rect -1964 1969 -938 1988
rect -1964 1935 -1948 1969
rect -1914 1935 -1756 1969
rect -1722 1935 -1564 1969
rect -1530 1935 -1372 1969
rect -1338 1935 -1180 1969
rect -1146 1935 -988 1969
rect -954 1935 -938 1969
rect -1964 1922 -938 1935
rect 7102 2116 7132 2142
rect 7198 2116 7228 2142
rect 7294 2116 7324 2142
rect 7390 2116 7420 2142
rect 7486 2116 7516 2142
rect 7582 2116 7612 2142
rect 7678 2116 7708 2142
rect 7774 2116 7804 2142
rect 7870 2116 7900 2142
rect 7966 2116 7996 2142
rect 7102 1988 7132 2010
rect 7198 1988 7228 2010
rect 7294 1988 7324 2010
rect 7390 1988 7420 2010
rect 7486 1988 7516 2010
rect 7582 1988 7612 2010
rect 7678 1988 7708 2010
rect 7774 1988 7804 2010
rect 7870 1988 7900 2010
rect 7966 1988 7996 2010
rect 7036 1969 8062 1988
rect 7036 1935 7052 1969
rect 7086 1935 7244 1969
rect 7278 1935 7436 1969
rect 7470 1935 7628 1969
rect 7662 1935 7820 1969
rect 7854 1935 8012 1969
rect 8046 1935 8062 1969
rect 7036 1922 8062 1935
rect -1964 976 -938 992
rect -1964 942 -1948 976
rect -1914 942 -1756 976
rect -1722 942 -1564 976
rect -1530 942 -1372 976
rect -1338 942 -1180 976
rect -1146 942 -988 976
rect -954 942 -938 976
rect -1964 926 -938 942
rect -1898 895 -1868 926
rect -1802 895 -1772 926
rect -1706 895 -1676 926
rect -1610 895 -1580 926
rect -1514 895 -1484 926
rect -1418 895 -1388 926
rect -1322 895 -1292 926
rect -1226 895 -1196 926
rect -1130 895 -1100 926
rect -1034 895 -1004 926
rect -1898 595 -1868 621
rect -1802 595 -1772 621
rect -1706 595 -1676 621
rect -1610 595 -1580 621
rect -1514 595 -1484 621
rect -1418 595 -1388 621
rect -1322 595 -1292 621
rect -1226 595 -1196 621
rect -1130 595 -1100 621
rect -1034 595 -1004 621
rect 7036 976 8062 992
rect 7036 942 7052 976
rect 7086 942 7244 976
rect 7278 942 7436 976
rect 7470 942 7628 976
rect 7662 942 7820 976
rect 7854 942 8012 976
rect 8046 942 8062 976
rect 7036 926 8062 942
rect 7102 895 7132 926
rect 7198 895 7228 926
rect 7294 895 7324 926
rect 7390 895 7420 926
rect 7486 895 7516 926
rect 7582 895 7612 926
rect 7678 895 7708 926
rect 7774 895 7804 926
rect 7870 895 7900 926
rect 7966 895 7996 926
rect 7102 595 7132 621
rect 7198 595 7228 621
rect 7294 595 7324 621
rect 7390 595 7420 621
rect 7486 595 7516 621
rect 7582 595 7612 621
rect 7678 595 7708 621
rect 7774 595 7804 621
rect 7870 595 7900 621
rect 7966 595 7996 621
rect -1898 316 -1868 342
rect -1802 316 -1772 342
rect -1706 316 -1676 342
rect -1610 316 -1580 342
rect -1514 316 -1484 342
rect -1418 316 -1388 342
rect -1322 316 -1292 342
rect -1226 316 -1196 342
rect -1130 316 -1100 342
rect -1034 316 -1004 342
rect -1898 188 -1868 210
rect -1802 188 -1772 210
rect -1706 188 -1676 210
rect -1610 188 -1580 210
rect -1514 188 -1484 210
rect -1418 188 -1388 210
rect -1322 188 -1292 210
rect -1226 188 -1196 210
rect -1130 188 -1100 210
rect -1034 188 -1004 210
rect -1964 169 -938 188
rect -1964 135 -1948 169
rect -1914 135 -1756 169
rect -1722 135 -1564 169
rect -1530 135 -1372 169
rect -1338 135 -1180 169
rect -1146 135 -988 169
rect -954 135 -938 169
rect -1964 122 -938 135
rect 7102 316 7132 342
rect 7198 316 7228 342
rect 7294 316 7324 342
rect 7390 316 7420 342
rect 7486 316 7516 342
rect 7582 316 7612 342
rect 7678 316 7708 342
rect 7774 316 7804 342
rect 7870 316 7900 342
rect 7966 316 7996 342
rect 7102 188 7132 210
rect 7198 188 7228 210
rect 7294 188 7324 210
rect 7390 188 7420 210
rect 7486 188 7516 210
rect 7582 188 7612 210
rect 7678 188 7708 210
rect 7774 188 7804 210
rect 7870 188 7900 210
rect 7966 188 7996 210
rect 7036 169 8062 188
rect 7036 135 7052 169
rect 7086 135 7244 169
rect 7278 135 7436 169
rect 7470 135 7628 169
rect 7662 135 7820 169
rect 7854 135 8012 169
rect 8046 135 8062 169
rect 7036 122 8062 135
rect -1964 -824 -938 -808
rect -1964 -858 -1948 -824
rect -1914 -858 -1756 -824
rect -1722 -858 -1564 -824
rect -1530 -858 -1372 -824
rect -1338 -858 -1180 -824
rect -1146 -858 -988 -824
rect -954 -858 -938 -824
rect -1964 -874 -938 -858
rect -1898 -905 -1868 -874
rect -1802 -905 -1772 -874
rect -1706 -905 -1676 -874
rect -1610 -905 -1580 -874
rect -1514 -905 -1484 -874
rect -1418 -905 -1388 -874
rect -1322 -905 -1292 -874
rect -1226 -905 -1196 -874
rect -1130 -905 -1100 -874
rect -1034 -905 -1004 -874
rect -1898 -1205 -1868 -1179
rect -1802 -1205 -1772 -1179
rect -1706 -1205 -1676 -1179
rect -1610 -1205 -1580 -1179
rect -1514 -1205 -1484 -1179
rect -1418 -1205 -1388 -1179
rect -1322 -1205 -1292 -1179
rect -1226 -1205 -1196 -1179
rect -1130 -1205 -1100 -1179
rect -1034 -1205 -1004 -1179
rect 7036 -824 8062 -808
rect 7036 -858 7052 -824
rect 7086 -858 7244 -824
rect 7278 -858 7436 -824
rect 7470 -858 7628 -824
rect 7662 -858 7820 -824
rect 7854 -858 8012 -824
rect 8046 -858 8062 -824
rect 7036 -874 8062 -858
rect 7102 -905 7132 -874
rect 7198 -905 7228 -874
rect 7294 -905 7324 -874
rect 7390 -905 7420 -874
rect 7486 -905 7516 -874
rect 7582 -905 7612 -874
rect 7678 -905 7708 -874
rect 7774 -905 7804 -874
rect 7870 -905 7900 -874
rect 7966 -905 7996 -874
rect 7102 -1205 7132 -1179
rect 7198 -1205 7228 -1179
rect 7294 -1205 7324 -1179
rect 7390 -1205 7420 -1179
rect 7486 -1205 7516 -1179
rect 7582 -1205 7612 -1179
rect 7678 -1205 7708 -1179
rect 7774 -1205 7804 -1179
rect 7870 -1205 7900 -1179
rect 7966 -1205 7996 -1179
rect -1898 -1484 -1868 -1458
rect -1802 -1484 -1772 -1458
rect -1706 -1484 -1676 -1458
rect -1610 -1484 -1580 -1458
rect -1514 -1484 -1484 -1458
rect -1418 -1484 -1388 -1458
rect -1322 -1484 -1292 -1458
rect -1226 -1484 -1196 -1458
rect -1130 -1484 -1100 -1458
rect -1034 -1484 -1004 -1458
rect -1898 -1612 -1868 -1590
rect -1802 -1612 -1772 -1590
rect -1706 -1612 -1676 -1590
rect -1610 -1612 -1580 -1590
rect -1514 -1612 -1484 -1590
rect -1418 -1612 -1388 -1590
rect -1322 -1612 -1292 -1590
rect -1226 -1612 -1196 -1590
rect -1130 -1612 -1100 -1590
rect -1034 -1612 -1004 -1590
rect -1964 -1631 -938 -1612
rect -1964 -1665 -1948 -1631
rect -1914 -1665 -1756 -1631
rect -1722 -1665 -1564 -1631
rect -1530 -1665 -1372 -1631
rect -1338 -1665 -1180 -1631
rect -1146 -1665 -988 -1631
rect -954 -1665 -938 -1631
rect -1964 -1678 -938 -1665
rect 7102 -1484 7132 -1458
rect 7198 -1484 7228 -1458
rect 7294 -1484 7324 -1458
rect 7390 -1484 7420 -1458
rect 7486 -1484 7516 -1458
rect 7582 -1484 7612 -1458
rect 7678 -1484 7708 -1458
rect 7774 -1484 7804 -1458
rect 7870 -1484 7900 -1458
rect 7966 -1484 7996 -1458
rect 7102 -1612 7132 -1590
rect 7198 -1612 7228 -1590
rect 7294 -1612 7324 -1590
rect 7390 -1612 7420 -1590
rect 7486 -1612 7516 -1590
rect 7582 -1612 7612 -1590
rect 7678 -1612 7708 -1590
rect 7774 -1612 7804 -1590
rect 7870 -1612 7900 -1590
rect 7966 -1612 7996 -1590
rect 7036 -1631 8062 -1612
rect 7036 -1665 7052 -1631
rect 7086 -1665 7244 -1631
rect 7278 -1665 7436 -1631
rect 7470 -1665 7628 -1631
rect 7662 -1665 7820 -1631
rect 7854 -1665 8012 -1631
rect 8046 -1665 8062 -1631
rect 7036 -1678 8062 -1665
<< polycont >>
rect -1948 8142 -1914 8176
rect -1756 8142 -1722 8176
rect -1564 8142 -1530 8176
rect -1372 8142 -1338 8176
rect -1180 8142 -1146 8176
rect -988 8142 -954 8176
rect 7052 8142 7086 8176
rect 7244 8142 7278 8176
rect 7436 8142 7470 8176
rect 7628 8142 7662 8176
rect 7820 8142 7854 8176
rect 8012 8142 8046 8176
rect -1948 7335 -1914 7369
rect -1756 7335 -1722 7369
rect -1564 7335 -1530 7369
rect -1372 7335 -1338 7369
rect -1180 7335 -1146 7369
rect -988 7335 -954 7369
rect 7052 7335 7086 7369
rect 7244 7335 7278 7369
rect 7436 7335 7470 7369
rect 7628 7335 7662 7369
rect 7820 7335 7854 7369
rect 8012 7335 8046 7369
rect -1948 6342 -1914 6376
rect -1756 6342 -1722 6376
rect -1564 6342 -1530 6376
rect -1372 6342 -1338 6376
rect -1180 6342 -1146 6376
rect -988 6342 -954 6376
rect 7052 6342 7086 6376
rect 7244 6342 7278 6376
rect 7436 6342 7470 6376
rect 7628 6342 7662 6376
rect 7820 6342 7854 6376
rect 8012 6342 8046 6376
rect -1948 5535 -1914 5569
rect -1756 5535 -1722 5569
rect -1564 5535 -1530 5569
rect -1372 5535 -1338 5569
rect -1180 5535 -1146 5569
rect -988 5535 -954 5569
rect 7052 5535 7086 5569
rect 7244 5535 7278 5569
rect 7436 5535 7470 5569
rect 7628 5535 7662 5569
rect 7820 5535 7854 5569
rect 8012 5535 8046 5569
rect -1948 4542 -1914 4576
rect -1756 4542 -1722 4576
rect -1564 4542 -1530 4576
rect -1372 4542 -1338 4576
rect -1180 4542 -1146 4576
rect -988 4542 -954 4576
rect 7052 4542 7086 4576
rect 7244 4542 7278 4576
rect 7436 4542 7470 4576
rect 7628 4542 7662 4576
rect 7820 4542 7854 4576
rect 8012 4542 8046 4576
rect -1948 3735 -1914 3769
rect -1756 3735 -1722 3769
rect -1564 3735 -1530 3769
rect -1372 3735 -1338 3769
rect -1180 3735 -1146 3769
rect -988 3735 -954 3769
rect 7052 3735 7086 3769
rect 7244 3735 7278 3769
rect 7436 3735 7470 3769
rect 7628 3735 7662 3769
rect 7820 3735 7854 3769
rect 8012 3735 8046 3769
rect -1948 2742 -1914 2776
rect -1756 2742 -1722 2776
rect -1564 2742 -1530 2776
rect -1372 2742 -1338 2776
rect -1180 2742 -1146 2776
rect -988 2742 -954 2776
rect 7052 2742 7086 2776
rect 7244 2742 7278 2776
rect 7436 2742 7470 2776
rect 7628 2742 7662 2776
rect 7820 2742 7854 2776
rect 8012 2742 8046 2776
rect -1948 1935 -1914 1969
rect -1756 1935 -1722 1969
rect -1564 1935 -1530 1969
rect -1372 1935 -1338 1969
rect -1180 1935 -1146 1969
rect -988 1935 -954 1969
rect 7052 1935 7086 1969
rect 7244 1935 7278 1969
rect 7436 1935 7470 1969
rect 7628 1935 7662 1969
rect 7820 1935 7854 1969
rect 8012 1935 8046 1969
rect -1948 942 -1914 976
rect -1756 942 -1722 976
rect -1564 942 -1530 976
rect -1372 942 -1338 976
rect -1180 942 -1146 976
rect -988 942 -954 976
rect 7052 942 7086 976
rect 7244 942 7278 976
rect 7436 942 7470 976
rect 7628 942 7662 976
rect 7820 942 7854 976
rect 8012 942 8046 976
rect -1948 135 -1914 169
rect -1756 135 -1722 169
rect -1564 135 -1530 169
rect -1372 135 -1338 169
rect -1180 135 -1146 169
rect -988 135 -954 169
rect 7052 135 7086 169
rect 7244 135 7278 169
rect 7436 135 7470 169
rect 7628 135 7662 169
rect 7820 135 7854 169
rect 8012 135 8046 169
rect -1948 -858 -1914 -824
rect -1756 -858 -1722 -824
rect -1564 -858 -1530 -824
rect -1372 -858 -1338 -824
rect -1180 -858 -1146 -824
rect -988 -858 -954 -824
rect 7052 -858 7086 -824
rect 7244 -858 7278 -824
rect 7436 -858 7470 -824
rect 7628 -858 7662 -824
rect 7820 -858 7854 -824
rect 8012 -858 8046 -824
rect -1948 -1665 -1914 -1631
rect -1756 -1665 -1722 -1631
rect -1564 -1665 -1530 -1631
rect -1372 -1665 -1338 -1631
rect -1180 -1665 -1146 -1631
rect -988 -1665 -954 -1631
rect 7052 -1665 7086 -1631
rect 7244 -1665 7278 -1631
rect 7436 -1665 7470 -1631
rect 7628 -1665 7662 -1631
rect 7820 -1665 7854 -1631
rect 8012 -1665 8046 -1631
<< locali >>
rect -2062 8244 -1966 8278
rect -936 8244 -840 8278
rect -2062 8182 -2028 8244
rect -874 8182 -840 8244
rect -1964 8142 -1948 8176
rect -1914 8142 -1898 8176
rect -1772 8142 -1756 8176
rect -1722 8142 -1706 8176
rect -1580 8142 -1564 8176
rect -1530 8142 -1514 8176
rect -1388 8142 -1372 8176
rect -1338 8142 -1322 8176
rect -1196 8142 -1180 8176
rect -1146 8142 -1130 8176
rect -1004 8142 -988 8176
rect -954 8142 -938 8176
rect -1948 8083 -1914 8099
rect -1948 7817 -1914 7833
rect -1852 8083 -1818 8099
rect -1852 7817 -1818 7833
rect -1756 8083 -1722 8099
rect -1756 7817 -1722 7833
rect -1660 8083 -1626 8099
rect -1660 7817 -1626 7833
rect -1564 8083 -1530 8099
rect -1564 7817 -1530 7833
rect -1468 8083 -1434 8099
rect -1468 7817 -1434 7833
rect -1372 8083 -1338 8099
rect -1372 7817 -1338 7833
rect -1276 8083 -1242 8099
rect -1276 7817 -1242 7833
rect -1180 8083 -1146 8099
rect -1180 7817 -1146 7833
rect -1084 8083 -1050 8099
rect -1084 7817 -1050 7833
rect -988 8083 -954 8099
rect -988 7817 -954 7833
rect -2062 7734 -2028 7796
rect -874 7734 -840 7796
rect -2062 7700 -1966 7734
rect -936 7700 -840 7734
rect 6938 8244 7034 8278
rect 8064 8244 8160 8278
rect 6938 8182 6972 8244
rect 8126 8182 8160 8244
rect 7036 8142 7052 8176
rect 7086 8142 7102 8176
rect 7228 8142 7244 8176
rect 7278 8142 7294 8176
rect 7420 8142 7436 8176
rect 7470 8142 7486 8176
rect 7612 8142 7628 8176
rect 7662 8142 7678 8176
rect 7804 8142 7820 8176
rect 7854 8142 7870 8176
rect 7996 8142 8012 8176
rect 8046 8142 8062 8176
rect 7052 8083 7086 8099
rect 7052 7817 7086 7833
rect 7148 8083 7182 8099
rect 7148 7817 7182 7833
rect 7244 8083 7278 8099
rect 7244 7817 7278 7833
rect 7340 8083 7374 8099
rect 7340 7817 7374 7833
rect 7436 8083 7470 8099
rect 7436 7817 7470 7833
rect 7532 8083 7566 8099
rect 7532 7817 7566 7833
rect 7628 8083 7662 8099
rect 7628 7817 7662 7833
rect 7724 8083 7758 8099
rect 7724 7817 7758 7833
rect 7820 8083 7854 8099
rect 7820 7817 7854 7833
rect 7916 8083 7950 8099
rect 7916 7817 7950 7833
rect 8012 8083 8046 8099
rect 8012 7817 8046 7833
rect 6938 7734 6972 7796
rect 8126 7734 8160 7796
rect 6938 7700 7034 7734
rect 8064 7700 8160 7734
rect -2062 7594 -1966 7628
rect -936 7594 -840 7628
rect -2062 7532 -2028 7594
rect -874 7532 -840 7594
rect -1948 7504 -1914 7520
rect -1948 7406 -1914 7422
rect -1852 7504 -1818 7520
rect -1852 7406 -1818 7422
rect -1756 7504 -1722 7520
rect -1756 7406 -1722 7422
rect -1660 7504 -1626 7520
rect -1660 7406 -1626 7422
rect -1564 7504 -1530 7520
rect -1564 7406 -1530 7422
rect -1468 7504 -1434 7520
rect -1468 7406 -1434 7422
rect -1372 7504 -1338 7520
rect -1372 7406 -1338 7422
rect -1276 7504 -1242 7520
rect -1276 7406 -1242 7422
rect -1180 7504 -1146 7520
rect -1180 7406 -1146 7422
rect -1084 7504 -1050 7520
rect -1084 7406 -1050 7422
rect -988 7504 -954 7520
rect -988 7406 -954 7422
rect -1964 7335 -1948 7369
rect -1914 7335 -1898 7369
rect -1772 7335 -1756 7369
rect -1722 7335 -1706 7369
rect -1580 7335 -1564 7369
rect -1530 7335 -1514 7369
rect -1388 7335 -1372 7369
rect -1338 7335 -1322 7369
rect -1196 7335 -1180 7369
rect -1146 7335 -1130 7369
rect -1004 7335 -988 7369
rect -954 7335 -938 7369
rect -2062 7270 -2028 7332
rect -874 7270 -840 7332
rect -2062 7236 -1966 7270
rect -936 7236 -840 7270
rect 6938 7594 7034 7628
rect 8064 7594 8160 7628
rect 6938 7532 6972 7594
rect 8126 7532 8160 7594
rect 7052 7504 7086 7520
rect 7052 7406 7086 7422
rect 7148 7504 7182 7520
rect 7148 7406 7182 7422
rect 7244 7504 7278 7520
rect 7244 7406 7278 7422
rect 7340 7504 7374 7520
rect 7340 7406 7374 7422
rect 7436 7504 7470 7520
rect 7436 7406 7470 7422
rect 7532 7504 7566 7520
rect 7532 7406 7566 7422
rect 7628 7504 7662 7520
rect 7628 7406 7662 7422
rect 7724 7504 7758 7520
rect 7724 7406 7758 7422
rect 7820 7504 7854 7520
rect 7820 7406 7854 7422
rect 7916 7504 7950 7520
rect 7916 7406 7950 7422
rect 8012 7504 8046 7520
rect 8012 7406 8046 7422
rect 7036 7335 7052 7369
rect 7086 7335 7102 7369
rect 7228 7335 7244 7369
rect 7278 7335 7294 7369
rect 7420 7335 7436 7369
rect 7470 7335 7486 7369
rect 7612 7335 7628 7369
rect 7662 7335 7678 7369
rect 7804 7335 7820 7369
rect 7854 7335 7870 7369
rect 7996 7335 8012 7369
rect 8046 7335 8062 7369
rect 6938 7270 6972 7332
rect 8126 7270 8160 7332
rect 6938 7236 7034 7270
rect 8064 7236 8160 7270
rect -2062 6444 -1966 6478
rect -936 6444 -840 6478
rect -2062 6382 -2028 6444
rect -874 6382 -840 6444
rect -1964 6342 -1948 6376
rect -1914 6342 -1898 6376
rect -1772 6342 -1756 6376
rect -1722 6342 -1706 6376
rect -1580 6342 -1564 6376
rect -1530 6342 -1514 6376
rect -1388 6342 -1372 6376
rect -1338 6342 -1322 6376
rect -1196 6342 -1180 6376
rect -1146 6342 -1130 6376
rect -1004 6342 -988 6376
rect -954 6342 -938 6376
rect -1948 6283 -1914 6299
rect -1948 6017 -1914 6033
rect -1852 6283 -1818 6299
rect -1852 6017 -1818 6033
rect -1756 6283 -1722 6299
rect -1756 6017 -1722 6033
rect -1660 6283 -1626 6299
rect -1660 6017 -1626 6033
rect -1564 6283 -1530 6299
rect -1564 6017 -1530 6033
rect -1468 6283 -1434 6299
rect -1468 6017 -1434 6033
rect -1372 6283 -1338 6299
rect -1372 6017 -1338 6033
rect -1276 6283 -1242 6299
rect -1276 6017 -1242 6033
rect -1180 6283 -1146 6299
rect -1180 6017 -1146 6033
rect -1084 6283 -1050 6299
rect -1084 6017 -1050 6033
rect -988 6283 -954 6299
rect -988 6017 -954 6033
rect -2062 5934 -2028 5996
rect -874 5934 -840 5996
rect -2062 5900 -1966 5934
rect -936 5900 -840 5934
rect 6938 6444 7034 6478
rect 8064 6444 8160 6478
rect 6938 6382 6972 6444
rect 8126 6382 8160 6444
rect 7036 6342 7052 6376
rect 7086 6342 7102 6376
rect 7228 6342 7244 6376
rect 7278 6342 7294 6376
rect 7420 6342 7436 6376
rect 7470 6342 7486 6376
rect 7612 6342 7628 6376
rect 7662 6342 7678 6376
rect 7804 6342 7820 6376
rect 7854 6342 7870 6376
rect 7996 6342 8012 6376
rect 8046 6342 8062 6376
rect 7052 6283 7086 6299
rect 7052 6017 7086 6033
rect 7148 6283 7182 6299
rect 7148 6017 7182 6033
rect 7244 6283 7278 6299
rect 7244 6017 7278 6033
rect 7340 6283 7374 6299
rect 7340 6017 7374 6033
rect 7436 6283 7470 6299
rect 7436 6017 7470 6033
rect 7532 6283 7566 6299
rect 7532 6017 7566 6033
rect 7628 6283 7662 6299
rect 7628 6017 7662 6033
rect 7724 6283 7758 6299
rect 7724 6017 7758 6033
rect 7820 6283 7854 6299
rect 7820 6017 7854 6033
rect 7916 6283 7950 6299
rect 7916 6017 7950 6033
rect 8012 6283 8046 6299
rect 8012 6017 8046 6033
rect 6938 5934 6972 5996
rect 8126 5934 8160 5996
rect 6938 5900 7034 5934
rect 8064 5900 8160 5934
rect -2062 5794 -1966 5828
rect -936 5794 -840 5828
rect -2062 5732 -2028 5794
rect -874 5732 -840 5794
rect -1948 5704 -1914 5720
rect -1948 5606 -1914 5622
rect -1852 5704 -1818 5720
rect -1852 5606 -1818 5622
rect -1756 5704 -1722 5720
rect -1756 5606 -1722 5622
rect -1660 5704 -1626 5720
rect -1660 5606 -1626 5622
rect -1564 5704 -1530 5720
rect -1564 5606 -1530 5622
rect -1468 5704 -1434 5720
rect -1468 5606 -1434 5622
rect -1372 5704 -1338 5720
rect -1372 5606 -1338 5622
rect -1276 5704 -1242 5720
rect -1276 5606 -1242 5622
rect -1180 5704 -1146 5720
rect -1180 5606 -1146 5622
rect -1084 5704 -1050 5720
rect -1084 5606 -1050 5622
rect -988 5704 -954 5720
rect -988 5606 -954 5622
rect -1964 5535 -1948 5569
rect -1914 5535 -1898 5569
rect -1772 5535 -1756 5569
rect -1722 5535 -1706 5569
rect -1580 5535 -1564 5569
rect -1530 5535 -1514 5569
rect -1388 5535 -1372 5569
rect -1338 5535 -1322 5569
rect -1196 5535 -1180 5569
rect -1146 5535 -1130 5569
rect -1004 5535 -988 5569
rect -954 5535 -938 5569
rect -2062 5470 -2028 5532
rect -874 5470 -840 5532
rect -2062 5436 -1966 5470
rect -936 5436 -840 5470
rect 6938 5794 7034 5828
rect 8064 5794 8160 5828
rect 6938 5732 6972 5794
rect 8126 5732 8160 5794
rect 7052 5704 7086 5720
rect 7052 5606 7086 5622
rect 7148 5704 7182 5720
rect 7148 5606 7182 5622
rect 7244 5704 7278 5720
rect 7244 5606 7278 5622
rect 7340 5704 7374 5720
rect 7340 5606 7374 5622
rect 7436 5704 7470 5720
rect 7436 5606 7470 5622
rect 7532 5704 7566 5720
rect 7532 5606 7566 5622
rect 7628 5704 7662 5720
rect 7628 5606 7662 5622
rect 7724 5704 7758 5720
rect 7724 5606 7758 5622
rect 7820 5704 7854 5720
rect 7820 5606 7854 5622
rect 7916 5704 7950 5720
rect 7916 5606 7950 5622
rect 8012 5704 8046 5720
rect 8012 5606 8046 5622
rect 7036 5535 7052 5569
rect 7086 5535 7102 5569
rect 7228 5535 7244 5569
rect 7278 5535 7294 5569
rect 7420 5535 7436 5569
rect 7470 5535 7486 5569
rect 7612 5535 7628 5569
rect 7662 5535 7678 5569
rect 7804 5535 7820 5569
rect 7854 5535 7870 5569
rect 7996 5535 8012 5569
rect 8046 5535 8062 5569
rect 6938 5470 6972 5532
rect 8126 5470 8160 5532
rect 6938 5436 7034 5470
rect 8064 5436 8160 5470
rect -2062 4644 -1966 4678
rect -936 4644 -840 4678
rect -2062 4582 -2028 4644
rect -874 4582 -840 4644
rect -1964 4542 -1948 4576
rect -1914 4542 -1898 4576
rect -1772 4542 -1756 4576
rect -1722 4542 -1706 4576
rect -1580 4542 -1564 4576
rect -1530 4542 -1514 4576
rect -1388 4542 -1372 4576
rect -1338 4542 -1322 4576
rect -1196 4542 -1180 4576
rect -1146 4542 -1130 4576
rect -1004 4542 -988 4576
rect -954 4542 -938 4576
rect -1948 4483 -1914 4499
rect -1948 4217 -1914 4233
rect -1852 4483 -1818 4499
rect -1852 4217 -1818 4233
rect -1756 4483 -1722 4499
rect -1756 4217 -1722 4233
rect -1660 4483 -1626 4499
rect -1660 4217 -1626 4233
rect -1564 4483 -1530 4499
rect -1564 4217 -1530 4233
rect -1468 4483 -1434 4499
rect -1468 4217 -1434 4233
rect -1372 4483 -1338 4499
rect -1372 4217 -1338 4233
rect -1276 4483 -1242 4499
rect -1276 4217 -1242 4233
rect -1180 4483 -1146 4499
rect -1180 4217 -1146 4233
rect -1084 4483 -1050 4499
rect -1084 4217 -1050 4233
rect -988 4483 -954 4499
rect -988 4217 -954 4233
rect -2062 4134 -2028 4196
rect -874 4134 -840 4196
rect -2062 4100 -1966 4134
rect -936 4100 -840 4134
rect 6938 4644 7034 4678
rect 8064 4644 8160 4678
rect 6938 4582 6972 4644
rect 8126 4582 8160 4644
rect 7036 4542 7052 4576
rect 7086 4542 7102 4576
rect 7228 4542 7244 4576
rect 7278 4542 7294 4576
rect 7420 4542 7436 4576
rect 7470 4542 7486 4576
rect 7612 4542 7628 4576
rect 7662 4542 7678 4576
rect 7804 4542 7820 4576
rect 7854 4542 7870 4576
rect 7996 4542 8012 4576
rect 8046 4542 8062 4576
rect 7052 4483 7086 4499
rect 7052 4217 7086 4233
rect 7148 4483 7182 4499
rect 7148 4217 7182 4233
rect 7244 4483 7278 4499
rect 7244 4217 7278 4233
rect 7340 4483 7374 4499
rect 7340 4217 7374 4233
rect 7436 4483 7470 4499
rect 7436 4217 7470 4233
rect 7532 4483 7566 4499
rect 7532 4217 7566 4233
rect 7628 4483 7662 4499
rect 7628 4217 7662 4233
rect 7724 4483 7758 4499
rect 7724 4217 7758 4233
rect 7820 4483 7854 4499
rect 7820 4217 7854 4233
rect 7916 4483 7950 4499
rect 7916 4217 7950 4233
rect 8012 4483 8046 4499
rect 8012 4217 8046 4233
rect 6938 4134 6972 4196
rect 8126 4134 8160 4196
rect 6938 4100 7034 4134
rect 8064 4100 8160 4134
rect -2062 3994 -1966 4028
rect -936 3994 -840 4028
rect -2062 3932 -2028 3994
rect -874 3932 -840 3994
rect -1948 3904 -1914 3920
rect -1948 3806 -1914 3822
rect -1852 3904 -1818 3920
rect -1852 3806 -1818 3822
rect -1756 3904 -1722 3920
rect -1756 3806 -1722 3822
rect -1660 3904 -1626 3920
rect -1660 3806 -1626 3822
rect -1564 3904 -1530 3920
rect -1564 3806 -1530 3822
rect -1468 3904 -1434 3920
rect -1468 3806 -1434 3822
rect -1372 3904 -1338 3920
rect -1372 3806 -1338 3822
rect -1276 3904 -1242 3920
rect -1276 3806 -1242 3822
rect -1180 3904 -1146 3920
rect -1180 3806 -1146 3822
rect -1084 3904 -1050 3920
rect -1084 3806 -1050 3822
rect -988 3904 -954 3920
rect -988 3806 -954 3822
rect -1964 3735 -1948 3769
rect -1914 3735 -1898 3769
rect -1772 3735 -1756 3769
rect -1722 3735 -1706 3769
rect -1580 3735 -1564 3769
rect -1530 3735 -1514 3769
rect -1388 3735 -1372 3769
rect -1338 3735 -1322 3769
rect -1196 3735 -1180 3769
rect -1146 3735 -1130 3769
rect -1004 3735 -988 3769
rect -954 3735 -938 3769
rect -2062 3670 -2028 3732
rect -874 3670 -840 3732
rect -2062 3636 -1966 3670
rect -936 3636 -840 3670
rect 6938 3994 7034 4028
rect 8064 3994 8160 4028
rect 6938 3932 6972 3994
rect 8126 3932 8160 3994
rect 7052 3904 7086 3920
rect 7052 3806 7086 3822
rect 7148 3904 7182 3920
rect 7148 3806 7182 3822
rect 7244 3904 7278 3920
rect 7244 3806 7278 3822
rect 7340 3904 7374 3920
rect 7340 3806 7374 3822
rect 7436 3904 7470 3920
rect 7436 3806 7470 3822
rect 7532 3904 7566 3920
rect 7532 3806 7566 3822
rect 7628 3904 7662 3920
rect 7628 3806 7662 3822
rect 7724 3904 7758 3920
rect 7724 3806 7758 3822
rect 7820 3904 7854 3920
rect 7820 3806 7854 3822
rect 7916 3904 7950 3920
rect 7916 3806 7950 3822
rect 8012 3904 8046 3920
rect 8012 3806 8046 3822
rect 7036 3735 7052 3769
rect 7086 3735 7102 3769
rect 7228 3735 7244 3769
rect 7278 3735 7294 3769
rect 7420 3735 7436 3769
rect 7470 3735 7486 3769
rect 7612 3735 7628 3769
rect 7662 3735 7678 3769
rect 7804 3735 7820 3769
rect 7854 3735 7870 3769
rect 7996 3735 8012 3769
rect 8046 3735 8062 3769
rect 6938 3670 6972 3732
rect 8126 3670 8160 3732
rect 6938 3636 7034 3670
rect 8064 3636 8160 3670
rect -2062 2844 -1966 2878
rect -936 2844 -840 2878
rect -2062 2782 -2028 2844
rect -874 2782 -840 2844
rect -1964 2742 -1948 2776
rect -1914 2742 -1898 2776
rect -1772 2742 -1756 2776
rect -1722 2742 -1706 2776
rect -1580 2742 -1564 2776
rect -1530 2742 -1514 2776
rect -1388 2742 -1372 2776
rect -1338 2742 -1322 2776
rect -1196 2742 -1180 2776
rect -1146 2742 -1130 2776
rect -1004 2742 -988 2776
rect -954 2742 -938 2776
rect -1948 2683 -1914 2699
rect -1948 2417 -1914 2433
rect -1852 2683 -1818 2699
rect -1852 2417 -1818 2433
rect -1756 2683 -1722 2699
rect -1756 2417 -1722 2433
rect -1660 2683 -1626 2699
rect -1660 2417 -1626 2433
rect -1564 2683 -1530 2699
rect -1564 2417 -1530 2433
rect -1468 2683 -1434 2699
rect -1468 2417 -1434 2433
rect -1372 2683 -1338 2699
rect -1372 2417 -1338 2433
rect -1276 2683 -1242 2699
rect -1276 2417 -1242 2433
rect -1180 2683 -1146 2699
rect -1180 2417 -1146 2433
rect -1084 2683 -1050 2699
rect -1084 2417 -1050 2433
rect -988 2683 -954 2699
rect -988 2417 -954 2433
rect -2062 2334 -2028 2396
rect -874 2334 -840 2396
rect -2062 2300 -1966 2334
rect -936 2300 -840 2334
rect 6938 2844 7034 2878
rect 8064 2844 8160 2878
rect 6938 2782 6972 2844
rect 8126 2782 8160 2844
rect 7036 2742 7052 2776
rect 7086 2742 7102 2776
rect 7228 2742 7244 2776
rect 7278 2742 7294 2776
rect 7420 2742 7436 2776
rect 7470 2742 7486 2776
rect 7612 2742 7628 2776
rect 7662 2742 7678 2776
rect 7804 2742 7820 2776
rect 7854 2742 7870 2776
rect 7996 2742 8012 2776
rect 8046 2742 8062 2776
rect 7052 2683 7086 2699
rect 7052 2417 7086 2433
rect 7148 2683 7182 2699
rect 7148 2417 7182 2433
rect 7244 2683 7278 2699
rect 7244 2417 7278 2433
rect 7340 2683 7374 2699
rect 7340 2417 7374 2433
rect 7436 2683 7470 2699
rect 7436 2417 7470 2433
rect 7532 2683 7566 2699
rect 7532 2417 7566 2433
rect 7628 2683 7662 2699
rect 7628 2417 7662 2433
rect 7724 2683 7758 2699
rect 7724 2417 7758 2433
rect 7820 2683 7854 2699
rect 7820 2417 7854 2433
rect 7916 2683 7950 2699
rect 7916 2417 7950 2433
rect 8012 2683 8046 2699
rect 8012 2417 8046 2433
rect 6938 2334 6972 2396
rect 8126 2334 8160 2396
rect 6938 2300 7034 2334
rect 8064 2300 8160 2334
rect -2062 2194 -1966 2228
rect -936 2194 -840 2228
rect -2062 2132 -2028 2194
rect -874 2132 -840 2194
rect -1948 2104 -1914 2120
rect -1948 2006 -1914 2022
rect -1852 2104 -1818 2120
rect -1852 2006 -1818 2022
rect -1756 2104 -1722 2120
rect -1756 2006 -1722 2022
rect -1660 2104 -1626 2120
rect -1660 2006 -1626 2022
rect -1564 2104 -1530 2120
rect -1564 2006 -1530 2022
rect -1468 2104 -1434 2120
rect -1468 2006 -1434 2022
rect -1372 2104 -1338 2120
rect -1372 2006 -1338 2022
rect -1276 2104 -1242 2120
rect -1276 2006 -1242 2022
rect -1180 2104 -1146 2120
rect -1180 2006 -1146 2022
rect -1084 2104 -1050 2120
rect -1084 2006 -1050 2022
rect -988 2104 -954 2120
rect -988 2006 -954 2022
rect -1964 1935 -1948 1969
rect -1914 1935 -1898 1969
rect -1772 1935 -1756 1969
rect -1722 1935 -1706 1969
rect -1580 1935 -1564 1969
rect -1530 1935 -1514 1969
rect -1388 1935 -1372 1969
rect -1338 1935 -1322 1969
rect -1196 1935 -1180 1969
rect -1146 1935 -1130 1969
rect -1004 1935 -988 1969
rect -954 1935 -938 1969
rect -2062 1870 -2028 1932
rect -874 1870 -840 1932
rect -2062 1836 -1966 1870
rect -936 1836 -840 1870
rect 6938 2194 7034 2228
rect 8064 2194 8160 2228
rect 6938 2132 6972 2194
rect 8126 2132 8160 2194
rect 7052 2104 7086 2120
rect 7052 2006 7086 2022
rect 7148 2104 7182 2120
rect 7148 2006 7182 2022
rect 7244 2104 7278 2120
rect 7244 2006 7278 2022
rect 7340 2104 7374 2120
rect 7340 2006 7374 2022
rect 7436 2104 7470 2120
rect 7436 2006 7470 2022
rect 7532 2104 7566 2120
rect 7532 2006 7566 2022
rect 7628 2104 7662 2120
rect 7628 2006 7662 2022
rect 7724 2104 7758 2120
rect 7724 2006 7758 2022
rect 7820 2104 7854 2120
rect 7820 2006 7854 2022
rect 7916 2104 7950 2120
rect 7916 2006 7950 2022
rect 8012 2104 8046 2120
rect 8012 2006 8046 2022
rect 7036 1935 7052 1969
rect 7086 1935 7102 1969
rect 7228 1935 7244 1969
rect 7278 1935 7294 1969
rect 7420 1935 7436 1969
rect 7470 1935 7486 1969
rect 7612 1935 7628 1969
rect 7662 1935 7678 1969
rect 7804 1935 7820 1969
rect 7854 1935 7870 1969
rect 7996 1935 8012 1969
rect 8046 1935 8062 1969
rect 6938 1870 6972 1932
rect 8126 1870 8160 1932
rect 6938 1836 7034 1870
rect 8064 1836 8160 1870
rect -2062 1044 -1966 1078
rect -936 1044 -840 1078
rect -2062 982 -2028 1044
rect -874 982 -840 1044
rect -1964 942 -1948 976
rect -1914 942 -1898 976
rect -1772 942 -1756 976
rect -1722 942 -1706 976
rect -1580 942 -1564 976
rect -1530 942 -1514 976
rect -1388 942 -1372 976
rect -1338 942 -1322 976
rect -1196 942 -1180 976
rect -1146 942 -1130 976
rect -1004 942 -988 976
rect -954 942 -938 976
rect -1948 883 -1914 899
rect -1948 617 -1914 633
rect -1852 883 -1818 899
rect -1852 617 -1818 633
rect -1756 883 -1722 899
rect -1756 617 -1722 633
rect -1660 883 -1626 899
rect -1660 617 -1626 633
rect -1564 883 -1530 899
rect -1564 617 -1530 633
rect -1468 883 -1434 899
rect -1468 617 -1434 633
rect -1372 883 -1338 899
rect -1372 617 -1338 633
rect -1276 883 -1242 899
rect -1276 617 -1242 633
rect -1180 883 -1146 899
rect -1180 617 -1146 633
rect -1084 883 -1050 899
rect -1084 617 -1050 633
rect -988 883 -954 899
rect -988 617 -954 633
rect -2062 534 -2028 596
rect -874 534 -840 596
rect -2062 500 -1966 534
rect -936 500 -840 534
rect 6938 1044 7034 1078
rect 8064 1044 8160 1078
rect 6938 982 6972 1044
rect 8126 982 8160 1044
rect 7036 942 7052 976
rect 7086 942 7102 976
rect 7228 942 7244 976
rect 7278 942 7294 976
rect 7420 942 7436 976
rect 7470 942 7486 976
rect 7612 942 7628 976
rect 7662 942 7678 976
rect 7804 942 7820 976
rect 7854 942 7870 976
rect 7996 942 8012 976
rect 8046 942 8062 976
rect 7052 883 7086 899
rect 7052 617 7086 633
rect 7148 883 7182 899
rect 7148 617 7182 633
rect 7244 883 7278 899
rect 7244 617 7278 633
rect 7340 883 7374 899
rect 7340 617 7374 633
rect 7436 883 7470 899
rect 7436 617 7470 633
rect 7532 883 7566 899
rect 7532 617 7566 633
rect 7628 883 7662 899
rect 7628 617 7662 633
rect 7724 883 7758 899
rect 7724 617 7758 633
rect 7820 883 7854 899
rect 7820 617 7854 633
rect 7916 883 7950 899
rect 7916 617 7950 633
rect 8012 883 8046 899
rect 8012 617 8046 633
rect 6938 534 6972 596
rect 8126 534 8160 596
rect 6938 500 7034 534
rect 8064 500 8160 534
rect -2062 394 -1966 428
rect -936 394 -840 428
rect -2062 332 -2028 394
rect -874 332 -840 394
rect -1948 304 -1914 320
rect -1948 206 -1914 222
rect -1852 304 -1818 320
rect -1852 206 -1818 222
rect -1756 304 -1722 320
rect -1756 206 -1722 222
rect -1660 304 -1626 320
rect -1660 206 -1626 222
rect -1564 304 -1530 320
rect -1564 206 -1530 222
rect -1468 304 -1434 320
rect -1468 206 -1434 222
rect -1372 304 -1338 320
rect -1372 206 -1338 222
rect -1276 304 -1242 320
rect -1276 206 -1242 222
rect -1180 304 -1146 320
rect -1180 206 -1146 222
rect -1084 304 -1050 320
rect -1084 206 -1050 222
rect -988 304 -954 320
rect -988 206 -954 222
rect -1964 135 -1948 169
rect -1914 135 -1898 169
rect -1772 135 -1756 169
rect -1722 135 -1706 169
rect -1580 135 -1564 169
rect -1530 135 -1514 169
rect -1388 135 -1372 169
rect -1338 135 -1322 169
rect -1196 135 -1180 169
rect -1146 135 -1130 169
rect -1004 135 -988 169
rect -954 135 -938 169
rect -2062 70 -2028 132
rect -874 70 -840 132
rect -2062 36 -1966 70
rect -936 36 -840 70
rect 6938 394 7034 428
rect 8064 394 8160 428
rect 6938 332 6972 394
rect 8126 332 8160 394
rect 7052 304 7086 320
rect 7052 206 7086 222
rect 7148 304 7182 320
rect 7148 206 7182 222
rect 7244 304 7278 320
rect 7244 206 7278 222
rect 7340 304 7374 320
rect 7340 206 7374 222
rect 7436 304 7470 320
rect 7436 206 7470 222
rect 7532 304 7566 320
rect 7532 206 7566 222
rect 7628 304 7662 320
rect 7628 206 7662 222
rect 7724 304 7758 320
rect 7724 206 7758 222
rect 7820 304 7854 320
rect 7820 206 7854 222
rect 7916 304 7950 320
rect 7916 206 7950 222
rect 8012 304 8046 320
rect 8012 206 8046 222
rect 7036 135 7052 169
rect 7086 135 7102 169
rect 7228 135 7244 169
rect 7278 135 7294 169
rect 7420 135 7436 169
rect 7470 135 7486 169
rect 7612 135 7628 169
rect 7662 135 7678 169
rect 7804 135 7820 169
rect 7854 135 7870 169
rect 7996 135 8012 169
rect 8046 135 8062 169
rect 6938 70 6972 132
rect 8126 70 8160 132
rect 6938 36 7034 70
rect 8064 36 8160 70
rect -2062 -756 -1966 -722
rect -936 -756 -840 -722
rect -2062 -818 -2028 -756
rect -874 -818 -840 -756
rect -1964 -858 -1948 -824
rect -1914 -858 -1898 -824
rect -1772 -858 -1756 -824
rect -1722 -858 -1706 -824
rect -1580 -858 -1564 -824
rect -1530 -858 -1514 -824
rect -1388 -858 -1372 -824
rect -1338 -858 -1322 -824
rect -1196 -858 -1180 -824
rect -1146 -858 -1130 -824
rect -1004 -858 -988 -824
rect -954 -858 -938 -824
rect -1948 -917 -1914 -901
rect -1948 -1183 -1914 -1167
rect -1852 -917 -1818 -901
rect -1852 -1183 -1818 -1167
rect -1756 -917 -1722 -901
rect -1756 -1183 -1722 -1167
rect -1660 -917 -1626 -901
rect -1660 -1183 -1626 -1167
rect -1564 -917 -1530 -901
rect -1564 -1183 -1530 -1167
rect -1468 -917 -1434 -901
rect -1468 -1183 -1434 -1167
rect -1372 -917 -1338 -901
rect -1372 -1183 -1338 -1167
rect -1276 -917 -1242 -901
rect -1276 -1183 -1242 -1167
rect -1180 -917 -1146 -901
rect -1180 -1183 -1146 -1167
rect -1084 -917 -1050 -901
rect -1084 -1183 -1050 -1167
rect -988 -917 -954 -901
rect -988 -1183 -954 -1167
rect -2062 -1266 -2028 -1204
rect -874 -1266 -840 -1204
rect -2062 -1300 -1966 -1266
rect -936 -1300 -840 -1266
rect 6938 -756 7034 -722
rect 8064 -756 8160 -722
rect 6938 -818 6972 -756
rect 8126 -818 8160 -756
rect 7036 -858 7052 -824
rect 7086 -858 7102 -824
rect 7228 -858 7244 -824
rect 7278 -858 7294 -824
rect 7420 -858 7436 -824
rect 7470 -858 7486 -824
rect 7612 -858 7628 -824
rect 7662 -858 7678 -824
rect 7804 -858 7820 -824
rect 7854 -858 7870 -824
rect 7996 -858 8012 -824
rect 8046 -858 8062 -824
rect 7052 -917 7086 -901
rect 7052 -1183 7086 -1167
rect 7148 -917 7182 -901
rect 7148 -1183 7182 -1167
rect 7244 -917 7278 -901
rect 7244 -1183 7278 -1167
rect 7340 -917 7374 -901
rect 7340 -1183 7374 -1167
rect 7436 -917 7470 -901
rect 7436 -1183 7470 -1167
rect 7532 -917 7566 -901
rect 7532 -1183 7566 -1167
rect 7628 -917 7662 -901
rect 7628 -1183 7662 -1167
rect 7724 -917 7758 -901
rect 7724 -1183 7758 -1167
rect 7820 -917 7854 -901
rect 7820 -1183 7854 -1167
rect 7916 -917 7950 -901
rect 7916 -1183 7950 -1167
rect 8012 -917 8046 -901
rect 8012 -1183 8046 -1167
rect 6938 -1266 6972 -1204
rect 8126 -1266 8160 -1204
rect 6938 -1300 7034 -1266
rect 8064 -1300 8160 -1266
rect -2062 -1406 -1966 -1372
rect -936 -1406 -840 -1372
rect -2062 -1468 -2028 -1406
rect -874 -1468 -840 -1406
rect -1948 -1496 -1914 -1480
rect -1948 -1594 -1914 -1578
rect -1852 -1496 -1818 -1480
rect -1852 -1594 -1818 -1578
rect -1756 -1496 -1722 -1480
rect -1756 -1594 -1722 -1578
rect -1660 -1496 -1626 -1480
rect -1660 -1594 -1626 -1578
rect -1564 -1496 -1530 -1480
rect -1564 -1594 -1530 -1578
rect -1468 -1496 -1434 -1480
rect -1468 -1594 -1434 -1578
rect -1372 -1496 -1338 -1480
rect -1372 -1594 -1338 -1578
rect -1276 -1496 -1242 -1480
rect -1276 -1594 -1242 -1578
rect -1180 -1496 -1146 -1480
rect -1180 -1594 -1146 -1578
rect -1084 -1496 -1050 -1480
rect -1084 -1594 -1050 -1578
rect -988 -1496 -954 -1480
rect -988 -1594 -954 -1578
rect -1964 -1665 -1948 -1631
rect -1914 -1665 -1898 -1631
rect -1772 -1665 -1756 -1631
rect -1722 -1665 -1706 -1631
rect -1580 -1665 -1564 -1631
rect -1530 -1665 -1514 -1631
rect -1388 -1665 -1372 -1631
rect -1338 -1665 -1322 -1631
rect -1196 -1665 -1180 -1631
rect -1146 -1665 -1130 -1631
rect -1004 -1665 -988 -1631
rect -954 -1665 -938 -1631
rect -2062 -1730 -2028 -1668
rect -874 -1730 -840 -1668
rect -2062 -1764 -1966 -1730
rect -936 -1764 -840 -1730
rect 6938 -1406 7034 -1372
rect 8064 -1406 8160 -1372
rect 6938 -1468 6972 -1406
rect 8126 -1468 8160 -1406
rect 7052 -1496 7086 -1480
rect 7052 -1594 7086 -1578
rect 7148 -1496 7182 -1480
rect 7148 -1594 7182 -1578
rect 7244 -1496 7278 -1480
rect 7244 -1594 7278 -1578
rect 7340 -1496 7374 -1480
rect 7340 -1594 7374 -1578
rect 7436 -1496 7470 -1480
rect 7436 -1594 7470 -1578
rect 7532 -1496 7566 -1480
rect 7532 -1594 7566 -1578
rect 7628 -1496 7662 -1480
rect 7628 -1594 7662 -1578
rect 7724 -1496 7758 -1480
rect 7724 -1594 7758 -1578
rect 7820 -1496 7854 -1480
rect 7820 -1594 7854 -1578
rect 7916 -1496 7950 -1480
rect 7916 -1594 7950 -1578
rect 8012 -1496 8046 -1480
rect 8012 -1594 8046 -1578
rect 7036 -1665 7052 -1631
rect 7086 -1665 7102 -1631
rect 7228 -1665 7244 -1631
rect 7278 -1665 7294 -1631
rect 7420 -1665 7436 -1631
rect 7470 -1665 7486 -1631
rect 7612 -1665 7628 -1631
rect 7662 -1665 7678 -1631
rect 7804 -1665 7820 -1631
rect 7854 -1665 7870 -1631
rect 7996 -1665 8012 -1631
rect 8046 -1665 8062 -1631
rect 6938 -1730 6972 -1668
rect 8126 -1730 8160 -1668
rect 6938 -1764 7034 -1730
rect 8064 -1764 8160 -1730
<< viali >>
rect -2062 7796 -2028 8182
rect -1948 8142 -1914 8176
rect -1756 8142 -1722 8176
rect -1564 8142 -1530 8176
rect -1372 8142 -1338 8176
rect -1180 8142 -1146 8176
rect -988 8142 -954 8176
rect -1948 7833 -1914 8083
rect -1852 7833 -1818 8083
rect -1756 7833 -1722 8083
rect -1660 7833 -1626 8083
rect -1564 7833 -1530 8083
rect -1468 7833 -1434 8083
rect -1372 7833 -1338 8083
rect -1276 7833 -1242 8083
rect -1180 7833 -1146 8083
rect -1084 7833 -1050 8083
rect -988 7833 -954 8083
rect 6938 7796 6972 8182
rect 7052 8142 7086 8176
rect 7244 8142 7278 8176
rect 7436 8142 7470 8176
rect 7628 8142 7662 8176
rect 7820 8142 7854 8176
rect 8012 8142 8046 8176
rect 7052 7833 7086 8083
rect 7148 7833 7182 8083
rect 7244 7833 7278 8083
rect 7340 7833 7374 8083
rect 7436 7833 7470 8083
rect 7532 7833 7566 8083
rect 7628 7833 7662 8083
rect 7724 7833 7758 8083
rect 7820 7833 7854 8083
rect 7916 7833 7950 8083
rect 8012 7833 8046 8083
rect -2062 7332 -2028 7532
rect -1948 7422 -1914 7504
rect -1852 7422 -1818 7504
rect -1756 7422 -1722 7504
rect -1660 7422 -1626 7504
rect -1564 7422 -1530 7504
rect -1468 7422 -1434 7504
rect -1372 7422 -1338 7504
rect -1276 7422 -1242 7504
rect -1180 7422 -1146 7504
rect -1084 7422 -1050 7504
rect -988 7422 -954 7504
rect -1948 7335 -1914 7369
rect -1756 7335 -1722 7369
rect -1564 7335 -1530 7369
rect -1372 7335 -1338 7369
rect -1180 7335 -1146 7369
rect -988 7335 -954 7369
rect 6938 7332 6972 7532
rect 7052 7422 7086 7504
rect 7148 7422 7182 7504
rect 7244 7422 7278 7504
rect 7340 7422 7374 7504
rect 7436 7422 7470 7504
rect 7532 7422 7566 7504
rect 7628 7422 7662 7504
rect 7724 7422 7758 7504
rect 7820 7422 7854 7504
rect 7916 7422 7950 7504
rect 8012 7422 8046 7504
rect 7052 7335 7086 7369
rect 7244 7335 7278 7369
rect 7436 7335 7470 7369
rect 7628 7335 7662 7369
rect 7820 7335 7854 7369
rect 8012 7335 8046 7369
rect -2062 5996 -2028 6382
rect -1948 6342 -1914 6376
rect -1756 6342 -1722 6376
rect -1564 6342 -1530 6376
rect -1372 6342 -1338 6376
rect -1180 6342 -1146 6376
rect -988 6342 -954 6376
rect -1948 6033 -1914 6283
rect -1852 6033 -1818 6283
rect -1756 6033 -1722 6283
rect -1660 6033 -1626 6283
rect -1564 6033 -1530 6283
rect -1468 6033 -1434 6283
rect -1372 6033 -1338 6283
rect -1276 6033 -1242 6283
rect -1180 6033 -1146 6283
rect -1084 6033 -1050 6283
rect -988 6033 -954 6283
rect 6938 5996 6972 6382
rect 7052 6342 7086 6376
rect 7244 6342 7278 6376
rect 7436 6342 7470 6376
rect 7628 6342 7662 6376
rect 7820 6342 7854 6376
rect 8012 6342 8046 6376
rect 7052 6033 7086 6283
rect 7148 6033 7182 6283
rect 7244 6033 7278 6283
rect 7340 6033 7374 6283
rect 7436 6033 7470 6283
rect 7532 6033 7566 6283
rect 7628 6033 7662 6283
rect 7724 6033 7758 6283
rect 7820 6033 7854 6283
rect 7916 6033 7950 6283
rect 8012 6033 8046 6283
rect -2062 5532 -2028 5732
rect -1948 5622 -1914 5704
rect -1852 5622 -1818 5704
rect -1756 5622 -1722 5704
rect -1660 5622 -1626 5704
rect -1564 5622 -1530 5704
rect -1468 5622 -1434 5704
rect -1372 5622 -1338 5704
rect -1276 5622 -1242 5704
rect -1180 5622 -1146 5704
rect -1084 5622 -1050 5704
rect -988 5622 -954 5704
rect -1948 5535 -1914 5569
rect -1756 5535 -1722 5569
rect -1564 5535 -1530 5569
rect -1372 5535 -1338 5569
rect -1180 5535 -1146 5569
rect -988 5535 -954 5569
rect 6938 5532 6972 5732
rect 7052 5622 7086 5704
rect 7148 5622 7182 5704
rect 7244 5622 7278 5704
rect 7340 5622 7374 5704
rect 7436 5622 7470 5704
rect 7532 5622 7566 5704
rect 7628 5622 7662 5704
rect 7724 5622 7758 5704
rect 7820 5622 7854 5704
rect 7916 5622 7950 5704
rect 8012 5622 8046 5704
rect 7052 5535 7086 5569
rect 7244 5535 7278 5569
rect 7436 5535 7470 5569
rect 7628 5535 7662 5569
rect 7820 5535 7854 5569
rect 8012 5535 8046 5569
rect -2062 4196 -2028 4582
rect -1948 4542 -1914 4576
rect -1756 4542 -1722 4576
rect -1564 4542 -1530 4576
rect -1372 4542 -1338 4576
rect -1180 4542 -1146 4576
rect -988 4542 -954 4576
rect -1948 4233 -1914 4483
rect -1852 4233 -1818 4483
rect -1756 4233 -1722 4483
rect -1660 4233 -1626 4483
rect -1564 4233 -1530 4483
rect -1468 4233 -1434 4483
rect -1372 4233 -1338 4483
rect -1276 4233 -1242 4483
rect -1180 4233 -1146 4483
rect -1084 4233 -1050 4483
rect -988 4233 -954 4483
rect 6938 4196 6972 4582
rect 7052 4542 7086 4576
rect 7244 4542 7278 4576
rect 7436 4542 7470 4576
rect 7628 4542 7662 4576
rect 7820 4542 7854 4576
rect 8012 4542 8046 4576
rect 7052 4233 7086 4483
rect 7148 4233 7182 4483
rect 7244 4233 7278 4483
rect 7340 4233 7374 4483
rect 7436 4233 7470 4483
rect 7532 4233 7566 4483
rect 7628 4233 7662 4483
rect 7724 4233 7758 4483
rect 7820 4233 7854 4483
rect 7916 4233 7950 4483
rect 8012 4233 8046 4483
rect -2062 3732 -2028 3932
rect -1948 3822 -1914 3904
rect -1852 3822 -1818 3904
rect -1756 3822 -1722 3904
rect -1660 3822 -1626 3904
rect -1564 3822 -1530 3904
rect -1468 3822 -1434 3904
rect -1372 3822 -1338 3904
rect -1276 3822 -1242 3904
rect -1180 3822 -1146 3904
rect -1084 3822 -1050 3904
rect -988 3822 -954 3904
rect -1948 3735 -1914 3769
rect -1756 3735 -1722 3769
rect -1564 3735 -1530 3769
rect -1372 3735 -1338 3769
rect -1180 3735 -1146 3769
rect -988 3735 -954 3769
rect 6938 3732 6972 3932
rect 7052 3822 7086 3904
rect 7148 3822 7182 3904
rect 7244 3822 7278 3904
rect 7340 3822 7374 3904
rect 7436 3822 7470 3904
rect 7532 3822 7566 3904
rect 7628 3822 7662 3904
rect 7724 3822 7758 3904
rect 7820 3822 7854 3904
rect 7916 3822 7950 3904
rect 8012 3822 8046 3904
rect 7052 3735 7086 3769
rect 7244 3735 7278 3769
rect 7436 3735 7470 3769
rect 7628 3735 7662 3769
rect 7820 3735 7854 3769
rect 8012 3735 8046 3769
rect -2062 2396 -2028 2782
rect -1948 2742 -1914 2776
rect -1756 2742 -1722 2776
rect -1564 2742 -1530 2776
rect -1372 2742 -1338 2776
rect -1180 2742 -1146 2776
rect -988 2742 -954 2776
rect -1948 2433 -1914 2683
rect -1852 2433 -1818 2683
rect -1756 2433 -1722 2683
rect -1660 2433 -1626 2683
rect -1564 2433 -1530 2683
rect -1468 2433 -1434 2683
rect -1372 2433 -1338 2683
rect -1276 2433 -1242 2683
rect -1180 2433 -1146 2683
rect -1084 2433 -1050 2683
rect -988 2433 -954 2683
rect 6938 2396 6972 2782
rect 7052 2742 7086 2776
rect 7244 2742 7278 2776
rect 7436 2742 7470 2776
rect 7628 2742 7662 2776
rect 7820 2742 7854 2776
rect 8012 2742 8046 2776
rect 7052 2433 7086 2683
rect 7148 2433 7182 2683
rect 7244 2433 7278 2683
rect 7340 2433 7374 2683
rect 7436 2433 7470 2683
rect 7532 2433 7566 2683
rect 7628 2433 7662 2683
rect 7724 2433 7758 2683
rect 7820 2433 7854 2683
rect 7916 2433 7950 2683
rect 8012 2433 8046 2683
rect -2062 1932 -2028 2132
rect -1948 2022 -1914 2104
rect -1852 2022 -1818 2104
rect -1756 2022 -1722 2104
rect -1660 2022 -1626 2104
rect -1564 2022 -1530 2104
rect -1468 2022 -1434 2104
rect -1372 2022 -1338 2104
rect -1276 2022 -1242 2104
rect -1180 2022 -1146 2104
rect -1084 2022 -1050 2104
rect -988 2022 -954 2104
rect -1948 1935 -1914 1969
rect -1756 1935 -1722 1969
rect -1564 1935 -1530 1969
rect -1372 1935 -1338 1969
rect -1180 1935 -1146 1969
rect -988 1935 -954 1969
rect 6938 1932 6972 2132
rect 7052 2022 7086 2104
rect 7148 2022 7182 2104
rect 7244 2022 7278 2104
rect 7340 2022 7374 2104
rect 7436 2022 7470 2104
rect 7532 2022 7566 2104
rect 7628 2022 7662 2104
rect 7724 2022 7758 2104
rect 7820 2022 7854 2104
rect 7916 2022 7950 2104
rect 8012 2022 8046 2104
rect 7052 1935 7086 1969
rect 7244 1935 7278 1969
rect 7436 1935 7470 1969
rect 7628 1935 7662 1969
rect 7820 1935 7854 1969
rect 8012 1935 8046 1969
rect -2062 596 -2028 982
rect -1948 942 -1914 976
rect -1756 942 -1722 976
rect -1564 942 -1530 976
rect -1372 942 -1338 976
rect -1180 942 -1146 976
rect -988 942 -954 976
rect -1948 633 -1914 883
rect -1852 633 -1818 883
rect -1756 633 -1722 883
rect -1660 633 -1626 883
rect -1564 633 -1530 883
rect -1468 633 -1434 883
rect -1372 633 -1338 883
rect -1276 633 -1242 883
rect -1180 633 -1146 883
rect -1084 633 -1050 883
rect -988 633 -954 883
rect 6938 596 6972 982
rect 7052 942 7086 976
rect 7244 942 7278 976
rect 7436 942 7470 976
rect 7628 942 7662 976
rect 7820 942 7854 976
rect 8012 942 8046 976
rect 7052 633 7086 883
rect 7148 633 7182 883
rect 7244 633 7278 883
rect 7340 633 7374 883
rect 7436 633 7470 883
rect 7532 633 7566 883
rect 7628 633 7662 883
rect 7724 633 7758 883
rect 7820 633 7854 883
rect 7916 633 7950 883
rect 8012 633 8046 883
rect -2062 132 -2028 332
rect -1948 222 -1914 304
rect -1852 222 -1818 304
rect -1756 222 -1722 304
rect -1660 222 -1626 304
rect -1564 222 -1530 304
rect -1468 222 -1434 304
rect -1372 222 -1338 304
rect -1276 222 -1242 304
rect -1180 222 -1146 304
rect -1084 222 -1050 304
rect -988 222 -954 304
rect -1948 135 -1914 169
rect -1756 135 -1722 169
rect -1564 135 -1530 169
rect -1372 135 -1338 169
rect -1180 135 -1146 169
rect -988 135 -954 169
rect 6938 132 6972 332
rect 7052 222 7086 304
rect 7148 222 7182 304
rect 7244 222 7278 304
rect 7340 222 7374 304
rect 7436 222 7470 304
rect 7532 222 7566 304
rect 7628 222 7662 304
rect 7724 222 7758 304
rect 7820 222 7854 304
rect 7916 222 7950 304
rect 8012 222 8046 304
rect 7052 135 7086 169
rect 7244 135 7278 169
rect 7436 135 7470 169
rect 7628 135 7662 169
rect 7820 135 7854 169
rect 8012 135 8046 169
rect -2062 -1204 -2028 -818
rect -1948 -858 -1914 -824
rect -1756 -858 -1722 -824
rect -1564 -858 -1530 -824
rect -1372 -858 -1338 -824
rect -1180 -858 -1146 -824
rect -988 -858 -954 -824
rect -1948 -1167 -1914 -917
rect -1852 -1167 -1818 -917
rect -1756 -1167 -1722 -917
rect -1660 -1167 -1626 -917
rect -1564 -1167 -1530 -917
rect -1468 -1167 -1434 -917
rect -1372 -1167 -1338 -917
rect -1276 -1167 -1242 -917
rect -1180 -1167 -1146 -917
rect -1084 -1167 -1050 -917
rect -988 -1167 -954 -917
rect 6938 -1204 6972 -818
rect 7052 -858 7086 -824
rect 7244 -858 7278 -824
rect 7436 -858 7470 -824
rect 7628 -858 7662 -824
rect 7820 -858 7854 -824
rect 8012 -858 8046 -824
rect 7052 -1167 7086 -917
rect 7148 -1167 7182 -917
rect 7244 -1167 7278 -917
rect 7340 -1167 7374 -917
rect 7436 -1167 7470 -917
rect 7532 -1167 7566 -917
rect 7628 -1167 7662 -917
rect 7724 -1167 7758 -917
rect 7820 -1167 7854 -917
rect 7916 -1167 7950 -917
rect 8012 -1167 8046 -917
rect -2062 -1668 -2028 -1468
rect -1948 -1578 -1914 -1496
rect -1852 -1578 -1818 -1496
rect -1756 -1578 -1722 -1496
rect -1660 -1578 -1626 -1496
rect -1564 -1578 -1530 -1496
rect -1468 -1578 -1434 -1496
rect -1372 -1578 -1338 -1496
rect -1276 -1578 -1242 -1496
rect -1180 -1578 -1146 -1496
rect -1084 -1578 -1050 -1496
rect -988 -1578 -954 -1496
rect -1948 -1665 -1914 -1631
rect -1756 -1665 -1722 -1631
rect -1564 -1665 -1530 -1631
rect -1372 -1665 -1338 -1631
rect -1180 -1665 -1146 -1631
rect -988 -1665 -954 -1631
rect 6938 -1668 6972 -1468
rect 7052 -1578 7086 -1496
rect 7148 -1578 7182 -1496
rect 7244 -1578 7278 -1496
rect 7340 -1578 7374 -1496
rect 7436 -1578 7470 -1496
rect 7532 -1578 7566 -1496
rect 7628 -1578 7662 -1496
rect 7724 -1578 7758 -1496
rect 7820 -1578 7854 -1496
rect 7916 -1578 7950 -1496
rect 8012 -1578 8046 -1496
rect 7052 -1665 7086 -1631
rect 7244 -1665 7278 -1631
rect 7436 -1665 7470 -1631
rect 7628 -1665 7662 -1631
rect 7820 -1665 7854 -1631
rect 8012 -1665 8046 -1631
<< metal1 >>
rect -2068 8182 -2022 8360
rect -1852 8244 -770 8278
rect -2068 7796 -2062 8182
rect -2028 7796 -2022 8182
rect -1967 8134 -1957 8186
rect -1905 8134 -1895 8186
rect -1852 8095 -1818 8244
rect -1775 8134 -1765 8186
rect -1713 8134 -1703 8186
rect -1660 8095 -1626 8244
rect -1583 8134 -1573 8186
rect -1521 8134 -1511 8186
rect -1468 8095 -1434 8244
rect -1391 8134 -1381 8186
rect -1329 8134 -1319 8186
rect -1276 8095 -1242 8244
rect -1200 8134 -1190 8186
rect -1138 8134 -1128 8186
rect -1084 8095 -1050 8244
rect -1007 8134 -997 8186
rect -945 8134 -935 8186
rect -1954 8083 -1908 8095
rect -1954 7833 -1948 8083
rect -1914 7833 -1908 8083
rect -1954 7821 -1908 7833
rect -1858 8083 -1812 8095
rect -1858 7833 -1852 8083
rect -1818 7833 -1812 8083
rect -1858 7821 -1812 7833
rect -1762 8083 -1716 8095
rect -1762 7833 -1756 8083
rect -1722 7833 -1716 8083
rect -1762 7821 -1716 7833
rect -1666 8083 -1620 8095
rect -1666 7833 -1660 8083
rect -1626 7833 -1620 8083
rect -1666 7821 -1620 7833
rect -1570 8083 -1524 8095
rect -1570 7833 -1564 8083
rect -1530 7833 -1524 8083
rect -1570 7821 -1524 7833
rect -1474 8083 -1428 8095
rect -1474 7833 -1468 8083
rect -1434 7833 -1428 8083
rect -1474 7821 -1428 7833
rect -1378 8083 -1332 8095
rect -1378 7833 -1372 8083
rect -1338 7833 -1332 8083
rect -1378 7821 -1332 7833
rect -1282 8083 -1236 8095
rect -1282 7833 -1276 8083
rect -1242 7833 -1236 8083
rect -1282 7821 -1236 7833
rect -1186 8083 -1140 8095
rect -1186 7833 -1180 8083
rect -1146 7833 -1140 8083
rect -1186 7821 -1140 7833
rect -1090 8083 -1044 8095
rect -1090 7833 -1084 8083
rect -1050 7833 -1044 8083
rect -1090 7821 -1044 7833
rect -994 8083 -948 8095
rect -994 7833 -988 8083
rect -954 7833 -948 8083
rect -994 7821 -948 7833
rect -2068 7784 -2022 7796
rect -1948 7681 -1914 7821
rect -1756 7681 -1722 7821
rect -1564 7681 -1530 7821
rect -1372 7681 -1338 7821
rect -1180 7681 -1146 7821
rect -988 7695 -954 7821
rect -1032 7681 -1022 7695
rect -3494 7647 -1022 7681
rect -3494 -1319 -3419 7647
rect -2068 7532 -2022 7544
rect -2068 7332 -2062 7532
rect -2028 7332 -2022 7532
rect -1948 7516 -1914 7647
rect -1756 7516 -1722 7647
rect -1564 7516 -1530 7647
rect -1372 7516 -1338 7647
rect -1180 7516 -1146 7647
rect -1032 7631 -1022 7647
rect -958 7631 -948 7695
rect -804 7681 -770 8244
rect -730 8134 -720 8186
rect -668 8134 -641 8186
rect 6932 8182 6978 8360
rect 7148 8244 8230 8278
rect 6932 7796 6938 8182
rect 6972 7796 6978 8182
rect 7033 8134 7043 8186
rect 7095 8134 7105 8186
rect 7148 8095 7182 8244
rect 7225 8134 7235 8186
rect 7287 8134 7297 8186
rect 7340 8095 7374 8244
rect 7417 8134 7427 8186
rect 7479 8134 7489 8186
rect 7532 8095 7566 8244
rect 7609 8134 7619 8186
rect 7671 8134 7681 8186
rect 7724 8095 7758 8244
rect 7800 8134 7810 8186
rect 7862 8134 7872 8186
rect 7916 8095 7950 8244
rect 7993 8134 8003 8186
rect 8055 8134 8065 8186
rect 7046 8083 7092 8095
rect 7046 7833 7052 8083
rect 7086 7833 7092 8083
rect 7046 7821 7092 7833
rect 7142 8083 7188 8095
rect 7142 7833 7148 8083
rect 7182 7833 7188 8083
rect 7142 7821 7188 7833
rect 7238 8083 7284 8095
rect 7238 7833 7244 8083
rect 7278 7833 7284 8083
rect 7238 7821 7284 7833
rect 7334 8083 7380 8095
rect 7334 7833 7340 8083
rect 7374 7833 7380 8083
rect 7334 7821 7380 7833
rect 7430 8083 7476 8095
rect 7430 7833 7436 8083
rect 7470 7833 7476 8083
rect 7430 7821 7476 7833
rect 7526 8083 7572 8095
rect 7526 7833 7532 8083
rect 7566 7833 7572 8083
rect 7526 7821 7572 7833
rect 7622 8083 7668 8095
rect 7622 7833 7628 8083
rect 7662 7833 7668 8083
rect 7622 7821 7668 7833
rect 7718 8083 7764 8095
rect 7718 7833 7724 8083
rect 7758 7833 7764 8083
rect 7718 7821 7764 7833
rect 7814 8083 7860 8095
rect 7814 7833 7820 8083
rect 7854 7833 7860 8083
rect 7814 7821 7860 7833
rect 7910 8083 7956 8095
rect 7910 7833 7916 8083
rect 7950 7833 7956 8083
rect 7910 7821 7956 7833
rect 8006 8083 8052 8095
rect 8006 7833 8012 8083
rect 8046 7833 8052 8083
rect 8006 7821 8052 7833
rect 6932 7784 6978 7796
rect -485 7681 2411 7697
rect -804 7647 2411 7681
rect -988 7516 -954 7631
rect -1954 7504 -1908 7516
rect -1954 7422 -1948 7504
rect -1914 7422 -1908 7504
rect -1954 7410 -1908 7422
rect -1858 7504 -1812 7516
rect -1858 7422 -1852 7504
rect -1818 7422 -1812 7504
rect -1858 7410 -1812 7422
rect -1762 7504 -1716 7516
rect -1762 7422 -1756 7504
rect -1722 7422 -1716 7504
rect -1762 7410 -1716 7422
rect -1666 7504 -1620 7516
rect -1666 7422 -1660 7504
rect -1626 7422 -1620 7504
rect -1666 7410 -1620 7422
rect -1570 7504 -1524 7516
rect -1570 7422 -1564 7504
rect -1530 7422 -1524 7504
rect -1570 7410 -1524 7422
rect -1474 7504 -1428 7516
rect -1474 7422 -1468 7504
rect -1434 7422 -1428 7504
rect -1474 7410 -1428 7422
rect -1378 7504 -1332 7516
rect -1378 7422 -1372 7504
rect -1338 7422 -1332 7504
rect -1378 7410 -1332 7422
rect -1282 7504 -1236 7516
rect -1282 7422 -1276 7504
rect -1242 7422 -1236 7504
rect -1282 7410 -1236 7422
rect -1186 7504 -1140 7516
rect -1186 7422 -1180 7504
rect -1146 7422 -1140 7504
rect -1186 7410 -1140 7422
rect -1090 7504 -1044 7516
rect -1090 7422 -1084 7504
rect -1050 7422 -1044 7504
rect -1090 7410 -1044 7422
rect -994 7504 -948 7516
rect -994 7422 -988 7504
rect -954 7422 -948 7504
rect -994 7410 -948 7422
rect -1964 7378 -1898 7382
rect -2068 7160 -2022 7332
rect -1967 7326 -1957 7378
rect -1905 7326 -1895 7378
rect -1964 7322 -1898 7326
rect -1852 7270 -1818 7410
rect -1772 7378 -1706 7382
rect -1775 7326 -1765 7378
rect -1713 7326 -1703 7378
rect -1772 7322 -1706 7326
rect -1660 7270 -1626 7410
rect -1580 7379 -1514 7382
rect -1582 7327 -1572 7379
rect -1520 7327 -1510 7379
rect -1580 7322 -1514 7327
rect -1468 7270 -1434 7410
rect -1388 7379 -1322 7382
rect -1390 7327 -1380 7379
rect -1328 7327 -1318 7379
rect -1388 7322 -1322 7327
rect -1276 7270 -1242 7410
rect -1196 7379 -1130 7382
rect -1198 7327 -1188 7379
rect -1136 7327 -1126 7379
rect -1196 7322 -1130 7327
rect -1084 7270 -1050 7410
rect -1004 7379 -938 7382
rect -1007 7327 -997 7379
rect -945 7327 -935 7379
rect -1004 7322 -938 7327
rect -804 7270 -770 7647
rect -485 7633 2411 7647
rect 6681 7633 6691 7697
rect 6755 7681 6765 7697
rect 7052 7681 7086 7821
rect 7244 7681 7278 7821
rect 7436 7681 7470 7821
rect 7628 7681 7662 7821
rect 7820 7681 7854 7821
rect 8012 7681 8046 7821
rect 6755 7647 8046 7681
rect 6755 7633 6765 7647
rect -730 7327 -720 7379
rect -668 7327 -641 7379
rect -1852 7236 -770 7270
rect -2068 6382 -2022 6560
rect -1852 6444 -770 6478
rect -2068 5996 -2062 6382
rect -2028 5996 -2022 6382
rect -1967 6334 -1957 6386
rect -1905 6334 -1895 6386
rect -1852 6295 -1818 6444
rect -1775 6334 -1765 6386
rect -1713 6334 -1703 6386
rect -1660 6295 -1626 6444
rect -1583 6334 -1573 6386
rect -1521 6334 -1511 6386
rect -1468 6295 -1434 6444
rect -1391 6334 -1381 6386
rect -1329 6334 -1319 6386
rect -1276 6295 -1242 6444
rect -1200 6334 -1190 6386
rect -1138 6334 -1128 6386
rect -1084 6295 -1050 6444
rect -1007 6334 -997 6386
rect -945 6334 -935 6386
rect -1954 6283 -1908 6295
rect -1954 6033 -1948 6283
rect -1914 6033 -1908 6283
rect -1954 6021 -1908 6033
rect -1858 6283 -1812 6295
rect -1858 6033 -1852 6283
rect -1818 6033 -1812 6283
rect -1858 6021 -1812 6033
rect -1762 6283 -1716 6295
rect -1762 6033 -1756 6283
rect -1722 6033 -1716 6283
rect -1762 6021 -1716 6033
rect -1666 6283 -1620 6295
rect -1666 6033 -1660 6283
rect -1626 6033 -1620 6283
rect -1666 6021 -1620 6033
rect -1570 6283 -1524 6295
rect -1570 6033 -1564 6283
rect -1530 6033 -1524 6283
rect -1570 6021 -1524 6033
rect -1474 6283 -1428 6295
rect -1474 6033 -1468 6283
rect -1434 6033 -1428 6283
rect -1474 6021 -1428 6033
rect -1378 6283 -1332 6295
rect -1378 6033 -1372 6283
rect -1338 6033 -1332 6283
rect -1378 6021 -1332 6033
rect -1282 6283 -1236 6295
rect -1282 6033 -1276 6283
rect -1242 6033 -1236 6283
rect -1282 6021 -1236 6033
rect -1186 6283 -1140 6295
rect -1186 6033 -1180 6283
rect -1146 6033 -1140 6283
rect -1186 6021 -1140 6033
rect -1090 6283 -1044 6295
rect -1090 6033 -1084 6283
rect -1050 6033 -1044 6283
rect -1090 6021 -1044 6033
rect -994 6283 -948 6295
rect -994 6033 -988 6283
rect -954 6033 -948 6283
rect -994 6021 -948 6033
rect -2068 5984 -2022 5996
rect -1948 5881 -1914 6021
rect -1756 5881 -1722 6021
rect -1564 5881 -1530 6021
rect -1372 5881 -1338 6021
rect -1180 5881 -1146 6021
rect -988 5895 -954 6021
rect -1038 5881 -1028 5895
rect -2886 5847 -1028 5881
rect -2886 481 -2811 5847
rect -2068 5732 -2022 5744
rect -2068 5532 -2062 5732
rect -2028 5532 -2022 5732
rect -1948 5716 -1914 5847
rect -1756 5716 -1722 5847
rect -1564 5716 -1530 5847
rect -1372 5716 -1338 5847
rect -1180 5716 -1146 5847
rect -1038 5831 -1028 5847
rect -964 5831 -954 5895
rect -988 5716 -954 5831
rect -804 5881 -770 6444
rect 1618 6412 1628 6476
rect 1692 6412 1702 6476
rect -730 6334 -720 6386
rect -668 6334 -641 6386
rect -487 5881 -477 5893
rect -804 5847 -477 5881
rect -1954 5704 -1908 5716
rect -1954 5622 -1948 5704
rect -1914 5622 -1908 5704
rect -1954 5610 -1908 5622
rect -1858 5704 -1812 5716
rect -1858 5622 -1852 5704
rect -1818 5622 -1812 5704
rect -1858 5610 -1812 5622
rect -1762 5704 -1716 5716
rect -1762 5622 -1756 5704
rect -1722 5622 -1716 5704
rect -1762 5610 -1716 5622
rect -1666 5704 -1620 5716
rect -1666 5622 -1660 5704
rect -1626 5622 -1620 5704
rect -1666 5610 -1620 5622
rect -1570 5704 -1524 5716
rect -1570 5622 -1564 5704
rect -1530 5622 -1524 5704
rect -1570 5610 -1524 5622
rect -1474 5704 -1428 5716
rect -1474 5622 -1468 5704
rect -1434 5622 -1428 5704
rect -1474 5610 -1428 5622
rect -1378 5704 -1332 5716
rect -1378 5622 -1372 5704
rect -1338 5622 -1332 5704
rect -1378 5610 -1332 5622
rect -1282 5704 -1236 5716
rect -1282 5622 -1276 5704
rect -1242 5622 -1236 5704
rect -1282 5610 -1236 5622
rect -1186 5704 -1140 5716
rect -1186 5622 -1180 5704
rect -1146 5622 -1140 5704
rect -1186 5610 -1140 5622
rect -1090 5704 -1044 5716
rect -1090 5622 -1084 5704
rect -1050 5622 -1044 5704
rect -1090 5610 -1044 5622
rect -994 5704 -948 5716
rect -994 5622 -988 5704
rect -954 5622 -948 5704
rect -994 5610 -948 5622
rect -1964 5578 -1898 5582
rect -2068 5360 -2022 5532
rect -1967 5526 -1957 5578
rect -1905 5526 -1895 5578
rect -1964 5522 -1898 5526
rect -1852 5470 -1818 5610
rect -1772 5578 -1706 5582
rect -1775 5526 -1765 5578
rect -1713 5526 -1703 5578
rect -1772 5522 -1706 5526
rect -1660 5470 -1626 5610
rect -1580 5579 -1514 5582
rect -1582 5527 -1572 5579
rect -1520 5527 -1510 5579
rect -1580 5522 -1514 5527
rect -1468 5470 -1434 5610
rect -1388 5579 -1322 5582
rect -1390 5527 -1380 5579
rect -1328 5527 -1318 5579
rect -1388 5522 -1322 5527
rect -1276 5470 -1242 5610
rect -1196 5579 -1130 5582
rect -1198 5527 -1188 5579
rect -1136 5527 -1126 5579
rect -1196 5522 -1130 5527
rect -1084 5470 -1050 5610
rect -1004 5579 -938 5582
rect -1007 5527 -997 5579
rect -945 5527 -935 5579
rect -1004 5522 -938 5527
rect -804 5470 -770 5847
rect -487 5829 -477 5847
rect -413 5829 -403 5893
rect -730 5527 -720 5579
rect -668 5527 -641 5579
rect -1852 5436 -770 5470
rect -2068 4582 -2022 4760
rect -1852 4644 -770 4678
rect -2068 4196 -2062 4582
rect -2028 4196 -2022 4582
rect -1967 4534 -1957 4586
rect -1905 4534 -1895 4586
rect -1852 4495 -1818 4644
rect -1775 4534 -1765 4586
rect -1713 4534 -1703 4586
rect -1660 4495 -1626 4644
rect -1583 4534 -1573 4586
rect -1521 4534 -1511 4586
rect -1468 4495 -1434 4644
rect -1391 4534 -1381 4586
rect -1329 4534 -1319 4586
rect -1276 4495 -1242 4644
rect -1200 4534 -1190 4586
rect -1138 4534 -1128 4586
rect -1084 4495 -1050 4644
rect -1007 4534 -997 4586
rect -945 4534 -935 4586
rect -1954 4483 -1908 4495
rect -1954 4233 -1948 4483
rect -1914 4233 -1908 4483
rect -1954 4221 -1908 4233
rect -1858 4483 -1812 4495
rect -1858 4233 -1852 4483
rect -1818 4233 -1812 4483
rect -1858 4221 -1812 4233
rect -1762 4483 -1716 4495
rect -1762 4233 -1756 4483
rect -1722 4233 -1716 4483
rect -1762 4221 -1716 4233
rect -1666 4483 -1620 4495
rect -1666 4233 -1660 4483
rect -1626 4233 -1620 4483
rect -1666 4221 -1620 4233
rect -1570 4483 -1524 4495
rect -1570 4233 -1564 4483
rect -1530 4233 -1524 4483
rect -1570 4221 -1524 4233
rect -1474 4483 -1428 4495
rect -1474 4233 -1468 4483
rect -1434 4233 -1428 4483
rect -1474 4221 -1428 4233
rect -1378 4483 -1332 4495
rect -1378 4233 -1372 4483
rect -1338 4233 -1332 4483
rect -1378 4221 -1332 4233
rect -1282 4483 -1236 4495
rect -1282 4233 -1276 4483
rect -1242 4233 -1236 4483
rect -1282 4221 -1236 4233
rect -1186 4483 -1140 4495
rect -1186 4233 -1180 4483
rect -1146 4233 -1140 4483
rect -1186 4221 -1140 4233
rect -1090 4483 -1044 4495
rect -1090 4233 -1084 4483
rect -1050 4233 -1044 4483
rect -1090 4221 -1044 4233
rect -994 4483 -948 4495
rect -994 4233 -988 4483
rect -954 4233 -948 4483
rect -994 4221 -948 4233
rect -2068 4184 -2022 4196
rect -1948 4081 -1914 4221
rect -1756 4081 -1722 4221
rect -1564 4081 -1530 4221
rect -1372 4081 -1338 4221
rect -1180 4081 -1146 4221
rect -988 4095 -954 4221
rect -1034 4081 -1024 4095
rect -2428 4047 -1024 4081
rect -2428 2281 -2353 4047
rect -2068 3932 -2022 3944
rect -2068 3732 -2062 3932
rect -2028 3732 -2022 3932
rect -1948 3916 -1914 4047
rect -1756 3916 -1722 4047
rect -1564 3916 -1530 4047
rect -1372 3916 -1338 4047
rect -1180 3916 -1146 4047
rect -1034 4031 -1024 4047
rect -960 4031 -950 4095
rect -804 4081 -770 4644
rect -730 4534 -720 4586
rect -668 4534 -641 4586
rect -444 4081 -434 4094
rect -804 4047 -434 4081
rect -988 3916 -954 4031
rect -1954 3904 -1908 3916
rect -1954 3822 -1948 3904
rect -1914 3822 -1908 3904
rect -1954 3810 -1908 3822
rect -1858 3904 -1812 3916
rect -1858 3822 -1852 3904
rect -1818 3822 -1812 3904
rect -1858 3810 -1812 3822
rect -1762 3904 -1716 3916
rect -1762 3822 -1756 3904
rect -1722 3822 -1716 3904
rect -1762 3810 -1716 3822
rect -1666 3904 -1620 3916
rect -1666 3822 -1660 3904
rect -1626 3822 -1620 3904
rect -1666 3810 -1620 3822
rect -1570 3904 -1524 3916
rect -1570 3822 -1564 3904
rect -1530 3822 -1524 3904
rect -1570 3810 -1524 3822
rect -1474 3904 -1428 3916
rect -1474 3822 -1468 3904
rect -1434 3822 -1428 3904
rect -1474 3810 -1428 3822
rect -1378 3904 -1332 3916
rect -1378 3822 -1372 3904
rect -1338 3822 -1332 3904
rect -1378 3810 -1332 3822
rect -1282 3904 -1236 3916
rect -1282 3822 -1276 3904
rect -1242 3822 -1236 3904
rect -1282 3810 -1236 3822
rect -1186 3904 -1140 3916
rect -1186 3822 -1180 3904
rect -1146 3822 -1140 3904
rect -1186 3810 -1140 3822
rect -1090 3904 -1044 3916
rect -1090 3822 -1084 3904
rect -1050 3822 -1044 3904
rect -1090 3810 -1044 3822
rect -994 3904 -948 3916
rect -994 3822 -988 3904
rect -954 3822 -948 3904
rect -994 3810 -948 3822
rect -1964 3778 -1898 3782
rect -2068 3560 -2022 3732
rect -1967 3726 -1957 3778
rect -1905 3726 -1895 3778
rect -1964 3722 -1898 3726
rect -1852 3670 -1818 3810
rect -1772 3778 -1706 3782
rect -1775 3726 -1765 3778
rect -1713 3726 -1703 3778
rect -1772 3722 -1706 3726
rect -1660 3670 -1626 3810
rect -1580 3779 -1514 3782
rect -1582 3727 -1572 3779
rect -1520 3727 -1510 3779
rect -1580 3722 -1514 3727
rect -1468 3670 -1434 3810
rect -1388 3779 -1322 3782
rect -1390 3727 -1380 3779
rect -1328 3727 -1318 3779
rect -1388 3722 -1322 3727
rect -1276 3670 -1242 3810
rect -1196 3779 -1130 3782
rect -1198 3727 -1188 3779
rect -1136 3727 -1126 3779
rect -1196 3722 -1130 3727
rect -1084 3670 -1050 3810
rect -1004 3779 -938 3782
rect -1007 3727 -997 3779
rect -945 3727 -935 3779
rect -1004 3722 -938 3727
rect -804 3670 -770 4047
rect -444 4030 -434 4047
rect -370 4030 -360 4094
rect 1628 3846 1692 6412
rect 2347 4563 2411 7633
rect 6932 7532 6978 7544
rect 6932 7332 6938 7532
rect 6972 7332 6978 7532
rect 7052 7516 7086 7647
rect 7244 7516 7278 7647
rect 7436 7516 7470 7647
rect 7628 7516 7662 7647
rect 7820 7516 7854 7647
rect 8012 7516 8046 7647
rect 8196 7681 8230 8244
rect 8270 8134 8280 8186
rect 8332 8134 8359 8186
rect 8196 7647 9310 7681
rect 7046 7504 7092 7516
rect 7046 7422 7052 7504
rect 7086 7422 7092 7504
rect 7046 7410 7092 7422
rect 7142 7504 7188 7516
rect 7142 7422 7148 7504
rect 7182 7422 7188 7504
rect 7142 7410 7188 7422
rect 7238 7504 7284 7516
rect 7238 7422 7244 7504
rect 7278 7422 7284 7504
rect 7238 7410 7284 7422
rect 7334 7504 7380 7516
rect 7334 7422 7340 7504
rect 7374 7422 7380 7504
rect 7334 7410 7380 7422
rect 7430 7504 7476 7516
rect 7430 7422 7436 7504
rect 7470 7422 7476 7504
rect 7430 7410 7476 7422
rect 7526 7504 7572 7516
rect 7526 7422 7532 7504
rect 7566 7422 7572 7504
rect 7526 7410 7572 7422
rect 7622 7504 7668 7516
rect 7622 7422 7628 7504
rect 7662 7422 7668 7504
rect 7622 7410 7668 7422
rect 7718 7504 7764 7516
rect 7718 7422 7724 7504
rect 7758 7422 7764 7504
rect 7718 7410 7764 7422
rect 7814 7504 7860 7516
rect 7814 7422 7820 7504
rect 7854 7422 7860 7504
rect 7814 7410 7860 7422
rect 7910 7504 7956 7516
rect 7910 7422 7916 7504
rect 7950 7422 7956 7504
rect 7910 7410 7956 7422
rect 8006 7504 8052 7516
rect 8006 7422 8012 7504
rect 8046 7422 8052 7504
rect 8006 7410 8052 7422
rect 7036 7378 7102 7382
rect 6932 7160 6978 7332
rect 7033 7326 7043 7378
rect 7095 7326 7105 7378
rect 7036 7322 7102 7326
rect 7148 7270 7182 7410
rect 7228 7378 7294 7382
rect 7225 7326 7235 7378
rect 7287 7326 7297 7378
rect 7228 7322 7294 7326
rect 7340 7270 7374 7410
rect 7420 7379 7486 7382
rect 7418 7327 7428 7379
rect 7480 7327 7490 7379
rect 7420 7322 7486 7327
rect 7532 7270 7566 7410
rect 7612 7379 7678 7382
rect 7610 7327 7620 7379
rect 7672 7327 7682 7379
rect 7612 7322 7678 7327
rect 7724 7270 7758 7410
rect 7804 7379 7870 7382
rect 7802 7327 7812 7379
rect 7864 7327 7874 7379
rect 7804 7322 7870 7327
rect 7916 7270 7950 7410
rect 7996 7379 8062 7382
rect 7993 7327 8003 7379
rect 8055 7327 8065 7379
rect 7996 7322 8062 7327
rect 8196 7270 8230 7647
rect 8270 7327 8280 7379
rect 8332 7327 8359 7379
rect 7148 7236 8230 7270
rect 6932 6382 6978 6560
rect 7148 6444 8230 6478
rect 6932 5996 6938 6382
rect 6972 5996 6978 6382
rect 7033 6334 7043 6386
rect 7095 6334 7105 6386
rect 7148 6295 7182 6444
rect 7225 6334 7235 6386
rect 7287 6334 7297 6386
rect 7340 6295 7374 6444
rect 7417 6334 7427 6386
rect 7479 6334 7489 6386
rect 7532 6295 7566 6444
rect 7609 6334 7619 6386
rect 7671 6334 7681 6386
rect 7724 6295 7758 6444
rect 7800 6334 7810 6386
rect 7862 6334 7872 6386
rect 7916 6295 7950 6444
rect 7993 6334 8003 6386
rect 8055 6334 8065 6386
rect 7046 6283 7092 6295
rect 7046 6033 7052 6283
rect 7086 6033 7092 6283
rect 7046 6021 7092 6033
rect 7142 6283 7188 6295
rect 7142 6033 7148 6283
rect 7182 6033 7188 6283
rect 7142 6021 7188 6033
rect 7238 6283 7284 6295
rect 7238 6033 7244 6283
rect 7278 6033 7284 6283
rect 7238 6021 7284 6033
rect 7334 6283 7380 6295
rect 7334 6033 7340 6283
rect 7374 6033 7380 6283
rect 7334 6021 7380 6033
rect 7430 6283 7476 6295
rect 7430 6033 7436 6283
rect 7470 6033 7476 6283
rect 7430 6021 7476 6033
rect 7526 6283 7572 6295
rect 7526 6033 7532 6283
rect 7566 6033 7572 6283
rect 7526 6021 7572 6033
rect 7622 6283 7668 6295
rect 7622 6033 7628 6283
rect 7662 6033 7668 6283
rect 7622 6021 7668 6033
rect 7718 6283 7764 6295
rect 7718 6033 7724 6283
rect 7758 6033 7764 6283
rect 7718 6021 7764 6033
rect 7814 6283 7860 6295
rect 7814 6033 7820 6283
rect 7854 6033 7860 6283
rect 7814 6021 7860 6033
rect 7910 6283 7956 6295
rect 7910 6033 7916 6283
rect 7950 6033 7956 6283
rect 7910 6021 7956 6033
rect 8006 6283 8052 6295
rect 8006 6033 8012 6283
rect 8046 6033 8052 6283
rect 8006 6021 8052 6033
rect 6932 5984 6978 5996
rect 6694 5831 6704 5895
rect 6768 5881 6778 5895
rect 7052 5881 7086 6021
rect 7244 5881 7278 6021
rect 7436 5881 7470 6021
rect 7628 5881 7662 6021
rect 7820 5881 7854 6021
rect 8012 5881 8046 6021
rect 6768 5847 8046 5881
rect 6768 5831 6778 5847
rect 6932 5732 6978 5744
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 6932 5532 6938 5732
rect 6972 5532 6978 5732
rect 7052 5716 7086 5847
rect 7244 5716 7278 5847
rect 7436 5716 7470 5847
rect 7628 5716 7662 5847
rect 7820 5716 7854 5847
rect 8012 5716 8046 5847
rect 8196 5881 8230 6444
rect 8270 6334 8280 6386
rect 8332 6334 8359 6386
rect 8196 5847 8799 5881
rect 7046 5704 7092 5716
rect 7046 5622 7052 5704
rect 7086 5622 7092 5704
rect 7046 5610 7092 5622
rect 7142 5704 7188 5716
rect 7142 5622 7148 5704
rect 7182 5622 7188 5704
rect 7142 5610 7188 5622
rect 7238 5704 7284 5716
rect 7238 5622 7244 5704
rect 7278 5622 7284 5704
rect 7238 5610 7284 5622
rect 7334 5704 7380 5716
rect 7334 5622 7340 5704
rect 7374 5622 7380 5704
rect 7334 5610 7380 5622
rect 7430 5704 7476 5716
rect 7430 5622 7436 5704
rect 7470 5622 7476 5704
rect 7430 5610 7476 5622
rect 7526 5704 7572 5716
rect 7526 5622 7532 5704
rect 7566 5622 7572 5704
rect 7526 5610 7572 5622
rect 7622 5704 7668 5716
rect 7622 5622 7628 5704
rect 7662 5622 7668 5704
rect 7622 5610 7668 5622
rect 7718 5704 7764 5716
rect 7718 5622 7724 5704
rect 7758 5622 7764 5704
rect 7718 5610 7764 5622
rect 7814 5704 7860 5716
rect 7814 5622 7820 5704
rect 7854 5622 7860 5704
rect 7814 5610 7860 5622
rect 7910 5704 7956 5716
rect 7910 5622 7916 5704
rect 7950 5622 7956 5704
rect 7910 5610 7956 5622
rect 8006 5704 8052 5716
rect 8006 5622 8012 5704
rect 8046 5622 8052 5704
rect 8006 5610 8052 5622
rect 7036 5578 7102 5582
rect 3157 5084 3221 5494
rect 6932 5360 6978 5532
rect 7033 5526 7043 5578
rect 7095 5526 7105 5578
rect 7036 5522 7102 5526
rect 7148 5470 7182 5610
rect 7228 5578 7294 5582
rect 7225 5526 7235 5578
rect 7287 5526 7297 5578
rect 7228 5522 7294 5526
rect 7340 5470 7374 5610
rect 7420 5579 7486 5582
rect 7418 5527 7428 5579
rect 7480 5527 7490 5579
rect 7420 5522 7486 5527
rect 7532 5470 7566 5610
rect 7612 5579 7678 5582
rect 7610 5527 7620 5579
rect 7672 5527 7682 5579
rect 7612 5522 7678 5527
rect 7724 5470 7758 5610
rect 7804 5579 7870 5582
rect 7802 5527 7812 5579
rect 7864 5527 7874 5579
rect 7804 5522 7870 5527
rect 7916 5470 7950 5610
rect 7996 5579 8062 5582
rect 7993 5527 8003 5579
rect 8055 5527 8065 5579
rect 7996 5522 8062 5527
rect 8196 5470 8230 5847
rect 8270 5527 8280 5579
rect 8332 5527 8359 5579
rect 7148 5436 8230 5470
rect 3147 5020 3157 5084
rect 3221 5020 3231 5084
rect 3831 4928 6166 4932
rect 3758 4864 3768 4928
rect 3832 4868 6166 4928
rect 6230 4868 6240 4932
rect 3832 4864 3842 4868
rect 6932 4582 6978 4760
rect 7148 4644 8230 4678
rect 2347 4499 3106 4563
rect 3170 4499 3180 4563
rect 4874 4326 5207 4390
rect 5271 4326 5281 4390
rect 3298 4148 3308 4212
rect 3372 4148 3382 4212
rect 3308 4085 3372 4148
rect 1628 3782 1866 3846
rect -730 3727 -720 3779
rect -668 3727 -641 3779
rect -1852 3636 -770 3670
rect 323 3419 333 3483
rect 397 3419 1631 3483
rect 1695 3419 1705 3483
rect 1802 3154 1866 3782
rect 323 3090 333 3154
rect 397 3090 1866 3154
rect -2068 2782 -2022 2960
rect -1852 2844 -770 2878
rect -2068 2396 -2062 2782
rect -2028 2396 -2022 2782
rect -1967 2734 -1957 2786
rect -1905 2734 -1895 2786
rect -1852 2695 -1818 2844
rect -1775 2734 -1765 2786
rect -1713 2734 -1703 2786
rect -1660 2695 -1626 2844
rect -1583 2734 -1573 2786
rect -1521 2734 -1511 2786
rect -1468 2695 -1434 2844
rect -1391 2734 -1381 2786
rect -1329 2734 -1319 2786
rect -1276 2695 -1242 2844
rect -1200 2734 -1190 2786
rect -1138 2734 -1128 2786
rect -1084 2695 -1050 2844
rect -1007 2734 -997 2786
rect -945 2734 -935 2786
rect -1954 2683 -1908 2695
rect -1954 2433 -1948 2683
rect -1914 2433 -1908 2683
rect -1954 2421 -1908 2433
rect -1858 2683 -1812 2695
rect -1858 2433 -1852 2683
rect -1818 2433 -1812 2683
rect -1858 2421 -1812 2433
rect -1762 2683 -1716 2695
rect -1762 2433 -1756 2683
rect -1722 2433 -1716 2683
rect -1762 2421 -1716 2433
rect -1666 2683 -1620 2695
rect -1666 2433 -1660 2683
rect -1626 2433 -1620 2683
rect -1666 2421 -1620 2433
rect -1570 2683 -1524 2695
rect -1570 2433 -1564 2683
rect -1530 2433 -1524 2683
rect -1570 2421 -1524 2433
rect -1474 2683 -1428 2695
rect -1474 2433 -1468 2683
rect -1434 2433 -1428 2683
rect -1474 2421 -1428 2433
rect -1378 2683 -1332 2695
rect -1378 2433 -1372 2683
rect -1338 2433 -1332 2683
rect -1378 2421 -1332 2433
rect -1282 2683 -1236 2695
rect -1282 2433 -1276 2683
rect -1242 2433 -1236 2683
rect -1282 2421 -1236 2433
rect -1186 2683 -1140 2695
rect -1186 2433 -1180 2683
rect -1146 2433 -1140 2683
rect -1186 2421 -1140 2433
rect -1090 2683 -1044 2695
rect -1090 2433 -1084 2683
rect -1050 2433 -1044 2683
rect -1090 2421 -1044 2433
rect -994 2683 -948 2695
rect -994 2433 -988 2683
rect -954 2433 -948 2683
rect -994 2421 -948 2433
rect -2068 2384 -2022 2396
rect -1948 2281 -1914 2421
rect -1756 2281 -1722 2421
rect -1564 2281 -1530 2421
rect -1372 2281 -1338 2421
rect -1180 2281 -1146 2421
rect -988 2295 -954 2421
rect -1037 2281 -1027 2295
rect -2428 2247 -1027 2281
rect -2068 2132 -2022 2144
rect -2068 1932 -2062 2132
rect -2028 1932 -2022 2132
rect -1948 2116 -1914 2247
rect -1756 2116 -1722 2247
rect -1564 2116 -1530 2247
rect -1372 2116 -1338 2247
rect -1180 2116 -1146 2247
rect -1037 2231 -1027 2247
rect -963 2231 -953 2295
rect -804 2281 -770 2844
rect -730 2734 -720 2786
rect -668 2734 -641 2786
rect -444 2281 -434 2291
rect -804 2247 -434 2281
rect -988 2116 -954 2231
rect -1954 2104 -1908 2116
rect -1954 2022 -1948 2104
rect -1914 2022 -1908 2104
rect -1954 2010 -1908 2022
rect -1858 2104 -1812 2116
rect -1858 2022 -1852 2104
rect -1818 2022 -1812 2104
rect -1858 2010 -1812 2022
rect -1762 2104 -1716 2116
rect -1762 2022 -1756 2104
rect -1722 2022 -1716 2104
rect -1762 2010 -1716 2022
rect -1666 2104 -1620 2116
rect -1666 2022 -1660 2104
rect -1626 2022 -1620 2104
rect -1666 2010 -1620 2022
rect -1570 2104 -1524 2116
rect -1570 2022 -1564 2104
rect -1530 2022 -1524 2104
rect -1570 2010 -1524 2022
rect -1474 2104 -1428 2116
rect -1474 2022 -1468 2104
rect -1434 2022 -1428 2104
rect -1474 2010 -1428 2022
rect -1378 2104 -1332 2116
rect -1378 2022 -1372 2104
rect -1338 2022 -1332 2104
rect -1378 2010 -1332 2022
rect -1282 2104 -1236 2116
rect -1282 2022 -1276 2104
rect -1242 2022 -1236 2104
rect -1282 2010 -1236 2022
rect -1186 2104 -1140 2116
rect -1186 2022 -1180 2104
rect -1146 2022 -1140 2104
rect -1186 2010 -1140 2022
rect -1090 2104 -1044 2116
rect -1090 2022 -1084 2104
rect -1050 2022 -1044 2104
rect -1090 2010 -1044 2022
rect -994 2104 -948 2116
rect -994 2022 -988 2104
rect -954 2022 -948 2104
rect -994 2010 -948 2022
rect -1964 1978 -1898 1982
rect -2068 1760 -2022 1932
rect -1967 1926 -1957 1978
rect -1905 1926 -1895 1978
rect -1964 1922 -1898 1926
rect -1852 1870 -1818 2010
rect -1772 1978 -1706 1982
rect -1775 1926 -1765 1978
rect -1713 1926 -1703 1978
rect -1772 1922 -1706 1926
rect -1660 1870 -1626 2010
rect -1580 1979 -1514 1982
rect -1582 1927 -1572 1979
rect -1520 1927 -1510 1979
rect -1580 1922 -1514 1927
rect -1468 1870 -1434 2010
rect -1388 1979 -1322 1982
rect -1390 1927 -1380 1979
rect -1328 1927 -1318 1979
rect -1388 1922 -1322 1927
rect -1276 1870 -1242 2010
rect -1196 1979 -1130 1982
rect -1198 1927 -1188 1979
rect -1136 1927 -1126 1979
rect -1196 1922 -1130 1927
rect -1084 1870 -1050 2010
rect -1004 1979 -938 1982
rect -1007 1927 -997 1979
rect -945 1927 -935 1979
rect -1004 1922 -938 1927
rect -804 1870 -770 2247
rect -444 2227 -434 2247
rect -370 2227 -360 2291
rect 3308 2223 3371 4085
rect 4874 3642 4938 4326
rect 6932 4196 6938 4582
rect 6972 4196 6978 4582
rect 7033 4534 7043 4586
rect 7095 4534 7105 4586
rect 7148 4495 7182 4644
rect 7225 4534 7235 4586
rect 7287 4534 7297 4586
rect 7340 4495 7374 4644
rect 7417 4534 7427 4586
rect 7479 4534 7489 4586
rect 7532 4495 7566 4644
rect 7609 4534 7619 4586
rect 7671 4534 7681 4586
rect 7724 4495 7758 4644
rect 7800 4534 7810 4586
rect 7862 4534 7872 4586
rect 7916 4495 7950 4644
rect 7993 4534 8003 4586
rect 8055 4534 8065 4586
rect 7046 4483 7092 4495
rect 7046 4233 7052 4483
rect 7086 4233 7092 4483
rect 7046 4221 7092 4233
rect 7142 4483 7188 4495
rect 7142 4233 7148 4483
rect 7182 4233 7188 4483
rect 7142 4221 7188 4233
rect 7238 4483 7284 4495
rect 7238 4233 7244 4483
rect 7278 4233 7284 4483
rect 7238 4221 7284 4233
rect 7334 4483 7380 4495
rect 7334 4233 7340 4483
rect 7374 4233 7380 4483
rect 7334 4221 7380 4233
rect 7430 4483 7476 4495
rect 7430 4233 7436 4483
rect 7470 4233 7476 4483
rect 7430 4221 7476 4233
rect 7526 4483 7572 4495
rect 7526 4233 7532 4483
rect 7566 4233 7572 4483
rect 7526 4221 7572 4233
rect 7622 4483 7668 4495
rect 7622 4233 7628 4483
rect 7662 4233 7668 4483
rect 7622 4221 7668 4233
rect 7718 4483 7764 4495
rect 7718 4233 7724 4483
rect 7758 4233 7764 4483
rect 7718 4221 7764 4233
rect 7814 4483 7860 4495
rect 7814 4233 7820 4483
rect 7854 4233 7860 4483
rect 7814 4221 7860 4233
rect 7910 4483 7956 4495
rect 7910 4233 7916 4483
rect 7950 4233 7956 4483
rect 7910 4221 7956 4233
rect 8006 4483 8052 4495
rect 8006 4233 8012 4483
rect 8046 4233 8052 4483
rect 8006 4221 8052 4233
rect 6932 4184 6978 4196
rect 6749 4031 6759 4095
rect 6823 4081 6833 4095
rect 7052 4081 7086 4221
rect 7244 4081 7278 4221
rect 7436 4081 7470 4221
rect 7628 4081 7662 4221
rect 7820 4081 7854 4221
rect 8012 4081 8046 4221
rect 6823 4047 8046 4081
rect 6823 4031 6833 4047
rect 6932 3932 6978 3944
rect 6932 3732 6938 3932
rect 6972 3732 6978 3932
rect 7052 3916 7086 4047
rect 7244 3916 7278 4047
rect 7436 3916 7470 4047
rect 7628 3916 7662 4047
rect 7820 3916 7854 4047
rect 8012 3916 8046 4047
rect 8196 4081 8230 4644
rect 8270 4534 8280 4586
rect 8332 4534 8359 4586
rect 8724 4081 8799 5847
rect 8196 4047 8799 4081
rect 7046 3904 7092 3916
rect 7046 3822 7052 3904
rect 7086 3822 7092 3904
rect 7046 3810 7092 3822
rect 7142 3904 7188 3916
rect 7142 3822 7148 3904
rect 7182 3822 7188 3904
rect 7142 3810 7188 3822
rect 7238 3904 7284 3916
rect 7238 3822 7244 3904
rect 7278 3822 7284 3904
rect 7238 3810 7284 3822
rect 7334 3904 7380 3916
rect 7334 3822 7340 3904
rect 7374 3822 7380 3904
rect 7334 3810 7380 3822
rect 7430 3904 7476 3916
rect 7430 3822 7436 3904
rect 7470 3822 7476 3904
rect 7430 3810 7476 3822
rect 7526 3904 7572 3916
rect 7526 3822 7532 3904
rect 7566 3822 7572 3904
rect 7526 3810 7572 3822
rect 7622 3904 7668 3916
rect 7622 3822 7628 3904
rect 7662 3822 7668 3904
rect 7622 3810 7668 3822
rect 7718 3904 7764 3916
rect 7718 3822 7724 3904
rect 7758 3822 7764 3904
rect 7718 3810 7764 3822
rect 7814 3904 7860 3916
rect 7814 3822 7820 3904
rect 7854 3822 7860 3904
rect 7814 3810 7860 3822
rect 7910 3904 7956 3916
rect 7910 3822 7916 3904
rect 7950 3822 7956 3904
rect 7910 3810 7956 3822
rect 8006 3904 8052 3916
rect 8006 3822 8012 3904
rect 8046 3822 8052 3904
rect 8006 3810 8052 3822
rect 7036 3778 7102 3782
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 6932 3560 6978 3732
rect 7033 3726 7043 3778
rect 7095 3726 7105 3778
rect 7036 3722 7102 3726
rect 7148 3670 7182 3810
rect 7228 3778 7294 3782
rect 7225 3726 7235 3778
rect 7287 3726 7297 3778
rect 7228 3722 7294 3726
rect 7340 3670 7374 3810
rect 7420 3779 7486 3782
rect 7418 3727 7428 3779
rect 7480 3727 7490 3779
rect 7420 3722 7486 3727
rect 7532 3670 7566 3810
rect 7612 3779 7678 3782
rect 7610 3727 7620 3779
rect 7672 3727 7682 3779
rect 7612 3722 7678 3727
rect 7724 3670 7758 3810
rect 7804 3779 7870 3782
rect 7802 3727 7812 3779
rect 7864 3727 7874 3779
rect 7804 3722 7870 3727
rect 7916 3670 7950 3810
rect 7996 3779 8062 3782
rect 7993 3727 8003 3779
rect 8055 3727 8065 3779
rect 7996 3722 8062 3727
rect 8196 3670 8230 4047
rect 8270 3727 8280 3779
rect 8332 3727 8359 3779
rect 7148 3636 8230 3670
rect 6932 2782 6978 2960
rect 7148 2844 8230 2878
rect 6932 2396 6938 2782
rect 6972 2396 6978 2782
rect 7033 2734 7043 2786
rect 7095 2734 7105 2786
rect 7148 2695 7182 2844
rect 7225 2734 7235 2786
rect 7287 2734 7297 2786
rect 7340 2695 7374 2844
rect 7417 2734 7427 2786
rect 7479 2734 7489 2786
rect 7532 2695 7566 2844
rect 7609 2734 7619 2786
rect 7671 2734 7681 2786
rect 7724 2695 7758 2844
rect 7800 2734 7810 2786
rect 7862 2734 7872 2786
rect 7916 2695 7950 2844
rect 7993 2734 8003 2786
rect 8055 2734 8065 2786
rect 7046 2683 7092 2695
rect 7046 2433 7052 2683
rect 7086 2433 7092 2683
rect 7046 2421 7092 2433
rect 7142 2683 7188 2695
rect 7142 2433 7148 2683
rect 7182 2433 7188 2683
rect 7142 2421 7188 2433
rect 7238 2683 7284 2695
rect 7238 2433 7244 2683
rect 7278 2433 7284 2683
rect 7238 2421 7284 2433
rect 7334 2683 7380 2695
rect 7334 2433 7340 2683
rect 7374 2433 7380 2683
rect 7334 2421 7380 2433
rect 7430 2683 7476 2695
rect 7430 2433 7436 2683
rect 7470 2433 7476 2683
rect 7430 2421 7476 2433
rect 7526 2683 7572 2695
rect 7526 2433 7532 2683
rect 7566 2433 7572 2683
rect 7526 2421 7572 2433
rect 7622 2683 7668 2695
rect 7622 2433 7628 2683
rect 7662 2433 7668 2683
rect 7622 2421 7668 2433
rect 7718 2683 7764 2695
rect 7718 2433 7724 2683
rect 7758 2433 7764 2683
rect 7718 2421 7764 2433
rect 7814 2683 7860 2695
rect 7814 2433 7820 2683
rect 7854 2433 7860 2683
rect 7814 2421 7860 2433
rect 7910 2683 7956 2695
rect 7910 2433 7916 2683
rect 7950 2433 7956 2683
rect 7910 2421 7956 2433
rect 8006 2683 8052 2695
rect 8006 2433 8012 2683
rect 8046 2433 8052 2683
rect 8006 2421 8052 2433
rect 6932 2384 6978 2396
rect 6754 2233 6764 2297
rect 6828 2281 6838 2297
rect 7052 2281 7086 2421
rect 7244 2281 7278 2421
rect 7436 2281 7470 2421
rect 7628 2281 7662 2421
rect 7820 2281 7854 2421
rect 8012 2281 8046 2421
rect 6828 2247 8046 2281
rect 6828 2233 6838 2247
rect 3298 2159 3308 2223
rect 3372 2159 3382 2223
rect 6932 2132 6978 2144
rect -730 1927 -720 1979
rect -668 1927 -641 1979
rect 6932 1932 6938 2132
rect 6972 1932 6978 2132
rect 7052 2116 7086 2247
rect 7244 2116 7278 2247
rect 7436 2116 7470 2247
rect 7628 2116 7662 2247
rect 7820 2116 7854 2247
rect 8012 2116 8046 2247
rect 8196 2281 8230 2844
rect 8270 2734 8280 2786
rect 8332 2734 8359 2786
rect 8724 2281 8799 4047
rect 8196 2247 8799 2281
rect 7046 2104 7092 2116
rect 7046 2022 7052 2104
rect 7086 2022 7092 2104
rect 7046 2010 7092 2022
rect 7142 2104 7188 2116
rect 7142 2022 7148 2104
rect 7182 2022 7188 2104
rect 7142 2010 7188 2022
rect 7238 2104 7284 2116
rect 7238 2022 7244 2104
rect 7278 2022 7284 2104
rect 7238 2010 7284 2022
rect 7334 2104 7380 2116
rect 7334 2022 7340 2104
rect 7374 2022 7380 2104
rect 7334 2010 7380 2022
rect 7430 2104 7476 2116
rect 7430 2022 7436 2104
rect 7470 2022 7476 2104
rect 7430 2010 7476 2022
rect 7526 2104 7572 2116
rect 7526 2022 7532 2104
rect 7566 2022 7572 2104
rect 7526 2010 7572 2022
rect 7622 2104 7668 2116
rect 7622 2022 7628 2104
rect 7662 2022 7668 2104
rect 7622 2010 7668 2022
rect 7718 2104 7764 2116
rect 7718 2022 7724 2104
rect 7758 2022 7764 2104
rect 7718 2010 7764 2022
rect 7814 2104 7860 2116
rect 7814 2022 7820 2104
rect 7854 2022 7860 2104
rect 7814 2010 7860 2022
rect 7910 2104 7956 2116
rect 7910 2022 7916 2104
rect 7950 2022 7956 2104
rect 7910 2010 7956 2022
rect 8006 2104 8052 2116
rect 8006 2022 8012 2104
rect 8046 2022 8052 2104
rect 8006 2010 8052 2022
rect 7036 1978 7102 1982
rect -1852 1836 -770 1870
rect 6932 1760 6978 1932
rect 7033 1926 7043 1978
rect 7095 1926 7105 1978
rect 7036 1922 7102 1926
rect 7148 1870 7182 2010
rect 7228 1978 7294 1982
rect 7225 1926 7235 1978
rect 7287 1926 7297 1978
rect 7228 1922 7294 1926
rect 7340 1870 7374 2010
rect 7420 1979 7486 1982
rect 7418 1927 7428 1979
rect 7480 1927 7490 1979
rect 7420 1922 7486 1927
rect 7532 1870 7566 2010
rect 7612 1979 7678 1982
rect 7610 1927 7620 1979
rect 7672 1927 7682 1979
rect 7612 1922 7678 1927
rect 7724 1870 7758 2010
rect 7804 1979 7870 1982
rect 7802 1927 7812 1979
rect 7864 1927 7874 1979
rect 7804 1922 7870 1927
rect 7916 1870 7950 2010
rect 7996 1979 8062 1982
rect 7993 1927 8003 1979
rect 8055 1927 8065 1979
rect 7996 1922 8062 1927
rect 8196 1870 8230 2247
rect 8270 1927 8280 1979
rect 8332 1927 8359 1979
rect 7148 1836 8230 1870
rect -364 1576 2330 1640
rect 2394 1576 2404 1640
rect -2068 982 -2022 1160
rect -1852 1044 -770 1078
rect -2068 596 -2062 982
rect -2028 596 -2022 982
rect -1967 934 -1957 986
rect -1905 934 -1895 986
rect -1852 895 -1818 1044
rect -1775 934 -1765 986
rect -1713 934 -1703 986
rect -1660 895 -1626 1044
rect -1583 934 -1573 986
rect -1521 934 -1511 986
rect -1468 895 -1434 1044
rect -1391 934 -1381 986
rect -1329 934 -1319 986
rect -1276 895 -1242 1044
rect -1200 934 -1190 986
rect -1138 934 -1128 986
rect -1084 895 -1050 1044
rect -1007 934 -997 986
rect -945 934 -935 986
rect -1954 883 -1908 895
rect -1954 633 -1948 883
rect -1914 633 -1908 883
rect -1954 621 -1908 633
rect -1858 883 -1812 895
rect -1858 633 -1852 883
rect -1818 633 -1812 883
rect -1858 621 -1812 633
rect -1762 883 -1716 895
rect -1762 633 -1756 883
rect -1722 633 -1716 883
rect -1762 621 -1716 633
rect -1666 883 -1620 895
rect -1666 633 -1660 883
rect -1626 633 -1620 883
rect -1666 621 -1620 633
rect -1570 883 -1524 895
rect -1570 633 -1564 883
rect -1530 633 -1524 883
rect -1570 621 -1524 633
rect -1474 883 -1428 895
rect -1474 633 -1468 883
rect -1434 633 -1428 883
rect -1474 621 -1428 633
rect -1378 883 -1332 895
rect -1378 633 -1372 883
rect -1338 633 -1332 883
rect -1378 621 -1332 633
rect -1282 883 -1236 895
rect -1282 633 -1276 883
rect -1242 633 -1236 883
rect -1282 621 -1236 633
rect -1186 883 -1140 895
rect -1186 633 -1180 883
rect -1146 633 -1140 883
rect -1186 621 -1140 633
rect -1090 883 -1044 895
rect -1090 633 -1084 883
rect -1050 633 -1044 883
rect -1090 621 -1044 633
rect -994 883 -948 895
rect -994 633 -988 883
rect -954 633 -948 883
rect -994 621 -948 633
rect -2068 584 -2022 596
rect -1948 481 -1914 621
rect -1756 481 -1722 621
rect -1564 481 -1530 621
rect -1372 481 -1338 621
rect -1180 481 -1146 621
rect -988 497 -954 621
rect -1030 481 -1020 497
rect -2886 447 -1020 481
rect -2068 332 -2022 344
rect -2068 132 -2062 332
rect -2028 132 -2022 332
rect -1948 316 -1914 447
rect -1756 316 -1722 447
rect -1564 316 -1530 447
rect -1372 316 -1338 447
rect -1180 316 -1146 447
rect -1030 433 -1020 447
rect -956 433 -946 497
rect -804 481 -770 1044
rect -730 934 -720 986
rect -668 934 -641 986
rect -364 481 -300 1576
rect 3592 1462 3602 1526
rect 3666 1462 6152 1526
rect 6216 1462 6226 1526
rect 160 1277 170 1341
rect 234 1277 4326 1341
rect 4390 1277 4400 1341
rect 6932 982 6978 1160
rect 7148 1044 8230 1078
rect 6932 596 6938 982
rect 6972 596 6978 982
rect 7033 934 7043 986
rect 7095 934 7105 986
rect 7148 895 7182 1044
rect 7225 934 7235 986
rect 7287 934 7297 986
rect 7340 895 7374 1044
rect 7417 934 7427 986
rect 7479 934 7489 986
rect 7532 895 7566 1044
rect 7609 934 7619 986
rect 7671 934 7681 986
rect 7724 895 7758 1044
rect 7800 934 7810 986
rect 7862 934 7872 986
rect 7916 895 7950 1044
rect 7993 934 8003 986
rect 8055 934 8065 986
rect 7046 883 7092 895
rect 7046 633 7052 883
rect 7086 633 7092 883
rect 7046 621 7092 633
rect 7142 883 7188 895
rect 7142 633 7148 883
rect 7182 633 7188 883
rect 7142 621 7188 633
rect 7238 883 7284 895
rect 7238 633 7244 883
rect 7278 633 7284 883
rect 7238 621 7284 633
rect 7334 883 7380 895
rect 7334 633 7340 883
rect 7374 633 7380 883
rect 7334 621 7380 633
rect 7430 883 7476 895
rect 7430 633 7436 883
rect 7470 633 7476 883
rect 7430 621 7476 633
rect 7526 883 7572 895
rect 7526 633 7532 883
rect 7566 633 7572 883
rect 7526 621 7572 633
rect 7622 883 7668 895
rect 7622 633 7628 883
rect 7662 633 7668 883
rect 7622 621 7668 633
rect 7718 883 7764 895
rect 7718 633 7724 883
rect 7758 633 7764 883
rect 7718 621 7764 633
rect 7814 883 7860 895
rect 7814 633 7820 883
rect 7854 633 7860 883
rect 7814 621 7860 633
rect 7910 883 7956 895
rect 7910 633 7916 883
rect 7950 633 7956 883
rect 7910 621 7956 633
rect 8006 883 8052 895
rect 8006 633 8012 883
rect 8046 633 8052 883
rect 8006 621 8052 633
rect 6932 584 6978 596
rect -804 447 -300 481
rect -988 316 -954 433
rect -1954 304 -1908 316
rect -1954 222 -1948 304
rect -1914 222 -1908 304
rect -1954 210 -1908 222
rect -1858 304 -1812 316
rect -1858 222 -1852 304
rect -1818 222 -1812 304
rect -1858 210 -1812 222
rect -1762 304 -1716 316
rect -1762 222 -1756 304
rect -1722 222 -1716 304
rect -1762 210 -1716 222
rect -1666 304 -1620 316
rect -1666 222 -1660 304
rect -1626 222 -1620 304
rect -1666 210 -1620 222
rect -1570 304 -1524 316
rect -1570 222 -1564 304
rect -1530 222 -1524 304
rect -1570 210 -1524 222
rect -1474 304 -1428 316
rect -1474 222 -1468 304
rect -1434 222 -1428 304
rect -1474 210 -1428 222
rect -1378 304 -1332 316
rect -1378 222 -1372 304
rect -1338 222 -1332 304
rect -1378 210 -1332 222
rect -1282 304 -1236 316
rect -1282 222 -1276 304
rect -1242 222 -1236 304
rect -1282 210 -1236 222
rect -1186 304 -1140 316
rect -1186 222 -1180 304
rect -1146 222 -1140 304
rect -1186 210 -1140 222
rect -1090 304 -1044 316
rect -1090 222 -1084 304
rect -1050 222 -1044 304
rect -1090 210 -1044 222
rect -994 304 -948 316
rect -994 222 -988 304
rect -954 222 -948 304
rect -994 210 -948 222
rect -1964 178 -1898 182
rect -2068 -40 -2022 132
rect -1967 126 -1957 178
rect -1905 126 -1895 178
rect -1964 122 -1898 126
rect -1852 70 -1818 210
rect -1772 178 -1706 182
rect -1775 126 -1765 178
rect -1713 126 -1703 178
rect -1772 122 -1706 126
rect -1660 70 -1626 210
rect -1580 179 -1514 182
rect -1582 127 -1572 179
rect -1520 127 -1510 179
rect -1580 122 -1514 127
rect -1468 70 -1434 210
rect -1388 179 -1322 182
rect -1390 127 -1380 179
rect -1328 127 -1318 179
rect -1388 122 -1322 127
rect -1276 70 -1242 210
rect -1196 179 -1130 182
rect -1198 127 -1188 179
rect -1136 127 -1126 179
rect -1196 122 -1130 127
rect -1084 70 -1050 210
rect -1004 179 -938 182
rect -1007 127 -997 179
rect -945 127 -935 179
rect -1004 122 -938 127
rect -804 70 -770 447
rect -364 446 -300 447
rect 6690 429 6700 493
rect 6764 481 6774 493
rect 7052 481 7086 621
rect 7244 481 7278 621
rect 7436 481 7470 621
rect 7628 481 7662 621
rect 7820 481 7854 621
rect 8012 481 8046 621
rect 6764 447 8046 481
rect 6764 429 6774 447
rect 6932 332 6978 344
rect -730 127 -720 179
rect -668 127 -641 179
rect 6932 132 6938 332
rect 6972 132 6978 332
rect 7052 316 7086 447
rect 7244 316 7278 447
rect 7436 316 7470 447
rect 7628 316 7662 447
rect 7820 316 7854 447
rect 8012 316 8046 447
rect 8196 481 8230 1044
rect 8270 934 8280 986
rect 8332 934 8359 986
rect 8724 481 8799 2247
rect 8196 447 8799 481
rect 7046 304 7092 316
rect 7046 222 7052 304
rect 7086 222 7092 304
rect 7046 210 7092 222
rect 7142 304 7188 316
rect 7142 222 7148 304
rect 7182 222 7188 304
rect 7142 210 7188 222
rect 7238 304 7284 316
rect 7238 222 7244 304
rect 7278 222 7284 304
rect 7238 210 7284 222
rect 7334 304 7380 316
rect 7334 222 7340 304
rect 7374 222 7380 304
rect 7334 210 7380 222
rect 7430 304 7476 316
rect 7430 222 7436 304
rect 7470 222 7476 304
rect 7430 210 7476 222
rect 7526 304 7572 316
rect 7526 222 7532 304
rect 7566 222 7572 304
rect 7526 210 7572 222
rect 7622 304 7668 316
rect 7622 222 7628 304
rect 7662 222 7668 304
rect 7622 210 7668 222
rect 7718 304 7764 316
rect 7718 222 7724 304
rect 7758 222 7764 304
rect 7718 210 7764 222
rect 7814 304 7860 316
rect 7814 222 7820 304
rect 7854 222 7860 304
rect 7814 210 7860 222
rect 7910 304 7956 316
rect 7910 222 7916 304
rect 7950 222 7956 304
rect 7910 210 7956 222
rect 8006 304 8052 316
rect 8006 222 8012 304
rect 8046 222 8052 304
rect 8006 210 8052 222
rect 7036 178 7102 182
rect -1852 36 -770 70
rect 6932 -40 6978 132
rect 7033 126 7043 178
rect 7095 126 7105 178
rect 7036 122 7102 126
rect 7148 70 7182 210
rect 7228 178 7294 182
rect 7225 126 7235 178
rect 7287 126 7297 178
rect 7228 122 7294 126
rect 7340 70 7374 210
rect 7420 179 7486 182
rect 7418 127 7428 179
rect 7480 127 7490 179
rect 7420 122 7486 127
rect 7532 70 7566 210
rect 7612 179 7678 182
rect 7610 127 7620 179
rect 7672 127 7682 179
rect 7612 122 7678 127
rect 7724 70 7758 210
rect 7804 179 7870 182
rect 7802 127 7812 179
rect 7864 127 7874 179
rect 7804 122 7870 127
rect 7916 70 7950 210
rect 7996 179 8062 182
rect 7993 127 8003 179
rect 8055 127 8065 179
rect 7996 122 8062 127
rect 8196 70 8230 447
rect 8270 127 8280 179
rect 8332 127 8359 179
rect 7148 36 8230 70
rect -2068 -818 -2022 -640
rect -1852 -756 -770 -722
rect -2068 -1204 -2062 -818
rect -2028 -1204 -2022 -818
rect -1967 -866 -1957 -814
rect -1905 -866 -1895 -814
rect -1852 -905 -1818 -756
rect -1775 -866 -1765 -814
rect -1713 -866 -1703 -814
rect -1660 -905 -1626 -756
rect -1583 -866 -1573 -814
rect -1521 -866 -1511 -814
rect -1468 -905 -1434 -756
rect -1391 -866 -1381 -814
rect -1329 -866 -1319 -814
rect -1276 -905 -1242 -756
rect -1200 -866 -1190 -814
rect -1138 -866 -1128 -814
rect -1084 -905 -1050 -756
rect -1007 -866 -997 -814
rect -945 -866 -935 -814
rect -1954 -917 -1908 -905
rect -1954 -1167 -1948 -917
rect -1914 -1167 -1908 -917
rect -1954 -1179 -1908 -1167
rect -1858 -917 -1812 -905
rect -1858 -1167 -1852 -917
rect -1818 -1167 -1812 -917
rect -1858 -1179 -1812 -1167
rect -1762 -917 -1716 -905
rect -1762 -1167 -1756 -917
rect -1722 -1167 -1716 -917
rect -1762 -1179 -1716 -1167
rect -1666 -917 -1620 -905
rect -1666 -1167 -1660 -917
rect -1626 -1167 -1620 -917
rect -1666 -1179 -1620 -1167
rect -1570 -917 -1524 -905
rect -1570 -1167 -1564 -917
rect -1530 -1167 -1524 -917
rect -1570 -1179 -1524 -1167
rect -1474 -917 -1428 -905
rect -1474 -1167 -1468 -917
rect -1434 -1167 -1428 -917
rect -1474 -1179 -1428 -1167
rect -1378 -917 -1332 -905
rect -1378 -1167 -1372 -917
rect -1338 -1167 -1332 -917
rect -1378 -1179 -1332 -1167
rect -1282 -917 -1236 -905
rect -1282 -1167 -1276 -917
rect -1242 -1167 -1236 -917
rect -1282 -1179 -1236 -1167
rect -1186 -917 -1140 -905
rect -1186 -1167 -1180 -917
rect -1146 -1167 -1140 -917
rect -1186 -1179 -1140 -1167
rect -1090 -917 -1044 -905
rect -1090 -1167 -1084 -917
rect -1050 -1167 -1044 -917
rect -1090 -1179 -1044 -1167
rect -994 -917 -948 -905
rect -994 -1167 -988 -917
rect -954 -1167 -948 -917
rect -994 -1179 -948 -1167
rect -2068 -1216 -2022 -1204
rect -1948 -1319 -1914 -1179
rect -1756 -1319 -1722 -1179
rect -1564 -1319 -1530 -1179
rect -1372 -1319 -1338 -1179
rect -1180 -1319 -1146 -1179
rect -988 -1304 -954 -1179
rect -1029 -1319 -1019 -1304
rect -3494 -1353 -1019 -1319
rect -2068 -1468 -2022 -1456
rect -2068 -1668 -2062 -1468
rect -2028 -1668 -2022 -1468
rect -1948 -1484 -1914 -1353
rect -1756 -1484 -1722 -1353
rect -1564 -1484 -1530 -1353
rect -1372 -1484 -1338 -1353
rect -1180 -1484 -1146 -1353
rect -1029 -1368 -1019 -1353
rect -955 -1368 -945 -1304
rect -804 -1319 -770 -756
rect -730 -866 -720 -814
rect -668 -866 -641 -814
rect 6932 -818 6978 -640
rect 7148 -756 8230 -722
rect 6932 -1204 6938 -818
rect 6972 -1204 6978 -818
rect 7033 -866 7043 -814
rect 7095 -866 7105 -814
rect 7148 -905 7182 -756
rect 7225 -866 7235 -814
rect 7287 -866 7297 -814
rect 7340 -905 7374 -756
rect 7417 -866 7427 -814
rect 7479 -866 7489 -814
rect 7532 -905 7566 -756
rect 7609 -866 7619 -814
rect 7671 -866 7681 -814
rect 7724 -905 7758 -756
rect 7800 -866 7810 -814
rect 7862 -866 7872 -814
rect 7916 -905 7950 -756
rect 7993 -866 8003 -814
rect 8055 -866 8065 -814
rect 7046 -917 7092 -905
rect 7046 -1167 7052 -917
rect 7086 -1167 7092 -917
rect 7046 -1179 7092 -1167
rect 7142 -917 7188 -905
rect 7142 -1167 7148 -917
rect 7182 -1167 7188 -917
rect 7142 -1179 7188 -1167
rect 7238 -917 7284 -905
rect 7238 -1167 7244 -917
rect 7278 -1167 7284 -917
rect 7238 -1179 7284 -1167
rect 7334 -917 7380 -905
rect 7334 -1167 7340 -917
rect 7374 -1167 7380 -917
rect 7334 -1179 7380 -1167
rect 7430 -917 7476 -905
rect 7430 -1167 7436 -917
rect 7470 -1167 7476 -917
rect 7430 -1179 7476 -1167
rect 7526 -917 7572 -905
rect 7526 -1167 7532 -917
rect 7566 -1167 7572 -917
rect 7526 -1179 7572 -1167
rect 7622 -917 7668 -905
rect 7622 -1167 7628 -917
rect 7662 -1167 7668 -917
rect 7622 -1179 7668 -1167
rect 7718 -917 7764 -905
rect 7718 -1167 7724 -917
rect 7758 -1167 7764 -917
rect 7718 -1179 7764 -1167
rect 7814 -917 7860 -905
rect 7814 -1167 7820 -917
rect 7854 -1167 7860 -917
rect 7814 -1179 7860 -1167
rect 7910 -917 7956 -905
rect 7910 -1167 7916 -917
rect 7950 -1167 7956 -917
rect 7910 -1179 7956 -1167
rect 8006 -917 8052 -905
rect 8006 -1167 8012 -917
rect 8046 -1167 8052 -917
rect 8006 -1179 8052 -1167
rect 6932 -1216 6978 -1204
rect -512 -1319 -502 -1301
rect -804 -1353 -502 -1319
rect -988 -1484 -954 -1368
rect -1954 -1496 -1908 -1484
rect -1954 -1578 -1948 -1496
rect -1914 -1578 -1908 -1496
rect -1954 -1590 -1908 -1578
rect -1858 -1496 -1812 -1484
rect -1858 -1578 -1852 -1496
rect -1818 -1578 -1812 -1496
rect -1858 -1590 -1812 -1578
rect -1762 -1496 -1716 -1484
rect -1762 -1578 -1756 -1496
rect -1722 -1578 -1716 -1496
rect -1762 -1590 -1716 -1578
rect -1666 -1496 -1620 -1484
rect -1666 -1578 -1660 -1496
rect -1626 -1578 -1620 -1496
rect -1666 -1590 -1620 -1578
rect -1570 -1496 -1524 -1484
rect -1570 -1578 -1564 -1496
rect -1530 -1578 -1524 -1496
rect -1570 -1590 -1524 -1578
rect -1474 -1496 -1428 -1484
rect -1474 -1578 -1468 -1496
rect -1434 -1578 -1428 -1496
rect -1474 -1590 -1428 -1578
rect -1378 -1496 -1332 -1484
rect -1378 -1578 -1372 -1496
rect -1338 -1578 -1332 -1496
rect -1378 -1590 -1332 -1578
rect -1282 -1496 -1236 -1484
rect -1282 -1578 -1276 -1496
rect -1242 -1578 -1236 -1496
rect -1282 -1590 -1236 -1578
rect -1186 -1496 -1140 -1484
rect -1186 -1578 -1180 -1496
rect -1146 -1578 -1140 -1496
rect -1186 -1590 -1140 -1578
rect -1090 -1496 -1044 -1484
rect -1090 -1578 -1084 -1496
rect -1050 -1578 -1044 -1496
rect -1090 -1590 -1044 -1578
rect -994 -1496 -948 -1484
rect -994 -1578 -988 -1496
rect -954 -1578 -948 -1496
rect -994 -1590 -948 -1578
rect -1964 -1622 -1898 -1618
rect -2068 -1840 -2022 -1668
rect -1967 -1674 -1957 -1622
rect -1905 -1674 -1895 -1622
rect -1964 -1678 -1898 -1674
rect -1852 -1730 -1818 -1590
rect -1772 -1622 -1706 -1618
rect -1775 -1674 -1765 -1622
rect -1713 -1674 -1703 -1622
rect -1772 -1678 -1706 -1674
rect -1660 -1730 -1626 -1590
rect -1580 -1621 -1514 -1618
rect -1582 -1673 -1572 -1621
rect -1520 -1673 -1510 -1621
rect -1580 -1678 -1514 -1673
rect -1468 -1730 -1434 -1590
rect -1388 -1621 -1322 -1618
rect -1390 -1673 -1380 -1621
rect -1328 -1673 -1318 -1621
rect -1388 -1678 -1322 -1673
rect -1276 -1730 -1242 -1590
rect -1196 -1621 -1130 -1618
rect -1198 -1673 -1188 -1621
rect -1136 -1673 -1126 -1621
rect -1196 -1678 -1130 -1673
rect -1084 -1730 -1050 -1590
rect -1004 -1621 -938 -1618
rect -1007 -1673 -997 -1621
rect -945 -1673 -935 -1621
rect -1004 -1678 -938 -1673
rect -804 -1730 -770 -1353
rect -512 -1365 -502 -1353
rect -438 -1365 -428 -1301
rect 6708 -1363 6718 -1299
rect 6782 -1319 6792 -1299
rect 7052 -1319 7086 -1179
rect 7244 -1319 7278 -1179
rect 7436 -1319 7470 -1179
rect 7628 -1319 7662 -1179
rect 7820 -1319 7854 -1179
rect 8012 -1319 8046 -1179
rect 6782 -1353 8046 -1319
rect 6782 -1363 6792 -1353
rect 6932 -1468 6978 -1456
rect -730 -1673 -720 -1621
rect -668 -1673 -641 -1621
rect 6932 -1668 6938 -1468
rect 6972 -1668 6978 -1468
rect 7052 -1484 7086 -1353
rect 7244 -1484 7278 -1353
rect 7436 -1484 7470 -1353
rect 7628 -1484 7662 -1353
rect 7820 -1484 7854 -1353
rect 8012 -1484 8046 -1353
rect 8196 -1319 8230 -756
rect 8270 -866 8280 -814
rect 8332 -866 8359 -814
rect 9235 -1319 9310 7647
rect 8196 -1353 9310 -1319
rect 7046 -1496 7092 -1484
rect 7046 -1578 7052 -1496
rect 7086 -1578 7092 -1496
rect 7046 -1590 7092 -1578
rect 7142 -1496 7188 -1484
rect 7142 -1578 7148 -1496
rect 7182 -1578 7188 -1496
rect 7142 -1590 7188 -1578
rect 7238 -1496 7284 -1484
rect 7238 -1578 7244 -1496
rect 7278 -1578 7284 -1496
rect 7238 -1590 7284 -1578
rect 7334 -1496 7380 -1484
rect 7334 -1578 7340 -1496
rect 7374 -1578 7380 -1496
rect 7334 -1590 7380 -1578
rect 7430 -1496 7476 -1484
rect 7430 -1578 7436 -1496
rect 7470 -1578 7476 -1496
rect 7430 -1590 7476 -1578
rect 7526 -1496 7572 -1484
rect 7526 -1578 7532 -1496
rect 7566 -1578 7572 -1496
rect 7526 -1590 7572 -1578
rect 7622 -1496 7668 -1484
rect 7622 -1578 7628 -1496
rect 7662 -1578 7668 -1496
rect 7622 -1590 7668 -1578
rect 7718 -1496 7764 -1484
rect 7718 -1578 7724 -1496
rect 7758 -1578 7764 -1496
rect 7718 -1590 7764 -1578
rect 7814 -1496 7860 -1484
rect 7814 -1578 7820 -1496
rect 7854 -1578 7860 -1496
rect 7814 -1590 7860 -1578
rect 7910 -1496 7956 -1484
rect 7910 -1578 7916 -1496
rect 7950 -1578 7956 -1496
rect 7910 -1590 7956 -1578
rect 8006 -1496 8052 -1484
rect 8006 -1578 8012 -1496
rect 8046 -1578 8052 -1496
rect 8006 -1590 8052 -1578
rect 7036 -1622 7102 -1618
rect -1852 -1764 -770 -1730
rect 6932 -1840 6978 -1668
rect 7033 -1674 7043 -1622
rect 7095 -1674 7105 -1622
rect 7036 -1678 7102 -1674
rect 7148 -1730 7182 -1590
rect 7228 -1622 7294 -1618
rect 7225 -1674 7235 -1622
rect 7287 -1674 7297 -1622
rect 7228 -1678 7294 -1674
rect 7340 -1730 7374 -1590
rect 7420 -1621 7486 -1618
rect 7418 -1673 7428 -1621
rect 7480 -1673 7490 -1621
rect 7420 -1678 7486 -1673
rect 7532 -1730 7566 -1590
rect 7612 -1621 7678 -1618
rect 7610 -1673 7620 -1621
rect 7672 -1673 7682 -1621
rect 7612 -1678 7678 -1673
rect 7724 -1730 7758 -1590
rect 7804 -1621 7870 -1618
rect 7802 -1673 7812 -1621
rect 7864 -1673 7874 -1621
rect 7804 -1678 7870 -1673
rect 7916 -1730 7950 -1590
rect 7996 -1621 8062 -1618
rect 7993 -1673 8003 -1621
rect 8055 -1673 8065 -1621
rect 7996 -1678 8062 -1673
rect 8196 -1730 8230 -1353
rect 8270 -1673 8280 -1621
rect 8332 -1673 8359 -1621
rect 7148 -1764 8230 -1730
<< via1 >>
rect -1957 8176 -1905 8186
rect -1957 8142 -1948 8176
rect -1948 8142 -1914 8176
rect -1914 8142 -1905 8176
rect -1957 8134 -1905 8142
rect -1765 8176 -1713 8186
rect -1765 8142 -1756 8176
rect -1756 8142 -1722 8176
rect -1722 8142 -1713 8176
rect -1765 8134 -1713 8142
rect -1573 8176 -1521 8186
rect -1573 8142 -1564 8176
rect -1564 8142 -1530 8176
rect -1530 8142 -1521 8176
rect -1573 8134 -1521 8142
rect -1381 8176 -1329 8186
rect -1381 8142 -1372 8176
rect -1372 8142 -1338 8176
rect -1338 8142 -1329 8176
rect -1381 8134 -1329 8142
rect -1190 8176 -1138 8186
rect -1190 8142 -1180 8176
rect -1180 8142 -1146 8176
rect -1146 8142 -1138 8176
rect -1190 8134 -1138 8142
rect -997 8176 -945 8186
rect -997 8142 -988 8176
rect -988 8142 -954 8176
rect -954 8142 -945 8176
rect -997 8134 -945 8142
rect -1022 7631 -958 7695
rect -720 8134 -668 8186
rect 7043 8176 7095 8186
rect 7043 8142 7052 8176
rect 7052 8142 7086 8176
rect 7086 8142 7095 8176
rect 7043 8134 7095 8142
rect 7235 8176 7287 8186
rect 7235 8142 7244 8176
rect 7244 8142 7278 8176
rect 7278 8142 7287 8176
rect 7235 8134 7287 8142
rect 7427 8176 7479 8186
rect 7427 8142 7436 8176
rect 7436 8142 7470 8176
rect 7470 8142 7479 8176
rect 7427 8134 7479 8142
rect 7619 8176 7671 8186
rect 7619 8142 7628 8176
rect 7628 8142 7662 8176
rect 7662 8142 7671 8176
rect 7619 8134 7671 8142
rect 7810 8176 7862 8186
rect 7810 8142 7820 8176
rect 7820 8142 7854 8176
rect 7854 8142 7862 8176
rect 7810 8134 7862 8142
rect 8003 8176 8055 8186
rect 8003 8142 8012 8176
rect 8012 8142 8046 8176
rect 8046 8142 8055 8176
rect 8003 8134 8055 8142
rect -1957 7369 -1905 7378
rect -1957 7335 -1948 7369
rect -1948 7335 -1914 7369
rect -1914 7335 -1905 7369
rect -1957 7326 -1905 7335
rect -1765 7369 -1713 7378
rect -1765 7335 -1756 7369
rect -1756 7335 -1722 7369
rect -1722 7335 -1713 7369
rect -1765 7326 -1713 7335
rect -1572 7369 -1520 7379
rect -1572 7335 -1564 7369
rect -1564 7335 -1530 7369
rect -1530 7335 -1520 7369
rect -1572 7327 -1520 7335
rect -1380 7369 -1328 7379
rect -1380 7335 -1372 7369
rect -1372 7335 -1338 7369
rect -1338 7335 -1328 7369
rect -1380 7327 -1328 7335
rect -1188 7369 -1136 7379
rect -1188 7335 -1180 7369
rect -1180 7335 -1146 7369
rect -1146 7335 -1136 7369
rect -1188 7327 -1136 7335
rect -997 7369 -945 7379
rect -997 7335 -988 7369
rect -988 7335 -954 7369
rect -954 7335 -945 7369
rect -997 7327 -945 7335
rect 6691 7633 6755 7697
rect -720 7327 -668 7379
rect -1957 6376 -1905 6386
rect -1957 6342 -1948 6376
rect -1948 6342 -1914 6376
rect -1914 6342 -1905 6376
rect -1957 6334 -1905 6342
rect -1765 6376 -1713 6386
rect -1765 6342 -1756 6376
rect -1756 6342 -1722 6376
rect -1722 6342 -1713 6376
rect -1765 6334 -1713 6342
rect -1573 6376 -1521 6386
rect -1573 6342 -1564 6376
rect -1564 6342 -1530 6376
rect -1530 6342 -1521 6376
rect -1573 6334 -1521 6342
rect -1381 6376 -1329 6386
rect -1381 6342 -1372 6376
rect -1372 6342 -1338 6376
rect -1338 6342 -1329 6376
rect -1381 6334 -1329 6342
rect -1190 6376 -1138 6386
rect -1190 6342 -1180 6376
rect -1180 6342 -1146 6376
rect -1146 6342 -1138 6376
rect -1190 6334 -1138 6342
rect -997 6376 -945 6386
rect -997 6342 -988 6376
rect -988 6342 -954 6376
rect -954 6342 -945 6376
rect -997 6334 -945 6342
rect -1028 5831 -964 5895
rect 1628 6412 1692 6476
rect -720 6334 -668 6386
rect -1957 5569 -1905 5578
rect -1957 5535 -1948 5569
rect -1948 5535 -1914 5569
rect -1914 5535 -1905 5569
rect -1957 5526 -1905 5535
rect -1765 5569 -1713 5578
rect -1765 5535 -1756 5569
rect -1756 5535 -1722 5569
rect -1722 5535 -1713 5569
rect -1765 5526 -1713 5535
rect -1572 5569 -1520 5579
rect -1572 5535 -1564 5569
rect -1564 5535 -1530 5569
rect -1530 5535 -1520 5569
rect -1572 5527 -1520 5535
rect -1380 5569 -1328 5579
rect -1380 5535 -1372 5569
rect -1372 5535 -1338 5569
rect -1338 5535 -1328 5569
rect -1380 5527 -1328 5535
rect -1188 5569 -1136 5579
rect -1188 5535 -1180 5569
rect -1180 5535 -1146 5569
rect -1146 5535 -1136 5569
rect -1188 5527 -1136 5535
rect -997 5569 -945 5579
rect -997 5535 -988 5569
rect -988 5535 -954 5569
rect -954 5535 -945 5569
rect -997 5527 -945 5535
rect -477 5829 -413 5893
rect -720 5527 -668 5579
rect -1957 4576 -1905 4586
rect -1957 4542 -1948 4576
rect -1948 4542 -1914 4576
rect -1914 4542 -1905 4576
rect -1957 4534 -1905 4542
rect -1765 4576 -1713 4586
rect -1765 4542 -1756 4576
rect -1756 4542 -1722 4576
rect -1722 4542 -1713 4576
rect -1765 4534 -1713 4542
rect -1573 4576 -1521 4586
rect -1573 4542 -1564 4576
rect -1564 4542 -1530 4576
rect -1530 4542 -1521 4576
rect -1573 4534 -1521 4542
rect -1381 4576 -1329 4586
rect -1381 4542 -1372 4576
rect -1372 4542 -1338 4576
rect -1338 4542 -1329 4576
rect -1381 4534 -1329 4542
rect -1190 4576 -1138 4586
rect -1190 4542 -1180 4576
rect -1180 4542 -1146 4576
rect -1146 4542 -1138 4576
rect -1190 4534 -1138 4542
rect -997 4576 -945 4586
rect -997 4542 -988 4576
rect -988 4542 -954 4576
rect -954 4542 -945 4576
rect -997 4534 -945 4542
rect -1024 4031 -960 4095
rect -720 4534 -668 4586
rect -1957 3769 -1905 3778
rect -1957 3735 -1948 3769
rect -1948 3735 -1914 3769
rect -1914 3735 -1905 3769
rect -1957 3726 -1905 3735
rect -1765 3769 -1713 3778
rect -1765 3735 -1756 3769
rect -1756 3735 -1722 3769
rect -1722 3735 -1713 3769
rect -1765 3726 -1713 3735
rect -1572 3769 -1520 3779
rect -1572 3735 -1564 3769
rect -1564 3735 -1530 3769
rect -1530 3735 -1520 3769
rect -1572 3727 -1520 3735
rect -1380 3769 -1328 3779
rect -1380 3735 -1372 3769
rect -1372 3735 -1338 3769
rect -1338 3735 -1328 3769
rect -1380 3727 -1328 3735
rect -1188 3769 -1136 3779
rect -1188 3735 -1180 3769
rect -1180 3735 -1146 3769
rect -1146 3735 -1136 3769
rect -1188 3727 -1136 3735
rect -997 3769 -945 3779
rect -997 3735 -988 3769
rect -988 3735 -954 3769
rect -954 3735 -945 3769
rect -997 3727 -945 3735
rect -434 4030 -370 4094
rect 8280 8134 8332 8186
rect 7043 7369 7095 7378
rect 7043 7335 7052 7369
rect 7052 7335 7086 7369
rect 7086 7335 7095 7369
rect 7043 7326 7095 7335
rect 7235 7369 7287 7378
rect 7235 7335 7244 7369
rect 7244 7335 7278 7369
rect 7278 7335 7287 7369
rect 7235 7326 7287 7335
rect 7428 7369 7480 7379
rect 7428 7335 7436 7369
rect 7436 7335 7470 7369
rect 7470 7335 7480 7369
rect 7428 7327 7480 7335
rect 7620 7369 7672 7379
rect 7620 7335 7628 7369
rect 7628 7335 7662 7369
rect 7662 7335 7672 7369
rect 7620 7327 7672 7335
rect 7812 7369 7864 7379
rect 7812 7335 7820 7369
rect 7820 7335 7854 7369
rect 7854 7335 7864 7369
rect 7812 7327 7864 7335
rect 8003 7369 8055 7379
rect 8003 7335 8012 7369
rect 8012 7335 8046 7369
rect 8046 7335 8055 7369
rect 8003 7327 8055 7335
rect 8280 7327 8332 7379
rect 7043 6376 7095 6386
rect 7043 6342 7052 6376
rect 7052 6342 7086 6376
rect 7086 6342 7095 6376
rect 7043 6334 7095 6342
rect 7235 6376 7287 6386
rect 7235 6342 7244 6376
rect 7244 6342 7278 6376
rect 7278 6342 7287 6376
rect 7235 6334 7287 6342
rect 7427 6376 7479 6386
rect 7427 6342 7436 6376
rect 7436 6342 7470 6376
rect 7470 6342 7479 6376
rect 7427 6334 7479 6342
rect 7619 6376 7671 6386
rect 7619 6342 7628 6376
rect 7628 6342 7662 6376
rect 7662 6342 7671 6376
rect 7619 6334 7671 6342
rect 7810 6376 7862 6386
rect 7810 6342 7820 6376
rect 7820 6342 7854 6376
rect 7854 6342 7862 6376
rect 7810 6334 7862 6342
rect 8003 6376 8055 6386
rect 8003 6342 8012 6376
rect 8012 6342 8046 6376
rect 8046 6342 8055 6376
rect 8003 6334 8055 6342
rect 6704 5831 6768 5895
rect 3157 5494 3221 5558
rect 8280 6334 8332 6386
rect 7043 5569 7095 5578
rect 7043 5535 7052 5569
rect 7052 5535 7086 5569
rect 7086 5535 7095 5569
rect 7043 5526 7095 5535
rect 7235 5569 7287 5578
rect 7235 5535 7244 5569
rect 7244 5535 7278 5569
rect 7278 5535 7287 5569
rect 7235 5526 7287 5535
rect 7428 5569 7480 5579
rect 7428 5535 7436 5569
rect 7436 5535 7470 5569
rect 7470 5535 7480 5569
rect 7428 5527 7480 5535
rect 7620 5569 7672 5579
rect 7620 5535 7628 5569
rect 7628 5535 7662 5569
rect 7662 5535 7672 5569
rect 7620 5527 7672 5535
rect 7812 5569 7864 5579
rect 7812 5535 7820 5569
rect 7820 5535 7854 5569
rect 7854 5535 7864 5569
rect 7812 5527 7864 5535
rect 8003 5569 8055 5579
rect 8003 5535 8012 5569
rect 8012 5535 8046 5569
rect 8046 5535 8055 5569
rect 8003 5527 8055 5535
rect 8280 5527 8332 5579
rect 3157 5020 3221 5084
rect 3768 4864 3832 4928
rect 6166 4868 6230 4932
rect 3106 4499 3170 4563
rect 5207 4326 5271 4390
rect 3308 4148 3372 4212
rect -720 3727 -668 3779
rect 333 3419 397 3483
rect 1631 3419 1695 3483
rect 333 3090 397 3154
rect -1957 2776 -1905 2786
rect -1957 2742 -1948 2776
rect -1948 2742 -1914 2776
rect -1914 2742 -1905 2776
rect -1957 2734 -1905 2742
rect -1765 2776 -1713 2786
rect -1765 2742 -1756 2776
rect -1756 2742 -1722 2776
rect -1722 2742 -1713 2776
rect -1765 2734 -1713 2742
rect -1573 2776 -1521 2786
rect -1573 2742 -1564 2776
rect -1564 2742 -1530 2776
rect -1530 2742 -1521 2776
rect -1573 2734 -1521 2742
rect -1381 2776 -1329 2786
rect -1381 2742 -1372 2776
rect -1372 2742 -1338 2776
rect -1338 2742 -1329 2776
rect -1381 2734 -1329 2742
rect -1190 2776 -1138 2786
rect -1190 2742 -1180 2776
rect -1180 2742 -1146 2776
rect -1146 2742 -1138 2776
rect -1190 2734 -1138 2742
rect -997 2776 -945 2786
rect -997 2742 -988 2776
rect -988 2742 -954 2776
rect -954 2742 -945 2776
rect -997 2734 -945 2742
rect -1027 2231 -963 2295
rect -720 2734 -668 2786
rect -1957 1969 -1905 1978
rect -1957 1935 -1948 1969
rect -1948 1935 -1914 1969
rect -1914 1935 -1905 1969
rect -1957 1926 -1905 1935
rect -1765 1969 -1713 1978
rect -1765 1935 -1756 1969
rect -1756 1935 -1722 1969
rect -1722 1935 -1713 1969
rect -1765 1926 -1713 1935
rect -1572 1969 -1520 1979
rect -1572 1935 -1564 1969
rect -1564 1935 -1530 1969
rect -1530 1935 -1520 1969
rect -1572 1927 -1520 1935
rect -1380 1969 -1328 1979
rect -1380 1935 -1372 1969
rect -1372 1935 -1338 1969
rect -1338 1935 -1328 1969
rect -1380 1927 -1328 1935
rect -1188 1969 -1136 1979
rect -1188 1935 -1180 1969
rect -1180 1935 -1146 1969
rect -1146 1935 -1136 1969
rect -1188 1927 -1136 1935
rect -997 1969 -945 1979
rect -997 1935 -988 1969
rect -988 1935 -954 1969
rect -954 1935 -945 1969
rect -997 1927 -945 1935
rect -434 2227 -370 2291
rect 7043 4576 7095 4586
rect 7043 4542 7052 4576
rect 7052 4542 7086 4576
rect 7086 4542 7095 4576
rect 7043 4534 7095 4542
rect 7235 4576 7287 4586
rect 7235 4542 7244 4576
rect 7244 4542 7278 4576
rect 7278 4542 7287 4576
rect 7235 4534 7287 4542
rect 7427 4576 7479 4586
rect 7427 4542 7436 4576
rect 7436 4542 7470 4576
rect 7470 4542 7479 4576
rect 7427 4534 7479 4542
rect 7619 4576 7671 4586
rect 7619 4542 7628 4576
rect 7628 4542 7662 4576
rect 7662 4542 7671 4576
rect 7619 4534 7671 4542
rect 7810 4576 7862 4586
rect 7810 4542 7820 4576
rect 7820 4542 7854 4576
rect 7854 4542 7862 4576
rect 7810 4534 7862 4542
rect 8003 4576 8055 4586
rect 8003 4542 8012 4576
rect 8012 4542 8046 4576
rect 8046 4542 8055 4576
rect 8003 4534 8055 4542
rect 6759 4031 6823 4095
rect 8280 4534 8332 4586
rect 4874 3578 4938 3642
rect 7043 3769 7095 3778
rect 7043 3735 7052 3769
rect 7052 3735 7086 3769
rect 7086 3735 7095 3769
rect 7043 3726 7095 3735
rect 7235 3769 7287 3778
rect 7235 3735 7244 3769
rect 7244 3735 7278 3769
rect 7278 3735 7287 3769
rect 7235 3726 7287 3735
rect 7428 3769 7480 3779
rect 7428 3735 7436 3769
rect 7436 3735 7470 3769
rect 7470 3735 7480 3769
rect 7428 3727 7480 3735
rect 7620 3769 7672 3779
rect 7620 3735 7628 3769
rect 7628 3735 7662 3769
rect 7662 3735 7672 3769
rect 7620 3727 7672 3735
rect 7812 3769 7864 3779
rect 7812 3735 7820 3769
rect 7820 3735 7854 3769
rect 7854 3735 7864 3769
rect 7812 3727 7864 3735
rect 8003 3769 8055 3779
rect 8003 3735 8012 3769
rect 8012 3735 8046 3769
rect 8046 3735 8055 3769
rect 8003 3727 8055 3735
rect 8280 3727 8332 3779
rect 7043 2776 7095 2786
rect 7043 2742 7052 2776
rect 7052 2742 7086 2776
rect 7086 2742 7095 2776
rect 7043 2734 7095 2742
rect 7235 2776 7287 2786
rect 7235 2742 7244 2776
rect 7244 2742 7278 2776
rect 7278 2742 7287 2776
rect 7235 2734 7287 2742
rect 7427 2776 7479 2786
rect 7427 2742 7436 2776
rect 7436 2742 7470 2776
rect 7470 2742 7479 2776
rect 7427 2734 7479 2742
rect 7619 2776 7671 2786
rect 7619 2742 7628 2776
rect 7628 2742 7662 2776
rect 7662 2742 7671 2776
rect 7619 2734 7671 2742
rect 7810 2776 7862 2786
rect 7810 2742 7820 2776
rect 7820 2742 7854 2776
rect 7854 2742 7862 2776
rect 7810 2734 7862 2742
rect 8003 2776 8055 2786
rect 8003 2742 8012 2776
rect 8012 2742 8046 2776
rect 8046 2742 8055 2776
rect 8003 2734 8055 2742
rect 6764 2233 6828 2297
rect 3308 2159 3372 2223
rect -720 1927 -668 1979
rect 8280 2734 8332 2786
rect 7043 1969 7095 1978
rect 7043 1935 7052 1969
rect 7052 1935 7086 1969
rect 7086 1935 7095 1969
rect 7043 1926 7095 1935
rect 7235 1969 7287 1978
rect 7235 1935 7244 1969
rect 7244 1935 7278 1969
rect 7278 1935 7287 1969
rect 7235 1926 7287 1935
rect 7428 1969 7480 1979
rect 7428 1935 7436 1969
rect 7436 1935 7470 1969
rect 7470 1935 7480 1969
rect 7428 1927 7480 1935
rect 7620 1969 7672 1979
rect 7620 1935 7628 1969
rect 7628 1935 7662 1969
rect 7662 1935 7672 1969
rect 7620 1927 7672 1935
rect 7812 1969 7864 1979
rect 7812 1935 7820 1969
rect 7820 1935 7854 1969
rect 7854 1935 7864 1969
rect 7812 1927 7864 1935
rect 8003 1969 8055 1979
rect 8003 1935 8012 1969
rect 8012 1935 8046 1969
rect 8046 1935 8055 1969
rect 8003 1927 8055 1935
rect 8280 1927 8332 1979
rect 2330 1576 2394 1640
rect -1957 976 -1905 986
rect -1957 942 -1948 976
rect -1948 942 -1914 976
rect -1914 942 -1905 976
rect -1957 934 -1905 942
rect -1765 976 -1713 986
rect -1765 942 -1756 976
rect -1756 942 -1722 976
rect -1722 942 -1713 976
rect -1765 934 -1713 942
rect -1573 976 -1521 986
rect -1573 942 -1564 976
rect -1564 942 -1530 976
rect -1530 942 -1521 976
rect -1573 934 -1521 942
rect -1381 976 -1329 986
rect -1381 942 -1372 976
rect -1372 942 -1338 976
rect -1338 942 -1329 976
rect -1381 934 -1329 942
rect -1190 976 -1138 986
rect -1190 942 -1180 976
rect -1180 942 -1146 976
rect -1146 942 -1138 976
rect -1190 934 -1138 942
rect -997 976 -945 986
rect -997 942 -988 976
rect -988 942 -954 976
rect -954 942 -945 976
rect -997 934 -945 942
rect -1020 433 -956 497
rect -720 934 -668 986
rect 3602 1462 3666 1526
rect 6152 1462 6216 1526
rect 170 1277 234 1341
rect 4326 1277 4390 1341
rect 7043 976 7095 986
rect 7043 942 7052 976
rect 7052 942 7086 976
rect 7086 942 7095 976
rect 7043 934 7095 942
rect 7235 976 7287 986
rect 7235 942 7244 976
rect 7244 942 7278 976
rect 7278 942 7287 976
rect 7235 934 7287 942
rect 7427 976 7479 986
rect 7427 942 7436 976
rect 7436 942 7470 976
rect 7470 942 7479 976
rect 7427 934 7479 942
rect 7619 976 7671 986
rect 7619 942 7628 976
rect 7628 942 7662 976
rect 7662 942 7671 976
rect 7619 934 7671 942
rect 7810 976 7862 986
rect 7810 942 7820 976
rect 7820 942 7854 976
rect 7854 942 7862 976
rect 7810 934 7862 942
rect 8003 976 8055 986
rect 8003 942 8012 976
rect 8012 942 8046 976
rect 8046 942 8055 976
rect 8003 934 8055 942
rect -1957 169 -1905 178
rect -1957 135 -1948 169
rect -1948 135 -1914 169
rect -1914 135 -1905 169
rect -1957 126 -1905 135
rect -1765 169 -1713 178
rect -1765 135 -1756 169
rect -1756 135 -1722 169
rect -1722 135 -1713 169
rect -1765 126 -1713 135
rect -1572 169 -1520 179
rect -1572 135 -1564 169
rect -1564 135 -1530 169
rect -1530 135 -1520 169
rect -1572 127 -1520 135
rect -1380 169 -1328 179
rect -1380 135 -1372 169
rect -1372 135 -1338 169
rect -1338 135 -1328 169
rect -1380 127 -1328 135
rect -1188 169 -1136 179
rect -1188 135 -1180 169
rect -1180 135 -1146 169
rect -1146 135 -1136 169
rect -1188 127 -1136 135
rect -997 169 -945 179
rect -997 135 -988 169
rect -988 135 -954 169
rect -954 135 -945 169
rect -997 127 -945 135
rect 6700 429 6764 493
rect -720 127 -668 179
rect 8280 934 8332 986
rect 7043 169 7095 178
rect 7043 135 7052 169
rect 7052 135 7086 169
rect 7086 135 7095 169
rect 7043 126 7095 135
rect 7235 169 7287 178
rect 7235 135 7244 169
rect 7244 135 7278 169
rect 7278 135 7287 169
rect 7235 126 7287 135
rect 7428 169 7480 179
rect 7428 135 7436 169
rect 7436 135 7470 169
rect 7470 135 7480 169
rect 7428 127 7480 135
rect 7620 169 7672 179
rect 7620 135 7628 169
rect 7628 135 7662 169
rect 7662 135 7672 169
rect 7620 127 7672 135
rect 7812 169 7864 179
rect 7812 135 7820 169
rect 7820 135 7854 169
rect 7854 135 7864 169
rect 7812 127 7864 135
rect 8003 169 8055 179
rect 8003 135 8012 169
rect 8012 135 8046 169
rect 8046 135 8055 169
rect 8003 127 8055 135
rect 8280 127 8332 179
rect -1957 -824 -1905 -814
rect -1957 -858 -1948 -824
rect -1948 -858 -1914 -824
rect -1914 -858 -1905 -824
rect -1957 -866 -1905 -858
rect -1765 -824 -1713 -814
rect -1765 -858 -1756 -824
rect -1756 -858 -1722 -824
rect -1722 -858 -1713 -824
rect -1765 -866 -1713 -858
rect -1573 -824 -1521 -814
rect -1573 -858 -1564 -824
rect -1564 -858 -1530 -824
rect -1530 -858 -1521 -824
rect -1573 -866 -1521 -858
rect -1381 -824 -1329 -814
rect -1381 -858 -1372 -824
rect -1372 -858 -1338 -824
rect -1338 -858 -1329 -824
rect -1381 -866 -1329 -858
rect -1190 -824 -1138 -814
rect -1190 -858 -1180 -824
rect -1180 -858 -1146 -824
rect -1146 -858 -1138 -824
rect -1190 -866 -1138 -858
rect -997 -824 -945 -814
rect -997 -858 -988 -824
rect -988 -858 -954 -824
rect -954 -858 -945 -824
rect -997 -866 -945 -858
rect -1019 -1368 -955 -1304
rect -720 -866 -668 -814
rect 7043 -824 7095 -814
rect 7043 -858 7052 -824
rect 7052 -858 7086 -824
rect 7086 -858 7095 -824
rect 7043 -866 7095 -858
rect 7235 -824 7287 -814
rect 7235 -858 7244 -824
rect 7244 -858 7278 -824
rect 7278 -858 7287 -824
rect 7235 -866 7287 -858
rect 7427 -824 7479 -814
rect 7427 -858 7436 -824
rect 7436 -858 7470 -824
rect 7470 -858 7479 -824
rect 7427 -866 7479 -858
rect 7619 -824 7671 -814
rect 7619 -858 7628 -824
rect 7628 -858 7662 -824
rect 7662 -858 7671 -824
rect 7619 -866 7671 -858
rect 7810 -824 7862 -814
rect 7810 -858 7820 -824
rect 7820 -858 7854 -824
rect 7854 -858 7862 -824
rect 7810 -866 7862 -858
rect 8003 -824 8055 -814
rect 8003 -858 8012 -824
rect 8012 -858 8046 -824
rect 8046 -858 8055 -824
rect 8003 -866 8055 -858
rect -1957 -1631 -1905 -1622
rect -1957 -1665 -1948 -1631
rect -1948 -1665 -1914 -1631
rect -1914 -1665 -1905 -1631
rect -1957 -1674 -1905 -1665
rect -1765 -1631 -1713 -1622
rect -1765 -1665 -1756 -1631
rect -1756 -1665 -1722 -1631
rect -1722 -1665 -1713 -1631
rect -1765 -1674 -1713 -1665
rect -1572 -1631 -1520 -1621
rect -1572 -1665 -1564 -1631
rect -1564 -1665 -1530 -1631
rect -1530 -1665 -1520 -1631
rect -1572 -1673 -1520 -1665
rect -1380 -1631 -1328 -1621
rect -1380 -1665 -1372 -1631
rect -1372 -1665 -1338 -1631
rect -1338 -1665 -1328 -1631
rect -1380 -1673 -1328 -1665
rect -1188 -1631 -1136 -1621
rect -1188 -1665 -1180 -1631
rect -1180 -1665 -1146 -1631
rect -1146 -1665 -1136 -1631
rect -1188 -1673 -1136 -1665
rect -997 -1631 -945 -1621
rect -997 -1665 -988 -1631
rect -988 -1665 -954 -1631
rect -954 -1665 -945 -1631
rect -997 -1673 -945 -1665
rect -502 -1365 -438 -1301
rect 6718 -1363 6782 -1299
rect -720 -1673 -668 -1621
rect 8280 -866 8332 -814
rect 7043 -1631 7095 -1622
rect 7043 -1665 7052 -1631
rect 7052 -1665 7086 -1631
rect 7086 -1665 7095 -1631
rect 7043 -1674 7095 -1665
rect 7235 -1631 7287 -1622
rect 7235 -1665 7244 -1631
rect 7244 -1665 7278 -1631
rect 7278 -1665 7287 -1631
rect 7235 -1674 7287 -1665
rect 7428 -1631 7480 -1621
rect 7428 -1665 7436 -1631
rect 7436 -1665 7470 -1631
rect 7470 -1665 7480 -1631
rect 7428 -1673 7480 -1665
rect 7620 -1631 7672 -1621
rect 7620 -1665 7628 -1631
rect 7628 -1665 7662 -1631
rect 7662 -1665 7672 -1631
rect 7620 -1673 7672 -1665
rect 7812 -1631 7864 -1621
rect 7812 -1665 7820 -1631
rect 7820 -1665 7854 -1631
rect 7854 -1665 7864 -1631
rect 7812 -1673 7864 -1665
rect 8003 -1631 8055 -1621
rect 8003 -1665 8012 -1631
rect 8012 -1665 8046 -1631
rect 8046 -1665 8055 -1631
rect 8003 -1673 8055 -1665
rect 8280 -1673 8332 -1621
<< metal2 >>
rect -2651 8198 -2587 8208
rect 8848 8198 8912 8208
rect -1957 8186 -1905 8196
rect -1765 8186 -1713 8196
rect -1573 8186 -1521 8196
rect -1381 8186 -1329 8196
rect -1190 8186 -1138 8196
rect -997 8186 -945 8196
rect -720 8186 -668 8196
rect 7043 8186 7095 8196
rect 7235 8186 7287 8196
rect 7427 8186 7479 8196
rect 7619 8186 7671 8196
rect 7810 8186 7862 8196
rect 8003 8186 8055 8196
rect 8280 8186 8332 8196
rect -2587 8134 -1957 8186
rect -1905 8134 -1765 8186
rect -1713 8134 -1573 8186
rect -1521 8134 -1381 8186
rect -1329 8134 -1190 8186
rect -1138 8134 -997 8186
rect -945 8134 -720 8186
rect 7036 8134 7043 8186
rect 7095 8134 7235 8186
rect 7287 8134 7427 8186
rect 7479 8134 7619 8186
rect 7671 8134 7810 8186
rect 7862 8134 8003 8186
rect 8055 8134 8280 8186
rect 8332 8134 8848 8186
rect -2651 8124 -2587 8134
rect -1957 8124 -1905 8134
rect -1765 8124 -1713 8134
rect -1573 8124 -1521 8134
rect -1381 8124 -1329 8134
rect -1190 8124 -1138 8134
rect -997 8124 -945 8134
rect -720 8124 -668 8134
rect 7043 8124 7095 8134
rect 7235 8124 7287 8134
rect 7427 8124 7479 8134
rect 7619 8124 7671 8134
rect 7810 8124 7862 8134
rect 8003 8124 8055 8134
rect 8280 8124 8332 8134
rect 8848 8124 8912 8134
rect -1022 7855 2060 7919
rect -1022 7695 -958 7855
rect -1022 7621 -958 7631
rect -2398 7390 -2334 7400
rect -1957 7379 -1905 7388
rect -1765 7379 -1713 7388
rect -1572 7379 -1520 7389
rect -1380 7379 -1328 7389
rect -1188 7379 -1136 7389
rect -997 7379 -945 7389
rect -720 7379 -668 7389
rect -1964 7378 -1572 7379
rect -2334 7326 -1957 7378
rect -1905 7327 -1765 7378
rect -2398 7316 -2334 7326
rect -1957 7316 -1905 7326
rect -1713 7327 -1572 7378
rect -1520 7327 -1380 7379
rect -1328 7327 -1188 7379
rect -1136 7327 -997 7379
rect -945 7327 -720 7379
rect -1765 7316 -1713 7326
rect -1572 7317 -1520 7327
rect -1380 7317 -1328 7327
rect -1188 7317 -1136 7327
rect -997 7317 -945 7327
rect -720 7317 -668 7327
rect 1996 6756 2060 7855
rect 6691 7697 6755 7707
rect 6691 7623 6755 7633
rect 8595 7391 8659 7401
rect 7043 7379 7095 7388
rect 7235 7379 7287 7388
rect 7428 7379 7480 7389
rect 7620 7379 7672 7389
rect 7812 7379 7864 7389
rect 8003 7379 8055 7389
rect 8280 7379 8332 7389
rect 7036 7378 7428 7379
rect 7036 7327 7043 7378
rect 7095 7327 7235 7378
rect 7043 7316 7095 7326
rect 7287 7327 7428 7378
rect 7480 7327 7620 7379
rect 7672 7327 7812 7379
rect 7864 7327 8003 7379
rect 8055 7327 8280 7379
rect 8332 7327 8595 7379
rect 7235 7316 7287 7326
rect 7428 7317 7480 7327
rect 7620 7317 7672 7327
rect 7812 7317 7864 7327
rect 8003 7317 8055 7327
rect 8280 7317 8332 7327
rect 8595 7317 8659 7327
rect 1996 6682 2060 6692
rect 1628 6476 1692 6486
rect -2651 6398 -2587 6408
rect 1628 6402 1692 6412
rect 8848 6398 8912 6408
rect -1957 6386 -1905 6396
rect -1765 6386 -1713 6396
rect -1573 6386 -1521 6396
rect -1381 6386 -1329 6396
rect -1190 6386 -1138 6396
rect -997 6386 -945 6396
rect -720 6386 -668 6396
rect 7043 6386 7095 6396
rect 7235 6386 7287 6396
rect 7427 6386 7479 6396
rect 7619 6386 7671 6396
rect 7810 6386 7862 6396
rect 8003 6386 8055 6396
rect 8280 6386 8332 6396
rect -2587 6334 -1957 6386
rect -1905 6334 -1765 6386
rect -1713 6334 -1573 6386
rect -1521 6334 -1381 6386
rect -1329 6334 -1190 6386
rect -1138 6334 -997 6386
rect -945 6334 -720 6386
rect 7036 6334 7043 6386
rect 7095 6334 7235 6386
rect 7287 6334 7427 6386
rect 7479 6334 7619 6386
rect 7671 6334 7810 6386
rect 7862 6334 8003 6386
rect 8055 6334 8280 6386
rect 8332 6334 8848 6386
rect -2651 6324 -2587 6334
rect -1957 6324 -1905 6334
rect -1765 6324 -1713 6334
rect -1573 6324 -1521 6334
rect -1381 6324 -1329 6334
rect -1190 6324 -1138 6334
rect -997 6324 -945 6334
rect -720 6324 -668 6334
rect 7043 6324 7095 6334
rect 7235 6324 7287 6334
rect 7427 6324 7479 6334
rect 7619 6324 7671 6334
rect 7810 6324 7862 6334
rect 8003 6324 8055 6334
rect 8280 6324 8332 6334
rect 8848 6324 8912 6334
rect -1028 5895 -964 5905
rect -1028 5726 -964 5831
rect -477 5893 -413 5903
rect -477 5819 -413 5829
rect 6704 5895 6768 5905
rect 6704 5821 6768 5831
rect 3410 5781 3474 5791
rect -1028 5662 -133 5726
rect -2398 5590 -2334 5600
rect -1957 5579 -1905 5588
rect -1765 5579 -1713 5588
rect -1572 5579 -1520 5589
rect -1380 5579 -1328 5589
rect -1188 5579 -1136 5589
rect -997 5579 -945 5589
rect -720 5579 -668 5589
rect -1964 5578 -1572 5579
rect -2334 5526 -1957 5578
rect -1905 5527 -1765 5578
rect -2398 5516 -2334 5526
rect -1957 5516 -1905 5526
rect -1713 5527 -1572 5578
rect -1520 5527 -1380 5579
rect -1328 5527 -1188 5579
rect -1136 5527 -997 5579
rect -945 5527 -720 5579
rect -1765 5516 -1713 5526
rect -1572 5517 -1520 5527
rect -1380 5517 -1328 5527
rect -1188 5517 -1136 5527
rect -997 5517 -945 5527
rect -720 5517 -668 5527
rect -197 5170 -133 5662
rect -197 5096 -133 5106
rect 1282 5612 1346 5622
rect -2651 4598 -2587 4608
rect -1957 4586 -1905 4596
rect -1765 4586 -1713 4596
rect -1573 4586 -1521 4596
rect -1381 4586 -1329 4596
rect -1190 4586 -1138 4596
rect -997 4586 -945 4596
rect -720 4586 -668 4596
rect -2587 4534 -1957 4586
rect -1905 4534 -1765 4586
rect -1713 4534 -1573 4586
rect -1521 4534 -1381 4586
rect -1329 4534 -1190 4586
rect -1138 4534 -997 4586
rect -945 4534 -720 4586
rect -2651 4524 -2587 4534
rect -1957 4524 -1905 4534
rect -1765 4524 -1713 4534
rect -1573 4524 -1521 4534
rect -1381 4524 -1329 4534
rect -1190 4524 -1138 4534
rect -997 4524 -945 4534
rect -720 4524 -668 4534
rect 1282 4219 1346 5548
rect 1630 5613 1694 5623
rect 1428 4219 1492 4229
rect -434 4155 1428 4219
rect -1024 4095 -960 4105
rect -1024 3923 -960 4031
rect -434 4094 -370 4155
rect 1428 4145 1492 4155
rect -434 4020 -370 4030
rect -1024 3859 -369 3923
rect -2398 3790 -2334 3800
rect -1957 3779 -1905 3788
rect -1765 3779 -1713 3788
rect -1572 3779 -1520 3789
rect -1380 3779 -1328 3789
rect -1188 3779 -1136 3789
rect -997 3779 -945 3789
rect -720 3779 -668 3789
rect -1964 3778 -1572 3779
rect -2334 3726 -1957 3778
rect -1905 3727 -1765 3778
rect -2398 3716 -2334 3726
rect -1957 3716 -1905 3726
rect -1713 3727 -1572 3778
rect -1520 3727 -1380 3779
rect -1328 3727 -1188 3779
rect -1136 3727 -997 3779
rect -945 3727 -720 3779
rect -1765 3716 -1713 3726
rect -1572 3717 -1520 3727
rect -1380 3717 -1328 3727
rect -1188 3717 -1136 3727
rect -997 3717 -945 3727
rect -720 3717 -668 3727
rect -433 3327 -369 3859
rect 1630 3843 1694 5549
rect 3157 5558 3221 5568
rect 3157 5484 3221 5494
rect 3410 5169 3474 5717
rect 8595 5591 8659 5601
rect 7043 5579 7095 5588
rect 7235 5579 7287 5588
rect 7428 5579 7480 5589
rect 7620 5579 7672 5589
rect 7812 5579 7864 5589
rect 8003 5579 8055 5589
rect 8280 5579 8332 5589
rect 7036 5578 7428 5579
rect 7036 5527 7043 5578
rect 7095 5527 7235 5578
rect 7043 5516 7095 5526
rect 7287 5527 7428 5578
rect 7480 5527 7620 5579
rect 7672 5527 7812 5579
rect 7864 5527 8003 5579
rect 8055 5527 8280 5579
rect 8332 5527 8595 5579
rect 7235 5516 7287 5526
rect 7428 5517 7480 5527
rect 7620 5517 7672 5527
rect 7812 5517 7864 5527
rect 8003 5517 8055 5527
rect 8280 5517 8332 5527
rect 8595 5517 8659 5527
rect 3410 5095 3474 5105
rect 4658 5106 4722 5116
rect 5418 5106 5482 5116
rect 3157 5084 3221 5094
rect 4722 5042 5418 5106
rect 4658 5032 4722 5042
rect 5418 5032 5482 5042
rect 3157 5010 3221 5020
rect 3768 4928 3832 4938
rect 3768 4854 3832 4864
rect 4084 4928 4148 4938
rect 5706 4928 5770 4938
rect 4148 4864 5706 4928
rect 4084 4854 4148 4864
rect 5706 4854 5770 4864
rect 6166 4932 6230 4942
rect 6166 4858 6230 4868
rect 8848 4598 8912 4608
rect 7043 4586 7095 4596
rect 7235 4586 7287 4596
rect 7427 4586 7479 4596
rect 7619 4586 7671 4596
rect 7810 4586 7862 4596
rect 8003 4586 8055 4596
rect 8280 4586 8332 4596
rect 3106 4563 3170 4573
rect 7036 4534 7043 4586
rect 7095 4534 7235 4586
rect 7287 4534 7427 4586
rect 7479 4534 7619 4586
rect 7671 4534 7810 4586
rect 7862 4534 8003 4586
rect 8055 4534 8280 4586
rect 8332 4534 8848 4586
rect 7043 4524 7095 4534
rect 7235 4524 7287 4534
rect 7427 4524 7479 4534
rect 7619 4524 7671 4534
rect 7810 4524 7862 4534
rect 8003 4524 8055 4534
rect 8280 4524 8332 4534
rect 8848 4524 8912 4534
rect 3106 4489 3170 4499
rect 5207 4390 5271 4400
rect 5207 4316 5271 4326
rect 3308 4212 3372 4222
rect 3308 4138 3372 4148
rect 6759 4095 6823 4105
rect 5952 4031 6759 4095
rect 4876 3980 4940 3990
rect 5206 3980 5270 3990
rect 4940 3916 5206 3980
rect 4876 3906 4940 3916
rect 5206 3906 5270 3916
rect 3306 3862 3370 3872
rect 1630 3779 1866 3843
rect 333 3483 397 3493
rect 333 3409 397 3419
rect 765 3483 829 3493
rect 1408 3483 1472 3493
rect 829 3419 1408 3483
rect 765 3409 829 3419
rect 1408 3409 1472 3419
rect 1631 3483 1695 3493
rect 1631 3409 1695 3419
rect 333 3327 397 3337
rect -433 3307 333 3327
rect -434 3263 333 3307
rect 397 3263 402 3327
rect -2651 2798 -2587 2808
rect -1957 2786 -1905 2796
rect -1765 2786 -1713 2796
rect -1573 2786 -1521 2796
rect -1381 2786 -1329 2796
rect -1190 2786 -1138 2796
rect -997 2786 -945 2796
rect -720 2786 -668 2796
rect -2587 2734 -1957 2786
rect -1905 2734 -1765 2786
rect -1713 2734 -1573 2786
rect -1521 2734 -1381 2786
rect -1329 2734 -1190 2786
rect -1138 2734 -997 2786
rect -945 2734 -720 2786
rect -2651 2724 -2587 2734
rect -1957 2724 -1905 2734
rect -1765 2724 -1713 2734
rect -1573 2724 -1521 2734
rect -1381 2724 -1329 2734
rect -1190 2724 -1138 2734
rect -997 2724 -945 2734
rect -720 2724 -668 2734
rect -434 2536 -370 3263
rect 333 3253 397 3263
rect 333 3154 397 3164
rect 333 3080 397 3090
rect 764 3153 828 3163
rect 1802 3153 1866 3779
rect 828 3089 1866 3153
rect 764 3079 828 3089
rect 3306 2623 3370 3798
rect 4874 3642 4938 3652
rect 4874 3568 4938 3578
rect 4510 3462 4574 3472
rect 5952 3462 6016 4031
rect 6759 4021 6823 4031
rect 8595 3791 8659 3801
rect 7043 3779 7095 3788
rect 7235 3779 7287 3788
rect 7428 3779 7480 3789
rect 7620 3779 7672 3789
rect 7812 3779 7864 3789
rect 8003 3779 8055 3789
rect 8280 3779 8332 3789
rect 7036 3778 7428 3779
rect 7036 3727 7043 3778
rect 7095 3727 7235 3778
rect 7043 3716 7095 3726
rect 7287 3727 7428 3778
rect 7480 3727 7620 3779
rect 7672 3727 7812 3779
rect 7864 3727 8003 3779
rect 8055 3727 8280 3779
rect 8332 3727 8595 3779
rect 7235 3716 7287 3726
rect 7428 3717 7480 3727
rect 7620 3717 7672 3727
rect 7812 3717 7864 3727
rect 8003 3717 8055 3727
rect 8280 3717 8332 3727
rect 8595 3717 8659 3727
rect 4574 3398 6016 3462
rect 4510 3388 4574 3398
rect 4508 3151 4572 3161
rect 4572 3087 6011 3151
rect 4508 3077 4572 3087
rect 3306 2549 3370 2559
rect -1027 2472 -370 2536
rect -1027 2295 -963 2472
rect -1027 2221 -963 2231
rect -434 2291 -370 2301
rect 5947 2297 6011 3087
rect 8848 2798 8912 2808
rect 7043 2786 7095 2796
rect 7235 2786 7287 2796
rect 7427 2786 7479 2796
rect 7619 2786 7671 2796
rect 7810 2786 7862 2796
rect 8003 2786 8055 2796
rect 8280 2786 8332 2796
rect 7036 2734 7043 2786
rect 7095 2734 7235 2786
rect 7287 2734 7427 2786
rect 7479 2734 7619 2786
rect 7671 2734 7810 2786
rect 7862 2734 8003 2786
rect 8055 2734 8280 2786
rect 8332 2734 8848 2786
rect 7043 2724 7095 2734
rect 7235 2724 7287 2734
rect 7427 2724 7479 2734
rect 7619 2724 7671 2734
rect 7810 2724 7862 2734
rect 8003 2724 8055 2734
rect 8280 2724 8332 2734
rect 8848 2724 8912 2734
rect 6764 2297 6828 2307
rect 5947 2233 6764 2297
rect -2398 1990 -2334 2000
rect -1957 1979 -1905 1988
rect -1765 1979 -1713 1988
rect -1572 1979 -1520 1989
rect -1380 1979 -1328 1989
rect -1188 1979 -1136 1989
rect -997 1979 -945 1989
rect -720 1979 -668 1989
rect -1964 1978 -1572 1979
rect -2334 1926 -1957 1978
rect -1905 1927 -1765 1978
rect -2398 1916 -2334 1926
rect -1957 1916 -1905 1926
rect -1713 1927 -1572 1978
rect -1520 1927 -1380 1979
rect -1328 1927 -1188 1979
rect -1136 1927 -997 1979
rect -945 1927 -720 1979
rect -1765 1916 -1713 1926
rect -1572 1917 -1520 1927
rect -1380 1917 -1328 1927
rect -1188 1917 -1136 1927
rect -997 1917 -945 1927
rect -720 1917 -668 1927
rect -434 1674 -370 2227
rect 3308 2223 3372 2233
rect 6764 2223 6828 2233
rect 3308 2149 3372 2159
rect 8595 1991 8659 2001
rect 7043 1979 7095 1988
rect 7235 1979 7287 1988
rect 7428 1979 7480 1989
rect 7620 1979 7672 1989
rect 7812 1979 7864 1989
rect 8003 1979 8055 1989
rect 8280 1979 8332 1989
rect 7036 1978 7428 1979
rect 7036 1927 7043 1978
rect 7095 1927 7235 1978
rect 7043 1916 7095 1926
rect 7287 1927 7428 1978
rect 7480 1927 7620 1979
rect 7672 1927 7812 1979
rect 7864 1927 8003 1979
rect 8055 1927 8280 1979
rect 8332 1927 8595 1979
rect 7235 1916 7287 1926
rect 7428 1917 7480 1927
rect 7620 1917 7672 1927
rect 7812 1917 7864 1927
rect 8003 1917 8055 1927
rect 8280 1917 8332 1927
rect 8595 1917 8659 1927
rect 4437 1704 4501 1714
rect 5426 1704 5490 1714
rect 540 1674 604 1684
rect 1830 1674 1894 1684
rect -434 1610 540 1674
rect 604 1610 1830 1674
rect 540 1600 604 1610
rect 1830 1600 1894 1610
rect 2330 1640 2394 1650
rect 4501 1640 5426 1704
rect 4437 1630 4501 1640
rect 5426 1630 5490 1640
rect 2330 1566 2394 1576
rect 3602 1526 3666 1536
rect 3602 1452 3666 1462
rect 3894 1522 3958 1532
rect 5736 1522 5800 1532
rect 3958 1458 5736 1522
rect 3894 1448 3958 1458
rect 5736 1448 5800 1458
rect 6152 1526 6216 1536
rect 6152 1452 6216 1462
rect 170 1341 234 1351
rect 170 1267 234 1277
rect 930 1341 994 1351
rect 3943 1341 4007 1351
rect 994 1277 3943 1341
rect 930 1267 994 1277
rect 3943 1267 4007 1277
rect 4326 1341 4390 1351
rect 4326 1267 4390 1277
rect -2651 998 -2587 1008
rect 8848 998 8912 1008
rect -1957 986 -1905 996
rect -1765 986 -1713 996
rect -1573 986 -1521 996
rect -1381 986 -1329 996
rect -1190 986 -1138 996
rect -997 986 -945 996
rect -720 986 -668 996
rect 7043 986 7095 996
rect 7235 986 7287 996
rect 7427 986 7479 996
rect 7619 986 7671 996
rect 7810 986 7862 996
rect 8003 986 8055 996
rect 8280 986 8332 996
rect -2587 934 -1957 986
rect -1905 934 -1765 986
rect -1713 934 -1573 986
rect -1521 934 -1381 986
rect -1329 934 -1190 986
rect -1138 934 -997 986
rect -945 934 -720 986
rect 7036 934 7043 986
rect 7095 934 7235 986
rect 7287 934 7427 986
rect 7479 934 7619 986
rect 7671 934 7810 986
rect 7862 934 8003 986
rect 8055 934 8280 986
rect 8332 934 8848 986
rect -2651 924 -2587 934
rect -1957 924 -1905 934
rect -1765 924 -1713 934
rect -1573 924 -1521 934
rect -1381 924 -1329 934
rect -1190 924 -1138 934
rect -997 924 -945 934
rect -720 924 -668 934
rect 7043 924 7095 934
rect 7235 924 7287 934
rect 7427 924 7479 934
rect 7619 924 7671 934
rect 7810 924 7862 934
rect 8003 924 8055 934
rect 8280 924 8332 934
rect 8848 924 8912 934
rect -1020 497 -956 507
rect -1020 348 -956 433
rect 6700 493 6764 503
rect 6700 419 6764 429
rect 1423 349 1487 359
rect -1020 285 1423 348
rect -1020 284 1487 285
rect 1423 275 1487 284
rect -2398 190 -2334 200
rect 8595 191 8659 201
rect -1957 179 -1905 188
rect -1765 179 -1713 188
rect -1572 179 -1520 189
rect -1380 179 -1328 189
rect -1188 179 -1136 189
rect -997 179 -945 189
rect -720 179 -668 189
rect 7043 179 7095 188
rect 7235 179 7287 188
rect 7428 179 7480 189
rect 7620 179 7672 189
rect 7812 179 7864 189
rect 8003 179 8055 189
rect 8280 179 8332 189
rect -1964 178 -1572 179
rect -2334 126 -1957 178
rect -1905 127 -1765 178
rect -2398 116 -2334 126
rect -1957 116 -1905 126
rect -1713 127 -1572 178
rect -1520 127 -1380 179
rect -1328 127 -1188 179
rect -1136 127 -997 179
rect -945 127 -720 179
rect 7036 178 7428 179
rect 7036 127 7043 178
rect -1765 116 -1713 126
rect -1572 117 -1520 127
rect -1380 117 -1328 127
rect -1188 117 -1136 127
rect -997 117 -945 127
rect -720 117 -668 127
rect 7095 127 7235 178
rect 7043 116 7095 126
rect 7287 127 7428 178
rect 7480 127 7620 179
rect 7672 127 7812 179
rect 7864 127 8003 179
rect 8055 127 8280 179
rect 8332 127 8595 179
rect 7235 116 7287 126
rect 7428 117 7480 127
rect 7620 117 7672 127
rect 7812 117 7864 127
rect 8003 117 8055 127
rect 8280 117 8332 127
rect 8595 117 8659 127
rect 160 -218 224 -208
rect -2651 -802 -2587 -792
rect -1957 -814 -1905 -804
rect -1765 -814 -1713 -804
rect -1573 -814 -1521 -804
rect -1381 -814 -1329 -804
rect -1190 -814 -1138 -804
rect -997 -814 -945 -804
rect -720 -814 -668 -804
rect -2587 -866 -1957 -814
rect -1905 -866 -1765 -814
rect -1713 -866 -1573 -814
rect -1521 -866 -1381 -814
rect -1329 -866 -1190 -814
rect -1138 -866 -997 -814
rect -945 -866 -720 -814
rect -2651 -876 -2587 -866
rect -1957 -876 -1905 -866
rect -1765 -876 -1713 -866
rect -1573 -876 -1521 -866
rect -1381 -876 -1329 -866
rect -1190 -876 -1138 -866
rect -997 -876 -945 -866
rect -720 -876 -668 -866
rect -364 -1074 -300 -1064
rect -1019 -1138 -364 -1074
rect -1019 -1304 -955 -1138
rect -364 -1148 -300 -1138
rect -1019 -1378 -955 -1368
rect -502 -1301 -438 -1291
rect 160 -1301 224 -282
rect 8848 -802 8912 -792
rect 7043 -814 7095 -804
rect 7235 -814 7287 -804
rect 7427 -814 7479 -804
rect 7619 -814 7671 -804
rect 7810 -814 7862 -804
rect 8003 -814 8055 -804
rect 8280 -814 8332 -804
rect 7036 -866 7043 -814
rect 7095 -866 7235 -814
rect 7287 -866 7427 -814
rect 7479 -866 7619 -814
rect 7671 -866 7810 -814
rect 7862 -866 8003 -814
rect 8055 -866 8280 -814
rect 8332 -866 8848 -814
rect 7043 -876 7095 -866
rect 7235 -876 7287 -866
rect 7427 -876 7479 -866
rect 7619 -876 7671 -866
rect 7810 -876 7862 -866
rect 8003 -876 8055 -866
rect 8280 -876 8332 -866
rect 8848 -876 8912 -866
rect -438 -1365 224 -1301
rect 6718 -1299 6782 -1289
rect -502 -1375 -438 -1365
rect 6718 -1373 6782 -1363
rect -2398 -1610 -2334 -1600
rect 8595 -1609 8659 -1599
rect -1957 -1621 -1905 -1612
rect -1765 -1621 -1713 -1612
rect -1572 -1621 -1520 -1611
rect -1380 -1621 -1328 -1611
rect -1188 -1621 -1136 -1611
rect -997 -1621 -945 -1611
rect -720 -1621 -668 -1611
rect 7043 -1621 7095 -1612
rect 7235 -1621 7287 -1612
rect 7428 -1621 7480 -1611
rect 7620 -1621 7672 -1611
rect 7812 -1621 7864 -1611
rect 8003 -1621 8055 -1611
rect 8280 -1621 8332 -1611
rect -1964 -1622 -1572 -1621
rect -2334 -1674 -1957 -1622
rect -1905 -1673 -1765 -1622
rect -2398 -1684 -2334 -1674
rect -1957 -1684 -1905 -1674
rect -1713 -1673 -1572 -1622
rect -1520 -1673 -1380 -1621
rect -1328 -1673 -1188 -1621
rect -1136 -1673 -997 -1621
rect -945 -1673 -720 -1621
rect 7036 -1622 7428 -1621
rect 7036 -1673 7043 -1622
rect -1765 -1684 -1713 -1674
rect -1572 -1683 -1520 -1673
rect -1380 -1683 -1328 -1673
rect -1188 -1683 -1136 -1673
rect -997 -1683 -945 -1673
rect -720 -1683 -668 -1673
rect 7095 -1673 7235 -1622
rect 7043 -1684 7095 -1674
rect 7287 -1673 7428 -1622
rect 7480 -1673 7620 -1621
rect 7672 -1673 7812 -1621
rect 7864 -1673 8003 -1621
rect 8055 -1673 8280 -1621
rect 8332 -1673 8595 -1621
rect 7235 -1684 7287 -1674
rect 7428 -1683 7480 -1673
rect 7620 -1683 7672 -1673
rect 7812 -1683 7864 -1673
rect 8003 -1683 8055 -1673
rect 8280 -1683 8332 -1673
rect 8595 -1683 8659 -1673
<< via2 >>
rect -2651 8134 -2587 8198
rect 8848 8134 8912 8198
rect -2398 7326 -2334 7390
rect 6691 7633 6755 7697
rect 8595 7327 8659 7391
rect 1996 6692 2060 6756
rect 1628 6412 1692 6476
rect -2651 6334 -2587 6398
rect 8848 6334 8912 6398
rect -477 5829 -413 5893
rect 6704 5831 6768 5895
rect -2398 5526 -2334 5590
rect 3410 5717 3474 5781
rect -197 5106 -133 5170
rect 1282 5548 1346 5612
rect -2651 4534 -2587 4598
rect 1630 5549 1694 5613
rect 1428 4155 1492 4219
rect -2398 3726 -2334 3790
rect 3157 5494 3221 5558
rect 8595 5527 8659 5591
rect 3410 5105 3474 5169
rect 3157 5020 3221 5084
rect 4658 5042 4722 5106
rect 5418 5042 5482 5106
rect 3768 4864 3832 4928
rect 4084 4864 4148 4928
rect 5706 4864 5770 4928
rect 6166 4868 6230 4932
rect 3106 4499 3170 4563
rect 8848 4534 8912 4598
rect 5207 4326 5271 4390
rect 3308 4148 3372 4212
rect 4876 3916 4940 3980
rect 5206 3916 5270 3980
rect 333 3419 397 3483
rect 765 3419 829 3483
rect 1408 3419 1472 3483
rect 1631 3419 1695 3483
rect 333 3263 397 3327
rect -2651 2734 -2587 2798
rect 333 3090 397 3154
rect 764 3089 828 3153
rect 3306 3798 3370 3862
rect 4874 3578 4938 3642
rect 8595 3727 8659 3791
rect 4510 3398 4574 3462
rect 4508 3087 4572 3151
rect 3306 2559 3370 2623
rect 8848 2734 8912 2798
rect -2398 1926 -2334 1990
rect 3308 2159 3372 2223
rect 8595 1927 8659 1991
rect 540 1610 604 1674
rect 1830 1610 1894 1674
rect 2330 1576 2394 1640
rect 4437 1640 4501 1704
rect 5426 1640 5490 1704
rect 3602 1462 3666 1526
rect 3894 1458 3958 1522
rect 5736 1458 5800 1522
rect 6152 1462 6216 1526
rect 170 1277 234 1341
rect 930 1277 994 1341
rect 3943 1277 4007 1341
rect 4326 1277 4390 1341
rect -2651 934 -2587 998
rect 8848 934 8912 998
rect 6700 429 6764 493
rect 1423 285 1487 349
rect -2398 126 -2334 190
rect 8595 127 8659 191
rect 160 -282 224 -218
rect -2651 -866 -2587 -802
rect -364 -1138 -300 -1074
rect 8848 -866 8912 -802
rect 6718 -1363 6782 -1299
rect -2398 -1674 -2334 -1610
rect 8595 -1673 8659 -1609
<< metal3 >>
rect -2651 8203 -2587 8208
rect -2661 8198 -2577 8203
rect -2661 8134 -2651 8198
rect -2587 8134 -2577 8198
rect -2661 8129 -2577 8134
rect -2651 6403 -2587 8129
rect -2398 7395 -2334 7400
rect -2408 7390 -2324 7395
rect -2408 7326 -2398 7390
rect -2334 7326 -2324 7390
rect -2408 7321 -2324 7326
rect -2661 6398 -2577 6403
rect -2661 6334 -2651 6398
rect -2587 6334 -2577 6398
rect -2661 6329 -2577 6334
rect -2651 4603 -2587 6329
rect -2398 5595 -2334 7321
rect -1800 7200 -641 8360
rect 0 7200 1159 8360
rect 1800 7200 2959 8360
rect 3600 7200 4759 8360
rect 5400 7200 6559 8360
rect 6681 7697 6765 7702
rect 6681 7633 6691 7697
rect 6755 7633 6765 7697
rect 6681 7628 6765 7633
rect 1975 6756 2080 6780
rect 6691 6779 6755 7628
rect 7200 7200 8359 8360
rect 8848 8203 8912 8208
rect 8838 8198 8922 8203
rect 8838 8134 8848 8198
rect 8912 8134 8922 8198
rect 8838 8129 8922 8134
rect 8595 7396 8659 7401
rect 8585 7391 8669 7396
rect 8585 7327 8595 7391
rect 8659 7327 8669 7391
rect 8585 7322 8669 7327
rect 1975 6692 1996 6756
rect 2060 6692 2080 6756
rect 1975 6669 2080 6692
rect 6191 6715 6755 6779
rect 6191 6560 6255 6715
rect -2408 5590 -2324 5595
rect -2408 5526 -2398 5590
rect -2334 5526 -2324 5590
rect -2408 5521 -2324 5526
rect -2661 4598 -2577 4603
rect -2661 4534 -2651 4598
rect -2587 4534 -2577 4598
rect -2661 4529 -2577 4534
rect -2651 4524 -2587 4529
rect -2398 3795 -2334 5521
rect -1800 5400 -641 6560
rect -497 5893 -391 5915
rect -497 5829 -477 5893
rect -413 5829 -391 5893
rect -497 5808 -391 5829
rect 0 5612 1159 6560
rect 1618 6476 1702 6481
rect 1800 6476 2959 6560
rect 1618 6412 1628 6476
rect 1692 6412 2959 6476
rect 1618 6407 1702 6412
rect 1272 5612 1356 5617
rect 0 5548 1282 5612
rect 1346 5548 1356 5612
rect 0 5400 1159 5548
rect 1272 5543 1356 5548
rect 1616 5613 1708 5646
rect 1616 5549 1630 5613
rect 1694 5549 1708 5613
rect 1616 5524 1708 5549
rect 1800 5400 2959 6412
rect 3600 6197 4759 6560
rect 3157 6133 4759 6197
rect 3157 5563 3221 6133
rect 3400 5781 3484 5810
rect 3400 5717 3410 5781
rect 3474 5717 3484 5781
rect 3400 5693 3484 5717
rect 3147 5558 3231 5563
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 3147 5489 3231 5494
rect 3600 5400 4759 6133
rect 5400 5400 6559 6560
rect 6686 5895 6784 5914
rect 6686 5831 6704 5895
rect 6768 5831 6784 5895
rect 6686 5814 6784 5831
rect 7200 5400 8359 6560
rect 8595 5596 8659 7322
rect 8848 6403 8912 8129
rect 8838 6398 8922 6403
rect 8838 6334 8848 6398
rect 8912 6334 8922 6398
rect 8838 6329 8922 6334
rect 8585 5591 8669 5596
rect 8585 5527 8595 5591
rect 8659 5527 8669 5591
rect 8585 5522 8669 5527
rect 544 5311 608 5400
rect 544 5247 5105 5311
rect -238 5170 -98 5201
rect -238 5106 -197 5170
rect -133 5106 -98 5170
rect -238 5072 -98 5106
rect 3379 5169 3508 5177
rect 3379 5105 3410 5169
rect 3474 5105 3508 5169
rect 3379 5097 3508 5105
rect 4648 5106 4732 5111
rect 3147 5084 3231 5089
rect 754 5020 3157 5084
rect 3221 5020 3231 5084
rect 4648 5042 4658 5106
rect 4722 5042 4732 5106
rect 4648 5037 4732 5042
rect 754 4760 818 5020
rect 3147 5015 3231 5020
rect 3758 4928 3842 4933
rect 1241 4864 3768 4928
rect 3832 4864 3842 4928
rect -2408 3790 -2324 3795
rect -2408 3726 -2398 3790
rect -2334 3726 -2324 3790
rect -2408 3721 -2324 3726
rect -1800 3600 -641 4760
rect 0 3600 1159 4760
rect 333 3488 397 3600
rect 323 3483 407 3488
rect 323 3419 333 3483
rect 397 3419 407 3483
rect 323 3414 407 3419
rect 743 3483 849 3501
rect 743 3419 765 3483
rect 829 3419 849 3483
rect 333 3332 397 3414
rect 743 3404 849 3419
rect 323 3327 407 3332
rect 323 3263 333 3327
rect 397 3263 407 3327
rect 323 3258 407 3263
rect 333 3159 397 3258
rect 323 3154 407 3159
rect 323 3090 333 3154
rect 397 3090 407 3154
rect 323 3085 407 3090
rect 745 3158 837 3183
rect 745 3153 838 3158
rect 745 3089 764 3153
rect 828 3089 838 3153
rect 333 2960 397 3085
rect 745 3084 838 3089
rect 745 3061 837 3084
rect -2651 2803 -2587 2808
rect -2661 2798 -2577 2803
rect -2661 2734 -2651 2798
rect -2587 2734 -2577 2798
rect -2661 2729 -2577 2734
rect -2651 1003 -2587 2729
rect -2398 1995 -2334 2000
rect -2408 1990 -2324 1995
rect -2408 1926 -2398 1990
rect -2334 1926 -2324 1990
rect -2408 1921 -2324 1926
rect -2661 998 -2577 1003
rect -2661 934 -2651 998
rect -2587 934 -2577 998
rect -2661 929 -2577 934
rect -2651 -797 -2587 929
rect -2398 195 -2334 1921
rect -1800 1800 -641 2960
rect 0 1800 1159 2960
rect 170 1346 234 1800
rect 530 1674 614 1679
rect 530 1610 540 1674
rect 604 1610 614 1674
rect 530 1605 614 1610
rect 160 1341 244 1346
rect 160 1277 170 1341
rect 234 1277 244 1341
rect 160 1272 244 1277
rect 540 1160 604 1605
rect 910 1341 1011 1357
rect 910 1277 930 1341
rect 994 1277 1011 1341
rect 910 1259 1011 1277
rect -2408 190 -2324 195
rect -2408 126 -2398 190
rect -2334 126 -2324 190
rect -2408 121 -2324 126
rect -2661 -802 -2577 -797
rect -2661 -866 -2651 -802
rect -2587 -866 -2577 -802
rect -2661 -871 -2577 -866
rect -2651 -876 -2587 -871
rect -2398 -1605 -2334 121
rect -1800 0 -641 1160
rect 0 354 1159 1160
rect 1241 354 1305 4864
rect 3758 4859 3842 4864
rect 4061 4928 4171 4944
rect 4061 4864 4084 4928
rect 4148 4864 4171 4928
rect 4061 4850 4171 4864
rect 4658 4760 4722 5037
rect 1418 4219 1502 4224
rect 1800 4219 2959 4760
rect 3081 4563 3190 4586
rect 3081 4499 3106 4563
rect 3170 4499 3190 4563
rect 3081 4479 3190 4499
rect 1418 4155 1428 4219
rect 1492 4155 2959 4219
rect 1418 4150 1502 4155
rect 1800 3600 2959 4155
rect 3298 4212 3382 4217
rect 3600 4212 4759 4760
rect 3298 4148 3308 4212
rect 3372 4148 4759 4212
rect 3298 4143 3382 4148
rect 3283 3862 3389 3885
rect 3283 3798 3306 3862
rect 3370 3798 3389 3862
rect 3283 3778 3389 3798
rect 3600 3600 4759 4148
rect 4862 3980 4953 4019
rect 4862 3916 4876 3980
rect 4940 3916 4953 3980
rect 4862 3879 4953 3916
rect 4864 3642 4948 3647
rect 1397 3483 1484 3517
rect 1397 3419 1408 3483
rect 1472 3419 1484 3483
rect 1397 3388 1484 3419
rect 1621 3483 1705 3488
rect 1621 3419 1631 3483
rect 1695 3419 1705 3483
rect 1621 3414 1705 3419
rect 2348 3432 2412 3600
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 4864 3573 4948 3578
rect 4479 3462 4604 3492
rect 0 290 1305 354
rect 1405 349 1503 380
rect 0 0 1159 290
rect 1405 285 1423 349
rect 1487 285 1503 349
rect 1631 365 1695 3414
rect 2348 3368 3912 3432
rect 4479 3398 4510 3462
rect 4574 3398 4604 3462
rect 4479 3371 4604 3398
rect 3848 2960 3912 3368
rect 4486 3151 4590 3171
rect 4486 3087 4508 3151
rect 4572 3087 4590 3151
rect 4486 3071 4590 3087
rect 1800 2223 2959 2960
rect 3284 2623 3390 2645
rect 3284 2559 3306 2623
rect 3370 2559 3390 2623
rect 3284 2538 3390 2559
rect 3298 2223 3382 2228
rect 1800 2159 3308 2223
rect 3372 2159 3382 2223
rect 1800 1800 2959 2159
rect 3298 2154 3382 2159
rect 3600 1800 4759 2960
rect 1830 1679 1894 1800
rect 4437 1709 4501 1800
rect 4427 1704 4511 1709
rect 1820 1674 1904 1679
rect 1820 1610 1830 1674
rect 1894 1610 1904 1674
rect 1820 1605 1904 1610
rect 2307 1640 2415 1666
rect 2307 1576 2330 1640
rect 2394 1576 2415 1640
rect 4427 1640 4437 1704
rect 4501 1640 4511 1704
rect 4427 1635 4511 1640
rect 2307 1553 2415 1576
rect 3592 1526 3676 1531
rect 3083 1462 3602 1526
rect 3666 1462 3676 1526
rect 1800 365 2959 1160
rect 1631 363 2959 365
rect 3083 363 3147 1462
rect 3592 1457 3676 1462
rect 3873 1522 3978 1546
rect 3873 1458 3894 1522
rect 3958 1458 3978 1522
rect 3873 1437 3978 1458
rect 3923 1341 4024 1360
rect 3923 1277 3943 1341
rect 4007 1277 4024 1341
rect 3923 1262 4024 1277
rect 4316 1341 4400 1346
rect 4316 1277 4326 1341
rect 4390 1277 4400 1341
rect 4316 1272 4400 1277
rect 4326 1160 4390 1272
rect 1631 301 3147 363
rect 1405 260 1503 285
rect 1800 299 3147 301
rect 3600 448 4759 1160
rect 4874 448 4938 3573
rect 5041 616 5105 5247
rect 5418 5111 5482 5400
rect 5408 5106 5492 5111
rect 5408 5042 5418 5106
rect 5482 5042 5492 5106
rect 5408 5037 5492 5042
rect 5683 4928 5793 4943
rect 6166 4937 6230 5400
rect 5683 4864 5706 4928
rect 5770 4864 5793 4928
rect 5683 4849 5793 4864
rect 6156 4932 6240 4937
rect 6156 4868 6166 4932
rect 6230 4868 6240 4932
rect 6156 4863 6240 4868
rect 5197 4390 5281 4395
rect 5400 4390 6559 4760
rect 5197 4326 5207 4390
rect 5271 4326 6559 4390
rect 5197 4321 5281 4326
rect 5193 3980 5284 4018
rect 5193 3916 5206 3980
rect 5270 3916 5284 3980
rect 5193 3878 5284 3916
rect 5400 3600 6559 4326
rect 7200 3600 8359 4760
rect 8595 3796 8659 5522
rect 8848 4603 8912 6329
rect 8838 4598 8922 4603
rect 8838 4534 8848 4598
rect 8912 4534 8922 4598
rect 8838 4529 8922 4534
rect 8585 3791 8669 3796
rect 8585 3727 8595 3791
rect 8659 3727 8669 3791
rect 8585 3722 8669 3727
rect 8595 3717 8659 3722
rect 5400 1800 6559 2960
rect 7200 1800 8359 2960
rect 8848 2803 8912 2808
rect 8838 2798 8922 2803
rect 8838 2734 8848 2798
rect 8912 2734 8922 2798
rect 8838 2729 8922 2734
rect 8595 1996 8659 2001
rect 8585 1991 8669 1996
rect 8585 1927 8595 1991
rect 8659 1927 8669 1991
rect 8585 1922 8669 1927
rect 5416 1704 5500 1709
rect 5416 1640 5426 1704
rect 5490 1640 5500 1704
rect 5416 1635 5500 1640
rect 5426 1160 5490 1635
rect 5715 1522 5820 1544
rect 6152 1531 6216 1800
rect 5715 1458 5736 1522
rect 5800 1458 5820 1522
rect 5715 1435 5820 1458
rect 6142 1526 6226 1531
rect 6142 1462 6152 1526
rect 6216 1462 6226 1526
rect 6142 1457 6226 1462
rect 5400 616 6559 1160
rect 5041 552 6559 616
rect 3600 384 4941 448
rect 1800 0 2959 299
rect 3600 0 4759 384
rect 5400 0 6559 552
rect 6683 493 6785 514
rect 6683 429 6700 493
rect 6764 429 6785 493
rect 6683 411 6785 429
rect 7200 0 8359 1160
rect 8595 196 8659 1922
rect 8848 1003 8912 2729
rect 8838 998 8922 1003
rect 8838 934 8848 998
rect 8912 934 8922 998
rect 8838 929 8922 934
rect 8585 191 8669 196
rect 8585 127 8595 191
rect 8659 127 8669 191
rect 8585 122 8669 127
rect 139 -218 245 -195
rect 139 -282 160 -218
rect 224 -282 245 -218
rect 139 -299 245 -282
rect 6179 -442 6243 0
rect 6179 -506 6782 -442
rect -2408 -1610 -2324 -1605
rect -2408 -1674 -2398 -1610
rect -2334 -1674 -2324 -1610
rect -2408 -1679 -2324 -1674
rect -2398 -1684 -2334 -1679
rect -1800 -1800 -641 -640
rect -378 -1074 -280 -1056
rect -378 -1138 -364 -1074
rect -300 -1138 -280 -1074
rect -378 -1159 -280 -1138
rect 0 -1800 1159 -640
rect 1800 -1800 2959 -640
rect 3600 -1800 4759 -640
rect 5400 -1800 6559 -640
rect 6718 -1294 6782 -506
rect 6708 -1299 6792 -1294
rect 6708 -1363 6718 -1299
rect 6782 -1363 6792 -1299
rect 6708 -1368 6792 -1363
rect 6718 -1372 6782 -1368
rect 7200 -1800 8359 -640
rect 8595 -1604 8659 122
rect 8848 -797 8912 929
rect 8838 -802 8922 -797
rect 8838 -866 8848 -802
rect 8912 -866 8922 -802
rect 8838 -871 8922 -866
rect 8585 -1609 8669 -1604
rect 8585 -1673 8595 -1609
rect 8659 -1673 8669 -1609
rect 8585 -1678 8669 -1673
rect 8595 -1683 8659 -1678
<< via3 >>
rect 1996 6692 2060 6756
rect -477 5829 -413 5893
rect 1630 5549 1694 5613
rect 3410 5717 3474 5781
rect 6704 5831 6768 5895
rect -197 5106 -133 5170
rect 3410 5105 3474 5169
rect 765 3419 829 3483
rect 764 3089 828 3153
rect 930 1277 994 1341
rect 4084 4864 4148 4928
rect 3106 4499 3170 4563
rect 3306 3798 3370 3862
rect 4876 3916 4940 3980
rect 1408 3419 1472 3483
rect 1423 285 1487 349
rect 4510 3398 4574 3462
rect 4508 3087 4572 3151
rect 3306 2559 3370 2623
rect 2330 1576 2394 1640
rect 3894 1458 3958 1522
rect 3943 1277 4007 1341
rect 5706 4864 5770 4928
rect 5206 3916 5270 3980
rect 5736 1458 5800 1522
rect 6700 429 6764 493
rect 160 -282 224 -218
rect -364 -1138 -300 -1074
<< mimcap >>
rect -1700 8220 -740 8260
rect -1700 7340 -1660 8220
rect -780 7340 -740 8220
rect -1700 7300 -740 7340
rect 100 8220 1060 8260
rect 100 7340 140 8220
rect 1020 7340 1060 8220
rect 100 7300 1060 7340
rect 1900 8220 2860 8260
rect 1900 7340 1940 8220
rect 2820 7340 2860 8220
rect 1900 7300 2860 7340
rect 3700 8220 4660 8260
rect 3700 7340 3740 8220
rect 4620 7340 4660 8220
rect 3700 7300 4660 7340
rect 5500 8220 6460 8260
rect 5500 7340 5540 8220
rect 6420 7340 6460 8220
rect 5500 7300 6460 7340
rect 7300 8220 8260 8260
rect 7300 7340 7340 8220
rect 8220 7340 8260 8220
rect 7300 7300 8260 7340
rect -1700 6420 -740 6460
rect -1700 5540 -1660 6420
rect -780 5540 -740 6420
rect -1700 5500 -740 5540
rect 100 6420 1060 6460
rect 100 5540 140 6420
rect 1020 5540 1060 6420
rect 100 5500 1060 5540
rect 1900 6420 2860 6460
rect 1900 5540 1940 6420
rect 2820 5540 2860 6420
rect 1900 5500 2860 5540
rect 3700 6420 4660 6460
rect 3700 5540 3740 6420
rect 4620 5540 4660 6420
rect 3700 5500 4660 5540
rect 5500 6420 6460 6460
rect 5500 5540 5540 6420
rect 6420 5540 6460 6420
rect 5500 5500 6460 5540
rect 7300 6420 8260 6460
rect 7300 5540 7340 6420
rect 8220 5540 8260 6420
rect 7300 5500 8260 5540
rect -1700 4620 -740 4660
rect -1700 3740 -1660 4620
rect -780 3740 -740 4620
rect -1700 3700 -740 3740
rect 100 4620 1060 4660
rect 100 3740 140 4620
rect 1020 3740 1060 4620
rect 100 3700 1060 3740
rect 1900 4620 2860 4660
rect 1900 3740 1940 4620
rect 2820 3740 2860 4620
rect 1900 3700 2860 3740
rect 3700 4620 4660 4660
rect 3700 3740 3740 4620
rect 4620 3740 4660 4620
rect 3700 3700 4660 3740
rect 5500 4620 6460 4660
rect 5500 3740 5540 4620
rect 6420 3740 6460 4620
rect 5500 3700 6460 3740
rect 7300 4620 8260 4660
rect 7300 3740 7340 4620
rect 8220 3740 8260 4620
rect 7300 3700 8260 3740
rect -1700 2820 -740 2860
rect -1700 1940 -1660 2820
rect -780 1940 -740 2820
rect -1700 1900 -740 1940
rect 100 2820 1060 2860
rect 100 1940 140 2820
rect 1020 1940 1060 2820
rect 100 1900 1060 1940
rect 1900 2820 2860 2860
rect 1900 1940 1940 2820
rect 2820 1940 2860 2820
rect 1900 1900 2860 1940
rect 3700 2820 4660 2860
rect 3700 1940 3740 2820
rect 4620 1940 4660 2820
rect 3700 1900 4660 1940
rect 5500 2820 6460 2860
rect 5500 1940 5540 2820
rect 6420 1940 6460 2820
rect 5500 1900 6460 1940
rect 7300 2820 8260 2860
rect 7300 1940 7340 2820
rect 8220 1940 8260 2820
rect 7300 1900 8260 1940
rect -1700 1020 -740 1060
rect -1700 140 -1660 1020
rect -780 140 -740 1020
rect -1700 100 -740 140
rect 100 1020 1060 1060
rect 100 140 140 1020
rect 1020 140 1060 1020
rect 100 100 1060 140
rect 1900 1020 2860 1060
rect 1900 140 1940 1020
rect 2820 140 2860 1020
rect 1900 100 2860 140
rect 3700 1020 4660 1060
rect 3700 140 3740 1020
rect 4620 140 4660 1020
rect 3700 100 4660 140
rect 5500 1020 6460 1060
rect 5500 140 5540 1020
rect 6420 140 6460 1020
rect 5500 100 6460 140
rect 7300 1020 8260 1060
rect 7300 140 7340 1020
rect 8220 140 8260 1020
rect 7300 100 8260 140
rect -1700 -780 -740 -740
rect -1700 -1660 -1660 -780
rect -780 -1660 -740 -780
rect -1700 -1700 -740 -1660
rect 100 -780 1060 -740
rect 100 -1660 140 -780
rect 1020 -1660 1060 -780
rect 100 -1700 1060 -1660
rect 1900 -780 2860 -740
rect 1900 -1660 1940 -780
rect 2820 -1660 2860 -780
rect 1900 -1700 2860 -1660
rect 3700 -780 4660 -740
rect 3700 -1660 3740 -780
rect 4620 -1660 4660 -780
rect 3700 -1700 4660 -1660
rect 5500 -780 6460 -740
rect 5500 -1660 5540 -780
rect 6420 -1660 6460 -780
rect 5500 -1700 6460 -1660
rect 7300 -780 8260 -740
rect 7300 -1660 7340 -780
rect 8220 -1660 8260 -780
rect 7300 -1700 8260 -1660
<< mimcapcontact >>
rect -1660 7340 -780 8220
rect 140 7340 1020 8220
rect 1940 7340 2820 8220
rect 3740 7340 4620 8220
rect 5540 7340 6420 8220
rect 7340 7340 8220 8220
rect -1660 5540 -780 6420
rect 140 5540 1020 6420
rect 1940 5540 2820 6420
rect 3740 5540 4620 6420
rect 5540 5540 6420 6420
rect 7340 5540 8220 6420
rect -1660 3740 -780 4620
rect 140 3740 1020 4620
rect 1940 3740 2820 4620
rect 3740 3740 4620 4620
rect 5540 3740 6420 4620
rect 7340 3740 8220 4620
rect -1660 1940 -780 2820
rect 140 1940 1020 2820
rect 1940 1940 2820 2820
rect 3740 1940 4620 2820
rect 5540 1940 6420 2820
rect 7340 1940 8220 2820
rect -1660 140 -780 1020
rect 140 140 1020 1020
rect 1940 140 2820 1020
rect 3740 140 4620 1020
rect 5540 140 6420 1020
rect 7340 140 8220 1020
rect -1660 -1660 -780 -780
rect 140 -1660 1020 -780
rect 1940 -1660 2820 -780
rect 3740 -1660 4620 -780
rect 5540 -1660 6420 -780
rect 7340 -1660 8220 -780
<< metal4 >>
rect -1661 8220 -779 8221
rect -1661 7340 -1660 8220
rect -780 7340 -779 8220
rect -1661 7339 -779 7340
rect 139 8220 1021 8221
rect 139 7340 140 8220
rect 1020 7340 1021 8220
rect 139 7339 1021 7340
rect 1939 8220 2821 8221
rect 1939 7340 1940 8220
rect 2820 7340 2821 8220
rect 1939 7339 2821 7340
rect 3739 8220 4621 8221
rect 3739 7340 3740 8220
rect 4620 7340 4621 8220
rect 3739 7339 4621 7340
rect 5539 8220 6421 8221
rect 5539 7340 5540 8220
rect 6420 7340 6421 8220
rect 5539 7339 6421 7340
rect 7339 8220 8221 8221
rect 7339 7340 7340 8220
rect 8220 7340 8221 8220
rect 7339 7339 8221 7340
rect 1995 6756 2061 6757
rect 1995 6692 1996 6756
rect 2060 6692 2061 6756
rect 1995 6691 2061 6692
rect 1996 6421 2060 6691
rect -1661 6420 -779 6421
rect -1661 5540 -1660 6420
rect -780 5540 -779 6420
rect 139 6420 1021 6421
rect -478 5893 -412 5894
rect 139 5893 140 6420
rect -478 5829 -477 5893
rect -413 5829 140 5893
rect -478 5828 -412 5829
rect -1661 5539 -779 5540
rect 139 5540 140 5829
rect 1020 5540 1021 6420
rect 1939 6420 2821 6421
rect 1629 5613 1695 5614
rect 1939 5613 1940 6420
rect 1629 5549 1630 5613
rect 1694 5549 1940 5613
rect 1629 5548 1695 5549
rect 139 5539 1021 5540
rect 1939 5540 1940 5549
rect 2820 5540 2821 6420
rect 3739 6420 4621 6421
rect 3409 5781 3475 5782
rect 3739 5781 3740 6420
rect 3409 5717 3410 5781
rect 3474 5717 3740 5781
rect 3409 5716 3475 5717
rect 1939 5539 2821 5540
rect 3739 5540 3740 5717
rect 4620 5540 4621 6420
rect 3739 5539 4621 5540
rect 5539 6420 6421 6421
rect 5539 5540 5540 6420
rect 6420 5895 6421 6420
rect 7339 6420 8221 6421
rect 6703 5895 6769 5896
rect 6420 5831 6704 5895
rect 6768 5831 6769 5895
rect 6420 5540 6421 5831
rect 6703 5830 6769 5831
rect 5539 5539 6421 5540
rect 7339 5540 7340 6420
rect 8220 5540 8221 6420
rect 7339 5539 8221 5540
rect 544 5311 608 5539
rect 544 5247 5105 5311
rect -198 5170 -132 5171
rect -198 5106 -197 5170
rect -133 5169 -132 5170
rect 3409 5169 3475 5170
rect -133 5106 3410 5169
rect -198 5105 3410 5106
rect 3474 5105 3475 5169
rect 320 4621 384 5105
rect 3409 5104 3475 5105
rect 4083 4928 4149 4929
rect 1242 4864 4084 4928
rect 4148 4864 4150 4928
rect -1661 4620 -779 4621
rect -1661 3740 -1660 4620
rect -780 3740 -779 4620
rect -1661 3739 -779 3740
rect 139 4620 1021 4621
rect 139 3740 140 4620
rect 1020 3740 1021 4620
rect 139 3739 1021 3740
rect 765 3484 829 3739
rect 764 3483 830 3484
rect 764 3419 765 3483
rect 829 3419 830 3483
rect 764 3418 830 3419
rect 763 3153 829 3154
rect 763 3089 764 3153
rect 828 3089 829 3153
rect 763 3088 829 3089
rect 764 2821 828 3088
rect -1661 2820 -779 2821
rect -1661 1940 -1660 2820
rect -780 1940 -779 2820
rect 139 2820 1021 2821
rect 139 2049 140 2820
rect -1661 1939 -779 1940
rect -364 1985 140 2049
rect -1661 1020 -779 1021
rect -1661 140 -1660 1020
rect -780 140 -779 1020
rect -1661 139 -779 140
rect -1661 -780 -779 -779
rect -1661 -1660 -1660 -780
rect -780 -1660 -779 -780
rect -364 -1073 -300 1985
rect 139 1940 140 1985
rect 1020 1940 1021 2820
rect 139 1939 1021 1940
rect 930 1342 994 1939
rect 929 1341 995 1342
rect 929 1277 930 1341
rect 994 1277 995 1341
rect 929 1276 995 1277
rect 139 1020 1021 1021
rect 139 140 140 1020
rect 1020 859 1021 1020
rect 1242 859 1306 4864
rect 4083 4863 4149 4864
rect 1939 4620 2821 4621
rect 1939 3740 1940 4620
rect 2820 4563 2821 4620
rect 3739 4620 4621 4621
rect 3105 4563 3171 4564
rect 2820 4499 3106 4563
rect 3170 4499 3171 4563
rect 2820 3740 2821 4499
rect 3105 4498 3171 4499
rect 3305 3862 3371 3863
rect 3739 3862 3740 4620
rect 3305 3798 3306 3862
rect 3370 3798 3740 3862
rect 3305 3797 3371 3798
rect 1939 3739 2821 3740
rect 3739 3740 3740 3798
rect 4620 3740 4621 4620
rect 4875 3980 4941 3981
rect 4875 3916 4876 3980
rect 4940 3916 4941 3980
rect 4875 3915 4941 3916
rect 3739 3739 4621 3740
rect 1407 3483 1473 3484
rect 1407 3419 1408 3483
rect 1472 3419 1473 3483
rect 1407 3418 1473 3419
rect 2348 3432 2412 3739
rect 4510 3463 4574 3739
rect 4509 3462 4575 3463
rect 1020 795 1306 859
rect 1408 813 1472 3418
rect 2348 3368 3912 3432
rect 4509 3398 4510 3462
rect 4574 3398 4575 3462
rect 4509 3397 4575 3398
rect 3848 2821 3912 3368
rect 4507 3151 4573 3152
rect 4507 3087 4508 3151
rect 4572 3087 4573 3151
rect 4507 3086 4573 3087
rect 4508 2821 4572 3086
rect 1939 2820 2821 2821
rect 1939 1940 1940 2820
rect 2820 2623 2821 2820
rect 3739 2820 4621 2821
rect 3305 2623 3371 2624
rect 2820 2559 3306 2623
rect 3370 2559 3371 2623
rect 2820 1940 2821 2559
rect 3305 2558 3371 2559
rect 1939 1939 2821 1940
rect 3739 1940 3740 2820
rect 4620 1940 4621 2820
rect 3739 1939 4621 1940
rect 2330 1641 2394 1939
rect 2329 1640 2395 1641
rect 2329 1576 2330 1640
rect 2394 1576 2395 1640
rect 2329 1575 2395 1576
rect 3893 1522 3959 1523
rect 3083 1458 3894 1522
rect 3958 1458 3959 1522
rect 1939 1020 2821 1021
rect 1939 813 1940 1020
rect 1020 140 1021 795
rect 1408 749 1940 813
rect 1422 349 1488 350
rect 1939 349 1940 749
rect 1420 285 1423 349
rect 1487 285 1940 349
rect 1422 284 1488 285
rect 139 139 1021 140
rect 1939 140 1940 285
rect 2820 812 2821 1020
rect 3083 812 3147 1458
rect 3893 1457 3959 1458
rect 3943 1342 4007 1345
rect 3942 1341 4008 1342
rect 3942 1277 3943 1341
rect 4007 1277 4008 1341
rect 3942 1276 4008 1277
rect 3943 1021 4007 1276
rect 2820 748 3147 812
rect 3739 1020 4621 1021
rect 2820 140 2821 748
rect 1939 139 2821 140
rect 3739 140 3740 1020
rect 4620 844 4621 1020
rect 4876 844 4940 3915
rect 4620 780 4940 844
rect 4620 140 4621 780
rect 5041 616 5105 5247
rect 5706 4929 5770 5539
rect 5705 4928 5771 4929
rect 5705 4864 5706 4928
rect 5770 4864 5771 4928
rect 5705 4863 5771 4864
rect 5539 4620 6421 4621
rect 5205 3980 5271 3981
rect 5539 3980 5540 4620
rect 5205 3916 5206 3980
rect 5270 3916 5540 3980
rect 5205 3915 5271 3916
rect 5539 3740 5540 3916
rect 6420 3740 6421 4620
rect 5539 3739 6421 3740
rect 7339 4620 8221 4621
rect 7339 3740 7340 4620
rect 8220 3740 8221 4620
rect 7339 3739 8221 3740
rect 5539 2820 6421 2821
rect 5539 1940 5540 2820
rect 6420 1940 6421 2820
rect 5539 1939 6421 1940
rect 7339 2820 8221 2821
rect 7339 1940 7340 2820
rect 8220 1940 8221 2820
rect 7339 1939 8221 1940
rect 5736 1523 5800 1939
rect 5735 1522 5801 1523
rect 5735 1458 5736 1522
rect 5800 1458 5801 1522
rect 5735 1457 5801 1458
rect 5539 1020 6421 1021
rect 5539 616 5540 1020
rect 5041 552 5540 616
rect 3739 139 4621 140
rect 5539 140 5540 552
rect 6420 493 6421 1020
rect 7339 1020 8221 1021
rect 6699 493 6765 494
rect 6420 429 6700 493
rect 6764 429 6766 493
rect 6420 140 6421 429
rect 6699 428 6765 429
rect 5539 139 6421 140
rect 7339 140 7340 1020
rect 8220 140 8221 1020
rect 7339 139 8221 140
rect 160 -217 224 139
rect 159 -218 225 -217
rect 159 -282 160 -218
rect 224 -282 225 -218
rect 159 -283 225 -282
rect 139 -780 1021 -779
rect -365 -1074 -299 -1073
rect -365 -1138 -364 -1074
rect -300 -1138 -299 -1074
rect -365 -1139 -299 -1138
rect -1661 -1661 -779 -1660
rect 139 -1660 140 -780
rect 1020 -1660 1021 -780
rect 139 -1661 1021 -1660
rect 1939 -780 2821 -779
rect 1939 -1660 1940 -780
rect 2820 -1660 2821 -780
rect 1939 -1661 2821 -1660
rect 3739 -780 4621 -779
rect 3739 -1660 3740 -780
rect 4620 -1660 4621 -780
rect 3739 -1661 4621 -1660
rect 5539 -780 6421 -779
rect 5539 -1660 5540 -780
rect 6420 -1660 6421 -780
rect 5539 -1661 6421 -1660
rect 7339 -780 8221 -779
rect 7339 -1660 7340 -780
rect 8220 -1660 8221 -780
rect 7339 -1661 8221 -1660
<< labels >>
flabel metal3 -2642 8019 -2642 8019 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal3 -2389 7236 -2389 7236 1 FreeSans 400 0 0 0 p2
port 7 n
flabel metal3 -2639 2626 -2639 2626 1 FreeSans 400 0 0 0 p1_b
port 8 n
flabel metal3 -2389 1840 -2389 1840 1 FreeSans 400 0 0 0 p1
port 9 n
flabel metal3 8645 -1537 8645 -1537 1 FreeSans 400 0 0 0 p1
port 9 n
flabel metal3 8898 -670 8898 -670 1 FreeSans 400 0 0 0 p1_b
port 8 n
flabel metal3 8648 7246 8648 7246 1 FreeSans 400 0 0 0 p2
port 7 n
flabel metal3 8904 8016 8904 8016 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal1 -3484 3369 -3484 3369 1 FreeSans 400 0 0 0 op
port 4 n
flabel metal1 -2872 3368 -2872 3368 1 FreeSans 400 0 0 0 on
port 1 n
flabel metal1 -2412 3371 -2412 3371 1 FreeSans 400 0 0 0 cmc
port 5 n
flabel metal1 8790 3295 8790 3295 1 FreeSans 400 0 0 0 cm
port 2 n
flabel metal1 9292 3298 9292 3298 1 FreeSans 400 0 0 0 bias_a
port 3 n
flabel metal1 -2046 8350 -2046 8350 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 7178 -2045 7178 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2043 6543 -2043 6543 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 5370 -2045 5370 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2043 4743 -2043 4743 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2047 3574 -2047 3574 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2047 2942 -2047 2942 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 1776 -2045 1776 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2043 1146 -2043 1146 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2047 -27 -2047 -27 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 -2045 -659 -2045 -659 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 -1822 -2045 -1822 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6957 -1822 6957 -1822 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6954 -659 6954 -659 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6957 -26 6957 -26 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6952 1141 6952 1141 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6952 1776 6952 1776 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6954 2944 6954 2944 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6954 3579 6954 3579 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6957 4740 6957 4740 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6954 5375 6954 5375 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6952 6547 6952 6547 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 6954 7180 6954 7180 1 FreeSans 400 0 0 0 VSS
port 11 n power bidirectional
flabel metal1 6954 8345 6954 8345 1 FreeSans 400 0 0 0 VDD
port 10 n power bidirectional
flabel metal1 -2045 -1797 -2045 -1797 1 FreeSans 400 0 0 0 transmission_gate_11/VSS
flabel metal1 -2045 -691 -2045 -691 5 FreeSans 400 0 0 0 transmission_gate_11/VDD
flabel metal1 -646 -840 -646 -840 7 FreeSans 400 0 0 0 transmission_gate_11/en_b
flabel metal1 -645 -1336 -645 -1336 7 FreeSans 400 0 0 0 transmission_gate_11/in
flabel metal1 -645 -1647 -645 -1647 7 FreeSans 400 0 0 0 transmission_gate_11/en
flabel metal1 -2136 -1337 -2136 -1337 3 FreeSans 400 0 0 0 transmission_gate_11/out
flabel metal1 6955 -1797 6955 -1797 1 FreeSans 400 0 0 0 transmission_gate_2/VSS
flabel metal1 6955 -691 6955 -691 5 FreeSans 400 0 0 0 transmission_gate_2/VDD
flabel metal1 8354 -840 8354 -840 7 FreeSans 400 0 0 0 transmission_gate_2/en_b
flabel metal1 8355 -1336 8355 -1336 7 FreeSans 400 0 0 0 transmission_gate_2/in
flabel metal1 8355 -1647 8355 -1647 7 FreeSans 400 0 0 0 transmission_gate_2/en
flabel metal1 6864 -1337 6864 -1337 3 FreeSans 400 0 0 0 transmission_gate_2/out
flabel metal1 -2045 3 -2045 3 1 FreeSans 400 0 0 0 transmission_gate_10/VSS
flabel metal1 -2045 1109 -2045 1109 5 FreeSans 400 0 0 0 transmission_gate_10/VDD
flabel metal1 -646 960 -646 960 7 FreeSans 400 0 0 0 transmission_gate_10/en_b
flabel metal1 -645 464 -645 464 7 FreeSans 400 0 0 0 transmission_gate_10/in
flabel metal1 -645 153 -645 153 7 FreeSans 400 0 0 0 transmission_gate_10/en
flabel metal1 -2136 463 -2136 463 3 FreeSans 400 0 0 0 transmission_gate_10/out
flabel metal1 6955 3 6955 3 1 FreeSans 400 0 0 0 transmission_gate_0/VSS
flabel metal1 6955 1109 6955 1109 5 FreeSans 400 0 0 0 transmission_gate_0/VDD
flabel metal1 8354 960 8354 960 7 FreeSans 400 0 0 0 transmission_gate_0/en_b
flabel metal1 8355 464 8355 464 7 FreeSans 400 0 0 0 transmission_gate_0/in
flabel metal1 8355 153 8355 153 7 FreeSans 400 0 0 0 transmission_gate_0/en
flabel metal1 6864 463 6864 463 3 FreeSans 400 0 0 0 transmission_gate_0/out
flabel metal1 -2045 1803 -2045 1803 1 FreeSans 400 0 0 0 transmission_gate_9/VSS
flabel metal1 -2045 2909 -2045 2909 5 FreeSans 400 0 0 0 transmission_gate_9/VDD
flabel metal1 -646 2760 -646 2760 7 FreeSans 400 0 0 0 transmission_gate_9/en_b
flabel metal1 -645 2264 -645 2264 7 FreeSans 400 0 0 0 transmission_gate_9/in
flabel metal1 -645 1953 -645 1953 7 FreeSans 400 0 0 0 transmission_gate_9/en
flabel metal1 -2136 2263 -2136 2263 3 FreeSans 400 0 0 0 transmission_gate_9/out
flabel metal1 6955 1803 6955 1803 1 FreeSans 400 0 0 0 transmission_gate_1/VSS
flabel metal1 6955 2909 6955 2909 5 FreeSans 400 0 0 0 transmission_gate_1/VDD
flabel metal1 8354 2760 8354 2760 7 FreeSans 400 0 0 0 transmission_gate_1/en_b
flabel metal1 8355 2264 8355 2264 7 FreeSans 400 0 0 0 transmission_gate_1/in
flabel metal1 8355 1953 8355 1953 7 FreeSans 400 0 0 0 transmission_gate_1/en
flabel metal1 6864 2263 6864 2263 3 FreeSans 400 0 0 0 transmission_gate_1/out
flabel metal1 -2045 3603 -2045 3603 1 FreeSans 400 0 0 0 transmission_gate_8/VSS
flabel metal1 -2045 4709 -2045 4709 5 FreeSans 400 0 0 0 transmission_gate_8/VDD
flabel metal1 -646 4560 -646 4560 7 FreeSans 400 0 0 0 transmission_gate_8/en_b
flabel metal1 -645 4064 -645 4064 7 FreeSans 400 0 0 0 transmission_gate_8/in
flabel metal1 -645 3753 -645 3753 7 FreeSans 400 0 0 0 transmission_gate_8/en
flabel metal1 -2136 4063 -2136 4063 3 FreeSans 400 0 0 0 transmission_gate_8/out
flabel metal1 6955 3603 6955 3603 1 FreeSans 400 0 0 0 transmission_gate_3/VSS
flabel metal1 6955 4709 6955 4709 5 FreeSans 400 0 0 0 transmission_gate_3/VDD
flabel metal1 8354 4560 8354 4560 7 FreeSans 400 0 0 0 transmission_gate_3/en_b
flabel metal1 8355 4064 8355 4064 7 FreeSans 400 0 0 0 transmission_gate_3/in
flabel metal1 8355 3753 8355 3753 7 FreeSans 400 0 0 0 transmission_gate_3/en
flabel metal1 6864 4063 6864 4063 3 FreeSans 400 0 0 0 transmission_gate_3/out
flabel metal1 -2045 5403 -2045 5403 1 FreeSans 400 0 0 0 transmission_gate_7/VSS
flabel metal1 -2045 6509 -2045 6509 5 FreeSans 400 0 0 0 transmission_gate_7/VDD
flabel metal1 -646 6360 -646 6360 7 FreeSans 400 0 0 0 transmission_gate_7/en_b
flabel metal1 -645 5864 -645 5864 7 FreeSans 400 0 0 0 transmission_gate_7/in
flabel metal1 -645 5553 -645 5553 7 FreeSans 400 0 0 0 transmission_gate_7/en
flabel metal1 -2136 5863 -2136 5863 3 FreeSans 400 0 0 0 transmission_gate_7/out
flabel metal1 6955 5403 6955 5403 1 FreeSans 400 0 0 0 transmission_gate_4/VSS
flabel metal1 6955 6509 6955 6509 5 FreeSans 400 0 0 0 transmission_gate_4/VDD
flabel metal1 8354 6360 8354 6360 7 FreeSans 400 0 0 0 transmission_gate_4/en_b
flabel metal1 8355 5864 8355 5864 7 FreeSans 400 0 0 0 transmission_gate_4/in
flabel metal1 8355 5553 8355 5553 7 FreeSans 400 0 0 0 transmission_gate_4/en
flabel metal1 6864 5863 6864 5863 3 FreeSans 400 0 0 0 transmission_gate_4/out
flabel metal1 -2045 7203 -2045 7203 1 FreeSans 400 0 0 0 transmission_gate_6/VSS
flabel metal1 -2045 8309 -2045 8309 5 FreeSans 400 0 0 0 transmission_gate_6/VDD
flabel metal1 -646 8160 -646 8160 7 FreeSans 400 0 0 0 transmission_gate_6/en_b
flabel metal1 -645 7664 -645 7664 7 FreeSans 400 0 0 0 transmission_gate_6/in
flabel metal1 -645 7353 -645 7353 7 FreeSans 400 0 0 0 transmission_gate_6/en
flabel metal1 -2136 7663 -2136 7663 3 FreeSans 400 0 0 0 transmission_gate_6/out
flabel metal1 6955 7203 6955 7203 1 FreeSans 400 0 0 0 transmission_gate_5/VSS
flabel metal1 6955 8309 6955 8309 5 FreeSans 400 0 0 0 transmission_gate_5/VDD
flabel metal1 8354 8160 8354 8160 7 FreeSans 400 0 0 0 transmission_gate_5/en_b
flabel metal1 8355 7664 8355 7664 7 FreeSans 400 0 0 0 transmission_gate_5/in
flabel metal1 8355 7353 8355 7353 7 FreeSans 400 0 0 0 transmission_gate_5/en
flabel metal1 6864 7663 6864 7663 3 FreeSans 400 0 0 0 transmission_gate_5/out
<< end >>
