magic
tech sky130A
magscale 1 2
timestamp 1654674269
<< nwell >>
rect 5734 5006 13811 6712
rect 7933 3685 13811 5006
<< pwell >>
rect 13904 3655 21142 4529
rect 5450 -332 21142 3655
<< psubdiff >>
rect 14053 4265 14171 4314
rect 20754 4265 20865 4314
rect 14053 4229 14102 4265
rect 14053 3599 14102 3625
rect 7667 3550 7797 3599
rect 14025 3550 14102 3599
rect 20816 4213 20865 4265
rect 20816 -264 20865 -186
rect 7566 -313 7821 -264
rect 20722 -313 20865 -264
<< nsubdiff >>
rect 6594 6622 6727 6656
rect 13581 6622 13716 6656
rect 13682 6517 13716 6622
rect 6562 5044 6762 5078
rect 7918 5044 8027 5078
rect 7993 4980 8027 5044
rect 7993 3789 8027 3886
rect 13682 3789 13716 3863
rect 7993 3755 8102 3789
rect 13573 3755 13716 3789
<< psubdiffcont >>
rect 14171 4265 20754 4314
rect 14053 3625 14102 4229
rect 7797 3550 14025 3599
rect 20816 -186 20865 4213
rect 7821 -313 20722 -264
<< nsubdiffcont >>
rect 6727 6622 13581 6656
rect 6762 5044 7918 5078
rect 7993 3886 8027 4980
rect 13682 3863 13716 6517
rect 8102 3755 13573 3789
<< locali >>
rect 7687 6656 13766 6712
rect 6559 6622 6727 6656
rect 13581 6622 13766 6656
rect 7687 6584 13766 6622
rect 8152 5335 8280 6584
rect 10768 6444 10973 6584
rect 10768 6249 10974 6444
rect 6562 5044 6762 5078
rect 7918 5044 8027 5078
rect 7993 4980 8027 5044
rect 2569 3157 2666 4903
rect 7451 4656 7588 4906
rect 7993 3789 8027 3886
rect 8521 3789 8629 4905
rect 10768 3789 10973 6249
rect 13451 5318 13579 6584
rect 13682 6517 13716 6584
rect 13093 3789 13221 4874
rect 13682 3789 13716 3863
rect 7993 3755 8102 3789
rect 13573 3755 13716 3789
rect 14053 4265 14171 4314
rect 20754 4265 20865 4314
rect 14053 4229 14102 4265
rect 13093 3748 13221 3755
rect 14053 3599 14102 3625
rect 7667 3550 7797 3599
rect 14025 3550 14102 3599
rect 15453 3574 15590 4265
rect 8132 -186 8269 3550
rect 10765 -186 10959 3550
rect 13447 -186 13584 3550
rect 13842 -186 13979 3550
rect 17183 -186 17377 4265
rect 18961 3593 19098 4265
rect 20816 4213 20865 4265
rect 20576 -186 20713 3176
rect 7740 -264 20950 -186
rect 7740 -313 7821 -264
rect 20722 -313 20950 -264
rect 7740 -314 20950 -313
<< viali >>
rect 6727 6622 13581 6656
rect 8436 6228 8470 6262
rect 8792 6228 8826 6262
rect 9148 6228 9182 6262
rect 9504 6228 9538 6262
rect 9860 6228 9894 6262
rect 10216 6228 10250 6262
rect 10572 6228 10606 6262
rect 8614 6006 8648 6040
rect 8970 6006 9004 6040
rect 9326 6006 9360 6040
rect 9682 6006 9716 6040
rect 10038 6006 10072 6040
rect 10394 6006 10428 6040
rect 8436 5651 8470 5685
rect 8792 5651 8826 5685
rect 9148 5651 9182 5685
rect 9504 5651 9538 5685
rect 9860 5651 9894 5685
rect 10216 5651 10250 5685
rect 10572 5651 10606 5685
rect 8614 5429 8648 5463
rect 8970 5429 9004 5463
rect 9326 5429 9360 5463
rect 9682 5429 9716 5463
rect 10038 5429 10072 5463
rect 10394 5429 10428 5463
rect 8792 4770 8826 4804
rect 9148 4770 9182 4804
rect 9504 4770 9538 4804
rect 9860 4770 9894 4804
rect 10216 4770 10250 4804
rect 10572 4770 10606 4804
rect 8970 4548 9004 4582
rect 9326 4548 9360 4582
rect 9682 4548 9716 4582
rect 10038 4548 10072 4582
rect 10394 4548 10428 4582
rect 8792 4200 8826 4234
rect 9148 4200 9182 4234
rect 9504 4200 9538 4234
rect 9860 4200 9894 4234
rect 10216 4200 10250 4234
rect 10572 4200 10606 4234
rect 8970 3978 9004 4012
rect 9326 3978 9360 4012
rect 9682 3978 9716 4012
rect 10038 3978 10072 4012
rect 10394 3978 10428 4012
rect 11122 6228 11156 6262
rect 11478 6228 11512 6262
rect 11834 6228 11868 6262
rect 12190 6228 12224 6262
rect 12546 6228 12580 6262
rect 12902 6228 12936 6262
rect 13258 6228 13292 6262
rect 11300 6006 11334 6040
rect 11656 6006 11690 6040
rect 12012 6006 12046 6040
rect 12368 6006 12402 6040
rect 12724 6006 12758 6040
rect 13080 6006 13114 6040
rect 11122 5650 11156 5684
rect 11478 5650 11512 5684
rect 11834 5650 11868 5684
rect 12190 5650 12224 5684
rect 12546 5650 12580 5684
rect 12902 5650 12936 5684
rect 13258 5650 13292 5684
rect 11300 5428 11334 5462
rect 11656 5428 11690 5462
rect 12012 5428 12046 5462
rect 12368 5428 12402 5462
rect 12724 5428 12758 5462
rect 13080 5428 13114 5462
rect 11122 4770 11156 4804
rect 11478 4770 11512 4804
rect 11834 4770 11868 4804
rect 12190 4770 12224 4804
rect 12546 4770 12580 4804
rect 12902 4770 12936 4804
rect 11300 4548 11334 4582
rect 11656 4548 11690 4582
rect 12012 4548 12046 4582
rect 12368 4548 12402 4582
rect 12724 4548 12758 4582
rect 11122 4200 11156 4234
rect 11478 4200 11512 4234
rect 11834 4200 11868 4234
rect 12190 4200 12224 4234
rect 12546 4200 12580 4234
rect 12902 4200 12936 4234
rect 11300 3978 11334 4012
rect 11656 3978 11690 4012
rect 12012 3978 12046 4012
rect 12368 3978 12402 4012
rect 12724 3978 12758 4012
rect 15792 3850 15826 3884
rect 16004 3850 16038 3884
rect 16216 3850 16250 3884
rect 16428 3850 16462 3884
rect 16640 3850 16674 3884
rect 16852 3850 16886 3884
rect 15890 3668 15924 3702
rect 16102 3668 16136 3702
rect 16314 3668 16348 3702
rect 16526 3668 16560 3702
rect 16738 3668 16772 3702
rect 16950 3668 16984 3702
rect 8434 3270 8468 3304
rect 8790 3270 8824 3304
rect 9146 3270 9180 3304
rect 9502 3270 9536 3304
rect 9858 3270 9892 3304
rect 10214 3270 10248 3304
rect 10570 3270 10604 3304
rect 8612 3048 8646 3082
rect 8968 3048 9002 3082
rect 9324 3048 9358 3082
rect 9680 3048 9714 3082
rect 10036 3048 10070 3082
rect 10392 3048 10426 3082
rect 8434 2770 8468 2804
rect 8790 2770 8824 2804
rect 9146 2770 9180 2804
rect 9502 2770 9536 2804
rect 9858 2770 9892 2804
rect 10214 2770 10248 2804
rect 10570 2770 10604 2804
rect 8612 2548 8646 2582
rect 8968 2548 9002 2582
rect 9324 2548 9358 2582
rect 9680 2548 9714 2582
rect 10036 2548 10070 2582
rect 10392 2548 10426 2582
rect 8434 2270 8468 2304
rect 8790 2270 8824 2304
rect 9146 2270 9180 2304
rect 9502 2270 9536 2304
rect 9858 2270 9892 2304
rect 10214 2270 10248 2304
rect 10570 2270 10604 2304
rect 8612 2048 8646 2082
rect 8968 2048 9002 2082
rect 9324 2048 9358 2082
rect 9680 2048 9714 2082
rect 10036 2048 10070 2082
rect 10392 2048 10426 2082
rect 8434 1570 8468 1604
rect 8790 1570 8824 1604
rect 9146 1570 9180 1604
rect 9502 1570 9536 1604
rect 9858 1570 9892 1604
rect 10214 1570 10248 1604
rect 10570 1570 10604 1604
rect 8612 1348 8646 1382
rect 8968 1348 9002 1382
rect 9324 1348 9358 1382
rect 9680 1348 9714 1382
rect 10036 1348 10070 1382
rect 10392 1348 10426 1382
rect 8434 1070 8468 1104
rect 8790 1070 8824 1104
rect 9146 1070 9180 1104
rect 9502 1070 9536 1104
rect 9858 1070 9892 1104
rect 10214 1070 10248 1104
rect 10570 1070 10604 1104
rect 8612 848 8646 882
rect 8968 848 9002 882
rect 9324 848 9358 882
rect 9680 848 9714 882
rect 10036 848 10070 882
rect 10392 848 10426 882
rect 8434 570 8468 604
rect 8790 570 8824 604
rect 9146 570 9180 604
rect 9502 570 9536 604
rect 9858 570 9892 604
rect 10214 570 10248 604
rect 10570 570 10604 604
rect 8612 348 8646 382
rect 8968 348 9002 382
rect 9324 348 9358 382
rect 9680 348 9714 382
rect 10036 348 10070 382
rect 10392 348 10426 382
rect 11121 3270 11155 3304
rect 11477 3270 11511 3304
rect 11833 3270 11867 3304
rect 12189 3270 12223 3304
rect 12545 3270 12579 3304
rect 12901 3270 12935 3304
rect 13257 3270 13291 3304
rect 11299 3048 11333 3082
rect 11655 3048 11689 3082
rect 12011 3048 12045 3082
rect 12367 3048 12401 3082
rect 12723 3048 12757 3082
rect 13079 3048 13113 3082
rect 11121 2770 11155 2804
rect 11477 2770 11511 2804
rect 11833 2770 11867 2804
rect 12189 2770 12223 2804
rect 12545 2770 12579 2804
rect 12901 2770 12935 2804
rect 13257 2770 13291 2804
rect 11299 2548 11333 2582
rect 11655 2548 11689 2582
rect 12011 2548 12045 2582
rect 12367 2548 12401 2582
rect 12723 2548 12757 2582
rect 13079 2548 13113 2582
rect 11121 2270 11155 2304
rect 11477 2270 11511 2304
rect 11833 2270 11867 2304
rect 12189 2270 12223 2304
rect 12545 2270 12579 2304
rect 12901 2270 12935 2304
rect 13257 2270 13291 2304
rect 11299 2048 11333 2082
rect 11655 2048 11689 2082
rect 12011 2048 12045 2082
rect 12367 2048 12401 2082
rect 12723 2048 12757 2082
rect 13079 2048 13113 2082
rect 11121 1570 11155 1604
rect 11477 1570 11511 1604
rect 11833 1570 11867 1604
rect 12189 1570 12223 1604
rect 12545 1570 12579 1604
rect 12901 1570 12935 1604
rect 13257 1570 13291 1604
rect 11299 1348 11333 1382
rect 11655 1348 11689 1382
rect 12011 1348 12045 1382
rect 12367 1348 12401 1382
rect 12723 1348 12757 1382
rect 13079 1348 13113 1382
rect 11121 1070 11155 1104
rect 11477 1070 11511 1104
rect 11833 1070 11867 1104
rect 12189 1070 12223 1104
rect 12545 1070 12579 1104
rect 12901 1070 12935 1104
rect 13257 1070 13291 1104
rect 11299 848 11333 882
rect 11655 848 11689 882
rect 12011 848 12045 882
rect 12367 848 12401 882
rect 12723 848 12757 882
rect 13079 848 13113 882
rect 11121 570 11155 604
rect 11477 570 11511 604
rect 11833 570 11867 604
rect 12189 570 12223 604
rect 12545 570 12579 604
rect 12901 570 12935 604
rect 13257 570 13291 604
rect 11299 348 11333 382
rect 11655 348 11689 382
rect 12011 348 12045 382
rect 12367 348 12401 382
rect 12723 348 12757 382
rect 13079 348 13113 382
rect 14138 3070 14172 3104
rect 14494 3070 14528 3104
rect 14850 3070 14884 3104
rect 15206 3070 15240 3104
rect 15562 3070 15596 3104
rect 15918 3070 15952 3104
rect 16274 3070 16308 3104
rect 16630 3070 16664 3104
rect 16986 3070 17020 3104
rect 14316 2848 14350 2882
rect 14672 2848 14706 2882
rect 15028 2848 15062 2882
rect 15384 2848 15418 2882
rect 15740 2848 15774 2882
rect 16096 2848 16130 2882
rect 16452 2848 16486 2882
rect 16808 2848 16842 2882
rect 14138 2570 14172 2604
rect 14494 2570 14528 2604
rect 14850 2570 14884 2604
rect 15206 2570 15240 2604
rect 15562 2570 15596 2604
rect 15918 2570 15952 2604
rect 16274 2570 16308 2604
rect 16630 2570 16664 2604
rect 16986 2570 17020 2604
rect 14316 2348 14350 2382
rect 14672 2348 14706 2382
rect 15028 2348 15062 2382
rect 15384 2348 15418 2382
rect 15740 2348 15774 2382
rect 16096 2348 16130 2382
rect 16452 2348 16486 2382
rect 16808 2348 16842 2382
rect 14138 2070 14172 2104
rect 14494 2070 14528 2104
rect 14850 2070 14884 2104
rect 15206 2070 15240 2104
rect 15562 2070 15596 2104
rect 15918 2070 15952 2104
rect 16274 2070 16308 2104
rect 16630 2070 16664 2104
rect 16986 2070 17020 2104
rect 14316 1848 14350 1882
rect 14672 1848 14706 1882
rect 15028 1848 15062 1882
rect 15384 1848 15418 1882
rect 15740 1848 15774 1882
rect 16096 1848 16130 1882
rect 16452 1848 16486 1882
rect 16808 1848 16842 1882
rect 14138 1570 14172 1604
rect 14494 1570 14528 1604
rect 14850 1570 14884 1604
rect 15206 1570 15240 1604
rect 15562 1570 15596 1604
rect 15918 1570 15952 1604
rect 16274 1570 16308 1604
rect 16630 1570 16664 1604
rect 16986 1570 17020 1604
rect 14316 1348 14350 1382
rect 14672 1348 14706 1382
rect 15028 1348 15062 1382
rect 15384 1348 15418 1382
rect 15740 1348 15774 1382
rect 16096 1348 16130 1382
rect 16452 1348 16486 1382
rect 16808 1348 16842 1382
rect 14138 1070 14172 1104
rect 14494 1070 14528 1104
rect 14850 1070 14884 1104
rect 15206 1070 15240 1104
rect 15562 1070 15596 1104
rect 15918 1070 15952 1104
rect 16274 1070 16308 1104
rect 16630 1070 16664 1104
rect 16986 1070 17020 1104
rect 14316 848 14350 882
rect 14672 848 14706 882
rect 15028 848 15062 882
rect 15384 848 15418 882
rect 15740 848 15774 882
rect 16096 848 16130 882
rect 16452 848 16486 882
rect 16808 848 16842 882
rect 14138 570 14172 604
rect 14494 570 14528 604
rect 14850 570 14884 604
rect 15206 570 15240 604
rect 15562 570 15596 604
rect 15918 570 15952 604
rect 16274 570 16308 604
rect 16630 570 16664 604
rect 16986 570 17020 604
rect 14316 348 14350 382
rect 14672 348 14706 382
rect 15028 348 15062 382
rect 15384 348 15418 382
rect 15740 348 15774 382
rect 16096 348 16130 382
rect 16452 348 16486 382
rect 16808 348 16842 382
rect 17572 3850 17606 3884
rect 17784 3850 17818 3884
rect 17996 3850 18030 3884
rect 18208 3850 18242 3884
rect 18420 3850 18454 3884
rect 18632 3850 18666 3884
rect 17670 3668 17704 3702
rect 17882 3668 17916 3702
rect 18094 3668 18128 3702
rect 18306 3668 18340 3702
rect 18518 3668 18552 3702
rect 18730 3668 18764 3702
rect 17538 3070 17572 3104
rect 17894 3070 17928 3104
rect 18250 3070 18284 3104
rect 18606 3070 18640 3104
rect 18962 3070 18996 3104
rect 19318 3070 19352 3104
rect 19674 3070 19708 3104
rect 20030 3070 20064 3104
rect 20386 3070 20420 3104
rect 17716 2848 17750 2882
rect 18072 2848 18106 2882
rect 18428 2848 18462 2882
rect 18784 2848 18818 2882
rect 19140 2848 19174 2882
rect 19496 2848 19530 2882
rect 19852 2848 19886 2882
rect 20208 2848 20242 2882
rect 17538 2570 17572 2604
rect 17894 2570 17928 2604
rect 18250 2570 18284 2604
rect 18606 2570 18640 2604
rect 18962 2570 18996 2604
rect 19318 2570 19352 2604
rect 19674 2570 19708 2604
rect 20030 2570 20064 2604
rect 20386 2570 20420 2604
rect 17716 2348 17750 2382
rect 18072 2348 18106 2382
rect 18428 2348 18462 2382
rect 18784 2348 18818 2382
rect 19140 2348 19174 2382
rect 19496 2348 19530 2382
rect 19852 2348 19886 2382
rect 20208 2348 20242 2382
rect 17538 2070 17572 2104
rect 17894 2070 17928 2104
rect 18250 2070 18284 2104
rect 18606 2070 18640 2104
rect 18962 2070 18996 2104
rect 19318 2070 19352 2104
rect 19674 2070 19708 2104
rect 20030 2070 20064 2104
rect 20386 2070 20420 2104
rect 17716 1848 17750 1882
rect 18072 1848 18106 1882
rect 18428 1848 18462 1882
rect 18784 1848 18818 1882
rect 19140 1848 19174 1882
rect 19496 1848 19530 1882
rect 19852 1848 19886 1882
rect 20208 1848 20242 1882
rect 17538 1570 17572 1604
rect 17894 1570 17928 1604
rect 18250 1570 18284 1604
rect 18606 1570 18640 1604
rect 18962 1570 18996 1604
rect 19318 1570 19352 1604
rect 19674 1570 19708 1604
rect 20030 1570 20064 1604
rect 20386 1570 20420 1604
rect 17716 1348 17750 1382
rect 18072 1348 18106 1382
rect 18428 1348 18462 1382
rect 18784 1348 18818 1382
rect 19140 1348 19174 1382
rect 19496 1348 19530 1382
rect 19852 1348 19886 1382
rect 20208 1348 20242 1382
rect 17538 1070 17572 1104
rect 17894 1070 17928 1104
rect 18250 1070 18284 1104
rect 18606 1070 18640 1104
rect 18962 1070 18996 1104
rect 19318 1070 19352 1104
rect 19674 1070 19708 1104
rect 20030 1070 20064 1104
rect 20386 1070 20420 1104
rect 17716 848 17750 882
rect 18072 848 18106 882
rect 18428 848 18462 882
rect 18784 848 18818 882
rect 19140 848 19174 882
rect 19496 848 19530 882
rect 19852 848 19886 882
rect 20208 848 20242 882
rect 17538 570 17572 604
rect 17894 570 17928 604
rect 18250 570 18284 604
rect 18606 570 18640 604
rect 18962 570 18996 604
rect 19318 570 19352 604
rect 19674 570 19708 604
rect 20030 570 20064 604
rect 20386 570 20420 604
rect 17716 348 17750 382
rect 18072 348 18106 382
rect 18428 348 18462 382
rect 18784 348 18818 382
rect 19140 348 19174 382
rect 19496 348 19530 382
rect 19852 348 19886 382
rect 20208 348 20242 382
rect 7821 -313 20722 -264
<< metal1 >>
rect -1037 6672 13788 6712
rect -1037 6656 8958 6672
rect 9016 6670 13788 6672
rect 9016 6667 11644 6670
rect 9016 6656 10026 6667
rect 10084 6656 11644 6667
rect 11702 6667 13788 6670
rect 11702 6656 12712 6667
rect 12770 6656 13788 6667
rect -1037 6622 6727 6656
rect 13581 6622 13788 6656
rect -1037 6614 8958 6622
rect 9016 6614 10026 6622
rect -1037 6609 10026 6614
rect 10084 6612 11644 6622
rect 11702 6612 12712 6622
rect 10084 6609 12712 6612
rect 12770 6609 13788 6622
rect -1037 6584 13788 6609
rect 8770 6268 8780 6269
rect 8424 6262 8780 6268
rect 8838 6268 8848 6269
rect 8838 6262 10618 6268
rect 8424 6228 8436 6262
rect 8470 6228 8780 6262
rect 8838 6228 9148 6262
rect 9182 6228 9504 6262
rect 9538 6228 9860 6262
rect 9894 6228 10204 6262
rect 10262 6228 10572 6262
rect 10606 6228 10618 6262
rect 8424 6222 8780 6228
rect 8770 6211 8780 6222
rect 8838 6222 10204 6228
rect 8838 6211 8848 6222
rect 10194 6204 10204 6222
rect 10262 6222 10618 6228
rect 11110 6262 11466 6268
rect 11524 6263 13304 6268
rect 11524 6262 12890 6263
rect 12948 6262 13304 6263
rect 11110 6228 11122 6262
rect 11156 6228 11466 6262
rect 11524 6228 11834 6262
rect 11868 6228 12190 6262
rect 12224 6228 12546 6262
rect 12580 6228 12890 6262
rect 12948 6228 13258 6262
rect 13292 6228 13304 6262
rect 11110 6222 11466 6228
rect 10262 6204 10272 6222
rect 11456 6210 11466 6222
rect 11524 6222 12890 6228
rect 11524 6210 11534 6222
rect 12880 6205 12890 6222
rect 12948 6222 13304 6228
rect 12948 6205 12958 6222
rect 8948 6046 8958 6058
rect 8602 6040 8958 6046
rect 9016 6046 9026 6058
rect 10016 6046 10026 6058
rect 9016 6040 10026 6046
rect 10084 6046 10094 6058
rect 11634 6046 11644 6058
rect 10084 6040 10440 6046
rect 8602 6006 8614 6040
rect 8648 6006 8958 6040
rect 9016 6006 9326 6040
rect 9360 6006 9682 6040
rect 9716 6006 10026 6040
rect 10084 6006 10394 6040
rect 10428 6006 10440 6040
rect 8602 6000 8958 6006
rect 9016 6000 10026 6006
rect 10084 6000 10440 6006
rect 11288 6040 11644 6046
rect 11702 6046 11712 6058
rect 12702 6046 12712 6058
rect 11702 6040 12712 6046
rect 12770 6046 12780 6058
rect 12770 6040 13126 6046
rect 11288 6006 11300 6040
rect 11334 6006 11644 6040
rect 11702 6006 12012 6040
rect 12046 6006 12368 6040
rect 12402 6006 12712 6040
rect 12770 6006 13080 6040
rect 13114 6006 13126 6040
rect 11288 6000 11644 6006
rect 11702 6000 12712 6006
rect 12770 6000 13126 6006
rect 8568 5945 10511 5947
rect 7518 5776 8069 5893
rect 8182 5776 8192 5893
rect 8491 5745 8501 5945
rect 8580 5944 10511 5945
rect 8580 5913 10538 5944
rect 11229 5937 13172 5947
rect 8580 5778 8590 5913
rect 10462 5874 10538 5913
rect 11190 5936 13172 5937
rect 11190 5913 13224 5936
rect 11190 5874 11266 5913
rect 10461 5816 10471 5874
rect 10529 5816 10539 5874
rect 11190 5816 11200 5874
rect 11258 5816 11268 5874
rect 10462 5778 10538 5816
rect 8580 5759 10538 5778
rect 11190 5777 11266 5816
rect 13148 5777 13224 5913
rect 8580 5745 10512 5759
rect 11190 5752 13224 5777
rect 8560 5744 10512 5745
rect 11234 5751 13224 5752
rect 11234 5743 13177 5751
rect 9416 5691 9426 5695
rect 8424 5685 8780 5691
rect 8838 5685 9426 5691
rect 9618 5691 9628 5695
rect 9618 5685 10204 5691
rect 10262 5685 10618 5691
rect 12102 5690 12112 5697
rect 8424 5651 8436 5685
rect 8470 5651 8780 5685
rect 8838 5651 9148 5685
rect 9182 5651 9426 5685
rect 9618 5651 9860 5685
rect 9894 5651 10204 5685
rect 10262 5651 10572 5685
rect 10606 5651 10618 5685
rect 8424 5645 8780 5651
rect 8770 5633 8780 5645
rect 8838 5645 9426 5651
rect 8838 5633 8848 5645
rect 9416 5637 9426 5645
rect 9618 5645 10204 5651
rect 9618 5637 9628 5645
rect 9482 5633 9492 5637
rect 9550 5633 9560 5637
rect 10194 5633 10204 5645
rect 10262 5645 10618 5651
rect 11110 5684 11466 5690
rect 11524 5684 12112 5690
rect 12304 5690 12314 5697
rect 12304 5684 12890 5690
rect 12948 5684 13304 5690
rect 11110 5650 11122 5684
rect 11156 5650 11466 5684
rect 11524 5650 11834 5684
rect 11868 5650 12112 5684
rect 12304 5650 12546 5684
rect 12580 5650 12890 5684
rect 12948 5650 13258 5684
rect 13292 5650 13304 5684
rect 10262 5633 10272 5645
rect 11110 5644 11466 5650
rect 11456 5632 11466 5644
rect 11524 5644 12112 5650
rect 11524 5632 11534 5644
rect 12102 5639 12112 5644
rect 12304 5644 12890 5650
rect 12304 5639 12314 5644
rect 12168 5632 12178 5639
rect 12236 5632 12246 5639
rect 12880 5632 12890 5644
rect 12948 5644 13304 5650
rect 12948 5632 12958 5644
rect 8948 5469 8958 5481
rect 8602 5463 8958 5469
rect 9016 5469 9026 5481
rect 10016 5469 10026 5481
rect 9016 5463 10026 5469
rect 10084 5469 10094 5481
rect 10084 5463 10440 5469
rect 11634 5468 11644 5480
rect 8602 5429 8614 5463
rect 8648 5429 8958 5463
rect 9016 5429 9326 5463
rect 9360 5429 9682 5463
rect 9716 5429 10026 5463
rect 10084 5429 10394 5463
rect 10428 5429 10440 5463
rect 8602 5423 8958 5429
rect 9016 5423 10026 5429
rect 10084 5423 10440 5429
rect 11288 5462 11644 5468
rect 11702 5468 11712 5480
rect 12702 5468 12712 5480
rect 11702 5462 12712 5468
rect 12770 5468 12780 5480
rect 12770 5462 13126 5468
rect 11288 5428 11300 5462
rect 11334 5428 11644 5462
rect 11702 5428 12012 5462
rect 12046 5428 12368 5462
rect 12402 5428 12712 5462
rect 12770 5428 13080 5462
rect 13114 5428 13126 5462
rect 11288 5422 11644 5428
rect 11702 5422 12712 5428
rect 12770 5422 13126 5428
rect 7617 5010 11266 5127
rect 10462 4903 10538 5010
rect 11190 4897 11266 5010
rect 8924 4863 9645 4897
rect 9762 4863 10512 4897
rect 11190 4864 11969 4897
rect 11229 4863 11969 4864
rect 12086 4863 12817 4897
rect 8770 4752 8780 4810
rect 8838 4804 10560 4810
rect 8838 4770 9148 4804
rect 9182 4770 9504 4804
rect 9538 4770 9860 4804
rect 9894 4770 10216 4804
rect 10250 4770 10560 4804
rect 8838 4764 10560 4770
rect 8838 4752 8848 4764
rect 10550 4752 10560 4764
rect 10618 4752 10628 4810
rect 11100 4752 11110 4810
rect 11168 4804 12890 4810
rect 11168 4770 11478 4804
rect 11512 4770 11834 4804
rect 11868 4770 12190 4804
rect 12224 4770 12546 4804
rect 12580 4770 12890 4804
rect 11168 4764 12890 4770
rect 11168 4752 11178 4764
rect 12880 4752 12890 4764
rect 12948 4752 12958 4810
rect 8948 4542 8958 4600
rect 9016 4588 9026 4600
rect 9482 4597 9492 4600
rect 9550 4597 9560 4600
rect 9420 4588 9430 4597
rect 9016 4582 9430 4588
rect 9016 4548 9326 4582
rect 9360 4548 9430 4582
rect 9016 4542 9430 4548
rect 9420 4539 9430 4542
rect 9622 4588 9632 4597
rect 10372 4588 10382 4600
rect 9622 4582 10382 4588
rect 9622 4548 9682 4582
rect 9716 4548 10038 4582
rect 10072 4548 10382 4582
rect 9622 4542 10382 4548
rect 10440 4542 10450 4600
rect 11278 4542 11288 4600
rect 11346 4588 11356 4600
rect 12168 4596 12178 4600
rect 12236 4596 12246 4600
rect 12099 4588 12109 4596
rect 11346 4582 12109 4588
rect 11346 4548 11656 4582
rect 11690 4548 12012 4582
rect 12046 4548 12109 4582
rect 11346 4542 12109 4548
rect 9622 4539 9632 4542
rect 12099 4538 12109 4542
rect 12301 4588 12311 4596
rect 12702 4588 12712 4600
rect 12301 4582 12712 4588
rect 12301 4548 12368 4582
rect 12402 4548 12712 4582
rect 12301 4542 12712 4548
rect 12770 4542 12780 4600
rect 12301 4538 12311 4542
rect 8860 4327 8936 4484
rect 10462 4327 10538 4483
rect 8860 4299 10538 4327
rect 8913 4298 10538 4299
rect 11190 4327 11266 4479
rect 12792 4327 12868 4485
rect 11190 4300 12868 4327
rect 8913 4293 10501 4298
rect 11190 4294 12832 4300
rect 11244 4293 12832 4294
rect 9418 4240 9428 4241
rect 8770 4182 8780 4240
rect 8838 4234 9428 4240
rect 9620 4240 9630 4241
rect 12099 4240 12109 4242
rect 9620 4234 10560 4240
rect 8838 4200 9148 4234
rect 9182 4200 9428 4234
rect 9620 4200 9860 4234
rect 9894 4200 10216 4234
rect 10250 4200 10560 4234
rect 8838 4194 9428 4200
rect 8838 4182 8848 4194
rect 9418 4183 9428 4194
rect 9620 4194 10560 4200
rect 9620 4183 9630 4194
rect 9480 4182 9490 4183
rect 9548 4182 9558 4183
rect 10550 4182 10560 4194
rect 10618 4182 10628 4240
rect 11100 4182 11110 4240
rect 11168 4234 12109 4240
rect 12301 4240 12311 4242
rect 12301 4234 12890 4240
rect 11168 4200 11478 4234
rect 11512 4200 11834 4234
rect 11868 4200 12109 4234
rect 12301 4200 12546 4234
rect 12580 4200 12890 4234
rect 11168 4194 12109 4200
rect 11168 4182 11178 4194
rect 12099 4184 12109 4194
rect 12301 4194 12890 4200
rect 12301 4184 12311 4194
rect 12168 4182 12178 4184
rect 12236 4182 12246 4184
rect 12880 4182 12890 4194
rect 12948 4182 12958 4240
rect 8948 3972 8958 4030
rect 9016 4018 9026 4030
rect 10372 4018 10382 4030
rect 9016 4012 10382 4018
rect 9016 3978 9326 4012
rect 9360 3978 9682 4012
rect 9716 3978 10038 4012
rect 10072 3978 10382 4012
rect 9016 3972 10382 3978
rect 10440 3972 10450 4030
rect 11278 3972 11288 4030
rect 11346 4018 11356 4030
rect 12702 4018 12712 4030
rect 11346 4012 12712 4018
rect 11346 3978 11656 4012
rect 11690 3978 12012 4012
rect 12046 3978 12368 4012
rect 12402 3978 12712 4012
rect 11346 3972 12712 3978
rect 12770 3972 12780 4030
rect 16250 3984 16306 4783
rect 16349 3984 16359 3986
rect 15825 3928 16359 3984
rect 16417 3984 16427 3986
rect 18033 3984 18089 4783
rect 18129 3984 18139 3986
rect 16417 3928 16739 3984
rect 17097 3928 17163 3984
rect 17605 3928 18139 3984
rect 18197 3984 18207 3986
rect 18197 3928 18519 3984
rect 18877 3928 18943 3984
rect 16723 3890 16733 3893
rect 15780 3884 16733 3890
rect 15780 3850 15792 3884
rect 15826 3850 16004 3884
rect 16038 3850 16216 3884
rect 16250 3850 16428 3884
rect 16462 3850 16640 3884
rect 16674 3850 16733 3884
rect 15780 3844 16733 3850
rect 16723 3839 16733 3844
rect 16898 3839 16908 3893
rect 17447 3838 17457 3892
rect 17622 3890 17632 3892
rect 17622 3884 18678 3890
rect 17622 3850 17784 3884
rect 17818 3850 17996 3884
rect 18030 3850 18208 3884
rect 18242 3850 18420 3884
rect 18454 3850 18632 3884
rect 18666 3850 18678 3884
rect 17622 3844 18678 3850
rect 17622 3838 17632 3844
rect 7687 3673 11265 3790
rect 10460 3388 10536 3673
rect 8566 3358 10536 3388
rect 11189 3388 11265 3673
rect 15866 3662 15876 3716
rect 16142 3708 16152 3716
rect 18494 3708 18504 3714
rect 16142 3702 16996 3708
rect 16142 3668 16314 3702
rect 16348 3668 16526 3702
rect 16560 3668 16738 3702
rect 16772 3668 16950 3702
rect 16984 3668 16996 3702
rect 16142 3662 16996 3668
rect 17658 3702 18504 3708
rect 17658 3668 17670 3702
rect 17704 3668 17882 3702
rect 17916 3668 18094 3702
rect 18128 3668 18306 3702
rect 18340 3668 18504 3702
rect 17658 3662 18504 3668
rect 18494 3660 18504 3662
rect 18770 3660 18780 3714
rect 16349 3624 16359 3626
rect 15613 3568 15679 3624
rect 16037 3568 16359 3624
rect 16417 3624 16427 3626
rect 18129 3624 18139 3626
rect 16417 3568 16951 3624
rect 17393 3568 17459 3624
rect 17817 3568 18139 3624
rect 18197 3624 18207 3626
rect 18197 3568 18731 3624
rect 11189 3369 13211 3388
rect 8566 3354 10524 3358
rect 11253 3354 13211 3369
rect 9410 3310 9420 3311
rect 8412 3252 8422 3310
rect 8480 3304 9420 3310
rect 9612 3310 9622 3311
rect 9612 3304 10558 3310
rect 8480 3270 8790 3304
rect 8824 3270 9146 3304
rect 9180 3270 9420 3304
rect 9612 3270 9858 3304
rect 9892 3270 10214 3304
rect 10248 3270 10558 3304
rect 8480 3264 9420 3270
rect 8480 3252 8490 3264
rect 9410 3253 9420 3264
rect 9612 3264 10558 3270
rect 9612 3253 9622 3264
rect 9480 3252 9490 3253
rect 9548 3252 9558 3253
rect 10548 3252 10558 3264
rect 10616 3252 10626 3310
rect 11099 3252 11109 3310
rect 11167 3304 12116 3310
rect 12308 3304 13245 3310
rect 11167 3270 11477 3304
rect 11511 3270 11833 3304
rect 11867 3270 12116 3304
rect 12308 3270 12545 3304
rect 12579 3270 12901 3304
rect 12935 3270 13245 3304
rect 11167 3264 12116 3270
rect 11167 3252 11177 3264
rect 12106 3252 12116 3264
rect 12308 3264 13245 3270
rect 12308 3252 12318 3264
rect 13235 3252 13245 3264
rect 13303 3252 13313 3310
rect 20276 3188 20352 3419
rect 14218 3154 16940 3188
rect 17664 3154 19030 3188
rect 19106 3155 20352 3188
rect 19106 3154 20346 3155
rect 15864 3110 15874 3113
rect 8946 3088 8956 3100
rect 8600 3082 8956 3088
rect 9014 3088 9024 3100
rect 10014 3088 10024 3100
rect 9014 3082 10024 3088
rect 10082 3088 10092 3100
rect 11633 3088 11643 3100
rect 10082 3082 10438 3088
rect 8600 3048 8612 3082
rect 8646 3048 8956 3082
rect 9014 3048 9324 3082
rect 9358 3048 9680 3082
rect 9714 3048 10024 3082
rect 10082 3048 10392 3082
rect 10426 3048 10438 3082
rect 8600 3042 8956 3048
rect 9014 3042 10024 3048
rect 10082 3042 10438 3048
rect 11287 3082 11643 3088
rect 11701 3088 11711 3100
rect 12701 3088 12711 3100
rect 11701 3082 12711 3088
rect 12769 3088 12779 3100
rect 12769 3082 13125 3088
rect 11287 3048 11299 3082
rect 11333 3048 11643 3082
rect 11701 3048 12011 3082
rect 12045 3048 12367 3082
rect 12401 3048 12711 3082
rect 12769 3048 13079 3082
rect 13113 3048 13125 3082
rect 14116 3052 14126 3110
rect 14184 3104 15550 3110
rect 14184 3070 14494 3104
rect 14528 3070 14850 3104
rect 14884 3070 15206 3104
rect 15240 3070 15550 3104
rect 14184 3064 15550 3070
rect 14184 3052 14194 3064
rect 15540 3052 15550 3064
rect 15608 3064 15874 3110
rect 16140 3110 16150 3113
rect 16140 3104 16974 3110
rect 16140 3070 16274 3104
rect 16308 3070 16630 3104
rect 16664 3070 16974 3104
rect 15608 3052 15618 3064
rect 15864 3059 15874 3064
rect 16140 3064 16974 3070
rect 16140 3059 16150 3064
rect 16964 3052 16974 3064
rect 17032 3064 17526 3110
rect 17584 3104 18504 3110
rect 17584 3070 17894 3104
rect 17928 3070 18250 3104
rect 18284 3070 18504 3104
rect 17032 3052 17042 3064
rect 17516 3052 17526 3064
rect 17584 3064 18504 3070
rect 17584 3052 17594 3064
rect 18494 3056 18504 3064
rect 18770 3064 18950 3110
rect 19008 3104 20374 3110
rect 19008 3070 19318 3104
rect 19352 3070 19674 3104
rect 19708 3070 20030 3104
rect 20064 3070 20374 3104
rect 18770 3056 18780 3064
rect 18940 3052 18950 3064
rect 19008 3064 20374 3070
rect 19008 3052 19018 3064
rect 20364 3052 20374 3064
rect 20432 3052 20442 3110
rect 11287 3042 11643 3048
rect 11701 3042 12711 3048
rect 12769 3042 13125 3048
rect 8502 2888 8578 2986
rect 10460 2888 10536 2985
rect 8502 2863 10536 2888
rect 11189 2888 11265 2986
rect 13147 2888 13223 2985
rect 15006 2888 15016 2900
rect 11189 2863 13223 2888
rect 8566 2862 10536 2863
rect 11253 2862 13223 2863
rect 14304 2882 15016 2888
rect 15074 2888 15084 2900
rect 16074 2888 16084 2900
rect 15074 2882 16084 2888
rect 16142 2888 16152 2900
rect 18406 2888 18416 2900
rect 16142 2882 16854 2888
rect 8566 2854 10519 2862
rect 11253 2854 13206 2862
rect 14304 2848 14316 2882
rect 14350 2848 14672 2882
rect 14706 2848 15016 2882
rect 15074 2848 15384 2882
rect 15418 2848 15740 2882
rect 15774 2848 16084 2882
rect 16142 2848 16452 2882
rect 16486 2848 16808 2882
rect 16842 2848 16854 2882
rect 14304 2842 15016 2848
rect 15074 2842 16084 2848
rect 16142 2842 16854 2848
rect 17704 2882 18416 2888
rect 18474 2888 18484 2900
rect 19474 2888 19484 2900
rect 18474 2882 19484 2888
rect 19542 2888 19552 2900
rect 19542 2882 20254 2888
rect 17704 2848 17716 2882
rect 17750 2848 18072 2882
rect 18106 2848 18416 2882
rect 18474 2848 18784 2882
rect 18818 2848 19140 2882
rect 19174 2848 19484 2882
rect 19542 2848 19852 2882
rect 19886 2848 20208 2882
rect 20242 2848 20254 2882
rect 17704 2842 18416 2848
rect 18474 2842 19484 2848
rect 19542 2842 20254 2848
rect 8412 2752 8422 2810
rect 8480 2804 9490 2810
rect 9548 2804 10558 2810
rect 8480 2770 8790 2804
rect 8824 2770 9146 2804
rect 9180 2770 9490 2804
rect 9548 2770 9858 2804
rect 9892 2770 10214 2804
rect 10248 2770 10558 2804
rect 8480 2764 9490 2770
rect 8480 2752 8490 2764
rect 9480 2752 9490 2764
rect 9548 2764 10558 2770
rect 9548 2752 9558 2764
rect 10548 2752 10558 2764
rect 10616 2752 10626 2810
rect 11099 2752 11109 2810
rect 11167 2804 12177 2810
rect 12235 2804 13245 2810
rect 11167 2770 11477 2804
rect 11511 2770 11833 2804
rect 11867 2770 12177 2804
rect 12235 2770 12545 2804
rect 12579 2770 12901 2804
rect 12935 2770 13245 2804
rect 11167 2764 12177 2770
rect 11167 2752 11177 2764
rect 12167 2752 12177 2764
rect 12235 2764 13245 2770
rect 12235 2752 12245 2764
rect 13235 2752 13245 2764
rect 13303 2752 13313 2810
rect 6105 2253 6163 2704
rect 14206 2691 14282 2765
rect 16876 2690 16952 2767
rect 17606 2690 17682 2770
rect 20276 2689 20352 2771
rect 14270 2654 16940 2688
rect 17660 2654 20342 2688
rect 8946 2588 8956 2600
rect 8600 2582 8956 2588
rect 9014 2588 9024 2600
rect 10014 2588 10024 2600
rect 9014 2582 10024 2588
rect 10082 2588 10092 2600
rect 11633 2588 11643 2600
rect 10082 2582 10438 2588
rect 8600 2548 8612 2582
rect 8646 2548 8956 2582
rect 9014 2548 9324 2582
rect 9358 2548 9680 2582
rect 9714 2548 10024 2582
rect 10082 2548 10392 2582
rect 10426 2548 10438 2582
rect 8600 2542 8956 2548
rect 9014 2542 10024 2548
rect 10082 2542 10438 2548
rect 11287 2582 11643 2588
rect 11701 2588 11711 2600
rect 12701 2588 12711 2600
rect 11701 2582 12711 2588
rect 12769 2588 12779 2600
rect 12769 2582 13125 2588
rect 11287 2548 11299 2582
rect 11333 2548 11643 2582
rect 11701 2548 12011 2582
rect 12045 2548 12367 2582
rect 12401 2548 12711 2582
rect 12769 2548 13079 2582
rect 13113 2548 13125 2582
rect 14116 2552 14126 2610
rect 14184 2604 15550 2610
rect 15608 2604 16974 2610
rect 14184 2570 14494 2604
rect 14528 2570 14850 2604
rect 14884 2570 15206 2604
rect 15240 2570 15550 2604
rect 15608 2570 15918 2604
rect 15952 2570 16274 2604
rect 16308 2570 16630 2604
rect 16664 2570 16974 2604
rect 14184 2564 15550 2570
rect 14184 2552 14194 2564
rect 15540 2552 15550 2564
rect 15608 2564 16974 2570
rect 15608 2552 15618 2564
rect 16964 2552 16974 2564
rect 17032 2552 17042 2610
rect 17516 2552 17526 2610
rect 17584 2604 18950 2610
rect 19008 2604 20374 2610
rect 17584 2570 17894 2604
rect 17928 2570 18250 2604
rect 18284 2570 18606 2604
rect 18640 2570 18950 2604
rect 19008 2570 19318 2604
rect 19352 2570 19674 2604
rect 19708 2570 20030 2604
rect 20064 2570 20374 2604
rect 17584 2564 18950 2570
rect 17584 2552 17594 2564
rect 18940 2552 18950 2564
rect 19008 2564 20374 2570
rect 19008 2552 19018 2564
rect 20364 2552 20374 2564
rect 20432 2552 20442 2610
rect 11287 2542 11643 2548
rect 11701 2542 12711 2548
rect 12769 2542 13125 2548
rect 8502 2388 8578 2481
rect 10460 2388 10536 2490
rect 8502 2367 10536 2388
rect 11189 2388 11265 2481
rect 13147 2388 13223 2490
rect 15006 2388 15016 2401
rect 11189 2367 13223 2388
rect 14304 2382 15016 2388
rect 15074 2388 15084 2401
rect 16074 2388 16084 2400
rect 15074 2382 16084 2388
rect 16142 2388 16152 2400
rect 18406 2388 18416 2400
rect 16142 2382 16854 2388
rect 8502 2358 10497 2367
rect 11189 2358 13184 2367
rect 8544 2354 10497 2358
rect 11231 2354 13184 2358
rect 14304 2348 14316 2382
rect 14350 2348 14672 2382
rect 14706 2348 15016 2382
rect 15074 2348 15384 2382
rect 15418 2348 15740 2382
rect 15774 2348 16084 2382
rect 16142 2348 16452 2382
rect 16486 2348 16808 2382
rect 16842 2348 16854 2382
rect 14304 2343 15016 2348
rect 15074 2343 16084 2348
rect 14304 2342 16084 2343
rect 16142 2342 16854 2348
rect 17704 2382 18416 2388
rect 18474 2388 18484 2400
rect 19474 2388 19484 2400
rect 18474 2382 19484 2388
rect 19542 2388 19552 2400
rect 19542 2382 20254 2388
rect 17704 2348 17716 2382
rect 17750 2348 18072 2382
rect 18106 2348 18416 2382
rect 18474 2348 18784 2382
rect 18818 2348 19140 2382
rect 19174 2348 19484 2382
rect 19542 2348 19852 2382
rect 19886 2348 20208 2382
rect 20242 2348 20254 2382
rect 17704 2342 18416 2348
rect 18474 2342 19484 2348
rect 19542 2342 20254 2348
rect 8412 2252 8422 2310
rect 8480 2304 9490 2310
rect 9548 2304 10558 2310
rect 8480 2270 8790 2304
rect 8824 2270 9146 2304
rect 9180 2270 9490 2304
rect 9548 2270 9858 2304
rect 9892 2270 10214 2304
rect 10248 2270 10558 2304
rect 8480 2264 9490 2270
rect 8480 2252 8490 2264
rect 9480 2252 9490 2264
rect 9548 2264 10558 2270
rect 9548 2252 9558 2264
rect 10548 2252 10558 2264
rect 10616 2252 10626 2310
rect 11099 2252 11109 2310
rect 11167 2304 12177 2310
rect 12235 2304 13245 2310
rect 11167 2270 11477 2304
rect 11511 2270 11833 2304
rect 11867 2270 12177 2304
rect 12235 2270 12545 2304
rect 12579 2270 12901 2304
rect 12935 2270 13245 2304
rect 11167 2264 12177 2270
rect 11167 2252 11177 2264
rect 12167 2252 12177 2264
rect 12235 2264 13245 2270
rect 12235 2252 12245 2264
rect 13235 2252 13245 2264
rect 13303 2252 13313 2310
rect 14206 2188 14282 2265
rect 16876 2191 16952 2268
rect 17606 2191 17682 2271
rect 20276 2188 20352 2270
rect 14257 2154 16939 2188
rect 17660 2154 20342 2188
rect 8946 2088 8956 2100
rect 8600 2082 8956 2088
rect 9014 2088 9024 2100
rect 9302 2092 9380 2100
rect 9270 2091 9482 2092
rect 9264 2088 9274 2091
rect 8600 2048 8612 2082
rect 8646 2048 8956 2082
rect 8600 2042 8956 2048
rect 9014 2042 9274 2088
rect 9480 2088 9490 2091
rect 10014 2088 10024 2100
rect 9480 2082 10024 2088
rect 10082 2088 10092 2100
rect 11633 2088 11643 2100
rect 10082 2082 10438 2088
rect 9480 2048 9680 2082
rect 9714 2048 10024 2082
rect 10082 2048 10392 2082
rect 10426 2048 10438 2082
rect 9264 2033 9274 2042
rect 9480 2042 10024 2048
rect 10082 2042 10438 2048
rect 11287 2082 11643 2088
rect 11701 2088 11711 2100
rect 12226 2091 12438 2096
rect 12216 2088 12226 2091
rect 11701 2082 12226 2088
rect 12417 2088 12438 2091
rect 12701 2088 12711 2100
rect 11287 2048 11299 2082
rect 11333 2048 11643 2082
rect 11701 2048 12011 2082
rect 12045 2048 12226 2082
rect 11287 2042 11643 2048
rect 11701 2042 12226 2048
rect 9480 2033 9490 2042
rect 12216 2038 12226 2042
rect 12417 2042 12711 2088
rect 12769 2088 12779 2100
rect 12769 2082 13125 2088
rect 12769 2048 13079 2082
rect 13113 2048 13125 2082
rect 14116 2052 14126 2110
rect 14184 2104 15550 2110
rect 15608 2104 16974 2110
rect 14184 2070 14494 2104
rect 14528 2070 14850 2104
rect 14884 2070 15206 2104
rect 15240 2070 15550 2104
rect 15608 2070 15918 2104
rect 15952 2070 16274 2104
rect 16308 2070 16630 2104
rect 16664 2070 16974 2104
rect 14184 2064 15550 2070
rect 14184 2052 14194 2064
rect 15540 2052 15550 2064
rect 15608 2064 16974 2070
rect 15608 2052 15618 2064
rect 16964 2052 16974 2064
rect 17032 2052 17042 2110
rect 17516 2052 17526 2110
rect 17584 2104 18950 2110
rect 19008 2104 20374 2110
rect 17584 2070 17894 2104
rect 17928 2070 18250 2104
rect 18284 2070 18606 2104
rect 18640 2070 18950 2104
rect 19008 2070 19318 2104
rect 19352 2070 19674 2104
rect 19708 2070 20030 2104
rect 20064 2070 20374 2104
rect 17584 2064 18950 2070
rect 17584 2052 17594 2064
rect 18940 2052 18950 2064
rect 19008 2064 20374 2070
rect 19008 2052 19018 2064
rect 20364 2052 20374 2064
rect 20432 2052 20442 2110
rect 12769 2042 13125 2048
rect 12417 2038 12438 2042
rect 15006 1888 15016 1900
rect 14304 1882 15016 1888
rect 15074 1888 15084 1900
rect 16074 1888 16084 1900
rect 15074 1882 16084 1888
rect 16142 1888 16152 1900
rect 18406 1888 18416 1900
rect 16142 1882 16854 1888
rect 14304 1848 14316 1882
rect 14350 1848 14672 1882
rect 14706 1848 15016 1882
rect 15074 1848 15384 1882
rect 15418 1848 15740 1882
rect 15774 1848 16084 1882
rect 16142 1848 16452 1882
rect 16486 1848 16808 1882
rect 16842 1848 16854 1882
rect 14304 1842 15016 1848
rect 15074 1842 16084 1848
rect 16142 1842 16854 1848
rect 17704 1882 18416 1888
rect 18474 1888 18484 1900
rect 19474 1888 19484 1900
rect 18474 1882 19484 1888
rect 19542 1888 19552 1900
rect 19542 1882 20254 1888
rect 17704 1848 17716 1882
rect 17750 1848 18072 1882
rect 18106 1848 18416 1882
rect 18474 1848 18784 1882
rect 18818 1848 19140 1882
rect 19174 1848 19484 1882
rect 19542 1848 19852 1882
rect 19886 1848 20208 1882
rect 20242 1848 20254 1882
rect 17704 1842 18416 1848
rect 18474 1842 19484 1848
rect 19542 1842 20254 1848
rect 14206 1689 14282 1766
rect 16876 1691 16952 1768
rect 17606 1690 17682 1770
rect 20276 1689 20352 1771
rect 8566 1654 10524 1688
rect 11253 1654 13211 1688
rect 14253 1654 16935 1688
rect 17659 1654 20341 1688
rect 9308 1610 9318 1611
rect 9524 1610 9534 1611
rect 12159 1610 12169 1611
rect 8412 1552 8422 1610
rect 8480 1604 9318 1610
rect 9548 1604 10558 1610
rect 8480 1570 8790 1604
rect 8824 1570 9146 1604
rect 9180 1570 9318 1604
rect 9548 1570 9858 1604
rect 9892 1570 10214 1604
rect 10248 1570 10558 1604
rect 8480 1564 9318 1570
rect 8480 1552 8490 1564
rect 9281 1552 9318 1564
rect 9548 1564 10558 1570
rect 9548 1552 9558 1564
rect 10548 1552 10558 1564
rect 10616 1552 10626 1610
rect 11099 1552 11109 1610
rect 11167 1604 12169 1610
rect 12433 1610 12443 1611
rect 12433 1604 13245 1610
rect 11167 1570 11477 1604
rect 11511 1570 11833 1604
rect 11867 1570 12169 1604
rect 12433 1570 12545 1604
rect 12579 1570 12901 1604
rect 12935 1570 13245 1604
rect 11167 1564 12169 1570
rect 11167 1552 11177 1564
rect 12159 1552 12169 1564
rect 12433 1564 13245 1570
rect 12433 1552 12443 1564
rect 13235 1552 13245 1564
rect 13303 1552 13313 1610
rect 14116 1552 14126 1610
rect 14184 1604 15550 1610
rect 15608 1604 16974 1610
rect 14184 1570 14494 1604
rect 14528 1570 14850 1604
rect 14884 1570 15206 1604
rect 15240 1570 15550 1604
rect 15608 1570 15918 1604
rect 15952 1570 16274 1604
rect 16308 1570 16630 1604
rect 16664 1570 16974 1604
rect 14184 1564 15550 1570
rect 14184 1552 14194 1564
rect 15540 1552 15550 1564
rect 15608 1564 16974 1570
rect 15608 1552 15618 1564
rect 16964 1552 16974 1564
rect 17032 1552 17042 1610
rect 17516 1552 17526 1610
rect 17584 1604 18950 1610
rect 19008 1604 20374 1610
rect 17584 1570 17894 1604
rect 17928 1570 18250 1604
rect 18284 1570 18606 1604
rect 18640 1570 18950 1604
rect 19008 1570 19318 1604
rect 19352 1570 19674 1604
rect 19708 1570 20030 1604
rect 20064 1570 20374 1604
rect 17584 1564 18950 1570
rect 17584 1552 17594 1564
rect 18940 1552 18950 1564
rect 19008 1564 20374 1570
rect 19008 1552 19018 1564
rect 20364 1552 20374 1564
rect 20432 1552 20442 1610
rect 9308 1551 9318 1552
rect 9524 1551 9534 1552
rect 8946 1388 8956 1400
rect 8600 1382 8956 1388
rect 9014 1388 9024 1400
rect 10014 1388 10024 1400
rect 9014 1382 10024 1388
rect 10082 1388 10092 1400
rect 11633 1388 11643 1400
rect 10082 1382 10438 1388
rect 8600 1348 8612 1382
rect 8646 1348 8956 1382
rect 9014 1348 9324 1382
rect 9358 1348 9680 1382
rect 9714 1348 10024 1382
rect 10082 1348 10392 1382
rect 10426 1348 10438 1382
rect 8600 1342 8956 1348
rect 9014 1342 10024 1348
rect 10082 1342 10438 1348
rect 11287 1382 11643 1388
rect 11701 1388 11711 1400
rect 12701 1388 12711 1400
rect 11701 1382 12711 1388
rect 12769 1388 12779 1400
rect 15006 1388 15016 1400
rect 12769 1382 13125 1388
rect 11287 1348 11299 1382
rect 11333 1348 11643 1382
rect 11701 1348 12011 1382
rect 12045 1348 12367 1382
rect 12401 1348 12711 1382
rect 12769 1348 13079 1382
rect 13113 1348 13125 1382
rect 11287 1342 11643 1348
rect 11701 1342 12711 1348
rect 12769 1342 13125 1348
rect 14304 1382 15016 1388
rect 15074 1388 15084 1400
rect 16074 1388 16084 1400
rect 15074 1382 16084 1388
rect 16142 1388 16152 1400
rect 18406 1388 18416 1400
rect 16142 1382 16854 1388
rect 14304 1348 14316 1382
rect 14350 1348 14672 1382
rect 14706 1348 15016 1382
rect 15074 1348 15384 1382
rect 15418 1348 15740 1382
rect 15774 1348 16084 1382
rect 16142 1348 16452 1382
rect 16486 1348 16808 1382
rect 16842 1348 16854 1382
rect 14304 1342 15016 1348
rect 15074 1342 16084 1348
rect 16142 1342 16854 1348
rect 17704 1382 18416 1388
rect 18474 1388 18484 1400
rect 19474 1388 19484 1400
rect 18474 1382 19484 1388
rect 19542 1388 19552 1400
rect 19542 1382 20254 1388
rect 17704 1348 17716 1382
rect 17750 1348 18072 1382
rect 18106 1348 18416 1382
rect 18474 1348 18784 1382
rect 18818 1348 19140 1382
rect 19174 1348 19484 1382
rect 19542 1348 19852 1382
rect 19886 1348 20208 1382
rect 20242 1348 20254 1382
rect 17704 1342 18416 1348
rect 18474 1342 19484 1348
rect 19542 1342 20254 1348
rect 8502 1188 8578 1286
rect 10460 1188 10536 1285
rect 8502 1163 10536 1188
rect 11189 1188 11265 1286
rect 13147 1188 13223 1285
rect 14206 1190 14282 1267
rect 16876 1190 16952 1267
rect 17606 1191 17682 1271
rect 20276 1189 20352 1271
rect 11189 1163 13223 1188
rect 8566 1162 10536 1163
rect 11253 1162 13223 1163
rect 8566 1154 10519 1162
rect 11253 1154 13206 1162
rect 14252 1154 16934 1188
rect 17662 1154 20344 1188
rect 8412 1052 8422 1110
rect 8480 1104 9490 1110
rect 9548 1104 10558 1110
rect 8480 1070 8790 1104
rect 8824 1070 9146 1104
rect 9180 1070 9490 1104
rect 9548 1070 9858 1104
rect 9892 1070 10214 1104
rect 10248 1070 10558 1104
rect 8480 1064 9490 1070
rect 8480 1052 8490 1064
rect 9480 1052 9490 1064
rect 9548 1064 10558 1070
rect 9548 1052 9558 1064
rect 10548 1052 10558 1064
rect 10616 1052 10626 1110
rect 11099 1052 11109 1110
rect 11167 1104 12177 1110
rect 12235 1104 13245 1110
rect 11167 1070 11477 1104
rect 11511 1070 11833 1104
rect 11867 1070 12177 1104
rect 12235 1070 12545 1104
rect 12579 1070 12901 1104
rect 12935 1070 13245 1104
rect 11167 1064 12177 1070
rect 11167 1052 11177 1064
rect 12167 1052 12177 1064
rect 12235 1064 13245 1070
rect 12235 1052 12245 1064
rect 13235 1052 13245 1064
rect 13303 1052 13313 1110
rect 14116 1052 14126 1110
rect 14184 1104 15550 1110
rect 15608 1104 16974 1110
rect 14184 1070 14494 1104
rect 14528 1070 14850 1104
rect 14884 1070 15206 1104
rect 15240 1070 15550 1104
rect 15608 1070 15918 1104
rect 15952 1070 16274 1104
rect 16308 1070 16630 1104
rect 16664 1070 16974 1104
rect 14184 1064 15550 1070
rect 14184 1052 14194 1064
rect 15540 1052 15550 1064
rect 15608 1064 16974 1070
rect 15608 1052 15618 1064
rect 16964 1052 16974 1064
rect 17032 1052 17042 1110
rect 17516 1052 17526 1110
rect 17584 1104 18950 1110
rect 19008 1104 20374 1110
rect 17584 1070 17894 1104
rect 17928 1070 18250 1104
rect 18284 1070 18606 1104
rect 18640 1070 18950 1104
rect 19008 1070 19318 1104
rect 19352 1070 19674 1104
rect 19708 1070 20030 1104
rect 20064 1070 20374 1104
rect 17584 1064 18950 1070
rect 17584 1052 17594 1064
rect 18940 1052 18950 1064
rect 19008 1064 20374 1070
rect 19008 1052 19018 1064
rect 20364 1052 20374 1064
rect 20432 1052 20442 1110
rect 8946 888 8956 900
rect -715 757 1417 885
rect 8600 882 8956 888
rect 9014 888 9024 900
rect 10014 888 10024 900
rect 9014 882 10024 888
rect 10082 888 10092 900
rect 11633 888 11643 900
rect 10082 882 10438 888
rect 8600 848 8612 882
rect 8646 848 8956 882
rect 9014 848 9324 882
rect 9358 848 9680 882
rect 9714 848 10024 882
rect 10082 848 10392 882
rect 10426 848 10438 882
rect 8600 842 8956 848
rect 9014 842 10024 848
rect 10082 842 10438 848
rect 11287 882 11643 888
rect 11701 888 11711 900
rect 12701 888 12711 900
rect 11701 882 12711 888
rect 12769 888 12779 900
rect 15006 888 15016 900
rect 12769 882 13125 888
rect 11287 848 11299 882
rect 11333 848 11643 882
rect 11701 848 12011 882
rect 12045 848 12367 882
rect 12401 848 12711 882
rect 12769 848 13079 882
rect 13113 848 13125 882
rect 11287 842 11643 848
rect 11701 842 12711 848
rect 12769 842 13125 848
rect 14304 882 15016 888
rect 15074 888 15084 900
rect 16074 888 16084 900
rect 15074 882 16084 888
rect 16142 888 16152 900
rect 18406 888 18416 900
rect 16142 882 16854 888
rect 14304 848 14316 882
rect 14350 848 14672 882
rect 14706 848 15016 882
rect 15074 848 15384 882
rect 15418 848 15740 882
rect 15774 848 16084 882
rect 16142 848 16452 882
rect 16486 848 16808 882
rect 16842 848 16854 882
rect 14304 842 15016 848
rect 15074 842 16084 848
rect 16142 842 16854 848
rect 17704 882 18416 888
rect 18474 888 18484 900
rect 19474 888 19484 900
rect 18474 882 19484 888
rect 19542 888 19552 900
rect 19542 882 20254 888
rect 17704 848 17716 882
rect 17750 848 18072 882
rect 18106 848 18416 882
rect 18474 848 18784 882
rect 18818 848 19140 882
rect 19174 848 19484 882
rect 19542 848 19852 882
rect 19886 848 20208 882
rect 20242 848 20254 882
rect 17704 842 18416 848
rect 18474 842 19484 848
rect 19542 842 20254 848
rect 8502 688 8578 781
rect 10460 688 10536 790
rect 8502 667 10536 688
rect 11189 688 11265 781
rect 13147 688 13223 790
rect 14206 690 14282 767
rect 16876 691 16952 768
rect 17606 690 17682 770
rect 20276 688 20352 770
rect 11189 667 13223 688
rect 8502 658 10497 667
rect 11189 658 13184 667
rect 8544 654 10497 658
rect 11231 654 13184 658
rect 14255 654 16937 688
rect 17659 654 20341 688
rect 8412 552 8422 610
rect 8480 604 9490 610
rect 9548 604 10558 610
rect 8480 570 8790 604
rect 8824 570 9146 604
rect 9180 570 9490 604
rect 9548 570 9858 604
rect 9892 570 10214 604
rect 10248 570 10558 604
rect 8480 564 9490 570
rect 8480 552 8490 564
rect 9480 552 9490 564
rect 9548 564 10558 570
rect 9548 552 9558 564
rect 10548 552 10558 564
rect 10616 552 10626 610
rect 11099 552 11109 610
rect 11167 604 12177 610
rect 12235 604 13245 610
rect 11167 570 11477 604
rect 11511 570 11833 604
rect 11867 570 12177 604
rect 12235 570 12545 604
rect 12579 570 12901 604
rect 12935 570 13245 604
rect 11167 564 12177 570
rect 11167 552 11177 564
rect 12167 552 12177 564
rect 12235 564 13245 570
rect 12235 552 12245 564
rect 13235 552 13245 564
rect 13303 552 13313 610
rect 14116 552 14126 610
rect 14184 604 15550 610
rect 15608 604 16974 610
rect 14184 570 14494 604
rect 14528 570 14850 604
rect 14884 570 15206 604
rect 15240 570 15550 604
rect 15608 570 15918 604
rect 15952 570 16274 604
rect 16308 570 16630 604
rect 16664 570 16974 604
rect 14184 564 15550 570
rect 14184 552 14194 564
rect 15540 552 15550 564
rect 15608 564 16974 570
rect 15608 552 15618 564
rect 16964 552 16974 564
rect 17032 564 17526 610
rect 17584 604 18950 610
rect 19008 604 20374 610
rect 17584 570 17894 604
rect 17928 570 18250 604
rect 18284 570 18606 604
rect 18640 570 18950 604
rect 19008 570 19318 604
rect 19352 570 19674 604
rect 19708 570 20030 604
rect 20064 570 20374 604
rect 17032 552 17042 564
rect 17516 552 17526 564
rect 17584 564 18950 570
rect 17584 552 17594 564
rect 18940 552 18950 564
rect 19008 564 20374 570
rect 19008 552 19018 564
rect 20364 552 20374 564
rect 20432 552 20442 610
rect 8946 388 8956 400
rect 8600 382 8956 388
rect 9014 388 9024 400
rect 10014 388 10024 400
rect 9014 382 10024 388
rect 10082 388 10092 400
rect 11633 388 11643 400
rect 10082 382 10438 388
rect 8600 348 8612 382
rect 8646 348 8956 382
rect 9014 348 9324 382
rect 9358 348 9680 382
rect 9714 348 10024 382
rect 10082 348 10392 382
rect 10426 348 10438 382
rect 8600 342 8956 348
rect 9014 342 10024 348
rect 10082 342 10438 348
rect 11287 382 11643 388
rect 11701 388 11711 400
rect 12701 388 12711 400
rect 11701 382 12711 388
rect 12769 388 12779 400
rect 15006 388 15016 400
rect 12769 382 13125 388
rect 11287 348 11299 382
rect 11333 348 11643 382
rect 11701 348 12011 382
rect 12045 348 12367 382
rect 12401 348 12711 382
rect 12769 348 13079 382
rect 13113 348 13125 382
rect 11287 342 11643 348
rect 11701 342 12711 348
rect 12769 342 13125 348
rect 14304 382 15016 388
rect 15074 388 15084 400
rect 16074 388 16084 400
rect 15074 382 16084 388
rect 16142 388 16152 400
rect 18406 388 18416 400
rect 16142 382 16854 388
rect 14304 348 14316 382
rect 14350 348 14672 382
rect 14706 348 15016 382
rect 15074 348 15384 382
rect 15418 348 15740 382
rect 15774 348 16084 382
rect 16142 348 16452 382
rect 16486 348 16808 382
rect 16842 348 16854 382
rect 14304 342 15016 348
rect 15074 342 16084 348
rect 16142 342 16854 348
rect 17704 382 18416 388
rect 18474 388 18484 400
rect 19474 388 19484 400
rect 18474 382 19484 388
rect 19542 388 19552 400
rect 19542 382 20254 388
rect 17704 348 17716 382
rect 17750 348 18072 382
rect 18106 348 18416 382
rect 18474 348 18784 382
rect 18818 348 19140 382
rect 19174 348 19484 382
rect 19542 348 19852 382
rect 19886 348 20208 382
rect 20242 348 20254 382
rect 17704 342 18416 348
rect 18474 342 19484 348
rect 19542 342 20254 348
rect 8560 264 10513 298
rect 11230 274 13183 298
rect 11188 264 13183 274
rect 14254 264 16936 298
rect 10460 75 10536 260
rect 11188 75 11264 264
rect 15630 75 15706 258
rect 7788 -42 15706 75
rect -1045 -194 20939 -186
rect -1045 -196 12671 -194
rect -1045 -213 9990 -196
rect -1045 -264 8929 -213
rect 9048 -264 9990 -213
rect 10116 -206 12671 -196
rect 10116 -264 11586 -206
rect 11753 -264 12671 -206
rect 12809 -196 16018 -194
rect 12809 -264 14955 -196
rect 15135 -264 16018 -196
rect 16208 -196 20939 -194
rect 16208 -264 18336 -196
rect 18526 -201 20939 -196
rect 18526 -264 19417 -201
rect 19607 -264 20939 -201
rect -1045 -313 7821 -264
rect 20722 -313 20939 -264
rect -1045 -314 11586 -313
rect 7809 -319 11586 -314
rect 11576 -322 11586 -319
rect 11753 -315 12671 -313
rect 12809 -314 20939 -313
rect 12809 -315 20734 -314
rect 11753 -319 20734 -315
rect 11753 -322 11763 -319
<< via1 >>
rect 8958 6656 9016 6672
rect 10026 6656 10084 6667
rect 11644 6656 11702 6670
rect 12712 6656 12770 6667
rect 8958 6622 9016 6656
rect 10026 6622 10084 6656
rect 11644 6622 11702 6656
rect 12712 6622 12770 6656
rect 8958 6614 9016 6622
rect 10026 6609 10084 6622
rect 11644 6612 11702 6622
rect 12712 6609 12770 6622
rect 8780 6262 8838 6269
rect 8780 6228 8792 6262
rect 8792 6228 8826 6262
rect 8826 6228 8838 6262
rect 10204 6228 10216 6262
rect 10216 6228 10250 6262
rect 10250 6228 10262 6262
rect 8780 6211 8838 6228
rect 10204 6204 10262 6228
rect 11466 6262 11524 6268
rect 12890 6262 12948 6263
rect 11466 6228 11478 6262
rect 11478 6228 11512 6262
rect 11512 6228 11524 6262
rect 12890 6228 12902 6262
rect 12902 6228 12936 6262
rect 12936 6228 12948 6262
rect 11466 6210 11524 6228
rect 12890 6205 12948 6228
rect 8958 6040 9016 6058
rect 10026 6040 10084 6058
rect 8958 6006 8970 6040
rect 8970 6006 9004 6040
rect 9004 6006 9016 6040
rect 10026 6006 10038 6040
rect 10038 6006 10072 6040
rect 10072 6006 10084 6040
rect 8958 6000 9016 6006
rect 10026 6000 10084 6006
rect 11644 6040 11702 6058
rect 12712 6040 12770 6058
rect 11644 6006 11656 6040
rect 11656 6006 11690 6040
rect 11690 6006 11702 6040
rect 12712 6006 12724 6040
rect 12724 6006 12758 6040
rect 12758 6006 12770 6040
rect 11644 6000 11702 6006
rect 12712 6000 12770 6006
rect 8069 5776 8182 5893
rect 8501 5745 8580 5945
rect 10471 5816 10529 5874
rect 11200 5816 11258 5874
rect 8780 5685 8838 5691
rect 9426 5685 9618 5695
rect 10204 5685 10262 5691
rect 8780 5651 8792 5685
rect 8792 5651 8826 5685
rect 8826 5651 8838 5685
rect 9426 5651 9504 5685
rect 9504 5651 9538 5685
rect 9538 5651 9618 5685
rect 10204 5651 10216 5685
rect 10216 5651 10250 5685
rect 10250 5651 10262 5685
rect 8780 5633 8838 5651
rect 9426 5637 9618 5651
rect 9492 5633 9550 5637
rect 10204 5633 10262 5651
rect 11466 5684 11524 5690
rect 12112 5684 12304 5697
rect 12890 5684 12948 5690
rect 11466 5650 11478 5684
rect 11478 5650 11512 5684
rect 11512 5650 11524 5684
rect 12112 5650 12190 5684
rect 12190 5650 12224 5684
rect 12224 5650 12304 5684
rect 12890 5650 12902 5684
rect 12902 5650 12936 5684
rect 12936 5650 12948 5684
rect 11466 5632 11524 5650
rect 12112 5639 12304 5650
rect 12178 5632 12236 5639
rect 12890 5632 12948 5650
rect 8958 5463 9016 5481
rect 10026 5463 10084 5481
rect 8958 5429 8970 5463
rect 8970 5429 9004 5463
rect 9004 5429 9016 5463
rect 10026 5429 10038 5463
rect 10038 5429 10072 5463
rect 10072 5429 10084 5463
rect 8958 5423 9016 5429
rect 10026 5423 10084 5429
rect 11644 5462 11702 5480
rect 12712 5462 12770 5480
rect 11644 5428 11656 5462
rect 11656 5428 11690 5462
rect 11690 5428 11702 5462
rect 12712 5428 12724 5462
rect 12724 5428 12758 5462
rect 12758 5428 12770 5462
rect 11644 5422 11702 5428
rect 12712 5422 12770 5428
rect 8780 4804 8838 4810
rect 10560 4804 10618 4810
rect 8780 4770 8792 4804
rect 8792 4770 8826 4804
rect 8826 4770 8838 4804
rect 10560 4770 10572 4804
rect 10572 4770 10606 4804
rect 10606 4770 10618 4804
rect 8780 4752 8838 4770
rect 10560 4752 10618 4770
rect 11110 4804 11168 4810
rect 12890 4804 12948 4810
rect 11110 4770 11122 4804
rect 11122 4770 11156 4804
rect 11156 4770 11168 4804
rect 12890 4770 12902 4804
rect 12902 4770 12936 4804
rect 12936 4770 12948 4804
rect 11110 4752 11168 4770
rect 12890 4752 12948 4770
rect 8958 4582 9016 4600
rect 9492 4597 9550 4600
rect 8958 4548 8970 4582
rect 8970 4548 9004 4582
rect 9004 4548 9016 4582
rect 8958 4542 9016 4548
rect 9430 4539 9622 4597
rect 10382 4582 10440 4600
rect 10382 4548 10394 4582
rect 10394 4548 10428 4582
rect 10428 4548 10440 4582
rect 10382 4542 10440 4548
rect 11288 4582 11346 4600
rect 12178 4596 12236 4600
rect 11288 4548 11300 4582
rect 11300 4548 11334 4582
rect 11334 4548 11346 4582
rect 11288 4542 11346 4548
rect 12109 4538 12301 4596
rect 12712 4582 12770 4600
rect 12712 4548 12724 4582
rect 12724 4548 12758 4582
rect 12758 4548 12770 4582
rect 12712 4542 12770 4548
rect 8780 4234 8838 4240
rect 9428 4234 9620 4241
rect 10560 4234 10618 4240
rect 8780 4200 8792 4234
rect 8792 4200 8826 4234
rect 8826 4200 8838 4234
rect 9428 4200 9504 4234
rect 9504 4200 9538 4234
rect 9538 4200 9620 4234
rect 10560 4200 10572 4234
rect 10572 4200 10606 4234
rect 10606 4200 10618 4234
rect 8780 4182 8838 4200
rect 9428 4183 9620 4200
rect 9490 4182 9548 4183
rect 10560 4182 10618 4200
rect 11110 4234 11168 4240
rect 12109 4234 12301 4242
rect 12890 4234 12948 4240
rect 11110 4200 11122 4234
rect 11122 4200 11156 4234
rect 11156 4200 11168 4234
rect 12109 4200 12190 4234
rect 12190 4200 12224 4234
rect 12224 4200 12301 4234
rect 12890 4200 12902 4234
rect 12902 4200 12936 4234
rect 12936 4200 12948 4234
rect 11110 4182 11168 4200
rect 12109 4184 12301 4200
rect 12178 4182 12236 4184
rect 12890 4182 12948 4200
rect 8958 4012 9016 4030
rect 10382 4012 10440 4030
rect 8958 3978 8970 4012
rect 8970 3978 9004 4012
rect 9004 3978 9016 4012
rect 10382 3978 10394 4012
rect 10394 3978 10428 4012
rect 10428 3978 10440 4012
rect 8958 3972 9016 3978
rect 10382 3972 10440 3978
rect 11288 4012 11346 4030
rect 12712 4012 12770 4030
rect 11288 3978 11300 4012
rect 11300 3978 11334 4012
rect 11334 3978 11346 4012
rect 12712 3978 12724 4012
rect 12724 3978 12758 4012
rect 12758 3978 12770 4012
rect 11288 3972 11346 3978
rect 12712 3972 12770 3978
rect 16359 3928 16417 3986
rect 18139 3928 18197 3986
rect 16733 3884 16898 3893
rect 16733 3850 16852 3884
rect 16852 3850 16886 3884
rect 16886 3850 16898 3884
rect 16733 3839 16898 3850
rect 17457 3884 17622 3892
rect 17457 3850 17572 3884
rect 17572 3850 17606 3884
rect 17606 3850 17622 3884
rect 17457 3838 17622 3850
rect 15876 3702 16142 3716
rect 15876 3668 15890 3702
rect 15890 3668 15924 3702
rect 15924 3668 16102 3702
rect 16102 3668 16136 3702
rect 16136 3668 16142 3702
rect 15876 3662 16142 3668
rect 18504 3702 18770 3714
rect 18504 3668 18518 3702
rect 18518 3668 18552 3702
rect 18552 3668 18730 3702
rect 18730 3668 18764 3702
rect 18764 3668 18770 3702
rect 18504 3660 18770 3668
rect 16359 3568 16417 3626
rect 18139 3568 18197 3626
rect 8422 3304 8480 3310
rect 9420 3304 9612 3311
rect 10558 3304 10616 3310
rect 8422 3270 8434 3304
rect 8434 3270 8468 3304
rect 8468 3270 8480 3304
rect 9420 3270 9502 3304
rect 9502 3270 9536 3304
rect 9536 3270 9612 3304
rect 10558 3270 10570 3304
rect 10570 3270 10604 3304
rect 10604 3270 10616 3304
rect 8422 3252 8480 3270
rect 9420 3253 9612 3270
rect 9490 3252 9548 3253
rect 10558 3252 10616 3270
rect 11109 3304 11167 3310
rect 12116 3304 12308 3310
rect 13245 3304 13303 3310
rect 11109 3270 11121 3304
rect 11121 3270 11155 3304
rect 11155 3270 11167 3304
rect 12116 3270 12189 3304
rect 12189 3270 12223 3304
rect 12223 3270 12308 3304
rect 13245 3270 13257 3304
rect 13257 3270 13291 3304
rect 13291 3270 13303 3304
rect 11109 3252 11167 3270
rect 12116 3252 12308 3270
rect 13245 3252 13303 3270
rect 8956 3082 9014 3100
rect 10024 3082 10082 3100
rect 8956 3048 8968 3082
rect 8968 3048 9002 3082
rect 9002 3048 9014 3082
rect 10024 3048 10036 3082
rect 10036 3048 10070 3082
rect 10070 3048 10082 3082
rect 8956 3042 9014 3048
rect 10024 3042 10082 3048
rect 11643 3082 11701 3100
rect 12711 3082 12769 3100
rect 11643 3048 11655 3082
rect 11655 3048 11689 3082
rect 11689 3048 11701 3082
rect 12711 3048 12723 3082
rect 12723 3048 12757 3082
rect 12757 3048 12769 3082
rect 14126 3104 14184 3110
rect 15550 3104 15608 3110
rect 14126 3070 14138 3104
rect 14138 3070 14172 3104
rect 14172 3070 14184 3104
rect 15550 3070 15562 3104
rect 15562 3070 15596 3104
rect 15596 3070 15608 3104
rect 14126 3052 14184 3070
rect 15550 3052 15608 3070
rect 15874 3104 16140 3113
rect 16974 3104 17032 3110
rect 15874 3070 15918 3104
rect 15918 3070 15952 3104
rect 15952 3070 16140 3104
rect 16974 3070 16986 3104
rect 16986 3070 17020 3104
rect 17020 3070 17032 3104
rect 15874 3059 16140 3070
rect 16974 3052 17032 3070
rect 17526 3104 17584 3110
rect 18504 3104 18770 3110
rect 17526 3070 17538 3104
rect 17538 3070 17572 3104
rect 17572 3070 17584 3104
rect 18504 3070 18606 3104
rect 18606 3070 18640 3104
rect 18640 3070 18770 3104
rect 17526 3052 17584 3070
rect 18504 3056 18770 3070
rect 18950 3104 19008 3110
rect 20374 3104 20432 3110
rect 18950 3070 18962 3104
rect 18962 3070 18996 3104
rect 18996 3070 19008 3104
rect 20374 3070 20386 3104
rect 20386 3070 20420 3104
rect 20420 3070 20432 3104
rect 18950 3052 19008 3070
rect 20374 3052 20432 3070
rect 11643 3042 11701 3048
rect 12711 3042 12769 3048
rect 15016 2882 15074 2900
rect 16084 2882 16142 2900
rect 15016 2848 15028 2882
rect 15028 2848 15062 2882
rect 15062 2848 15074 2882
rect 16084 2848 16096 2882
rect 16096 2848 16130 2882
rect 16130 2848 16142 2882
rect 15016 2842 15074 2848
rect 16084 2842 16142 2848
rect 18416 2882 18474 2900
rect 19484 2882 19542 2900
rect 18416 2848 18428 2882
rect 18428 2848 18462 2882
rect 18462 2848 18474 2882
rect 19484 2848 19496 2882
rect 19496 2848 19530 2882
rect 19530 2848 19542 2882
rect 18416 2842 18474 2848
rect 19484 2842 19542 2848
rect 8422 2804 8480 2810
rect 9490 2804 9548 2810
rect 10558 2804 10616 2810
rect 8422 2770 8434 2804
rect 8434 2770 8468 2804
rect 8468 2770 8480 2804
rect 9490 2770 9502 2804
rect 9502 2770 9536 2804
rect 9536 2770 9548 2804
rect 10558 2770 10570 2804
rect 10570 2770 10604 2804
rect 10604 2770 10616 2804
rect 8422 2752 8480 2770
rect 9490 2752 9548 2770
rect 10558 2752 10616 2770
rect 11109 2804 11167 2810
rect 12177 2804 12235 2810
rect 13245 2804 13303 2810
rect 11109 2770 11121 2804
rect 11121 2770 11155 2804
rect 11155 2770 11167 2804
rect 12177 2770 12189 2804
rect 12189 2770 12223 2804
rect 12223 2770 12235 2804
rect 13245 2770 13257 2804
rect 13257 2770 13291 2804
rect 13291 2770 13303 2804
rect 11109 2752 11167 2770
rect 12177 2752 12235 2770
rect 13245 2752 13303 2770
rect 8956 2582 9014 2600
rect 10024 2582 10082 2600
rect 8956 2548 8968 2582
rect 8968 2548 9002 2582
rect 9002 2548 9014 2582
rect 10024 2548 10036 2582
rect 10036 2548 10070 2582
rect 10070 2548 10082 2582
rect 8956 2542 9014 2548
rect 10024 2542 10082 2548
rect 11643 2582 11701 2600
rect 12711 2582 12769 2600
rect 11643 2548 11655 2582
rect 11655 2548 11689 2582
rect 11689 2548 11701 2582
rect 12711 2548 12723 2582
rect 12723 2548 12757 2582
rect 12757 2548 12769 2582
rect 14126 2604 14184 2610
rect 15550 2604 15608 2610
rect 16974 2604 17032 2610
rect 14126 2570 14138 2604
rect 14138 2570 14172 2604
rect 14172 2570 14184 2604
rect 15550 2570 15562 2604
rect 15562 2570 15596 2604
rect 15596 2570 15608 2604
rect 16974 2570 16986 2604
rect 16986 2570 17020 2604
rect 17020 2570 17032 2604
rect 14126 2552 14184 2570
rect 15550 2552 15608 2570
rect 16974 2552 17032 2570
rect 17526 2604 17584 2610
rect 18950 2604 19008 2610
rect 20374 2604 20432 2610
rect 17526 2570 17538 2604
rect 17538 2570 17572 2604
rect 17572 2570 17584 2604
rect 18950 2570 18962 2604
rect 18962 2570 18996 2604
rect 18996 2570 19008 2604
rect 20374 2570 20386 2604
rect 20386 2570 20420 2604
rect 20420 2570 20432 2604
rect 17526 2552 17584 2570
rect 18950 2552 19008 2570
rect 20374 2552 20432 2570
rect 11643 2542 11701 2548
rect 12711 2542 12769 2548
rect 15016 2382 15074 2401
rect 16084 2382 16142 2400
rect 15016 2348 15028 2382
rect 15028 2348 15062 2382
rect 15062 2348 15074 2382
rect 16084 2348 16096 2382
rect 16096 2348 16130 2382
rect 16130 2348 16142 2382
rect 15016 2343 15074 2348
rect 16084 2342 16142 2348
rect 18416 2382 18474 2400
rect 19484 2382 19542 2400
rect 18416 2348 18428 2382
rect 18428 2348 18462 2382
rect 18462 2348 18474 2382
rect 19484 2348 19496 2382
rect 19496 2348 19530 2382
rect 19530 2348 19542 2382
rect 18416 2342 18474 2348
rect 19484 2342 19542 2348
rect 8422 2304 8480 2310
rect 9490 2304 9548 2310
rect 10558 2304 10616 2310
rect 8422 2270 8434 2304
rect 8434 2270 8468 2304
rect 8468 2270 8480 2304
rect 9490 2270 9502 2304
rect 9502 2270 9536 2304
rect 9536 2270 9548 2304
rect 10558 2270 10570 2304
rect 10570 2270 10604 2304
rect 10604 2270 10616 2304
rect 8422 2252 8480 2270
rect 9490 2252 9548 2270
rect 10558 2252 10616 2270
rect 11109 2304 11167 2310
rect 12177 2304 12235 2310
rect 13245 2304 13303 2310
rect 11109 2270 11121 2304
rect 11121 2270 11155 2304
rect 11155 2270 11167 2304
rect 12177 2270 12189 2304
rect 12189 2270 12223 2304
rect 12223 2270 12235 2304
rect 13245 2270 13257 2304
rect 13257 2270 13291 2304
rect 13291 2270 13303 2304
rect 11109 2252 11167 2270
rect 12177 2252 12235 2270
rect 13245 2252 13303 2270
rect 8956 2082 9014 2100
rect 8956 2048 8968 2082
rect 8968 2048 9002 2082
rect 9002 2048 9014 2082
rect 8956 2042 9014 2048
rect 9274 2082 9480 2091
rect 10024 2082 10082 2100
rect 9274 2048 9324 2082
rect 9324 2048 9358 2082
rect 9358 2048 9480 2082
rect 10024 2048 10036 2082
rect 10036 2048 10070 2082
rect 10070 2048 10082 2082
rect 9274 2033 9480 2048
rect 10024 2042 10082 2048
rect 11643 2082 11701 2100
rect 12226 2082 12417 2091
rect 11643 2048 11655 2082
rect 11655 2048 11689 2082
rect 11689 2048 11701 2082
rect 12226 2048 12367 2082
rect 12367 2048 12401 2082
rect 12401 2048 12417 2082
rect 11643 2042 11701 2048
rect 12226 2038 12417 2048
rect 12711 2082 12769 2100
rect 12711 2048 12723 2082
rect 12723 2048 12757 2082
rect 12757 2048 12769 2082
rect 14126 2104 14184 2110
rect 15550 2104 15608 2110
rect 16974 2104 17032 2110
rect 14126 2070 14138 2104
rect 14138 2070 14172 2104
rect 14172 2070 14184 2104
rect 15550 2070 15562 2104
rect 15562 2070 15596 2104
rect 15596 2070 15608 2104
rect 16974 2070 16986 2104
rect 16986 2070 17020 2104
rect 17020 2070 17032 2104
rect 14126 2052 14184 2070
rect 15550 2052 15608 2070
rect 16974 2052 17032 2070
rect 17526 2104 17584 2110
rect 18950 2104 19008 2110
rect 20374 2104 20432 2110
rect 17526 2070 17538 2104
rect 17538 2070 17572 2104
rect 17572 2070 17584 2104
rect 18950 2070 18962 2104
rect 18962 2070 18996 2104
rect 18996 2070 19008 2104
rect 20374 2070 20386 2104
rect 20386 2070 20420 2104
rect 20420 2070 20432 2104
rect 17526 2052 17584 2070
rect 18950 2052 19008 2070
rect 20374 2052 20432 2070
rect 12711 2042 12769 2048
rect 15016 1882 15074 1900
rect 16084 1882 16142 1900
rect 15016 1848 15028 1882
rect 15028 1848 15062 1882
rect 15062 1848 15074 1882
rect 16084 1848 16096 1882
rect 16096 1848 16130 1882
rect 16130 1848 16142 1882
rect 15016 1842 15074 1848
rect 16084 1842 16142 1848
rect 18416 1882 18474 1900
rect 19484 1882 19542 1900
rect 18416 1848 18428 1882
rect 18428 1848 18462 1882
rect 18462 1848 18474 1882
rect 19484 1848 19496 1882
rect 19496 1848 19530 1882
rect 19530 1848 19542 1882
rect 18416 1842 18474 1848
rect 19484 1842 19542 1848
rect 9318 1610 9524 1611
rect 8422 1604 8480 1610
rect 9318 1604 9548 1610
rect 10558 1604 10616 1610
rect 8422 1570 8434 1604
rect 8434 1570 8468 1604
rect 8468 1570 8480 1604
rect 9318 1570 9502 1604
rect 9502 1570 9536 1604
rect 9536 1570 9548 1604
rect 10558 1570 10570 1604
rect 10570 1570 10604 1604
rect 10604 1570 10616 1604
rect 8422 1552 8480 1570
rect 9318 1552 9548 1570
rect 10558 1552 10616 1570
rect 11109 1604 11167 1610
rect 12169 1604 12433 1611
rect 13245 1604 13303 1610
rect 11109 1570 11121 1604
rect 11121 1570 11155 1604
rect 11155 1570 11167 1604
rect 12169 1570 12189 1604
rect 12189 1570 12223 1604
rect 12223 1570 12433 1604
rect 13245 1570 13257 1604
rect 13257 1570 13291 1604
rect 13291 1570 13303 1604
rect 11109 1552 11167 1570
rect 12169 1552 12433 1570
rect 13245 1552 13303 1570
rect 14126 1604 14184 1610
rect 15550 1604 15608 1610
rect 16974 1604 17032 1610
rect 14126 1570 14138 1604
rect 14138 1570 14172 1604
rect 14172 1570 14184 1604
rect 15550 1570 15562 1604
rect 15562 1570 15596 1604
rect 15596 1570 15608 1604
rect 16974 1570 16986 1604
rect 16986 1570 17020 1604
rect 17020 1570 17032 1604
rect 14126 1552 14184 1570
rect 15550 1552 15608 1570
rect 16974 1552 17032 1570
rect 17526 1604 17584 1610
rect 18950 1604 19008 1610
rect 20374 1604 20432 1610
rect 17526 1570 17538 1604
rect 17538 1570 17572 1604
rect 17572 1570 17584 1604
rect 18950 1570 18962 1604
rect 18962 1570 18996 1604
rect 18996 1570 19008 1604
rect 20374 1570 20386 1604
rect 20386 1570 20420 1604
rect 20420 1570 20432 1604
rect 17526 1552 17584 1570
rect 18950 1552 19008 1570
rect 20374 1552 20432 1570
rect 9318 1551 9524 1552
rect 8956 1382 9014 1400
rect 10024 1382 10082 1400
rect 8956 1348 8968 1382
rect 8968 1348 9002 1382
rect 9002 1348 9014 1382
rect 10024 1348 10036 1382
rect 10036 1348 10070 1382
rect 10070 1348 10082 1382
rect 8956 1342 9014 1348
rect 10024 1342 10082 1348
rect 11643 1382 11701 1400
rect 12711 1382 12769 1400
rect 11643 1348 11655 1382
rect 11655 1348 11689 1382
rect 11689 1348 11701 1382
rect 12711 1348 12723 1382
rect 12723 1348 12757 1382
rect 12757 1348 12769 1382
rect 11643 1342 11701 1348
rect 12711 1342 12769 1348
rect 15016 1382 15074 1400
rect 16084 1382 16142 1400
rect 15016 1348 15028 1382
rect 15028 1348 15062 1382
rect 15062 1348 15074 1382
rect 16084 1348 16096 1382
rect 16096 1348 16130 1382
rect 16130 1348 16142 1382
rect 15016 1342 15074 1348
rect 16084 1342 16142 1348
rect 18416 1382 18474 1400
rect 19484 1382 19542 1400
rect 18416 1348 18428 1382
rect 18428 1348 18462 1382
rect 18462 1348 18474 1382
rect 19484 1348 19496 1382
rect 19496 1348 19530 1382
rect 19530 1348 19542 1382
rect 18416 1342 18474 1348
rect 19484 1342 19542 1348
rect 8422 1104 8480 1110
rect 9490 1104 9548 1110
rect 10558 1104 10616 1110
rect 8422 1070 8434 1104
rect 8434 1070 8468 1104
rect 8468 1070 8480 1104
rect 9490 1070 9502 1104
rect 9502 1070 9536 1104
rect 9536 1070 9548 1104
rect 10558 1070 10570 1104
rect 10570 1070 10604 1104
rect 10604 1070 10616 1104
rect 8422 1052 8480 1070
rect 9490 1052 9548 1070
rect 10558 1052 10616 1070
rect 11109 1104 11167 1110
rect 12177 1104 12235 1110
rect 13245 1104 13303 1110
rect 11109 1070 11121 1104
rect 11121 1070 11155 1104
rect 11155 1070 11167 1104
rect 12177 1070 12189 1104
rect 12189 1070 12223 1104
rect 12223 1070 12235 1104
rect 13245 1070 13257 1104
rect 13257 1070 13291 1104
rect 13291 1070 13303 1104
rect 11109 1052 11167 1070
rect 12177 1052 12235 1070
rect 13245 1052 13303 1070
rect 14126 1104 14184 1110
rect 15550 1104 15608 1110
rect 16974 1104 17032 1110
rect 14126 1070 14138 1104
rect 14138 1070 14172 1104
rect 14172 1070 14184 1104
rect 15550 1070 15562 1104
rect 15562 1070 15596 1104
rect 15596 1070 15608 1104
rect 16974 1070 16986 1104
rect 16986 1070 17020 1104
rect 17020 1070 17032 1104
rect 14126 1052 14184 1070
rect 15550 1052 15608 1070
rect 16974 1052 17032 1070
rect 17526 1104 17584 1110
rect 18950 1104 19008 1110
rect 20374 1104 20432 1110
rect 17526 1070 17538 1104
rect 17538 1070 17572 1104
rect 17572 1070 17584 1104
rect 18950 1070 18962 1104
rect 18962 1070 18996 1104
rect 18996 1070 19008 1104
rect 20374 1070 20386 1104
rect 20386 1070 20420 1104
rect 20420 1070 20432 1104
rect 17526 1052 17584 1070
rect 18950 1052 19008 1070
rect 20374 1052 20432 1070
rect 8956 882 9014 900
rect 10024 882 10082 900
rect 8956 848 8968 882
rect 8968 848 9002 882
rect 9002 848 9014 882
rect 10024 848 10036 882
rect 10036 848 10070 882
rect 10070 848 10082 882
rect 8956 842 9014 848
rect 10024 842 10082 848
rect 11643 882 11701 900
rect 12711 882 12769 900
rect 11643 848 11655 882
rect 11655 848 11689 882
rect 11689 848 11701 882
rect 12711 848 12723 882
rect 12723 848 12757 882
rect 12757 848 12769 882
rect 11643 842 11701 848
rect 12711 842 12769 848
rect 15016 882 15074 900
rect 16084 882 16142 900
rect 15016 848 15028 882
rect 15028 848 15062 882
rect 15062 848 15074 882
rect 16084 848 16096 882
rect 16096 848 16130 882
rect 16130 848 16142 882
rect 15016 842 15074 848
rect 16084 842 16142 848
rect 18416 882 18474 900
rect 19484 882 19542 900
rect 18416 848 18428 882
rect 18428 848 18462 882
rect 18462 848 18474 882
rect 19484 848 19496 882
rect 19496 848 19530 882
rect 19530 848 19542 882
rect 18416 842 18474 848
rect 19484 842 19542 848
rect 8422 604 8480 610
rect 9490 604 9548 610
rect 10558 604 10616 610
rect 8422 570 8434 604
rect 8434 570 8468 604
rect 8468 570 8480 604
rect 9490 570 9502 604
rect 9502 570 9536 604
rect 9536 570 9548 604
rect 10558 570 10570 604
rect 10570 570 10604 604
rect 10604 570 10616 604
rect 8422 552 8480 570
rect 9490 552 9548 570
rect 10558 552 10616 570
rect 11109 604 11167 610
rect 12177 604 12235 610
rect 13245 604 13303 610
rect 11109 570 11121 604
rect 11121 570 11155 604
rect 11155 570 11167 604
rect 12177 570 12189 604
rect 12189 570 12223 604
rect 12223 570 12235 604
rect 13245 570 13257 604
rect 13257 570 13291 604
rect 13291 570 13303 604
rect 11109 552 11167 570
rect 12177 552 12235 570
rect 13245 552 13303 570
rect 14126 604 14184 610
rect 15550 604 15608 610
rect 16974 604 17032 610
rect 14126 570 14138 604
rect 14138 570 14172 604
rect 14172 570 14184 604
rect 15550 570 15562 604
rect 15562 570 15596 604
rect 15596 570 15608 604
rect 16974 570 16986 604
rect 16986 570 17020 604
rect 17020 570 17032 604
rect 14126 552 14184 570
rect 15550 552 15608 570
rect 16974 552 17032 570
rect 17526 604 17584 610
rect 18950 604 19008 610
rect 20374 604 20432 610
rect 17526 570 17538 604
rect 17538 570 17572 604
rect 17572 570 17584 604
rect 18950 570 18962 604
rect 18962 570 18996 604
rect 18996 570 19008 604
rect 20374 570 20386 604
rect 20386 570 20420 604
rect 20420 570 20432 604
rect 17526 552 17584 570
rect 18950 552 19008 570
rect 20374 552 20432 570
rect 8956 382 9014 400
rect 10024 382 10082 400
rect 8956 348 8968 382
rect 8968 348 9002 382
rect 9002 348 9014 382
rect 10024 348 10036 382
rect 10036 348 10070 382
rect 10070 348 10082 382
rect 8956 342 9014 348
rect 10024 342 10082 348
rect 11643 382 11701 400
rect 12711 382 12769 400
rect 11643 348 11655 382
rect 11655 348 11689 382
rect 11689 348 11701 382
rect 12711 348 12723 382
rect 12723 348 12757 382
rect 12757 348 12769 382
rect 11643 342 11701 348
rect 12711 342 12769 348
rect 15016 382 15074 400
rect 16084 382 16142 400
rect 15016 348 15028 382
rect 15028 348 15062 382
rect 15062 348 15074 382
rect 16084 348 16096 382
rect 16096 348 16130 382
rect 16130 348 16142 382
rect 15016 342 15074 348
rect 16084 342 16142 348
rect 18416 382 18474 400
rect 19484 382 19542 400
rect 18416 348 18428 382
rect 18428 348 18462 382
rect 18462 348 18474 382
rect 19484 348 19496 382
rect 19496 348 19530 382
rect 19530 348 19542 382
rect 18416 342 18474 348
rect 19484 342 19542 348
rect 8929 -264 9048 -213
rect 9990 -264 10116 -196
rect 11586 -264 11753 -206
rect 12671 -264 12809 -194
rect 14955 -264 15135 -196
rect 16018 -264 16208 -194
rect 18336 -264 18526 -196
rect 19417 -264 19607 -201
rect 8929 -310 9048 -264
rect 9990 -310 10116 -264
rect 11586 -313 11753 -264
rect 12671 -313 12809 -264
rect 14955 -312 15135 -264
rect 16018 -305 16208 -264
rect 18336 -307 18526 -264
rect 19417 -312 19607 -264
rect 11586 -322 11753 -313
rect 12671 -315 12809 -313
<< metal2 >>
rect 8958 6672 9016 6682
rect 8780 6269 8838 6279
rect 8501 5945 8580 5955
rect 8069 5893 8182 5903
rect 8182 5776 8501 5893
rect 8069 5766 8182 5776
rect 8501 5735 8580 5745
rect 8780 5691 8838 6211
rect 8780 5623 8838 5633
rect 8958 6058 9016 6614
rect 8958 5481 9016 6000
rect 10026 6667 10084 6677
rect 10026 6058 10084 6609
rect 11644 6670 11702 6680
rect 9426 5695 9618 5705
rect 9426 5633 9492 5637
rect 9550 5633 9618 5637
rect 9426 5627 9618 5633
rect 8958 5413 9016 5423
rect 9471 5010 9581 5627
rect 10026 5481 10084 6000
rect 10204 6262 10262 6272
rect 10204 5691 10262 6204
rect 11466 6268 11524 6278
rect 10471 5874 10529 5884
rect 11200 5874 11258 5884
rect 10529 5816 11200 5874
rect 10471 5806 10529 5816
rect 11200 5806 11258 5816
rect 10204 5623 10262 5633
rect 11466 5690 11524 6210
rect 11466 5622 11524 5632
rect 11644 6058 11702 6612
rect 10026 5413 10084 5423
rect 11644 5480 11702 6000
rect 12712 6667 12770 6677
rect 12712 6058 12770 6609
rect 12112 5697 12304 5707
rect 12112 5632 12178 5639
rect 12236 5632 12304 5639
rect 12112 5629 12304 5632
rect 11644 5412 11702 5422
rect 9553 4928 9581 5010
rect 8780 4810 8838 4820
rect 8780 4240 8838 4752
rect 8780 4172 8838 4182
rect 8958 4600 9016 4610
rect 9471 4607 9581 4928
rect 12151 5395 12261 5629
rect 12712 5480 12770 6000
rect 12890 6263 12948 6273
rect 12890 5690 12948 6205
rect 12890 5622 12948 5632
rect 12712 5412 12770 5422
rect 12151 5313 12155 5395
rect 12237 5313 12261 5395
rect 10560 4810 10618 4820
rect 8958 4030 9016 4542
rect 9430 4600 9622 4607
rect 9430 4597 9492 4600
rect 9550 4597 9622 4600
rect 9430 4529 9622 4539
rect 10382 4600 10440 4610
rect 9428 4241 9620 4251
rect 9428 4182 9490 4183
rect 9548 4182 9620 4183
rect 9428 4173 9620 4182
rect 8958 3962 9016 3972
rect 9466 3321 9576 4173
rect 10382 4120 10440 4542
rect 10560 4240 10618 4752
rect 10560 4172 10618 4182
rect 11110 4810 11168 4820
rect 11110 4240 11168 4752
rect 11288 4600 11346 4610
rect 12151 4606 12261 5313
rect 17477 5308 17486 5400
rect 17578 5308 17587 5400
rect 16768 5015 16860 5030
rect 12890 4810 12948 4820
rect 11288 4346 11346 4542
rect 12109 4600 12301 4606
rect 12109 4596 12178 4600
rect 12236 4596 12301 4600
rect 12109 4528 12301 4538
rect 12712 4600 12770 4610
rect 11274 4234 11366 4346
rect 12109 4242 12301 4252
rect 11110 4172 11168 4182
rect 10364 4030 10456 4120
rect 10364 4008 10382 4030
rect 10440 4008 10456 4030
rect 11288 4030 11346 4234
rect 12109 4182 12178 4184
rect 12236 4182 12301 4184
rect 12109 4174 12301 4182
rect 10382 3962 10440 3972
rect 11288 3962 11346 3972
rect 8422 3310 8480 3320
rect 8422 2810 8480 3252
rect 9420 3311 9612 3321
rect 12153 3320 12263 4174
rect 12712 4030 12770 4542
rect 12890 4240 12948 4752
rect 12890 4172 12948 4182
rect 12712 3962 12770 3972
rect 16359 3986 16417 3996
rect 15876 3716 16142 3726
rect 15876 3652 16142 3662
rect 9420 3252 9490 3253
rect 9548 3252 9612 3253
rect 9420 3243 9612 3252
rect 10558 3310 10616 3320
rect 8422 2310 8480 2752
rect 8422 2242 8480 2252
rect 8956 3100 9014 3110
rect 8956 2600 9014 3042
rect 8956 2100 9014 2542
rect 9490 2810 9548 3243
rect 9490 2310 9548 2752
rect 9490 2242 9548 2252
rect 10024 3100 10082 3110
rect 10024 2600 10082 3042
rect 9325 2101 9435 2104
rect 8956 2032 9014 2042
rect 9274 2091 9480 2101
rect 9274 2023 9480 2033
rect 10024 2100 10082 2542
rect 10558 2810 10616 3252
rect 10558 2310 10616 2752
rect 10558 2242 10616 2252
rect 11109 3310 11167 3320
rect 11109 2810 11167 3252
rect 12116 3310 12308 3320
rect 12116 3242 12308 3252
rect 13245 3310 13303 3320
rect 12177 3201 12236 3242
rect 11109 2310 11167 2752
rect 11109 2242 11167 2252
rect 11643 3100 11701 3110
rect 11643 2600 11701 3042
rect 10024 2032 10082 2042
rect 11643 2100 11701 2542
rect 12177 2810 12235 3201
rect 12177 2310 12235 2752
rect 12177 2242 12235 2252
rect 12711 3100 12769 3110
rect 12711 2600 12769 3042
rect 11643 2032 11701 2042
rect 12226 2091 12417 2101
rect 12226 2028 12417 2038
rect 12711 2100 12769 2542
rect 13245 2810 13303 3252
rect 15973 3123 16065 3652
rect 16359 3626 16417 3928
rect 16768 3903 16860 4923
rect 17486 4341 17578 5308
rect 17485 4229 17578 4341
rect 16733 3893 16898 3903
rect 17486 3902 17578 4229
rect 18139 3986 18197 3996
rect 16733 3829 16898 3839
rect 17457 3892 17622 3902
rect 17457 3828 17622 3838
rect 16359 3560 16417 3568
rect 18139 3626 18197 3928
rect 18504 3714 18770 3724
rect 18504 3650 18770 3660
rect 18139 3557 18197 3568
rect 13245 2310 13303 2752
rect 13245 2242 13303 2252
rect 14126 3110 14184 3120
rect 14126 2610 14184 3052
rect 15550 3110 15608 3120
rect 12711 2032 12769 2042
rect 14126 2110 14184 2552
rect 9325 1621 9435 2023
rect 12246 1621 12356 2028
rect 9318 1620 9526 1621
rect 8422 1610 8480 1620
rect 8422 1110 8480 1552
rect 9318 1611 9548 1620
rect 9524 1610 9548 1611
rect 9524 1551 9548 1552
rect 9318 1541 9548 1551
rect 8422 610 8480 1052
rect 8422 542 8480 552
rect 8956 1400 9014 1410
rect 8956 900 9014 1342
rect 8956 400 9014 842
rect 9490 1110 9548 1541
rect 10558 1610 10616 1620
rect 9490 610 9548 1052
rect 9490 542 9548 552
rect 10024 1400 10082 1410
rect 10024 900 10082 1342
rect 8956 -203 9014 342
rect 10024 400 10082 842
rect 10558 1110 10616 1552
rect 10558 610 10616 1052
rect 10558 542 10616 552
rect 11109 1610 11167 1620
rect 11109 1110 11167 1552
rect 12169 1611 12433 1621
rect 12169 1542 12433 1552
rect 13245 1610 13303 1620
rect 11109 610 11167 1052
rect 11109 542 11167 552
rect 11643 1400 11701 1410
rect 11643 900 11701 1342
rect 10024 -186 10082 342
rect 11643 400 11701 842
rect 12177 1110 12235 1542
rect 12177 610 12235 1052
rect 12177 542 12235 552
rect 12711 1400 12769 1410
rect 12711 900 12769 1342
rect 9990 -196 10116 -186
rect 11643 -196 11701 342
rect 12711 400 12769 842
rect 13245 1110 13303 1552
rect 13245 610 13303 1052
rect 13245 542 13303 552
rect 14126 1610 14184 2052
rect 14126 1110 14184 1552
rect 14126 610 14184 1052
rect 14126 542 14184 552
rect 15016 2900 15074 2910
rect 15016 2401 15074 2842
rect 15016 1900 15074 2343
rect 15016 1400 15074 1842
rect 15016 900 15074 1342
rect 12711 -184 12769 342
rect 15016 400 15074 842
rect 15550 2610 15608 3052
rect 15874 3113 16140 3123
rect 18596 3120 18688 3650
rect 15874 3049 16140 3059
rect 16974 3110 17032 3120
rect 15550 2110 15608 2552
rect 15550 1610 15608 2052
rect 15550 1110 15608 1552
rect 15550 610 15608 1052
rect 15550 542 15608 552
rect 16084 2900 16142 2910
rect 16084 2400 16142 2842
rect 16084 1900 16142 2342
rect 16084 1400 16142 1842
rect 16084 900 16142 1342
rect 12671 -194 12809 -184
rect 15016 -186 15074 342
rect 16084 400 16142 842
rect 16974 2610 17032 3052
rect 16974 2110 17032 2552
rect 16974 1610 17032 2052
rect 16974 1110 17032 1552
rect 16974 610 17032 1052
rect 16974 542 17032 552
rect 17526 3110 17584 3120
rect 17526 2610 17584 3052
rect 18504 3110 18770 3120
rect 18504 3046 18770 3056
rect 18950 3110 19008 3120
rect 17526 2110 17584 2552
rect 17526 1610 17584 2052
rect 17526 1110 17584 1552
rect 17526 610 17584 1052
rect 17526 542 17584 552
rect 18416 2900 18474 2910
rect 18416 2400 18474 2842
rect 18416 1900 18474 2342
rect 18416 1400 18474 1842
rect 18416 900 18474 1342
rect 16084 -184 16142 342
rect 18416 400 18474 842
rect 18950 2610 19008 3052
rect 20374 3110 20432 3120
rect 18950 2110 19008 2552
rect 18950 1610 19008 2052
rect 18950 1110 19008 1552
rect 18950 610 19008 1052
rect 18950 542 19008 552
rect 19484 2900 19542 2910
rect 19484 2400 19542 2842
rect 19484 1900 19542 2342
rect 19484 1400 19542 1842
rect 19484 900 19542 1342
rect 8929 -213 9048 -203
rect 8929 -320 9048 -310
rect 9990 -320 10116 -310
rect 11586 -206 11753 -196
rect 11586 -332 11753 -322
rect 12671 -325 12809 -315
rect 14955 -196 15135 -186
rect 14955 -322 15135 -312
rect 16018 -194 16208 -184
rect 18416 -186 18474 342
rect 19484 400 19542 842
rect 20374 2610 20432 3052
rect 20374 2110 20432 2552
rect 20374 1610 20432 2052
rect 20374 1110 20432 1552
rect 20374 610 20432 1052
rect 20374 542 20432 552
rect 16018 -315 16208 -305
rect 18336 -196 18526 -186
rect 19484 -191 19542 342
rect 18336 -317 18526 -307
rect 19417 -201 19607 -191
rect 19417 -322 19607 -312
<< via2 >>
rect 9471 4928 9553 5010
rect 12155 5313 12237 5395
rect 17486 5308 17578 5400
rect 16768 4923 16860 5015
<< metal3 >>
rect 17481 5400 17583 5405
rect 12150 5395 17486 5400
rect 12150 5313 12155 5395
rect 12237 5313 17486 5395
rect 12150 5308 17486 5313
rect 17578 5308 17583 5400
rect 17481 5303 17583 5308
rect 16763 5015 16865 5020
rect 9466 5010 16768 5015
rect 9466 4928 9471 5010
rect 9553 4928 16768 5010
rect 9466 4923 16768 4928
rect 16860 4923 16865 5015
rect 16763 4918 16865 4923
use bias_circuit  bias_circuit_0
timestamp 1654674269
transform 1 0 -615 0 1 276
box -430 -610 8656 6437
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_0
timestamp 1654674269
transform 1 0 9519 0 1 476
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_1
timestamp 1654674269
transform 1 0 9519 0 1 976
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_2
timestamp 1654674269
transform 1 0 9519 0 1 1476
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_3
timestamp 1654674269
transform 1 0 12206 0 1 1476
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_4
timestamp 1654674269
transform 1 0 12206 0 1 976
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_5
timestamp 1654674269
transform 1 0 12206 0 1 476
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_6
timestamp 1654674269
transform 1 0 9519 0 1 2176
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_7
timestamp 1654674269
transform 1 0 9519 0 1 2676
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_8
timestamp 1654674269
transform 1 0 9519 0 1 3176
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_9
timestamp 1654674269
transform 1 0 12206 0 1 3176
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_10
timestamp 1654674269
transform 1 0 12206 0 1 2676
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_AKSJZW  sky130_fd_pr__nfet_01v8_AKSJZW_11
timestamp 1654674269
transform 1 0 12206 0 1 2176
box -1275 -228 1275 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_0
timestamp 1654674269
transform 1 0 15579 0 1 2476
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_1
timestamp 1654674269
transform 1 0 18979 0 1 476
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_2
timestamp 1654674269
transform 1 0 18979 0 1 976
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_3
timestamp 1654674269
transform 1 0 18979 0 1 1476
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_4
timestamp 1654674269
transform 1 0 18979 0 1 1976
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_5
timestamp 1654674269
transform 1 0 18979 0 1 2476
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_6
timestamp 1654674269
transform 1 0 18979 0 1 2976
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_7
timestamp 1654674269
transform 1 0 15579 0 1 2976
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_8
timestamp 1654674269
transform 1 0 15579 0 1 1976
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_9
timestamp 1654674269
transform 1 0 15579 0 1 1476
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_10
timestamp 1654674269
transform 1 0 15579 0 1 976
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_S6RQQZ  sky130_fd_pr__nfet_01v8_S6RQQZ_11
timestamp 1654674269
transform 1 0 15579 0 1 476
box -1631 -228 1631 228
use sky130_fd_pr__nfet_01v8_lvt_K7HVMB  sky130_fd_pr__nfet_01v8_lvt_K7HVMB_0
timestamp 1654674269
transform 1 0 16388 0 1 3776
box -820 -208 820 208
use sky130_fd_pr__nfet_01v8_lvt_K7HVMB  sky130_fd_pr__nfet_01v8_lvt_K7HVMB_1
timestamp 1654674269
transform 1 0 18168 0 1 3776
box -820 -208 820 208
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_0
timestamp 1654674269
transform 1 0 9699 0 1 4106
box -1133 -241 1133 241
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_1
timestamp 1654674269
transform 1 0 9699 0 1 4676
box -1133 -241 1133 241
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_2
timestamp 1654674269
transform 1 0 12029 0 1 4676
box -1133 -241 1133 241
use sky130_fd_pr__pfet_01v8_YVTMSC  sky130_fd_pr__pfet_01v8_YVTMSC_3
timestamp 1654674269
transform 1 0 12029 0 1 4106
box -1133 -241 1133 241
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_0
timestamp 1654674269
transform 1 0 9521 0 1 5557
box -1311 -241 1311 241
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_1
timestamp 1654674269
transform 1 0 12207 0 1 5556
box -1311 -241 1311 241
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_2
timestamp 1654674269
transform 1 0 9521 0 1 6134
box -1311 -241 1311 241
use sky130_fd_pr__pfet_01v8_lvt_YVTR7C  sky130_fd_pr__pfet_01v8_lvt_YVTR7C_3
timestamp 1654674269
transform 1 0 12207 0 1 6134
box -1311 -241 1311 241
<< labels >>
flabel metal1 20312 3383 20312 3383 1 FreeSans 800 0 0 0 cmc
flabel metal1 16275 4764 16275 4764 1 FreeSans 800 0 0 0 ip
flabel metal1 18061 4759 18061 4759 1 FreeSans 800 0 0 0 in
flabel metal1 6138 2598 6138 2598 1 FreeSans 800 0 0 0 bias_e
flabel metal1 -539 773 -539 773 1 FreeSans 800 0 0 0 i_bias
flabel metal1 -1030 -255 -1030 -255 1 FreeSans 800 0 0 0 VSS
flabel metal1 -842 6648 -842 6648 1 FreeSans 800 0 0 0 VDD
flabel metal1 15652 13 15652 13 1 FreeSans 800 0 0 0 bias_a
flabel metal2 9517 3665 9517 3665 1 FreeSans 800 0 0 0 on
flabel metal2 12208 3672 12208 3672 1 FreeSans 800 0 0 0 op
<< end >>
