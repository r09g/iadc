* NGSPICE file created from esd_cell.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_BRTJC6 a_n345_n500# a_1135_n588# a_n603_n588#
+ a_n1393_n588# a_n1609_n500# a_661_n588# a_n1135_n500# a_n977_n500# a_1293_n588#
+ a_n761_n588# a_n503_n500# a_n1551_n588# a_129_n500# a_n1293_n500# a_287_n500# a_n661_n500#
+ a_1451_n588# a_n1451_n500# a_919_n500# a_445_n500# a_1077_n500# a_29_n588# a_n129_n588#
+ a_603_n500# a_187_n588# a_1235_n500# a_n287_n588# a_761_n500# a_819_n588# a_345_n588#
+ a_n1077_n588# a_n29_n500# a_1393_n500# a_n919_n588# a_n1743_n722# a_n187_n500# a_977_n588#
+ a_n445_n588# a_503_n588# a_n1235_n588# a_1551_n500# a_n819_n500#
X0 a_n819_n500# a_n919_n588# a_n977_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n588# a_n819_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n588# a_761_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n588# a_n345_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n588# a_603_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n588# a_129_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n588# a_n1451_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n588# a_1235_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n588# a_n503_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n588# a_n29_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n588# a_287_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n588# a_n1609_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n588# a_1393_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n588# a_n1135_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_n503_n500# a_n603_n588# a_n661_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_1077_n500# a_977_n588# a_919_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n588# a_n187_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n588# a_445_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n588# a_n1293_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n588# a_1077_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_287_n500# a_n187_n500# 0.15fF
C1 a_n345_n500# a_129_n500# 0.15fF
C2 a_n187_n500# a_445_n500# 0.11fF
C3 a_n187_n500# a_129_n500# 0.24fF
C4 a_761_n500# a_n503_n500# 0.05fF
C5 a_n503_n500# a_603_n500# 0.06fF
C6 a_919_n500# a_n503_n500# 0.05fF
C7 a_287_n500# a_n503_n500# 0.09fF
C8 a_603_n500# a_n661_n500# 0.05fF
C9 a_445_n500# a_n503_n500# 0.07fF
C10 a_761_n500# a_n661_n500# 0.05fF
C11 a_919_n500# a_n661_n500# 0.04fF
C12 a_129_n500# a_n503_n500# 0.11fF
C13 a_287_n500# a_n661_n500# 0.07fF
C14 a_445_n500# a_n661_n500# 0.06fF
C15 a_n819_n500# a_603_n500# 0.05fF
C16 a_761_n500# a_n819_n500# 0.04fF
C17 a_129_n500# a_n661_n500# 0.09fF
C18 a_287_n500# a_n819_n500# 0.06fF
C19 a_445_n500# a_n819_n500# 0.05fF
C20 a_129_n500# a_n819_n500# 0.07fF
C21 a_n29_n500# a_n345_n500# 0.24fF
C22 a_n29_n500# a_n187_n500# 0.56fF
C23 a_603_n500# a_n977_n500# 0.04fF
C24 a_n345_n500# a_n187_n500# 0.56fF
C25 a_445_n500# a_n1135_n500# 0.04fF
C26 a_287_n500# a_n1135_n500# 0.05fF
C27 a_445_n500# a_n977_n500# 0.05fF
C28 a_287_n500# a_n977_n500# 0.05fF
C29 a_n1135_n500# a_129_n500# 0.05fF
C30 a_129_n500# a_n977_n500# 0.06fF
C31 a_287_n500# a_n1293_n500# 0.04fF
C32 a_n29_n500# a_n503_n500# 0.15fF
C33 a_n345_n500# a_n503_n500# 0.56fF
C34 a_129_n500# a_n1293_n500# 0.05fF
C35 a_n1451_n500# a_129_n500# 0.04fF
C36 a_n187_n500# a_n503_n500# 0.24fF
C37 a_n29_n500# a_n661_n500# 0.11fF
C38 a_n345_n500# a_n661_n500# 0.24fF
C39 a_n187_n500# a_n661_n500# 0.15fF
C40 a_n29_n500# a_n819_n500# 0.09fF
C41 a_n345_n500# a_n819_n500# 0.15fF
C42 a_n187_n500# a_n819_n500# 0.11fF
C43 a_n503_n500# a_n661_n500# 0.56fF
C44 a_n29_n500# a_n1135_n500# 0.06fF
C45 a_n29_n500# a_n977_n500# 0.07fF
C46 a_n345_n500# a_n1135_n500# 0.09fF
C47 a_n345_n500# a_n977_n500# 0.11fF
C48 a_n503_n500# a_n819_n500# 0.24fF
C49 a_n187_n500# a_n1135_n500# 0.07fF
C50 a_n187_n500# a_n977_n500# 0.09fF
C51 a_n29_n500# a_n1293_n500# 0.05fF
C52 a_n29_n500# a_n1451_n500# 0.05fF
C53 a_n345_n500# a_n1293_n500# 0.07fF
C54 a_n29_n500# a_n1609_n500# 0.04fF
C55 a_n345_n500# a_n1451_n500# 0.06fF
C56 a_n819_n500# a_n661_n500# 0.56fF
C57 a_n187_n500# a_n1293_n500# 0.06fF
C58 a_n345_n500# a_n1609_n500# 0.05fF
C59 a_n187_n500# a_n1451_n500# 0.05fF
C60 a_n187_n500# a_n1609_n500# 0.05fF
C61 a_n1135_n500# a_n503_n500# 0.11fF
C62 a_n503_n500# a_n977_n500# 0.15fF
C63 a_n503_n500# a_n1293_n500# 0.09fF
C64 a_n1135_n500# a_n661_n500# 0.15fF
C65 a_n977_n500# a_n661_n500# 0.24fF
C66 a_n1451_n500# a_n503_n500# 0.07fF
C67 a_n503_n500# a_n1609_n500# 0.06fF
C68 a_n1293_n500# a_n661_n500# 0.11fF
C69 a_n1451_n500# a_n661_n500# 0.09fF
C70 a_n1135_n500# a_n819_n500# 0.24fF
C71 a_n819_n500# a_n977_n500# 0.56fF
C72 a_n661_n500# a_n1609_n500# 0.07fF
C73 a_n819_n500# a_n1293_n500# 0.15fF
C74 a_n1451_n500# a_n819_n500# 0.11fF
C75 a_n819_n500# a_n1609_n500# 0.09fF
C76 a_n1135_n500# a_n977_n500# 0.56fF
C77 a_n1135_n500# a_n1293_n500# 0.56fF
C78 a_n977_n500# a_n1293_n500# 0.24fF
C79 a_n1451_n500# a_n1135_n500# 0.24fF
C80 a_n1451_n500# a_n977_n500# 0.15fF
C81 a_n1135_n500# a_n1609_n500# 0.15fF
C82 a_n977_n500# a_n1609_n500# 0.11fF
C83 a_n1451_n500# a_n1293_n500# 0.56fF
C84 a_n1293_n500# a_n1609_n500# 0.24fF
C85 a_n1451_n500# a_n1609_n500# 0.56fF
C86 a_1451_n588# a_1135_n588# 0.04fF
C87 a_1293_n588# a_1135_n588# 0.12fF
C88 a_1293_n588# a_1451_n588# 0.12fF
C89 a_977_n588# a_1135_n588# 0.12fF
C90 a_977_n588# a_1451_n588# 0.02fF
C91 a_1293_n588# a_977_n588# 0.04fF
C92 a_819_n588# a_1135_n588# 0.04fF
C93 a_1451_n588# a_819_n588# 0.02fF
C94 a_1293_n588# a_819_n588# 0.02fF
C95 a_977_n588# a_819_n588# 0.12fF
C96 a_1451_n588# a_661_n588# 0.01fF
C97 a_661_n588# a_1135_n588# 0.02fF
C98 a_1293_n588# a_661_n588# 0.02fF
C99 a_977_n588# a_661_n588# 0.04fF
C100 a_187_n588# a_1135_n588# 0.01fF
C101 a_1451_n588# a_187_n588# 0.01fF
C102 a_1293_n588# a_187_n588# 0.01fF
C103 a_1451_n588# a_345_n588# 0.01fF
C104 a_345_n588# a_1135_n588# 0.01fF
C105 a_661_n588# a_819_n588# 0.12fF
C106 a_977_n588# a_187_n588# 0.01fF
C107 a_1293_n588# a_345_n588# 0.01fF
C108 a_503_n588# a_1135_n588# 0.02fF
C109 a_1451_n588# a_503_n588# 0.01fF
C110 a_977_n588# a_345_n588# 0.02fF
C111 a_1293_n588# a_503_n588# 0.01fF
C112 a_187_n588# a_819_n588# 0.02fF
C113 a_977_n588# a_503_n588# 0.02fF
C114 a_345_n588# a_819_n588# 0.02fF
C115 a_503_n588# a_819_n588# 0.04fF
C116 a_29_n588# a_1135_n588# 0.01fF
C117 a_1451_n588# a_29_n588# 0.01fF
C118 a_1293_n588# a_29_n588# 0.01fF
C119 a_187_n588# a_661_n588# 0.02fF
C120 a_345_n588# a_661_n588# 0.04fF
C121 a_977_n588# a_29_n588# 0.01fF
C122 a_503_n588# a_661_n588# 0.12fF
C123 a_29_n588# a_819_n588# 0.01fF
C124 a_345_n588# a_187_n588# 0.12fF
C125 a_503_n588# a_187_n588# 0.04fF
C126 a_345_n588# a_503_n588# 0.12fF
C127 a_n129_n588# a_1135_n588# 0.01fF
C128 a_1451_n588# a_n129_n588# 0.01fF
C129 a_1293_n588# a_n129_n588# 0.01fF
C130 a_977_n588# a_n129_n588# 0.01fF
C131 a_n287_n588# a_1135_n588# 0.01fF
C132 a_n445_n588# a_1135_n588# 0.01fF
C133 a_1293_n588# a_n287_n588# 0.01fF
C134 a_29_n588# a_661_n588# 0.02fF
C135 a_977_n588# a_n287_n588# 0.01fF
C136 a_n445_n588# a_977_n588# 0.01fF
C137 a_n129_n588# a_819_n588# 0.01fF
C138 a_187_n588# a_29_n588# 0.12fF
C139 a_n287_n588# a_819_n588# 0.01fF
C140 a_345_n588# a_29_n588# 0.04fF
C141 a_n445_n588# a_819_n588# 0.01fF
C142 a_503_n588# a_29_n588# 0.02fF
C143 a_977_n588# a_n603_n588# 0.01fF
C144 a_n129_n588# a_661_n588# 0.01fF
C145 a_819_n588# a_n603_n588# 0.01fF
C146 a_n761_n588# a_819_n588# 0.01fF
C147 a_n287_n588# a_661_n588# 0.01fF
C148 a_n129_n588# a_187_n588# 0.04fF
C149 a_n445_n588# a_661_n588# 0.01fF
C150 a_345_n588# a_n129_n588# 0.02fF
C151 a_187_n588# a_n287_n588# 0.02fF
C152 a_n445_n588# a_187_n588# 0.02fF
C153 a_503_n588# a_n129_n588# 0.02fF
C154 a_345_n588# a_n287_n588# 0.02fF
C155 a_n445_n588# a_345_n588# 0.01fF
C156 a_661_n588# a_n919_n588# 0.01fF
C157 a_503_n588# a_n287_n588# 0.01fF
C158 a_n761_n588# a_661_n588# 0.01fF
C159 a_661_n588# a_n603_n588# 0.01fF
C160 a_n445_n588# a_503_n588# 0.01fF
C161 a_187_n588# a_n919_n588# 0.01fF
C162 a_187_n588# a_n603_n588# 0.01fF
C163 a_n761_n588# a_187_n588# 0.01fF
C164 a_345_n588# a_n919_n588# 0.01fF
C165 a_n761_n588# a_345_n588# 0.01fF
C166 a_345_n588# a_n603_n588# 0.01fF
C167 a_503_n588# a_n919_n588# 0.01fF
C168 a_187_n588# a_n1077_n588# 0.01fF
C169 a_n129_n588# a_29_n588# 0.12fF
C170 a_503_n588# a_n603_n588# 0.01fF
C171 a_345_n588# a_n1077_n588# 0.01fF
C172 a_n761_n588# a_503_n588# 0.01fF
C173 a_29_n588# a_n287_n588# 0.04fF
C174 a_n445_n588# a_29_n588# 0.02fF
C175 a_503_n588# a_n1077_n588# 0.01fF
C176 a_n1235_n588# a_187_n588# 0.01fF
C177 a_29_n588# a_n919_n588# 0.01fF
C178 a_n1235_n588# a_345_n588# 0.01fF
C179 a_29_n588# a_n603_n588# 0.02fF
C180 a_n761_n588# a_29_n588# 0.01fF
C181 a_n1393_n588# a_187_n588# 0.01fF
C182 a_29_n588# a_n1077_n588# 0.01fF
C183 a_n129_n588# a_n287_n588# 0.12fF
C184 a_n445_n588# a_n129_n588# 0.04fF
C185 a_n445_n588# a_n287_n588# 0.12fF
C186 a_n129_n588# a_n919_n588# 0.01fF
C187 a_n129_n588# a_n603_n588# 0.02fF
C188 a_n1235_n588# a_29_n588# 0.01fF
C189 a_n761_n588# a_n129_n588# 0.02fF
C190 a_n287_n588# a_n919_n588# 0.02fF
C191 a_n129_n588# a_n1077_n588# 0.01fF
C192 a_n445_n588# a_n919_n588# 0.02fF
C193 a_n287_n588# a_n603_n588# 0.04fF
C194 a_n761_n588# a_n287_n588# 0.02fF
C195 a_n445_n588# a_n603_n588# 0.12fF
C196 a_n445_n588# a_n761_n588# 0.04fF
C197 a_n1393_n588# a_29_n588# 0.01fF
C198 a_n287_n588# a_n1077_n588# 0.01fF
C199 a_n445_n588# a_n1077_n588# 0.02fF
C200 a_n603_n588# a_n919_n588# 0.04fF
C201 a_n761_n588# a_n919_n588# 0.12fF
C202 a_n761_n588# a_n603_n588# 0.12fF
C203 a_29_n588# a_n1551_n588# 0.01fF
C204 a_n1235_n588# a_n129_n588# 0.01fF
C205 a_n919_n588# a_n1077_n588# 0.12fF
C206 a_n761_n588# a_n1077_n588# 0.04fF
C207 a_n603_n588# a_n1077_n588# 0.02fF
C208 a_n1235_n588# a_n287_n588# 0.01fF
C209 a_n445_n588# a_n1235_n588# 0.01fF
C210 a_n1393_n588# a_n129_n588# 0.01fF
C211 a_n1393_n588# a_n287_n588# 0.01fF
C212 a_n445_n588# a_n1393_n588# 0.01fF
C213 a_n1235_n588# a_n919_n588# 0.04fF
C214 a_n1235_n588# a_n603_n588# 0.02fF
C215 a_n129_n588# a_n1551_n588# 0.01fF
C216 a_n761_n588# a_n1235_n588# 0.02fF
C217 a_n1235_n588# a_n1077_n588# 0.12fF
C218 a_n287_n588# a_n1551_n588# 0.01fF
C219 a_n445_n588# a_n1551_n588# 0.01fF
C220 a_n1393_n588# a_n919_n588# 0.02fF
C221 a_n1393_n588# a_n603_n588# 0.01fF
C222 a_n761_n588# a_n1393_n588# 0.02fF
C223 a_n1393_n588# a_n1077_n588# 0.04fF
C224 a_n919_n588# a_n1551_n588# 0.02fF
C225 a_n761_n588# a_n1551_n588# 0.01fF
C226 a_n603_n588# a_n1551_n588# 0.01fF
C227 a_n1077_n588# a_n1551_n588# 0.02fF
C228 a_n1393_n588# a_n1235_n588# 0.12fF
C229 a_n1235_n588# a_n1551_n588# 0.04fF
C230 a_n1393_n588# a_n1551_n588# 0.12fF
C231 a_1551_n500# a_1393_n500# 0.56fF
C232 a_1551_n500# a_1077_n500# 0.15fF
C233 a_1077_n500# a_1393_n500# 0.24fF
C234 a_1235_n500# a_1393_n500# 0.56fF
C235 a_1551_n500# a_1235_n500# 0.24fF
C236 a_1551_n500# a_603_n500# 0.07fF
C237 a_761_n500# a_1551_n500# 0.09fF
C238 a_603_n500# a_1393_n500# 0.09fF
C239 a_919_n500# a_1551_n500# 0.11fF
C240 a_761_n500# a_1393_n500# 0.11fF
C241 a_919_n500# a_1393_n500# 0.15fF
C242 a_1077_n500# a_1235_n500# 0.56fF
C243 a_445_n500# a_1551_n500# 0.06fF
C244 a_287_n500# a_1393_n500# 0.06fF
C245 a_287_n500# a_1551_n500# 0.05fF
C246 a_445_n500# a_1393_n500# 0.07fF
C247 a_1551_n500# a_129_n500# 0.05fF
C248 a_129_n500# a_1393_n500# 0.05fF
C249 a_1077_n500# a_603_n500# 0.15fF
C250 a_919_n500# a_1077_n500# 0.56fF
C251 a_761_n500# a_1077_n500# 0.24fF
C252 a_761_n500# a_1235_n500# 0.15fF
C253 a_1235_n500# a_603_n500# 0.11fF
C254 a_919_n500# a_1235_n500# 0.24fF
C255 a_287_n500# a_1077_n500# 0.09fF
C256 a_445_n500# a_1077_n500# 0.11fF
C257 a_1077_n500# a_129_n500# 0.07fF
C258 a_445_n500# a_1235_n500# 0.09fF
C259 a_287_n500# a_1235_n500# 0.07fF
C260 a_1235_n500# a_129_n500# 0.06fF
C261 a_761_n500# a_603_n500# 0.56fF
C262 a_919_n500# a_603_n500# 0.24fF
C263 a_919_n500# a_761_n500# 0.56fF
C264 a_287_n500# a_761_n500# 0.15fF
C265 a_287_n500# a_603_n500# 0.24fF
C266 a_761_n500# a_445_n500# 0.24fF
C267 a_445_n500# a_603_n500# 0.56fF
C268 a_287_n500# a_919_n500# 0.11fF
C269 a_919_n500# a_445_n500# 0.15fF
C270 a_761_n500# a_129_n500# 0.11fF
C271 a_129_n500# a_603_n500# 0.15fF
C272 a_919_n500# a_129_n500# 0.09fF
C273 a_n29_n500# a_1551_n500# 0.04fF
C274 a_n29_n500# a_1393_n500# 0.05fF
C275 a_287_n500# a_445_n500# 0.56fF
C276 a_287_n500# a_129_n500# 0.56fF
C277 a_445_n500# a_129_n500# 0.24fF
C278 a_n187_n500# a_1393_n500# 0.04fF
C279 a_n29_n500# a_1077_n500# 0.06fF
C280 a_n345_n500# a_1077_n500# 0.05fF
C281 a_n29_n500# a_1235_n500# 0.05fF
C282 a_n187_n500# a_1077_n500# 0.05fF
C283 a_n345_n500# a_1235_n500# 0.04fF
C284 a_n187_n500# a_1235_n500# 0.05fF
C285 a_n29_n500# a_603_n500# 0.11fF
C286 a_n29_n500# a_761_n500# 0.09fF
C287 a_n29_n500# a_919_n500# 0.07fF
C288 a_n345_n500# a_761_n500# 0.06fF
C289 a_n345_n500# a_603_n500# 0.07fF
C290 a_n345_n500# a_919_n500# 0.05fF
C291 a_1077_n500# a_n503_n500# 0.04fF
C292 a_n187_n500# a_603_n500# 0.09fF
C293 a_761_n500# a_n187_n500# 0.07fF
C294 a_919_n500# a_n187_n500# 0.06fF
C295 a_n29_n500# a_287_n500# 0.24fF
C296 a_n29_n500# a_445_n500# 0.15fF
C297 a_n345_n500# a_287_n500# 0.11fF
C298 a_n29_n500# a_129_n500# 0.56fF
C299 a_n345_n500# a_445_n500# 0.09fF
C300 a_1551_n500# a_n1743_n722# 0.30fF
C301 a_1393_n500# a_n1743_n722# 0.13fF
C302 a_1235_n500# a_n1743_n722# 0.09fF
C303 a_1077_n500# a_n1743_n722# 0.07fF
C304 a_919_n500# a_n1743_n722# 0.06fF
C305 a_761_n500# a_n1743_n722# 0.05fF
C306 a_603_n500# a_n1743_n722# 0.05fF
C307 a_445_n500# a_n1743_n722# 0.04fF
C308 a_287_n500# a_n1743_n722# 0.04fF
C309 a_129_n500# a_n1743_n722# 0.04fF
C310 a_n29_n500# a_n1743_n722# 0.02fF
C311 a_n187_n500# a_n1743_n722# 0.04fF
C312 a_n345_n500# a_n1743_n722# 0.04fF
C313 a_n503_n500# a_n1743_n722# 0.04fF
C314 a_n661_n500# a_n1743_n722# 0.05fF
C315 a_n819_n500# a_n1743_n722# 0.05fF
C316 a_n977_n500# a_n1743_n722# 0.06fF
C317 a_n1135_n500# a_n1743_n722# 0.07fF
C318 a_n1293_n500# a_n1743_n722# 0.09fF
C319 a_n1451_n500# a_n1743_n722# 0.13fF
C320 a_n1609_n500# a_n1743_n722# 0.30fF
C321 a_1451_n588# a_n1743_n722# 0.28fF
C322 a_1293_n588# a_n1743_n722# 0.23fF
C323 a_1135_n588# a_n1743_n722# 0.24fF
C324 a_977_n588# a_n1743_n722# 0.25fF
C325 a_819_n588# a_n1743_n722# 0.26fF
C326 a_661_n588# a_n1743_n722# 0.26fF
C327 a_503_n588# a_n1743_n722# 0.27fF
C328 a_345_n588# a_n1743_n722# 0.28fF
C329 a_187_n588# a_n1743_n722# 0.28fF
C330 a_29_n588# a_n1743_n722# 0.28fF
C331 a_n129_n588# a_n1743_n722# 0.28fF
C332 a_n287_n588# a_n1743_n722# 0.28fF
C333 a_n445_n588# a_n1743_n722# 0.28fF
C334 a_n603_n588# a_n1743_n722# 0.28fF
C335 a_n761_n588# a_n1743_n722# 0.28fF
C336 a_n919_n588# a_n1743_n722# 0.28fF
C337 a_n1077_n588# a_n1743_n722# 0.28fF
C338 a_n1235_n588# a_n1743_n722# 0.29fF
C339 a_n1393_n588# a_n1743_n722# 0.29fF
C340 a_n1551_n588# a_n1743_n722# 0.34fF
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CADZ46 a_n345_n500# a_n1609_n500# a_n1135_n500#
+ a_29_n597# a_n977_n500# a_n129_n597# a_187_n597# a_n503_n500# a_129_n500# a_n1293_n500#
+ a_n287_n597# a_819_n597# a_n1077_n597# a_287_n500# a_n661_n500# a_345_n597# a_n919_n597#
+ a_n1451_n500# a_977_n597# a_n445_n597# a_919_n500# a_n1235_n597# a_445_n500# a_503_n597#
+ w_n1809_n797# a_n603_n597# a_1077_n500# a_1135_n597# a_661_n597# a_n1393_n597# a_603_n500#
+ a_1293_n597# a_n761_n597# a_1235_n500# a_n1551_n597# a_761_n500# a_n29_n500# a_1451_n597#
+ a_1393_n500# a_n187_n500# a_1551_n500# a_n819_n500# VSUBS
X0 a_n819_n500# a_n919_n597# a_n977_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n597# a_n819_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n597# a_761_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n597# a_n345_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n597# a_603_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n597# a_129_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n597# a_n1451_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n597# a_1235_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n597# a_n503_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n597# a_n29_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n597# a_287_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n597# a_n1609_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n597# a_1393_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n597# a_n1135_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_1077_n500# a_977_n597# a_919_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X15 a_n503_n500# a_n603_n597# a_n661_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n597# a_n187_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n597# a_445_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n597# a_n1293_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n597# a_1077_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_n603_n597# a_n129_n597# 0.02fF
C1 a_29_n597# a_n445_n597# 0.02fF
C2 a_n129_n597# a_n761_n597# 0.02fF
C3 a_n129_n597# a_n445_n597# 0.04fF
C4 a_819_n597# w_n1809_n797# 0.21fF
C5 a_661_n597# w_n1809_n797# 0.22fF
C6 a_n1077_n597# a_187_n597# 0.01fF
C7 a_187_n597# a_n919_n597# 0.01fF
C8 a_n1235_n597# a_187_n597# 0.01fF
C9 a_977_n597# w_n1809_n797# 0.20fF
C10 a_n603_n597# a_187_n597# 0.01fF
C11 a_n919_n597# a_345_n597# 0.01fF
C12 a_1135_n597# w_n1809_n797# 0.20fF
C13 a_n761_n597# a_187_n597# 0.01fF
C14 a_n1077_n597# a_345_n597# 0.01fF
C15 a_n1235_n597# a_345_n597# 0.01fF
C16 w_n1809_n797# a_1293_n597# 0.19fF
C17 a_n445_n597# a_187_n597# 0.02fF
C18 a_n603_n597# a_345_n597# 0.01fF
C19 a_n761_n597# a_345_n597# 0.01fF
C20 a_n1077_n597# a_503_n597# 0.01fF
C21 a_503_n597# a_n919_n597# 0.01fF
C22 a_n445_n597# a_345_n597# 0.01fF
C23 a_n603_n597# a_503_n597# 0.01fF
C24 a_n761_n597# a_503_n597# 0.01fF
C25 a_1451_n597# w_n1809_n797# 0.24fF
C26 a_n1451_n500# w_n1809_n797# 0.13fF
C27 a_n1609_n500# w_n1809_n797# 0.30fF
C28 a_n445_n597# a_503_n597# 0.01fF
C29 a_n287_n597# a_29_n597# 0.04fF
C30 a_n1293_n500# w_n1809_n797# 0.09fF
C31 a_n287_n597# a_n129_n597# 0.12fF
C32 a_n1135_n500# w_n1809_n797# 0.07fF
C33 a_n919_n597# a_661_n597# 0.01fF
C34 a_29_n597# a_n129_n597# 0.12fF
C35 a_n761_n597# a_819_n597# 0.01fF
C36 a_n603_n597# a_819_n597# 0.01fF
C37 a_n761_n597# a_661_n597# 0.01fF
C38 a_n603_n597# a_661_n597# 0.01fF
C39 a_819_n597# a_n445_n597# 0.01fF
C40 a_n977_n500# w_n1809_n797# 0.06fF
C41 a_n445_n597# a_661_n597# 0.01fF
C42 a_n603_n597# a_977_n597# 0.01fF
C43 a_n287_n597# a_187_n597# 0.02fF
C44 a_n503_n500# w_n1809_n797# 0.04fF
C45 a_29_n597# a_187_n597# 0.12fF
C46 a_n445_n597# a_977_n597# 0.01fF
C47 a_n661_n500# w_n1809_n797# 0.05fF
C48 a_1135_n597# a_n445_n597# 0.01fF
C49 a_n129_n597# a_187_n597# 0.04fF
C50 a_n819_n500# w_n1809_n797# 0.05fF
C51 a_n287_n597# a_345_n597# 0.02fF
C52 a_29_n597# a_345_n597# 0.04fF
C53 a_n129_n597# a_345_n597# 0.02fF
C54 a_n287_n597# a_503_n597# 0.01fF
C55 a_1551_n500# a_n29_n500# 0.04fF
C56 a_n345_n500# w_n1809_n797# 0.04fF
C57 a_129_n500# a_1551_n500# 0.05fF
C58 a_29_n597# a_503_n597# 0.02fF
C59 a_n129_n597# a_503_n597# 0.02fF
C60 a_1551_n500# a_603_n500# 0.07fF
C61 a_445_n500# a_1551_n500# 0.06fF
C62 a_n187_n500# a_1393_n500# 0.04fF
C63 a_1551_n500# a_287_n500# 0.05fF
C64 a_187_n597# a_345_n597# 0.12fF
C65 a_1551_n500# a_761_n500# 0.09fF
C66 a_n29_n500# a_1393_n500# 0.05fF
C67 a_129_n500# a_1393_n500# 0.05fF
C68 a_n187_n500# w_n1809_n797# 0.04fF
C69 a_n287_n597# a_819_n597# 0.01fF
C70 a_n287_n597# a_661_n597# 0.01fF
C71 a_n29_n500# w_n1809_n797# 0.02fF
C72 a_29_n597# a_819_n597# 0.01fF
C73 a_129_n500# w_n1809_n797# 0.04fF
C74 a_29_n597# a_661_n597# 0.02fF
C75 a_187_n597# a_503_n597# 0.04fF
C76 a_n129_n597# a_819_n597# 0.01fF
C77 a_n129_n597# a_661_n597# 0.01fF
C78 a_n287_n597# a_977_n597# 0.01fF
C79 a_603_n500# a_1393_n500# 0.09fF
C80 a_287_n500# a_1393_n500# 0.06fF
C81 a_445_n500# a_1393_n500# 0.07fF
C82 a_919_n500# a_1551_n500# 0.11fF
C83 a_n287_n597# a_1135_n597# 0.01fF
C84 a_29_n597# a_977_n597# 0.01fF
C85 a_603_n500# w_n1809_n797# 0.05fF
C86 a_761_n500# a_1393_n500# 0.11fF
C87 a_n287_n597# a_1293_n597# 0.01fF
C88 a_29_n597# a_1135_n597# 0.01fF
C89 a_445_n500# w_n1809_n797# 0.04fF
C90 a_287_n500# w_n1809_n797# 0.04fF
C91 a_n129_n597# a_977_n597# 0.01fF
C92 a_503_n597# a_345_n597# 0.12fF
C93 a_29_n597# a_1293_n597# 0.01fF
C94 a_1077_n500# a_1551_n500# 0.15fF
C95 a_n129_n597# a_1135_n597# 0.01fF
C96 a_761_n500# w_n1809_n797# 0.05fF
C97 a_n129_n597# a_1293_n597# 0.01fF
C98 a_819_n597# a_187_n597# 0.02fF
C99 a_187_n597# a_661_n597# 0.02fF
C100 a_919_n500# a_1393_n500# 0.15fF
C101 a_1551_n500# a_1235_n500# 0.24fF
C102 a_919_n500# w_n1809_n797# 0.06fF
C103 a_187_n597# a_977_n597# 0.01fF
C104 a_1077_n500# a_1393_n500# 0.24fF
C105 a_819_n597# a_345_n597# 0.02fF
C106 a_29_n597# a_1451_n597# 0.01fF
C107 a_661_n597# a_345_n597# 0.04fF
C108 a_1135_n597# a_187_n597# 0.01fF
C109 a_187_n597# a_1293_n597# 0.01fF
C110 a_1077_n500# w_n1809_n797# 0.07fF
C111 a_1451_n597# a_n129_n597# 0.01fF
C112 a_1235_n500# a_1393_n500# 0.56fF
C113 a_977_n597# a_345_n597# 0.02fF
C114 a_1135_n597# a_345_n597# 0.01fF
C115 a_819_n597# a_503_n597# 0.04fF
C116 a_503_n597# a_661_n597# 0.12fF
C117 a_1235_n500# w_n1809_n797# 0.09fF
C118 a_345_n597# a_1293_n597# 0.01fF
C119 a_503_n597# a_977_n597# 0.02fF
C120 a_1135_n597# a_503_n597# 0.02fF
C121 a_1451_n597# a_187_n597# 0.01fF
C122 a_503_n597# a_1293_n597# 0.01fF
C123 a_819_n597# a_661_n597# 0.12fF
C124 a_1451_n597# a_345_n597# 0.01fF
C125 a_819_n597# a_977_n597# 0.12fF
C126 a_661_n597# a_977_n597# 0.04fF
C127 a_1135_n597# a_819_n597# 0.04fF
C128 a_1135_n597# a_661_n597# 0.02fF
C129 a_819_n597# a_1293_n597# 0.02fF
C130 a_1451_n597# a_503_n597# 0.01fF
C131 a_661_n597# a_1293_n597# 0.02fF
C132 a_1135_n597# a_977_n597# 0.12fF
C133 a_977_n597# a_1293_n597# 0.04fF
C134 a_1135_n597# a_1293_n597# 0.12fF
C135 a_1451_n597# a_819_n597# 0.02fF
C136 a_1451_n597# a_661_n597# 0.01fF
C137 a_1451_n597# a_977_n597# 0.02fF
C138 a_1451_n597# a_1135_n597# 0.04fF
C139 a_1451_n597# a_1293_n597# 0.12fF
C140 a_n1609_n500# a_n1451_n500# 0.56fF
C141 a_n1293_n500# a_n1451_n500# 0.56fF
C142 a_n1609_n500# a_n1293_n500# 0.24fF
C143 a_n1135_n500# a_n1451_n500# 0.24fF
C144 a_n1609_n500# a_n1135_n500# 0.15fF
C145 a_n1293_n500# a_n1135_n500# 0.56fF
C146 a_n977_n500# a_n1451_n500# 0.15fF
C147 a_n1609_n500# a_n977_n500# 0.11fF
C148 a_n1293_n500# a_n977_n500# 0.24fF
C149 a_n503_n500# a_n1451_n500# 0.07fF
C150 a_n1609_n500# a_n503_n500# 0.06fF
C151 a_n661_n500# a_n1451_n500# 0.09fF
C152 a_n977_n500# a_n1135_n500# 0.56fF
C153 a_n1609_n500# a_n661_n500# 0.07fF
C154 a_n1293_n500# a_n503_n500# 0.09fF
C155 a_n819_n500# a_n1451_n500# 0.11fF
C156 a_n1293_n500# a_n661_n500# 0.11fF
C157 a_n1609_n500# a_n819_n500# 0.09fF
C158 a_n1293_n500# a_n819_n500# 0.15fF
C159 a_n503_n500# a_n1135_n500# 0.11fF
C160 a_n661_n500# a_n1135_n500# 0.15fF
C161 a_n819_n500# a_n1135_n500# 0.24fF
C162 a_n345_n500# a_n1451_n500# 0.06fF
C163 a_n1609_n500# a_n345_n500# 0.05fF
C164 a_n503_n500# a_n977_n500# 0.15fF
C165 a_n1293_n500# a_n345_n500# 0.07fF
C166 a_n661_n500# a_n977_n500# 0.24fF
C167 a_n819_n500# a_n977_n500# 0.56fF
C168 a_n345_n500# a_n1135_n500# 0.09fF
C169 a_n661_n500# a_n503_n500# 0.56fF
C170 a_n819_n500# a_n503_n500# 0.24fF
C171 a_n661_n500# a_n819_n500# 0.56fF
C172 a_n187_n500# a_n1451_n500# 0.05fF
C173 a_n1609_n500# a_n187_n500# 0.05fF
C174 a_n1293_n500# a_n187_n500# 0.06fF
C175 a_n29_n500# a_n1451_n500# 0.05fF
C176 a_129_n500# a_n1451_n500# 0.04fF
C177 a_n1609_n500# a_n29_n500# 0.04fF
C178 a_n345_n500# a_n977_n500# 0.11fF
C179 a_n1293_n500# a_n29_n500# 0.05fF
C180 a_n187_n500# a_n1135_n500# 0.07fF
C181 a_129_n500# a_n1293_n500# 0.05fF
C182 a_n503_n500# a_n345_n500# 0.56fF
C183 a_n29_n500# a_n1135_n500# 0.06fF
C184 a_n661_n500# a_n345_n500# 0.24fF
C185 a_129_n500# a_n1135_n500# 0.05fF
C186 a_n819_n500# a_n345_n500# 0.15fF
C187 a_n1293_n500# a_287_n500# 0.04fF
C188 a_n187_n500# a_n977_n500# 0.09fF
C189 a_445_n500# a_n1135_n500# 0.04fF
C190 a_n1135_n500# a_287_n500# 0.05fF
C191 a_n29_n500# a_n977_n500# 0.07fF
C192 a_129_n500# a_n977_n500# 0.06fF
C193 a_n187_n500# a_n503_n500# 0.24fF
C194 a_n661_n500# a_n187_n500# 0.15fF
C195 a_n503_n500# a_n29_n500# 0.15fF
C196 a_129_n500# a_n503_n500# 0.11fF
C197 a_n819_n500# a_n187_n500# 0.11fF
C198 a_n661_n500# a_n29_n500# 0.11fF
C199 a_n977_n500# a_603_n500# 0.04fF
C200 a_129_n500# a_n661_n500# 0.09fF
C201 a_n819_n500# a_n29_n500# 0.09fF
C202 a_n977_n500# a_287_n500# 0.05fF
C203 a_445_n500# a_n977_n500# 0.05fF
C204 a_129_n500# a_n819_n500# 0.07fF
C205 a_n503_n500# a_603_n500# 0.06fF
C206 a_445_n500# a_n503_n500# 0.07fF
C207 a_n503_n500# a_287_n500# 0.09fF
C208 a_n661_n500# a_603_n500# 0.05fF
C209 a_445_n500# a_n661_n500# 0.06fF
C210 a_n661_n500# a_287_n500# 0.07fF
C211 a_n503_n500# a_761_n500# 0.05fF
C212 a_n819_n500# a_603_n500# 0.05fF
C213 a_n187_n500# a_n345_n500# 0.56fF
C214 a_n819_n500# a_287_n500# 0.06fF
C215 a_n661_n500# a_761_n500# 0.05fF
C216 a_445_n500# a_n819_n500# 0.05fF
C217 a_n345_n500# a_n29_n500# 0.24fF
C218 a_n819_n500# a_761_n500# 0.04fF
C219 a_129_n500# a_n345_n500# 0.15fF
C220 a_919_n500# a_n503_n500# 0.05fF
C221 a_n345_n500# a_603_n500# 0.07fF
C222 a_919_n500# a_n661_n500# 0.04fF
C223 a_445_n500# a_n345_n500# 0.09fF
C224 a_n345_n500# a_287_n500# 0.11fF
C225 a_n345_n500# a_761_n500# 0.06fF
C226 a_1077_n500# a_n503_n500# 0.04fF
C227 a_n187_n500# a_n29_n500# 0.56fF
C228 a_129_n500# a_n187_n500# 0.24fF
C229 a_129_n500# a_n29_n500# 0.56fF
C230 a_n187_n500# a_603_n500# 0.09fF
C231 a_n187_n500# a_287_n500# 0.15fF
C232 a_445_n500# a_n187_n500# 0.11fF
C233 a_919_n500# a_n345_n500# 0.05fF
C234 a_n29_n500# a_603_n500# 0.11fF
C235 a_129_n500# a_603_n500# 0.15fF
C236 a_n187_n500# a_761_n500# 0.07fF
C237 a_445_n500# a_n29_n500# 0.15fF
C238 a_n29_n500# a_287_n500# 0.24fF
C239 a_129_n500# a_287_n500# 0.56fF
C240 a_129_n500# a_445_n500# 0.24fF
C241 a_n29_n500# a_761_n500# 0.09fF
C242 a_1077_n500# a_n345_n500# 0.05fF
C243 a_129_n500# a_761_n500# 0.11fF
C244 a_445_n500# a_603_n500# 0.56fF
C245 a_287_n500# a_603_n500# 0.24fF
C246 a_n345_n500# a_1235_n500# 0.04fF
C247 a_445_n500# a_287_n500# 0.56fF
C248 a_919_n500# a_n187_n500# 0.06fF
C249 a_603_n500# a_761_n500# 0.56fF
C250 a_287_n500# a_761_n500# 0.15fF
C251 a_445_n500# a_761_n500# 0.24fF
C252 a_919_n500# a_n29_n500# 0.07fF
C253 a_129_n500# a_919_n500# 0.09fF
C254 a_1077_n500# a_n187_n500# 0.05fF
C255 a_1077_n500# a_n29_n500# 0.06fF
C256 a_129_n500# a_1077_n500# 0.07fF
C257 a_919_n500# a_603_n500# 0.24fF
C258 a_n187_n500# a_1235_n500# 0.05fF
C259 a_445_n500# a_919_n500# 0.15fF
C260 a_919_n500# a_287_n500# 0.11fF
C261 a_919_n500# a_761_n500# 0.56fF
C262 a_n29_n500# a_1235_n500# 0.05fF
C263 a_1077_n500# a_603_n500# 0.15fF
C264 a_129_n500# a_1235_n500# 0.06fF
C265 a_445_n500# a_1077_n500# 0.11fF
C266 a_1077_n500# a_287_n500# 0.09fF
C267 a_1077_n500# a_761_n500# 0.24fF
C268 a_603_n500# a_1235_n500# 0.11fF
C269 a_445_n500# a_1235_n500# 0.09fF
C270 a_287_n500# a_1235_n500# 0.07fF
C271 a_761_n500# a_1235_n500# 0.15fF
C272 a_1077_n500# a_919_n500# 0.56fF
C273 a_919_n500# a_1235_n500# 0.24fF
C274 a_1077_n500# a_1235_n500# 0.56fF
C275 a_1551_n500# a_1393_n500# 0.56fF
C276 a_1551_n500# w_n1809_n797# 0.30fF
C277 w_n1809_n797# a_1393_n500# 0.13fF
C278 a_n1393_n597# w_n1809_n797# 0.25fF
C279 a_n1551_n597# w_n1809_n797# 0.30fF
C280 a_n1077_n597# w_n1809_n797# 0.24fF
C281 a_n919_n597# w_n1809_n797# 0.24fF
C282 a_n1235_n597# w_n1809_n797# 0.24fF
C283 a_n1393_n597# a_n1551_n597# 0.12fF
C284 a_n603_n597# w_n1809_n797# 0.24fF
C285 a_n761_n597# w_n1809_n797# 0.24fF
C286 a_n445_n597# w_n1809_n797# 0.24fF
C287 a_n1393_n597# a_n919_n597# 0.02fF
C288 a_n1235_n597# a_n1393_n597# 0.12fF
C289 a_n1077_n597# a_n1393_n597# 0.04fF
C290 a_n1077_n597# a_n1551_n597# 0.02fF
C291 a_n1551_n597# a_n919_n597# 0.02fF
C292 a_n1235_n597# a_n1551_n597# 0.04fF
C293 a_n603_n597# a_n1393_n597# 0.01fF
C294 a_n761_n597# a_n1393_n597# 0.02fF
C295 a_n1393_n597# a_n445_n597# 0.01fF
C296 a_n603_n597# a_n1551_n597# 0.01fF
C297 a_n761_n597# a_n1551_n597# 0.01fF
C298 a_n1551_n597# a_n445_n597# 0.01fF
C299 a_n1077_n597# a_n919_n597# 0.12fF
C300 a_n1235_n597# a_n919_n597# 0.04fF
C301 a_n1235_n597# a_n1077_n597# 0.12fF
C302 a_n603_n597# a_n1077_n597# 0.02fF
C303 a_n603_n597# a_n919_n597# 0.04fF
C304 a_n1077_n597# a_n761_n597# 0.04fF
C305 a_n761_n597# a_n919_n597# 0.12fF
C306 a_n603_n597# a_n1235_n597# 0.02fF
C307 a_n1235_n597# a_n761_n597# 0.02fF
C308 a_n1077_n597# a_n445_n597# 0.02fF
C309 a_n445_n597# a_n919_n597# 0.02fF
C310 a_n1235_n597# a_n445_n597# 0.01fF
C311 a_n287_n597# w_n1809_n797# 0.24fF
C312 a_n603_n597# a_n761_n597# 0.12fF
C313 a_29_n597# w_n1809_n797# 0.24fF
C314 a_n603_n597# a_n445_n597# 0.12fF
C315 a_n761_n597# a_n445_n597# 0.04fF
C316 a_n129_n597# w_n1809_n797# 0.24fF
C317 a_n287_n597# a_n1393_n597# 0.01fF
C318 a_29_n597# a_n1393_n597# 0.01fF
C319 a_187_n597# w_n1809_n797# 0.24fF
C320 a_n287_n597# a_n1551_n597# 0.01fF
C321 a_n129_n597# a_n1393_n597# 0.01fF
C322 a_29_n597# a_n1551_n597# 0.01fF
C323 a_n129_n597# a_n1551_n597# 0.01fF
C324 w_n1809_n797# a_345_n597# 0.23fF
C325 a_n287_n597# a_n919_n597# 0.02fF
C326 a_n287_n597# a_n1077_n597# 0.01fF
C327 a_n287_n597# a_n1235_n597# 0.01fF
C328 a_29_n597# a_n1077_n597# 0.01fF
C329 a_29_n597# a_n919_n597# 0.01fF
C330 a_503_n597# w_n1809_n797# 0.23fF
C331 a_n1393_n597# a_187_n597# 0.01fF
C332 a_29_n597# a_n1235_n597# 0.01fF
C333 a_n129_n597# a_n919_n597# 0.01fF
C334 a_n1077_n597# a_n129_n597# 0.01fF
C335 a_n1235_n597# a_n129_n597# 0.01fF
C336 a_n287_n597# a_n603_n597# 0.04fF
C337 a_n287_n597# a_n761_n597# 0.02fF
C338 a_29_n597# a_n603_n597# 0.02fF
C339 a_29_n597# a_n761_n597# 0.01fF
C340 a_n287_n597# a_n445_n597# 0.12fF
C341 w_n1809_n797# VSUBS 17.30fF
.ends

.subckt esd_cell esd VDD VSS
Xsky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0 VSS VSS VSS VSS VSS VSS esd VSS VSS VSS esd
+ VSS esd VSS VSS VSS VSS esd VSS esd esd VSS VSS VSS VSS VSS VSS esd VSS VSS VSS
+ VSS esd VSS VSS esd VSS VSS VSS VSS VSS esd sky130_fd_pr__nfet_g5v0d10v5_BRTJC6
Xsky130_fd_pr__pfet_g5v0d10v5_CADZ46_0 VDD VDD esd VDD VDD VDD VDD esd esd VDD VDD
+ VDD VDD VDD VDD VDD VDD esd VDD VDD VDD VDD esd VDD VDD VDD esd VDD VDD VDD VDD
+ VDD VDD VDD VDD esd VDD VDD esd esd VDD esd VSS sky130_fd_pr__pfet_g5v0d10v5_CADZ46
C0 esd VDD 7.39fF
C1 VDD VSS -181.47fF
C2 esd VSS 8.04fF
.ends

