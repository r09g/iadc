magic
tech sky130A
magscale 1 2
timestamp 1654572275
<< nwell >>
rect 1089 2796 1135 2842
rect 1405 2796 1451 2842
rect 1721 2796 1767 2842
rect 2037 2796 2083 2842
rect 2353 2796 2399 2842
rect 2669 2796 2715 2842
rect 2985 2796 3031 2842
rect 3301 2796 3347 2842
rect 141 1711 187 1814
rect 3301 1757 3347 1798
rect 3140 1501 3192 1544
<< pwell >>
rect 3140 1440 3192 1451
rect 3301 1189 3347 1234
rect 141 115 187 205
rect 457 115 503 205
rect 773 115 819 205
rect 1089 115 1135 205
rect 1405 115 1451 205
rect 1721 115 1767 205
rect 2037 115 2083 205
rect 2353 115 2399 205
rect 2669 115 2715 205
rect 2985 115 3031 205
rect 3301 158 3347 204
<< mvndiff >>
rect 141 193 187 205
rect 457 193 503 205
rect 773 193 819 205
rect 1089 193 1135 205
rect 1405 193 1451 205
rect 1721 193 1767 205
rect 2037 193 2083 205
rect 2353 193 2399 205
rect 2669 193 2715 205
rect 2985 193 3031 205
<< mvpdiff >>
rect 1089 2796 1135 2798
rect 1405 2796 1451 2798
rect 1721 2796 1767 2798
rect 2037 2796 2083 2798
rect 2353 2796 2399 2798
rect 2669 2796 2715 2798
rect 2985 2796 3031 2798
rect 3301 2796 3347 2798
<< locali >>
rect 1095 2796 1129 2802
rect 1411 2796 1445 2802
rect 1727 2796 1761 2802
rect 2043 2796 2077 2802
rect 2359 2796 2393 2802
rect 2675 2796 2709 2802
rect 2991 2796 3025 2802
rect 3307 2796 3341 2802
rect 147 189 181 205
rect 463 189 497 205
rect 779 189 813 205
rect 1095 189 1129 205
rect 1411 189 1445 205
rect 1727 189 1761 205
rect 2043 189 2077 205
rect 2359 189 2393 205
rect 2675 189 2709 205
rect 2991 189 3025 205
<< viali >>
rect 109 2983 3379 3017
rect 13 1675 47 2921
rect 3441 1675 3475 2921
rect 13 79 47 1307
rect 3441 79 3475 1307
rect 109 -17 3379 17
<< metal1 >>
rect 7 3017 3481 3023
rect 7 2983 109 3017
rect 3379 2983 3481 3017
rect 7 2921 3481 2983
rect 7 1675 13 2921
rect 47 2839 3441 2921
rect 47 1757 59 2839
rect 141 2789 187 2839
rect 457 2795 503 2839
rect 773 2796 819 2839
rect 1089 2796 1135 2839
rect 1405 2796 1451 2839
rect 1721 2796 1767 2839
rect 2037 2796 2083 2839
rect 2353 2796 2399 2839
rect 2669 2796 2715 2839
rect 2985 2796 3031 2839
rect 3301 2796 3347 2839
rect 141 1757 187 1814
rect 286 1810 296 2786
rect 348 1810 358 2786
rect 602 1810 612 2786
rect 664 1810 674 2786
rect 918 1810 928 2786
rect 980 1810 990 2786
rect 1234 1810 1244 2786
rect 1296 1810 1306 2786
rect 1550 1810 1560 2786
rect 1612 1810 1622 2786
rect 1866 1810 1876 2786
rect 1928 1810 1938 2786
rect 2182 1810 2192 2786
rect 2244 1810 2254 2786
rect 2498 1810 2508 2786
rect 2560 1810 2570 2786
rect 2814 1810 2824 2786
rect 2876 1810 2886 2786
rect 3130 1810 3140 2786
rect 3192 1810 3202 2786
rect 3301 1757 3347 1798
rect 3429 1757 3441 2839
rect 47 1711 3441 1757
rect 47 1675 53 1711
rect 7 1663 53 1675
rect 3435 1675 3441 1711
rect 3475 1675 3481 2921
rect 3435 1663 3481 1675
rect -65 1544 3553 1555
rect -65 1440 296 1544
rect 348 1440 612 1544
rect 664 1440 928 1544
rect 980 1440 1244 1544
rect 1296 1440 1560 1544
rect 1612 1440 1876 1544
rect 1928 1440 2192 1544
rect 2244 1440 2508 1544
rect 2560 1440 2824 1544
rect 2876 1440 3140 1544
rect 3192 1440 3553 1544
rect -65 1427 3553 1440
rect 7 1307 53 1319
rect 7 79 13 1307
rect 47 1271 53 1307
rect 3435 1307 3481 1319
rect 3435 1271 3441 1307
rect 47 1225 3441 1271
rect 47 161 53 1225
rect 3301 1189 3347 1225
rect 286 205 296 1181
rect 348 205 358 1181
rect 602 205 612 1181
rect 664 205 674 1181
rect 918 205 928 1181
rect 980 205 990 1181
rect 1234 205 1244 1181
rect 1296 205 1306 1181
rect 1550 205 1560 1181
rect 1612 205 1622 1181
rect 1866 205 1876 1181
rect 1928 205 1938 1181
rect 2182 205 2192 1181
rect 2244 205 2254 1181
rect 2498 205 2508 1181
rect 2560 205 2570 1181
rect 2814 205 2824 1181
rect 2876 205 2886 1181
rect 3130 205 3140 1181
rect 3192 205 3202 1181
rect 141 161 187 205
rect 457 161 503 205
rect 773 161 819 205
rect 1089 161 1135 205
rect 1405 161 1451 205
rect 1721 161 1767 205
rect 2037 161 2083 205
rect 2353 161 2399 205
rect 2669 161 2715 205
rect 2985 161 3031 205
rect 3301 161 3347 204
rect 3435 161 3441 1225
rect 47 79 3441 161
rect 3475 79 3481 1307
rect 7 17 3481 79
rect 7 -17 109 17
rect 3379 -17 3481 17
rect 7 -23 3481 -17
<< via1 >>
rect 296 1810 348 2786
rect 612 1810 664 2786
rect 928 1810 980 2786
rect 1244 1810 1296 2786
rect 1560 1810 1612 2786
rect 1876 1810 1928 2786
rect 2192 1810 2244 2786
rect 2508 1810 2560 2786
rect 2824 1810 2876 2786
rect 3140 1810 3192 2786
rect 296 1440 348 1544
rect 612 1440 664 1544
rect 928 1440 980 1544
rect 1244 1440 1296 1544
rect 1560 1440 1612 1544
rect 1876 1440 1928 1544
rect 2192 1440 2244 1544
rect 2508 1440 2560 1544
rect 2824 1440 2876 1544
rect 3140 1440 3192 1544
rect 296 205 348 1181
rect 612 205 664 1181
rect 928 205 980 1181
rect 1244 205 1296 1181
rect 1560 205 1612 1181
rect 1876 205 1928 1181
rect 2192 205 2244 1181
rect 2508 205 2560 1181
rect 2824 205 2876 1181
rect 3140 205 3192 1181
<< metal2 >>
rect 296 2786 348 2796
rect 296 1544 348 1810
rect 296 1181 348 1440
rect 296 195 348 205
rect 612 2786 664 2796
rect 612 1544 664 1810
rect 612 1181 664 1440
rect 612 195 664 205
rect 928 2786 980 2796
rect 928 1544 980 1810
rect 928 1181 980 1440
rect 928 195 980 205
rect 1244 2786 1296 2796
rect 1244 1544 1296 1810
rect 1244 1181 1296 1440
rect 1244 195 1296 205
rect 1560 2786 1612 2796
rect 1560 1544 1612 1810
rect 1560 1181 1612 1440
rect 1560 195 1612 205
rect 1876 2786 1928 2796
rect 1876 1544 1928 1810
rect 1876 1181 1928 1440
rect 1876 195 1928 205
rect 2192 2786 2244 2796
rect 2192 1544 2244 1810
rect 2192 1181 2244 1440
rect 2192 195 2244 205
rect 2508 2786 2560 2796
rect 2508 1544 2560 1810
rect 2508 1181 2560 1440
rect 2508 195 2560 205
rect 2824 2786 2876 2796
rect 2824 1544 2876 1810
rect 2824 1181 2876 1440
rect 2824 195 2876 205
rect 3140 2786 3192 2796
rect 3140 1544 3192 1810
rect 3140 1181 3192 1440
rect 3140 195 3192 205
use sky130_fd_pr__nfet_g5v0d10v5_BRTJC6  sky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0
timestamp 1654572275
transform 1 0 1744 0 1 693
box -1779 -758 1779 758
use sky130_fd_pr__pfet_g5v0d10v5_CADZ46  sky130_fd_pr__pfet_g5v0d10v5_CADZ46_0
timestamp 1654572275
transform 1 0 1744 0 1 2298
box -1809 -797 1809 797
<< labels >>
flabel metal1 -54 1487 -54 1487 1 FreeSans 400 0 0 0 esd
flabel metal1 30 2927 30 2927 1 FreeSans 400 0 0 0 VDD
flabel metal1 30 71 30 71 1 FreeSans 400 0 0 0 VSS
<< end >>
