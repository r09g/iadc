* NGSPICE file created from clock_flat.ext - technology: sky130A

.subckt clock_flat clk p2d_b p2d p2_b p2 p1d_b p1d p1_b p1 Ad_b Ad A_b A Bd_b Bd B_b
+ B VDD VSS
X0 VSS a_6941_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS sky130_fd_pr__nfet_01v8 ad=2.2138e+14p pd=2.39592e+09u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1 VDD a_5653_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD sky130_fd_pr__pfet_01v8_hvt ad=3.8151e+14p pd=3.51993e+09u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2 a_9876_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8162_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X5 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6 VSS a_501_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X7 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X8 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X9 a_n1738_n6671# a_n2602_n7037# a_n1995_n6925# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X10 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X11 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X12 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X13 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X14 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X15 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_4661_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X16 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X17 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X18 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X19 a_9876_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X20 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X21 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X22 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X23 a_3077_n1909# a_3176_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X24 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u
X25 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X26 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_7237_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_9517_n4709# a_9616_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X28 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X29 VDD a_2148_n3799# a_1888_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X30 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X31 VDD a_7130_n10301# a_7237_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X32 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X33 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6874_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X34 VDD sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X35 VDD a_8418_n6493# a_8525_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X36 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X37 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X38 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X39 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X40 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X41 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X42 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X43 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X44 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X45 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 a_6012_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X47 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X48 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X49 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X50 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X51 VSS a_3436_n9783# a_3176_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X52 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X53 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X54 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X55 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X56 a_9706_n8125# a_9450_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X57 a_8418_n1597# a_8162_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X58 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X59 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X60 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X61 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X62 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_3373_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X63 a_3077_n3621# a_3176_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X64 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X65 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X67 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X68 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X69 VSS sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X70 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X71 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X72 VSS sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X73 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X74 VDD a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X75 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X76 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X77 VSS a_501_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X78 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X79 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X80 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X81 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X82 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X84 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X85 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X86 VSS sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X87 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X88 VDD sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X89 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X90 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X91 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X92 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X93 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X95 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X96 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X97 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 a_11164_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X99 VSS sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_1_0/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X100 VDD clk sky130_fd_sc_hd__clkinv_1_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X101 a_7130_n509# a_6874_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X102 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X103 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X104 VDD a_3436_n13591# a_3176_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X105 a_5842_n11933# a_5586_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X106 VDD sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X107 a_3077_n8437# a_3176_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X108 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X109 VDD a_9706_n5405# a_9813_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X110 a_3266_n10301# a_3010_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X111 VDD a_6012_n8695# a_5752_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X112 VSS a_7130_n8125# a_7237_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X113 a_10805_n5797# a_10904_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X114 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X115 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X116 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X117 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 VDD a_8588_n8695# a_8328_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X119 VDD a_501_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X120 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X121 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X122 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X123 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X124 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_3373_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X125 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X126 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X127 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4298_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X128 VSS a_n1995_n6925# a_n2037_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X129 VSS a_5842_n13021# a_5949_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X130 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X131 a_5653_n12325# a_5752_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X132 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X133 sky130_fd_sc_hd__nand2_4_2/B a_9813_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X134 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X135 a_501_n3621# a_600_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X136 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_8525_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X137 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X138 VDD a_5653_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X139 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_10738_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X140 a_4365_n11237# a_4464_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X141 VDD a_4554_n10301# a_4661_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X142 VSS a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X143 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X144 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X145 VDD a_9706_n2685# a_9813_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X146 a_8418_n5405# a_8162_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X147 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X148 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=9.408e+11p pd=1.12e+07u as=0p ps=0u w=420000u l=150000u
X149 a_7130_n4317# a_6874_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X150 VDD a_3436_n12503# a_3176_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X151 VDD a_690_n10301# a_797_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X152 a_8229_n821# a_8328_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X153 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_6874_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X154 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_3373_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X155 VDD sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 VSS a_6012_n13591# a_5752_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X157 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_2085_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X158 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X159 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_9813_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X160 VDD a_4554_n5405# a_4661_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X161 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u
X162 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X163 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X164 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X165 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X166 a_860_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X167 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_797_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X168 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X169 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_8525_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X171 VSS sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X173 VDD a_3436_n8695# a_3176_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X174 VDD sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X175 a_1978_n10301# a_1722_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X176 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_9813_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X177 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_8525_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X178 VDD a_3077_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X179 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X180 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X181 a_8418_n14109# a_8162_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X182 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X183 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X184 a_8588_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X185 a_2622_n509# a_2366_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X186 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X187 VSS sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X188 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X189 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_1722_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X190 VDD a_4554_n2685# a_4661_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X191 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X192 a_7300_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X193 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_9813_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X194 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X195 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X196 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X197 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X198 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X199 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X200 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X201 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X202 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_5949_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X203 VDD a_690_n4317# a_797_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X204 a_690_n9213# a_434_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X205 VDD sky130_fd_sc_hd__clkinv_1_0/Y a_2366_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X206 a_4554_n4317# a_4298_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X207 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X208 VSS a_5842_n4317# a_5949_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X209 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X210 VSS a_501_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X211 VDD a_3077_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X212 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_6006_n7607# a_6101_n7254# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X214 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X216 a_5842_n2685# a_5586_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X217 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 a_n2436_n7037# a_n2602_n7037# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X219 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X220 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X221 VSS a_8418_n4317# a_8525_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X222 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X223 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X224 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X225 VSS sky130_fd_sc_hd__nand2_4_0/B a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X226 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X227 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X228 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X229 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X230 VDD a_4365_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X231 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X232 a_10994_n5405# a_10738_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X233 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_8525_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X234 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X235 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X236 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X237 a_n2436_n7037# a_n2602_n7037# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X238 a_4724_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X239 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_7237_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X240 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X241 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 VDD a_10994_n9213# a_11101_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X243 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9450_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X244 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X245 VDD a_5842_n11933# a_5949_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X246 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X247 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X248 VSS a_n428_n4887# a_n688_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X249 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_434_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X250 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X251 VDD a_7300_n3799# a_7040_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X252 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_797_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X253 VSS a_501_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_59/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X254 a_n787_n12325# a_n688_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X255 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X256 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X257 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X258 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X259 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X260 a_1789_n11237# a_1888_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X261 VDD a_9876_n3799# a_9616_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X262 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X263 VDD sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X264 a_5653_n2997# a_5752_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X265 VDD a_8588_n13591# a_8328_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X266 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X267 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X268 a_1978_n4317# a_1722_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X269 a_10994_n2685# a_10738_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X270 VSS a_3266_n4317# a_3373_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X271 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_9706_n9213# a_9450_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X273 VDD a_7300_n11415# a_7040_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X274 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X275 a_1789_n10613# a_1888_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X276 VSS a_3077_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X277 sky130_fd_sc_hd__dfxbp_1_1/D a_n1139_n6715# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X278 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_9450_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X279 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X280 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X281 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X282 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X283 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X284 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X285 VSS a_7130_n14109# a_7237_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X286 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X287 VDD a_6006_n7607# sky130_fd_sc_hd__dfxbp_1_0/Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X288 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X289 VSS a_n428_n9783# a_n688_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X290 VDD a_501_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_59/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X291 a_11164_n5975# sky130_fd_sc_hd__clkinv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X292 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X293 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_11101_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X294 VSS a_7300_n10871# a_7040_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X295 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X296 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X297 VDD a_10994_n10301# a_11101_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X298 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X299 VDD a_9706_n10301# a_9813_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X300 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X301 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_3373_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X302 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X303 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X304 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X305 VDD sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X306 sky130_fd_sc_hd__nand2_4_2/B a_9813_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X307 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X308 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6874_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X309 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X310 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_8525_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X311 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X312 a_5653_n1909# a_5752_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X313 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X314 VDD a_8588_n12503# a_8328_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X315 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X317 VDD a_4724_n3799# a_4464_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X318 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X319 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X320 VSS sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X321 VDD a_6012_n5975# a_5752_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X322 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_7237_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X323 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X324 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X325 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X326 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X327 VSS sky130_fd_sc_hd__nand2_4_3/B a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X328 VSS sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X329 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X330 VDD sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X331 a_8588_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X332 VDD sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X333 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_5949_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X334 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1722_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X335 VDD a_7130_n9213# a_7237_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X336 VDD a_4623_n7349# sky130_fd_sc_hd__mux2_1_0/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X337 VSS sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X338 VDD a_8588_n5975# a_8328_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X339 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X340 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X341 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X342 a_11164_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X343 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_10738_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X344 VDD sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X345 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X346 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X347 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X348 VSS sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X349 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_3373_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X350 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 VSS a_5842_n9213# a_5949_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X352 a_5653_n3621# a_5752_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X353 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X354 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X355 a_6794_n7203# a_6658_n7363# a_6373_n7349# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X356 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X357 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X358 VSS a_3077_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X359 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X360 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_3373_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X361 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X362 VSS a_8418_n9213# a_8525_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X363 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X364 a_7130_n1597# a_6874_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X365 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X366 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X367 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X368 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X369 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X370 VDD sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X371 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X372 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X373 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X374 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X375 VDD sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X376 a_n860_n6173# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X377 a_1978_n13021# a_1722_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X378 a_6941_n10613# a_7040_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X379 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_3010_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X380 a_11164_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X381 a_7300_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X382 VDD a_3436_n5975# a_3176_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X383 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X386 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X387 a_10805_n13413# a_10904_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X388 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X389 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X390 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X391 VDD a_2622_n8125# a_2729_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X392 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X393 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 a_5653_n8437# a_5752_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X395 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X396 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X397 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X398 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X399 a_8418_n5405# a_8162_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X400 a_8588_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X401 VSS a_n1738_n6671# a_n1570_n6769# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X402 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X403 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X404 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_11101_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X405 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X406 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5586_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X407 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X408 VSS a_1978_n2685# a_2085_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X409 a_n428_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X410 VSS a_5653_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X411 VSS a_3266_n9213# a_3373_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X412 VSS a_9517_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X413 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X414 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X415 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X416 VSS a_1789_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X417 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X418 VSS a_4365_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X419 VDD a_501_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X420 VDD a_690_n1597# a_797_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X421 VDD a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X422 a_11164_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X423 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X424 a_n2037_n7037# a_n2436_n7037# a_n2163_n6671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X425 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X426 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X427 a_4554_n1597# a_4298_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X428 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X429 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X430 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X431 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X432 a_8418_n10301# a_8162_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X433 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X434 VDD a_2148_n10871# a_1888_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X435 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X436 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X437 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_9450_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X438 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X439 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X440 a_8418_n2685# a_8162_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X441 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X442 VSS a_n787_n12325# sky130_fd_sc_hd__nand2_1_4/B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X443 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X444 a_3077_n4709# a_3176_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X445 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X446 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X447 VDD sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X448 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X449 sky130_fd_sc_hd__clkdlybuf4s50_1_31/X a_11101_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X450 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X452 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X453 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X454 a_n428_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X455 VDD a_5653_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X456 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X457 VDD a_9517_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X458 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X460 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X461 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X462 a_n787_n1909# a_n688_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X463 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X464 VSS a_11164_n5975# a_10904_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X465 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X466 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X467 VDD a_2148_n3255# a_1888_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X468 VDD a_4365_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X469 a_6941_n2997# a_7040_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X470 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_434_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X471 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X472 a_11164_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X473 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X474 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X475 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X476 a_7300_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X477 VDD a_4365_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X478 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4298_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X479 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X480 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X481 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X482 VDD a_n787_n12325# sky130_fd_sc_hd__nand2_1_4/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X483 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.24e+12p pd=2.048e+07u as=0p ps=0u w=1e+06u l=150000u
X484 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X485 a_2148_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X486 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_5949_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X487 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X488 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_4661_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X489 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X490 a_2622_n6493# a_2366_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X491 VDD sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X492 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X493 a_9517_n5797# a_9616_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X494 a_6941_n821# a_7040_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X495 a_1978_n1597# a_1722_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X496 a_4724_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X497 a_501_n10613# a_600_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X498 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X499 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X500 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7237_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X501 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_6874_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X502 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_8525_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X503 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X504 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X505 VSS sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X506 a_2622_n14109# a_2366_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X507 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9813_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X508 VSS a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X509 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X510 VSS a_11164_n4887# a_10904_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X511 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8162_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X512 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_1_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X513 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X515 a_13765_n1597# sky130_fd_sc_hd__clkinv_4_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X516 VDD a_2148_n2167# a_1888_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X517 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X518 a_11164_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X519 a_6941_n1909# a_7040_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X520 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X521 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=0p ps=0u w=840000u l=150000u
X522 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X523 a_5653_n13413# a_5752_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X524 a_6941_n9525# a_7040_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X525 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X526 VSS a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X527 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X528 a_2148_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X529 VDD a_9706_n8125# a_9813_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X530 VSS sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X531 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X532 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X533 VSS a_860_n3255# a_600_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X534 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X535 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__mux2_1_0/X a_3832_n7261# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X536 a_7130_n509# a_6874_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X537 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X539 a_8229_n11237# a_8328_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X540 a_4365_n2997# a_4464_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X541 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X542 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X543 a_4724_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X544 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_7237_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X545 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X546 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X547 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X548 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_797_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X549 a_9517_n4709# a_9616_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X550 VDD sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X551 VSS a_2148_n3799# a_1888_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X552 VSS a_7130_n10301# a_7237_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X553 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X554 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X555 VDD a_4365_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X556 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X557 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X558 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_8525_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X559 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9450_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X560 a_8229_n10613# a_8328_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X561 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X562 a_7130_n11933# a_6874_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X563 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X564 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X565 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_2085_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X566 VSS a_11164_n9783# a_10904_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X567 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X568 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X569 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X570 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X571 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X572 a_5653_n12325# a_5752_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X573 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_4661_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X574 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X575 a_501_n2997# a_600_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X576 a_8229_n3621# a_8328_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X577 VSS a_9706_n14109# a_9813_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X578 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X579 a_6941_n12325# a_7040_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X580 VDD a_n787_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X581 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X582 VSS a_860_n2167# a_600_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X583 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X584 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_7237_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X585 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X586 a_4365_n1909# a_4464_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X587 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X588 VDD a_860_n9783# a_600_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X589 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X590 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X591 VDD a_5842_n10301# a_5949_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X592 a_4365_n9525# a_4464_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X593 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X595 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X596 a_9517_n9525# a_9616_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X597 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9450_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X598 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 VSS a_2148_n8695# a_1888_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X600 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X601 VSS a_3266_n13021# a_3373_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X602 sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_2085_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X603 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X604 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X605 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X606 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X607 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X608 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X609 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X610 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6874_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X611 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X612 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X613 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X614 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X615 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_8162_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X616 a_1789_n2997# a_1888_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X617 a_8418_n14109# a_8162_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X618 a_1789_n11237# a_1888_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X619 a_7300_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X620 VSS a_n1570_n6769# a_n1612_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X621 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_11101_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X622 VSS a_1978_n11933# a_2085_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X623 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X625 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X626 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X627 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X628 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_4661_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X629 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X630 a_n2248_n7037# sky130_fd_sc_hd__dfxbp_1_1/D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X631 VSS sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X633 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X634 a_501_n1909# a_600_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X635 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_9450_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X636 VSS a_4365_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X637 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6874_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X638 VSS a_2622_n6493# a_2729_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X639 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X640 VSS a_3436_n13591# a_3176_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X641 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X642 VSS a_7300_n11415# a_7040_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X643 a_2622_n509# a_2366_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X644 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X645 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X646 a_3266_n10301# a_3010_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X647 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X648 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X649 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X650 VDD sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X651 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X652 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_5586_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X653 a_9706_n6493# a_9450_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X654 VSS a_2148_n12503# a_1888_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X655 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X656 VSS sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X657 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X658 a_n860_n509# sky130_fd_sc_hd__nand2_1_0/B VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X659 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X660 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X661 VSS a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X662 VDD a_5842_n4317# a_5949_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X663 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X664 VDD a_10805_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X665 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X666 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X667 VSS a_3077_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X668 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X669 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X670 a_1789_n1909# a_1888_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X671 a_501_n3621# a_600_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X672 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X673 a_8418_n13021# a_8162_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X674 VDD a_8418_n4317# a_8525_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X675 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X676 VSS a_4554_n10301# a_4661_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X677 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X678 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X679 a_1789_n9525# a_1888_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X680 a_2148_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X681 VSS a_9706_n2685# a_9813_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X682 VDD a_9517_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X683 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X684 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_3373_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X685 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X686 VDD a_8229_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X687 a_4724_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X688 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X689 a_9517_n10613# a_9616_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X690 VSS a_690_n10301# a_797_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X691 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X692 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X693 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_2729_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X694 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X695 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X696 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X697 a_4724_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X698 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3010_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X699 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X700 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X702 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X703 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A a_5949_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X704 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X705 VDD a_11164_n8695# a_10904_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X706 VSS a_1789_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X707 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X708 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_4298_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X709 VSS sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X710 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_5586_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X711 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_6874_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X712 VDD a_10805_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X713 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X714 VDD a_7130_n6493# a_7237_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X715 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X716 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X717 VSS sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X718 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X719 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X720 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X721 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X722 VDD sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X723 a_501_n12325# a_600_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X724 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 a_501_n8437# a_600_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X726 a_2148_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X727 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_434_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X728 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X729 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X730 sky130_fd_sc_hd__clkinv_1_6/Y clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X731 VDD a_7300_n3255# a_7040_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X732 a_7130_n1597# a_6874_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X733 VDD a_3266_n4317# a_3373_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X734 a_3266_n9213# a_3010_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X735 VDD a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X736 VDD a_6101_n7254# sky130_fd_sc_hd__dfxbp_1_0/Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X737 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X738 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X739 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_2085_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X740 VDD a_9876_n3255# a_9616_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X741 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X742 a_6865_n7304# a_6665_n7459# a_7014_n7215# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.392e+11p ps=1.53e+06u w=360000u l=150000u
X743 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X744 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X745 VSS a_4554_n2685# a_4661_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X746 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X747 a_9517_n8437# a_9616_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X748 VSS a_10805_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X749 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X750 VDD a_7130_n14109# a_7237_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X751 VDD a_3266_n11933# a_3373_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X752 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X753 VDD a_1789_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X754 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_4298_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X755 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X756 a_3077_n11237# a_3176_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X757 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X758 VDD a_6941_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X759 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X760 VDD a_5653_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X761 a_10994_n13021# a_10738_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X762 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X763 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_797_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X764 VSS a_9517_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X765 a_3077_n10613# a_3176_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X766 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X768 VDD a_7300_n2167# a_7040_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X769 a_10805_n2997# a_10904_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X770 a_5653_n4709# a_5752_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X771 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X772 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X773 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1722_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X774 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X775 a_690_n4317# a_434_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X776 VSS a_9706_n6493# a_9813_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X777 VSS sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X778 VSS a_9517_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X779 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X780 VDD a_4724_n11415# a_4464_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X781 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X782 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X783 VDD a_9876_n2167# a_9616_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X784 VDD a_10805_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X785 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_6874_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X786 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X787 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X789 VDD a_7130_n13021# a_7237_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X790 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X791 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X792 VSS a_690_n1597# a_797_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X793 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X794 VDD a_4724_n3255# a_4464_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X795 VDD a_860_n11415# a_600_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X796 a_4554_n1597# a_4298_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X797 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X798 VSS a_8418_n13021# a_8525_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X799 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X800 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_797_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X801 VSS a_4724_n10871# a_4464_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X802 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_9813_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X803 VDD a_6941_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X804 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_8525_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X805 VSS a_7300_n3799# a_7040_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X806 VDD sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X807 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X808 VDD a_9517_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X809 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4298_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X810 VSS a_8229_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X811 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X812 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X813 VSS a_860_n10871# a_600_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X814 VDD sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X815 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_1722_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X816 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X817 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_8525_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X818 VSS a_10994_n4317# a_11101_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X819 a_10805_n1909# a_10904_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X820 VSS a_9876_n3799# a_9616_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X821 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_3010_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X822 a_7130_n5405# a_6874_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X823 VSS a_8588_n13591# a_8328_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X824 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X825 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_5949_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X826 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_4661_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X827 a_10805_n9525# a_10904_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X828 a_10994_n2685# a_10738_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X829 VDD sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X830 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X831 a_6941_n821# a_7040_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X832 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X833 VSS a_6941_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X834 a_6373_n7349# a_6665_n7459# a_6616_n7581# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X835 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X836 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9450_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X837 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X838 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X839 VDD a_4724_n2167# a_4464_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X840 sky130_fd_sc_hd__nand2_4_1/B a_9813_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X841 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X842 a_9876_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X843 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X844 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X845 a_9706_n4317# a_9450_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X846 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X847 VSS a_7300_n8695# a_7040_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X848 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X849 VSS a_10805_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X850 a_13765_n5405# sky130_fd_sc_hd__clkinv_4_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X851 VSS a_10994_n10301# a_11101_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X852 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X853 VSS a_9706_n10301# a_9813_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X854 a_8418_n8125# a_8162_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X855 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X856 a_9706_n11933# a_9450_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X857 VSS sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X858 a_1978_n1597# a_1722_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X859 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_5/A a_n860_n6173# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X860 VSS a_9876_n8695# a_9616_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X861 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X862 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nand2_1_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=0p ps=0u w=840000u l=150000u
X863 a_3266_n13021# a_3010_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X864 a_n860_n8125# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X865 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X866 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X867 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X868 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X869 VSS a_4724_n3799# a_4464_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X870 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X871 VDD a_6941_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X872 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_797_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X873 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X874 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_9450_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X875 VSS a_9517_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X876 VDD a_1789_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X877 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X878 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X879 a_4365_n10613# a_4464_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X880 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X881 a_10994_n11933# a_10738_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X882 VSS a_690_n5405# a_797_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X883 a_9517_n12325# a_9616_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X884 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X885 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A a_5949_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X886 VDD a_5842_n1597# a_5949_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X887 a_9876_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X888 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_3010_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X889 a_4554_n5405# a_4298_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X890 VSS sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X891 VSS clk a_n2602_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X892 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X893 VDD a_860_n1079# a_600_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X894 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X895 VSS a_n1570_n6769# a_n1139_n6715# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X896 a_4365_n821# a_4464_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X897 VDD sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_1_0/B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.268e+11p ps=2.22e+06u w=840000u l=150000u
X898 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X899 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X900 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X901 VDD a_4554_n13021# a_4661_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X902 a_8229_n11237# a_8328_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X903 a_7300_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X904 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X905 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X906 VDD a_8418_n1597# a_8525_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X907 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6874_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X908 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X909 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X910 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X911 VSS a_7130_n4317# a_7237_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X912 VDD a_690_n13021# a_797_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X913 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X914 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_7237_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X915 VDD clk a_n2602_n7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X916 a_13765_n13565# sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X917 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X918 VSS a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X919 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X920 a_n787_n4709# a_n688_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X921 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X922 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X923 a_690_n9213# a_434_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X924 VSS a_4724_n8695# a_4464_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X925 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X926 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X927 VDD a_8418_n11933# a_8525_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X928 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X929 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X931 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X932 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X933 a_6012_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X934 VDD a_11164_n5975# a_10904_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X935 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X936 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X937 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X938 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X939 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X940 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X941 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_797_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X942 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X943 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_6874_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X944 VSS a_6941_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X945 a_3436_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X946 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X947 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X948 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X949 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X950 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X951 a_3077_n5797# a_3176_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X952 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X953 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_2085_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X954 a_1978_n5405# a_1722_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X955 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X956 VSS a_n787_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X957 VDD a_3266_n1597# a_3373_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X958 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X959 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X960 VDD a_11164_n11415# a_10904_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X961 VDD a_6941_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X962 VSS a_10994_n9213# a_11101_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X963 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X964 a_2622_n14109# a_2366_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X965 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X966 VDD a_9876_n11415# a_9616_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X967 a_2148_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X968 a_1789_n821# a_1888_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X969 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X970 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X971 a_9876_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X972 a_9517_n5797# a_9616_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X973 VDD a_2148_n4887# a_1888_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X974 a_n2163_n6671# a_n2436_n7037# a_n2248_n7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X975 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X976 a_860_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X977 VDD sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X978 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X979 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X980 VSS a_11164_n10871# a_10904_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X981 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X982 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A a_5949_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X983 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_133/A a_1722_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X984 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X985 VSS a_9876_n10871# a_9616_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X986 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_10738_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X987 a_6012_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X988 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X989 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X990 a_860_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X991 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X992 a_8418_n2685# a_8162_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X993 VDD sky130_fd_sc_hd__clkinv_1_5/A a_7212_n7203# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X994 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X995 sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_3373_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X996 a_9706_n9213# a_9450_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X997 VSS a_6012_n3255# a_5752_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X998 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_5586_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X999 a_3077_n4709# a_3176_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1000 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1001 a_6941_n13413# a_7040_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1002 VSS sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1003 VSS sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1004 VSS a_4724_n1079# a_4464_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1005 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1006 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3010_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1007 VSS a_8588_n3255# a_8328_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1008 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A a_8525_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1009 VDD a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1010 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1011 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_434_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1012 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1013 a_3832_n7261# sky130_fd_sc_hd__nand2_1_4/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1014 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1015 VSS a_501_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1016 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1017 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1018 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1019 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1020 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1021 VSS a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1022 VSS a_n787_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1023 VDD a_9706_n14109# a_9813_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1024 a_5842_n9213# a_5586_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1025 a_860_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1026 a_9876_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1027 sky130_fd_sc_hd__nand2_4_0/B a_9813_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1028 VSS a_3436_n1079# a_3176_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1029 VSS a_6012_n2167# a_5752_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1030 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1031 a_5842_n13021# a_5586_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1032 VDD sky130_fd_sc_hd__clkinv_4_7/A a_13765_n13565# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1034 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1035 a_3077_n9525# a_3176_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1036 a_8229_n2997# a_8328_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1037 a_6941_n12325# a_7040_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1038 VDD a_6012_n9783# a_5752_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1039 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1040 VSS a_7130_n9213# a_7237_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1041 a_n1995_n6925# a_n2163_n6671# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X1042 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1043 VSS a_8588_n2167# a_8328_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1044 VDD a_2148_n13591# a_1888_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1045 a_4554_n11933# a_4298_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1046 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1047 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1048 a_6012_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1049 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1050 VDD a_501_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_78/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1051 VDD a_8588_n9783# a_8328_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1052 VSS a_3436_n3255# a_3176_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1053 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1055 VDD a_501_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1056 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1057 VSS a_2148_n1079# a_1888_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1058 a_690_n11933# a_434_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1059 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1060 a_860_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1061 VDD sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1062 a_5653_n13413# a_5752_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1063 a_7041_n7581# a_6794_n7203# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X1064 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_3010_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1065 VDD a_10994_n13021# a_11101_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1066 a_501_n4709# a_600_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1067 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1068 VDD a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1069 VDD a_9706_n13021# a_9813_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1070 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1071 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1072 a_4365_n12325# a_4464_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1073 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_5949_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1074 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_7237_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1075 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1076 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_7237_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1077 a_8418_n6493# a_8162_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1078 a_8588_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1079 a_7130_n5405# a_6874_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1080 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1081 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1082 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1083 a_3077_n11237# a_3176_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1084 VDD a_3266_n10301# a_3373_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1085 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1086 a_8229_n1909# a_8328_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1087 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6874_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1088 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1089 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1090 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1091 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_9813_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1092 VDD a_2148_n12503# a_1888_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1093 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1094 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1095 VSS sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1096 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/X a_434_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1097 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 a_10805_n821# a_10904_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1099 VSS a_3436_n2167# a_3176_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1100 a_6865_n7304# a_6658_n7363# a_7041_n7581# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1101 VSS a_2622_n8125# a_2729_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1102 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_797_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1103 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1104 VSS a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1105 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1106 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1107 a_860_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1108 VSS sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1109 VDD a_3436_n9783# a_3176_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1110 VDD a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1111 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1112 a_501_n13413# a_600_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1113 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1114 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8162_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1115 VSS a_4724_n11415# a_4464_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1116 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A a_5949_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1117 a_6012_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1118 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_8525_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1119 a_8229_n3621# a_8328_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1120 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1121 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1122 a_7130_n2685# a_6874_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1123 a_8588_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1124 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1125 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_7237_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1126 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1127 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1128 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1129 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1130 VSS a_860_n11415# a_600_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1131 a_n2163_n6671# a_n2602_n7037# a_n2248_n7037# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X1132 VDD a_n1570_n6769# a_n1139_n6715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1133 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1134 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_797_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1135 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1136 VSS sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1137 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1138 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1139 a_7300_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1140 a_3436_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1141 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_9813_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1142 VSS a_5842_n10301# a_5949_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1143 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1144 VDD sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkinv_1_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1145 a_11164_n5975# sky130_fd_sc_hd__clkinv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1146 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1147 VSS sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1148 a_6012_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1149 VDD a_1789_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1150 VDD a_690_n5405# a_797_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1151 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1152 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1153 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1154 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1155 a_4554_n5405# a_4298_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1156 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1157 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1158 VDD a_3077_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1159 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1160 a_501_n12325# a_600_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1161 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1162 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1163 a_5842_n11933# a_5586_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1164 VDD a_9517_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1165 a_3077_n8437# a_3176_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1166 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1167 a_8229_n8437# a_8328_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1168 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1169 sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_797_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1170 a_860_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1171 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1172 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9450_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1173 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1174 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1175 a_11164_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1176 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1177 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1178 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_5586_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1179 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_8525_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1180 VDD sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 VDD a_690_n2685# a_797_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1182 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1183 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1184 a_4554_n2685# a_4298_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1185 VSS a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1186 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_9450_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1187 sky130_fd_sc_hd__clkdlybuf4s50_1_157/A a_11101_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1188 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1189 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_8162_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1190 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=0p ps=0u w=1e+06u l=150000u
X1191 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1192 VSS a_10805_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1193 VSS a_4365_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1194 a_n1995_n6925# a_n2163_n6671# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1195 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1196 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1197 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_59/A a_434_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1198 VDD a_7300_n4887# a_7040_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1199 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1200 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1201 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1202 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1203 a_690_n4317# a_434_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1204 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1205 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1206 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1207 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1208 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1209 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1210 VDD a_9876_n4887# a_9616_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1211 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1212 VSS a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1213 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1214 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1215 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X1216 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1217 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1218 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1219 a_1978_n5405# a_1722_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1220 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1221 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1222 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1223 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 a_3436_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1225 VSS a_5842_n1597# a_5949_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1226 a_10994_n10301# a_10738_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1227 VDD a_1978_n9213# a_2085_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1228 a_8588_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1229 VDD a_3077_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1230 a_7300_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1231 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1232 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1233 VDD a_10805_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1234 VDD a_6012_n11415# a_5752_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1235 VSS a_8418_n1597# a_8525_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1236 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1237 VSS a_9706_n8125# a_9813_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1238 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1239 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_8162_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1240 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1241 VDD a_10994_n4317# a_11101_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1242 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1243 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1244 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_2729_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1245 VDD sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1246 VSS sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1247 a_5653_n5797# a_5752_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1248 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_3373_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1249 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X1250 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1251 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 a_3436_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1254 VSS sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1255 VSS a_6012_n10871# a_5752_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1256 a_6941_n3621# a_7040_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1257 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_5586_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1258 a_1978_n2685# a_1722_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1259 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_6874_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1260 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1261 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1262 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3010_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1263 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1264 VDD a_8418_n10301# a_8525_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1265 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1266 VDD a_4724_n4887# a_4464_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1267 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1268 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1269 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_7237_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1270 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1272 a_8588_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1273 a_3266_n4317# a_3010_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1274 a_9706_n4317# a_9450_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1275 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1276 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_1722_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1277 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_5949_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1278 a_9517_n13413# a_9616_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1279 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1280 VDD a_8229_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1281 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1282 a_2148_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1283 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X1284 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1285 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10738_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1286 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1287 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1288 VSS a_3266_n1597# a_3373_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1289 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A a_3373_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1290 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X1291 VSS a_11164_n11415# a_10904_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1292 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1293 VSS a_9876_n11415# a_9616_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1294 a_3436_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1295 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1296 a_5653_n4709# a_5752_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1297 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1298 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1299 a_4724_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1300 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1301 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_3010_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1302 VSS a_3077_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1303 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5586_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1304 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1305 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1306 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1307 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1308 VSS a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1309 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1310 a_8588_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1311 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1312 VDD sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1313 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_434_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1314 VSS a_5842_n5405# a_5949_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1315 VDD a_860_n3799# a_600_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1316 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1317 VSS sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1318 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1319 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1320 a_4365_n3621# a_4464_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1321 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1322 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1323 VDD a_6012_n1079# a_5752_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1324 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1326 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_4/Y a_n860_n8125# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1327 a_9517_n12325# a_9616_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1328 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1329 VSS a_8418_n5405# a_8525_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1330 VDD a_7130_n4317# a_7237_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1331 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1332 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1333 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1334 VDD a_8588_n1079# a_8328_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1335 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1336 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1337 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1338 a_5653_n9525# a_5752_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1339 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1340 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1341 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9450_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1342 VDD a_5653_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1343 a_8588_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1344 a_n2248_n7037# sky130_fd_sc_hd__dfxbp_1_1/D VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1345 VDD a_5842_n13021# a_5949_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1346 a_1789_n10613# a_1888_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1347 VSS a_8229_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1348 VSS a_n428_n2167# a_n688_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1349 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=0p ps=0u w=420000u l=150000u
X1350 VSS a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1351 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1352 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1353 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_89/A a_2366_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1354 VSS sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1355 VDD a_n428_n9783# a_n688_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1356 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_5586_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1357 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1358 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4298_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1359 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1360 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1361 VDD a_7300_n10871# a_7040_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1362 VSS sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1363 VSS a_4365_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1364 VSS a_8229_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1365 a_4724_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1366 VDD a_501_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1367 a_6101_n7254# a_6373_n7349# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1368 a_11164_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1369 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1370 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_8525_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1371 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/X a_434_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1373 VSS a_3266_n5405# a_3373_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1374 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1375 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_4661_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1376 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1377 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1378 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1379 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1380 VDD a_3436_n1079# a_3176_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1381 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1382 a_1789_n3621# a_1888_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1383 VSS sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1384 a_3077_n5797# a_3176_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1385 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1386 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1387 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_9450_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1388 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1389 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1390 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_8525_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1391 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1392 VDD a_9517_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1393 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1394 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1395 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1396 VSS a_10805_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1397 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A a_11101_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1398 VSS a_4365_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1399 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1400 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1401 VDD a_4365_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1402 VDD a_8229_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1403 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1404 a_7212_n7203# a_6658_n7363# a_6865_n7304# VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=360000u l=150000u
X1405 VDD sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1406 a_11164_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1407 a_3266_n9213# a_3010_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1408 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1409 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1410 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1411 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A a_8525_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1412 a_8588_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1413 VSS a_5653_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1414 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1415 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_7237_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1416 a_9876_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1417 VSS a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1418 VSS a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1419 a_690_n1597# a_434_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1420 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_3010_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1421 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1422 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1423 VDD sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1424 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A a_5949_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1425 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1426 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1427 a_n787_n4709# a_n688_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1428 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1429 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_6874_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1430 VSS a_2148_n5975# a_1888_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1431 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1432 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1433 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1434 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1435 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1436 VSS a_4365_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1437 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1438 a_13765_n9757# sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1439 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_8162_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1440 a_13765_n2685# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1441 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1442 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1443 a_11164_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1444 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1445 a_5653_n8437# a_5752_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1446 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1447 VDD a_10994_n1597# a_11101_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1448 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1449 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1450 a_4365_n13413# a_4464_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1451 VDD a_9706_n9213# a_9813_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1452 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1453 VSS sky130_fd_sc_hd__nand2_4_2/B a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X1454 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1455 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1456 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1457 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1458 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1459 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_0/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1460 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1461 VDD a_1789_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1462 VSS a_8229_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1463 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 a_10805_n11237# a_10904_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1465 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1466 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1467 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1468 a_n787_n9525# a_n688_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1469 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1470 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_797_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1471 VSS a_2148_n4887# a_1888_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1472 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1473 VSS a_5653_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1474 VDD a_4365_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1475 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1476 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1477 VSS a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1478 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9450_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1479 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1480 a_7130_n13021# a_6874_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1481 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1482 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1483 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1484 a_10805_n10613# a_10904_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1485 a_9706_n1597# a_9450_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1486 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1487 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1488 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1489 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1490 a_5842_n10301# a_5586_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1491 VSS sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1492 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1493 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1494 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A a_2729_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1495 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1496 a_7130_n8125# a_6874_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1497 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1498 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1499 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1500 a_8229_n4709# a_8328_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1501 a_4365_n12325# a_4464_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1502 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1503 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1504 a_6941_n13413# a_7040_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1505 a_1978_n11933# a_1722_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1506 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X1507 sky130_fd_sc_hd__nand2_4_3/A clk VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1508 VDD a_4554_n9213# a_4661_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1509 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1510 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1511 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1512 VSS a_8418_n14109# a_8525_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1513 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1514 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1515 a_10805_n3621# a_10904_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1516 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1517 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1518 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_103/A a_9450_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1519 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1520 sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkinv_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1521 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1522 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1523 VSS a_2148_n9783# a_1888_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1524 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1525 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1526 a_8418_n8125# a_8162_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1527 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1528 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1529 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8162_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1530 VSS a_9706_n509# a_9813_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1531 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1532 a_501_n5797# a_600_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1533 VSS a_1978_n13021# a_2085_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1534 a_1789_n12325# a_1888_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1535 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1536 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1537 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1538 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1539 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1540 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1541 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_2085_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1542 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1543 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1544 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1545 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1546 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1547 VDD a_7130_n1597# a_7237_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1548 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5586_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1549 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1550 VSS sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1551 VSS a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1552 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6874_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1553 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1554 VSS a_7300_n12503# a_7040_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1555 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1556 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1557 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1558 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1559 VSS sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X1560 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1561 VSS a_11164_n3255# a_10904_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1562 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1563 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_42/X a_434_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1564 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1565 VSS a_2148_n13591# a_1888_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1566 VSS a_6012_n11415# a_5752_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1567 a_5842_n4317# a_5586_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1568 VSS a_8418_n509# a_8525_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1569 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_10738_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1570 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1571 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1572 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1573 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1574 VDD a_5842_n5405# a_5949_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1575 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_4298_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1576 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1577 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1578 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1579 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1580 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1581 a_501_n4709# a_600_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1582 VDD a_8418_n5405# a_8525_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1583 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1584 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1585 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1586 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_4661_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1587 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_5586_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1588 a_2148_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1589 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1590 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1591 VDD sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1592 VDD a_3077_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1593 a_9517_n2997# a_9616_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1594 a_4724_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1595 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1596 VSS a_3266_n10301# a_3373_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1597 a_10994_n9213# a_10738_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1598 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1599 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/X a_434_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1600 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1601 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_3010_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1602 VSS a_10805_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1603 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1604 VSS a_11164_n2167# a_10904_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1605 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1606 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1607 VDD a_5842_n2685# a_5949_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1608 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1610 a_7130_n11933# a_6874_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1611 a_8229_n10613# a_8328_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1612 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1613 VDD a_4365_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1614 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1615 VDD a_11164_n9783# a_10904_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1616 VSS sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1617 VSS sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1618 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1619 VDD a_8418_n2685# a_8525_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1620 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1621 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1622 a_7014_n7215# a_6794_n7203# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1623 VSS a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1624 VDD a_6941_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1625 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1626 a_501_n13413# a_600_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1627 a_501_n9525# a_600_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1628 sky130_fd_sc_hd__nand2_4_3/B a_9813_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1629 a_7130_n2685# a_6874_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1630 VDD a_3266_n5405# a_3373_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1631 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1632 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6874_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1633 VDD a_501_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1634 a_860_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1635 a_9517_n1909# a_9616_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1636 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1637 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1638 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1639 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1640 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1641 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1642 a_9517_n9525# a_9616_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1643 VSS a_10805_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1644 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_7237_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1645 VDD sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__clkinv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1646 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1647 VDD a_2148_n8695# a_1888_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1648 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_797_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1649 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9450_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1650 VDD sky130_fd_sc_hd__clkinv_4_1/Y a_13765_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1651 VSS a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1652 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1653 a_6012_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1654 VDD a_1978_n11933# a_2085_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1655 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1656 VSS a_7300_n5975# a_7040_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1657 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1658 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1659 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1660 VSS a_9517_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1661 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1662 a_1789_n821# a_1888_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1663 VDD a_3266_n2685# a_3373_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1664 VDD a_2622_n6493# a_2729_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1665 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1666 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1667 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1668 a_5653_n5797# a_5752_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1669 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1670 VSS a_9876_n5975# a_9616_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1671 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1672 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8162_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1673 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1674 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1675 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1676 a_6941_n2997# a_7040_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1677 VDD a_10805_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1678 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1679 a_3266_n4317# a_3010_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1680 VSS a_6941_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1681 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1682 VDD a_3436_n11415# a_3176_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1683 VSS a_690_n2685# a_797_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1684 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1685 a_4554_n2685# a_4298_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1686 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1687 a_5842_n9213# a_5586_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1688 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1689 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1690 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_1_6/Y a_n860_n13789# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1691 VSS a_501_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1692 VSS a_7300_n4887# a_7040_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1693 VDD a_9517_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1694 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1695 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1696 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1697 VSS a_3436_n10871# a_3176_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1698 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_7237_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1699 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1700 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.4e+11p ps=7.68e+06u w=1e+06u l=150000u
X1701 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1702 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1703 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1704 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1705 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1706 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A a_8525_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1707 VSS a_6658_n7363# a_6665_n7459# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1708 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3010_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1709 VSS a_9876_n4887# a_9616_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1710 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A a_7237_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1711 a_11164_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1712 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1713 a_7130_n6493# a_6874_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1714 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9813_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1715 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_8525_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1716 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1717 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8162_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1718 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1719 VSS a_4724_n5975# a_4464_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1720 sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nand2_1_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1721 a_6941_n1909# a_7040_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1722 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1723 sky130_fd_sc_hd__clkinv_1_5/A a_n1570_n6769# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1724 a_10994_n10301# a_10738_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1725 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1726 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1727 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1728 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1729 VDD a_6012_n3799# a_5752_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1730 VSS a_6941_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1731 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1732 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1733 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9450_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1734 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1735 a_13765_n13021# sky130_fd_sc_hd__clkinv_4_7/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1736 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1737 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1738 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1739 VSS a_n428_n12503# a_n688_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1740 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1741 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1742 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1743 VDD a_860_n3255# a_600_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1744 VDD a_8588_n3799# a_8328_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1745 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1746 a_501_n8437# a_600_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1747 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1748 a_690_n1597# a_434_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1749 a_4365_n2997# a_4464_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1750 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_10738_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1751 VSS a_7300_n9783# a_7040_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1752 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1753 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1754 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1755 VSS a_1978_n4317# a_2085_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1756 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1757 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1758 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1759 a_8418_n9213# a_8162_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1760 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1761 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1762 a_6941_n3621# a_7040_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1763 a_9706_n13021# a_9450_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1764 a_1978_n2685# a_1722_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1765 VSS a_9876_n9783# a_9616_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1766 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1767 VSS a_8418_n10301# a_8525_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1768 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1769 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1770 VSS a_4724_n4887# a_4464_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1771 a_8418_n11933# a_8162_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1772 VDD a_6941_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1773 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1774 VSS a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1775 a_9876_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1776 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_9450_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1777 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1778 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1779 VDD a_1789_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1780 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1781 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1782 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1783 VDD a_n787_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_49/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1784 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1785 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1786 a_9517_n13413# a_9616_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1787 VSS a_10994_n1597# a_11101_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1788 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1789 VDD a_860_n2167# a_600_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1790 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1791 a_3077_n10613# a_3176_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1792 a_11164_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1793 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1794 a_4365_n1909# a_4464_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1795 a_8229_n12325# a_8328_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1796 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1797 VDD a_3436_n3799# a_3176_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1798 VSS sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1799 a_10805_n11237# a_10904_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1800 VSS sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1801 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6874_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1802 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1803 VDD a_9706_n6493# a_9813_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1804 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_6874_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1805 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1806 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1807 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1808 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1809 VDD a_3266_n13021# a_3373_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1810 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1811 a_6941_n8437# a_7040_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1812 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1813 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1814 a_7300_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1815 a_6012_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1816 VDD a_1789_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1817 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1818 VDD a_10805_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1819 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1820 VSS a_6941_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1821 a_1789_n2997# a_1888_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1822 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1823 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1824 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1825 VSS a_4724_n9783# a_4464_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1826 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1827 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1828 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_5949_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1829 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1722_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1830 a_9706_n1597# a_9450_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1831 VDD a_4724_n10871# a_4464_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1832 VSS a_860_n3799# a_600_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1833 VSS a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1834 a_4365_n3621# a_4464_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1835 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1836 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1837 VSS sky130_fd_sc_hd__nand2_4_1/B a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X1838 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1839 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1840 sky130_fd_sc_hd__nand2_4_0/B a_9813_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1841 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1842 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1843 VSS a_3077_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1844 VDD a_860_n10871# a_600_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1845 VSS a_2622_n14109# a_2729_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1846 VDD a_9517_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1847 a_690_n5405# a_434_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1848 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1849 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_6874_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1850 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1851 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_6874_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1852 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1853 sky130_fd_sc_hd__clkdlybuf4s50_1_100/A sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=0p ps=0u w=840000u l=150000u
X1854 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1855 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1856 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1857 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1858 VDD a_6941_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1859 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1860 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1861 a_2148_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1862 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_797_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X1863 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1864 a_2148_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1865 a_1789_n1909# a_1888_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1866 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1867 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1868 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1869 a_9876_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1870 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1871 a_n428_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1872 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10738_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1873 a_6012_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1874 VDD sky130_fd_sc_hd__clkinv_4_7/Y a_13765_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1875 VDD a_8588_n11415# a_8328_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1876 VDD a_5653_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1877 VDD a_2148_n5975# a_1888_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1878 a_860_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1879 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1880 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1881 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1882 VSS a_860_n8695# a_600_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1883 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1884 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1885 a_4365_n8437# a_4464_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1886 VDD a_7300_n8695# a_7040_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1887 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1888 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1889 VSS a_7130_n1597# a_7237_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1890 VSS a_10994_n5405# a_11101_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1891 a_7300_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1892 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1893 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1894 VSS a_8588_n10871# a_8328_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1895 VDD a_11164_n1079# a_10904_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1896 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1897 a_9706_n11933# a_9450_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1898 VSS a_7130_n11933# a_7237_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1899 VDD sky130_fd_sc_hd__clkinv_1_5/A sky130_fd_sc_hd__nand2_4_1/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1900 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1901 VDD a_9876_n8695# a_9616_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1902 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_11101_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1903 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1904 VSS a_1978_n9213# a_2085_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1905 a_1789_n3621# a_1888_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1906 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_5586_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1907 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10738_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1908 VDD a_n1570_n6769# a_n1654_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X1909 VDD sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1910 VDD a_10805_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1911 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1912 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1913 a_4724_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1914 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1915 VDD a_6941_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X1916 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1917 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1918 a_3266_n1597# a_3010_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1919 a_6012_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1920 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/A a_434_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1921 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1922 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_8162_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1923 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_3373_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1924 a_9706_n5405# a_9450_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1925 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1926 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1927 a_3436_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1928 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1929 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1930 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1931 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1932 a_9517_n821# a_9616_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1933 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1934 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1935 a_n1612_n7037# a_n2602_n7037# a_n1738_n6671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X1936 a_1789_n13413# a_1888_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1937 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1938 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_10738_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1939 a_2148_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1940 a_n428_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1941 VSS a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X1942 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1943 VDD a_8418_n14109# a_8525_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1944 VSS clk sky130_fd_sc_hd__clkinv_1_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1945 VSS a_9876_n1079# a_9616_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1946 a_1789_n8437# a_1888_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1947 VDD a_7300_n13591# a_7040_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1948 VDD a_4724_n8695# a_4464_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1949 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1950 a_10994_n13021# a_10738_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1951 a_7130_n10301# a_6874_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1952 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1953 a_4724_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1954 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1955 VDD a_13765_n13021# p1_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1956 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1957 a_4554_n13021# a_4298_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1958 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1959 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1960 a_6012_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1961 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1962 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1963 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1964 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1965 a_10805_n2997# a_10904_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1966 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1967 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1968 VDD sky130_fd_sc_hd__clkinv_1_4/Y sky130_fd_sc_hd__nand2_4_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1969 a_3266_n11933# a_3010_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1970 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1971 a_690_n13021# a_434_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X1972 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1973 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1974 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1975 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1976 VDD sky130_fd_sc_hd__clkinv_4_4/Y a_13765_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1977 VSS a_8588_n1079# a_8328_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X1978 VSS a_7130_n5405# a_7237_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X1979 VDD a_9706_n509# a_9813_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1980 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1981 a_501_n5797# a_600_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1982 a_1789_n12325# a_1888_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1983 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1984 a_8229_n5797# a_8328_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1985 a_4365_n13413# a_4464_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1986 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_9450_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1987 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_5949_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1988 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_7237_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X1989 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1990 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1991 VDD a_8418_n13021# a_8525_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1992 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1993 a_5842_n4317# a_5586_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X1994 VDD a_7300_n12503# a_7040_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X1995 a_3077_n12325# a_3176_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X1996 a_2148_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_10/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1997 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_6874_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1998 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_0/A a_n860_n509# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1999 sky130_fd_sc_hd__clkdlybuf4s50_1_157/A a_11101_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2000 a_9876_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2001 a_7300_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2002 VSS a_4554_n11933# a_4661_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2003 VDD a_11164_n10871# a_10904_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2004 VDD a_1978_n10301# a_2085_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2005 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2006 VSS a_860_n1079# a_600_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2007 VSS a_9706_n4317# a_9813_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2008 VDD a_9876_n10871# a_9616_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2009 VDD a_8418_n509# a_8525_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2010 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2011 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2012 a_10805_n1909# a_10904_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2013 VDD a_8418_n8125# a_8525_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2014 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2015 VSS a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2016 VSS a_690_n11933# a_797_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2017 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2018 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2019 a_860_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2020 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2021 a_5842_n10301# a_5586_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2022 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2023 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2024 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2025 a_3077_n2997# a_3176_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2026 a_860_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2027 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2028 a_4724_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2029 VSS a_4724_n12503# a_4464_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2030 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A a_5949_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2031 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_8525_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2032 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2033 VDD sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2034 a_8229_n4709# a_8328_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2035 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_434_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2036 VDD sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2037 VSS a_7300_n1079# a_7040_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2038 VDD a_6658_n7363# a_6665_n7459# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X2039 VSS sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_7/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2040 VSS a_3436_n11415# a_3176_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2041 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8162_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2042 VSS a_860_n12503# a_600_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2043 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2044 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_797_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2045 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_2085_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2046 a_7300_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2047 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2048 a_10805_n3621# a_10904_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2049 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2050 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_114/A a_1722_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2051 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A a_5949_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2052 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2053 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2054 B a_13765_n1053# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2055 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2056 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__nand2_1_4/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2057 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_2729_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2058 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2059 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2060 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2061 VSS a_3077_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2062 a_6012_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2063 VDD a_1789_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2064 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_4661_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2065 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2066 VDD a_13765_n9757# p2d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2067 VSS a_6012_n1079# a_5752_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2068 VSS a_4554_n4317# a_4661_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2069 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2070 VDD a_1789_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2071 VDD sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 a_3077_n1909# a_3176_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2073 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2074 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2075 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2076 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2077 a_3077_n9525# a_3176_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2078 a_4765_n7542# sky130_fd_sc_hd__dfxbp_1_0/Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X2079 a_8229_n9525# a_8328_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2080 sky130_fd_sc_hd__clkdlybuf4s50_1_45/A a_797_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2081 a_4554_n11933# a_4298_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2082 VDD a_8229_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2083 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2084 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2085 a_4765_n7215# sky130_fd_sc_hd__dfxbp_1_0/Q VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2086 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2087 a_6012_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2088 a_10805_n8437# a_10904_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2089 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2090 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2091 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2092 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2093 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2094 a_690_n11933# a_434_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2095 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2096 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8162_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2097 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2098 a_9876_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2099 VSS a_3077_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2100 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_8162_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2101 VSS a_10805_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2102 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2103 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2104 VDD a_7300_n5975# a_7040_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2105 a_6593_n7215# a_6101_n7254# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X2106 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2107 a_4623_n7349# Ad_b a_4765_n7542# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X2108 a_690_n5405# a_434_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2109 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2110 a_8418_n6493# a_8162_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2111 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2112 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2113 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2114 a_5653_n11237# a_5752_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2115 VDD a_9876_n5975# a_9616_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2116 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2117 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2118 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2119 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2120 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2121 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2122 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10738_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2123 a_3436_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2124 VSS a_5842_n2685# a_5949_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2125 VSS a_1789_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2126 a_5653_n10613# a_5752_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2127 VDD sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2128 VDD sky130_fd_sc_hd__clkinv_1_6/Y sky130_fd_sc_hd__nand2_4_2/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2129 VDD a_3077_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2130 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2131 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2132 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2133 a_860_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2134 VDD a_10805_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2135 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2136 VSS a_8418_n2685# a_8525_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2137 VDD a_8229_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2138 a_10994_n4317# a_10738_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2139 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2140 VSS a_9706_n9213# a_9813_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2141 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2142 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2143 a_690_n2685# a_434_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2144 VDD a_10994_n5405# a_11101_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2145 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2146 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2147 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2148 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2149 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2150 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2151 VDD sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2152 a_5082_n7542# Bd_b a_4623_n7349# VDD sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X2153 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2154 VSS sky130_fd_sc_hd__clkinv_1_3/Y a_2366_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2155 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2156 a_3436_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2157 a_6941_n4709# a_7040_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2158 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2159 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2160 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2161 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2162 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_4298_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2163 a_10738_n509# sky130_fd_sc_hd__nand2_4_0/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2164 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3010_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2165 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2166 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/A a_10738_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2167 VSS a_5052_n7283# a_4986_n7215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2168 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2169 a_8588_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2170 VDD a_4724_n5975# a_4464_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2171 VSS a_10994_n11933# a_11101_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2172 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_161/A a_4298_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2173 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2174 VSS a_9706_n11933# a_9813_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2175 VSS sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2176 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2177 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2178 VDD a_6012_n3255# a_5752_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2179 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11101_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2180 a_9706_n5405# a_9450_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2181 VDD a_n428_n12503# a_n688_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2182 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5586_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2183 VDD a_1978_n4317# a_2085_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2184 a_7130_n8125# a_6874_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2185 VDD a_10994_n2685# a_11101_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2186 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A a_4661_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2187 VDD a_8229_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2188 a_4986_n7215# Ad_b a_4623_n7349# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X2189 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2190 VDD a_8588_n3255# a_8328_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2191 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2192 VSS a_11164_n12503# a_10904_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2193 VSS a_4554_n9213# a_4661_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2194 VSS a_3266_n2685# a_3373_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2195 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2196 a_8229_n13413# a_8328_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2197 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2198 a_8229_n8437# a_8328_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2199 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2200 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2201 VSS a_9876_n12503# a_9616_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2202 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2203 a_3436_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2204 VSS a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2205 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2206 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/A a_3010_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2207 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2208 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2209 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2210 VSS a_8588_n11415# a_8328_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2211 VDD a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2212 a_10805_n821# a_10904_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2213 VDD a_4365_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2214 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2215 a_5842_n1597# a_5586_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2216 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2217 a_7130_n14109# a_6874_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2218 sky130_fd_sc_hd__nand2_4_1/B a_9813_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2219 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2220 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2221 VDD sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2222 a_9706_n2685# a_9450_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2223 VSS a_8229_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2224 VDD a_860_n4887# a_600_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2225 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2226 VDD a_6012_n2167# a_5752_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2227 VDD sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2228 a_4365_n4709# a_4464_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2229 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2230 a_5842_n13021# a_5586_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2231 a_9706_n10301# a_9450_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2232 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_1722_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2233 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2234 VSS a_8418_n6493# a_8525_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2235 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2236 VDD a_7130_n5405# a_7237_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2237 VDD a_8588_n2167# a_8328_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2238 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2239 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2240 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2241 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2242 a_8229_n12325# a_8328_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2243 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2244 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2245 VDD a_3436_n3255# a_3176_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2246 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2247 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2248 a_3266_n1597# a_3010_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2249 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2250 a_6616_n7581# a_6101_n7254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2251 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2252 VDD a_5653_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2253 a_8588_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2254 a_6101_n7254# a_6373_n7349# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2255 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2256 VSS a_6012_n3799# a_5752_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2257 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8162_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2258 VDD a_8229_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2259 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2260 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2261 VSS a_9517_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2262 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2263 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2264 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2265 VDD a_3077_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2266 VDD a_2622_n14109# a_2729_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2267 VDD a_3077_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2268 a_3436_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2269 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_7237_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2270 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2271 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2272 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2273 VSS a_8588_n3799# a_8328_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2274 VDD a_7130_n2685# a_7237_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2275 VSS a_8229_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2276 a_11164_n13591# sky130_fd_sc_hd__clkinv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2277 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3010_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2278 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_8525_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2279 VSS sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__clkinv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2280 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2281 a_10994_n9213# a_10738_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2282 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2283 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2284 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2285 VDD a_5052_n7283# a_5082_n7542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 VDD a_6012_n10871# a_5752_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2287 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2288 a_13765_n2141# sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2289 VSS a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2290 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2291 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8162_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2292 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2293 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2294 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2295 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9450_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2296 sky130_fd_sc_hd__nand2_4_3/B a_9813_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2297 a_1789_n4709# a_1888_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2298 VDD a_3436_n2167# a_3176_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2299 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2300 VSS sky130_fd_sc_hd__nand2_4_3/B a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2301 a_n1738_n6671# a_n2436_n7037# a_n1995_n6925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2302 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2303 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2304 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2305 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2306 VDD a_9517_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2307 VSS a_6012_n8695# a_5752_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2308 a_8418_n4317# a_8162_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2309 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/X a_8162_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2310 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2311 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2312 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2313 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2314 a_5653_n2997# a_5752_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2315 VDD a_8229_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2316 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2317 VDD sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2318 VDD a_11164_n3799# a_10904_n3799# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2319 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2320 a_11164_n13591# sky130_fd_sc_hd__clkinv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2321 VSS a_8588_n8695# a_8328_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2322 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2323 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2324 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2325 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2326 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A a_8525_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2327 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2328 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_2085_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2329 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2330 VSS a_3436_n3799# a_3176_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2331 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2332 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2333 VDD a_5653_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2334 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_8162_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2335 VSS a_8229_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2336 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2337 a_9876_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2338 VDD a_13765_n1053# B VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2339 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2340 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2341 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2342 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2343 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_4661_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2344 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2345 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_9813_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2346 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2347 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_8525_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2348 a_3266_n5405# a_3010_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2349 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2350 a_13765_n10301# sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2351 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2352 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2353 a_3077_n821# a_3176_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2354 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2355 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2356 a_9517_n3621# a_9616_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2357 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2358 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2359 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2360 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2361 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6874_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2362 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2363 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2364 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2365 a_5653_n1909# a_5752_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2366 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2367 a_6658_n7363# p2 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2368 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2369 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2370 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2371 VSS a_13765_n2685# Bd_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2372 a_5653_n9525# a_5752_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2373 sky130_fd_sc_hd__clkdlybuf4s50_1_58/A a_11101_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2374 VSS a_3436_n8695# a_3176_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2375 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2376 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2377 VDD a_n1738_n6671# a_n1570_n6769# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2378 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2379 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2380 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2381 a_8588_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2382 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2383 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2384 a_3077_n13413# a_3176_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2385 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2386 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2387 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2388 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2389 VSS sky130_fd_sc_hd__nand2_4_0/B a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2390 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2391 VSS sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2392 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2393 VSS a_11164_n1079# a_10904_n1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2394 VSS a_5653_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2395 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2396 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2397 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2398 VSS a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2399 VSS a_13765_n9757# p2d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2400 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2401 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2402 VDD a_1978_n1597# a_2085_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2403 VDD a_13765_n2685# Bd_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2404 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2405 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2406 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2407 VSS sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2408 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2409 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2410 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2411 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2412 VDD a_4724_n13591# a_4464_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2413 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2414 a_7130_n9213# a_6874_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2415 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2416 a_8229_n5797# a_8328_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2417 VDD a_10805_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2418 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2419 a_4554_n10301# a_4298_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2420 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2421 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2422 a_4623_n7349# Bd_b a_4765_n7215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2423 VSS a_6101_n7254# sky130_fd_sc_hd__dfxbp_1_0/Q VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2424 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2425 a_1978_n13021# a_1722_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2426 VDD a_860_n13591# a_600_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2427 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2428 VDD a_9706_n4317# a_9813_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2429 a_3077_n12325# a_3176_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2430 VSS a_7130_n509# a_7237_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2431 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2432 a_690_n10301# a_434_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2433 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2434 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2435 a_10805_n4709# a_10904_n4887# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2436 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2437 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2438 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2439 VDD a_9517_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2440 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2441 a_9706_n509# a_9450_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2442 VDD a_501_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2443 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2444 a_8418_n9213# a_8162_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2445 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2446 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2447 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_102/A a_8162_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2448 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2449 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2450 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2451 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2452 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2453 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4298_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2454 a_1789_n13413# a_1888_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2455 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2456 VSS a_5842_n11933# a_5949_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2457 a_5653_n11237# a_5752_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2458 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2459 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_6874_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2460 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2461 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2462 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2463 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A a_7237_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2464 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2465 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5586_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2466 VDD a_4724_n12503# a_4464_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2467 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2468 VSS a_3077_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2469 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2470 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2471 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2472 VSS a_7300_n13591# a_7040_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2473 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_797_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2474 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/A a_9450_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2475 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2476 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2477 a_7130_n10301# a_6874_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2478 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2479 a_8418_n509# a_8162_n509# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2480 VDD a_860_n12503# a_600_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2481 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/A a_13765_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2482 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2483 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2484 VSS a_13765_n2141# Bd VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2485 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_434_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2486 a_2622_n8125# a_2366_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2487 VSS a_6012_n12503# a_5752_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2488 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_2085_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2489 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_10738_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2490 VDD a_690_n9213# a_797_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2491 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2492 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2493 VDD a_4554_n4317# a_4661_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2494 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2495 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2496 a_4554_n9213# a_4298_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2497 sky130_fd_sc_hd__clkdlybuf4s50_1_77/A a_11101_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2498 VDD a_6865_n7304# a_6794_n7203# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2499 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2500 VDD sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2501 VDD a_13765_n4317# Ad_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2502 VDD sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2503 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/A a_3010_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2504 a_9706_n14109# a_9450_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2505 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/A a_8162_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2506 VDD sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2507 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2508 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2509 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2510 VSS a_6006_n7607# sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2511 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2512 a_11164_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2513 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/A a_5586_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2514 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2515 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2516 VDD a_3077_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2517 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2518 a_n787_n1909# a_n688_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2519 VDD a_501_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2520 VDD a_6941_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2521 a_4724_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2522 a_8588_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2523 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2524 VSS a_2148_n3255# a_1888_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2525 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A a_2085_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2526 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/A a_10738_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2527 VSS a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2528 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2529 a_n787_n9525# a_n688_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2530 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2531 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/X a_434_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2532 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1722_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2533 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2534 VSS a_2622_n509# a_2729_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2535 VSS a_10805_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2536 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2537 VSS a_1978_n10301# a_2085_n10301# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2538 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A a_4661_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2539 VSS a_13765_n5949# A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2540 VDD a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2541 a_10805_n10613# a_10904_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2542 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_3373_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2543 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2544 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2545 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2546 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2547 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2548 a_9876_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2549 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2550 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2551 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2552 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2553 VSS a_4623_n7349# sky130_fd_sc_hd__mux2_1_0/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2554 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2555 VDD a_n428_n2167# a_n688_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2556 a_5842_n1597# a_5586_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2557 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2558 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_9813_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2559 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X a_11101_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2560 a_1978_n11933# a_1722_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2561 VDD a_5653_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2562 a_1978_n9213# a_1722_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2563 VDD a_13765_n10301# p2d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2564 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2565 VDD a_501_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2566 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2567 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2568 VSS a_2148_n2167# a_1888_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2569 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2570 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2571 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2572 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2573 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2574 VDD a_2148_n9783# a_1888_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2575 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2576 a_10994_n4317# a_10738_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2577 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2578 VSS sky130_fd_sc_hd__nand2_4_3/Y a_13765_n9757# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2579 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/A a_13765_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2580 VSS a_13765_n4861# Ad VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2581 a_6941_n11237# a_7040_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2582 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_7237_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2583 a_n428_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2584 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2585 a_6794_n7203# a_6665_n7459# a_6373_n7349# VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X2586 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2587 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2588 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2589 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2590 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2591 VSS a_501_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2592 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2366_n14109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2593 VDD a_11164_n13591# a_10904_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2594 a_6941_n10613# a_7040_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2595 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2596 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2597 VDD a_9876_n13591# a_9616_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2598 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2599 a_11164_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2600 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2601 VDD sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2602 a_9876_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2603 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X2604 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_2729_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2605 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2606 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2607 a_3266_n5405# a_3010_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2608 a_n1654_n6671# a_n2436_n7037# a_n1738_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2609 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2610 a_9706_n8125# a_9450_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2611 VSS sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2612 VDD a_13765_n4861# Ad VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2613 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2614 a_501_n2997# a_600_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2615 sky130_fd_sc_hd__clkdlybuf4s50_1_5/A sky130_fd_sc_hd__nand2_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2616 a_n428_n12503# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2617 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2618 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2619 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2620 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2621 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2622 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2623 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_2729_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2624 VDD a_2148_n11415# a_1888_n11415# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2625 a_5052_n7283# sky130_fd_sc_hd__dfxbp_1_0/Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2626 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2627 VDD a_501_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_50/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2628 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_2085_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2629 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2630 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2631 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2632 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2633 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2634 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2635 VDD a_11164_n12503# a_10904_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2636 VSS sky130_fd_sc_hd__clkinv_1_0/Y a_2366_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2637 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2638 a_6941_n5797# a_7040_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2639 a_5052_n7283# sky130_fd_sc_hd__dfxbp_1_0/Q VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X2640 VDD a_9876_n12503# a_9616_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2641 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/A a_434_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2642 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_4298_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2643 a_5842_n5405# a_5586_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2644 a_7130_n14109# a_6874_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2645 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A a_7237_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2646 VSS sky130_fd_sc_hd__nand2_4_0/Y a_13765_n2141# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2647 a_11164_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2648 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A a_4661_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2649 VSS a_2148_n10871# a_1888_n10871# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2650 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_9813_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2651 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A a_5949_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2652 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_160/A a_1722_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2653 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A a_8525_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2654 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2655 a_3266_n2685# a_3010_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2656 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_8162_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2657 a_5653_n821# a_5752_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2658 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2659 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2660 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2661 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2662 p2d a_13765_n9757# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2663 VDD a_9706_n1597# a_9813_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2664 VSS sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2665 VDD a_6012_n4887# a_5752_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2666 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2667 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A a_7237_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2668 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2669 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2670 a_501_n1909# a_600_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2671 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2672 VDD a_7130_n8125# a_7237_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2673 VDD a_8588_n4887# a_8328_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2674 a_6658_n7363# p2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2675 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2676 a_501_n9525# a_600_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2677 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2678 a_690_n2685# a_434_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2679 VSS sky130_fd_sc_hd__nand2_4_2/B a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2680 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2681 VDD a_13765_n13565# p1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2682 a_11164_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2683 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2684 a_n860_n13789# sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2685 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2686 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2687 a_5653_n821# a_5752_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2688 VSS a_13765_n4317# Ad_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2689 a_6941_n4709# a_7040_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2690 p2d_b a_13765_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2691 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2692 a_7300_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2693 a_7130_n13021# a_6874_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2694 a_6012_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2695 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2696 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2697 a_501_n11237# a_600_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2698 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A a_2085_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2699 a_8418_n13021# a_8162_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2700 VSS a_8418_n8125# a_8525_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2701 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2702 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2703 VSS a_501_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2704 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2705 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2706 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_2729_n8125# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2707 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2708 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2709 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2710 VSS a_860_n5975# a_600_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2711 a_2622_n6493# a_2366_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2712 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2713 a_4365_n5797# a_4464_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2714 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2715 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_60/A a_1722_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2716 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_3373_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2717 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A a_4661_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2718 VDD a_4554_n1597# a_4661_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2719 a_501_n10613# a_600_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2720 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2721 VSS a_10994_n2685# a_11101_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2722 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2723 a_4365_n821# a_4464_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2724 a_n428_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2725 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2726 a_11164_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_58/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2727 a_8229_n13413# a_8328_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2728 VDD a_13765_n2141# Bd VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2729 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2730 VDD a_3436_n4887# a_3176_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2731 a_10805_n12325# a_10904_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2732 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2733 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2734 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2735 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2736 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2737 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2738 VDD sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2739 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2740 a_6941_n9525# a_7040_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2741 a_7300_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2742 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2743 a_8418_n4317# a_8162_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2744 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2745 VDD a_10805_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2746 VSS a_6941_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2747 VSS sky130_fd_sc_hd__clkinv_4_10/Y a_13765_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2748 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2749 VSS a_n787_n4709# sky130_fd_sc_hd__nand2_1_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2750 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/A a_2366_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2751 VDD a_1978_n13021# a_2085_n13021# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2752 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2753 a_860_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2754 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2755 a_3077_n821# a_3176_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2756 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11101_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2757 VSS a_13765_n13021# p1_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2758 VDD a_13765_n8669# p2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2759 a_9706_n2685# a_9450_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2760 VSS a_7300_n3255# a_7040_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2761 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2762 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2763 VSS a_1978_n1597# a_2085_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2764 VSS a_860_n4887# a_600_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2765 VSS a_5653_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2766 a_4365_n4709# a_4464_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2767 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2768 Bd a_13765_n2141# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2769 a_860_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2770 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2771 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2772 a_9706_n10301# a_9450_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2773 B_b a_13765_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2774 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_81/A a_4298_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2775 VDD a_3436_n10871# a_3176_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2776 VSS a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2777 VDD a_9517_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2778 VSS a_9876_n3255# a_9616_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2779 VDD a_11164_n3255# a_10904_n3255# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2780 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2781 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2782 a_7300_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2783 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2784 a_7130_n6493# a_6874_n6493# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2785 a_1789_n5797# a_1888_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2786 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2787 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_100/A a_2366_n14109# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2788 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2789 a_3077_n3621# a_3176_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2790 VDD a_6941_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2791 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2792 VDD a_n787_n4709# sky130_fd_sc_hd__nand2_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2793 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X a_11101_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2794 a_2148_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_11/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2795 a_11164_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_31/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2796 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2797 VDD a_5653_n12325# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2798 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2799 VSS a_7300_n2167# a_7040_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2800 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2801 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2802 a_860_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2803 VSS a_860_n9783# a_600_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2804 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2805 a_10994_n1597# a_10738_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2806 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A a_2729_n14109# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2807 a_4365_n9525# a_4464_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2808 B_b a_13765_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2809 a_9517_n2997# a_9616_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2810 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_5586_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2811 VDD a_7300_n9783# a_7040_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2812 a_4724_n2167# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2813 VSS a_7130_n2685# a_7237_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2814 VSS a_13765_n5405# A_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2815 VDD a_4365_n11237# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2816 VSS a_9876_n2167# a_9616_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2817 a_7300_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2818 VDD a_4365_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2819 VDD a_11164_n2167# a_10904_n2167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2820 VSS a_7130_n13021# a_7237_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2821 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2822 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2823 VSS a_4724_n3255# a_4464_n3255# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2824 VDD a_9876_n9783# a_9616_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2825 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2826 VDD sky130_fd_sc_hd__clkinv_1_3/Y a_2366_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2827 VDD sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2828 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2829 a_1789_n4709# a_1888_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2830 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2831 p2 a_13765_n8669# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2832 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_121/A a_10738_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2833 a_8418_n11933# a_8162_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2834 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_181/A a_4298_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2835 VSS sky130_fd_sc_hd__clkinv_1_5/A a_7212_n7203# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2836 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2837 a_3436_n8695# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2838 VSS a_1789_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_41/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2839 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_79/A a_1722_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2840 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2841 VDD a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2842 VDD sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2843 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2844 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2845 a_13765_n1053# sky130_fd_sc_hd__clkinv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2846 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_7237_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2847 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_8525_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2848 a_9706_n6493# a_9450_n6493# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2849 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X a_3373_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2850 VSS sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_9813_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2852 VSS a_1978_n5405# a_2085_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2853 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2854 VSS a_11164_n3799# a_10904_n3799# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2855 a_9517_n1909# a_9616_n2167# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2856 VDD a_2148_n1079# a_1888_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2857 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2858 VSS a_13765_n12477# p1d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2859 VSS sky130_fd_sc_hd__clkinv_1_3/A a_13765_n8669# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2860 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2861 a_9517_n821# a_9616_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2862 a_6941_n8437# a_7040_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2863 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2864 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2865 a_9517_n11237# a_9616_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2866 VSS a_4724_n2167# a_4464_n2167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2867 a_2148_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2868 sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2869 a_1789_n9525# a_1888_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2870 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2871 VDD a_4724_n9783# a_4464_n9783# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2872 VDD a_13765_n9213# p2_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2873 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2874 VSS a_4365_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_145/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2875 VDD a_3077_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2876 a_13765_n9213# sky130_fd_sc_hd__clkinv_4_10/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2877 VDD a_7130_n509# a_7237_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2878 a_4724_n3799# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2879 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/A a_9450_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2880 VDD a_6012_n13591# a_5752_n13591# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2881 a_9517_n10613# a_9616_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2882 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A a_7237_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2883 a_7300_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2884 a_9517_n3621# a_9616_n3799# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2885 VDD sky130_fd_sc_hd__clkinv_4_8/A a_13765_n12477# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2886 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2887 sky130_fd_sc_hd__dfxbp_1_1/D a_n1139_n6715# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2888 VSS a_4365_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2889 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2890 a_n2068_n6671# a_n2602_n7037# a_n2163_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X2891 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2892 a_8229_n821# a_8328_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2893 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2894 VSS a_8229_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2895 a_3266_n13021# a_3010_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2896 a_9706_n509# a_9450_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2897 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_2085_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2898 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2899 VDD a_13765_n12477# p1d VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2900 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2901 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2902 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_179/A a_1722_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2903 VSS a_11164_n8695# a_10904_n8695# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2904 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2905 VSS a_7130_n6493# a_7237_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2906 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2907 a_1978_n10301# a_1722_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2908 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2909 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2910 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_4661_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2911 a_5842_n5405# a_5586_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2912 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2913 sky130_fd_sc_hd__clkdlybuf4s50_1_89/A sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2914 a_3077_n13413# a_3176_n13591# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2915 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2916 a_6941_n11237# a_7040_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2917 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/A a_8162_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2918 a_10805_n5797# a_10904_n5975# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2919 VDD a_5842_n9213# a_5949_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2920 a_501_n821# a_600_n1079# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2921 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2922 a_9876_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X2923 a_8418_n509# a_8162_n509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2924 a_8588_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2925 VSS a_4554_n13021# a_4661_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2926 p2d_b a_13765_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2927 VDD a_860_n8695# a_600_n8695# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2928 a_6006_n7607# a_6101_n7254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X2929 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2930 VDD a_6012_n12503# a_5752_n12503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2931 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2932 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2933 a_4365_n8437# a_4464_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2934 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_139/A a_9450_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2935 a_9517_n8437# a_9616_n8695# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2936 a_9706_n14109# a_9450_n14109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2937 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2938 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2939 VSS a_3266_n11933# a_3373_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2940 sky130_fd_sc_hd__clkdlybuf4s50_1_18/A a_2085_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2941 a_2148_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_32/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2942 VSS a_690_n13021# a_797_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X2943 VSS a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2944 a_6012_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2945 VDD a_8418_n9213# a_8525_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2946 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2947 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2948 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2949 VDD a_8588_n10871# a_8328_n10871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2950 B a_13765_n1053# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2951 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2952 VDD a_1789_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X2953 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2954 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2955 VDD a_7130_n11933# a_7237_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2956 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2957 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A a_11101_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X2958 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2959 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2960 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A a_6874_n6493# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2961 VSS a_4724_n13591# a_4464_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2962 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2963 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A a_4661_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X2964 a_4724_n3255# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2965 VSS a_6865_n7304# a_6794_n7203# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2966 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_113/A a_434_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2967 a_4554_n10301# a_4298_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2968 a_7300_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X2969 a_5842_n2685# a_5586_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2970 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2971 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2972 VSS sky130_fd_sc_hd__clkinv_4_8/Y a_13765_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2973 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2974 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/A a_9450_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2975 a_501_n821# a_600_n1079# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2976 VSS a_4365_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2977 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2978 VSS a_5653_n8437# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2979 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2980 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_95/A a_8162_n6493# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X2981 VDD sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkinv_4_8/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2982 VSS a_3436_n12503# a_3176_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2983 VSS a_860_n13591# a_600_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2984 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2985 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2986 VSS a_13765_n11933# p1d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2987 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2988 a_690_n10301# a_434_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X2989 a_8418_n1597# a_8162_n1597# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X2990 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2991 a_10805_n4709# a_10904_n4887# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X2992 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2993 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2994 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2995 VDD a_2622_n509# a_2729_n509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X2996 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2997 VSS a_2148_n11415# a_1888_n11415# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X2998 VSS a_6941_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X2999 a_7130_n4317# a_6874_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3000 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3001 Bd_b a_13765_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3002 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3003 VDD a_1789_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3004 a_6012_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3005 a_9706_n13021# a_9450_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3006 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3007 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3008 a_6012_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3009 VDD a_n428_n4887# a_n688_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3010 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3011 p1d a_13765_n12477# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3012 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X3013 VDD a_1789_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_46/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3014 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3015 VDD a_3266_n9213# a_3373_n9213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3016 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3017 VDD sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3018 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3019 a_8588_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3020 a_1789_n8437# a_1888_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3021 VSS sky130_fd_sc_hd__clkinv_1_0/A sky130_fd_sc_hd__clkinv_1_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3022 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3023 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3024 VSS a_9706_n1597# a_9813_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3025 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3026 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3027 VSS a_5653_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3028 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_3373_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3029 Ad_b a_13765_n4317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3030 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3031 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3032 p2d a_13765_n9757# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3033 a_6012_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3034 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3035 a_10805_n9525# a_10904_n9783# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3036 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3037 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3038 Bd_b a_13765_n2685# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3039 a_3266_n11933# a_3010_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3040 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3041 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3042 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3043 VSS a_1789_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3044 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4298_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3045 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3046 sky130_fd_sc_hd__clkinv_1_5/A a_n1570_n6769# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3047 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/A a_6874_n8125# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3048 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3049 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3050 VDD a_10805_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3051 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3052 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3053 p1d a_13765_n12477# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3054 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3055 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3056 VSS a_10805_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3057 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X3058 a_6373_n7349# a_6658_n7363# a_6593_n7215# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3059 VSS a_4365_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_10/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3060 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3061 VSS a_690_n4317# a_797_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3062 VDD sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3063 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3064 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A a_9813_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3065 a_501_n11237# a_600_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3066 A a_13765_n5949# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3067 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3068 a_4554_n4317# a_4298_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3069 a_3436_n5975# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3070 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3071 VSS a_13765_n9213# p2_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3072 VDD a_9517_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_4/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3073 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3074 VDD a_4554_n11933# a_4661_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3075 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3076 a_10738_n8125# sky130_fd_sc_hd__nand2_4_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3077 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10738_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3078 a_4365_n11237# a_4464_n11415# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3079 VSS a_4554_n1597# a_4661_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3080 A a_13765_n5949# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3081 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3082 VDD a_690_n11933# a_797_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3083 VDD a_1789_n3621# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3084 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3085 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_19/A a_4298_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3086 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3087 VSS a_13765_n1597# B_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3088 a_860_n9783# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3089 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3090 VSS sky130_fd_sc_hd__clkinv_4_4/A a_13765_n5949# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3091 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A a_10738_n8125# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3092 VDD a_10805_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3093 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3094 VDD sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3095 a_4365_n10613# a_4464_n10871# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3096 a_8229_n2997# a_8328_n3255# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3097 a_13765_n11933# sky130_fd_sc_hd__clkinv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3098 a_10994_n11933# a_10738_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3099 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3100 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3101 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3102 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3103 a_n787_n12325# a_n688_n12503# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3104 VDD sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3105 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3106 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3107 Bd a_13765_n2141# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3108 Ad a_13765_n4861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3109 a_3436_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_106/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3110 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3111 VDD a_7300_n1079# a_7040_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3112 a_5653_n3621# a_5752_n3799# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3113 a_3436_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3114 a_6941_n5797# a_7040_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3115 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3116 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1722_n1597# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3117 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3118 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3119 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3120 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3121 VSS a_9706_n5405# a_9813_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3122 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/A a_10738_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3123 p1d_b a_13765_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3124 VSS a_10805_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3125 VSS a_10994_n13021# a_11101_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3126 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3127 VSS sky130_fd_sc_hd__clkinv_1_0/A a_13765_n1053# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3128 VDD a_9876_n1079# a_9616_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3129 VSS a_9706_n13021# a_9813_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3130 VSS a_8229_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3131 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A a_2085_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3132 VDD a_13765_n1597# B_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3133 a_1978_n4317# a_1722_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3134 VDD a_13765_n11933# p1d_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3135 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3136 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3137 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/A a_3010_n10301# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3138 sky130_fd_sc_hd__clkdlybuf4s50_1_77/A a_11101_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3139 VSS a_8418_n11933# a_8525_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3140 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_117/A a_5586_n13021# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3141 a_7130_n9213# a_6874_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3142 VSS sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3143 VDD a_1978_n5405# a_2085_n5405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3144 VDD a_6941_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_7/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3145 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3146 a_8229_n1909# a_8328_n2167# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3147 VSS a_9517_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3148 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3149 A_b a_13765_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3150 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_135/A a_4298_n11933# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3151 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3152 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3153 VSS a_11164_n13591# a_10904_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3154 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3155 a_8229_n9525# a_8328_n9783# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3156 Ad a_13765_n4861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3157 VSS a_9876_n13591# a_9616_n13591# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3158 VSS sky130_fd_sc_hd__nand2_4_1/B a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3159 a_10805_n13413# a_10904_n13591# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3160 a_3436_n4887# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3161 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_43/A a_1722_n1597# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3162 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3163 VSS a_1789_n2997# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3164 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3165 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3166 VSS a_8588_n12503# a_8328_n12503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3167 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3168 VSS a_13765_n10301# p2d_b VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3169 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X3170 VSS sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkdlybuf4s50_1_89/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X3171 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A a_4661_n11933# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3172 VDD a_501_n10613# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3173 p1 a_13765_n13565# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3174 a_10805_n8437# a_10904_n8695# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3175 a_10994_n1597# a_10738_n1597# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3176 p1_b a_13765_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3177 sky130_fd_sc_hd__clkinv_4_8/A sky130_fd_sc_hd__nand2_4_2/A a_10738_n13789# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3178 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3179 VSS a_6012_n5975# a_5752_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3180 A_b a_13765_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3181 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3182 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3183 VDD sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3184 VSS a_4554_n5405# a_4661_n5405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3185 VSS a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3186 VDD a_1978_n2685# a_2085_n2685# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3187 VDD a_860_n5975# a_600_n5975# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3188 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3189 VDD a_4724_n1079# a_4464_n1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3190 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A a_9813_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3191 VDD sky130_fd_sc_hd__clkinv_4_3/A a_13765_n4861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3192 VDD sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__clkinv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3193 a_4365_n5797# a_4464_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3194 VSS a_13765_n8669# p2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3195 VSS a_8588_n5975# a_8328_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3196 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3197 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3198 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3199 VSS a_10805_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3200 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3201 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3202 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3203 a_4554_n13021# a_4298_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3204 a_8418_n10301# a_8162_n10301# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3205 VSS a_5653_n5797# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3206 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3207 a_2622_n8125# a_2366_n8125# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3208 a_10805_n12325# a_10904_n12503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3209 VSS a_690_n9213# a_797_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X3210 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3211 a_3266_n2685# a_3010_n2685# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3212 a_690_n13021# a_434_n13021# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3213 p1 a_13765_n13565# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3214 a_4554_n9213# a_4298_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3215 p2_b a_13765_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3216 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3217 VSS a_6941_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3218 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3219 a_10738_n13789# sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_4_8/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3220 a_5653_n10613# a_5752_n10871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3221 VSS a_6012_n4887# a_5752_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3222 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3223 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3224 VSS a_9517_n1909# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3225 VDD a_8229_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3226 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A a_3373_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3227 a_13765_n4317# sky130_fd_sc_hd__clkinv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3228 VDD a_13765_n5949# A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3229 Ad_b a_13765_n4317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3230 VDD a_3077_n9525# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3231 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3232 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3233 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A a_7237_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3234 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3235 VSS a_8588_n4887# a_8328_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3236 a_13765_n5949# sky130_fd_sc_hd__clkinv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3237 a_9517_n11237# a_9616_n11415# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u w=650000u l=500000u
X3238 a_9876_n1079# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3239 VSS a_8229_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3240 a_8588_n10871# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3241 sky130_fd_sc_hd__clkinv_4_4/A sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3242 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3243 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3244 sky130_fd_sc_hd__clkdlybuf4s50_1_195/A sky130_fd_sc_hd__nand2_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3245 p2_b a_13765_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3246 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3247 VSS a_3436_n5975# a_3176_n5975# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3248 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3249 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3250 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A a_9813_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3251 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A a_8525_n10301# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
X3252 VSS a_5653_n4709# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3253 a_9876_n13591# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3254 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_29/A a_8162_n2685# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3255 VDD a_n1995_n6925# a_n2068_n6671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3256 VSS sky130_fd_sc_hd__clkdlybuf4s50_1_185/A a_9450_n9213# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X3257 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A a_9813_n9213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3258 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3259 a_1789_n5797# a_1888_n5975# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3260 a_7212_n7203# a_6665_n7459# a_6865_n7304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3261 VSS a_13765_n13565# p1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3262 VDD a_10994_n11933# a_11101_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3263 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3264 VSS sky130_fd_sc_hd__clkinv_4_3/Y a_13765_n4317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3265 a_13765_n12477# sky130_fd_sc_hd__clkinv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3266 VDD a_9706_n11933# a_9813_n11933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3267 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3268 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X3269 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3270 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3271 a_3077_n2997# a_3176_n3255# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=0p ps=0u w=820000u l=500000u
X3272 a_10994_n5405# a_10738_n5405# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3273 sky130_fd_sc_hd__clkinv_4_3/A sky130_fd_sc_hd__nand2_4_1/A a_10738_n6173# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3274 a_2148_n11415# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VSS sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X3275 VSS a_6012_n9783# a_5752_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3276 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3277 VSS a_501_n821# sky130_fd_sc_hd__clkdlybuf4s50_1_42/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.491e+11p ps=1.55e+06u w=420000u l=150000u
X3278 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3279 p1d_b a_13765_n11933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3280 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X3281 VDD a_8229_n13413# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.55e+11p ps=2.71e+06u w=1e+06u l=150000u
X3282 VDD a_11164_n4887# a_10904_n4887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3283 a_1978_n9213# a_1722_n9213# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X3284 VSS a_13765_n1053# B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3285 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3286 a_13765_n4861# sky130_fd_sc_hd__clkinv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3287 VSS a_8588_n9783# a_8328_n9783# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3288 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A a_10738_n509# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3289 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3290 a_10738_n6173# sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3291 p1_b a_13765_n13021# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3292 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3293 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X3294 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A a_2085_n5405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X3295 a_13765_n8669# sky130_fd_sc_hd__clkinv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3296 VSS a_3436_n4887# a_3176_n4887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=500000u
X3297 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X3298 p2 a_13765_n8669# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3299 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X3300 VDD a_13765_n5405# A_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

