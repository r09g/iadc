magic
tech sky130A
magscale 1 2
timestamp 1654716000
<< nwell >>
rect -777 -240 777 240
<< pmoslvt >>
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
<< pdiff >>
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
<< pdiffc >>
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
<< poly >>
rect -665 221 -581 237
rect -665 204 -649 221
rect -683 187 -649 204
rect -597 204 -581 221
rect -487 221 -403 237
rect -487 204 -471 221
rect -597 187 -563 204
rect -683 140 -563 187
rect -505 187 -471 204
rect -419 204 -403 221
rect -309 221 -225 237
rect -309 204 -293 221
rect -419 187 -385 204
rect -505 140 -385 187
rect -327 187 -293 204
rect -241 204 -225 221
rect -131 221 -47 237
rect -131 204 -115 221
rect -241 187 -207 204
rect -327 140 -207 187
rect -149 187 -115 204
rect -63 204 -47 221
rect 47 221 131 237
rect 47 204 63 221
rect -63 187 -29 204
rect -149 140 -29 187
rect 29 187 63 204
rect 115 204 131 221
rect 225 221 309 237
rect 225 204 241 221
rect 115 187 149 204
rect 29 140 149 187
rect 207 187 241 204
rect 293 204 309 221
rect 403 221 487 237
rect 403 204 419 221
rect 293 187 327 204
rect 207 140 327 187
rect 385 187 419 204
rect 471 204 487 221
rect 581 221 665 237
rect 581 204 597 221
rect 471 187 505 204
rect 385 140 505 187
rect 563 187 597 204
rect 649 204 665 221
rect 649 187 683 204
rect 563 140 683 187
rect -683 -187 -563 -140
rect -683 -204 -649 -187
rect -665 -221 -649 -204
rect -597 -204 -563 -187
rect -505 -187 -385 -140
rect -505 -204 -471 -187
rect -597 -221 -581 -204
rect -665 -237 -581 -221
rect -487 -221 -471 -204
rect -419 -204 -385 -187
rect -327 -187 -207 -140
rect -327 -204 -293 -187
rect -419 -221 -403 -204
rect -487 -237 -403 -221
rect -309 -221 -293 -204
rect -241 -204 -207 -187
rect -149 -187 -29 -140
rect -149 -204 -115 -187
rect -241 -221 -225 -204
rect -309 -237 -225 -221
rect -131 -221 -115 -204
rect -63 -204 -29 -187
rect 29 -187 149 -140
rect 29 -204 63 -187
rect -63 -221 -47 -204
rect -131 -237 -47 -221
rect 47 -221 63 -204
rect 115 -204 149 -187
rect 207 -187 327 -140
rect 207 -204 241 -187
rect 115 -221 131 -204
rect 47 -237 131 -221
rect 225 -221 241 -204
rect 293 -204 327 -187
rect 385 -187 505 -140
rect 385 -204 419 -187
rect 293 -221 309 -204
rect 225 -237 309 -221
rect 403 -221 419 -204
rect 471 -204 505 -187
rect 563 -187 683 -140
rect 563 -204 597 -187
rect 471 -221 487 -204
rect 403 -237 487 -221
rect 581 -221 597 -204
rect 649 -204 683 -187
rect 649 -221 665 -204
rect 581 -237 665 -221
<< polycont >>
rect -649 187 -597 221
rect -471 187 -419 221
rect -293 187 -241 221
rect -115 187 -63 221
rect 63 187 115 221
rect 241 187 293 221
rect 419 187 471 221
rect 597 187 649 221
rect -649 -221 -597 -187
rect -471 -221 -419 -187
rect -293 -221 -241 -187
rect -115 -221 -63 -187
rect 63 -221 115 -187
rect 241 -221 293 -187
rect 419 -221 471 -187
rect 597 -221 649 -187
<< locali >>
rect -729 187 -649 221
rect -597 187 -581 221
rect -487 187 -471 221
rect -419 187 -403 221
rect -309 187 -293 221
rect -241 187 -225 221
rect -131 187 -115 221
rect -63 187 -47 221
rect 47 187 63 221
rect 115 187 131 221
rect 225 187 241 221
rect 293 187 309 221
rect 403 187 419 221
rect 471 187 487 221
rect 581 187 597 221
rect 649 187 729 221
rect -729 128 -695 187
rect -729 -187 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 187
rect 695 -187 729 -128
rect -729 -221 -649 -187
rect -597 -221 -581 -187
rect -487 -221 -471 -187
rect -419 -221 -403 -187
rect -309 -221 -293 -187
rect -241 -221 -225 -187
rect -131 -221 -115 -187
rect -63 -221 -47 -187
rect 47 -221 63 -187
rect 115 -221 131 -187
rect 225 -221 241 -187
rect 293 -221 309 -187
rect 403 -221 419 -187
rect 471 -221 487 -187
rect 581 -221 597 -187
rect 649 -221 729 -187
<< viali >>
rect -471 187 -419 221
rect -293 187 -241 221
rect -115 187 -63 221
rect 63 187 115 221
rect 241 187 293 221
rect 419 187 471 221
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect -471 -221 -419 -187
rect -293 -221 -241 -187
rect -115 -221 -63 -187
rect 63 -221 115 -187
rect 241 -221 293 -187
rect 419 -221 471 -187
<< metal1 >>
rect -483 221 -407 227
rect -483 187 -471 221
rect -419 187 -407 221
rect -483 181 -407 187
rect -305 221 -229 227
rect -305 187 -293 221
rect -241 187 -229 221
rect -305 181 -229 187
rect -127 221 -51 227
rect -127 187 -115 221
rect -63 187 -51 221
rect -127 181 -51 187
rect 51 221 127 227
rect 51 187 63 221
rect 115 187 127 221
rect 51 181 127 187
rect 229 221 305 227
rect 229 187 241 221
rect 293 187 305 221
rect 229 181 305 187
rect 407 221 483 227
rect 407 187 419 221
rect 471 187 483 221
rect 407 181 483 187
rect -557 128 -511 140
rect -557 -128 -551 128
rect -517 -128 -511 128
rect -557 -140 -511 -128
rect -379 128 -333 140
rect -379 -128 -373 128
rect -339 -128 -333 128
rect -379 -140 -333 -128
rect -201 128 -155 140
rect -201 -128 -195 128
rect -161 -128 -155 128
rect -201 -140 -155 -128
rect -23 128 23 140
rect -23 -128 -17 128
rect 17 -128 23 128
rect -23 -140 23 -128
rect 155 128 201 140
rect 155 -128 161 128
rect 195 -128 201 128
rect 155 -140 201 -128
rect 333 128 379 140
rect 333 -128 339 128
rect 373 -128 379 128
rect 333 -140 379 -128
rect 511 128 557 140
rect 511 -128 517 128
rect 551 -128 557 128
rect 511 -140 557 -128
rect -483 -187 -407 -181
rect -483 -221 -471 -187
rect -419 -221 -407 -187
rect -483 -227 -407 -221
rect -305 -187 -229 -181
rect -305 -221 -293 -187
rect -241 -221 -229 -187
rect -305 -227 -229 -221
rect -127 -187 -51 -181
rect -127 -221 -115 -187
rect -63 -221 -51 -187
rect -127 -227 -51 -221
rect 51 -187 127 -181
rect 51 -221 63 -187
rect 115 -221 127 -187
rect 51 -227 127 -221
rect 229 -187 305 -181
rect 229 -221 241 -187
rect 293 -221 305 -187
rect 229 -227 305 -221
rect 407 -187 483 -181
rect 407 -221 419 -187
rect 471 -221 483 -187
rect 407 -227 483 -221
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 8 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
