magic
tech sky130A
magscale 1 2
timestamp 1654408082
<< error_p >>
rect -29 136 29 142
rect -29 102 -17 136
rect -29 96 29 102
rect -29 -102 29 -96
rect -29 -136 -17 -102
rect -29 -142 29 -136
<< pwell >>
rect -311 -274 311 274
<< nmos >>
rect -111 -64 -81 64
rect -15 -64 15 64
rect 81 -64 111 64
<< ndiff >>
rect -173 52 -111 64
rect -173 -52 -161 52
rect -127 -52 -111 52
rect -173 -64 -111 -52
rect -81 52 -15 64
rect -81 -52 -65 52
rect -31 -52 -15 52
rect -81 -64 -15 -52
rect 15 52 81 64
rect 15 -52 31 52
rect 65 -52 81 52
rect 15 -64 81 -52
rect 111 52 173 64
rect 111 -52 127 52
rect 161 -52 173 52
rect 111 -64 173 -52
<< ndiffc >>
rect -161 -52 -127 52
rect -65 -52 -31 52
rect 31 -52 65 52
rect 127 -52 161 52
<< psubdiff >>
rect -275 204 -179 238
rect 179 204 275 238
rect -275 142 -241 204
rect 241 142 275 204
rect -275 -204 -241 -142
rect 241 -204 275 -142
rect -275 -238 -179 -204
rect 179 -238 275 -204
<< psubdiffcont >>
rect -179 204 179 238
rect -275 -142 -241 142
rect 241 -142 275 142
rect -179 -238 179 -204
<< poly >>
rect -129 136 129 152
rect -129 102 -17 136
rect 17 102 129 136
rect -129 86 129 102
rect -111 64 -81 86
rect -15 64 15 86
rect 81 64 111 86
rect -111 -86 -81 -64
rect -15 -86 15 -64
rect 81 -86 111 -64
rect -129 -102 129 -86
rect -129 -136 -17 -102
rect 17 -136 129 -102
rect -129 -152 129 -136
<< polycont >>
rect -17 102 17 136
rect -17 -136 17 -102
<< locali >>
rect -275 204 -179 238
rect 179 204 275 238
rect -275 142 -241 204
rect 241 142 275 204
rect -33 102 -17 136
rect 17 102 33 136
rect -161 52 -127 68
rect -161 -68 -127 -52
rect -65 52 -31 68
rect -65 -68 -31 -52
rect 31 52 65 68
rect 31 -68 65 -52
rect 127 52 161 68
rect 127 -68 161 -52
rect -33 -136 -17 -102
rect 17 -136 33 -102
rect -275 -204 -241 -142
rect 241 -204 275 -142
rect -275 -238 -179 -204
rect 179 -238 275 -204
<< viali >>
rect -17 102 17 136
rect -161 -52 -127 52
rect -65 -52 -31 52
rect 31 -52 65 52
rect 127 -52 161 52
rect -17 -136 17 -102
<< metal1 >>
rect -29 136 29 142
rect -29 102 -17 136
rect 17 102 29 136
rect -29 96 29 102
rect -167 52 -121 64
rect -167 16 -161 52
rect -276 -18 -161 16
rect -167 -52 -161 -18
rect -127 16 -121 52
rect -71 52 -25 64
rect -71 16 -65 52
rect -127 -18 -65 16
rect -127 -52 -121 -18
rect -167 -64 -121 -52
rect -71 -52 -65 -18
rect -31 16 -25 52
rect 25 52 71 64
rect 25 16 31 52
rect -31 -18 31 16
rect -31 -52 -25 -18
rect -71 -64 -25 -52
rect 25 -52 31 -18
rect 65 16 71 52
rect 121 52 167 64
rect 121 16 127 52
rect 65 -18 127 16
rect 65 -52 71 -18
rect 25 -64 71 -52
rect 121 -52 127 -18
rect 161 16 167 52
rect 161 -18 276 16
rect 161 -52 167 -18
rect 121 -64 167 -52
rect -29 -102 29 -96
rect -29 -136 -17 -102
rect 17 -136 29 -102
rect -29 -142 29 -136
<< properties >>
string FIXED_BBOX -258 -222 258 222
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.65 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
