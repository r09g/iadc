magic
tech sky130A
magscale 1 2
timestamp 1655484843
<< nwell >>
rect 64797 61228 64861 61613
rect 65883 61347 65953 61600
rect 66973 61263 67044 61642
rect 74797 61228 74861 61613
rect 75883 61347 75953 61600
rect 76973 61263 77044 61642
rect 61973 41581 62325 42706
rect 62860 41583 63140 42706
rect 96488 41588 96840 42713
rect 97375 41590 97655 42713
<< pwell >>
rect 94938 47035 96094 47329
rect 133030 -495 141582 -360
rect 133030 -1812 141582 -1677
rect 66954 -6624 67089 -2026
rect 133030 -3459 141582 -3324
rect 133030 -4706 141582 -4571
rect 144962 -11687 153514 -11552
<< psubdiff >>
rect 60515 47140 60539 47278
rect 61454 47140 61478 47278
rect 95022 47131 95046 47253
rect 96035 47131 96059 47253
<< nsubdiff >>
rect 62063 42598 62235 42622
rect 62063 41635 62235 41659
rect 62908 42595 63080 42619
rect 62908 41632 63080 41656
rect 96578 42605 96750 42629
rect 96578 41642 96750 41666
rect 97423 42602 97595 42626
rect 97423 41639 97595 41663
<< psubdiffcont >>
rect 60539 47140 61454 47278
rect 95046 47131 96035 47253
<< nsubdiffcont >>
rect 62063 41659 62235 42598
rect 62908 41656 63080 42595
rect 96578 41666 96750 42605
rect 97423 41663 97595 42602
<< locali >>
rect 85076 63849 85353 63920
rect 85076 63757 85128 63849
rect 85318 63757 85353 63849
rect 86412 63858 86692 63906
rect 85076 63752 85353 63757
rect 86412 63764 86485 63858
rect 86629 63764 86692 63858
rect 102730 63849 103007 63920
rect 86412 63758 86692 63764
rect 102730 63757 102782 63849
rect 102972 63757 103007 63849
rect 104066 63858 104346 63906
rect 102730 63752 103007 63757
rect 104066 63764 104139 63858
rect 104283 63764 104346 63858
rect 104066 63758 104346 63764
rect 63373 62146 63774 62315
rect 63373 62033 63429 62146
rect 63542 62033 63774 62146
rect 63373 62018 63774 62033
rect 64216 62159 64511 62302
rect 64216 62045 64378 62159
rect 64491 62045 64511 62159
rect 64216 62024 64511 62045
rect 64710 62177 65111 62327
rect 64710 62064 64721 62177
rect 64834 62064 65111 62177
rect 64710 62030 65111 62064
rect 66095 62151 66496 62315
rect 66095 62038 66175 62151
rect 66288 62038 66496 62151
rect 67464 62151 67865 62318
rect 66095 62018 66496 62038
rect 67464 62038 67543 62151
rect 67656 62038 67865 62151
rect 73373 62146 73774 62315
rect 67464 62021 67865 62038
rect 73373 62033 73429 62146
rect 73542 62033 73774 62146
rect 73373 62018 73774 62033
rect 74216 62159 74511 62302
rect 74216 62045 74378 62159
rect 74491 62045 74511 62159
rect 74216 62024 74511 62045
rect 74710 62177 75111 62327
rect 74710 62064 74721 62177
rect 74834 62064 75111 62177
rect 74710 62030 75111 62064
rect 76095 62151 76496 62315
rect 76095 62038 76175 62151
rect 76288 62038 76496 62151
rect 77464 62151 77865 62318
rect 76095 62018 76496 62038
rect 77464 62038 77543 62151
rect 77656 62038 77865 62151
rect 77464 62021 77865 62038
rect 84916 59636 85101 59656
rect 84916 59523 84943 59636
rect 85056 59555 85101 59636
rect 102570 59636 102755 59656
rect 85056 59523 85065 59555
rect 84916 59497 85065 59523
rect 102570 59523 102597 59636
rect 102710 59555 102755 59636
rect 102710 59523 102719 59555
rect 102570 59497 102719 59523
rect 67919 59416 68307 59439
rect 63838 59351 64074 59385
rect 63838 59238 63937 59351
rect 64050 59238 64074 59351
rect 63838 59221 64074 59238
rect 65175 59363 65433 59393
rect 65175 59250 65298 59363
rect 65411 59250 65433 59363
rect 65175 59228 65433 59250
rect 66556 59381 66783 59410
rect 66556 59268 66660 59381
rect 66773 59268 66783 59381
rect 67919 59303 68044 59416
rect 68157 59303 68307 59416
rect 77919 59416 78307 59439
rect 67919 59284 68307 59303
rect 73838 59351 74074 59385
rect 66556 59239 66783 59268
rect 73838 59238 73937 59351
rect 74050 59238 74074 59351
rect 73838 59221 74074 59238
rect 75175 59363 75433 59393
rect 75175 59250 75298 59363
rect 75411 59250 75433 59363
rect 75175 59228 75433 59250
rect 76556 59381 76783 59410
rect 76556 59268 76660 59381
rect 76773 59268 76783 59381
rect 77919 59303 78044 59416
rect 78157 59303 78307 59416
rect 77919 59284 78307 59303
rect 76556 59239 76783 59268
rect 87203 59030 87482 59051
rect 87203 58917 87336 59030
rect 87449 58917 87482 59030
rect 87203 58893 87482 58917
rect 104857 59030 105136 59051
rect 104857 58917 104990 59030
rect 105103 58917 105136 59030
rect 104857 58893 105136 58917
rect 116643 52514 116993 52566
rect 116643 52386 116738 52514
rect 116866 52386 116993 52514
rect 46128 52282 46394 52310
rect 46128 51695 46153 52282
rect 46271 51695 46394 52282
rect 46128 51177 46394 51695
rect 47396 51852 47633 52332
rect 47396 51229 47493 51852
rect 47608 51229 47633 51852
rect 47396 51188 47633 51229
rect 48181 52230 48392 52319
rect 48181 51690 48197 52230
rect 48307 51690 48392 52230
rect 48181 51209 48392 51690
rect 49392 51907 49686 52344
rect 116643 52159 116993 52386
rect 120617 52467 121009 52490
rect 120617 52363 120662 52467
rect 120933 52363 121009 52467
rect 120617 52148 121009 52363
rect 49392 51249 49511 51907
rect 49654 51249 49686 51907
rect 115349 51725 115474 52126
rect 115385 51273 115474 51725
rect 49392 51203 49686 51249
rect 115349 51000 115474 51273
rect 117639 51778 117775 52133
rect 117639 51316 117729 51778
rect 117639 51031 117775 51316
rect 119407 51003 119486 52129
rect 121638 52123 121792 52134
rect 121638 51027 121709 52123
rect 121638 51008 121792 51027
rect 115930 50861 116239 50980
rect 119929 50958 120507 50993
rect 115930 50709 115989 50861
rect 116141 50709 116239 50861
rect 119930 50944 120507 50958
rect 119930 50832 119936 50944
rect 119929 50772 119936 50832
rect 120225 50772 120507 50944
rect 119929 50752 120507 50772
rect 115930 50690 116239 50709
rect 36194 49927 36347 50298
rect 37349 50285 37571 50315
rect 36194 49483 36202 49927
rect 36285 49483 36347 49927
rect 36194 49210 36347 49483
rect 37349 49792 37447 50285
rect 37567 49792 37571 50285
rect 37349 49202 37571 49792
rect 38141 49857 38346 50330
rect 39354 50313 39617 50339
rect 38141 49278 38144 49857
rect 38243 49278 38346 49857
rect 39354 49780 39493 50313
rect 39608 49780 39617 50313
rect 65977 49946 66106 50155
rect 66426 49946 66540 50155
rect 65977 49817 66540 49946
rect 67886 49987 67970 50150
rect 69607 50200 70000 50263
rect 68198 49987 68374 50150
rect 67886 49821 68374 49987
rect 69607 49968 69664 50200
rect 69892 49968 70000 50200
rect 69607 49821 70000 49968
rect 71399 50211 71833 50291
rect 71399 49979 71483 50211
rect 71711 49979 71833 50211
rect 71399 49821 71833 49979
rect 73190 50208 73708 50291
rect 73190 49976 73267 50208
rect 73495 49976 73708 50208
rect 73190 49825 73708 49976
rect 74980 50206 75427 50279
rect 74980 49974 75052 50206
rect 75280 49974 75427 50206
rect 74980 49824 75427 49974
rect 100501 49952 100630 50161
rect 100950 49952 101064 50161
rect 38141 49199 38346 49278
rect 39354 49174 39617 49780
rect 96364 49481 97874 49834
rect 100501 49823 101064 49952
rect 102410 49993 102494 50156
rect 104131 50206 104524 50269
rect 102722 49993 102898 50156
rect 102410 49827 102898 49993
rect 104131 49974 104188 50206
rect 104416 49974 104524 50206
rect 104131 49827 104524 49974
rect 105923 50217 106357 50297
rect 105923 49985 106007 50217
rect 106235 49985 106357 50217
rect 105923 49827 106357 49985
rect 107714 50214 108232 50297
rect 107714 49982 107791 50214
rect 108019 49982 108232 50214
rect 107714 49831 108232 49982
rect 109504 50212 109951 50285
rect 109504 49980 109576 50212
rect 109804 49980 109951 50212
rect 109504 49830 109951 49980
rect 96364 49447 96390 49481
rect 97826 49447 97874 49481
rect 96364 49432 97874 49447
rect 60309 47309 61584 47469
rect 60309 47109 60492 47309
rect 61496 47109 61584 47309
rect 60309 46941 61584 47109
rect 94850 47253 96125 47460
rect 94850 47131 95046 47253
rect 96035 47131 96125 47253
rect 94850 46932 96125 47131
rect 62063 42598 62235 42614
rect 62063 41643 62235 41659
rect 62908 42595 63080 42611
rect 84499 42609 84708 43024
rect 84499 42267 84505 42609
rect 84628 42267 84708 42609
rect 84499 41849 84708 42267
rect 86528 42646 86708 43021
rect 86528 42262 86529 42646
rect 86618 42262 86708 42646
rect 86528 41878 86708 42262
rect 96578 42605 96750 42621
rect 62908 41640 63080 41656
rect 96578 41650 96750 41666
rect 97423 42602 97595 42618
rect 97423 41647 97595 41663
rect 79901 40739 80108 41177
rect 79901 40461 79904 40739
rect 79983 40461 80108 40739
rect 79901 40079 80108 40461
rect 81965 40703 82114 41189
rect 82045 40420 82114 40703
rect 81965 40056 82114 40420
rect 66873 37203 67174 37279
rect 66873 37088 66934 37203
rect 68727 37106 68833 37245
rect 70491 37290 70780 37309
rect 66873 36911 67174 37088
rect 68727 36908 69023 37106
rect 70491 37090 70550 37290
rect 72312 37285 72635 37309
rect 70491 36904 70780 37090
rect 72312 37085 72364 37285
rect 72608 37085 72635 37285
rect 72312 36900 72635 37085
rect 101389 37196 101690 37272
rect 101389 37081 101450 37196
rect 103243 37099 103349 37238
rect 105007 37283 105296 37302
rect 101389 36904 101690 37081
rect 103243 36901 103539 37099
rect 105007 37083 105066 37283
rect 106828 37278 107151 37302
rect 105007 36897 105296 37083
rect 106828 37078 106880 37278
rect 107124 37078 107151 37278
rect 106828 36893 107151 37078
rect 85494 24870 86377 24976
rect 86495 24870 86637 24976
rect 85494 24786 86637 24870
rect 40305 23742 41228 23862
rect 41356 23742 41450 23862
rect 40305 23654 41450 23742
rect 50980 23721 51068 23836
rect 51186 23721 52123 23836
rect 50980 23646 52123 23721
rect 62890 23722 62988 23839
rect 63106 23722 64033 23839
rect 62890 23649 64033 23722
rect 71474 23719 71557 23837
rect 71675 23719 72617 23837
rect 71474 23647 72617 23719
rect 82154 23772 83297 23784
rect 82154 23654 83055 23772
rect 83173 23654 83297 23772
rect 82154 23594 83297 23654
rect 85506 23722 86649 23783
rect 85506 23604 85591 23722
rect 85709 23604 86649 23722
rect 85506 23593 86649 23604
rect 91748 23670 92590 23782
rect 92708 23670 92891 23782
rect 91748 23592 92891 23670
rect 105662 23300 106372 23418
rect 106500 23300 106805 23418
rect 105662 23228 106805 23300
rect 40292 22578 41437 22649
rect 40292 22450 40383 22578
rect 40511 22450 41437 22578
rect 50992 22587 52135 22643
rect 50992 22469 51940 22587
rect 52058 22469 52135 22587
rect 50992 22453 52135 22469
rect 62902 22582 64045 22646
rect 62902 22464 63860 22582
rect 63978 22464 64045 22582
rect 62902 22456 64045 22464
rect 71486 22578 72629 22644
rect 71486 22460 72435 22578
rect 72553 22460 72629 22578
rect 71486 22454 72629 22460
rect 82166 22522 83309 22591
rect 40292 22441 41437 22450
rect 82166 22404 82256 22522
rect 82374 22404 83309 22522
rect 82166 22401 83309 22404
rect 91760 22528 92903 22589
rect 91760 22410 91882 22528
rect 92000 22410 92903 22528
rect 91760 22399 92903 22410
rect 105674 22156 106817 22225
rect 105674 22035 105796 22156
rect 105924 22035 106817 22156
rect 36746 21755 36843 21870
rect 36971 21755 37891 21870
rect 36746 21662 37891 21755
rect 47662 21719 47795 21843
rect 47923 21719 48805 21843
rect 43338 21534 43434 21652
rect 47662 21653 48805 21719
rect 60161 21753 60239 21840
rect 60357 21753 61304 21840
rect 43562 21534 44481 21652
rect 60161 21650 61304 21753
rect 43338 21462 44481 21534
rect 66614 20832 67099 20835
rect 36733 20579 37878 20657
rect 36733 20451 37638 20579
rect 37766 20451 37878 20579
rect 47674 20577 48817 20650
rect 47674 20460 48603 20577
rect 36733 20449 37878 20451
rect 43350 20397 44493 20459
rect 48731 20460 48817 20577
rect 60173 20579 61316 20647
rect 60173 20461 61061 20579
rect 61179 20461 61316 20579
rect 60173 20457 61316 20461
rect 43350 20269 44260 20397
rect 44388 20269 44493 20397
rect 66537 20332 67099 20832
rect 66537 20214 66649 20332
rect 66767 20214 67099 20332
rect 36735 19757 36843 19859
rect 36971 19757 37880 19859
rect 36735 19651 37880 19757
rect 47662 19714 47791 19842
rect 47919 19714 48805 19842
rect 43344 19526 43415 19654
rect 43543 19526 44487 19654
rect 47662 19652 48805 19714
rect 60158 19723 60241 19836
rect 60359 19723 61301 19836
rect 60158 19646 61301 19723
rect 66537 19703 67099 20214
rect 68106 20324 68577 20840
rect 73798 20585 73980 20586
rect 68106 20206 68386 20324
rect 68504 20206 68577 20324
rect 68106 19705 68577 20206
rect 73418 20070 73980 20585
rect 73418 19952 73565 20070
rect 73683 19952 73980 20070
rect 43344 19464 44487 19526
rect 73418 19467 73980 19952
rect 74987 20093 75458 20586
rect 74987 19975 75276 20093
rect 75394 19975 75458 20093
rect 74987 19469 75458 19975
rect 74987 19467 75169 19469
rect 36722 18578 37867 18646
rect 36722 18450 37633 18578
rect 37761 18450 37867 18578
rect 47674 18578 48817 18649
rect 47674 18459 48603 18578
rect 36722 18438 37867 18450
rect 43356 18389 44499 18456
rect 48731 18459 48817 18578
rect 60170 18583 61313 18643
rect 60170 18465 61055 18583
rect 61173 18465 61313 18583
rect 60170 18453 61313 18465
rect 43356 18266 44259 18389
rect 44387 18266 44499 18389
rect 40306 17738 40397 17850
rect 40525 17738 41449 17850
rect 71484 17844 72627 17847
rect 40306 17660 41449 17738
rect 50965 17722 51104 17835
rect 51222 17722 52108 17835
rect 50965 17645 52108 17722
rect 62893 17715 63015 17830
rect 63133 17715 64036 17830
rect 62893 17640 64036 17715
rect 71484 17726 71584 17844
rect 71702 17726 72627 17844
rect 71484 17657 72627 17726
rect 82147 17695 82968 17808
rect 83086 17695 83290 17808
rect 82147 17618 83290 17695
rect 91775 17701 92566 17814
rect 92684 17701 92918 17814
rect 91775 17624 92918 17701
rect 85495 16844 86412 16962
rect 86530 16844 86638 16962
rect 85495 16772 86638 16844
rect 40303 16563 41446 16659
rect 50977 16582 52120 16642
rect 40303 16542 41448 16563
rect 40303 16414 41211 16542
rect 41339 16414 41448 16542
rect 50977 16464 51817 16582
rect 51935 16464 52120 16582
rect 50977 16452 52120 16464
rect 62905 16573 64048 16637
rect 62905 16455 63827 16573
rect 63945 16455 64048 16573
rect 71496 16582 72639 16654
rect 71496 16464 72296 16582
rect 72414 16464 72639 16582
rect 82159 16561 83302 16615
rect 62905 16447 64048 16455
rect 82159 16443 82296 16561
rect 82414 16443 83302 16561
rect 82159 16425 83302 16443
rect 91787 16547 92930 16621
rect 91787 16431 91859 16547
rect 91977 16431 92930 16547
rect 40303 16335 41448 16414
rect 85507 15695 86650 15769
rect 85507 15579 85624 15695
rect 85742 15579 86650 15695
<< viali >>
rect 62920 64987 63118 65021
rect 63684 64989 63797 65102
rect 64254 64987 64452 65021
rect 65058 64998 65171 65111
rect 65632 64987 65830 65021
rect 66421 64998 66534 65111
rect 67010 64987 67208 65021
rect 67770 64999 67883 65112
rect 72920 64987 73118 65021
rect 73684 64989 73797 65102
rect 74254 64987 74452 65021
rect 75058 64998 75171 65111
rect 75632 64987 75830 65021
rect 76421 64998 76534 65111
rect 77010 64987 77208 65021
rect 77770 64999 77883 65112
rect 85128 63757 85318 63849
rect 85590 63746 85976 63780
rect 86485 63764 86629 63858
rect 86924 63746 87310 63780
rect 102782 63757 102972 63849
rect 103244 63746 103630 63780
rect 104139 63764 104283 63858
rect 104578 63746 104964 63780
rect 62731 62076 62844 62189
rect 63429 62033 63542 62146
rect 64378 62045 64491 62159
rect 64721 62064 64834 62177
rect 65456 62056 65569 62169
rect 66175 62038 66288 62151
rect 66828 62030 66941 62143
rect 67543 62038 67656 62151
rect 72731 62076 72844 62189
rect 73429 62033 73542 62146
rect 74378 62045 74491 62159
rect 74721 62064 74834 62177
rect 75456 62056 75569 62169
rect 76175 62038 76288 62151
rect 76828 62030 76941 62143
rect 77543 62038 77656 62151
rect 63052 59916 63305 59993
rect 64372 59915 64680 60000
rect 65760 59918 66042 59989
rect 67132 59920 67414 59991
rect 73052 59916 73305 59993
rect 74372 59915 74680 60000
rect 75760 59918 76042 59989
rect 77132 59920 77414 59991
rect 84943 59523 85056 59636
rect 102597 59523 102710 59636
rect 63937 59238 64050 59351
rect 65298 59250 65411 59363
rect 66660 59268 66773 59381
rect 68044 59303 68157 59416
rect 73937 59238 74050 59351
rect 75298 59250 75411 59363
rect 76660 59268 76773 59381
rect 78044 59303 78157 59416
rect 87336 58917 87449 59030
rect 104990 58917 105103 59030
rect 116738 52386 116866 52514
rect 46153 51695 46271 52282
rect 46469 52217 46503 52251
rect 47280 52217 47314 52251
rect 46469 51257 46503 51291
rect 47280 51257 47314 51291
rect 47493 51229 47608 51852
rect 48197 51690 48307 52230
rect 48469 52227 48503 52261
rect 49280 52227 49314 52261
rect 120662 52363 120933 52467
rect 48469 51267 48503 51301
rect 49280 51267 49314 51301
rect 49511 51249 49654 51907
rect 115289 51273 115385 51725
rect 117729 51316 117832 51778
rect 119326 51001 119407 52130
rect 121709 51027 121804 52123
rect 115989 50709 116141 50861
rect 119936 50772 120225 50944
rect 36423 50220 36457 50254
rect 37234 50220 37268 50254
rect 36202 49483 36285 49927
rect 37447 49792 37567 50285
rect 36423 49260 36457 49294
rect 37234 49260 37268 49294
rect 38423 50220 38457 50254
rect 39234 50220 39268 50254
rect 38144 49278 38243 49857
rect 39493 49780 39608 50313
rect 66106 49946 66426 50266
rect 67970 49987 68198 50219
rect 69664 49968 69892 50200
rect 71483 49979 71711 50211
rect 73267 49976 73495 50208
rect 75052 49974 75280 50206
rect 100630 49952 100950 50272
rect 38423 49260 38457 49294
rect 39234 49260 39268 49294
rect 61874 49454 63310 49488
rect 102494 49993 102722 50225
rect 104188 49974 104416 50206
rect 106007 49985 106235 50217
rect 107791 49982 108019 50214
rect 109576 49980 109804 50212
rect 96390 49447 97826 49481
rect 65284 48532 65560 48632
rect 67176 48617 67374 48651
rect 68976 48617 69174 48651
rect 70776 48617 70974 48651
rect 72576 48617 72774 48651
rect 74376 48617 74574 48651
rect 99808 48538 100084 48638
rect 101700 48623 101898 48657
rect 103500 48623 103698 48657
rect 105300 48623 105498 48657
rect 107100 48623 107298 48657
rect 108900 48623 109098 48657
rect 60492 47278 61496 47309
rect 60492 47140 60539 47278
rect 60539 47140 61454 47278
rect 61454 47140 61496 47278
rect 60492 47109 61496 47140
rect 62063 41659 62235 42598
rect 62908 41656 63080 42595
rect 84789 42901 84823 42935
rect 85600 42901 85634 42935
rect 84505 42267 84628 42609
rect 86789 42901 86823 42935
rect 87600 42901 87634 42935
rect 86529 42262 86618 42646
rect 84789 41941 84823 41975
rect 85600 41941 85634 41975
rect 86789 41941 86823 41975
rect 87600 41941 87634 41975
rect 85433 41827 85631 41861
rect 87433 41827 87631 41861
rect 96578 41666 96750 42605
rect 97423 41663 97595 42602
rect 80196 41097 80230 41131
rect 81007 41097 81041 41131
rect 79904 40461 79983 40739
rect 82196 41097 82230 41131
rect 83007 41097 83041 41131
rect 81965 40420 82045 40703
rect 80196 40137 80230 40171
rect 81007 40137 81041 40171
rect 80840 40023 81038 40057
rect 82196 40137 82230 40171
rect 83007 40137 83041 40171
rect 82840 40023 83038 40057
rect 65330 37034 65572 37149
rect 66934 37088 67176 37203
rect 68833 37106 69077 37306
rect 70550 37090 70794 37290
rect 72364 37085 72608 37285
rect 74336 37079 74580 37279
rect 99846 37027 100088 37142
rect 101450 37081 101692 37196
rect 103349 37099 103593 37299
rect 105066 37083 105310 37283
rect 106880 37078 107124 37278
rect 108852 37072 109096 37272
rect 96849 35740 97596 35851
rect 65846 35700 66232 35734
rect 67646 35700 68032 35734
rect 69446 35700 69832 35734
rect 71246 35700 71632 35734
rect 73046 35700 73432 35734
rect 74846 35700 75232 35734
rect 100362 35693 100748 35727
rect 102162 35693 102548 35727
rect 103962 35693 104348 35727
rect 105762 35693 106148 35727
rect 107562 35693 107948 35727
rect 109362 35693 109748 35727
rect 127227 33664 127585 33698
rect 127647 33228 127681 33602
rect 127647 32677 127681 32963
rect 127227 32581 127585 32615
rect 95427 30789 95711 31246
rect 60986 29648 61191 30188
rect 59363 28460 61033 28687
rect 95203 28464 95762 28684
rect 86377 24870 86495 24988
rect 85595 24671 85629 24705
rect 86555 24671 86589 24705
rect 41228 23742 41356 23870
rect 85595 23860 85629 23894
rect 86555 23860 86589 23894
rect 51068 23721 51186 23839
rect 62988 23722 63106 23840
rect 71557 23719 71675 23837
rect 83055 23654 83173 23772
rect 85591 23604 85709 23722
rect 92590 23670 92708 23788
rect 40384 23533 40418 23567
rect 41344 23533 41378 23567
rect 51062 23528 51096 23562
rect 52022 23528 52056 23562
rect 62992 23528 63026 23562
rect 63952 23528 63986 23562
rect 71556 23529 71590 23563
rect 72516 23529 72550 23563
rect 82235 23481 82269 23515
rect 83195 23481 83229 23515
rect 91836 23481 91870 23515
rect 92796 23481 92830 23515
rect 106372 23300 106500 23428
rect 105759 23108 105793 23142
rect 106719 23108 106753 23142
rect 40384 22722 40418 22756
rect 41344 22722 41378 22756
rect 51062 22717 51096 22751
rect 52022 22717 52056 22751
rect 62992 22717 63026 22751
rect 63952 22717 63986 22751
rect 71556 22718 71590 22752
rect 72516 22718 72550 22752
rect 82235 22670 82269 22704
rect 83195 22670 83229 22704
rect 91836 22670 91870 22704
rect 92796 22670 92830 22704
rect 40383 22450 40511 22578
rect 51940 22469 52058 22587
rect 63860 22464 63978 22582
rect 72435 22460 72553 22578
rect 82256 22404 82374 22522
rect 91882 22410 92000 22528
rect 105759 22297 105793 22331
rect 106719 22297 106753 22331
rect 105796 22028 105924 22156
rect 36843 21755 36971 21883
rect 47795 21719 47923 21847
rect 36809 21535 36843 21569
rect 37769 21535 37803 21569
rect 43434 21534 43562 21662
rect 60239 21753 60357 21871
rect 47752 21528 47786 21562
rect 48712 21528 48746 21562
rect 60272 21528 60306 21562
rect 61232 21528 61266 21562
rect 43427 21348 43461 21382
rect 44387 21348 44421 21382
rect 36809 20724 36843 20758
rect 37769 20724 37803 20758
rect 47752 20717 47786 20751
rect 48712 20717 48746 20751
rect 60272 20717 60306 20751
rect 61232 20717 61266 20751
rect 37638 20451 37766 20579
rect 43427 20537 43461 20571
rect 44387 20537 44421 20571
rect 48603 20449 48731 20577
rect 61061 20461 61179 20579
rect 44260 20269 44388 20397
rect 67183 20738 67217 20772
rect 67994 20738 68028 20772
rect 66649 20214 66767 20332
rect 36843 19757 36971 19885
rect 47791 19714 47919 19842
rect 36809 19535 36843 19569
rect 37769 19535 37803 19569
rect 43415 19526 43543 19654
rect 60241 19723 60359 19841
rect 68386 20206 68504 20324
rect 67183 19778 67217 19812
rect 67994 19778 68028 19812
rect 74056 20493 74090 20527
rect 74867 20493 74901 20527
rect 73565 19952 73683 20070
rect 47752 19528 47786 19562
rect 48712 19528 48746 19562
rect 60272 19528 60306 19562
rect 61232 19528 61266 19562
rect 75276 19975 75394 20093
rect 74056 19533 74090 19567
rect 74867 19533 74901 19567
rect 43427 19348 43461 19382
rect 44387 19348 44421 19382
rect 36809 18724 36843 18758
rect 37769 18724 37803 18758
rect 47752 18717 47786 18751
rect 48712 18717 48746 18751
rect 60272 18717 60306 18751
rect 61232 18717 61266 18751
rect 37633 18450 37761 18578
rect 43427 18537 43461 18571
rect 44387 18537 44421 18571
rect 48603 18450 48731 18578
rect 61055 18465 61173 18583
rect 44259 18261 44387 18389
rect 40397 17738 40525 17866
rect 51104 17722 51222 17840
rect 63015 17715 63133 17833
rect 71584 17726 71702 17844
rect 82968 17695 83086 17813
rect 92566 17701 92684 17819
rect 40384 17533 40418 17567
rect 41344 17533 41378 17567
rect 51062 17528 51096 17562
rect 52022 17528 52056 17562
rect 62992 17528 63026 17562
rect 63952 17528 63986 17562
rect 71556 17539 71590 17573
rect 72516 17539 72550 17573
rect 82235 17511 82269 17545
rect 83195 17511 83229 17545
rect 91836 17511 91870 17545
rect 92796 17511 92830 17545
rect 86412 16844 86530 16962
rect 40384 16722 40418 16756
rect 41344 16722 41378 16756
rect 51062 16717 51096 16751
rect 52022 16717 52056 16751
rect 62992 16717 63026 16751
rect 63952 16717 63986 16751
rect 71556 16728 71590 16762
rect 72516 16728 72550 16762
rect 82235 16700 82269 16734
rect 83195 16700 83229 16734
rect 91836 16700 91870 16734
rect 92796 16700 92830 16734
rect 85595 16661 85629 16695
rect 86555 16661 86589 16695
rect 41211 16414 41339 16542
rect 51817 16464 51935 16582
rect 63827 16455 63945 16573
rect 72296 16464 72414 16582
rect 82296 16443 82414 16561
rect 91859 16429 91977 16547
rect 85595 15850 85629 15884
rect 86555 15850 86589 15884
rect 85624 15577 85742 15695
rect 133786 -193 133820 -159
rect 134074 -271 134128 -220
rect 134205 -269 134259 -218
rect 133157 -330 133211 -279
rect 133296 -330 133350 -279
rect 134350 -325 134384 -291
rect 134984 -399 135030 -146
rect 136360 -328 136769 -289
rect 136824 -390 136868 -228
rect 138302 -236 138336 -202
rect 138474 -236 138508 -202
rect 138646 -236 138680 -202
rect 138818 -236 138852 -202
rect 138990 -236 139024 -202
rect 139195 -236 139229 -202
rect 139372 -236 139406 -202
rect 139544 -236 139578 -202
rect 139716 -236 139750 -202
rect 139888 -236 139922 -202
rect 140060 -236 140094 -202
rect 140232 -236 140266 -202
rect 138261 -339 138381 -293
rect 133786 -1510 133820 -1476
rect 134074 -1588 134128 -1537
rect 134205 -1586 134259 -1535
rect 133157 -1647 133211 -1596
rect 133296 -1647 133350 -1596
rect 134350 -1642 134384 -1608
rect 134984 -1716 135030 -1463
rect 136360 -1645 136769 -1606
rect 136824 -1707 136868 -1545
rect 138302 -1553 138336 -1519
rect 138474 -1553 138508 -1519
rect 138646 -1553 138680 -1519
rect 138818 -1553 138852 -1519
rect 138990 -1553 139024 -1519
rect 139195 -1553 139229 -1519
rect 139372 -1553 139406 -1519
rect 139544 -1553 139578 -1519
rect 139716 -1553 139750 -1519
rect 139888 -1553 139922 -1519
rect 140060 -1553 140094 -1519
rect 140232 -1553 140266 -1519
rect 138261 -1656 138381 -1610
rect 133786 -3157 133820 -3123
rect 134074 -3235 134128 -3184
rect 134205 -3233 134259 -3182
rect 133157 -3294 133211 -3243
rect 133296 -3294 133350 -3243
rect 134350 -3289 134384 -3255
rect 66796 -3376 66830 -3342
rect 134984 -3363 135030 -3110
rect 136360 -3292 136769 -3253
rect 136824 -3354 136868 -3192
rect 138302 -3200 138336 -3166
rect 138474 -3200 138508 -3166
rect 138646 -3200 138680 -3166
rect 138818 -3200 138852 -3166
rect 138990 -3200 139024 -3166
rect 139195 -3200 139229 -3166
rect 139372 -3200 139406 -3166
rect 139544 -3200 139578 -3166
rect 139716 -3200 139750 -3166
rect 139888 -3200 139922 -3166
rect 140060 -3200 140094 -3166
rect 140232 -3200 140266 -3166
rect 138261 -3303 138381 -3257
rect 66796 -3548 66830 -3514
rect 66796 -3720 66830 -3686
rect 66796 -3892 66830 -3858
rect 66796 -4064 66830 -4030
rect 66796 -4236 66830 -4202
rect 66796 -4413 66830 -4379
rect 133786 -4404 133820 -4370
rect 134074 -4482 134128 -4431
rect 134205 -4480 134259 -4429
rect 133157 -4541 133211 -4490
rect 133296 -4541 133350 -4490
rect 134350 -4536 134384 -4502
rect 66796 -4618 66830 -4584
rect 134984 -4610 135030 -4357
rect 136360 -4539 136769 -4500
rect 136824 -4601 136868 -4439
rect 138302 -4447 138336 -4413
rect 138474 -4447 138508 -4413
rect 138646 -4447 138680 -4413
rect 138818 -4447 138852 -4413
rect 138990 -4447 139024 -4413
rect 139195 -4447 139229 -4413
rect 139372 -4447 139406 -4413
rect 139544 -4447 139578 -4413
rect 139716 -4447 139750 -4413
rect 139888 -4447 139922 -4413
rect 140060 -4447 140094 -4413
rect 140232 -4447 140266 -4413
rect 138261 -4550 138381 -4504
rect 66796 -4790 66830 -4756
rect 66796 -4962 66830 -4928
rect 66796 -5134 66830 -5100
rect 66796 -5306 66830 -5272
rect 66881 -5360 66946 -5204
rect 145718 -11385 145752 -11351
rect 146006 -11463 146060 -11412
rect 146137 -11461 146191 -11410
rect 145089 -11522 145143 -11471
rect 145228 -11522 145282 -11471
rect 146282 -11517 146316 -11483
rect 146916 -11591 146962 -11338
rect 148292 -11520 148701 -11481
rect 148756 -11582 148800 -11420
rect 150234 -11428 150268 -11394
rect 150406 -11428 150440 -11394
rect 150578 -11428 150612 -11394
rect 150750 -11428 150784 -11394
rect 150922 -11428 150956 -11394
rect 151127 -11428 151161 -11394
rect 151304 -11428 151338 -11394
rect 151476 -11428 151510 -11394
rect 151648 -11428 151682 -11394
rect 151820 -11428 151854 -11394
rect 151992 -11428 152026 -11394
rect 152164 -11428 152198 -11394
rect 150193 -11531 150313 -11485
<< metal1 >>
rect 103391 71867 104426 71889
rect 36352 71835 37396 71862
rect 36352 70835 36373 71835
rect 37373 70835 37396 71835
rect 36352 70810 37396 70835
rect 43351 71817 44375 71828
rect 43351 70817 43364 71817
rect 44364 70817 44375 71817
rect 36795 70435 36923 70810
rect 43351 70806 44375 70817
rect 57794 71821 58825 71840
rect 57794 70821 57809 71821
rect 58809 70821 58825 71821
rect 74871 71807 75895 71820
rect 43795 70435 43923 70806
rect 57794 70802 58825 70821
rect 64867 71771 65896 71786
rect 58215 70435 58343 70802
rect 64867 70771 64881 71771
rect 65881 70771 65896 71771
rect 74871 70807 74883 71807
rect 75883 70807 75895 71807
rect 94051 71783 95086 71805
rect 74871 70796 75895 70807
rect 85741 71759 86776 71781
rect 64867 70758 65896 70771
rect 65315 70435 65443 70758
rect 75315 70435 75443 70796
rect 85741 70759 85758 71759
rect 86758 70759 86776 71759
rect 94051 70783 94068 71783
rect 95068 70783 95086 71783
rect 103391 70867 103408 71867
rect 104408 70867 104426 71867
rect 103391 70852 104426 70867
rect 94051 70768 95086 70783
rect 85741 70744 86776 70759
rect 86185 70435 86313 70744
rect 94495 70563 94623 70768
rect 103835 70435 103963 70852
rect 35275 67107 35285 70423
rect 35410 67107 35420 70423
rect 38284 67113 38294 70399
rect 38442 67113 38452 70399
rect 42285 67110 42295 70392
rect 42410 67110 42420 70392
rect 36795 66876 36923 67015
rect 36795 66742 36923 66748
rect 43795 66816 43923 67196
rect 45267 67092 45277 70421
rect 45431 67092 45441 70421
rect 56690 67113 56700 70393
rect 56848 67113 56858 70393
rect 59702 67113 59712 70398
rect 59864 67113 59874 70398
rect 63778 67105 63788 70396
rect 63951 67105 63961 70396
rect 58215 66906 58343 67073
rect 65315 66932 65443 67121
rect 66794 67117 66804 70395
rect 66952 67117 66962 70395
rect 73784 67107 73794 70398
rect 73935 67107 73945 70398
rect 76789 67113 76799 70396
rect 76934 67113 76944 70396
rect 84660 67112 84670 70393
rect 84798 67112 84808 70393
rect 87653 67108 87663 70406
rect 87817 67108 87827 70406
rect 92967 67100 92977 70406
rect 93119 67100 93129 70406
rect 95975 67112 95985 70403
rect 96113 67112 96123 70403
rect 102307 67100 102317 70406
rect 102459 67100 102469 70406
rect 105315 67112 105325 70403
rect 105453 67112 105463 70403
rect 75315 66959 75443 67085
rect 75315 66825 75443 66831
rect 86185 66913 86313 67073
rect 65315 66798 65443 66804
rect 86185 66779 86313 66785
rect 58215 66772 58343 66778
rect 43795 66682 43923 66688
rect 94495 66751 94623 67092
rect 103835 66870 103963 67073
rect 103835 66736 103963 66742
rect 94495 66617 94623 66623
rect 65309 65245 65315 65373
rect 65443 65245 65449 65373
rect 75309 65245 75315 65373
rect 75443 65245 75449 65373
rect 65046 65111 65183 65117
rect 63672 65102 63809 65108
rect 62898 64980 62908 65047
rect 63133 64980 63143 65047
rect 63672 64989 63684 65102
rect 63797 64989 63809 65102
rect 63672 64983 63809 64989
rect 64222 64976 64232 65055
rect 64460 64976 64470 65055
rect 65046 64998 65058 65111
rect 65171 64998 65183 65111
rect 66409 65111 66546 65117
rect 65046 64992 65183 64998
rect 65606 64980 65616 65055
rect 65843 64980 65853 65055
rect 66409 64998 66421 65111
rect 66534 64998 66546 65111
rect 67758 65112 67895 65118
rect 66409 64992 66546 64998
rect 66987 64982 66997 65054
rect 67225 64982 67235 65054
rect 67758 64999 67770 65112
rect 67883 64999 67895 65112
rect 75046 65111 75183 65117
rect 73672 65102 73809 65108
rect 67758 64993 67895 64999
rect 66998 64981 67220 64982
rect 72898 64980 72908 65047
rect 73133 64980 73143 65047
rect 73672 64989 73684 65102
rect 73797 64989 73809 65102
rect 73672 64983 73809 64989
rect 74222 64976 74232 65055
rect 74460 64976 74470 65055
rect 75046 64998 75058 65111
rect 75171 64998 75183 65111
rect 76409 65111 76546 65117
rect 75046 64992 75183 64998
rect 75606 64980 75616 65055
rect 75843 64980 75853 65055
rect 76409 64998 76421 65111
rect 76534 64998 76546 65111
rect 77758 65112 77895 65118
rect 76409 64992 76546 64998
rect 76987 64982 76997 65054
rect 77225 64982 77235 65054
rect 77758 64999 77770 65112
rect 77883 64999 77895 65112
rect 77758 64993 77895 64999
rect 76998 64981 77220 64982
rect 86178 64108 86328 64111
rect 86178 63980 86185 64108
rect 86313 63980 86328 64108
rect 86178 63964 86328 63980
rect 103832 64108 103982 64111
rect 103832 63980 103839 64108
rect 103967 63980 103982 64108
rect 103832 63964 103982 63980
rect 86473 63858 86641 63864
rect 85116 63849 85330 63855
rect 85116 63757 85128 63849
rect 85318 63757 85330 63849
rect 85116 63751 85330 63757
rect 85558 63736 85568 63823
rect 86002 63736 86012 63823
rect 86473 63764 86485 63858
rect 86629 63764 86641 63858
rect 104127 63858 104295 63864
rect 102770 63849 102984 63855
rect 86473 63758 86641 63764
rect 86894 63732 86904 63809
rect 87328 63732 87338 63809
rect 102770 63757 102782 63849
rect 102972 63757 102984 63849
rect 102770 63751 102984 63757
rect 103212 63736 103222 63823
rect 103656 63736 103666 63823
rect 104127 63764 104139 63858
rect 104283 63764 104295 63858
rect 104127 63758 104295 63764
rect 104548 63732 104558 63809
rect 104982 63732 104992 63809
rect 85209 62237 85219 62346
rect 85311 62237 85321 62346
rect 86540 62232 86550 62341
rect 86642 62232 86652 62341
rect 102863 62237 102873 62346
rect 102965 62237 102975 62346
rect 104194 62232 104204 62341
rect 104296 62232 104306 62341
rect 62719 62189 62856 62195
rect 62719 62076 62731 62189
rect 62844 62076 62856 62189
rect 72719 62189 72856 62195
rect 64709 62177 64846 62183
rect 64372 62159 64497 62171
rect 62719 62070 62856 62076
rect 63417 62146 63554 62152
rect 63417 62033 63429 62146
rect 63542 62033 63554 62146
rect 64368 62045 64378 62159
rect 64491 62045 64501 62159
rect 64709 62064 64721 62177
rect 64834 62064 64846 62177
rect 64709 62058 64846 62064
rect 65444 62169 65581 62175
rect 65444 62056 65456 62169
rect 65569 62056 65581 62169
rect 65444 62050 65581 62056
rect 66163 62151 66300 62157
rect 64372 62033 64497 62045
rect 66163 62038 66175 62151
rect 66288 62038 66300 62151
rect 67531 62151 67668 62157
rect 63417 62027 63554 62033
rect 66163 62032 66300 62038
rect 66816 62143 66953 62149
rect 66816 62030 66828 62143
rect 66941 62030 66953 62143
rect 67531 62038 67543 62151
rect 67656 62038 67668 62151
rect 72719 62076 72731 62189
rect 72844 62076 72856 62189
rect 74709 62177 74846 62183
rect 74372 62159 74497 62171
rect 72719 62070 72856 62076
rect 73417 62146 73554 62152
rect 67531 62032 67668 62038
rect 73417 62033 73429 62146
rect 73542 62033 73554 62146
rect 74368 62045 74378 62159
rect 74491 62045 74501 62159
rect 74709 62064 74721 62177
rect 74834 62064 74846 62177
rect 74709 62058 74846 62064
rect 75444 62169 75581 62175
rect 75444 62056 75456 62169
rect 75569 62056 75581 62169
rect 75444 62050 75581 62056
rect 76163 62151 76300 62157
rect 74372 62033 74497 62045
rect 76163 62038 76175 62151
rect 76288 62038 76300 62151
rect 77531 62151 77668 62157
rect 66816 62024 66953 62030
rect 73417 62027 73554 62033
rect 76163 62032 76300 62038
rect 76816 62143 76953 62149
rect 76816 62030 76828 62143
rect 76941 62030 76953 62143
rect 77531 62038 77543 62151
rect 77656 62038 77668 62151
rect 77531 62032 77668 62038
rect 76816 62024 76953 62030
rect 63153 61245 63163 61352
rect 63234 61245 63244 61352
rect 65874 61349 65884 61473
rect 65952 61349 65962 61473
rect 63695 61242 63705 61346
rect 63776 61242 63786 61346
rect 64241 61184 64251 61330
rect 64320 61184 64330 61330
rect 64788 61191 64798 61321
rect 64862 61191 64872 61321
rect 66416 61207 66426 61364
rect 66494 61207 66504 61364
rect 66961 61261 66971 61383
rect 67043 61261 67053 61383
rect 67504 61202 67514 61356
rect 67580 61202 67590 61356
rect 73153 61245 73163 61352
rect 73234 61245 73244 61352
rect 75874 61349 75884 61473
rect 75952 61349 75962 61473
rect 73695 61242 73705 61346
rect 73776 61242 73786 61346
rect 74241 61184 74251 61330
rect 74320 61184 74330 61330
rect 74788 61191 74798 61321
rect 74862 61191 74872 61321
rect 76416 61207 76426 61364
rect 76494 61207 76504 61364
rect 76961 61261 76971 61383
rect 77043 61261 77053 61383
rect 77504 61202 77514 61356
rect 77580 61202 77590 61356
rect 65333 60862 65343 61015
rect 65410 60862 65420 61015
rect 75333 60862 75343 61015
rect 75410 60862 75420 61015
rect 86084 60357 86094 60499
rect 86159 60357 86169 60499
rect 103738 60357 103748 60499
rect 103813 60357 103823 60499
rect 85534 60170 85544 60274
rect 85615 60170 85625 60274
rect 86626 60170 86636 60280
rect 86704 60170 86714 60280
rect 103188 60170 103198 60274
rect 103269 60170 103279 60274
rect 104280 60170 104290 60280
rect 104358 60170 104368 60280
rect 64360 60000 64692 60006
rect 63040 59993 63317 59999
rect 63040 59916 63052 59993
rect 63305 59916 63317 59993
rect 63040 59910 63317 59916
rect 64360 59915 64372 60000
rect 64680 59915 64692 60000
rect 74360 60000 74692 60006
rect 64360 59909 64692 59915
rect 65748 59989 66054 59995
rect 65748 59918 65760 59989
rect 66042 59918 66054 59989
rect 65748 59912 66054 59918
rect 67120 59991 67426 59997
rect 67120 59920 67132 59991
rect 67414 59920 67426 59991
rect 67120 59914 67426 59920
rect 73040 59993 73317 59999
rect 73040 59916 73052 59993
rect 73305 59916 73317 59993
rect 73040 59910 73317 59916
rect 74360 59915 74372 60000
rect 74680 59915 74692 60000
rect 74360 59909 74692 59915
rect 75748 59989 76054 59995
rect 75748 59918 75760 59989
rect 76042 59918 76054 59989
rect 75748 59912 76054 59918
rect 77120 59991 77426 59997
rect 77120 59920 77132 59991
rect 77414 59920 77426 59991
rect 77120 59914 77426 59920
rect 84931 59636 85068 59642
rect 84931 59523 84943 59636
rect 85056 59523 85068 59636
rect 84931 59517 85068 59523
rect 102585 59636 102722 59642
rect 102585 59523 102597 59636
rect 102710 59523 102722 59636
rect 102585 59517 102722 59523
rect 68032 59416 68169 59422
rect 66648 59381 66785 59387
rect 65286 59363 65423 59369
rect 63925 59351 64062 59357
rect 63925 59238 63937 59351
rect 64050 59238 64062 59351
rect 65286 59250 65298 59363
rect 65411 59250 65423 59363
rect 66648 59268 66660 59381
rect 66773 59268 66785 59381
rect 68032 59303 68044 59416
rect 68157 59303 68169 59416
rect 78032 59416 78169 59422
rect 76648 59381 76785 59387
rect 75286 59363 75423 59369
rect 68032 59297 68169 59303
rect 73925 59351 74062 59357
rect 66648 59262 66785 59268
rect 65286 59244 65423 59250
rect 63925 59232 64062 59238
rect 73925 59238 73937 59351
rect 74050 59238 74062 59351
rect 75286 59250 75298 59363
rect 75411 59250 75423 59363
rect 76648 59268 76660 59381
rect 76773 59268 76785 59381
rect 78032 59303 78044 59416
rect 78157 59303 78169 59416
rect 78032 59297 78169 59303
rect 76648 59262 76785 59268
rect 75286 59244 75423 59250
rect 73925 59232 74062 59238
rect 87324 59030 87461 59036
rect 87324 58917 87336 59030
rect 87449 58917 87461 59030
rect 87324 58911 87461 58917
rect 104978 59030 105115 59036
rect 104978 58917 104990 59030
rect 105103 58917 105115 59030
rect 104978 58911 105115 58917
rect 64706 58709 64837 58715
rect 63306 58495 63312 58701
rect 63518 58495 63524 58701
rect 64706 58572 64837 58578
rect 66033 58713 66239 58719
rect 73366 58714 73513 58723
rect 73366 58578 73373 58714
rect 73504 58578 73513 58714
rect 74721 58710 74838 58716
rect 76069 58685 76191 58730
rect 76069 58625 76105 58685
rect 76165 58625 76191 58685
rect 76069 58613 76191 58625
rect 74721 58587 74838 58593
rect 73366 58563 73513 58578
rect 66033 58501 66239 58507
rect 85378 58068 85384 58196
rect 85512 58068 85518 58196
rect 86722 58042 86728 58170
rect 86856 58042 86862 58170
rect 103032 58068 103038 58196
rect 103166 58068 103172 58196
rect 104376 58042 104382 58170
rect 104510 58042 104516 58170
rect 58762 57890 58822 57896
rect 76105 57890 76165 57896
rect 58822 57830 76105 57890
rect 58762 57824 58822 57830
rect 76105 57824 76165 57830
rect 38709 57231 38837 57237
rect 43795 57231 43923 57237
rect 82647 57231 82775 57237
rect 38837 57103 43795 57231
rect 43923 57103 82647 57231
rect 38709 57097 38837 57103
rect 43795 57097 43923 57103
rect 82647 57097 82775 57103
rect 104386 56792 104504 56798
rect 114081 56792 114199 56798
rect 104504 56674 114081 56792
rect 104386 56668 104504 56674
rect 114081 56668 114199 56674
rect 36795 56295 36923 56301
rect 80625 56295 80753 56301
rect 36923 56167 80625 56295
rect 36795 56161 36923 56167
rect 80625 56161 80753 56167
rect 92026 55627 92154 55633
rect 94495 55627 94623 55633
rect 64706 55604 64837 55610
rect 61612 55473 61618 55604
rect 61749 55473 64706 55604
rect 64706 55467 64837 55473
rect 78620 55566 78748 55572
rect 78748 55438 86730 55566
rect 86858 55438 86864 55566
rect 92154 55499 94495 55627
rect 92026 55493 92154 55499
rect 94495 55493 94623 55499
rect 103041 55499 103159 55505
rect 112911 55499 113054 55509
rect 78620 55432 78748 55438
rect 103159 55381 112927 55499
rect 113045 55381 113054 55499
rect 103041 55375 103159 55381
rect 112911 55370 113054 55381
rect 85378 54966 85384 54968
rect 79364 54838 79370 54966
rect 79498 54840 85384 54966
rect 85512 54966 85518 54968
rect 85512 54840 85536 54966
rect 79498 54838 85536 54840
rect 48941 53961 49059 53967
rect 48934 53843 48941 53961
rect 49059 53960 120608 53961
rect 49059 53843 87250 53960
rect 48941 53837 49059 53843
rect 87244 53842 87250 53843
rect 87368 53843 120608 53960
rect 87368 53842 87374 53843
rect 85345 53410 85463 53416
rect 46935 53292 85345 53410
rect 85463 53292 116623 53410
rect 46935 52387 47053 53292
rect 85345 53286 85463 53292
rect 48935 52399 48941 52517
rect 49059 52399 49065 52517
rect 46147 52282 46277 52294
rect 46143 51695 46153 52282
rect 46271 51695 46281 52282
rect 46439 52205 46449 52265
rect 46509 52205 46519 52265
rect 47261 52201 47271 52271
rect 47341 52201 47351 52271
rect 48191 52230 48313 52242
rect 47487 51852 47614 51864
rect 46147 51683 46277 51695
rect 46439 51242 46449 51302
rect 46509 51242 46519 51302
rect 46745 51153 46751 51281
rect 46879 51153 46885 51281
rect 47262 51240 47272 51310
rect 47342 51240 47352 51310
rect 47483 51229 47493 51852
rect 47608 51229 47618 51852
rect 48187 51690 48197 52230
rect 48307 51690 48317 52230
rect 48439 52215 48449 52275
rect 48509 52215 48519 52275
rect 49264 52215 49274 52275
rect 49334 52215 49344 52275
rect 116505 52230 116623 53292
rect 116726 52514 116878 52520
rect 116726 52386 116738 52514
rect 116866 52386 116878 52514
rect 116726 52380 116878 52386
rect 120490 52241 120608 53843
rect 120650 52467 120945 52473
rect 120650 52363 120662 52467
rect 120933 52363 120945 52467
rect 120650 52357 120945 52363
rect 119320 52130 119413 52142
rect 49505 51907 49660 51919
rect 48191 51678 48313 51690
rect 48440 51253 48450 51313
rect 48510 51253 48520 51313
rect 48730 51289 48873 51297
rect 47487 51217 47614 51229
rect 48730 51161 48737 51289
rect 48865 51161 48873 51289
rect 49266 51255 49276 51315
rect 49336 51255 49346 51315
rect 49501 51249 49511 51907
rect 49654 51249 49664 51907
rect 117723 51778 117838 51790
rect 115283 51725 115391 51737
rect 58215 51393 58343 51399
rect 57478 51265 58215 51393
rect 115279 51273 115289 51725
rect 115385 51273 115395 51725
rect 117719 51316 117729 51778
rect 117832 51316 117842 51778
rect 117723 51304 117838 51316
rect 49505 51237 49660 51249
rect 48730 51154 48873 51161
rect 57478 50702 57606 51265
rect 58215 51259 58343 51265
rect 115283 51261 115391 51273
rect 73367 50990 73373 51121
rect 73504 50990 73510 51121
rect 119316 51001 119326 52130
rect 119407 51001 119417 52130
rect 121703 52123 121810 52135
rect 121699 51027 121709 52123
rect 121804 51027 121814 52123
rect 121703 51015 121810 51027
rect 119320 50989 119413 51001
rect 36789 50498 36795 50626
rect 36923 50498 36929 50626
rect 38703 50500 38709 50628
rect 38837 50500 38843 50628
rect 91952 50598 91962 50845
rect 92205 50598 92215 50845
rect 115569 50800 115579 50928
rect 115707 50800 115717 50928
rect 117386 50869 117396 50953
rect 117553 50869 117563 50953
rect 119924 50944 120237 50950
rect 115977 50861 116153 50867
rect 115977 50709 115989 50861
rect 116141 50709 116153 50861
rect 119924 50772 119936 50944
rect 120225 50772 120237 50944
rect 121186 50888 121196 50958
rect 121516 50888 121526 50958
rect 119924 50766 120237 50772
rect 115977 50703 116153 50709
rect 36795 50381 36923 50498
rect 38709 50376 38837 50500
rect 39487 50313 39614 50325
rect 37441 50285 37573 50297
rect 36398 50207 36408 50263
rect 36464 50207 36474 50263
rect 37218 50211 37228 50271
rect 37288 50211 37298 50271
rect 36196 49927 36291 49939
rect 36192 49483 36202 49927
rect 36285 49483 36295 49927
rect 37437 49792 37447 50285
rect 37567 49792 37577 50285
rect 38394 50209 38404 50269
rect 38464 50209 38474 50269
rect 39217 50205 39227 50265
rect 39287 50205 39297 50265
rect 38138 49857 38249 49869
rect 37441 49780 37573 49792
rect 36196 49471 36291 49483
rect 36398 49248 36408 49304
rect 36464 49248 36474 49304
rect 36683 49210 36693 49338
rect 36821 49210 36831 49338
rect 37217 49249 37227 49309
rect 37287 49249 37297 49309
rect 38134 49278 38144 49857
rect 38243 49278 38253 49857
rect 39483 49780 39493 50313
rect 39608 49780 39618 50313
rect 100618 50272 100962 50278
rect 66094 50266 66438 50272
rect 66094 49946 66106 50266
rect 66426 49946 66438 50266
rect 67964 50219 68204 50231
rect 67960 49987 67970 50219
rect 68198 49987 68208 50219
rect 69658 50200 69898 50212
rect 71477 50211 71717 50223
rect 67964 49975 68204 49987
rect 69654 49968 69664 50200
rect 69892 49968 69902 50200
rect 71473 49979 71483 50211
rect 71711 49979 71721 50211
rect 73261 50208 73501 50220
rect 69658 49956 69898 49968
rect 71477 49967 71717 49979
rect 73257 49976 73267 50208
rect 73495 49976 73505 50208
rect 75046 50206 75286 50218
rect 73261 49964 73501 49976
rect 75042 49974 75052 50206
rect 75280 49974 75290 50206
rect 75046 49962 75286 49974
rect 100618 49952 100630 50272
rect 100950 49952 100962 50272
rect 102488 50225 102728 50237
rect 116873 50236 116991 50242
rect 120884 50236 121002 50242
rect 126619 50236 126751 50243
rect 102484 49993 102494 50225
rect 102722 49993 102732 50225
rect 104182 50206 104422 50218
rect 106001 50217 106241 50229
rect 102488 49981 102728 49993
rect 104178 49974 104188 50206
rect 104416 49974 104426 50206
rect 105997 49985 106007 50217
rect 106235 49985 106245 50217
rect 107785 50214 108025 50226
rect 104182 49962 104422 49974
rect 106001 49973 106241 49985
rect 107781 49982 107791 50214
rect 108019 49982 108029 50214
rect 109570 50212 109810 50224
rect 107785 49970 108025 49982
rect 109566 49980 109576 50212
rect 109804 49980 109814 50212
rect 116991 50118 120884 50236
rect 121002 50118 126626 50236
rect 126744 50118 126751 50236
rect 116873 50112 116991 50118
rect 120884 50112 121002 50118
rect 126619 50111 126751 50118
rect 109570 49968 109810 49980
rect 100618 49946 100962 49952
rect 66094 49940 66438 49946
rect 39487 49768 39614 49780
rect 62838 49494 62848 49622
rect 61862 49488 62848 49494
rect 61862 49454 61874 49488
rect 63380 49465 63390 49622
rect 63310 49454 63322 49465
rect 61862 49448 63322 49454
rect 96354 49432 96364 49834
rect 97874 49432 97884 49834
rect 116334 49381 116452 49387
rect 120328 49381 120460 49387
rect 125957 49381 126075 49387
rect 38138 49266 38249 49278
rect 38395 49248 38405 49308
rect 38465 49248 38475 49308
rect 38682 49225 38692 49353
rect 38820 49225 38830 49353
rect 39217 49247 39227 49307
rect 39287 49247 39297 49307
rect 116452 49263 120335 49381
rect 120453 49263 125957 49381
rect 116334 49257 116452 49263
rect 120328 49256 120460 49263
rect 125957 49257 126075 49263
rect 65272 48632 65572 48638
rect 65272 48532 65284 48632
rect 65560 48532 65572 48632
rect 67144 48584 67154 48662
rect 67390 48584 67400 48662
rect 68964 48655 69186 48657
rect 68949 48576 68959 48655
rect 69193 48576 69203 48655
rect 70764 48651 70986 48657
rect 72564 48655 72786 48657
rect 70755 48570 70765 48651
rect 70984 48570 70994 48651
rect 72541 48571 72551 48655
rect 72791 48571 72801 48655
rect 74364 48651 74586 48657
rect 74342 48586 74352 48651
rect 74604 48586 74614 48651
rect 99796 48638 100096 48644
rect 99796 48538 99808 48638
rect 100084 48538 100096 48638
rect 101668 48590 101678 48668
rect 101914 48590 101924 48668
rect 103488 48661 103710 48663
rect 103473 48582 103483 48661
rect 103717 48582 103727 48661
rect 105288 48657 105510 48663
rect 107088 48661 107310 48663
rect 105279 48576 105289 48657
rect 105508 48576 105518 48657
rect 107065 48577 107075 48661
rect 107315 48577 107325 48661
rect 108888 48657 109110 48663
rect 108866 48592 108876 48657
rect 109128 48592 109138 48657
rect 99796 48532 100096 48538
rect 65272 48526 65572 48532
rect 36693 48424 36821 48430
rect 46751 48424 46879 48430
rect 36821 48296 46751 48424
rect 36693 48290 36821 48296
rect 46751 48290 46879 48296
rect 56036 47379 56533 47392
rect 48737 47288 48865 47294
rect 38674 47160 38680 47288
rect 38808 47160 48737 47288
rect 48737 47154 48865 47160
rect 56036 46741 56046 47379
rect 56330 46741 56533 47379
rect 60480 47309 61508 47315
rect 60480 47109 60492 47309
rect 61496 47109 61508 47309
rect 61728 47276 61862 47284
rect 61728 47154 61736 47276
rect 61853 47154 61862 47276
rect 61728 47145 61862 47154
rect 60480 47103 61508 47109
rect 90786 46782 90796 47320
rect 91108 46782 91118 47320
rect 94977 47083 94987 47300
rect 96094 47083 96104 47300
rect 56036 46736 56533 46741
rect 38686 45429 38692 45557
rect 38820 45429 44965 45557
rect 45093 45429 45099 45557
rect 85345 43190 85463 43196
rect 85345 43066 85463 43072
rect 87250 43186 87368 43192
rect 87250 43062 87368 43068
rect 84757 42886 84767 42950
rect 84831 42886 84841 42950
rect 85582 42887 85592 42951
rect 85656 42887 85666 42951
rect 86757 42886 86767 42950
rect 86831 42886 86841 42950
rect 87583 42891 87593 42955
rect 87657 42891 87667 42955
rect 62000 41599 62010 42674
rect 62280 41599 62290 42674
rect 62847 41596 62857 42671
rect 63127 41596 63137 42671
rect 86523 42646 86624 42658
rect 84499 42609 84634 42621
rect 63402 41747 63412 42335
rect 63617 41747 63627 42335
rect 84495 42267 84505 42609
rect 84628 42267 84638 42609
rect 84499 42255 84634 42267
rect 86519 42262 86529 42646
rect 86618 42262 86628 42646
rect 86523 42250 86624 42262
rect 84756 41925 84766 41989
rect 84830 41925 84840 41989
rect 85234 41840 85240 41968
rect 85368 41840 85374 41968
rect 85582 41928 85592 41992
rect 85656 41928 85666 41992
rect 86756 41925 86766 41989
rect 86830 41925 86840 41989
rect 85421 41866 85643 41867
rect 85421 41861 85647 41866
rect 85421 41827 85433 41861
rect 85631 41827 85647 41861
rect 87241 41829 87247 41957
rect 87375 41829 87381 41957
rect 87584 41926 87594 41990
rect 87658 41926 87668 41990
rect 87421 41861 87643 41867
rect 85421 41817 85647 41827
rect 87421 41827 87433 41861
rect 87631 41827 87643 41861
rect 87421 41821 87643 41827
rect 85421 41591 86114 41817
rect 80619 41245 80625 41373
rect 80753 41245 80759 41373
rect 82641 41261 82647 41389
rect 82775 41261 82781 41389
rect 85888 41252 86114 41591
rect 87433 41766 87633 41821
rect 87433 41719 87634 41766
rect 87433 41518 88014 41719
rect 96515 41606 96525 42681
rect 96795 41606 96805 42681
rect 97362 41603 97372 42678
rect 97642 41603 97652 42678
rect 97954 41682 97972 42396
rect 98218 41682 98228 42396
rect 85864 41236 86138 41252
rect 87813 41236 88014 41518
rect 80164 41089 80174 41153
rect 80238 41089 80248 41153
rect 80990 41086 81000 41150
rect 81064 41086 81074 41150
rect 82156 41078 82166 41152
rect 82240 41078 82250 41152
rect 82990 41084 83000 41148
rect 83064 41084 83074 41148
rect 85864 41010 85888 41236
rect 86114 41010 86138 41236
rect 85864 40988 86138 41010
rect 87796 41218 88032 41236
rect 87796 41017 87813 41218
rect 88014 41017 88032 41218
rect 87796 41000 88032 41017
rect 79898 40739 79989 40751
rect 79894 40461 79904 40739
rect 79983 40461 79993 40739
rect 81959 40703 82051 40715
rect 79898 40449 79989 40461
rect 81955 40420 81965 40703
rect 82045 40420 82055 40703
rect 81959 40408 82051 40420
rect 80165 40118 80175 40182
rect 80239 40118 80249 40182
rect 80633 40168 80780 40176
rect 80633 40040 80643 40168
rect 80771 40040 80780 40168
rect 80990 40124 81000 40188
rect 81064 40124 81074 40188
rect 82156 40117 82166 40191
rect 82240 40117 82250 40191
rect 82645 40162 82773 40168
rect 80633 40033 80780 40040
rect 80828 40057 81050 40063
rect 80828 40023 80840 40057
rect 81038 40023 81050 40057
rect 82988 40116 82998 40190
rect 83072 40116 83082 40190
rect 82645 40028 82773 40034
rect 82828 40057 83050 40063
rect 80828 40017 81050 40023
rect 82828 40023 82840 40057
rect 83038 40023 83050 40057
rect 82828 40017 83050 40023
rect 80890 39699 81008 40017
rect 82884 39719 83008 40017
rect 117040 39736 117158 39742
rect 81151 39699 81299 39719
rect 80890 39581 81167 39699
rect 81285 39581 81299 39699
rect 82884 39595 83018 39719
rect 83142 39595 83152 39719
rect 114075 39618 114081 39736
rect 114199 39618 117040 39736
rect 117040 39612 117158 39618
rect 80890 39575 81008 39581
rect 81151 39557 81299 39581
rect 86311 39407 86317 39417
rect 56010 39355 56510 39386
rect 56010 38731 56027 39355
rect 56167 38731 56510 39355
rect 82639 39279 82645 39407
rect 82773 39289 86317 39407
rect 86445 39407 86451 39417
rect 87247 39407 87375 39413
rect 86445 39289 87247 39407
rect 82773 39279 87247 39289
rect 87247 39273 87375 39279
rect 56010 38714 56510 38731
rect 82310 38567 82438 38573
rect 85240 38567 85368 38573
rect 80637 38439 80643 38567
rect 80771 38439 82310 38567
rect 82438 38439 85240 38567
rect 82310 38433 82438 38439
rect 85240 38433 85368 38439
rect 90773 38091 90783 38958
rect 91030 38091 91040 38958
rect 114699 38737 114709 39378
rect 115008 38737 115018 39378
rect 85321 37663 85449 37669
rect 85449 37535 86317 37663
rect 86445 37535 86451 37663
rect 85321 37529 85449 37535
rect 68821 37306 69089 37312
rect 65318 37035 65328 37235
rect 65572 37155 65582 37235
rect 65318 37034 65330 37035
rect 65572 37034 65584 37155
rect 66920 37046 66930 37246
rect 67174 37209 67184 37246
rect 67174 37203 67188 37209
rect 67176 37088 67188 37203
rect 68821 37106 68833 37306
rect 69077 37106 69089 37306
rect 103337 37299 103605 37305
rect 68821 37100 69089 37106
rect 70538 37290 70806 37296
rect 67174 37082 67188 37088
rect 70538 37090 70550 37290
rect 70794 37090 70806 37290
rect 70538 37084 70806 37090
rect 72352 37285 72620 37291
rect 72352 37085 72364 37285
rect 72608 37085 72620 37285
rect 67174 37046 67184 37082
rect 72352 37079 72620 37085
rect 74324 37279 74592 37285
rect 74324 37079 74336 37279
rect 74580 37079 74592 37279
rect 74324 37073 74592 37079
rect 65318 37028 65584 37034
rect 99834 37028 99844 37228
rect 100088 37148 100098 37228
rect 99834 37027 99846 37028
rect 100088 37027 100100 37148
rect 101436 37039 101446 37239
rect 101690 37202 101700 37239
rect 101690 37196 101704 37202
rect 101692 37081 101704 37196
rect 103337 37099 103349 37299
rect 103593 37099 103605 37299
rect 103337 37093 103605 37099
rect 105054 37283 105322 37289
rect 101690 37075 101704 37081
rect 105054 37083 105066 37283
rect 105310 37083 105322 37283
rect 105054 37077 105322 37083
rect 106868 37278 107136 37284
rect 106868 37078 106880 37278
rect 107124 37078 107136 37278
rect 101690 37039 101700 37075
rect 106868 37072 107136 37078
rect 108840 37272 109108 37278
rect 108840 37072 108852 37272
rect 109096 37072 109108 37272
rect 108840 37066 109108 37072
rect 123001 37052 123011 38345
rect 123095 37052 123105 38345
rect 99834 37021 100100 37027
rect 89487 36058 89693 36064
rect 86373 36022 86501 36028
rect 86501 35894 89487 36022
rect 86373 35888 86501 35894
rect 89487 35846 89693 35852
rect 96837 35851 97608 35857
rect 65834 35734 66244 35740
rect 65834 35700 65846 35734
rect 65834 35694 65850 35700
rect 65840 35656 65850 35694
rect 66234 35656 66244 35734
rect 67631 35667 67641 35741
rect 68041 35667 68051 35741
rect 69437 35740 69447 35741
rect 69434 35734 69447 35740
rect 69434 35700 69446 35734
rect 69434 35694 69447 35700
rect 69437 35667 69447 35694
rect 69835 35667 69845 35741
rect 96837 35740 96849 35851
rect 97596 35740 97608 35851
rect 71234 35734 71644 35740
rect 71234 35706 71246 35734
rect 71234 35632 71244 35706
rect 71632 35694 71644 35734
rect 73034 35734 73444 35740
rect 73034 35694 73046 35734
rect 73432 35706 73444 35734
rect 71632 35632 71642 35694
rect 73036 35628 73046 35694
rect 73433 35694 73444 35706
rect 74834 35734 75244 35740
rect 96837 35734 97608 35740
rect 74834 35702 74846 35734
rect 75232 35702 75244 35734
rect 100350 35727 100760 35733
rect 73433 35628 73443 35694
rect 74830 35625 74840 35702
rect 75235 35625 75245 35702
rect 100350 35693 100362 35727
rect 100350 35687 100366 35693
rect 100356 35649 100366 35687
rect 100750 35649 100760 35727
rect 102147 35660 102157 35734
rect 102557 35660 102567 35734
rect 103953 35733 103963 35734
rect 103950 35727 103963 35733
rect 103950 35693 103962 35727
rect 103950 35687 103963 35693
rect 103953 35660 103963 35687
rect 104351 35660 104361 35734
rect 105750 35727 106160 35733
rect 105750 35699 105762 35727
rect 105750 35625 105760 35699
rect 106148 35687 106160 35727
rect 107550 35727 107960 35733
rect 107550 35687 107562 35727
rect 107948 35699 107960 35727
rect 106148 35625 106158 35687
rect 107552 35621 107562 35687
rect 107949 35687 107960 35699
rect 109350 35727 109760 35733
rect 109350 35695 109362 35727
rect 109748 35695 109760 35727
rect 107949 35621 107959 35687
rect 109346 35618 109356 35695
rect 109751 35618 109761 35695
rect 123001 35592 123011 36885
rect 123095 35592 123105 36885
rect 108106 35018 108313 35023
rect 83771 34890 83928 34908
rect 88533 34890 88556 34918
rect 83771 34762 83785 34890
rect 83913 34762 88556 34890
rect 83771 34736 83928 34762
rect 88533 34712 88556 34762
rect 88762 34712 88768 34918
rect 106842 34811 107906 35018
rect 108113 35017 108394 35018
rect 110831 35017 111038 35023
rect 107887 34810 108106 34811
rect 108441 34810 108447 35017
rect 111038 34810 114007 35017
rect 114214 34810 114220 35017
rect 108106 34804 108313 34810
rect 110831 34804 111038 34810
rect 67532 33421 67681 33440
rect 60673 33204 63007 33322
rect 67532 33303 67550 33421
rect 67668 33303 67681 33421
rect 67532 33291 67681 33303
rect 60702 33185 60712 33204
rect 60676 31414 61695 31532
rect 60699 31382 60712 31414
rect 55929 31354 56514 31378
rect 33486 31121 33614 31127
rect 35188 31121 35332 31130
rect 33614 30993 35195 31121
rect 35323 30993 35332 31121
rect 33486 30987 33614 30993
rect 35188 30986 35332 30993
rect 55929 30754 55952 31354
rect 56299 30754 56514 31354
rect 55929 30734 56514 30754
rect 60980 30188 61197 30200
rect 60976 29648 60986 30188
rect 61191 29648 61201 30188
rect 60980 29636 61197 29648
rect 59351 28687 61045 28693
rect 59351 28460 59363 28687
rect 61033 28460 61045 28687
rect 59351 28454 61045 28460
rect 61569 28056 61687 31414
rect 61568 27997 61687 28056
rect 35202 27752 35320 27758
rect 35320 27634 44800 27752
rect 44918 27634 44924 27752
rect 35202 27628 35320 27634
rect 61568 27103 61686 27997
rect 53287 26985 53293 27103
rect 53411 26985 61686 27103
rect 50234 26459 50240 26577
rect 50358 26459 58216 26577
rect 58334 26459 58340 26577
rect 54501 25989 54619 25995
rect 62889 25990 63007 33204
rect 67550 27921 67668 33291
rect 67544 27803 67550 27921
rect 67668 27803 67674 27921
rect 68703 27908 68821 34294
rect 83645 33674 83651 33792
rect 83769 33674 88643 33792
rect 88761 33674 88767 33792
rect 72420 33654 72548 33660
rect 72548 33526 78620 33654
rect 78748 33526 78754 33654
rect 72420 33520 72548 33526
rect 95208 33207 97247 33325
rect 95223 33112 95228 33207
rect 73792 32906 73920 32912
rect 73920 32778 79370 32906
rect 79498 32778 79504 32906
rect 73792 32772 73920 32778
rect 77070 31877 77188 31883
rect 77188 31759 81964 31877
rect 82082 31759 82088 31877
rect 77070 31753 77188 31759
rect 86660 31701 86666 31819
rect 86784 31701 87767 31819
rect 87885 31701 87891 31819
rect 95177 31414 96047 31532
rect 95219 31382 95228 31414
rect 95421 31246 95717 31258
rect 95417 30789 95427 31246
rect 95711 30789 95721 31246
rect 95421 30777 95717 30789
rect 90804 30288 90814 30752
rect 91056 30288 91066 30752
rect 77953 29370 78071 29376
rect 84866 29370 84984 29376
rect 77950 29252 77953 29370
rect 78071 29252 84866 29370
rect 77953 29246 78071 29252
rect 84866 29246 84984 29252
rect 95191 28684 95774 28690
rect 95191 28464 95203 28684
rect 95762 28464 95774 28684
rect 95191 28458 95774 28464
rect 82222 28351 82355 28361
rect 79184 28233 79190 28351
rect 79308 28233 82231 28351
rect 82349 28233 82355 28351
rect 82222 28226 82355 28233
rect 68697 27790 68703 27908
rect 68821 27790 68827 27908
rect 69638 27190 69766 27196
rect 69766 27062 72420 27190
rect 72548 27062 72554 27190
rect 69638 27056 69766 27062
rect 80123 27024 80129 27142
rect 80247 27024 85794 27142
rect 85912 27024 85918 27142
rect 88643 26607 88761 26613
rect 95929 26607 96047 31414
rect 88761 26489 96047 26607
rect 88643 26483 88761 26489
rect 61176 25989 63007 25990
rect 54619 25872 63007 25989
rect 54619 25871 61191 25872
rect 54501 25865 54619 25871
rect 40655 25324 40661 25442
rect 40779 25324 55642 25442
rect 55760 25324 55766 25442
rect 56914 25335 57032 25341
rect 67550 25335 67668 25341
rect 57032 25217 67550 25335
rect 56914 25211 57032 25217
rect 67550 25211 67668 25217
rect 97129 25170 97247 33207
rect 104350 27172 104557 34406
rect 109057 34199 112881 34406
rect 113088 34199 113094 34406
rect 123002 34387 123012 35405
rect 123095 34387 123105 35405
rect 128011 34932 129048 34952
rect 125957 34488 126075 34494
rect 125632 34370 125957 34382
rect 128011 34425 128026 34932
rect 127075 34382 128026 34425
rect 126075 34370 128026 34382
rect 125632 34348 128026 34370
rect 127075 34297 128026 34348
rect 125018 33811 125028 34131
rect 125348 33811 125358 34131
rect 128011 33932 128026 34297
rect 129026 33932 129048 34932
rect 128011 33908 129048 33932
rect 127205 33739 127729 33743
rect 126626 33700 126744 33706
rect 104350 27054 104393 27172
rect 104511 27054 104557 27172
rect 104350 27028 104557 27054
rect 107906 32601 108113 32691
rect 123000 32643 123010 33617
rect 123097 32643 123107 33617
rect 125624 33582 126626 33597
rect 127205 33666 127217 33739
rect 127594 33666 127729 33739
rect 127205 33664 127227 33666
rect 127585 33664 127729 33666
rect 127205 33657 127729 33664
rect 127639 33602 127725 33657
rect 126744 33582 127505 33597
rect 125624 33563 127505 33582
rect 126900 33268 126934 33563
rect 127639 33431 127647 33602
rect 127191 33399 127647 33431
rect 126900 33234 127488 33268
rect 126900 32957 126934 33234
rect 127639 33228 127647 33399
rect 127681 33228 127725 33602
rect 127639 33213 127725 33228
rect 127641 32963 127707 32976
rect 126900 32923 127487 32957
rect 126900 32717 126934 32923
rect 126900 32683 127487 32717
rect 127641 32677 127647 32963
rect 127681 32677 127707 32963
rect 127215 32617 127597 32621
rect 127209 32552 127219 32617
rect 127591 32614 127601 32617
rect 127641 32614 127707 32677
rect 127591 32552 127707 32614
rect 127526 32548 127707 32552
rect 107906 27185 108113 32394
rect 114706 30726 114716 31367
rect 115015 30726 115025 31367
rect 122997 31104 123007 32470
rect 123097 31104 123107 32470
rect 124319 30866 124329 31186
rect 124649 30866 124659 31186
rect 122998 29606 123008 30864
rect 123099 29606 123109 30864
rect 112927 28430 113045 28436
rect 113045 28422 113859 28430
rect 113045 28312 117180 28422
rect 112927 28306 113045 28312
rect 113559 28304 117180 28312
rect 117298 28304 117304 28422
rect 107906 27067 107956 27185
rect 108074 27067 108113 27185
rect 107906 27012 108113 27067
rect 94994 25052 95000 25170
rect 95118 25052 97247 25170
rect 86365 24988 86507 24994
rect 86365 24870 86377 24988
rect 86495 24870 86507 24988
rect 86365 24864 86507 24870
rect 70426 24748 70554 24754
rect 70554 24620 73792 24748
rect 73920 24620 73926 24748
rect 85571 24663 85581 24727
rect 85645 24663 85655 24727
rect 86534 24664 86544 24728
rect 86608 24664 86618 24728
rect 70426 24614 70554 24620
rect 36513 24596 36631 24602
rect 36631 24478 43018 24596
rect 43136 24478 43142 24596
rect 36513 24472 36631 24478
rect 88643 24435 88761 24441
rect 81509 24422 81627 24428
rect 68703 24414 68821 24420
rect 59549 24296 59555 24414
rect 59673 24296 68703 24414
rect 81627 24304 85469 24422
rect 86575 24317 88643 24435
rect 88643 24311 88761 24317
rect 81509 24298 81627 24304
rect 68703 24290 68821 24296
rect 41216 23870 41368 23876
rect 41216 23742 41228 23870
rect 41356 23742 41368 23870
rect 41216 23736 41368 23742
rect 51056 23839 51198 23845
rect 51056 23721 51068 23839
rect 51186 23721 51198 23839
rect 51056 23715 51198 23721
rect 62976 23840 63118 23846
rect 62976 23722 62988 23840
rect 63106 23722 63118 23840
rect 62976 23716 63118 23722
rect 71545 23837 71687 23843
rect 85571 23838 85581 23902
rect 85645 23838 85655 23902
rect 86533 23837 86543 23901
rect 86607 23837 86617 23901
rect 71545 23719 71557 23837
rect 71675 23719 71687 23837
rect 92578 23788 92720 23794
rect 71545 23713 71687 23719
rect 83043 23772 83185 23778
rect 83043 23654 83055 23772
rect 83173 23654 83185 23772
rect 83043 23648 83185 23654
rect 85579 23722 85721 23728
rect 85579 23604 85591 23722
rect 85709 23604 85721 23722
rect 92578 23670 92590 23788
rect 92708 23670 92720 23788
rect 92578 23664 92720 23670
rect 85579 23598 85721 23604
rect 40358 23526 40368 23590
rect 40432 23526 40442 23590
rect 41319 23520 41329 23584
rect 41393 23520 41403 23584
rect 51036 23516 51046 23580
rect 51110 23516 51120 23580
rect 52002 23516 52012 23580
rect 52076 23516 52086 23580
rect 62967 23519 62977 23583
rect 63041 23519 63051 23583
rect 63930 23519 63940 23583
rect 64004 23519 64014 23583
rect 71531 23520 71541 23584
rect 71605 23520 71615 23584
rect 72497 23523 72507 23587
rect 72571 23523 72581 23587
rect 82211 23475 82221 23539
rect 82285 23475 82295 23539
rect 83173 23472 83183 23536
rect 83247 23472 83257 23536
rect 91810 23474 91820 23538
rect 91884 23474 91894 23538
rect 92770 23472 92780 23536
rect 92844 23472 92854 23536
rect 106360 23428 106512 23434
rect 106360 23300 106372 23428
rect 106500 23300 106512 23428
rect 106360 23294 106512 23300
rect 88643 23243 88761 23249
rect 33479 23142 33619 23148
rect 33479 23014 33485 23142
rect 33613 23014 40241 23142
rect 41355 23112 46206 23116
rect 33479 23008 33619 23014
rect 41355 22998 43018 23112
rect 43012 22994 43018 22998
rect 43136 22998 46206 23112
rect 46324 22998 50941 23116
rect 53293 23110 53411 23116
rect 43136 22994 43142 22998
rect 52041 22992 53293 23110
rect 59549 23015 59555 23133
rect 59673 23015 62867 23133
rect 70420 23110 70426 23126
rect 63971 23105 67640 23110
rect 63971 22992 65692 23105
rect 53293 22986 53411 22992
rect 65686 22987 65692 22992
rect 65810 22992 67640 23105
rect 67758 22998 70426 23110
rect 70554 23110 70560 23126
rect 83214 23123 83768 23241
rect 83886 23123 83892 23241
rect 88761 23125 91858 23243
rect 93279 23241 93397 23247
rect 70554 22998 71434 23110
rect 77064 23108 77070 23123
rect 67758 22992 71434 22998
rect 65810 22987 65816 22992
rect 72533 22990 74332 23108
rect 74450 23005 77070 23108
rect 77188 23108 77194 23123
rect 79190 23117 79308 23123
rect 88643 23119 88761 23125
rect 92956 23123 93279 23241
rect 93279 23117 93397 23123
rect 77188 23005 77218 23108
rect 74450 22990 77218 23005
rect 79166 22999 79190 23108
rect 81509 23108 81627 23114
rect 79308 22999 81509 23108
rect 79166 22990 81509 22999
rect 81627 22990 82101 23108
rect 105734 23102 105744 23166
rect 105808 23102 105818 23166
rect 106696 23098 106706 23162
rect 106770 23098 106780 23162
rect 81509 22984 81627 22990
rect 40361 22709 40371 22773
rect 40435 22709 40445 22773
rect 41322 22708 41332 22772
rect 41396 22708 41406 22772
rect 51037 22702 51047 22766
rect 51111 22702 51121 22766
rect 51999 22699 52009 22763
rect 52073 22699 52083 22763
rect 62968 22697 62978 22761
rect 63042 22697 63052 22761
rect 63927 22697 63937 22761
rect 64001 22697 64011 22761
rect 71533 22698 71543 22762
rect 71607 22698 71617 22762
rect 72499 22701 72509 22765
rect 72573 22701 72583 22765
rect 82210 22647 82220 22711
rect 82284 22647 82294 22711
rect 83171 22646 83181 22710
rect 83245 22646 83255 22710
rect 91809 22648 91819 22712
rect 91883 22648 91893 22712
rect 92771 22650 92781 22714
rect 92845 22650 92855 22714
rect 107979 22694 108097 22700
rect 104384 22675 104518 22682
rect 51928 22587 52070 22593
rect 40371 22578 40523 22584
rect 40371 22450 40383 22578
rect 40511 22450 40523 22578
rect 51928 22469 51940 22587
rect 52058 22469 52070 22587
rect 51928 22463 52070 22469
rect 63848 22582 63990 22588
rect 63848 22464 63860 22582
rect 63978 22464 63990 22582
rect 63848 22458 63990 22464
rect 72423 22578 72565 22584
rect 72423 22460 72435 22578
rect 72553 22460 72565 22578
rect 104384 22557 104393 22675
rect 104511 22557 105773 22675
rect 106876 22576 107979 22694
rect 107979 22570 108097 22576
rect 104384 22544 104518 22557
rect 91870 22528 92012 22534
rect 72423 22454 72565 22460
rect 82244 22522 82386 22528
rect 40371 22444 40523 22450
rect 82244 22404 82256 22522
rect 82374 22404 82386 22522
rect 91870 22410 91882 22528
rect 92000 22410 92012 22528
rect 91870 22404 92012 22410
rect 82244 22398 82386 22404
rect 105730 22274 105740 22338
rect 105804 22274 105814 22338
rect 106696 22275 106706 22339
rect 106770 22275 106780 22339
rect 58216 22221 58334 22227
rect 63203 22221 63321 22227
rect 58334 22103 63203 22221
rect 58216 22097 58334 22103
rect 63203 22097 63321 22103
rect 105784 22156 105936 22162
rect 105784 22028 105796 22156
rect 105924 22028 105936 22156
rect 105784 22022 105936 22028
rect 36831 21883 36983 21889
rect 36831 21755 36843 21883
rect 36971 21755 36983 21883
rect 60227 21871 60369 21877
rect 36831 21749 36983 21755
rect 47783 21847 47935 21853
rect 47783 21719 47795 21847
rect 47923 21719 47935 21847
rect 60227 21753 60239 21871
rect 60357 21753 60369 21871
rect 60227 21747 60369 21753
rect 47783 21713 47935 21719
rect 43422 21662 43574 21668
rect 36779 21522 36789 21586
rect 36853 21522 36863 21586
rect 37748 21523 37758 21587
rect 37822 21523 37832 21587
rect 43422 21534 43434 21662
rect 43562 21534 43574 21662
rect 43422 21528 43574 21534
rect 47729 21518 47739 21582
rect 47803 21518 47813 21582
rect 48692 21519 48702 21583
rect 48766 21519 48776 21583
rect 60247 21520 60257 21584
rect 60321 21520 60331 21584
rect 61209 21519 61219 21583
rect 61283 21519 61293 21583
rect 43401 21339 43411 21403
rect 43475 21339 43485 21403
rect 44361 21339 44371 21403
rect 44435 21339 44445 21403
rect 33474 21115 33620 21124
rect 33474 20987 33485 21115
rect 33613 20987 36676 21115
rect 38492 21108 38610 21114
rect 44815 21109 44933 21115
rect 37778 20990 38492 21108
rect 43012 20990 43018 21108
rect 43136 20990 43437 21108
rect 44549 20991 44815 21109
rect 47044 21009 47050 21127
rect 47168 21009 47629 21127
rect 53293 21113 53411 21119
rect 48725 20995 53293 21113
rect 59549 20996 59555 21114
rect 59673 20996 60152 21114
rect 63203 21111 63321 21117
rect 64422 21111 64540 21117
rect 33474 20977 33620 20987
rect 38492 20984 38610 20990
rect 44815 20985 44933 20991
rect 53293 20989 53411 20995
rect 61241 20993 63203 21111
rect 63321 20993 64422 21111
rect 63203 20987 63321 20993
rect 64422 20987 64540 20993
rect 36786 20707 36796 20771
rect 36860 20707 36870 20771
rect 37745 20708 37755 20772
rect 37819 20708 37829 20772
rect 47727 20703 47737 20767
rect 47801 20703 47811 20767
rect 48688 20704 48698 20768
rect 48762 20704 48772 20768
rect 60245 20697 60255 20761
rect 60319 20697 60329 20761
rect 61209 20699 61219 20763
rect 61283 20699 61293 20763
rect 67151 20731 67161 20795
rect 67225 20731 67235 20795
rect 67630 20753 67640 20871
rect 67758 20753 67768 20871
rect 67979 20728 67989 20792
rect 68053 20728 68063 20792
rect 37626 20579 37778 20585
rect 37626 20451 37638 20579
rect 37766 20451 37778 20579
rect 43403 20519 43413 20583
rect 43477 20519 43487 20583
rect 44366 20521 44376 20585
rect 44440 20521 44450 20585
rect 48591 20577 48743 20583
rect 37626 20445 37778 20451
rect 48591 20449 48603 20577
rect 48731 20449 48743 20577
rect 61049 20579 61191 20585
rect 61049 20461 61061 20579
rect 61179 20461 61191 20579
rect 74018 20481 74028 20545
rect 74092 20481 74102 20545
rect 74322 20507 74332 20625
rect 74450 20507 74460 20625
rect 74848 20487 74856 20551
rect 74920 20487 74930 20551
rect 61049 20455 61191 20461
rect 48591 20443 48743 20449
rect 44248 20397 44400 20403
rect 44248 20269 44260 20397
rect 44388 20269 44400 20397
rect 44248 20263 44400 20269
rect 66637 20332 66779 20338
rect 66637 20214 66649 20332
rect 66767 20214 66779 20332
rect 66637 20208 66779 20214
rect 68374 20324 68516 20330
rect 68374 20206 68386 20324
rect 68504 20206 68516 20324
rect 93830 20242 94036 20248
rect 68374 20200 68516 20206
rect 83758 20208 83896 20218
rect 93231 20208 93830 20242
rect 44815 20171 44933 20172
rect 45524 20171 45642 20177
rect 44748 20166 45524 20171
rect 38486 20048 38492 20166
rect 38610 20048 44815 20166
rect 44933 20053 45524 20166
rect 75264 20093 75406 20099
rect 44933 20048 44942 20053
rect 44815 20042 44933 20048
rect 45524 20047 45642 20053
rect 73553 20070 73695 20076
rect 73553 19952 73565 20070
rect 73683 19952 73695 20070
rect 75264 19975 75276 20093
rect 75394 19975 75406 20093
rect 83758 20090 83768 20208
rect 83886 20090 93279 20208
rect 93397 20090 93830 20208
rect 83758 20084 83896 20090
rect 93231 20036 93830 20090
rect 93830 20030 94036 20036
rect 75264 19969 75406 19975
rect 73553 19946 73695 19952
rect 36831 19885 36983 19891
rect 36831 19757 36843 19885
rect 36971 19757 36983 19885
rect 36831 19751 36983 19757
rect 47779 19842 47931 19848
rect 47779 19714 47791 19842
rect 47919 19714 47931 19842
rect 60229 19841 60371 19847
rect 60229 19723 60241 19841
rect 60359 19723 60371 19841
rect 67153 19761 67163 19825
rect 67227 19761 67237 19825
rect 67975 19762 67985 19826
rect 68049 19762 68059 19826
rect 60229 19717 60371 19723
rect 47779 19708 47931 19714
rect 43403 19654 43555 19660
rect 36786 19525 36796 19589
rect 36860 19525 36870 19589
rect 37748 19529 37758 19593
rect 37822 19529 37832 19593
rect 43403 19526 43415 19654
rect 43543 19526 43555 19654
rect 43403 19520 43555 19526
rect 47729 19519 47739 19583
rect 47803 19519 47813 19583
rect 48685 19519 48695 19583
rect 48759 19519 48769 19583
rect 60244 19518 60254 19582
rect 60318 19518 60328 19582
rect 61209 19519 61219 19583
rect 61283 19519 61293 19583
rect 67627 19527 67637 19645
rect 67755 19527 67765 19645
rect 74024 19519 74034 19583
rect 74098 19519 74108 19583
rect 74850 19518 74860 19582
rect 74924 19518 74934 19582
rect 74330 19411 74448 19417
rect 43397 19338 43407 19402
rect 43471 19338 43481 19402
rect 44357 19335 44367 19399
rect 44431 19335 44441 19399
rect 74330 19287 74448 19293
rect 46206 19143 46324 19149
rect 35205 19128 35323 19134
rect 35323 19010 36683 19128
rect 38492 19118 38610 19124
rect 35205 19004 35323 19010
rect 37789 19000 38492 19118
rect 38492 18994 38610 19000
rect 42143 19116 42261 19122
rect 42261 18998 43009 19116
rect 43127 18998 43438 19116
rect 44815 19109 44933 19115
rect 42143 18992 42261 18998
rect 44539 18991 44815 19109
rect 46324 19025 47608 19143
rect 53306 19112 53424 19118
rect 46206 19019 46324 19025
rect 48729 18994 53306 19112
rect 56908 18995 56914 19113
rect 57032 18995 60137 19113
rect 63202 19112 63337 19122
rect 61249 18994 63210 19112
rect 63328 18994 65692 19112
rect 65810 18994 65816 19112
rect 44815 18985 44933 18991
rect 53306 18988 53424 18994
rect 63202 18987 63337 18994
rect 95000 18837 95118 18843
rect 36786 18708 36796 18772
rect 36860 18708 36870 18772
rect 37746 18707 37756 18771
rect 37820 18707 37830 18771
rect 47727 18697 47737 18761
rect 47801 18697 47811 18761
rect 48687 18696 48697 18760
rect 48761 18696 48771 18760
rect 60247 18699 60257 18763
rect 60321 18699 60331 18763
rect 61211 18701 61221 18765
rect 61285 18701 61295 18765
rect 87761 18719 87767 18837
rect 87885 18719 88626 18837
rect 88744 18719 95000 18837
rect 95000 18713 95118 18719
rect 37621 18578 37773 18584
rect 37621 18450 37633 18578
rect 37761 18450 37773 18578
rect 43401 18518 43411 18582
rect 43475 18518 43485 18582
rect 44362 18517 44372 18581
rect 44436 18517 44446 18581
rect 48591 18578 48743 18584
rect 37621 18444 37773 18450
rect 48591 18450 48603 18578
rect 48731 18450 48743 18578
rect 61043 18583 61185 18589
rect 61043 18465 61055 18583
rect 61173 18465 61185 18583
rect 61043 18459 61185 18465
rect 48591 18444 48743 18450
rect 44247 18389 44399 18395
rect 44247 18261 44259 18389
rect 44387 18261 44399 18389
rect 44247 18255 44399 18261
rect 55642 18168 55760 18174
rect 54501 18089 54619 18095
rect 53300 17971 53306 18089
rect 53424 17971 54501 18089
rect 55760 18050 63210 18168
rect 63328 18050 63334 18168
rect 55642 18044 55760 18050
rect 54501 17965 54619 17971
rect 40385 17866 40537 17872
rect 40385 17738 40397 17866
rect 40525 17738 40537 17866
rect 40385 17732 40537 17738
rect 51092 17840 51234 17846
rect 51092 17722 51104 17840
rect 51222 17722 51234 17840
rect 71572 17844 71714 17850
rect 51092 17716 51234 17722
rect 63003 17833 63145 17839
rect 63003 17715 63015 17833
rect 63133 17715 63145 17833
rect 71572 17726 71584 17844
rect 71702 17726 71714 17844
rect 92554 17819 92696 17825
rect 71572 17720 71714 17726
rect 82956 17813 83098 17819
rect 63003 17709 63145 17715
rect 82956 17695 82968 17813
rect 83086 17695 83098 17813
rect 92554 17701 92566 17819
rect 92684 17701 92696 17819
rect 92554 17695 92696 17701
rect 82956 17689 83098 17695
rect 40357 17523 40367 17587
rect 40431 17523 40441 17587
rect 41323 17522 41333 17586
rect 41397 17522 41407 17586
rect 51034 17518 51044 17582
rect 51108 17518 51118 17582
rect 52001 17519 52011 17583
rect 52075 17519 52085 17583
rect 62970 17517 62980 17581
rect 63044 17517 63054 17581
rect 63932 17518 63942 17582
rect 64006 17518 64016 17582
rect 71533 17529 71543 17593
rect 71607 17529 71617 17593
rect 72491 17530 72501 17594
rect 72565 17530 72575 17594
rect 82213 17503 82223 17567
rect 82287 17503 82297 17567
rect 83176 17503 83186 17567
rect 83250 17503 83260 17567
rect 91818 17503 91828 17567
rect 91892 17503 91902 17567
rect 92770 17501 92780 17565
rect 92844 17501 92854 17565
rect 56914 17157 57032 17163
rect 83205 17161 83768 17279
rect 83886 17161 83892 17279
rect 93279 17274 93397 17280
rect 43003 17115 43009 17127
rect 35205 17093 35323 17099
rect 35323 16975 40252 17093
rect 41359 17009 43009 17115
rect 43127 17115 43133 17127
rect 43127 17009 47050 17115
rect 41359 16997 47050 17009
rect 47168 16997 50925 17115
rect 53306 17109 53424 17115
rect 52034 16991 53306 17109
rect 57032 17039 62853 17157
rect 88620 17155 88626 17273
rect 88744 17155 91851 17273
rect 92953 17156 93279 17274
rect 93279 17150 93397 17156
rect 80123 17123 80129 17124
rect 67628 17112 67638 17113
rect 56914 17033 57032 17039
rect 63964 16994 64422 17112
rect 64540 16995 67638 17112
rect 67756 17112 67766 17113
rect 67756 17086 71417 17112
rect 67756 16995 69638 17086
rect 64540 16994 69638 16995
rect 53306 16985 53424 16991
rect 35205 16969 35323 16975
rect 69632 16958 69638 16994
rect 69766 16994 71417 17086
rect 72540 17005 74330 17123
rect 74448 17121 78096 17123
rect 74448 17005 77953 17121
rect 77947 17003 77953 17005
rect 78071 17005 78096 17121
rect 80111 17006 80129 17123
rect 80247 17123 80253 17124
rect 81500 17123 81640 17137
rect 80247 17006 81510 17123
rect 80111 17005 81510 17006
rect 81628 17005 82093 17123
rect 78071 17003 78077 17005
rect 69766 16958 69772 16994
rect 81500 16993 81640 17005
rect 86400 16962 86542 16968
rect 86400 16844 86412 16962
rect 86530 16844 86542 16962
rect 86400 16838 86542 16844
rect 40360 16701 40370 16765
rect 40434 16701 40444 16765
rect 41318 16698 41328 16762
rect 41392 16698 41402 16762
rect 51038 16696 51048 16760
rect 51112 16696 51122 16760
rect 51998 16696 52008 16760
rect 52072 16696 52082 16760
rect 62968 16698 62978 16762
rect 63042 16698 63052 16762
rect 63928 16699 63938 16763
rect 64002 16699 64012 16763
rect 71534 16710 71544 16774
rect 71608 16710 71618 16774
rect 72495 16711 72505 16775
rect 72569 16711 72579 16775
rect 82210 16678 82220 16742
rect 82284 16678 82294 16742
rect 83176 16678 83186 16742
rect 83250 16678 83260 16742
rect 85569 16653 85579 16717
rect 85643 16653 85653 16717
rect 86532 16655 86542 16719
rect 86606 16655 86616 16719
rect 91813 16678 91823 16742
rect 91887 16678 91897 16742
rect 92771 16681 92781 16745
rect 92845 16681 92855 16745
rect 51805 16582 51947 16588
rect 41199 16542 41351 16548
rect 41199 16414 41211 16542
rect 41339 16414 41351 16542
rect 51805 16464 51817 16582
rect 51935 16464 51947 16582
rect 72284 16582 72426 16588
rect 51805 16458 51947 16464
rect 63815 16573 63957 16579
rect 63815 16455 63827 16573
rect 63945 16455 63957 16573
rect 72284 16464 72296 16582
rect 72414 16464 72426 16582
rect 72284 16458 72426 16464
rect 82284 16561 82426 16567
rect 63815 16449 63957 16455
rect 82284 16443 82296 16561
rect 82414 16443 82426 16561
rect 82284 16437 82426 16443
rect 91847 16547 91989 16553
rect 91847 16429 91859 16547
rect 91977 16429 91989 16547
rect 88626 16423 88744 16429
rect 91847 16423 91989 16429
rect 41199 16408 41351 16414
rect 81510 16379 81628 16385
rect 81628 16261 85454 16379
rect 86574 16305 88626 16423
rect 88626 16299 88744 16305
rect 81510 16255 81628 16261
rect 85569 15829 85579 15893
rect 85643 15829 85653 15893
rect 86531 15827 86541 15891
rect 86605 15827 86615 15891
rect 85612 15695 85754 15701
rect 85612 15577 85624 15695
rect 85742 15577 85754 15695
rect 85612 15571 85754 15577
rect 135392 -36 135402 33
rect 135875 -36 135885 33
rect 134978 -146 135036 -134
rect 133767 -203 133777 -151
rect 133829 -203 133839 -151
rect 133141 -332 133151 -264
rect 133217 -332 133227 -264
rect 133145 -336 133223 -332
rect 133280 -340 133290 -272
rect 133356 -340 133366 -272
rect 134057 -282 134067 -214
rect 134133 -282 134143 -214
rect 134193 -216 134271 -212
rect 134190 -284 134200 -216
rect 134266 -284 134276 -216
rect 134333 -274 134404 -260
rect 134333 -326 134345 -274
rect 134397 -326 134404 -274
rect 134333 -331 134404 -326
rect 134978 -399 134984 -146
rect 135030 -283 135036 -146
rect 141777 -196 141783 -192
rect 138290 -202 141783 -196
rect 136818 -228 136874 -216
rect 135030 -289 136781 -283
rect 135030 -328 136360 -289
rect 136769 -328 136781 -289
rect 135030 -334 136781 -328
rect 135030 -338 136780 -334
rect 135030 -399 135036 -338
rect 134978 -411 135036 -399
rect 136818 -390 136824 -228
rect 136868 -279 136874 -228
rect 138290 -236 138302 -202
rect 138336 -236 138474 -202
rect 138508 -236 138646 -202
rect 138680 -236 138818 -202
rect 138852 -236 138990 -202
rect 139024 -236 139195 -202
rect 139229 -236 139372 -202
rect 139406 -236 139544 -202
rect 139578 -236 139716 -202
rect 139750 -236 139888 -202
rect 139922 -236 140060 -202
rect 140094 -236 140232 -202
rect 140266 -236 141783 -202
rect 138290 -240 141783 -236
rect 138290 -242 138348 -240
rect 138462 -242 138520 -240
rect 138634 -242 138692 -240
rect 138806 -242 138864 -240
rect 138978 -242 139036 -240
rect 139183 -242 139241 -240
rect 139360 -242 139418 -240
rect 139532 -242 139590 -240
rect 139704 -242 139762 -240
rect 139876 -242 139934 -240
rect 140048 -242 140106 -240
rect 140220 -242 140278 -240
rect 141777 -244 141783 -240
rect 141835 -244 141841 -192
rect 136868 -287 138379 -279
rect 136868 -293 138393 -287
rect 136868 -333 138261 -293
rect 136868 -390 136874 -333
rect 138249 -339 138261 -333
rect 138381 -339 138393 -293
rect 138249 -345 138393 -339
rect 136818 -402 136874 -390
rect 139072 -577 139082 -513
rect 139544 -577 139554 -513
rect 135395 -1351 135405 -1282
rect 135878 -1351 135888 -1282
rect 134978 -1463 135036 -1451
rect 133767 -1520 133777 -1468
rect 133829 -1520 133839 -1468
rect 133141 -1649 133151 -1581
rect 133217 -1649 133227 -1581
rect 133145 -1653 133223 -1649
rect 133280 -1657 133290 -1589
rect 133356 -1657 133366 -1589
rect 134057 -1599 134067 -1531
rect 134133 -1599 134143 -1531
rect 134193 -1533 134271 -1529
rect 134190 -1601 134200 -1533
rect 134266 -1601 134276 -1533
rect 134333 -1591 134404 -1577
rect 134333 -1643 134345 -1591
rect 134397 -1643 134404 -1591
rect 134333 -1648 134404 -1643
rect 134978 -1716 134984 -1463
rect 135030 -1600 135036 -1463
rect 141777 -1513 141783 -1509
rect 138290 -1519 141783 -1513
rect 136818 -1545 136874 -1533
rect 135030 -1606 136781 -1600
rect 135030 -1645 136360 -1606
rect 136769 -1645 136781 -1606
rect 135030 -1651 136781 -1645
rect 135030 -1655 136780 -1651
rect 135030 -1716 135036 -1655
rect 134978 -1728 135036 -1716
rect 136818 -1707 136824 -1545
rect 136868 -1596 136874 -1545
rect 138290 -1553 138302 -1519
rect 138336 -1553 138474 -1519
rect 138508 -1553 138646 -1519
rect 138680 -1553 138818 -1519
rect 138852 -1553 138990 -1519
rect 139024 -1553 139195 -1519
rect 139229 -1553 139372 -1519
rect 139406 -1553 139544 -1519
rect 139578 -1553 139716 -1519
rect 139750 -1553 139888 -1519
rect 139922 -1553 140060 -1519
rect 140094 -1553 140232 -1519
rect 140266 -1553 141783 -1519
rect 138290 -1557 141783 -1553
rect 138290 -1559 138348 -1557
rect 138462 -1559 138520 -1557
rect 138634 -1559 138692 -1557
rect 138806 -1559 138864 -1557
rect 138978 -1559 139036 -1557
rect 139183 -1559 139241 -1557
rect 139360 -1559 139418 -1557
rect 139532 -1559 139590 -1557
rect 139704 -1559 139762 -1557
rect 139876 -1559 139934 -1557
rect 140048 -1559 140106 -1557
rect 140220 -1559 140278 -1557
rect 141777 -1561 141783 -1557
rect 141835 -1561 141841 -1509
rect 136868 -1604 138379 -1596
rect 136868 -1610 138393 -1604
rect 136868 -1650 138261 -1610
rect 136868 -1707 136874 -1650
rect 138249 -1656 138261 -1650
rect 138381 -1656 138393 -1610
rect 138249 -1662 138393 -1656
rect 136818 -1719 136874 -1707
rect 66754 -1842 66882 -1836
rect 139082 -1891 139092 -1827
rect 139554 -1891 139564 -1827
rect 66754 -1976 66882 -1970
rect 66792 -3336 66834 -1976
rect 67093 -2665 67103 -2039
rect 67170 -2665 67180 -2039
rect 71858 -2165 71868 -2037
rect 71996 -2165 72006 -2037
rect 72400 -2172 72410 -2044
rect 72538 -2172 72548 -2044
rect 72944 -2175 72954 -2047
rect 73082 -2175 73092 -2047
rect 73488 -2176 73498 -2048
rect 73626 -2176 73636 -2048
rect 75114 -2164 75124 -2036
rect 75252 -2164 75262 -2036
rect 75659 -2159 75669 -2031
rect 75797 -2159 75807 -2031
rect 76201 -2161 76211 -2033
rect 76339 -2161 76349 -2033
rect 76748 -2161 76758 -2033
rect 76886 -2161 76896 -2033
rect 79466 -2157 79476 -2029
rect 79604 -2157 79614 -2029
rect 80010 -2159 80020 -2031
rect 80148 -2159 80158 -2031
rect 80553 -2157 80563 -2029
rect 80691 -2157 80701 -2029
rect 81096 -2159 81106 -2031
rect 81234 -2159 81244 -2031
rect 82739 -2150 82749 -2022
rect 82877 -2150 82887 -2022
rect 83279 -2155 83289 -2027
rect 83417 -2155 83427 -2027
rect 83820 -2157 83830 -2029
rect 83958 -2157 83968 -2029
rect 84360 -2150 84370 -2022
rect 84498 -2150 84508 -2022
rect 135387 -2997 135397 -2928
rect 135870 -2997 135880 -2928
rect 134978 -3110 135036 -3098
rect 133767 -3167 133777 -3115
rect 133829 -3167 133839 -3115
rect 133141 -3296 133151 -3228
rect 133217 -3296 133227 -3228
rect 133145 -3300 133223 -3296
rect 133280 -3304 133290 -3236
rect 133356 -3304 133366 -3236
rect 134057 -3246 134067 -3178
rect 134133 -3246 134143 -3178
rect 134193 -3180 134271 -3176
rect 134190 -3248 134200 -3180
rect 134266 -3248 134276 -3180
rect 134333 -3238 134404 -3224
rect 134333 -3290 134345 -3238
rect 134397 -3290 134404 -3238
rect 134333 -3295 134404 -3290
rect 66784 -3342 66842 -3336
rect 66784 -3376 66796 -3342
rect 66830 -3376 66842 -3342
rect 134978 -3363 134984 -3110
rect 135030 -3247 135036 -3110
rect 141777 -3160 141783 -3156
rect 138290 -3166 141783 -3160
rect 136818 -3192 136874 -3180
rect 135030 -3253 136781 -3247
rect 135030 -3292 136360 -3253
rect 136769 -3292 136781 -3253
rect 135030 -3298 136781 -3292
rect 135030 -3302 136780 -3298
rect 135030 -3363 135036 -3302
rect 134978 -3375 135036 -3363
rect 136818 -3354 136824 -3192
rect 136868 -3243 136874 -3192
rect 138290 -3200 138302 -3166
rect 138336 -3200 138474 -3166
rect 138508 -3200 138646 -3166
rect 138680 -3200 138818 -3166
rect 138852 -3200 138990 -3166
rect 139024 -3200 139195 -3166
rect 139229 -3200 139372 -3166
rect 139406 -3200 139544 -3166
rect 139578 -3200 139716 -3166
rect 139750 -3200 139888 -3166
rect 139922 -3200 140060 -3166
rect 140094 -3200 140232 -3166
rect 140266 -3200 141783 -3166
rect 138290 -3204 141783 -3200
rect 138290 -3206 138348 -3204
rect 138462 -3206 138520 -3204
rect 138634 -3206 138692 -3204
rect 138806 -3206 138864 -3204
rect 138978 -3206 139036 -3204
rect 139183 -3206 139241 -3204
rect 139360 -3206 139418 -3204
rect 139532 -3206 139590 -3204
rect 139704 -3206 139762 -3204
rect 139876 -3206 139934 -3204
rect 140048 -3206 140106 -3204
rect 140220 -3206 140278 -3204
rect 141777 -3208 141783 -3204
rect 141835 -3208 141841 -3156
rect 136868 -3251 138379 -3243
rect 136868 -3257 138393 -3251
rect 136868 -3297 138261 -3257
rect 136868 -3354 136874 -3297
rect 138249 -3303 138261 -3297
rect 138381 -3303 138393 -3257
rect 138249 -3309 138393 -3303
rect 136818 -3366 136874 -3354
rect 66784 -3382 66842 -3376
rect 66792 -3508 66834 -3382
rect 66784 -3514 66842 -3508
rect 66784 -3548 66796 -3514
rect 66830 -3548 66842 -3514
rect 139072 -3541 139082 -3477
rect 139544 -3541 139554 -3477
rect 66784 -3554 66842 -3548
rect 66792 -3680 66834 -3554
rect 66784 -3686 66842 -3680
rect 66784 -3720 66796 -3686
rect 66830 -3720 66842 -3686
rect 66784 -3726 66842 -3720
rect 66792 -3852 66834 -3726
rect 66784 -3858 66842 -3852
rect 66784 -3892 66796 -3858
rect 66830 -3892 66842 -3858
rect 66784 -3898 66842 -3892
rect 66792 -4024 66834 -3898
rect 66784 -4030 66842 -4024
rect 66784 -4064 66796 -4030
rect 66830 -4064 66842 -4030
rect 66784 -4070 66842 -4064
rect 66792 -4196 66834 -4070
rect 66784 -4202 66842 -4196
rect 66784 -4236 66796 -4202
rect 66830 -4236 66842 -4202
rect 66784 -4242 66842 -4236
rect 66792 -4373 66834 -4242
rect 135389 -4247 135399 -4178
rect 135872 -4247 135882 -4178
rect 134978 -4357 135036 -4345
rect 66784 -4379 66842 -4373
rect 66784 -4413 66796 -4379
rect 66830 -4413 66842 -4379
rect 66784 -4419 66842 -4413
rect 133767 -4414 133777 -4362
rect 133829 -4414 133839 -4362
rect 66792 -4578 66834 -4419
rect 133141 -4543 133151 -4475
rect 133217 -4543 133227 -4475
rect 133145 -4547 133223 -4543
rect 133280 -4551 133290 -4483
rect 133356 -4551 133366 -4483
rect 134057 -4493 134067 -4425
rect 134133 -4493 134143 -4425
rect 134193 -4427 134271 -4423
rect 134190 -4495 134200 -4427
rect 134266 -4495 134276 -4427
rect 134333 -4485 134404 -4471
rect 134333 -4537 134345 -4485
rect 134397 -4537 134404 -4485
rect 134333 -4542 134404 -4537
rect 66784 -4584 66842 -4578
rect 66784 -4618 66796 -4584
rect 66830 -4618 66842 -4584
rect 66784 -4624 66842 -4618
rect 134978 -4610 134984 -4357
rect 135030 -4494 135036 -4357
rect 141777 -4407 141783 -4403
rect 138290 -4413 141783 -4407
rect 136818 -4439 136874 -4427
rect 135030 -4500 136781 -4494
rect 135030 -4539 136360 -4500
rect 136769 -4539 136781 -4500
rect 135030 -4545 136781 -4539
rect 135030 -4549 136780 -4545
rect 135030 -4610 135036 -4549
rect 134978 -4622 135036 -4610
rect 136818 -4601 136824 -4439
rect 136868 -4490 136874 -4439
rect 138290 -4447 138302 -4413
rect 138336 -4447 138474 -4413
rect 138508 -4447 138646 -4413
rect 138680 -4447 138818 -4413
rect 138852 -4447 138990 -4413
rect 139024 -4447 139195 -4413
rect 139229 -4447 139372 -4413
rect 139406 -4447 139544 -4413
rect 139578 -4447 139716 -4413
rect 139750 -4447 139888 -4413
rect 139922 -4447 140060 -4413
rect 140094 -4447 140232 -4413
rect 140266 -4447 141783 -4413
rect 138290 -4451 141783 -4447
rect 138290 -4453 138348 -4451
rect 138462 -4453 138520 -4451
rect 138634 -4453 138692 -4451
rect 138806 -4453 138864 -4451
rect 138978 -4453 139036 -4451
rect 139183 -4453 139241 -4451
rect 139360 -4453 139418 -4451
rect 139532 -4453 139590 -4451
rect 139704 -4453 139762 -4451
rect 139876 -4453 139934 -4451
rect 140048 -4453 140106 -4451
rect 140220 -4453 140278 -4451
rect 141777 -4455 141783 -4451
rect 141835 -4455 141841 -4403
rect 136868 -4498 138379 -4490
rect 136868 -4504 138393 -4498
rect 136868 -4544 138261 -4504
rect 136868 -4601 136874 -4544
rect 138249 -4550 138261 -4544
rect 138381 -4550 138393 -4504
rect 138249 -4556 138393 -4550
rect 136818 -4613 136874 -4601
rect 66792 -4750 66834 -4624
rect 66784 -4756 66842 -4750
rect 66784 -4790 66796 -4756
rect 66830 -4790 66842 -4756
rect 139087 -4788 139097 -4724
rect 139559 -4788 139569 -4724
rect 66784 -4796 66842 -4790
rect 66792 -4922 66834 -4796
rect 66784 -4928 66842 -4922
rect 66784 -4962 66796 -4928
rect 66830 -4962 66842 -4928
rect 66784 -4968 66842 -4962
rect 66792 -5094 66834 -4968
rect 66784 -5100 66842 -5094
rect 66784 -5134 66796 -5100
rect 66830 -5134 66842 -5100
rect 66784 -5140 66842 -5134
rect 66792 -5266 66834 -5140
rect 66875 -5204 66952 -5192
rect 66784 -5272 66842 -5266
rect 66784 -5306 66796 -5272
rect 66830 -5306 66842 -5272
rect 66784 -5312 66842 -5306
rect 66792 -5316 66834 -5312
rect 66875 -5360 66881 -5204
rect 66946 -5360 66952 -5204
rect 66875 -5372 66952 -5360
rect 66550 -6253 66560 -5627
rect 66627 -6253 66637 -5627
rect 66881 -6677 66946 -5372
rect 71071 -6267 71081 -5629
rect 71140 -6267 71150 -5629
rect 74335 -6267 74345 -5629
rect 74404 -6267 74414 -5629
rect 77599 -6267 77609 -5629
rect 77668 -6267 77678 -5629
rect 78687 -6267 78697 -5629
rect 78756 -6267 78766 -5629
rect 81951 -6267 81961 -5629
rect 82020 -6267 82030 -5629
rect 85215 -6267 85225 -5629
rect 85284 -6267 85294 -5629
rect 66846 -6683 66974 -6677
rect 66846 -6817 66974 -6811
rect 71618 -9265 71628 -8627
rect 71687 -9265 71697 -8627
rect 72706 -9265 72716 -8627
rect 72775 -9265 72785 -8627
rect 73794 -9265 73804 -8627
rect 73863 -9265 73873 -8627
rect 74882 -9265 74892 -8627
rect 74951 -9265 74961 -8627
rect 75970 -9265 75980 -8627
rect 76039 -9265 76049 -8627
rect 77058 -9265 77068 -8627
rect 77127 -9265 77137 -8627
rect 78146 -9265 78156 -8627
rect 78215 -9265 78225 -8627
rect 79234 -9265 79244 -8627
rect 79303 -9265 79313 -8627
rect 80322 -9265 80332 -8627
rect 80391 -9265 80401 -8627
rect 81410 -9265 81420 -8627
rect 81479 -9265 81489 -8627
rect 82498 -9265 82508 -8627
rect 82567 -9265 82577 -8627
rect 83586 -9265 83596 -8627
rect 83655 -9265 83665 -8627
rect 84674 -9265 84684 -8627
rect 84743 -9265 84753 -8627
rect 147319 -11225 147329 -11156
rect 147802 -11225 147812 -11156
rect 146910 -11338 146968 -11326
rect 145699 -11395 145709 -11343
rect 145761 -11395 145771 -11343
rect 145073 -11524 145083 -11456
rect 145149 -11524 145159 -11456
rect 145077 -11528 145155 -11524
rect 145212 -11532 145222 -11464
rect 145288 -11532 145298 -11464
rect 145989 -11474 145999 -11406
rect 146065 -11474 146075 -11406
rect 146125 -11408 146203 -11404
rect 146122 -11476 146132 -11408
rect 146198 -11476 146208 -11408
rect 146265 -11466 146336 -11452
rect 146265 -11518 146277 -11466
rect 146329 -11518 146336 -11466
rect 146265 -11523 146336 -11518
rect 146910 -11591 146916 -11338
rect 146962 -11475 146968 -11338
rect 153842 -11388 153848 -11384
rect 150222 -11394 153848 -11388
rect 148750 -11420 148806 -11408
rect 146962 -11481 148713 -11475
rect 146962 -11520 148292 -11481
rect 148701 -11520 148713 -11481
rect 146962 -11526 148713 -11520
rect 146962 -11530 148712 -11526
rect 146962 -11591 146968 -11530
rect 146910 -11603 146968 -11591
rect 148750 -11582 148756 -11420
rect 148800 -11471 148806 -11420
rect 150222 -11428 150234 -11394
rect 150268 -11428 150406 -11394
rect 150440 -11428 150578 -11394
rect 150612 -11428 150750 -11394
rect 150784 -11428 150922 -11394
rect 150956 -11428 151127 -11394
rect 151161 -11428 151304 -11394
rect 151338 -11428 151476 -11394
rect 151510 -11428 151648 -11394
rect 151682 -11428 151820 -11394
rect 151854 -11428 151992 -11394
rect 152026 -11428 152164 -11394
rect 152198 -11428 153848 -11394
rect 150222 -11432 153848 -11428
rect 150222 -11434 150280 -11432
rect 150394 -11434 150452 -11432
rect 150566 -11434 150624 -11432
rect 150738 -11434 150796 -11432
rect 150910 -11434 150968 -11432
rect 151115 -11434 151173 -11432
rect 151292 -11434 151350 -11432
rect 151464 -11434 151522 -11432
rect 151636 -11434 151694 -11432
rect 151808 -11434 151866 -11432
rect 151980 -11434 152038 -11432
rect 152152 -11434 152210 -11432
rect 153842 -11436 153848 -11432
rect 153900 -11436 153906 -11384
rect 148800 -11479 150311 -11471
rect 148800 -11485 150325 -11479
rect 148800 -11525 150193 -11485
rect 148800 -11582 148806 -11525
rect 150181 -11531 150193 -11525
rect 150313 -11531 150325 -11485
rect 150181 -11537 150325 -11531
rect 148750 -11594 148806 -11582
rect 151004 -11769 151014 -11705
rect 151476 -11769 151486 -11705
rect 71069 -14265 71079 -13627
rect 71138 -14265 71148 -13627
rect 72157 -14265 72167 -13627
rect 72226 -14265 72236 -13627
rect 73245 -14265 73255 -13627
rect 73314 -14265 73324 -13627
rect 74333 -14265 74343 -13627
rect 74402 -14265 74412 -13627
rect 75421 -14265 75431 -13627
rect 75490 -14265 75500 -13627
rect 76509 -14265 76519 -13627
rect 76578 -14265 76588 -13627
rect 77597 -14265 77607 -13627
rect 77666 -14265 77676 -13627
rect 78685 -14265 78695 -13627
rect 78754 -14265 78764 -13627
rect 79773 -14265 79783 -13627
rect 79842 -14265 79852 -13627
rect 80861 -14265 80871 -13627
rect 80930 -14265 80940 -13627
rect 81949 -14265 81959 -13627
rect 82018 -14265 82028 -13627
rect 83037 -14265 83047 -13627
rect 83106 -14265 83116 -13627
rect 84125 -14265 84135 -13627
rect 84194 -14265 84204 -13627
rect 85213 -14265 85223 -13627
rect 85282 -14265 85292 -13627
rect 71611 -17271 71621 -16617
rect 71685 -17271 71695 -16617
rect 72699 -17271 72709 -16617
rect 72773 -17271 72783 -16617
rect 73787 -17271 73797 -16617
rect 73861 -17271 73871 -16617
rect 74875 -17271 74885 -16617
rect 74949 -17271 74959 -16617
rect 75963 -17271 75973 -16617
rect 76037 -17271 76047 -16617
rect 77051 -17271 77061 -16617
rect 77125 -17271 77135 -16617
rect 78139 -17271 78149 -16617
rect 78213 -17271 78223 -16617
rect 79227 -17271 79237 -16617
rect 79301 -17271 79311 -16617
rect 80315 -17271 80325 -16617
rect 80389 -17271 80399 -16617
rect 81403 -17271 81413 -16617
rect 81477 -17271 81487 -16617
rect 82491 -17271 82501 -16617
rect 82565 -17271 82575 -16617
rect 83579 -17271 83589 -16617
rect 83653 -17271 83663 -16617
rect 84667 -17271 84677 -16617
rect 84741 -17271 84751 -16617
rect 71065 -22006 71075 -21612
rect 71142 -22006 71152 -21612
rect 72155 -22012 72165 -21618
rect 72232 -22012 72242 -21618
rect 73243 -22012 73253 -21618
rect 73320 -22012 73330 -21618
rect 74331 -22012 74341 -21618
rect 74408 -22012 74418 -21618
rect 75419 -22012 75429 -21618
rect 75496 -22012 75506 -21618
rect 76507 -22012 76517 -21618
rect 76584 -22012 76594 -21618
rect 77595 -22012 77605 -21618
rect 77672 -22012 77682 -21618
rect 81947 -22012 81957 -21618
rect 82024 -22012 82034 -21618
rect 83035 -22012 83045 -21618
rect 83112 -22012 83122 -21618
rect 84123 -22012 84133 -21618
rect 84200 -22012 84210 -21618
rect 85211 -22012 85221 -21618
rect 85288 -22012 85298 -21618
rect 77469 -22175 78509 -22160
rect 77469 -23175 77491 -22175
rect 78491 -23175 78509 -22175
rect 77469 -23196 78509 -23175
<< via1 >>
rect 36373 70835 37373 71835
rect 43364 70817 44364 71817
rect 57809 70821 58809 71821
rect 64881 70771 65881 71771
rect 74883 70807 75883 71807
rect 85758 70759 86758 71759
rect 94068 70783 95068 71783
rect 103408 70867 104408 71867
rect 35285 67107 35410 70423
rect 38294 67113 38442 70399
rect 42295 67110 42410 70392
rect 36795 66748 36923 66876
rect 45277 67092 45431 70421
rect 56700 67113 56848 70393
rect 59712 67113 59864 70398
rect 63788 67105 63951 70396
rect 43795 66688 43923 66816
rect 58215 66778 58343 66906
rect 66804 67117 66952 70395
rect 73794 67107 73935 70398
rect 76799 67113 76934 70396
rect 84670 67112 84798 70393
rect 87663 67108 87817 70406
rect 92977 67100 93119 70406
rect 95985 67112 96113 70403
rect 102317 67100 102459 70406
rect 105325 67112 105453 70403
rect 65315 66804 65443 66932
rect 75315 66831 75443 66959
rect 86185 66785 86313 66913
rect 94495 66623 94623 66751
rect 103835 66742 103963 66870
rect 65315 65245 65443 65373
rect 75315 65245 75443 65373
rect 62908 65021 63133 65047
rect 62908 64987 62920 65021
rect 62920 64987 63118 65021
rect 63118 64987 63133 65021
rect 62908 64980 63133 64987
rect 63684 64989 63797 65102
rect 64232 65021 64460 65055
rect 64232 64987 64254 65021
rect 64254 64987 64452 65021
rect 64452 64987 64460 65021
rect 64232 64976 64460 64987
rect 65058 64998 65171 65111
rect 65616 65021 65843 65055
rect 65616 64987 65632 65021
rect 65632 64987 65830 65021
rect 65830 64987 65843 65021
rect 65616 64980 65843 64987
rect 66421 64998 66534 65111
rect 66997 65021 67225 65054
rect 66997 64987 67010 65021
rect 67010 64987 67208 65021
rect 67208 64987 67225 65021
rect 66997 64982 67225 64987
rect 67770 64999 67883 65112
rect 72908 65021 73133 65047
rect 72908 64987 72920 65021
rect 72920 64987 73118 65021
rect 73118 64987 73133 65021
rect 72908 64980 73133 64987
rect 73684 64989 73797 65102
rect 74232 65021 74460 65055
rect 74232 64987 74254 65021
rect 74254 64987 74452 65021
rect 74452 64987 74460 65021
rect 74232 64976 74460 64987
rect 75058 64998 75171 65111
rect 75616 65021 75843 65055
rect 75616 64987 75632 65021
rect 75632 64987 75830 65021
rect 75830 64987 75843 65021
rect 75616 64980 75843 64987
rect 76421 64998 76534 65111
rect 76997 65021 77225 65054
rect 76997 64987 77010 65021
rect 77010 64987 77208 65021
rect 77208 64987 77225 65021
rect 76997 64982 77225 64987
rect 77770 64999 77883 65112
rect 86185 63980 86313 64108
rect 103839 63980 103967 64108
rect 85128 63757 85318 63849
rect 85568 63780 86002 63823
rect 85568 63746 85590 63780
rect 85590 63746 85976 63780
rect 85976 63746 86002 63780
rect 85568 63736 86002 63746
rect 86485 63764 86629 63858
rect 86904 63780 87328 63809
rect 86904 63746 86924 63780
rect 86924 63746 87310 63780
rect 87310 63746 87328 63780
rect 86904 63732 87328 63746
rect 102782 63757 102972 63849
rect 103222 63780 103656 63823
rect 103222 63746 103244 63780
rect 103244 63746 103630 63780
rect 103630 63746 103656 63780
rect 103222 63736 103656 63746
rect 104139 63764 104283 63858
rect 104558 63780 104982 63809
rect 104558 63746 104578 63780
rect 104578 63746 104964 63780
rect 104964 63746 104982 63780
rect 104558 63732 104982 63746
rect 85219 62237 85311 62346
rect 86550 62232 86642 62341
rect 102873 62237 102965 62346
rect 104204 62232 104296 62341
rect 62731 62076 62844 62189
rect 63429 62033 63542 62146
rect 64378 62045 64491 62159
rect 64721 62064 64834 62177
rect 65456 62056 65569 62169
rect 66175 62038 66288 62151
rect 66828 62030 66941 62143
rect 67543 62038 67656 62151
rect 72731 62076 72844 62189
rect 73429 62033 73542 62146
rect 74378 62045 74491 62159
rect 74721 62064 74834 62177
rect 75456 62056 75569 62169
rect 76175 62038 76288 62151
rect 76828 62030 76941 62143
rect 77543 62038 77656 62151
rect 63163 61245 63234 61352
rect 65884 61349 65952 61473
rect 63705 61242 63776 61346
rect 64251 61184 64320 61330
rect 64798 61191 64862 61321
rect 66426 61207 66494 61364
rect 66971 61261 67043 61383
rect 67514 61202 67580 61356
rect 73163 61245 73234 61352
rect 75884 61349 75952 61473
rect 73705 61242 73776 61346
rect 74251 61184 74320 61330
rect 74798 61191 74862 61321
rect 76426 61207 76494 61364
rect 76971 61261 77043 61383
rect 77514 61202 77580 61356
rect 65343 60862 65410 61015
rect 75343 60862 75410 61015
rect 86094 60357 86159 60499
rect 103748 60357 103813 60499
rect 85544 60170 85615 60274
rect 86636 60170 86704 60280
rect 103198 60170 103269 60274
rect 104290 60170 104358 60280
rect 63052 59916 63305 59993
rect 64372 59915 64680 60000
rect 65760 59918 66042 59989
rect 67132 59920 67414 59991
rect 73052 59916 73305 59993
rect 74372 59915 74680 60000
rect 75760 59918 76042 59989
rect 77132 59920 77414 59991
rect 84943 59523 85056 59636
rect 102597 59523 102710 59636
rect 63937 59238 64050 59351
rect 65298 59250 65411 59363
rect 66660 59268 66773 59381
rect 68044 59303 68157 59416
rect 73937 59238 74050 59351
rect 75298 59250 75411 59363
rect 76660 59268 76773 59381
rect 78044 59303 78157 59416
rect 87336 58917 87449 59030
rect 104990 58917 105103 59030
rect 63312 58495 63518 58701
rect 64706 58578 64837 58709
rect 66033 58507 66239 58713
rect 73373 58578 73504 58714
rect 74721 58593 74838 58710
rect 76105 58625 76165 58685
rect 85384 58068 85512 58196
rect 86728 58042 86856 58170
rect 103038 58068 103166 58196
rect 104382 58042 104510 58170
rect 58762 57830 58822 57890
rect 76105 57830 76165 57890
rect 38709 57103 38837 57231
rect 43795 57103 43923 57231
rect 82647 57103 82775 57231
rect 104386 56674 104504 56792
rect 114081 56674 114199 56792
rect 36795 56167 36923 56295
rect 80625 56167 80753 56295
rect 61618 55473 61749 55604
rect 64706 55473 64837 55604
rect 78620 55438 78748 55566
rect 86730 55438 86858 55566
rect 92026 55499 92154 55627
rect 94495 55499 94623 55627
rect 103041 55381 103159 55499
rect 112927 55381 113045 55499
rect 79370 54838 79498 54966
rect 85384 54840 85512 54968
rect 48941 53843 49059 53961
rect 87250 53842 87368 53960
rect 85345 53292 85463 53410
rect 48941 52399 49059 52517
rect 46153 51695 46271 52282
rect 46449 52251 46509 52265
rect 46449 52217 46469 52251
rect 46469 52217 46503 52251
rect 46503 52217 46509 52251
rect 46449 52205 46509 52217
rect 47271 52251 47341 52271
rect 47271 52217 47280 52251
rect 47280 52217 47314 52251
rect 47314 52217 47341 52251
rect 47271 52201 47341 52217
rect 46449 51291 46509 51302
rect 46449 51257 46469 51291
rect 46469 51257 46503 51291
rect 46503 51257 46509 51291
rect 46449 51242 46509 51257
rect 46751 51153 46879 51281
rect 47272 51291 47342 51310
rect 47272 51257 47280 51291
rect 47280 51257 47314 51291
rect 47314 51257 47342 51291
rect 47272 51240 47342 51257
rect 47493 51229 47608 51852
rect 48197 51690 48307 52230
rect 48449 52261 48509 52275
rect 48449 52227 48469 52261
rect 48469 52227 48503 52261
rect 48503 52227 48509 52261
rect 48449 52215 48509 52227
rect 49274 52261 49334 52275
rect 49274 52227 49280 52261
rect 49280 52227 49314 52261
rect 49314 52227 49334 52261
rect 49274 52215 49334 52227
rect 116738 52386 116866 52514
rect 120662 52363 120933 52467
rect 48450 51301 48510 51313
rect 48450 51267 48469 51301
rect 48469 51267 48503 51301
rect 48503 51267 48510 51301
rect 48450 51253 48510 51267
rect 48737 51161 48865 51289
rect 49276 51301 49336 51315
rect 49276 51267 49280 51301
rect 49280 51267 49314 51301
rect 49314 51267 49336 51301
rect 49276 51255 49336 51267
rect 49511 51249 49654 51907
rect 58215 51265 58343 51393
rect 115289 51273 115385 51725
rect 117729 51316 117832 51778
rect 73373 50990 73504 51121
rect 119326 51001 119407 52130
rect 121709 51027 121804 52123
rect 36795 50498 36923 50626
rect 38709 50500 38837 50628
rect 91962 50598 92205 50845
rect 115579 50800 115707 50928
rect 117396 50869 117553 50953
rect 115989 50709 116141 50861
rect 119936 50772 120225 50944
rect 121196 50888 121516 50958
rect 36408 50254 36464 50263
rect 36408 50220 36423 50254
rect 36423 50220 36457 50254
rect 36457 50220 36464 50254
rect 36408 50207 36464 50220
rect 37228 50254 37288 50271
rect 37228 50220 37234 50254
rect 37234 50220 37268 50254
rect 37268 50220 37288 50254
rect 37228 50211 37288 50220
rect 36202 49483 36285 49927
rect 37447 49792 37567 50285
rect 38404 50254 38464 50269
rect 38404 50220 38423 50254
rect 38423 50220 38457 50254
rect 38457 50220 38464 50254
rect 38404 50209 38464 50220
rect 39227 50254 39287 50265
rect 39227 50220 39234 50254
rect 39234 50220 39268 50254
rect 39268 50220 39287 50254
rect 39227 50205 39287 50220
rect 36408 49294 36464 49304
rect 36408 49260 36423 49294
rect 36423 49260 36457 49294
rect 36457 49260 36464 49294
rect 36408 49248 36464 49260
rect 36693 49210 36821 49338
rect 37227 49294 37287 49309
rect 37227 49260 37234 49294
rect 37234 49260 37268 49294
rect 37268 49260 37287 49294
rect 37227 49249 37287 49260
rect 38144 49278 38243 49857
rect 39493 49780 39608 50313
rect 66174 50013 66362 50207
rect 67970 49987 68198 50219
rect 69664 49968 69892 50200
rect 71483 49979 71711 50211
rect 73267 49976 73495 50208
rect 75052 49974 75280 50206
rect 100698 50019 100886 50213
rect 102494 49993 102722 50225
rect 104188 49974 104416 50206
rect 106007 49985 106235 50217
rect 107791 49982 108019 50214
rect 109576 49980 109804 50212
rect 116873 50118 116991 50236
rect 120884 50118 121002 50236
rect 126626 50118 126744 50236
rect 62848 49488 63380 49622
rect 62848 49465 63310 49488
rect 63310 49465 63380 49488
rect 96364 49481 97874 49834
rect 96364 49447 96390 49481
rect 96390 49447 97826 49481
rect 97826 49447 97874 49481
rect 96364 49432 97874 49447
rect 38405 49294 38465 49308
rect 38405 49260 38423 49294
rect 38423 49260 38457 49294
rect 38457 49260 38465 49294
rect 38405 49248 38465 49260
rect 38692 49225 38820 49353
rect 39227 49294 39287 49307
rect 39227 49260 39234 49294
rect 39234 49260 39268 49294
rect 39268 49260 39287 49294
rect 39227 49247 39287 49260
rect 116334 49263 116452 49381
rect 120335 49263 120453 49381
rect 125957 49263 126075 49381
rect 65284 48532 65560 48632
rect 67154 48651 67390 48662
rect 67154 48617 67176 48651
rect 67176 48617 67374 48651
rect 67374 48617 67390 48651
rect 67154 48584 67390 48617
rect 68959 48651 69193 48655
rect 68959 48617 68976 48651
rect 68976 48617 69174 48651
rect 69174 48617 69193 48651
rect 68959 48576 69193 48617
rect 70765 48617 70776 48651
rect 70776 48617 70974 48651
rect 70974 48617 70984 48651
rect 70765 48570 70984 48617
rect 72551 48651 72791 48655
rect 72551 48617 72576 48651
rect 72576 48617 72774 48651
rect 72774 48617 72791 48651
rect 72551 48571 72791 48617
rect 74352 48617 74376 48651
rect 74376 48617 74574 48651
rect 74574 48617 74604 48651
rect 74352 48586 74604 48617
rect 99808 48538 100084 48638
rect 101678 48657 101914 48668
rect 101678 48623 101700 48657
rect 101700 48623 101898 48657
rect 101898 48623 101914 48657
rect 101678 48590 101914 48623
rect 103483 48657 103717 48661
rect 103483 48623 103500 48657
rect 103500 48623 103698 48657
rect 103698 48623 103717 48657
rect 103483 48582 103717 48623
rect 105289 48623 105300 48657
rect 105300 48623 105498 48657
rect 105498 48623 105508 48657
rect 105289 48576 105508 48623
rect 107075 48657 107315 48661
rect 107075 48623 107100 48657
rect 107100 48623 107298 48657
rect 107298 48623 107315 48657
rect 107075 48577 107315 48623
rect 108876 48623 108900 48657
rect 108900 48623 109098 48657
rect 109098 48623 109128 48657
rect 108876 48592 109128 48623
rect 36693 48296 36821 48424
rect 46751 48296 46879 48424
rect 38680 47160 38808 47288
rect 48737 47160 48865 47288
rect 56046 46741 56330 47379
rect 60492 47109 61496 47309
rect 61736 47154 61853 47276
rect 90796 46782 91108 47320
rect 94987 47083 96094 47300
rect 38692 45429 38820 45557
rect 44965 45429 45093 45557
rect 85345 43072 85463 43190
rect 87250 43068 87368 43186
rect 84767 42935 84831 42950
rect 84767 42901 84789 42935
rect 84789 42901 84823 42935
rect 84823 42901 84831 42935
rect 84767 42886 84831 42901
rect 85592 42935 85656 42951
rect 85592 42901 85600 42935
rect 85600 42901 85634 42935
rect 85634 42901 85656 42935
rect 85592 42887 85656 42901
rect 86767 42935 86831 42950
rect 86767 42901 86789 42935
rect 86789 42901 86823 42935
rect 86823 42901 86831 42935
rect 86767 42886 86831 42901
rect 87593 42935 87657 42955
rect 87593 42901 87600 42935
rect 87600 42901 87634 42935
rect 87634 42901 87657 42935
rect 87593 42891 87657 42901
rect 62010 42598 62280 42674
rect 62010 41659 62063 42598
rect 62063 41659 62235 42598
rect 62235 41659 62280 42598
rect 62010 41599 62280 41659
rect 62857 42595 63127 42671
rect 62857 41656 62908 42595
rect 62908 41656 63080 42595
rect 63080 41656 63127 42595
rect 62857 41596 63127 41656
rect 63412 41747 63617 42335
rect 84505 42267 84628 42609
rect 86529 42262 86618 42646
rect 84766 41975 84830 41989
rect 84766 41941 84789 41975
rect 84789 41941 84823 41975
rect 84823 41941 84830 41975
rect 84766 41925 84830 41941
rect 85240 41840 85368 41968
rect 85592 41975 85656 41992
rect 85592 41941 85600 41975
rect 85600 41941 85634 41975
rect 85634 41941 85656 41975
rect 85592 41928 85656 41941
rect 86766 41975 86830 41989
rect 86766 41941 86789 41975
rect 86789 41941 86823 41975
rect 86823 41941 86830 41975
rect 86766 41925 86830 41941
rect 87247 41829 87375 41957
rect 87594 41975 87658 41990
rect 87594 41941 87600 41975
rect 87600 41941 87634 41975
rect 87634 41941 87658 41975
rect 87594 41926 87658 41941
rect 80625 41245 80753 41373
rect 82647 41261 82775 41389
rect 96525 42605 96795 42681
rect 96525 41666 96578 42605
rect 96578 41666 96750 42605
rect 96750 41666 96795 42605
rect 96525 41606 96795 41666
rect 97372 42602 97642 42678
rect 97372 41663 97423 42602
rect 97423 41663 97595 42602
rect 97595 41663 97642 42602
rect 97372 41603 97642 41663
rect 97972 41682 98218 42396
rect 80174 41131 80238 41153
rect 80174 41097 80196 41131
rect 80196 41097 80230 41131
rect 80230 41097 80238 41131
rect 80174 41089 80238 41097
rect 81000 41131 81064 41150
rect 81000 41097 81007 41131
rect 81007 41097 81041 41131
rect 81041 41097 81064 41131
rect 81000 41086 81064 41097
rect 82166 41131 82240 41152
rect 82166 41097 82196 41131
rect 82196 41097 82230 41131
rect 82230 41097 82240 41131
rect 82166 41078 82240 41097
rect 83000 41131 83064 41148
rect 83000 41097 83007 41131
rect 83007 41097 83041 41131
rect 83041 41097 83064 41131
rect 83000 41084 83064 41097
rect 85888 41010 86114 41236
rect 87813 41017 88014 41218
rect 79904 40461 79983 40739
rect 81965 40420 82045 40703
rect 80175 40171 80239 40182
rect 80175 40137 80196 40171
rect 80196 40137 80230 40171
rect 80230 40137 80239 40171
rect 80175 40118 80239 40137
rect 80643 40040 80771 40168
rect 81000 40171 81064 40188
rect 81000 40137 81007 40171
rect 81007 40137 81041 40171
rect 81041 40137 81064 40171
rect 81000 40124 81064 40137
rect 82166 40171 82240 40191
rect 82166 40137 82196 40171
rect 82196 40137 82230 40171
rect 82230 40137 82240 40171
rect 82166 40117 82240 40137
rect 82645 40034 82773 40162
rect 82998 40171 83072 40190
rect 82998 40137 83007 40171
rect 83007 40137 83041 40171
rect 83041 40137 83072 40171
rect 82998 40116 83072 40137
rect 81167 39581 81285 39699
rect 83018 39595 83142 39719
rect 114081 39618 114199 39736
rect 117040 39618 117158 39736
rect 56027 38731 56167 39355
rect 82645 39279 82773 39407
rect 86317 39289 86445 39417
rect 87247 39279 87375 39407
rect 80643 38439 80771 38567
rect 82310 38439 82438 38567
rect 85240 38439 85368 38567
rect 90783 38091 91030 38958
rect 114709 38737 115008 39378
rect 85321 37535 85449 37663
rect 86317 37535 86445 37663
rect 65328 37149 65572 37235
rect 65328 37035 65330 37149
rect 65330 37035 65572 37149
rect 66930 37203 67174 37246
rect 66930 37088 66934 37203
rect 66934 37088 67174 37203
rect 68833 37106 69077 37306
rect 66930 37046 67174 37088
rect 70550 37090 70794 37290
rect 72364 37085 72608 37285
rect 74336 37079 74580 37279
rect 99844 37142 100088 37228
rect 99844 37028 99846 37142
rect 99846 37028 100088 37142
rect 101446 37196 101690 37239
rect 101446 37081 101450 37196
rect 101450 37081 101690 37196
rect 103349 37099 103593 37299
rect 101446 37039 101690 37081
rect 105066 37083 105310 37283
rect 106880 37078 107124 37278
rect 108852 37072 109096 37272
rect 123011 37052 123095 38345
rect 86373 35894 86501 36022
rect 89487 35852 89693 36058
rect 65850 35700 66232 35734
rect 66232 35700 66234 35734
rect 65850 35656 66234 35700
rect 67641 35734 68041 35741
rect 67641 35700 67646 35734
rect 67646 35700 68032 35734
rect 68032 35700 68041 35734
rect 67641 35667 68041 35700
rect 69447 35734 69835 35741
rect 69447 35700 69832 35734
rect 69832 35700 69835 35734
rect 69447 35667 69835 35700
rect 96849 35740 97596 35851
rect 71244 35700 71246 35706
rect 71246 35700 71632 35706
rect 71244 35632 71632 35700
rect 73046 35700 73432 35706
rect 73432 35700 73433 35706
rect 73046 35628 73433 35700
rect 74840 35700 74846 35702
rect 74846 35700 75232 35702
rect 75232 35700 75235 35702
rect 74840 35625 75235 35700
rect 100366 35693 100748 35727
rect 100748 35693 100750 35727
rect 100366 35649 100750 35693
rect 102157 35727 102557 35734
rect 102157 35693 102162 35727
rect 102162 35693 102548 35727
rect 102548 35693 102557 35727
rect 102157 35660 102557 35693
rect 103963 35727 104351 35734
rect 103963 35693 104348 35727
rect 104348 35693 104351 35727
rect 103963 35660 104351 35693
rect 105760 35693 105762 35699
rect 105762 35693 106148 35699
rect 105760 35625 106148 35693
rect 107562 35693 107948 35699
rect 107948 35693 107949 35699
rect 107562 35621 107949 35693
rect 109356 35693 109362 35695
rect 109362 35693 109748 35695
rect 109748 35693 109751 35695
rect 109356 35618 109751 35693
rect 123011 35592 123095 36885
rect 83785 34762 83913 34890
rect 88556 34712 88762 34918
rect 107906 35017 108113 35018
rect 107906 34811 108441 35017
rect 108106 34810 108441 34811
rect 110831 34810 111038 35017
rect 114007 34810 114214 35017
rect 67550 33303 67668 33421
rect 33486 30993 33614 31121
rect 35195 30993 35323 31121
rect 55952 30754 56299 31354
rect 60986 29648 61191 30188
rect 59363 28460 61033 28687
rect 35202 27634 35320 27752
rect 44800 27634 44918 27752
rect 53293 26985 53411 27103
rect 50240 26459 50358 26577
rect 58216 26459 58334 26577
rect 67550 27803 67668 27921
rect 83651 33674 83769 33792
rect 88643 33674 88761 33792
rect 72420 33526 72548 33654
rect 78620 33526 78748 33654
rect 73792 32778 73920 32906
rect 79370 32778 79498 32906
rect 77070 31759 77188 31877
rect 81964 31759 82082 31877
rect 86666 31701 86784 31819
rect 87767 31701 87885 31819
rect 95427 30789 95711 31246
rect 90814 30288 91056 30752
rect 77953 29252 78071 29370
rect 84866 29252 84984 29370
rect 95203 28464 95762 28684
rect 79190 28233 79308 28351
rect 82231 28233 82349 28351
rect 68703 27790 68821 27908
rect 69638 27062 69766 27190
rect 72420 27062 72548 27190
rect 80129 27024 80247 27142
rect 85794 27024 85912 27142
rect 88643 26489 88761 26607
rect 54501 25871 54619 25989
rect 40661 25324 40779 25442
rect 55642 25324 55760 25442
rect 56914 25217 57032 25335
rect 67550 25217 67668 25335
rect 112881 34199 113088 34406
rect 123012 34387 123095 35405
rect 125957 34370 126075 34488
rect 125028 33811 125348 34131
rect 128026 33932 129026 34932
rect 104393 27054 104511 27172
rect 123010 32643 123097 33617
rect 126626 33582 126744 33700
rect 127217 33698 127594 33739
rect 127217 33666 127227 33698
rect 127227 33666 127585 33698
rect 127585 33666 127594 33698
rect 107906 32394 108113 32601
rect 127219 32615 127591 32617
rect 127219 32581 127227 32615
rect 127227 32581 127585 32615
rect 127585 32581 127591 32615
rect 127219 32552 127591 32581
rect 114716 30726 115015 31367
rect 123007 31104 123097 32470
rect 124329 30866 124649 31186
rect 123008 29606 123099 30864
rect 112927 28312 113045 28430
rect 117180 28304 117298 28422
rect 107956 27067 108074 27185
rect 95000 25052 95118 25170
rect 86377 24870 86495 24988
rect 70426 24620 70554 24748
rect 73792 24620 73920 24748
rect 85581 24705 85645 24727
rect 85581 24671 85595 24705
rect 85595 24671 85629 24705
rect 85629 24671 85645 24705
rect 85581 24663 85645 24671
rect 86544 24705 86608 24728
rect 86544 24671 86555 24705
rect 86555 24671 86589 24705
rect 86589 24671 86608 24705
rect 86544 24664 86608 24671
rect 36513 24478 36631 24596
rect 43018 24478 43136 24596
rect 59555 24296 59673 24414
rect 68703 24296 68821 24414
rect 81509 24304 81627 24422
rect 88643 24317 88761 24435
rect 41228 23742 41356 23870
rect 51068 23721 51186 23839
rect 62988 23722 63106 23840
rect 85581 23894 85645 23902
rect 85581 23860 85595 23894
rect 85595 23860 85629 23894
rect 85629 23860 85645 23894
rect 85581 23838 85645 23860
rect 86543 23894 86607 23901
rect 86543 23860 86555 23894
rect 86555 23860 86589 23894
rect 86589 23860 86607 23894
rect 86543 23837 86607 23860
rect 71557 23719 71675 23837
rect 83055 23654 83173 23772
rect 85591 23604 85709 23722
rect 92590 23670 92708 23788
rect 40368 23567 40432 23590
rect 40368 23533 40384 23567
rect 40384 23533 40418 23567
rect 40418 23533 40432 23567
rect 40368 23526 40432 23533
rect 41329 23567 41393 23584
rect 41329 23533 41344 23567
rect 41344 23533 41378 23567
rect 41378 23533 41393 23567
rect 41329 23520 41393 23533
rect 51046 23562 51110 23580
rect 51046 23528 51062 23562
rect 51062 23528 51096 23562
rect 51096 23528 51110 23562
rect 51046 23516 51110 23528
rect 52012 23562 52076 23580
rect 52012 23528 52022 23562
rect 52022 23528 52056 23562
rect 52056 23528 52076 23562
rect 52012 23516 52076 23528
rect 62977 23562 63041 23583
rect 62977 23528 62992 23562
rect 62992 23528 63026 23562
rect 63026 23528 63041 23562
rect 62977 23519 63041 23528
rect 63940 23562 64004 23583
rect 63940 23528 63952 23562
rect 63952 23528 63986 23562
rect 63986 23528 64004 23562
rect 63940 23519 64004 23528
rect 71541 23563 71605 23584
rect 71541 23529 71556 23563
rect 71556 23529 71590 23563
rect 71590 23529 71605 23563
rect 71541 23520 71605 23529
rect 72507 23563 72571 23587
rect 72507 23529 72516 23563
rect 72516 23529 72550 23563
rect 72550 23529 72571 23563
rect 72507 23523 72571 23529
rect 82221 23515 82285 23539
rect 82221 23481 82235 23515
rect 82235 23481 82269 23515
rect 82269 23481 82285 23515
rect 82221 23475 82285 23481
rect 83183 23515 83247 23536
rect 83183 23481 83195 23515
rect 83195 23481 83229 23515
rect 83229 23481 83247 23515
rect 83183 23472 83247 23481
rect 91820 23515 91884 23538
rect 91820 23481 91836 23515
rect 91836 23481 91870 23515
rect 91870 23481 91884 23515
rect 91820 23474 91884 23481
rect 92780 23515 92844 23536
rect 92780 23481 92796 23515
rect 92796 23481 92830 23515
rect 92830 23481 92844 23515
rect 92780 23472 92844 23481
rect 106372 23300 106500 23428
rect 33485 23014 33613 23142
rect 43018 22994 43136 23112
rect 46206 22998 46324 23116
rect 53293 22992 53411 23110
rect 59555 23015 59673 23133
rect 65692 22987 65810 23105
rect 67640 22992 67758 23110
rect 70426 22998 70554 23126
rect 83768 23123 83886 23241
rect 88643 23125 88761 23243
rect 74332 22990 74450 23108
rect 77070 23005 77188 23123
rect 93279 23123 93397 23241
rect 79190 22999 79308 23117
rect 81509 22990 81627 23108
rect 105744 23142 105808 23166
rect 105744 23108 105759 23142
rect 105759 23108 105793 23142
rect 105793 23108 105808 23142
rect 105744 23102 105808 23108
rect 106706 23142 106770 23162
rect 106706 23108 106719 23142
rect 106719 23108 106753 23142
rect 106753 23108 106770 23142
rect 106706 23098 106770 23108
rect 40371 22756 40435 22773
rect 40371 22722 40384 22756
rect 40384 22722 40418 22756
rect 40418 22722 40435 22756
rect 40371 22709 40435 22722
rect 41332 22756 41396 22772
rect 41332 22722 41344 22756
rect 41344 22722 41378 22756
rect 41378 22722 41396 22756
rect 41332 22708 41396 22722
rect 51047 22751 51111 22766
rect 51047 22717 51062 22751
rect 51062 22717 51096 22751
rect 51096 22717 51111 22751
rect 51047 22702 51111 22717
rect 52009 22751 52073 22763
rect 52009 22717 52022 22751
rect 52022 22717 52056 22751
rect 52056 22717 52073 22751
rect 52009 22699 52073 22717
rect 62978 22751 63042 22761
rect 62978 22717 62992 22751
rect 62992 22717 63026 22751
rect 63026 22717 63042 22751
rect 62978 22697 63042 22717
rect 63937 22751 64001 22761
rect 63937 22717 63952 22751
rect 63952 22717 63986 22751
rect 63986 22717 64001 22751
rect 63937 22697 64001 22717
rect 71543 22752 71607 22762
rect 71543 22718 71556 22752
rect 71556 22718 71590 22752
rect 71590 22718 71607 22752
rect 71543 22698 71607 22718
rect 72509 22752 72573 22765
rect 72509 22718 72516 22752
rect 72516 22718 72550 22752
rect 72550 22718 72573 22752
rect 72509 22701 72573 22718
rect 82220 22704 82284 22711
rect 82220 22670 82235 22704
rect 82235 22670 82269 22704
rect 82269 22670 82284 22704
rect 82220 22647 82284 22670
rect 83181 22704 83245 22710
rect 83181 22670 83195 22704
rect 83195 22670 83229 22704
rect 83229 22670 83245 22704
rect 83181 22646 83245 22670
rect 91819 22704 91883 22712
rect 91819 22670 91836 22704
rect 91836 22670 91870 22704
rect 91870 22670 91883 22704
rect 91819 22648 91883 22670
rect 92781 22704 92845 22714
rect 92781 22670 92796 22704
rect 92796 22670 92830 22704
rect 92830 22670 92845 22704
rect 92781 22650 92845 22670
rect 40383 22450 40511 22578
rect 51940 22469 52058 22587
rect 63860 22464 63978 22582
rect 72435 22460 72553 22578
rect 104393 22557 104511 22675
rect 107979 22576 108097 22694
rect 82256 22404 82374 22522
rect 91882 22410 92000 22528
rect 105740 22331 105804 22338
rect 105740 22297 105759 22331
rect 105759 22297 105793 22331
rect 105793 22297 105804 22331
rect 105740 22274 105804 22297
rect 106706 22331 106770 22339
rect 106706 22297 106719 22331
rect 106719 22297 106753 22331
rect 106753 22297 106770 22331
rect 106706 22275 106770 22297
rect 58216 22103 58334 22221
rect 63203 22103 63321 22221
rect 105796 22028 105924 22156
rect 36843 21755 36971 21883
rect 47795 21719 47923 21847
rect 60239 21753 60357 21871
rect 36789 21569 36853 21586
rect 36789 21535 36809 21569
rect 36809 21535 36843 21569
rect 36843 21535 36853 21569
rect 36789 21522 36853 21535
rect 37758 21569 37822 21587
rect 37758 21535 37769 21569
rect 37769 21535 37803 21569
rect 37803 21535 37822 21569
rect 37758 21523 37822 21535
rect 43434 21534 43562 21662
rect 47739 21562 47803 21582
rect 47739 21528 47752 21562
rect 47752 21528 47786 21562
rect 47786 21528 47803 21562
rect 47739 21518 47803 21528
rect 48702 21562 48766 21583
rect 48702 21528 48712 21562
rect 48712 21528 48746 21562
rect 48746 21528 48766 21562
rect 48702 21519 48766 21528
rect 60257 21562 60321 21584
rect 60257 21528 60272 21562
rect 60272 21528 60306 21562
rect 60306 21528 60321 21562
rect 60257 21520 60321 21528
rect 61219 21562 61283 21583
rect 61219 21528 61232 21562
rect 61232 21528 61266 21562
rect 61266 21528 61283 21562
rect 61219 21519 61283 21528
rect 43411 21382 43475 21403
rect 43411 21348 43427 21382
rect 43427 21348 43461 21382
rect 43461 21348 43475 21382
rect 43411 21339 43475 21348
rect 44371 21382 44435 21403
rect 44371 21348 44387 21382
rect 44387 21348 44421 21382
rect 44421 21348 44435 21382
rect 44371 21339 44435 21348
rect 33485 20987 33613 21115
rect 38492 20990 38610 21108
rect 43018 20990 43136 21108
rect 44815 20991 44933 21109
rect 47050 21009 47168 21127
rect 53293 20995 53411 21113
rect 59555 20996 59673 21114
rect 63203 20993 63321 21111
rect 64422 20993 64540 21111
rect 36796 20758 36860 20771
rect 36796 20724 36809 20758
rect 36809 20724 36843 20758
rect 36843 20724 36860 20758
rect 36796 20707 36860 20724
rect 37755 20758 37819 20772
rect 37755 20724 37769 20758
rect 37769 20724 37803 20758
rect 37803 20724 37819 20758
rect 37755 20708 37819 20724
rect 47737 20751 47801 20767
rect 47737 20717 47752 20751
rect 47752 20717 47786 20751
rect 47786 20717 47801 20751
rect 47737 20703 47801 20717
rect 48698 20751 48762 20768
rect 48698 20717 48712 20751
rect 48712 20717 48746 20751
rect 48746 20717 48762 20751
rect 48698 20704 48762 20717
rect 60255 20751 60319 20761
rect 60255 20717 60272 20751
rect 60272 20717 60306 20751
rect 60306 20717 60319 20751
rect 60255 20697 60319 20717
rect 61219 20751 61283 20763
rect 61219 20717 61232 20751
rect 61232 20717 61266 20751
rect 61266 20717 61283 20751
rect 61219 20699 61283 20717
rect 67161 20772 67225 20795
rect 67161 20738 67183 20772
rect 67183 20738 67217 20772
rect 67217 20738 67225 20772
rect 67161 20731 67225 20738
rect 67640 20753 67758 20871
rect 67989 20772 68053 20792
rect 67989 20738 67994 20772
rect 67994 20738 68028 20772
rect 68028 20738 68053 20772
rect 67989 20728 68053 20738
rect 37638 20451 37766 20579
rect 43413 20571 43477 20583
rect 43413 20537 43427 20571
rect 43427 20537 43461 20571
rect 43461 20537 43477 20571
rect 43413 20519 43477 20537
rect 44376 20571 44440 20585
rect 44376 20537 44387 20571
rect 44387 20537 44421 20571
rect 44421 20537 44440 20571
rect 44376 20521 44440 20537
rect 48603 20449 48731 20577
rect 61061 20461 61179 20579
rect 74028 20527 74092 20545
rect 74028 20493 74056 20527
rect 74056 20493 74090 20527
rect 74090 20493 74092 20527
rect 74028 20481 74092 20493
rect 74332 20507 74450 20625
rect 74856 20527 74920 20551
rect 74856 20493 74867 20527
rect 74867 20493 74901 20527
rect 74901 20493 74920 20527
rect 74856 20487 74920 20493
rect 44260 20269 44388 20397
rect 66649 20214 66767 20332
rect 68386 20206 68504 20324
rect 38492 20048 38610 20166
rect 44815 20048 44933 20166
rect 45524 20053 45642 20171
rect 73565 19952 73683 20070
rect 75276 19975 75394 20093
rect 83768 20090 83886 20208
rect 93279 20090 93397 20208
rect 93830 20036 94036 20242
rect 36843 19757 36971 19885
rect 47791 19714 47919 19842
rect 60241 19723 60359 19841
rect 67163 19812 67227 19825
rect 67163 19778 67183 19812
rect 67183 19778 67217 19812
rect 67217 19778 67227 19812
rect 67163 19761 67227 19778
rect 67985 19812 68049 19826
rect 67985 19778 67994 19812
rect 67994 19778 68028 19812
rect 68028 19778 68049 19812
rect 67985 19762 68049 19778
rect 36796 19569 36860 19589
rect 36796 19535 36809 19569
rect 36809 19535 36843 19569
rect 36843 19535 36860 19569
rect 36796 19525 36860 19535
rect 37758 19569 37822 19593
rect 37758 19535 37769 19569
rect 37769 19535 37803 19569
rect 37803 19535 37822 19569
rect 37758 19529 37822 19535
rect 43415 19526 43543 19654
rect 47739 19562 47803 19583
rect 47739 19528 47752 19562
rect 47752 19528 47786 19562
rect 47786 19528 47803 19562
rect 47739 19519 47803 19528
rect 48695 19562 48759 19583
rect 48695 19528 48712 19562
rect 48712 19528 48746 19562
rect 48746 19528 48759 19562
rect 48695 19519 48759 19528
rect 60254 19562 60318 19582
rect 60254 19528 60272 19562
rect 60272 19528 60306 19562
rect 60306 19528 60318 19562
rect 60254 19518 60318 19528
rect 61219 19562 61283 19583
rect 61219 19528 61232 19562
rect 61232 19528 61266 19562
rect 61266 19528 61283 19562
rect 61219 19519 61283 19528
rect 67637 19527 67755 19645
rect 74034 19567 74098 19583
rect 74034 19533 74056 19567
rect 74056 19533 74090 19567
rect 74090 19533 74098 19567
rect 74034 19519 74098 19533
rect 74860 19567 74924 19582
rect 74860 19533 74867 19567
rect 74867 19533 74901 19567
rect 74901 19533 74924 19567
rect 74860 19518 74924 19533
rect 43407 19382 43471 19402
rect 43407 19348 43427 19382
rect 43427 19348 43461 19382
rect 43461 19348 43471 19382
rect 43407 19338 43471 19348
rect 44367 19382 44431 19399
rect 44367 19348 44387 19382
rect 44387 19348 44421 19382
rect 44421 19348 44431 19382
rect 44367 19335 44431 19348
rect 74330 19293 74448 19411
rect 35205 19010 35323 19128
rect 38492 19000 38610 19118
rect 42143 18998 42261 19116
rect 43009 18998 43127 19116
rect 44815 18991 44933 19109
rect 46206 19025 46324 19143
rect 53306 18994 53424 19112
rect 56914 18995 57032 19113
rect 63210 18994 63328 19112
rect 65692 18994 65810 19112
rect 36796 18758 36860 18772
rect 36796 18724 36809 18758
rect 36809 18724 36843 18758
rect 36843 18724 36860 18758
rect 36796 18708 36860 18724
rect 37756 18758 37820 18771
rect 37756 18724 37769 18758
rect 37769 18724 37803 18758
rect 37803 18724 37820 18758
rect 37756 18707 37820 18724
rect 47737 18751 47801 18761
rect 47737 18717 47752 18751
rect 47752 18717 47786 18751
rect 47786 18717 47801 18751
rect 47737 18697 47801 18717
rect 48697 18751 48761 18760
rect 48697 18717 48712 18751
rect 48712 18717 48746 18751
rect 48746 18717 48761 18751
rect 48697 18696 48761 18717
rect 60257 18751 60321 18763
rect 60257 18717 60272 18751
rect 60272 18717 60306 18751
rect 60306 18717 60321 18751
rect 60257 18699 60321 18717
rect 61221 18751 61285 18765
rect 61221 18717 61232 18751
rect 61232 18717 61266 18751
rect 61266 18717 61285 18751
rect 61221 18701 61285 18717
rect 87767 18719 87885 18837
rect 88626 18719 88744 18837
rect 95000 18719 95118 18837
rect 37633 18450 37761 18578
rect 43411 18571 43475 18582
rect 43411 18537 43427 18571
rect 43427 18537 43461 18571
rect 43461 18537 43475 18571
rect 43411 18518 43475 18537
rect 44372 18571 44436 18581
rect 44372 18537 44387 18571
rect 44387 18537 44421 18571
rect 44421 18537 44436 18571
rect 44372 18517 44436 18537
rect 48603 18450 48731 18578
rect 61055 18465 61173 18583
rect 44259 18261 44387 18389
rect 53306 17971 53424 18089
rect 54501 17971 54619 18089
rect 55642 18050 55760 18168
rect 63210 18050 63328 18168
rect 40397 17738 40525 17866
rect 51104 17722 51222 17840
rect 63015 17715 63133 17833
rect 71584 17726 71702 17844
rect 82968 17695 83086 17813
rect 92566 17701 92684 17819
rect 40367 17567 40431 17587
rect 40367 17533 40384 17567
rect 40384 17533 40418 17567
rect 40418 17533 40431 17567
rect 40367 17523 40431 17533
rect 41333 17567 41397 17586
rect 41333 17533 41344 17567
rect 41344 17533 41378 17567
rect 41378 17533 41397 17567
rect 41333 17522 41397 17533
rect 51044 17562 51108 17582
rect 51044 17528 51062 17562
rect 51062 17528 51096 17562
rect 51096 17528 51108 17562
rect 51044 17518 51108 17528
rect 52011 17562 52075 17583
rect 52011 17528 52022 17562
rect 52022 17528 52056 17562
rect 52056 17528 52075 17562
rect 52011 17519 52075 17528
rect 62980 17562 63044 17581
rect 62980 17528 62992 17562
rect 62992 17528 63026 17562
rect 63026 17528 63044 17562
rect 62980 17517 63044 17528
rect 63942 17562 64006 17582
rect 63942 17528 63952 17562
rect 63952 17528 63986 17562
rect 63986 17528 64006 17562
rect 63942 17518 64006 17528
rect 71543 17573 71607 17593
rect 71543 17539 71556 17573
rect 71556 17539 71590 17573
rect 71590 17539 71607 17573
rect 71543 17529 71607 17539
rect 72501 17573 72565 17594
rect 72501 17539 72516 17573
rect 72516 17539 72550 17573
rect 72550 17539 72565 17573
rect 72501 17530 72565 17539
rect 82223 17545 82287 17567
rect 82223 17511 82235 17545
rect 82235 17511 82269 17545
rect 82269 17511 82287 17545
rect 82223 17503 82287 17511
rect 83186 17545 83250 17567
rect 83186 17511 83195 17545
rect 83195 17511 83229 17545
rect 83229 17511 83250 17545
rect 83186 17503 83250 17511
rect 91828 17545 91892 17567
rect 91828 17511 91836 17545
rect 91836 17511 91870 17545
rect 91870 17511 91892 17545
rect 91828 17503 91892 17511
rect 92780 17545 92844 17565
rect 92780 17511 92796 17545
rect 92796 17511 92830 17545
rect 92830 17511 92844 17545
rect 92780 17501 92844 17511
rect 83768 17161 83886 17279
rect 35205 16975 35323 17093
rect 43009 17009 43127 17127
rect 47050 16997 47168 17115
rect 53306 16991 53424 17109
rect 56914 17039 57032 17157
rect 88626 17155 88744 17273
rect 93279 17156 93397 17274
rect 64422 16994 64540 17112
rect 67638 16995 67756 17113
rect 69638 16958 69766 17086
rect 74330 17005 74448 17123
rect 77953 17003 78071 17121
rect 80129 17006 80247 17124
rect 81510 17005 81628 17123
rect 86412 16844 86530 16962
rect 40370 16756 40434 16765
rect 40370 16722 40384 16756
rect 40384 16722 40418 16756
rect 40418 16722 40434 16756
rect 40370 16701 40434 16722
rect 41328 16756 41392 16762
rect 41328 16722 41344 16756
rect 41344 16722 41378 16756
rect 41378 16722 41392 16756
rect 41328 16698 41392 16722
rect 51048 16751 51112 16760
rect 51048 16717 51062 16751
rect 51062 16717 51096 16751
rect 51096 16717 51112 16751
rect 51048 16696 51112 16717
rect 52008 16751 52072 16760
rect 52008 16717 52022 16751
rect 52022 16717 52056 16751
rect 52056 16717 52072 16751
rect 52008 16696 52072 16717
rect 62978 16751 63042 16762
rect 62978 16717 62992 16751
rect 62992 16717 63026 16751
rect 63026 16717 63042 16751
rect 62978 16698 63042 16717
rect 63938 16751 64002 16763
rect 63938 16717 63952 16751
rect 63952 16717 63986 16751
rect 63986 16717 64002 16751
rect 63938 16699 64002 16717
rect 71544 16762 71608 16774
rect 71544 16728 71556 16762
rect 71556 16728 71590 16762
rect 71590 16728 71608 16762
rect 71544 16710 71608 16728
rect 72505 16762 72569 16775
rect 72505 16728 72516 16762
rect 72516 16728 72550 16762
rect 72550 16728 72569 16762
rect 72505 16711 72569 16728
rect 82220 16734 82284 16742
rect 82220 16700 82235 16734
rect 82235 16700 82269 16734
rect 82269 16700 82284 16734
rect 82220 16678 82284 16700
rect 83186 16734 83250 16742
rect 83186 16700 83195 16734
rect 83195 16700 83229 16734
rect 83229 16700 83250 16734
rect 83186 16678 83250 16700
rect 85579 16695 85643 16717
rect 85579 16661 85595 16695
rect 85595 16661 85629 16695
rect 85629 16661 85643 16695
rect 85579 16653 85643 16661
rect 86542 16695 86606 16719
rect 86542 16661 86555 16695
rect 86555 16661 86589 16695
rect 86589 16661 86606 16695
rect 86542 16655 86606 16661
rect 91823 16734 91887 16742
rect 91823 16700 91836 16734
rect 91836 16700 91870 16734
rect 91870 16700 91887 16734
rect 91823 16678 91887 16700
rect 92781 16734 92845 16745
rect 92781 16700 92796 16734
rect 92796 16700 92830 16734
rect 92830 16700 92845 16734
rect 92781 16681 92845 16700
rect 41211 16414 41339 16542
rect 51817 16464 51935 16582
rect 63827 16455 63945 16573
rect 72296 16464 72414 16582
rect 82296 16443 82414 16561
rect 91859 16429 91977 16547
rect 81510 16261 81628 16379
rect 88626 16305 88744 16423
rect 85579 15884 85643 15893
rect 85579 15850 85595 15884
rect 85595 15850 85629 15884
rect 85629 15850 85643 15884
rect 85579 15829 85643 15850
rect 86541 15884 86605 15891
rect 86541 15850 86555 15884
rect 86555 15850 86589 15884
rect 86589 15850 86605 15884
rect 86541 15827 86605 15850
rect 85624 15577 85742 15695
rect 135402 -36 135875 33
rect 133777 -159 133829 -151
rect 133777 -193 133786 -159
rect 133786 -193 133820 -159
rect 133820 -193 133829 -159
rect 133777 -203 133829 -193
rect 133151 -279 133217 -264
rect 133151 -330 133157 -279
rect 133157 -330 133211 -279
rect 133211 -330 133217 -279
rect 133151 -332 133217 -330
rect 133290 -279 133356 -272
rect 133290 -330 133296 -279
rect 133296 -330 133350 -279
rect 133350 -330 133356 -279
rect 133290 -340 133356 -330
rect 134067 -220 134133 -214
rect 134067 -271 134074 -220
rect 134074 -271 134128 -220
rect 134128 -271 134133 -220
rect 134067 -282 134133 -271
rect 134200 -218 134266 -216
rect 134200 -269 134205 -218
rect 134205 -269 134259 -218
rect 134259 -269 134266 -218
rect 134200 -284 134266 -269
rect 134345 -291 134397 -274
rect 134345 -325 134350 -291
rect 134350 -325 134384 -291
rect 134384 -325 134397 -291
rect 134345 -326 134397 -325
rect 141783 -244 141835 -192
rect 139082 -577 139544 -513
rect 135405 -1351 135878 -1282
rect 133777 -1476 133829 -1468
rect 133777 -1510 133786 -1476
rect 133786 -1510 133820 -1476
rect 133820 -1510 133829 -1476
rect 133777 -1520 133829 -1510
rect 133151 -1596 133217 -1581
rect 133151 -1647 133157 -1596
rect 133157 -1647 133211 -1596
rect 133211 -1647 133217 -1596
rect 133151 -1649 133217 -1647
rect 133290 -1596 133356 -1589
rect 133290 -1647 133296 -1596
rect 133296 -1647 133350 -1596
rect 133350 -1647 133356 -1596
rect 133290 -1657 133356 -1647
rect 134067 -1537 134133 -1531
rect 134067 -1588 134074 -1537
rect 134074 -1588 134128 -1537
rect 134128 -1588 134133 -1537
rect 134067 -1599 134133 -1588
rect 134200 -1535 134266 -1533
rect 134200 -1586 134205 -1535
rect 134205 -1586 134259 -1535
rect 134259 -1586 134266 -1535
rect 134200 -1601 134266 -1586
rect 134345 -1608 134397 -1591
rect 134345 -1642 134350 -1608
rect 134350 -1642 134384 -1608
rect 134384 -1642 134397 -1608
rect 134345 -1643 134397 -1642
rect 141783 -1561 141835 -1509
rect 66754 -1970 66882 -1842
rect 139092 -1891 139554 -1827
rect 67103 -2665 67170 -2039
rect 71868 -2165 71996 -2037
rect 72410 -2172 72538 -2044
rect 72954 -2175 73082 -2047
rect 73498 -2176 73626 -2048
rect 75124 -2164 75252 -2036
rect 75669 -2159 75797 -2031
rect 76211 -2161 76339 -2033
rect 76758 -2161 76886 -2033
rect 79476 -2157 79604 -2029
rect 80020 -2159 80148 -2031
rect 80563 -2157 80691 -2029
rect 81106 -2159 81234 -2031
rect 82749 -2150 82877 -2022
rect 83289 -2155 83417 -2027
rect 83830 -2157 83958 -2029
rect 84370 -2150 84498 -2022
rect 135397 -2997 135870 -2928
rect 133777 -3123 133829 -3115
rect 133777 -3157 133786 -3123
rect 133786 -3157 133820 -3123
rect 133820 -3157 133829 -3123
rect 133777 -3167 133829 -3157
rect 133151 -3243 133217 -3228
rect 133151 -3294 133157 -3243
rect 133157 -3294 133211 -3243
rect 133211 -3294 133217 -3243
rect 133151 -3296 133217 -3294
rect 133290 -3243 133356 -3236
rect 133290 -3294 133296 -3243
rect 133296 -3294 133350 -3243
rect 133350 -3294 133356 -3243
rect 133290 -3304 133356 -3294
rect 134067 -3184 134133 -3178
rect 134067 -3235 134074 -3184
rect 134074 -3235 134128 -3184
rect 134128 -3235 134133 -3184
rect 134067 -3246 134133 -3235
rect 134200 -3182 134266 -3180
rect 134200 -3233 134205 -3182
rect 134205 -3233 134259 -3182
rect 134259 -3233 134266 -3182
rect 134200 -3248 134266 -3233
rect 134345 -3255 134397 -3238
rect 134345 -3289 134350 -3255
rect 134350 -3289 134384 -3255
rect 134384 -3289 134397 -3255
rect 134345 -3290 134397 -3289
rect 141783 -3208 141835 -3156
rect 139082 -3541 139544 -3477
rect 135399 -4247 135872 -4178
rect 133777 -4370 133829 -4362
rect 133777 -4404 133786 -4370
rect 133786 -4404 133820 -4370
rect 133820 -4404 133829 -4370
rect 133777 -4414 133829 -4404
rect 133151 -4490 133217 -4475
rect 133151 -4541 133157 -4490
rect 133157 -4541 133211 -4490
rect 133211 -4541 133217 -4490
rect 133151 -4543 133217 -4541
rect 133290 -4490 133356 -4483
rect 133290 -4541 133296 -4490
rect 133296 -4541 133350 -4490
rect 133350 -4541 133356 -4490
rect 133290 -4551 133356 -4541
rect 134067 -4431 134133 -4425
rect 134067 -4482 134074 -4431
rect 134074 -4482 134128 -4431
rect 134128 -4482 134133 -4431
rect 134067 -4493 134133 -4482
rect 134200 -4429 134266 -4427
rect 134200 -4480 134205 -4429
rect 134205 -4480 134259 -4429
rect 134259 -4480 134266 -4429
rect 134200 -4495 134266 -4480
rect 134345 -4502 134397 -4485
rect 134345 -4536 134350 -4502
rect 134350 -4536 134384 -4502
rect 134384 -4536 134397 -4502
rect 134345 -4537 134397 -4536
rect 141783 -4455 141835 -4403
rect 139097 -4788 139559 -4724
rect 66560 -6253 66627 -5627
rect 71081 -6267 71140 -5629
rect 74345 -6267 74404 -5629
rect 77609 -6267 77668 -5629
rect 78697 -6267 78756 -5629
rect 81961 -6267 82020 -5629
rect 85225 -6267 85284 -5629
rect 66846 -6811 66974 -6683
rect 71628 -9265 71687 -8627
rect 72716 -9265 72775 -8627
rect 73804 -9265 73863 -8627
rect 74892 -9265 74951 -8627
rect 75980 -9265 76039 -8627
rect 77068 -9265 77127 -8627
rect 78156 -9265 78215 -8627
rect 79244 -9265 79303 -8627
rect 80332 -9265 80391 -8627
rect 81420 -9265 81479 -8627
rect 82508 -9265 82567 -8627
rect 83596 -9265 83655 -8627
rect 84684 -9265 84743 -8627
rect 147329 -11225 147802 -11156
rect 145709 -11351 145761 -11343
rect 145709 -11385 145718 -11351
rect 145718 -11385 145752 -11351
rect 145752 -11385 145761 -11351
rect 145709 -11395 145761 -11385
rect 145083 -11471 145149 -11456
rect 145083 -11522 145089 -11471
rect 145089 -11522 145143 -11471
rect 145143 -11522 145149 -11471
rect 145083 -11524 145149 -11522
rect 145222 -11471 145288 -11464
rect 145222 -11522 145228 -11471
rect 145228 -11522 145282 -11471
rect 145282 -11522 145288 -11471
rect 145222 -11532 145288 -11522
rect 145999 -11412 146065 -11406
rect 145999 -11463 146006 -11412
rect 146006 -11463 146060 -11412
rect 146060 -11463 146065 -11412
rect 145999 -11474 146065 -11463
rect 146132 -11410 146198 -11408
rect 146132 -11461 146137 -11410
rect 146137 -11461 146191 -11410
rect 146191 -11461 146198 -11410
rect 146132 -11476 146198 -11461
rect 146277 -11483 146329 -11466
rect 146277 -11517 146282 -11483
rect 146282 -11517 146316 -11483
rect 146316 -11517 146329 -11483
rect 146277 -11518 146329 -11517
rect 153848 -11436 153900 -11384
rect 151014 -11769 151476 -11705
rect 71079 -14265 71138 -13627
rect 72167 -14265 72226 -13627
rect 73255 -14265 73314 -13627
rect 74343 -14265 74402 -13627
rect 75431 -14265 75490 -13627
rect 76519 -14265 76578 -13627
rect 77607 -14265 77666 -13627
rect 78695 -14265 78754 -13627
rect 79783 -14265 79842 -13627
rect 80871 -14265 80930 -13627
rect 81959 -14265 82018 -13627
rect 83047 -14265 83106 -13627
rect 84135 -14265 84194 -13627
rect 85223 -14265 85282 -13627
rect 71621 -17271 71685 -16617
rect 72709 -17271 72773 -16617
rect 73797 -17271 73861 -16617
rect 74885 -17271 74949 -16617
rect 75973 -17271 76037 -16617
rect 77061 -17271 77125 -16617
rect 78149 -17271 78213 -16617
rect 79237 -17271 79301 -16617
rect 80325 -17271 80389 -16617
rect 81413 -17271 81477 -16617
rect 82501 -17271 82565 -16617
rect 83589 -17271 83653 -16617
rect 84677 -17271 84741 -16617
rect 71075 -22006 71142 -21612
rect 72165 -22012 72232 -21618
rect 73253 -22012 73320 -21618
rect 74341 -22012 74408 -21618
rect 75429 -22012 75496 -21618
rect 76517 -22012 76584 -21618
rect 77605 -22012 77672 -21618
rect 81957 -22012 82024 -21618
rect 83045 -22012 83112 -21618
rect 84133 -22012 84200 -21618
rect 85221 -22012 85288 -21618
rect 77491 -23175 78491 -22175
<< metal2 >>
rect 103391 71867 104426 71889
rect 36373 71835 37373 71844
rect 36373 70826 37373 70835
rect 43351 71817 44375 71828
rect 43351 70817 43364 71817
rect 44364 70817 44375 71817
rect 43351 70806 44375 70817
rect 57794 71821 58825 71840
rect 57794 70821 57809 71821
rect 58809 70821 58825 71821
rect 74871 71807 75895 71820
rect 57794 70802 58825 70821
rect 64867 71771 65896 71786
rect 64867 70771 64881 71771
rect 65881 70771 65896 71771
rect 74871 70807 74883 71807
rect 75883 70807 75895 71807
rect 94051 71783 95086 71805
rect 74871 70796 75895 70807
rect 85741 71759 86776 71781
rect 64867 70758 65896 70771
rect 85741 70759 85758 71759
rect 86758 70759 86776 71759
rect 94051 70783 94068 71783
rect 95068 70783 95086 71783
rect 103391 70867 103408 71867
rect 104408 70867 104426 71867
rect 103391 70852 104426 70867
rect 94051 70768 95086 70783
rect 85741 70744 86776 70759
rect 35285 70423 35410 70433
rect 45277 70421 45431 70431
rect 35285 67097 35410 67107
rect 38294 70399 38442 70409
rect 38294 67103 38442 67113
rect 42295 70392 42410 70402
rect 42295 67100 42410 67110
rect 56700 70393 56848 70403
rect 56700 67103 56848 67113
rect 59712 70398 59864 70408
rect 59712 67103 59864 67113
rect 63788 70396 63951 70406
rect 66804 70395 66952 70405
rect 66804 67107 66952 67117
rect 73794 70398 73935 70408
rect 87663 70406 87817 70416
rect 63788 67095 63951 67105
rect 73794 67097 73935 67107
rect 76799 70396 76934 70406
rect 76799 67103 76934 67113
rect 84670 70393 84798 70403
rect 84670 67102 84798 67112
rect 87663 67098 87817 67108
rect 92977 70406 93119 70416
rect 95985 70403 96113 70413
rect 95985 67102 96113 67112
rect 102317 70406 102459 70416
rect 45277 67082 45431 67092
rect 92977 67090 93119 67100
rect 105325 70403 105453 70413
rect 105325 67102 105453 67112
rect 102317 67090 102459 67100
rect 36789 66748 36795 66876
rect 36923 66748 36929 66876
rect 36795 56295 36923 66748
rect 43789 66688 43795 66816
rect 43923 66688 43929 66816
rect 58209 66778 58215 66906
rect 58343 66778 58349 66906
rect 65309 66804 65315 66932
rect 65443 66804 65449 66932
rect 75309 66831 75315 66959
rect 75443 66831 75449 66959
rect 43795 57231 43923 66688
rect 38703 57103 38709 57231
rect 38837 57103 38843 57231
rect 43789 57103 43795 57231
rect 43923 57103 43929 57231
rect 36789 56167 36795 56295
rect 36923 56167 36929 56295
rect 36795 50626 36923 56167
rect 36406 50593 36466 50602
rect 36406 50524 36466 50533
rect 36408 50263 36464 50524
rect 38709 50628 38837 57103
rect 48935 53843 48941 53961
rect 49059 53843 49065 53961
rect 46449 52636 46509 52645
rect 46153 52282 46271 52292
rect 46153 51685 46271 51695
rect 46449 52265 46509 52576
rect 48449 52633 48509 52642
rect 46449 51302 46509 52205
rect 47271 52276 47341 52281
rect 47271 52271 47343 52276
rect 47341 52201 47343 52271
rect 48449 52275 48509 52573
rect 48941 52517 49059 53843
rect 48941 52393 49059 52399
rect 47271 52191 47343 52201
rect 47273 51320 47343 52191
rect 48197 52230 48307 52240
rect 47272 51310 47343 51320
rect 46449 51232 46509 51242
rect 46751 51281 46879 51287
rect 36795 50492 36923 50498
rect 38404 50595 38464 50604
rect 37447 50285 37567 50295
rect 36202 49927 36285 49937
rect 36202 49473 36285 49483
rect 36408 49304 36464 50207
rect 37227 50271 37288 50281
rect 37227 50211 37228 50271
rect 37227 50201 37288 50211
rect 36408 49238 36464 49248
rect 36693 49338 36821 49348
rect 36693 48424 36821 49210
rect 37227 49309 37287 50201
rect 38404 50269 38464 50535
rect 38709 50494 38837 50500
rect 47342 51240 47343 51310
rect 47272 51230 47343 51240
rect 39493 50313 39608 50323
rect 37447 49782 37567 49792
rect 38144 49857 38243 49867
rect 38144 49268 38243 49278
rect 38404 49318 38464 50209
rect 39227 50265 39287 50277
rect 38692 49353 38820 49363
rect 38404 49308 38465 49318
rect 37227 49027 37287 49249
rect 38404 49248 38405 49308
rect 38404 49247 38465 49248
rect 38405 49238 38465 49247
rect 37227 48958 37287 48967
rect 36687 48296 36693 48424
rect 36821 48296 36827 48424
rect 36693 40605 36821 48296
rect 38692 47294 38820 49225
rect 39227 49307 39287 50205
rect 39493 49770 39608 49780
rect 39227 49016 39287 49247
rect 39227 48947 39287 48956
rect 46751 48424 46879 51153
rect 47273 50892 47343 51230
rect 47493 51852 47608 51862
rect 48197 51680 48307 51690
rect 48449 51323 48509 52215
rect 49271 52285 49331 52290
rect 49271 52275 49334 52285
rect 49271 52215 49274 52275
rect 49271 52205 49334 52215
rect 49271 51325 49331 52205
rect 49511 51907 49654 51917
rect 48449 51313 48510 51323
rect 48449 51253 48450 51313
rect 49271 51315 49336 51325
rect 48449 51247 48510 51253
rect 48450 51243 48510 51247
rect 48730 51289 48873 51297
rect 47493 51219 47608 51229
rect 48730 51161 48737 51289
rect 48865 51161 48873 51289
rect 48730 51154 48873 51161
rect 49271 51255 49276 51315
rect 49271 51245 49336 51255
rect 58215 51393 58343 66778
rect 65315 65373 65443 66804
rect 65315 65239 65443 65245
rect 75315 65373 75443 66831
rect 86179 66785 86185 66913
rect 86313 66785 86319 66913
rect 75315 65239 75443 65245
rect 63684 65102 63797 65112
rect 62908 65047 63133 65057
rect 62908 64970 63133 64980
rect 65058 65111 65171 65121
rect 63684 64979 63797 64989
rect 64232 65055 64460 65065
rect 66421 65111 66534 65121
rect 65058 64988 65171 64998
rect 65616 65055 65843 65065
rect 64232 64966 64460 64976
rect 67770 65112 67883 65122
rect 66421 64988 66534 64998
rect 66997 65054 67225 65064
rect 65616 64970 65843 64980
rect 73684 65102 73797 65112
rect 67770 64989 67883 64999
rect 72908 65047 73133 65057
rect 66997 64972 67225 64982
rect 72908 64970 73133 64980
rect 75058 65111 75171 65121
rect 73684 64979 73797 64989
rect 74232 65055 74460 65065
rect 76421 65111 76534 65121
rect 75058 64988 75171 64998
rect 75616 65055 75843 65065
rect 74232 64966 74460 64976
rect 77770 65112 77883 65122
rect 76421 64988 76534 64998
rect 76997 65054 77225 65064
rect 75616 64970 75843 64980
rect 77770 64989 77883 64999
rect 76997 64972 77225 64982
rect 61524 64144 61642 64153
rect 60896 62929 61014 62934
rect 60892 62821 60901 62929
rect 61009 62821 61018 62929
rect 60896 60424 61014 62821
rect 61524 60755 61642 64026
rect 71637 64136 71755 64145
rect 84175 64129 84293 64134
rect 84171 64021 84180 64129
rect 84288 64021 84297 64129
rect 86185 64108 86313 66785
rect 94489 66623 94495 66751
rect 94623 66623 94629 66751
rect 103829 66742 103835 66870
rect 103963 66742 103969 66870
rect 62129 63540 62247 63549
rect 62129 60994 62247 63422
rect 71105 62929 71223 62934
rect 71101 62821 71110 62929
rect 71218 62821 71227 62929
rect 62731 62189 62844 62199
rect 64721 62177 64834 62187
rect 64378 62159 64491 62169
rect 62731 62066 62844 62076
rect 63429 62146 63542 62156
rect 64721 62054 64834 62064
rect 65456 62169 65569 62179
rect 65456 62046 65569 62056
rect 66175 62151 66288 62161
rect 64378 62035 64491 62045
rect 63429 62023 63542 62033
rect 66175 62028 66288 62038
rect 66828 62143 66941 62153
rect 66828 62020 66941 62030
rect 67543 62151 67656 62161
rect 67543 62028 67656 62038
rect 65884 61473 65952 61483
rect 63163 61352 63234 61362
rect 63163 61235 63234 61245
rect 63705 61346 63776 61356
rect 66971 61383 67043 61393
rect 63705 61232 63776 61242
rect 64251 61330 64320 61340
rect 65884 61339 65952 61349
rect 66426 61364 66494 61374
rect 64251 61174 64320 61184
rect 64798 61321 64862 61331
rect 66971 61251 67043 61261
rect 67514 61356 67580 61366
rect 66426 61197 66494 61207
rect 67514 61192 67580 61202
rect 64798 61181 64862 61191
rect 65343 61015 65410 61025
rect 62129 60876 62625 60994
rect 65343 60852 65410 60862
rect 61524 60637 62754 60755
rect 71105 60447 71223 62821
rect 71637 60771 71755 64018
rect 72122 63539 72240 63548
rect 72122 60986 72240 63421
rect 72731 62189 72844 62199
rect 74721 62177 74834 62187
rect 74378 62159 74491 62169
rect 72731 62066 72844 62076
rect 73429 62146 73542 62156
rect 74721 62054 74834 62064
rect 75456 62169 75569 62179
rect 75456 62046 75569 62056
rect 76175 62151 76288 62161
rect 74378 62035 74491 62045
rect 73429 62023 73542 62033
rect 76175 62028 76288 62038
rect 76828 62143 76941 62153
rect 76828 62020 76941 62030
rect 77543 62151 77656 62161
rect 77543 62028 77656 62038
rect 75884 61473 75952 61483
rect 73163 61352 73234 61362
rect 73163 61235 73234 61245
rect 73705 61346 73776 61356
rect 76971 61383 77043 61393
rect 73705 61232 73776 61242
rect 74251 61330 74320 61340
rect 75884 61339 75952 61349
rect 76426 61364 76494 61374
rect 74251 61174 74320 61184
rect 74798 61321 74862 61331
rect 76971 61251 77043 61261
rect 77514 61356 77580 61366
rect 76426 61197 76494 61207
rect 77514 61192 77580 61202
rect 74798 61181 74862 61191
rect 75343 61015 75410 61025
rect 72122 60868 72682 60986
rect 75343 60852 75410 60862
rect 71637 60653 72671 60771
rect 60896 60306 62699 60424
rect 71105 60329 72652 60447
rect 84175 60403 84293 64021
rect 86185 63974 86313 63980
rect 85128 63849 85318 63859
rect 86485 63858 86629 63868
rect 85128 63747 85318 63757
rect 85568 63823 86002 63833
rect 86485 63754 86629 63764
rect 86904 63809 87328 63819
rect 85568 63726 86002 63736
rect 86904 63722 87328 63732
rect 88033 62929 88151 62934
rect 88029 62821 88038 62929
rect 88146 62821 88155 62929
rect 85219 62346 85311 62356
rect 85219 62227 85311 62237
rect 86550 62341 86642 62351
rect 86550 62222 86642 62232
rect 86094 60499 86159 60509
rect 84175 60285 84991 60403
rect 88033 60412 88151 62821
rect 86094 60347 86159 60357
rect 87327 60294 88151 60412
rect 85544 60274 85615 60284
rect 85544 60160 85615 60170
rect 86636 60280 86704 60290
rect 86636 60160 86704 60170
rect 63052 59993 63305 60003
rect 63052 59906 63305 59916
rect 64372 60000 64680 60010
rect 64372 59905 64680 59915
rect 65760 59989 66042 59999
rect 65760 59908 66042 59918
rect 67132 59991 67414 60001
rect 67132 59910 67414 59920
rect 73052 59993 73305 60003
rect 73052 59906 73305 59916
rect 74372 60000 74680 60010
rect 74372 59905 74680 59915
rect 75760 59989 76042 59999
rect 75760 59908 76042 59918
rect 77132 59991 77414 60001
rect 77132 59910 77414 59920
rect 84943 59636 85056 59646
rect 84943 59513 85056 59523
rect 68044 59416 68157 59426
rect 66660 59381 66773 59391
rect 65298 59363 65411 59373
rect 63937 59351 64050 59361
rect 78044 59416 78157 59426
rect 76660 59381 76773 59391
rect 75298 59363 75411 59373
rect 68044 59293 68157 59303
rect 73937 59351 74050 59361
rect 66660 59258 66773 59268
rect 65298 59240 65411 59250
rect 63937 59228 64050 59238
rect 78044 59293 78157 59303
rect 76660 59258 76773 59268
rect 75298 59240 75411 59250
rect 73937 59228 74050 59238
rect 87336 59030 87449 59040
rect 87336 58907 87449 58917
rect 73366 58714 73513 58723
rect 63312 58701 63518 58707
rect 64700 58578 64706 58709
rect 64837 58578 64843 58709
rect 58756 57830 58762 57890
rect 58822 57830 58828 57890
rect 58762 52159 58822 57830
rect 61618 55604 61749 55610
rect 58755 52103 58764 52159
rect 58820 52103 58829 52159
rect 58762 52101 58822 52103
rect 61618 51650 61749 55473
rect 62492 54651 62501 54768
rect 62618 54651 62627 54768
rect 62501 51663 62618 54651
rect 63312 52174 63518 58495
rect 64706 55604 64837 58578
rect 66027 58507 66033 58713
rect 66239 58507 66245 58713
rect 73366 58578 73373 58714
rect 73504 58578 73513 58714
rect 74715 58593 74721 58710
rect 74838 58593 74844 58710
rect 76105 58685 76165 58691
rect 73366 58563 73513 58578
rect 64700 55473 64706 55604
rect 64837 55473 64843 55604
rect 63312 51978 63317 52174
rect 63513 51978 63518 52174
rect 63312 51973 63518 51978
rect 63317 51969 63513 51973
rect 66033 51678 66239 58507
rect 61614 51529 61623 51650
rect 61744 51529 61753 51650
rect 62497 51556 62506 51663
rect 62613 51556 62622 51663
rect 62501 51551 62618 51556
rect 61618 51524 61749 51529
rect 66029 51482 66038 51678
rect 66234 51482 66243 51678
rect 66033 51477 66239 51482
rect 58209 51265 58215 51393
rect 58343 51265 58349 51393
rect 47273 50813 47343 50822
rect 46745 48296 46751 48424
rect 46879 48296 46885 48424
rect 38680 47288 38820 47294
rect 48737 47288 48865 51154
rect 49271 50890 49331 51245
rect 49511 51239 49654 51249
rect 73373 51121 73504 58563
rect 74721 54763 74838 58593
rect 76105 57890 76165 58625
rect 85384 58196 85512 58202
rect 76099 57830 76105 57890
rect 76165 57830 76171 57890
rect 82641 57103 82647 57231
rect 82775 57103 82781 57231
rect 80619 56167 80625 56295
rect 80753 56167 80759 56295
rect 78620 55566 78748 55575
rect 78614 55438 78620 55566
rect 78748 55438 78754 55566
rect 74717 54656 74726 54763
rect 74833 54656 74842 54763
rect 74721 54651 74838 54656
rect 73373 50984 73504 50990
rect 49271 50821 49331 50830
rect 61618 50387 61749 50396
rect 61618 48842 61749 50256
rect 67970 50219 68198 50229
rect 66174 50207 66362 50217
rect 66174 50003 66362 50013
rect 71483 50211 71711 50221
rect 67970 49977 68198 49987
rect 69664 50200 69892 50210
rect 71483 49969 71711 49979
rect 73267 50208 73495 50218
rect 69664 49958 69892 49968
rect 73267 49966 73495 49976
rect 75052 50206 75280 50216
rect 75052 49964 75280 49974
rect 62848 49622 63380 49632
rect 62848 49455 63380 49465
rect 67154 48662 67390 48672
rect 65284 48632 65560 48642
rect 67154 48574 67390 48584
rect 68959 48655 69193 48665
rect 68959 48566 69193 48576
rect 70765 48651 70984 48661
rect 70765 48560 70984 48570
rect 72551 48655 72791 48665
rect 74352 48651 74604 48661
rect 74352 48576 74604 48586
rect 72551 48561 72791 48571
rect 65284 48522 65560 48532
rect 56046 47379 56330 47389
rect 38808 47160 38820 47288
rect 48731 47160 48737 47288
rect 48865 47160 48871 47288
rect 38680 47154 38820 47160
rect 38692 45557 38820 47154
rect 60492 47309 61496 47319
rect 61728 47276 61862 47284
rect 61728 47154 61736 47276
rect 61853 47274 61862 47276
rect 61853 47157 62501 47274
rect 62618 47157 62627 47274
rect 61853 47154 61862 47157
rect 61728 47145 61862 47154
rect 60492 47099 61496 47109
rect 56046 46731 56330 46741
rect 58762 45842 58822 45851
rect 58762 45773 58822 45782
rect 38692 45423 38820 45429
rect 44965 45557 45093 45563
rect 44965 40528 45093 45429
rect 62010 42674 62280 42684
rect 62010 41589 62280 41599
rect 62857 42671 63127 42681
rect 63412 42335 63617 42345
rect 63412 41737 63617 41747
rect 62857 41586 63127 41596
rect 36693 40468 36821 40477
rect 44956 40400 44965 40528
rect 45093 40400 45102 40528
rect 56027 39355 56167 39365
rect 56027 38721 56167 38731
rect 68833 37306 69077 37316
rect 66930 37246 67174 37256
rect 65328 37235 65572 37245
rect 68833 37096 69077 37106
rect 70550 37290 70794 37300
rect 70550 37080 70794 37090
rect 72364 37285 72608 37295
rect 72364 37075 72608 37085
rect 74336 37279 74580 37289
rect 74336 37069 74580 37079
rect 66930 37036 67174 37046
rect 65328 37025 65572 37035
rect 65850 35734 66234 35744
rect 67641 35741 68041 35751
rect 67641 35657 68041 35667
rect 69447 35741 69835 35751
rect 69447 35657 69835 35667
rect 71244 35706 71632 35716
rect 65850 35646 66234 35656
rect 71244 35622 71632 35632
rect 73046 35706 73433 35716
rect 73046 35618 73433 35628
rect 74840 35702 75235 35712
rect 74840 35615 75235 35625
rect 67546 34952 67555 35060
rect 67663 34952 67672 35060
rect 35195 34277 35323 34282
rect 35191 34159 35200 34277
rect 35318 34159 35327 34277
rect 44800 34263 44918 34268
rect 35195 31130 35323 34159
rect 44796 34155 44805 34263
rect 44913 34155 44922 34263
rect 40652 32525 40661 32643
rect 40779 32525 40788 32643
rect 36513 31145 36631 31154
rect 35188 31121 35332 31130
rect 33480 30993 33486 31121
rect 33614 30993 33620 31121
rect 35188 30993 35195 31121
rect 35323 30993 35332 31121
rect 33486 26643 33614 30993
rect 35188 30986 35332 30993
rect 35196 27634 35202 27752
rect 35320 27634 35326 27752
rect 35202 26862 35320 27634
rect 35202 26817 35323 26862
rect 33485 26617 33614 26643
rect 33485 23148 33613 26617
rect 33479 23142 33619 23148
rect 33479 23014 33485 23142
rect 33613 23014 33619 23142
rect 33479 23008 33619 23014
rect 33485 21124 33613 23008
rect 33474 21115 33620 21124
rect 33474 20987 33485 21115
rect 33613 20987 33620 21115
rect 33474 20977 33620 20987
rect 35205 19128 35323 26817
rect 36513 24596 36631 31027
rect 40661 25442 40779 32525
rect 40661 25318 40779 25324
rect 42143 31066 42261 31075
rect 36507 24478 36513 24596
rect 36631 24478 36637 24596
rect 41228 23870 41356 23880
rect 41228 23732 41356 23742
rect 40368 23590 40432 23600
rect 41329 23590 41393 23594
rect 41701 23590 41765 23600
rect 40432 23584 41701 23590
rect 40432 23526 41329 23584
rect 40368 23516 40432 23526
rect 41393 23526 41701 23584
rect 41329 23510 41393 23520
rect 41701 23516 41765 23526
rect 39914 22775 39978 22785
rect 40371 22775 40435 22783
rect 41332 22775 41396 22782
rect 39978 22773 41396 22775
rect 39978 22711 40371 22773
rect 39914 22701 39978 22711
rect 40435 22772 41396 22773
rect 40435 22711 41332 22772
rect 40371 22699 40435 22709
rect 41332 22698 41396 22708
rect 40383 22578 40511 22588
rect 40383 22440 40511 22450
rect 36843 21883 36971 21893
rect 36843 21745 36971 21755
rect 36789 21586 36853 21596
rect 37758 21587 37822 21597
rect 36784 21522 36789 21586
rect 36853 21523 37758 21586
rect 37822 21523 38308 21586
rect 36853 21522 38308 21523
rect 38372 21522 38381 21586
rect 36789 21512 36853 21522
rect 37758 21513 37822 21522
rect 38486 20990 38492 21108
rect 38610 20990 38616 21108
rect 36278 20773 36342 20783
rect 36796 20773 36860 20781
rect 37755 20773 37819 20782
rect 36342 20772 37822 20773
rect 36342 20771 37755 20772
rect 36342 20709 36796 20771
rect 36278 20699 36342 20709
rect 36860 20709 37755 20771
rect 36796 20697 36860 20707
rect 37819 20709 37822 20772
rect 37755 20698 37819 20708
rect 37638 20579 37766 20589
rect 37638 20441 37766 20451
rect 38492 20166 38610 20990
rect 36843 19885 36971 19895
rect 36843 19747 36971 19757
rect 36796 19592 36860 19599
rect 37758 19593 37822 19603
rect 36792 19589 37758 19592
rect 36792 19528 36796 19589
rect 36860 19529 37758 19589
rect 38307 19592 38371 19602
rect 37822 19529 38307 19592
rect 36860 19528 38307 19529
rect 36796 19515 36860 19525
rect 37758 19519 37822 19528
rect 38307 19518 38371 19528
rect 35199 19010 35205 19128
rect 35323 19010 35329 19128
rect 38492 19118 38610 20048
rect 35205 17093 35323 19010
rect 38486 19000 38492 19118
rect 38610 19000 38616 19118
rect 42143 19116 42261 30948
rect 44800 27752 44918 34155
rect 78620 33654 78748 55438
rect 72414 33526 72420 33654
rect 72548 33526 72554 33654
rect 67532 33421 67681 33440
rect 67532 33303 67550 33421
rect 67668 33303 67681 33421
rect 67532 33291 67681 33303
rect 50229 32549 50238 32667
rect 50356 32549 50365 32667
rect 45534 27636 45652 27638
rect 44800 27628 44918 27634
rect 45524 27628 45652 27636
rect 45524 27510 45534 27628
rect 45524 27096 45652 27510
rect 50238 27224 50356 32549
rect 55952 31354 56299 31364
rect 55952 30744 56299 30754
rect 60986 30188 61191 30198
rect 60986 29638 61191 29648
rect 64046 29330 64252 29339
rect 64046 29115 64252 29124
rect 59363 28687 61033 28697
rect 59363 28450 61033 28460
rect 67550 27921 67668 27927
rect 50238 27096 50358 27224
rect 43018 24596 43136 24602
rect 43018 23112 43136 24478
rect 43018 21108 43136 22994
rect 43434 21662 43562 21672
rect 43434 21524 43562 21534
rect 43411 21403 43475 21413
rect 44371 21403 44435 21413
rect 43475 21339 44371 21403
rect 43411 21329 43475 21339
rect 44371 21329 44435 21339
rect 44809 20991 44815 21109
rect 44933 20991 44939 21109
rect 43018 20984 43136 20990
rect 43010 20582 43074 20592
rect 43413 20583 43477 20593
rect 43074 20519 43413 20582
rect 44376 20585 44440 20595
rect 43477 20521 44376 20582
rect 44440 20521 44445 20582
rect 43477 20519 44445 20521
rect 43074 20518 44445 20519
rect 43010 20508 43074 20518
rect 43413 20509 43477 20518
rect 44376 20511 44440 20518
rect 44260 20397 44388 20407
rect 44260 20259 44388 20269
rect 44815 20166 44933 20991
rect 45524 20171 45642 27096
rect 50240 26577 50358 27096
rect 50240 26453 50358 26459
rect 53293 27103 53411 27109
rect 51068 23839 51186 23849
rect 51068 23711 51186 23721
rect 51046 23580 51110 23590
rect 52012 23580 52076 23590
rect 52551 23580 52615 23590
rect 51110 23516 52012 23580
rect 52076 23516 52551 23580
rect 51046 23506 51110 23516
rect 52012 23506 52076 23516
rect 52551 23506 52615 23516
rect 46206 23116 46324 23122
rect 53293 23110 53411 26985
rect 58216 26577 58334 26583
rect 54495 25871 54501 25989
rect 54619 25871 54625 25989
rect 44809 20048 44815 20166
rect 44933 20048 44939 20166
rect 45518 20053 45524 20171
rect 45642 20053 45648 20171
rect 43415 19654 43543 19664
rect 43415 19516 43543 19526
rect 43407 19402 43471 19412
rect 44369 19409 44433 19412
rect 44367 19402 44433 19409
rect 43471 19399 44369 19402
rect 43471 19338 44367 19399
rect 44433 19338 44434 19402
rect 43407 19328 43471 19338
rect 44431 19335 44433 19338
rect 44367 19328 44433 19335
rect 44367 19325 44431 19328
rect 43009 19116 43127 19122
rect 42137 18998 42143 19116
rect 42261 18998 42267 19116
rect 44815 19109 44933 20048
rect 46206 19143 46324 22998
rect 53287 22992 53293 23110
rect 53411 22992 53417 23110
rect 50506 22768 50570 22778
rect 51047 22768 51111 22776
rect 52009 22768 52073 22773
rect 50570 22766 52074 22768
rect 50570 22704 51047 22766
rect 50506 22694 50570 22704
rect 51111 22763 52074 22766
rect 51111 22704 52009 22763
rect 51047 22692 51111 22702
rect 52073 22704 52074 22763
rect 52009 22689 52073 22699
rect 51940 22587 52058 22597
rect 51940 22459 52058 22469
rect 47795 21847 47923 21857
rect 47795 21709 47923 21719
rect 48704 21593 48768 21594
rect 47739 21584 47803 21592
rect 48702 21584 48768 21593
rect 47739 21583 48704 21584
rect 47739 21582 48702 21583
rect 47803 21520 48702 21582
rect 47739 21508 47803 21518
rect 48766 21519 48768 21520
rect 48702 21510 48768 21519
rect 48702 21509 48766 21510
rect 47050 21127 47168 21133
rect 53293 21113 53411 22992
rect 36280 18771 36344 18781
rect 36796 18772 36860 18782
rect 36344 18708 36796 18771
rect 37756 18771 37820 18781
rect 36860 18708 37756 18771
rect 36344 18707 37756 18708
rect 36280 18697 36344 18707
rect 36796 18698 36860 18707
rect 37756 18697 37820 18707
rect 37633 18578 37761 18588
rect 37633 18440 37761 18450
rect 40397 17866 40525 17876
rect 40397 17728 40525 17738
rect 40367 17587 40431 17597
rect 41333 17587 41397 17596
rect 41702 17587 41766 17597
rect 40363 17523 40367 17587
rect 40431 17586 41702 17587
rect 40431 17523 41333 17586
rect 40367 17513 40431 17523
rect 41397 17523 41702 17586
rect 41766 17523 41781 17587
rect 41333 17512 41397 17522
rect 41702 17513 41766 17523
rect 43009 17127 43127 18998
rect 44809 18991 44815 19109
rect 44933 18991 44939 19109
rect 46200 19025 46206 19143
rect 46324 19025 46330 19143
rect 43411 18582 43475 18592
rect 44372 18582 44436 18591
rect 43409 18518 43411 18582
rect 43475 18581 44436 18582
rect 43475 18518 44372 18581
rect 43411 18508 43475 18518
rect 44372 18507 44436 18517
rect 44259 18389 44387 18399
rect 44259 18251 44387 18261
rect 35199 16975 35205 17093
rect 35323 16975 35329 17093
rect 43009 17003 43127 17009
rect 47050 17115 47168 21009
rect 53287 20995 53293 21113
rect 53411 20995 53417 21113
rect 47737 20767 47801 20777
rect 48698 20768 48762 20778
rect 47801 20704 48698 20765
rect 48762 20704 48764 20765
rect 47801 20703 48764 20704
rect 47737 20701 48764 20703
rect 47737 20693 47801 20701
rect 48698 20694 48762 20701
rect 48603 20577 48731 20587
rect 48603 20439 48731 20449
rect 47791 19842 47919 19852
rect 47791 19704 47919 19714
rect 47739 19583 47803 19593
rect 48695 19583 48759 19593
rect 47803 19519 48695 19582
rect 49357 19582 49421 19592
rect 48759 19519 49357 19582
rect 47739 19518 49357 19519
rect 47739 19509 47803 19518
rect 48695 19509 48759 19518
rect 49357 19508 49421 19518
rect 53300 18994 53306 19112
rect 53424 18994 53430 19112
rect 47735 18761 47801 18771
rect 48697 18761 48761 18770
rect 47801 18760 48761 18761
rect 47801 18697 48697 18760
rect 47735 18687 47801 18697
rect 48697 18686 48761 18696
rect 48603 18578 48731 18588
rect 48603 18440 48731 18450
rect 53306 18089 53424 18994
rect 54501 18089 54619 25871
rect 55642 25442 55760 25448
rect 55642 18168 55760 25324
rect 56908 25217 56914 25335
rect 57032 25217 57038 25335
rect 56914 19113 57032 25217
rect 58216 22221 58334 26459
rect 67550 25335 67668 27803
rect 68703 27908 68821 27914
rect 67544 25217 67550 25335
rect 67668 25217 67674 25335
rect 59555 24414 59673 24420
rect 68703 24414 68821 27790
rect 72420 27190 72548 33526
rect 78620 33520 78748 33526
rect 79370 54966 79498 54972
rect 79370 32906 79498 54838
rect 80625 41373 80753 56167
rect 80625 41239 80753 41245
rect 81000 41431 81064 41440
rect 80174 41159 80238 41163
rect 80174 41153 80239 41159
rect 80238 41089 80239 41153
rect 80174 41079 80239 41089
rect 79904 40739 79983 40749
rect 79904 40451 79983 40461
rect 80175 40182 80239 41079
rect 81000 41150 81064 41367
rect 82647 41389 82775 57103
rect 85384 54968 85512 58068
rect 86728 58170 86856 58176
rect 86728 55572 86856 58042
rect 94495 55627 94623 66623
rect 103835 64910 103963 66742
rect 103835 64862 103967 64910
rect 101829 64129 101947 64134
rect 101825 64021 101834 64129
rect 101942 64021 101951 64129
rect 103839 64108 103967 64862
rect 101829 60403 101947 64021
rect 103839 63974 103967 63980
rect 102782 63849 102972 63859
rect 104139 63858 104283 63868
rect 102782 63747 102972 63757
rect 103222 63823 103656 63833
rect 104139 63754 104283 63764
rect 104558 63809 104982 63819
rect 103222 63726 103656 63736
rect 104558 63722 104982 63732
rect 105687 62929 105805 62934
rect 105683 62821 105692 62929
rect 105800 62821 105809 62929
rect 102873 62346 102965 62356
rect 102873 62227 102965 62237
rect 104204 62341 104296 62351
rect 104204 62222 104296 62232
rect 103748 60499 103813 60509
rect 101829 60285 102645 60403
rect 105687 60412 105805 62821
rect 103748 60347 103813 60357
rect 104981 60294 105805 60412
rect 103198 60274 103269 60284
rect 103198 60160 103269 60170
rect 104290 60280 104358 60290
rect 104290 60160 104358 60170
rect 102597 59636 102710 59646
rect 102597 59513 102710 59523
rect 104990 59030 105103 59040
rect 104990 58907 105103 58917
rect 103038 58196 103166 58202
rect 86728 55566 86858 55572
rect 86728 55438 86730 55566
rect 92020 55499 92026 55627
rect 92154 55499 92160 55627
rect 94489 55499 94495 55627
rect 94623 55499 94629 55627
rect 103038 55499 103166 58068
rect 104382 58170 104510 58176
rect 104382 56792 104510 58042
rect 104380 56674 104386 56792
rect 104504 56674 104510 56792
rect 114075 56674 114081 56792
rect 114199 56674 114205 56792
rect 112927 55509 113045 55515
rect 86728 55432 86858 55438
rect 86728 55406 86856 55432
rect 85384 54834 85512 54840
rect 87250 53960 87368 53966
rect 85339 53292 85345 53410
rect 85463 53292 85469 53410
rect 85345 43190 85463 53292
rect 85593 43237 85657 43246
rect 85339 43072 85345 43190
rect 85463 43072 85469 43190
rect 87250 43186 87368 53842
rect 92026 50855 92154 55499
rect 103035 55381 103041 55499
rect 103159 55405 103166 55499
rect 112911 55499 113054 55509
rect 103159 55381 103165 55405
rect 112911 55381 112927 55499
rect 113045 55381 113054 55499
rect 112911 55370 113054 55381
rect 91962 50845 92205 50855
rect 91962 50588 92205 50598
rect 102494 50225 102722 50235
rect 100698 50213 100886 50223
rect 100698 50009 100886 50019
rect 106007 50217 106235 50227
rect 102494 49983 102722 49993
rect 104188 50206 104416 50216
rect 106007 49975 106235 49985
rect 107791 50214 108019 50224
rect 104188 49964 104416 49974
rect 107791 49972 108019 49982
rect 109576 50212 109804 50222
rect 109576 49970 109804 49980
rect 96364 49834 97874 49844
rect 96364 49422 97874 49432
rect 101678 48668 101914 48678
rect 99808 48638 100084 48648
rect 101678 48580 101914 48590
rect 103483 48661 103717 48671
rect 103483 48572 103717 48582
rect 105289 48657 105508 48667
rect 105289 48566 105508 48576
rect 107075 48661 107315 48671
rect 108876 48657 109128 48667
rect 108876 48582 109128 48592
rect 107075 48567 107315 48577
rect 99808 48528 100084 48538
rect 90796 47320 91108 47330
rect 94987 47300 96094 47310
rect 94987 47073 96094 47083
rect 90796 46772 91108 46782
rect 87594 43237 87658 43246
rect 85593 42961 85657 43173
rect 87244 43068 87250 43186
rect 87368 43068 87374 43186
rect 87594 42965 87658 43173
rect 84767 42950 84831 42961
rect 84505 42609 84628 42619
rect 84505 42257 84628 42267
rect 84767 41999 84831 42886
rect 85592 42951 85657 42961
rect 86767 42959 86831 42960
rect 85656 42887 85657 42951
rect 85592 42877 85657 42887
rect 85593 42002 85657 42877
rect 86765 42950 86831 42959
rect 86765 42886 86767 42950
rect 86765 42876 86831 42886
rect 87593 42955 87658 42965
rect 87657 42891 87658 42955
rect 87593 42881 87658 42891
rect 86529 42646 86618 42656
rect 86529 42252 86618 42262
rect 84766 41989 84831 41999
rect 84830 41925 84831 41989
rect 85592 41992 85657 42002
rect 84766 41915 84831 41925
rect 84767 41728 84831 41915
rect 84767 41653 84831 41664
rect 85240 41968 85368 41974
rect 85656 41928 85657 41992
rect 86765 41999 86829 42876
rect 86765 41989 86830 41999
rect 85592 41918 85656 41928
rect 86765 41925 86766 41989
rect 87594 41990 87658 42881
rect 82647 41255 82775 41261
rect 83000 41440 83064 41449
rect 81000 40188 81064 41086
rect 82166 41152 82240 41168
rect 81965 40703 82045 40713
rect 81965 40410 82045 40420
rect 80175 39921 80239 40118
rect 80633 40168 80780 40176
rect 80633 40040 80643 40168
rect 80771 40040 80780 40168
rect 81000 40114 81064 40124
rect 82166 40191 82240 41078
rect 83000 41148 83064 41376
rect 83000 40200 83064 41084
rect 82998 40190 83072 40200
rect 80633 40033 80780 40040
rect 80175 39848 80239 39857
rect 80643 38567 80771 40033
rect 82166 39931 82240 40117
rect 82639 40034 82645 40162
rect 82773 40034 82779 40162
rect 82998 40106 83072 40116
rect 82156 39923 82245 39931
rect 82156 39849 82166 39923
rect 82240 39849 82245 39923
rect 82156 39836 82245 39849
rect 81151 39699 81299 39719
rect 81151 39581 81167 39699
rect 81285 39581 81299 39699
rect 81151 39557 81299 39581
rect 82645 39407 82773 40034
rect 83018 39719 83142 39729
rect 83018 39585 83142 39595
rect 82645 39273 82773 39279
rect 85240 38567 85368 41840
rect 86765 41915 86830 41925
rect 87247 41957 87375 41963
rect 86765 41731 86829 41915
rect 86765 41658 86829 41667
rect 87594 41916 87658 41926
rect 96525 42681 96795 42691
rect 85864 41236 86138 41252
rect 85864 41010 85888 41236
rect 86114 41010 86138 41236
rect 85864 40988 86138 41010
rect 86317 39417 86445 39423
rect 87247 39407 87375 41829
rect 96525 41596 96795 41606
rect 97372 42678 97642 42688
rect 97972 42396 98218 42406
rect 97972 41672 98218 41682
rect 97372 41593 97642 41603
rect 87796 41218 88032 41236
rect 87796 41017 87813 41218
rect 88014 41017 88032 41218
rect 87796 41000 88032 41017
rect 82304 38439 82310 38567
rect 82438 38439 82444 38567
rect 85234 38439 85240 38567
rect 85368 38439 85374 38567
rect 80643 38433 80771 38439
rect 82310 33160 82438 38439
rect 86317 37663 86445 39289
rect 87241 39279 87247 39407
rect 87375 39279 87381 39407
rect 90783 38958 91030 38968
rect 90783 38081 91030 38091
rect 85315 37535 85321 37663
rect 85449 37535 85455 37663
rect 83771 34890 83928 34908
rect 83771 34762 83785 34890
rect 83913 34762 83928 34890
rect 83771 34736 83928 34762
rect 83635 33792 83781 33808
rect 83635 33674 83651 33792
rect 83769 33674 83781 33792
rect 83635 33661 83781 33674
rect 82676 33515 82740 33519
rect 82671 33459 82680 33515
rect 82736 33459 82745 33515
rect 85007 33512 85071 33516
rect 82310 33023 82438 33032
rect 73786 32778 73792 32906
rect 73920 32778 73926 32906
rect 69632 27062 69638 27190
rect 69766 27062 69772 27190
rect 68697 24296 68703 24414
rect 68821 24296 68827 24414
rect 59555 23133 59673 24296
rect 62988 23840 63106 23850
rect 62988 23712 63106 23722
rect 62977 23583 63041 23593
rect 63940 23583 64004 23593
rect 62973 23519 62977 23583
rect 63041 23519 63940 23583
rect 64004 23519 64445 23583
rect 64509 23519 64518 23583
rect 62977 23509 63041 23519
rect 63940 23509 64004 23519
rect 58210 22103 58216 22221
rect 58334 22103 58340 22221
rect 59555 21114 59673 23015
rect 65692 23105 65810 23111
rect 62978 22761 63042 22771
rect 62411 22696 62420 22760
rect 62484 22697 62978 22760
rect 63937 22761 64001 22771
rect 63042 22697 63937 22760
rect 64001 22697 64004 22760
rect 62484 22696 64004 22697
rect 62978 22687 63042 22696
rect 63937 22687 64001 22696
rect 63860 22582 63978 22592
rect 63860 22454 63978 22464
rect 63197 22103 63203 22221
rect 63321 22103 63327 22221
rect 60239 21871 60357 21881
rect 60239 21743 60357 21753
rect 60257 21584 60321 21594
rect 61219 21584 61283 21593
rect 60321 21583 61664 21584
rect 60321 21520 61219 21583
rect 60257 21510 60321 21520
rect 61283 21520 61664 21583
rect 61728 21520 61737 21584
rect 61219 21509 61283 21519
rect 63203 21111 63321 22103
rect 59555 20990 59673 20996
rect 63197 20993 63203 21111
rect 63321 20993 63327 21111
rect 64416 20993 64422 21111
rect 64540 20993 64546 21111
rect 60255 20763 60319 20771
rect 61219 20763 61283 20773
rect 59689 20699 59698 20763
rect 59762 20761 61219 20763
rect 59762 20699 60255 20761
rect 60319 20699 61219 20761
rect 60255 20687 60319 20697
rect 61219 20689 61283 20699
rect 61061 20579 61179 20589
rect 61061 20451 61179 20461
rect 60241 19841 60359 19851
rect 60241 19713 60359 19723
rect 60254 19582 60318 19592
rect 60251 19518 60254 19581
rect 61219 19583 61283 19593
rect 60318 19519 61219 19581
rect 61283 19519 61667 19581
rect 60318 19518 61667 19519
rect 60251 19517 61667 19518
rect 61731 19517 61740 19581
rect 60254 19508 60318 19517
rect 61219 19509 61283 19517
rect 54495 17971 54501 18089
rect 54619 17971 54625 18089
rect 55636 18050 55642 18168
rect 55760 18050 55766 18168
rect 51104 17840 51222 17850
rect 51104 17712 51222 17722
rect 51044 17582 51108 17592
rect 51038 17518 51044 17580
rect 52011 17583 52075 17593
rect 51108 17519 52011 17580
rect 52547 17580 52611 17590
rect 52075 17519 52547 17580
rect 51108 17518 52547 17519
rect 51038 17516 52547 17518
rect 51044 17508 51108 17516
rect 52011 17509 52075 17516
rect 52547 17506 52611 17516
rect 53306 17109 53424 17971
rect 56914 17157 57032 18995
rect 63202 19112 63337 19122
rect 63202 18994 63210 19112
rect 63328 18994 63337 19112
rect 63202 18987 63337 18994
rect 59710 18764 59774 18774
rect 60257 18764 60321 18773
rect 61221 18765 61285 18775
rect 59774 18763 61221 18764
rect 59774 18700 60257 18763
rect 59710 18690 59774 18700
rect 60321 18701 61221 18763
rect 60321 18700 61285 18701
rect 60257 18689 60321 18699
rect 61221 18691 61285 18700
rect 61055 18583 61173 18593
rect 61055 18455 61173 18465
rect 63210 18168 63328 18987
rect 63210 18044 63328 18050
rect 63015 17833 63133 17843
rect 63015 17705 63133 17715
rect 62980 17583 63044 17591
rect 63942 17583 64006 17592
rect 62980 17582 64018 17583
rect 62980 17581 63942 17582
rect 63044 17519 63942 17581
rect 62980 17507 63044 17517
rect 64006 17519 64018 17582
rect 63942 17508 64006 17518
rect 47050 16991 47168 16997
rect 53300 16991 53306 17109
rect 53424 16991 53430 17109
rect 56908 17039 56914 17157
rect 57032 17039 57038 17157
rect 64422 17112 64540 20993
rect 65692 19112 65810 22987
rect 67640 23110 67758 23120
rect 67640 20871 67758 22992
rect 67161 20795 67225 20805
rect 67640 20743 67758 20753
rect 67989 20792 68053 20802
rect 67161 20721 67225 20731
rect 67989 20718 68053 20728
rect 66649 20332 66767 20342
rect 66649 20204 66767 20214
rect 68386 20324 68504 20334
rect 68386 20196 68504 20206
rect 67163 19825 67227 19835
rect 67163 19751 67227 19761
rect 67985 19826 68049 19836
rect 67985 19752 68049 19762
rect 65692 18988 65810 18994
rect 67637 19645 67755 19655
rect 64422 16988 64540 16994
rect 67637 17123 67755 19527
rect 67637 17113 67756 17123
rect 67637 16995 67638 17113
rect 67637 16990 67756 16995
rect 67638 16985 67756 16990
rect 69638 17086 69766 27062
rect 72420 27056 72548 27062
rect 73792 24748 73920 32778
rect 79370 32772 79498 32778
rect 82676 32063 82740 33459
rect 85002 33456 85011 33512
rect 85067 33456 85076 33512
rect 82676 31990 82740 31999
rect 81950 31877 82093 31890
rect 77064 31759 77070 31877
rect 77188 31759 77194 31877
rect 81950 31759 81964 31877
rect 82082 31759 82093 31877
rect 85007 31814 85071 33456
rect 85321 33167 85449 37535
rect 86317 37529 86445 37535
rect 103349 37299 103593 37309
rect 101446 37239 101690 37249
rect 99844 37228 100088 37238
rect 103349 37089 103593 37099
rect 105066 37283 105310 37293
rect 105066 37073 105310 37083
rect 106880 37278 107124 37288
rect 106880 37068 107124 37078
rect 108852 37272 109096 37282
rect 108852 37062 109096 37072
rect 101446 37029 101690 37039
rect 99844 37018 100088 37028
rect 86367 35894 86373 36022
rect 86501 35894 86507 36022
rect 86373 35338 86501 35894
rect 89481 35852 89487 36058
rect 89693 35852 89699 36058
rect 89487 35532 89693 35852
rect 96849 35851 97596 35861
rect 96849 35730 97596 35740
rect 100366 35727 100750 35737
rect 102157 35734 102557 35744
rect 102157 35650 102557 35660
rect 103963 35734 104351 35744
rect 103963 35650 104351 35660
rect 105760 35699 106148 35709
rect 100366 35639 100750 35649
rect 105760 35615 106148 35625
rect 107562 35699 107949 35709
rect 107562 35611 107949 35621
rect 109356 35695 109751 35705
rect 109356 35608 109751 35618
rect 86360 35325 86514 35338
rect 89483 35336 89492 35532
rect 89688 35336 89697 35532
rect 89487 35331 89693 35336
rect 86360 35197 86373 35325
rect 86501 35197 86514 35325
rect 86360 35183 86514 35197
rect 107906 35018 108113 35024
rect 108234 35017 108441 35023
rect 110866 35017 110984 35020
rect 88556 34918 88762 34924
rect 88556 34379 88762 34712
rect 107906 34810 108106 34811
rect 108441 34810 110831 35017
rect 111038 34810 111044 35017
rect 95270 34384 95466 34388
rect 95265 34379 95893 34384
rect 88552 34183 88561 34379
rect 88757 34183 88766 34379
rect 95265 34183 95270 34379
rect 95466 34183 95893 34379
rect 88556 34178 88762 34183
rect 95265 34178 95893 34183
rect 95270 34174 95466 34178
rect 85321 33030 85449 33039
rect 88643 33792 88761 33798
rect 85787 31831 85919 31850
rect 70420 24620 70426 24748
rect 70554 24620 70560 24748
rect 70426 23126 70554 24620
rect 73792 24614 73920 24620
rect 71557 23837 71675 23847
rect 71557 23709 71675 23719
rect 71541 23587 71605 23594
rect 72507 23587 72571 23597
rect 71541 23584 72507 23587
rect 71605 23523 72507 23584
rect 72571 23523 72875 23587
rect 72939 23523 72948 23587
rect 71541 23510 71605 23520
rect 72507 23513 72571 23523
rect 77070 23123 77188 31759
rect 81950 31747 82093 31759
rect 84866 31696 84971 31814
rect 85089 31696 85098 31814
rect 85787 31723 85799 31831
rect 85907 31723 85919 31831
rect 85787 31709 85919 31723
rect 86655 31819 86797 31833
rect 82222 31330 82358 31343
rect 82222 31222 82236 31330
rect 82344 31222 82358 31330
rect 82222 31211 82358 31222
rect 77947 29252 77953 29370
rect 78071 29252 78077 29370
rect 70426 22992 70554 22998
rect 74332 23108 74450 23118
rect 77070 22999 77188 23005
rect 71543 22762 71607 22772
rect 71177 22697 71186 22761
rect 71250 22698 71543 22761
rect 72509 22765 72573 22775
rect 71607 22701 72509 22761
rect 71607 22698 72573 22701
rect 71250 22697 72573 22698
rect 71543 22688 71607 22697
rect 72509 22691 72573 22697
rect 72435 22578 72553 22588
rect 72435 22450 72553 22460
rect 74332 20625 74450 22990
rect 74028 20545 74092 20555
rect 74332 20497 74450 20507
rect 74856 20551 74920 20561
rect 74028 20471 74092 20481
rect 74856 20477 74920 20487
rect 75276 20093 75394 20103
rect 73565 20070 73683 20080
rect 75276 19965 75394 19975
rect 73565 19942 73683 19952
rect 74034 19583 74098 19593
rect 74034 19509 74098 19519
rect 74860 19582 74924 19592
rect 74860 19508 74924 19518
rect 74324 19293 74330 19411
rect 74448 19293 74454 19411
rect 71584 17844 71702 17854
rect 71584 17716 71702 17726
rect 71543 17594 71607 17603
rect 72501 17594 72565 17604
rect 71541 17593 72501 17594
rect 71541 17530 71543 17593
rect 71607 17530 72501 17593
rect 72565 17530 72882 17594
rect 72946 17530 72955 17594
rect 71543 17519 71607 17529
rect 72501 17520 72565 17530
rect 74330 17123 74448 19293
rect 74330 16999 74448 17005
rect 77953 17121 78071 29252
rect 82231 28361 82349 31211
rect 84866 29370 84984 31696
rect 84860 29252 84866 29370
rect 84984 29252 84990 29370
rect 79190 28351 79308 28357
rect 79190 23117 79308 28233
rect 82222 28351 82355 28361
rect 82222 28233 82231 28351
rect 82349 28233 82355 28351
rect 82222 28226 82355 28233
rect 82231 28220 82349 28226
rect 80129 27142 80247 27148
rect 79184 22999 79190 23117
rect 79308 22999 79314 23117
rect 77953 16997 78071 17003
rect 80129 17124 80247 27024
rect 85794 27142 85912 31709
rect 86655 31701 86666 31819
rect 86784 31701 86797 31819
rect 86655 31685 86797 31701
rect 87767 31819 87885 31825
rect 85794 27018 85912 27024
rect 86377 24988 86495 24998
rect 86377 24860 86495 24870
rect 85581 24727 85645 24737
rect 86544 24728 86608 24738
rect 85203 24663 85212 24727
rect 85276 24663 85581 24727
rect 85645 24664 86544 24727
rect 86608 24664 86612 24727
rect 85645 24663 86612 24664
rect 85581 24653 85645 24663
rect 86544 24654 86608 24663
rect 81503 24304 81509 24422
rect 81627 24304 81633 24422
rect 81509 23108 81627 24304
rect 85581 23902 85645 23912
rect 86543 23902 86607 23911
rect 85645 23901 87019 23902
rect 85645 23838 86543 23901
rect 85581 23828 85645 23838
rect 86607 23838 87019 23901
rect 87083 23838 87092 23902
rect 86543 23827 86607 23837
rect 83055 23772 83173 23782
rect 83055 23644 83173 23654
rect 85591 23722 85709 23732
rect 85591 23594 85709 23604
rect 82221 23539 82285 23549
rect 81868 23474 81877 23538
rect 81941 23475 82221 23538
rect 83183 23538 83247 23546
rect 82285 23536 83247 23538
rect 82285 23475 83183 23536
rect 81941 23474 83183 23475
rect 82221 23465 82285 23474
rect 83183 23462 83247 23472
rect 83768 23241 83886 23247
rect 81503 22990 81509 23108
rect 81627 22990 81633 23108
rect 82220 22711 82284 22721
rect 83181 22711 83245 22720
rect 82217 22647 82220 22711
rect 82284 22710 83459 22711
rect 82284 22647 83181 22710
rect 82220 22637 82284 22647
rect 83245 22647 83459 22710
rect 83523 22647 83532 22711
rect 83181 22636 83245 22646
rect 82256 22522 82374 22532
rect 82256 22394 82374 22404
rect 83768 20218 83886 23123
rect 83758 20208 83896 20218
rect 83758 20090 83768 20208
rect 83886 20090 83896 20208
rect 83758 20084 83896 20090
rect 82968 17813 83086 17823
rect 82968 17685 83086 17695
rect 82223 17567 82287 17577
rect 83186 17567 83250 17577
rect 81873 17503 81882 17567
rect 81946 17503 82223 17567
rect 82287 17503 83186 17567
rect 82223 17493 82287 17503
rect 83186 17493 83250 17503
rect 83768 17279 83886 20084
rect 87767 18837 87885 31701
rect 88643 26607 88761 33674
rect 107906 32601 108113 34810
rect 108234 34804 108441 34810
rect 112927 34412 113045 55370
rect 114081 39736 114199 56674
rect 116738 52514 116866 52524
rect 116738 52376 116866 52386
rect 120662 52467 120933 52477
rect 120662 52353 120933 52363
rect 119326 52130 119407 52140
rect 117729 51778 117832 51788
rect 115289 51725 115385 51735
rect 117729 51306 117832 51316
rect 115289 51263 115385 51273
rect 121709 52123 121804 52133
rect 121709 51017 121804 51027
rect 119326 50991 119407 51001
rect 117396 50953 117553 50963
rect 121196 50958 121516 50968
rect 115579 50928 115707 50938
rect 115579 50790 115707 50800
rect 115989 50861 116141 50871
rect 116367 50862 116419 50910
rect 115989 50699 116141 50709
rect 116334 49381 116452 50862
rect 116911 50850 116963 50914
rect 117396 50859 117553 50869
rect 119936 50944 120225 50954
rect 116873 50236 116991 50850
rect 121196 50878 121516 50888
rect 119936 50762 120225 50772
rect 116867 50118 116873 50236
rect 116991 50118 116997 50236
rect 120335 49387 120453 50858
rect 120884 50236 121002 50864
rect 126619 50236 126751 50243
rect 120878 50118 120884 50236
rect 121002 50118 121008 50236
rect 126619 50118 126626 50236
rect 126744 50118 126751 50236
rect 126619 50111 126751 50118
rect 120328 49381 120460 49387
rect 116328 49263 116334 49381
rect 116452 49263 116458 49381
rect 120328 49263 120335 49381
rect 120453 49263 120460 49381
rect 125951 49263 125957 49381
rect 126075 49263 126081 49381
rect 120328 49256 120460 49263
rect 117034 39618 117040 39736
rect 117158 39618 117164 39736
rect 114081 35221 114199 39618
rect 117040 39470 117167 39618
rect 114709 39378 115008 39388
rect 114709 38727 115008 38737
rect 117049 38289 117167 39470
rect 123011 38345 123095 38355
rect 123011 37042 123095 37052
rect 123011 36885 123095 36895
rect 123011 35582 123095 35592
rect 114079 35023 114199 35221
rect 123012 35405 123095 35415
rect 114007 35017 114214 35023
rect 114007 34804 114214 34810
rect 112881 34406 113088 34412
rect 125957 34488 126075 49263
rect 123012 34377 123095 34387
rect 125951 34370 125957 34488
rect 126075 34370 126081 34488
rect 112881 34193 113088 34199
rect 107900 32394 107906 32601
rect 108113 32394 108119 32601
rect 95427 31246 95711 31256
rect 95427 30779 95711 30789
rect 90814 30752 91056 30762
rect 90814 30278 91056 30288
rect 95203 28684 95762 28694
rect 95203 28454 95762 28464
rect 112927 28430 113045 34193
rect 125028 34131 125348 34141
rect 125028 33801 125348 33811
rect 126626 33700 126744 50111
rect 128011 34932 129048 34952
rect 128011 33932 128026 34932
rect 129026 33932 129048 34932
rect 128011 33908 129048 33932
rect 127217 33739 127594 33749
rect 123010 33617 123097 33627
rect 126620 33582 126626 33700
rect 126744 33582 126750 33700
rect 127217 33656 127594 33666
rect 123010 32633 123097 32643
rect 127219 32617 127591 32627
rect 127219 32542 127591 32552
rect 123007 32470 123097 32480
rect 114716 31367 115015 31377
rect 123007 31094 123097 31104
rect 124329 31186 124649 31196
rect 114716 30716 115015 30726
rect 123008 30864 123099 30874
rect 112921 28312 112927 28430
rect 113045 28312 113051 28430
rect 117180 28422 117298 29684
rect 124329 30856 124649 30866
rect 123008 29596 123099 29606
rect 117180 28298 117298 28304
rect 107956 27185 108074 27191
rect 104393 27172 104511 27181
rect 104387 27054 104393 27172
rect 104511 27054 104517 27172
rect 107947 27067 107956 27185
rect 108074 27067 108083 27185
rect 107956 27061 108074 27067
rect 104393 27045 104511 27054
rect 93830 27016 94036 27033
rect 93830 26820 93840 27016
rect 94036 26820 94045 27016
rect 88637 26489 88643 26607
rect 88761 26489 88767 26607
rect 88643 24435 88761 26489
rect 88637 24317 88643 24435
rect 88761 24317 88767 24435
rect 88643 23243 88761 24317
rect 92590 23788 92708 23798
rect 92590 23660 92708 23670
rect 91820 23538 91884 23548
rect 91818 23474 91820 23537
rect 92780 23537 92844 23546
rect 91884 23536 93136 23537
rect 91884 23474 92780 23536
rect 91818 23473 92780 23474
rect 91820 23464 91884 23473
rect 92844 23473 93136 23536
rect 93200 23473 93209 23537
rect 92780 23462 92844 23472
rect 88637 23125 88643 23243
rect 88761 23125 88767 23243
rect 93273 23123 93279 23241
rect 93397 23123 93403 23241
rect 91819 22712 91883 22722
rect 92781 22714 92845 22724
rect 91383 22648 91392 22712
rect 91456 22648 91819 22712
rect 91883 22650 92781 22712
rect 91883 22648 92845 22650
rect 91819 22638 91883 22648
rect 92781 22640 92845 22648
rect 91882 22528 92000 22538
rect 91882 22400 92000 22410
rect 93279 20208 93397 23123
rect 93830 20242 94036 26820
rect 95000 25170 95118 25176
rect 93273 20090 93279 20208
rect 93397 20090 93403 20208
rect 87767 18713 87885 18719
rect 88626 18837 88744 18843
rect 83768 17155 83886 17161
rect 88626 17273 88744 18719
rect 92566 17819 92684 17829
rect 92566 17691 92684 17701
rect 91828 17567 91892 17577
rect 92780 17567 92844 17575
rect 91824 17503 91828 17567
rect 91892 17565 92782 17567
rect 91892 17503 92780 17565
rect 92846 17503 92855 17567
rect 91828 17493 91892 17503
rect 92780 17491 92844 17501
rect 93279 17274 93397 20090
rect 93824 20036 93830 20242
rect 94036 20036 94042 20242
rect 95000 18837 95118 25052
rect 106372 23428 106500 23438
rect 106372 23290 106500 23300
rect 105744 23166 105808 23176
rect 105413 23096 105422 23160
rect 105486 23102 105744 23160
rect 106706 23162 106770 23172
rect 105808 23102 106706 23160
rect 105486 23098 106706 23102
rect 105486 23096 106770 23098
rect 105744 23092 105808 23096
rect 106706 23088 106770 23096
rect 107984 22694 108092 22698
rect 104384 22675 104518 22682
rect 104384 22557 104393 22675
rect 104511 22557 104518 22675
rect 107973 22576 107979 22694
rect 108097 22576 108103 22694
rect 107984 22572 108092 22576
rect 104384 22544 104518 22557
rect 105741 22348 107095 22350
rect 105740 22339 107095 22348
rect 105740 22338 106706 22339
rect 105804 22276 106706 22338
rect 105740 22264 105804 22274
rect 106770 22276 107095 22339
rect 107169 22276 107178 22350
rect 106706 22265 106770 22275
rect 105796 22156 105924 22166
rect 105796 22018 105924 22028
rect 94994 18719 95000 18837
rect 95118 18719 95124 18837
rect 93273 17156 93279 17274
rect 93397 17156 93403 17274
rect 80129 17000 80247 17006
rect 81500 17123 81640 17137
rect 81500 17005 81510 17123
rect 81628 17005 81640 17123
rect 81500 16993 81640 17005
rect 69638 16952 69766 16958
rect 39911 16765 39975 16775
rect 40370 16765 40434 16775
rect 71544 16774 71608 16784
rect 72505 16775 72569 16785
rect 39975 16701 40370 16764
rect 41328 16764 41392 16772
rect 40434 16762 41396 16764
rect 40434 16701 41328 16762
rect 39911 16700 41328 16701
rect 39911 16691 39975 16700
rect 40370 16691 40434 16700
rect 41392 16700 41396 16762
rect 50503 16762 50567 16772
rect 51048 16762 51112 16770
rect 52008 16762 52072 16770
rect 62978 16763 63042 16772
rect 63938 16763 64002 16773
rect 41328 16688 41392 16698
rect 50567 16760 52072 16762
rect 50567 16698 51048 16760
rect 50503 16688 50567 16698
rect 51112 16698 52008 16760
rect 51048 16686 51112 16696
rect 62412 16699 62421 16763
rect 62485 16762 63938 16763
rect 62485 16699 62978 16762
rect 52008 16686 52072 16696
rect 63042 16699 63938 16762
rect 71181 16710 71190 16774
rect 71254 16710 71544 16774
rect 71608 16711 72505 16774
rect 71608 16710 72569 16711
rect 71544 16700 71608 16710
rect 72505 16701 72569 16710
rect 62978 16688 63042 16698
rect 63938 16689 64002 16699
rect 51817 16582 51935 16592
rect 41211 16542 41339 16552
rect 51817 16454 51935 16464
rect 63827 16573 63945 16583
rect 63827 16445 63945 16455
rect 72296 16582 72414 16592
rect 72296 16454 72414 16464
rect 41211 16404 41339 16414
rect 81510 16379 81628 16993
rect 86412 16962 86530 16972
rect 86412 16834 86530 16844
rect 82220 16747 82284 16752
rect 83186 16747 83250 16752
rect 82213 16742 83455 16747
rect 82213 16683 82220 16742
rect 82284 16683 83186 16742
rect 82220 16668 82284 16678
rect 83250 16683 83455 16742
rect 83519 16683 83528 16747
rect 85579 16717 85643 16727
rect 86542 16719 86606 16729
rect 83186 16668 83250 16678
rect 85201 16653 85210 16717
rect 85274 16653 85579 16717
rect 85643 16655 86542 16717
rect 86606 16655 86609 16717
rect 85643 16653 86609 16655
rect 85579 16643 85643 16653
rect 86542 16645 86606 16653
rect 82296 16561 82414 16571
rect 82296 16433 82414 16443
rect 88626 16423 88744 17155
rect 91823 16743 91887 16752
rect 92781 16745 92845 16755
rect 91393 16679 91402 16743
rect 91466 16742 92781 16743
rect 91466 16679 91823 16742
rect 91887 16681 92781 16742
rect 92845 16681 92847 16743
rect 91887 16679 92847 16681
rect 91823 16668 91887 16678
rect 92781 16671 92845 16679
rect 91859 16547 91977 16557
rect 81504 16261 81510 16379
rect 81628 16261 81634 16379
rect 88620 16305 88626 16423
rect 88744 16305 88750 16423
rect 91859 16419 91977 16429
rect 85579 15893 85643 15903
rect 85578 15829 85579 15892
rect 86541 15892 86605 15901
rect 85643 15891 87016 15892
rect 85643 15829 86541 15891
rect 85578 15828 86541 15829
rect 85579 15819 85643 15828
rect 86605 15828 87016 15891
rect 87080 15828 87089 15892
rect 86541 15817 86605 15827
rect 85624 15695 85742 15705
rect 85624 15567 85742 15577
rect 67431 14533 67559 14542
rect 66754 13990 66882 13999
rect 66754 -1842 66882 13862
rect 66748 -1970 66754 -1842
rect 66882 -1970 66888 -1842
rect 67103 -2039 67170 -2029
rect 67103 -2675 67170 -2665
rect 66560 -5627 66627 -5617
rect 66560 -6263 66627 -6253
rect 67121 -6683 67249 -6674
rect 67431 -6683 67559 14405
rect 71868 12348 71996 12357
rect 71868 -2037 71996 12220
rect 71868 -2175 71996 -2165
rect 72410 11809 72538 11818
rect 72410 -2044 72538 11681
rect 72410 -2182 72538 -2172
rect 72954 11260 73082 11269
rect 72954 -2047 73082 11132
rect 72954 -2185 73082 -2175
rect 73498 10738 73626 10747
rect 73498 -2048 73626 10610
rect 75124 9086 75252 9095
rect 75124 -2036 75252 8958
rect 75670 8552 75798 8561
rect 75670 -2021 75798 8424
rect 75124 -2174 75252 -2164
rect 75669 -2031 75798 -2021
rect 75797 -2090 75798 -2031
rect 76211 8003 76339 8012
rect 76211 -2033 76339 7875
rect 76759 7464 76887 7473
rect 76759 -2023 76887 7336
rect 75669 -2169 75797 -2159
rect 76211 -2171 76339 -2161
rect 76758 -2033 76887 -2023
rect 76886 -2118 76887 -2033
rect 79476 5833 79604 5842
rect 79476 -2029 79604 5705
rect 76758 -2171 76886 -2161
rect 79476 -2167 79604 -2157
rect 80020 5294 80148 5303
rect 80020 -2031 80148 5166
rect 80562 4742 80690 4751
rect 80562 -2019 80690 4614
rect 81106 4194 81234 4203
rect 80562 -2029 80691 -2019
rect 80562 -2100 80563 -2029
rect 80020 -2169 80148 -2159
rect 80563 -2167 80691 -2157
rect 81106 -2031 81234 4066
rect 82748 2566 82876 2575
rect 82748 -2012 82876 2438
rect 83289 2016 83417 2025
rect 82748 -2022 82877 -2012
rect 82748 -2136 82749 -2022
rect 81106 -2169 81234 -2159
rect 82749 -2160 82877 -2150
rect 83289 -2027 83417 1888
rect 83289 -2165 83417 -2155
rect 83830 1471 83958 1480
rect 83830 -2029 83958 1343
rect 84369 948 84497 957
rect 84369 -2012 84497 820
rect 133764 627 133773 687
rect 133833 627 133842 687
rect 132897 -49 132953 -45
rect 132572 -54 132958 -49
rect 132572 -101 132897 -54
rect 132456 -167 132465 -101
rect 132531 -110 132897 -101
rect 132953 -110 132958 -54
rect 132531 -115 132958 -110
rect 132531 -167 132638 -115
rect 132897 -119 132953 -115
rect 133777 -151 133829 627
rect 134341 350 134401 359
rect 134341 281 134401 290
rect 133151 -264 133217 -254
rect 133078 -266 133151 -264
rect 132572 -332 133151 -266
rect 132572 -399 132638 -332
rect 133151 -342 133217 -332
rect 133290 -272 133356 -262
rect 133290 -376 133356 -340
rect 132458 -465 132467 -399
rect 132533 -465 132638 -399
rect 132812 -442 133356 -376
rect 132812 -666 132878 -442
rect 132458 -732 132467 -666
rect 132533 -732 132878 -666
rect 132897 -1366 132953 -1362
rect 132572 -1371 132958 -1366
rect 132572 -1418 132897 -1371
rect 132456 -1484 132465 -1418
rect 132531 -1427 132897 -1418
rect 132953 -1427 132958 -1371
rect 132531 -1432 132958 -1427
rect 132531 -1484 132638 -1432
rect 132897 -1436 132953 -1432
rect 133777 -1468 133829 -203
rect 134067 -214 134133 -204
rect 134067 -292 134133 -282
rect 134200 -216 134313 -206
rect 134200 -294 134313 -284
rect 134345 -274 134397 281
rect 135402 33 135875 43
rect 135402 -46 135875 -36
rect 141764 -188 141853 -171
rect 141764 -248 141779 -188
rect 141839 -248 141853 -188
rect 143472 -190 143532 -188
rect 143465 -246 143474 -190
rect 143530 -246 143539 -190
rect 141764 -263 141853 -248
rect 133777 -1530 133829 -1520
rect 134067 -1531 134133 -1521
rect 133151 -1581 133217 -1571
rect 133078 -1583 133151 -1581
rect 132572 -1649 133151 -1583
rect 132572 -1716 132638 -1649
rect 133151 -1659 133217 -1649
rect 133290 -1589 133356 -1579
rect 134067 -1609 134133 -1599
rect 134200 -1533 134313 -1523
rect 134200 -1611 134313 -1601
rect 134345 -1591 134397 -326
rect 139082 -513 139544 -503
rect 139082 -587 139544 -577
rect 135405 -1282 135878 -1272
rect 135405 -1361 135878 -1351
rect 141764 -1505 141853 -1488
rect 141764 -1565 141779 -1505
rect 141839 -1565 141853 -1505
rect 143166 -1507 143226 -1505
rect 143159 -1563 143168 -1507
rect 143224 -1563 143233 -1507
rect 141764 -1580 141853 -1565
rect 134345 -1653 134397 -1643
rect 133290 -1693 133356 -1657
rect 132458 -1782 132467 -1716
rect 132533 -1782 132638 -1716
rect 132812 -1759 133356 -1693
rect 132812 -1983 132878 -1759
rect 139092 -1827 139554 -1817
rect 139092 -1901 139554 -1891
rect 84369 -2022 84498 -2012
rect 84369 -2088 84370 -2022
rect 83830 -2167 83958 -2157
rect 132458 -2049 132467 -1983
rect 132533 -2049 132878 -1983
rect 84370 -2160 84498 -2150
rect 73498 -2186 73626 -2176
rect 133764 -2337 133773 -2277
rect 133833 -2337 133842 -2277
rect 132897 -3013 132953 -3009
rect 132572 -3018 132958 -3013
rect 132572 -3065 132897 -3018
rect 132456 -3131 132465 -3065
rect 132531 -3074 132897 -3065
rect 132953 -3074 132958 -3018
rect 132531 -3079 132958 -3074
rect 132531 -3131 132638 -3079
rect 132897 -3083 132953 -3079
rect 133777 -3115 133829 -2337
rect 134341 -2614 134401 -2605
rect 134341 -2683 134401 -2674
rect 133151 -3228 133217 -3218
rect 133078 -3230 133151 -3228
rect 132572 -3296 133151 -3230
rect 132572 -3363 132638 -3296
rect 133151 -3306 133217 -3296
rect 133290 -3236 133356 -3226
rect 133290 -3340 133356 -3304
rect 132458 -3429 132467 -3363
rect 132533 -3429 132638 -3363
rect 132812 -3406 133356 -3340
rect 132812 -3630 132878 -3406
rect 132458 -3696 132467 -3630
rect 132533 -3696 132878 -3630
rect 132897 -4260 132953 -4256
rect 132572 -4265 132958 -4260
rect 132572 -4312 132897 -4265
rect 132456 -4378 132465 -4312
rect 132531 -4321 132897 -4312
rect 132953 -4321 132958 -4265
rect 132531 -4326 132958 -4321
rect 132531 -4378 132638 -4326
rect 132897 -4330 132953 -4326
rect 133777 -4362 133829 -3167
rect 134067 -3178 134133 -3168
rect 134067 -3256 134133 -3246
rect 134200 -3180 134313 -3170
rect 134200 -3258 134313 -3248
rect 134345 -3238 134397 -2683
rect 135397 -2928 135870 -2918
rect 135397 -3007 135870 -2997
rect 141764 -3152 141853 -3135
rect 141764 -3212 141779 -3152
rect 141839 -3212 141853 -3152
rect 142774 -3154 142834 -3152
rect 142767 -3210 142776 -3154
rect 142832 -3210 142841 -3154
rect 141764 -3227 141853 -3212
rect 133777 -4424 133829 -4414
rect 134067 -4425 134133 -4415
rect 133151 -4475 133217 -4465
rect 133078 -4477 133151 -4475
rect 132572 -4543 133151 -4477
rect 132572 -4610 132638 -4543
rect 133151 -4553 133217 -4543
rect 133290 -4483 133356 -4473
rect 134067 -4503 134133 -4493
rect 134200 -4427 134313 -4417
rect 134200 -4505 134313 -4495
rect 134345 -4485 134397 -3290
rect 139082 -3477 139544 -3467
rect 139082 -3551 139544 -3541
rect 135399 -4178 135872 -4168
rect 135399 -4257 135872 -4247
rect 141764 -4399 141853 -4382
rect 141764 -4459 141779 -4399
rect 141839 -4459 141853 -4399
rect 142368 -4401 142428 -4399
rect 142361 -4457 142370 -4401
rect 142426 -4457 142435 -4401
rect 141764 -4474 141853 -4459
rect 134345 -4547 134397 -4537
rect 133290 -4587 133356 -4551
rect 132458 -4676 132467 -4610
rect 132533 -4676 132638 -4610
rect 132812 -4653 133356 -4587
rect 132812 -4877 132878 -4653
rect 139097 -4724 139559 -4714
rect 139097 -4798 139559 -4788
rect 132458 -4943 132467 -4877
rect 132533 -4943 132878 -4877
rect 71081 -5629 71140 -5619
rect 71081 -6277 71140 -6267
rect 74345 -5629 74404 -5619
rect 74345 -6277 74404 -6267
rect 77609 -5629 77668 -5619
rect 77609 -6277 77668 -6267
rect 78697 -5629 78756 -5619
rect 78697 -6277 78756 -6267
rect 81961 -5629 82020 -5619
rect 81961 -6277 82020 -6267
rect 85225 -5629 85284 -5619
rect 85225 -6277 85284 -6267
rect 66840 -6811 66846 -6683
rect 66974 -6811 67121 -6683
rect 67249 -6811 67559 -6683
rect 67121 -6820 67249 -6811
rect 71628 -8627 71687 -8617
rect 71628 -9275 71687 -9265
rect 72716 -8627 72775 -8617
rect 72716 -9275 72775 -9265
rect 73804 -8627 73863 -8617
rect 73804 -9275 73863 -9265
rect 74892 -8627 74951 -8617
rect 74892 -9275 74951 -9265
rect 75980 -8627 76039 -8617
rect 75980 -9275 76039 -9265
rect 77068 -8627 77127 -8617
rect 77068 -9275 77127 -9265
rect 78156 -8627 78215 -8617
rect 78156 -9275 78215 -9265
rect 79244 -8627 79303 -8617
rect 79244 -9275 79303 -9265
rect 80332 -8627 80391 -8617
rect 80332 -9275 80391 -9265
rect 81420 -8627 81479 -8617
rect 81420 -9275 81479 -9265
rect 82508 -8627 82567 -8617
rect 82508 -9275 82567 -9265
rect 83596 -8627 83655 -8617
rect 83596 -9275 83655 -9265
rect 84684 -8627 84743 -8617
rect 84684 -9275 84743 -9265
rect 142368 -11863 142428 -4457
rect 142774 -11597 142834 -3210
rect 143166 -11297 143226 -1563
rect 143472 -11030 143532 -246
rect 143472 -11039 143534 -11030
rect 143472 -11046 143478 -11039
rect 143478 -11104 143534 -11095
rect 147329 -11156 147802 -11146
rect 144829 -11241 144885 -11237
rect 144504 -11246 144890 -11241
rect 144504 -11293 144829 -11246
rect 143166 -11353 143168 -11297
rect 143224 -11353 143226 -11297
rect 143166 -11364 143226 -11353
rect 144388 -11359 144397 -11293
rect 144463 -11302 144829 -11293
rect 144885 -11302 144890 -11246
rect 144463 -11307 144890 -11302
rect 144463 -11359 144570 -11307
rect 144829 -11311 144885 -11307
rect 145709 -11343 145761 -11208
rect 145083 -11456 145149 -11446
rect 145010 -11458 145083 -11456
rect 144504 -11524 145083 -11458
rect 144504 -11591 144570 -11524
rect 145083 -11534 145149 -11524
rect 145222 -11464 145288 -11454
rect 145222 -11568 145288 -11532
rect 142774 -11638 142778 -11597
rect 142778 -11662 142834 -11653
rect 144390 -11657 144399 -11591
rect 144465 -11657 144570 -11591
rect 144744 -11634 145288 -11568
rect 144744 -11858 144810 -11634
rect 142424 -11919 142428 -11863
rect 142368 -11928 142428 -11919
rect 144390 -11924 144399 -11858
rect 144465 -11924 144810 -11858
rect 145709 -12190 145761 -11395
rect 145999 -11406 146065 -11396
rect 145999 -11484 146065 -11474
rect 146132 -11408 146245 -11398
rect 146132 -11486 146245 -11476
rect 146277 -11466 146329 -11208
rect 147329 -11235 147802 -11225
rect 153848 -11380 153900 -11378
rect 153835 -11440 153844 -11380
rect 153904 -11440 153913 -11380
rect 153848 -11442 153900 -11440
rect 145696 -12250 145705 -12190
rect 145765 -12250 145774 -12190
rect 146277 -12620 146329 -11518
rect 151014 -11705 151476 -11695
rect 151014 -11779 151476 -11769
rect 146264 -12680 146273 -12620
rect 146333 -12680 146342 -12620
rect 71079 -13627 71138 -13617
rect 71079 -14275 71138 -14265
rect 72167 -13627 72226 -13617
rect 72167 -14275 72226 -14265
rect 73255 -13627 73314 -13617
rect 73255 -14275 73314 -14265
rect 74343 -13627 74402 -13617
rect 74343 -14275 74402 -14265
rect 75431 -13627 75490 -13617
rect 75431 -14275 75490 -14265
rect 76519 -13627 76578 -13617
rect 76519 -14275 76578 -14265
rect 77607 -13627 77666 -13617
rect 77607 -14275 77666 -14265
rect 78695 -13627 78754 -13617
rect 78695 -14275 78754 -14265
rect 79783 -13627 79842 -13617
rect 79783 -14275 79842 -14265
rect 80871 -13627 80930 -13617
rect 80871 -14275 80930 -14265
rect 81959 -13627 82018 -13617
rect 81959 -14275 82018 -14265
rect 83047 -13627 83106 -13617
rect 83047 -14275 83106 -14265
rect 84135 -13627 84194 -13617
rect 84135 -14275 84194 -14265
rect 85223 -13627 85282 -13617
rect 85223 -14275 85282 -14265
rect 71621 -16617 71685 -16607
rect 71621 -17281 71685 -17271
rect 72709 -16617 72773 -16607
rect 72709 -17281 72773 -17271
rect 73797 -16617 73861 -16607
rect 73797 -17281 73861 -17271
rect 74885 -16617 74949 -16607
rect 74885 -17281 74949 -17271
rect 75973 -16617 76037 -16607
rect 75973 -17281 76037 -17271
rect 77061 -16617 77125 -16607
rect 77061 -17281 77125 -17271
rect 78149 -16617 78213 -16607
rect 78149 -17281 78213 -17271
rect 79237 -16617 79301 -16607
rect 79237 -17281 79301 -17271
rect 80325 -16617 80389 -16607
rect 80325 -17281 80389 -17271
rect 81413 -16617 81477 -16607
rect 81413 -17281 81477 -17271
rect 82501 -16617 82565 -16607
rect 82501 -17281 82565 -17271
rect 83589 -16617 83653 -16607
rect 83589 -17281 83653 -17271
rect 84677 -16617 84741 -16607
rect 84677 -17281 84741 -17271
rect 71075 -21612 71142 -21602
rect 71075 -22016 71142 -22006
rect 72165 -21618 72232 -21608
rect 72165 -22022 72232 -22012
rect 73253 -21618 73320 -21608
rect 73253 -22022 73320 -22012
rect 74341 -21618 74408 -21608
rect 74341 -22022 74408 -22012
rect 75429 -21618 75496 -21608
rect 75429 -22022 75496 -22012
rect 76517 -21618 76584 -21608
rect 76517 -22022 76584 -22012
rect 77605 -21618 77672 -21608
rect 77605 -22022 77672 -22012
rect 81957 -21618 82024 -21608
rect 81957 -22022 82024 -22012
rect 83045 -21618 83112 -21608
rect 83045 -22022 83112 -22012
rect 84133 -21618 84200 -21608
rect 84133 -22022 84200 -22012
rect 85221 -21618 85288 -21608
rect 85221 -22022 85288 -22012
rect 77469 -22175 78509 -22160
rect 77469 -23175 77491 -22175
rect 78491 -23175 78509 -22175
rect 77469 -23196 78509 -23175
<< via2 >>
rect 36373 70835 37373 71835
rect 43364 70817 44364 71817
rect 57809 70821 58809 71821
rect 64881 70771 65881 71771
rect 74883 70807 75883 71807
rect 85758 70759 86758 71759
rect 94068 70783 95068 71783
rect 103408 70867 104408 71867
rect 35285 67107 35410 70423
rect 38294 67113 38442 70399
rect 42295 67110 42410 70392
rect 45277 67092 45431 70421
rect 56700 67113 56848 70393
rect 59712 67113 59864 70398
rect 63788 67105 63951 70396
rect 66804 67117 66952 70395
rect 73794 67107 73935 70398
rect 76799 67113 76934 70396
rect 84670 67112 84798 70393
rect 87663 67108 87817 70406
rect 92977 67100 93119 70406
rect 95985 67112 96113 70403
rect 102317 67100 102459 70406
rect 105325 67112 105453 70403
rect 36406 50533 36466 50593
rect 46449 52576 46509 52636
rect 46153 51695 46271 52282
rect 48449 52573 48509 52633
rect 38404 50535 38464 50595
rect 36202 49483 36285 49927
rect 37447 49792 37567 50285
rect 38144 49278 38243 49857
rect 37227 48967 37287 49027
rect 39493 49780 39608 50313
rect 39227 48956 39287 49016
rect 47493 51229 47608 51852
rect 48197 51690 48307 52230
rect 49511 51249 49654 51907
rect 62908 64980 63133 65047
rect 63684 64989 63797 65102
rect 64232 64976 64460 65055
rect 65058 64998 65171 65111
rect 65616 64980 65843 65055
rect 66421 64998 66534 65111
rect 66997 64982 67225 65054
rect 67770 64999 67883 65112
rect 72908 64980 73133 65047
rect 73684 64989 73797 65102
rect 74232 64976 74460 65055
rect 75058 64998 75171 65111
rect 75616 64980 75843 65055
rect 76421 64998 76534 65111
rect 76997 64982 77225 65054
rect 77770 64999 77883 65112
rect 61524 64026 61642 64144
rect 60901 62821 61009 62929
rect 71637 64018 71755 64136
rect 84180 64021 84288 64129
rect 62129 63422 62247 63540
rect 71110 62821 71218 62929
rect 62731 62076 62844 62189
rect 63429 62033 63542 62146
rect 64378 62045 64491 62159
rect 64721 62064 64834 62177
rect 65456 62056 65569 62169
rect 66175 62038 66288 62151
rect 66828 62030 66941 62143
rect 67543 62038 67656 62151
rect 63163 61245 63234 61352
rect 63705 61242 63776 61346
rect 65884 61349 65952 61473
rect 64251 61184 64320 61330
rect 64798 61191 64862 61321
rect 66426 61207 66494 61364
rect 66971 61261 67043 61383
rect 67514 61202 67580 61356
rect 65343 60862 65410 61015
rect 72122 63421 72240 63539
rect 72731 62076 72844 62189
rect 73429 62033 73542 62146
rect 74378 62045 74491 62159
rect 74721 62064 74834 62177
rect 75456 62056 75569 62169
rect 76175 62038 76288 62151
rect 76828 62030 76941 62143
rect 77543 62038 77656 62151
rect 73163 61245 73234 61352
rect 73705 61242 73776 61346
rect 75884 61349 75952 61473
rect 74251 61184 74320 61330
rect 74798 61191 74862 61321
rect 76426 61207 76494 61364
rect 76971 61261 77043 61383
rect 77514 61202 77580 61356
rect 75343 60862 75410 61015
rect 85128 63757 85318 63849
rect 85568 63736 86002 63823
rect 86485 63764 86629 63858
rect 86904 63732 87328 63809
rect 88038 62821 88146 62929
rect 85219 62237 85311 62346
rect 86550 62232 86642 62341
rect 86094 60357 86159 60499
rect 85544 60170 85615 60274
rect 86636 60170 86704 60280
rect 63052 59916 63305 59993
rect 64372 59915 64680 60000
rect 65760 59918 66042 59989
rect 67132 59920 67414 59991
rect 73052 59916 73305 59993
rect 74372 59915 74680 60000
rect 75760 59918 76042 59989
rect 77132 59920 77414 59991
rect 84943 59523 85056 59636
rect 63937 59238 64050 59351
rect 65298 59250 65411 59363
rect 66660 59268 66773 59381
rect 68044 59303 68157 59416
rect 73937 59238 74050 59351
rect 75298 59250 75411 59363
rect 76660 59268 76773 59381
rect 78044 59303 78157 59416
rect 87336 58917 87449 59030
rect 58764 52103 58820 52159
rect 62501 54651 62618 54768
rect 63317 51978 63513 52174
rect 61623 51529 61744 51650
rect 62506 51556 62613 51663
rect 66038 51482 66234 51678
rect 47273 50822 47343 50892
rect 74726 54656 74833 54763
rect 49271 50830 49331 50890
rect 61618 50256 61749 50387
rect 66174 50013 66362 50207
rect 67970 49987 68198 50219
rect 69664 49968 69892 50200
rect 71483 49979 71711 50211
rect 73267 49976 73495 50208
rect 75052 49974 75280 50206
rect 62848 49465 63380 49622
rect 65284 48532 65560 48632
rect 67154 48584 67390 48662
rect 68959 48576 69193 48655
rect 70765 48570 70984 48651
rect 72551 48571 72791 48655
rect 74352 48586 74604 48651
rect 56046 46741 56330 47379
rect 60492 47109 61496 47309
rect 62501 47157 62618 47274
rect 58762 45782 58822 45842
rect 36693 40477 36821 40605
rect 62010 41599 62280 42674
rect 62857 41596 63127 42671
rect 63412 41747 63617 42335
rect 44965 40400 45093 40528
rect 56027 38731 56167 39355
rect 65328 37035 65572 37235
rect 66930 37046 67174 37246
rect 68833 37106 69077 37306
rect 70550 37090 70794 37290
rect 72364 37085 72608 37285
rect 74336 37079 74580 37279
rect 65850 35656 66234 35734
rect 67641 35667 68041 35741
rect 69447 35667 69835 35741
rect 71244 35632 71632 35706
rect 73046 35628 73433 35706
rect 74840 35625 75235 35702
rect 67555 34952 67663 35060
rect 35200 34159 35318 34277
rect 44805 34155 44913 34263
rect 40661 32525 40779 32643
rect 36513 31027 36631 31145
rect 42143 30948 42261 31066
rect 41228 23742 41356 23870
rect 41701 23526 41765 23590
rect 39914 22711 39978 22775
rect 40383 22450 40511 22578
rect 36843 21755 36971 21883
rect 38308 21522 38372 21586
rect 36278 20709 36342 20773
rect 37638 20451 37766 20579
rect 36843 19757 36971 19885
rect 38307 19528 38371 19592
rect 67550 33303 67668 33421
rect 50238 32549 50356 32667
rect 45534 27510 45652 27628
rect 55952 30754 56299 31354
rect 60986 29648 61191 30188
rect 64046 29124 64252 29330
rect 59363 28460 61033 28687
rect 43434 21534 43562 21662
rect 44375 21343 44431 21399
rect 43010 20518 43074 20582
rect 44260 20269 44388 20397
rect 51068 23721 51186 23839
rect 52551 23516 52615 23580
rect 43415 19526 43543 19654
rect 44369 19399 44433 19402
rect 44369 19338 44431 19399
rect 44431 19338 44433 19399
rect 50506 22704 50570 22768
rect 51940 22469 52058 22587
rect 47795 21719 47923 21847
rect 48704 21583 48768 21584
rect 48704 21520 48766 21583
rect 48766 21520 48768 21583
rect 36280 18707 36344 18771
rect 37633 18450 37761 18578
rect 40397 17738 40525 17866
rect 41702 17523 41766 17587
rect 43413 18522 43469 18578
rect 44259 18261 44387 18389
rect 47737 20703 47801 20767
rect 48603 20449 48731 20577
rect 47791 19714 47919 19842
rect 49357 19518 49421 19582
rect 47735 18697 47737 18761
rect 47737 18697 47799 18761
rect 48603 18450 48731 18578
rect 81000 41367 81064 41431
rect 79904 40461 79983 40739
rect 101834 64021 101942 64129
rect 102782 63757 102972 63849
rect 103222 63736 103656 63823
rect 104139 63764 104283 63858
rect 104558 63732 104982 63809
rect 105692 62821 105800 62929
rect 102873 62237 102965 62346
rect 104204 62232 104296 62341
rect 103748 60357 103813 60499
rect 103198 60170 103269 60274
rect 104290 60170 104358 60280
rect 102597 59523 102710 59636
rect 104990 58917 105103 59030
rect 85593 43173 85657 43237
rect 100698 50019 100886 50213
rect 102494 49993 102722 50225
rect 104188 49974 104416 50206
rect 106007 49985 106235 50217
rect 107791 49982 108019 50214
rect 109576 49980 109804 50212
rect 96364 49432 97874 49834
rect 99808 48538 100084 48638
rect 101678 48590 101914 48668
rect 103483 48582 103717 48661
rect 105289 48576 105508 48657
rect 107075 48577 107315 48661
rect 108876 48592 109128 48657
rect 90796 46782 91108 47320
rect 94987 47083 96094 47300
rect 87594 43173 87658 43237
rect 84505 42267 84628 42609
rect 86529 42262 86618 42646
rect 84767 41664 84831 41728
rect 83000 41376 83064 41440
rect 81965 40420 82045 40703
rect 80175 39857 80239 39921
rect 82166 39849 82240 39923
rect 81167 39581 81285 39699
rect 83018 39595 83142 39719
rect 86765 41667 86829 41731
rect 85888 41010 86114 41236
rect 96525 41606 96795 42681
rect 97372 41603 97642 42678
rect 97972 41682 98218 42396
rect 87813 41017 88014 41218
rect 90783 38091 91030 38958
rect 83785 34762 83913 34890
rect 83651 33674 83769 33792
rect 82680 33459 82736 33515
rect 82310 33032 82438 33160
rect 62988 23722 63106 23840
rect 64445 23519 64509 23583
rect 62420 22696 62484 22760
rect 63860 22464 63978 22582
rect 60239 21753 60357 21871
rect 61664 21520 61728 21584
rect 59698 20699 59762 20763
rect 61061 20461 61179 20579
rect 60241 19723 60359 19841
rect 61667 19517 61731 19581
rect 51104 17722 51222 17840
rect 52547 17516 52611 17580
rect 59710 18700 59774 18764
rect 61055 18465 61173 18583
rect 63015 17715 63133 17833
rect 63942 17518 64006 17582
rect 67161 20731 67225 20795
rect 67989 20728 68053 20792
rect 66649 20214 66767 20332
rect 68386 20206 68504 20324
rect 67163 19761 67227 19825
rect 67985 19762 68049 19826
rect 85011 33456 85067 33512
rect 82676 31999 82740 32063
rect 81964 31759 82082 31877
rect 99844 37028 100088 37228
rect 101446 37039 101690 37239
rect 103349 37099 103593 37299
rect 105066 37083 105310 37283
rect 106880 37078 107124 37278
rect 108852 37072 109096 37272
rect 96849 35740 97596 35851
rect 100366 35649 100750 35727
rect 102157 35660 102557 35734
rect 103963 35660 104351 35734
rect 105760 35625 106148 35699
rect 107562 35621 107949 35699
rect 109356 35618 109751 35695
rect 89492 35336 89688 35532
rect 86373 35197 86501 35325
rect 88561 34183 88757 34379
rect 95270 34183 95466 34379
rect 85321 33039 85449 33167
rect 71557 23719 71675 23837
rect 72875 23523 72939 23587
rect 84971 31696 85089 31814
rect 85799 31723 85907 31831
rect 82236 31222 82344 31330
rect 71186 22697 71250 22761
rect 72435 22460 72553 22578
rect 74028 20481 74092 20545
rect 74856 20487 74920 20551
rect 73565 19952 73683 20070
rect 75276 19975 75394 20093
rect 74034 19519 74098 19583
rect 74860 19518 74924 19582
rect 71584 17726 71702 17844
rect 72882 17530 72946 17594
rect 86666 31701 86784 31819
rect 86377 24870 86495 24988
rect 85212 24663 85276 24727
rect 87019 23838 87083 23902
rect 83055 23654 83173 23772
rect 85591 23604 85709 23722
rect 81877 23474 81941 23538
rect 83459 22647 83523 22711
rect 82256 22404 82374 22522
rect 82968 17695 83086 17813
rect 81882 17503 81946 17567
rect 116738 52386 116866 52514
rect 120662 52363 120933 52467
rect 115289 51273 115385 51725
rect 117729 51316 117832 51778
rect 119326 51001 119407 52130
rect 121709 51027 121804 52123
rect 115579 50800 115707 50928
rect 115989 50709 116141 50861
rect 117396 50869 117553 50953
rect 119936 50772 120225 50944
rect 121196 50888 121516 50958
rect 114709 38737 115008 39378
rect 123011 37052 123095 38345
rect 123011 35592 123095 36885
rect 123012 34387 123095 35405
rect 95427 30789 95711 31246
rect 90814 30288 91056 30752
rect 95203 28464 95762 28684
rect 125028 33811 125348 34131
rect 128031 33937 129021 34927
rect 123010 32643 123097 33617
rect 127217 33666 127594 33739
rect 127219 32552 127591 32617
rect 114716 30726 115015 31367
rect 123007 31104 123097 32470
rect 123008 29606 123099 30864
rect 124329 30866 124649 31186
rect 104393 27054 104511 27172
rect 107956 27067 108074 27185
rect 93840 26820 94036 27016
rect 92590 23670 92708 23788
rect 93136 23473 93200 23537
rect 91392 22648 91456 22712
rect 91882 22410 92000 22528
rect 92566 17701 92684 17819
rect 92782 17565 92846 17567
rect 92782 17503 92844 17565
rect 92844 17503 92846 17565
rect 106372 23300 106500 23428
rect 105422 23096 105486 23160
rect 104398 22562 104506 22670
rect 107984 22581 108092 22689
rect 107095 22276 107169 22350
rect 105796 22028 105924 22156
rect 39911 16701 39975 16765
rect 50503 16698 50567 16762
rect 62421 16699 62485 16763
rect 71190 16710 71254 16774
rect 41211 16414 41339 16542
rect 51817 16464 51935 16582
rect 63827 16455 63945 16573
rect 72296 16464 72414 16582
rect 86412 16844 86530 16962
rect 83455 16683 83519 16747
rect 85210 16653 85274 16717
rect 82296 16443 82414 16561
rect 91402 16679 91466 16743
rect 91859 16429 91977 16547
rect 87016 15828 87080 15892
rect 85624 15577 85742 15695
rect 67431 14405 67559 14533
rect 66754 13862 66882 13990
rect 67103 -2665 67170 -2039
rect 66560 -6253 66627 -5627
rect 71868 12220 71996 12348
rect 72410 11681 72538 11809
rect 72954 11132 73082 11260
rect 73498 10610 73626 10738
rect 75124 8958 75252 9086
rect 75670 8424 75798 8552
rect 76211 7875 76339 8003
rect 76759 7336 76887 7464
rect 79476 5705 79604 5833
rect 80020 5166 80148 5294
rect 80562 4614 80690 4742
rect 81106 4066 81234 4194
rect 82748 2438 82876 2566
rect 83289 1888 83417 2016
rect 83830 1343 83958 1471
rect 84369 820 84497 948
rect 133773 627 133833 687
rect 132465 -167 132531 -101
rect 132897 -110 132953 -54
rect 134341 290 134401 350
rect 132467 -465 132533 -399
rect 132467 -732 132533 -666
rect 132465 -1484 132531 -1418
rect 132897 -1427 132953 -1371
rect 134067 -282 134133 -214
rect 134247 -284 134266 -216
rect 134266 -284 134313 -216
rect 135402 -36 135875 33
rect 141779 -192 141839 -188
rect 141779 -244 141783 -192
rect 141783 -244 141835 -192
rect 141835 -244 141839 -192
rect 141779 -248 141839 -244
rect 143474 -246 143530 -190
rect 134067 -1599 134133 -1531
rect 134247 -1601 134266 -1533
rect 134266 -1601 134313 -1533
rect 139082 -577 139544 -513
rect 135405 -1351 135878 -1282
rect 141779 -1509 141839 -1505
rect 141779 -1561 141783 -1509
rect 141783 -1561 141835 -1509
rect 141835 -1561 141839 -1509
rect 141779 -1565 141839 -1561
rect 143168 -1563 143224 -1507
rect 132467 -1782 132533 -1716
rect 139092 -1891 139554 -1827
rect 132467 -2049 132533 -1983
rect 133773 -2337 133833 -2277
rect 132465 -3131 132531 -3065
rect 132897 -3074 132953 -3018
rect 134341 -2674 134401 -2614
rect 132467 -3429 132533 -3363
rect 132467 -3696 132533 -3630
rect 132465 -4378 132531 -4312
rect 132897 -4321 132953 -4265
rect 134067 -3246 134133 -3178
rect 134247 -3248 134266 -3180
rect 134266 -3248 134313 -3180
rect 135397 -2997 135870 -2928
rect 141779 -3156 141839 -3152
rect 141779 -3208 141783 -3156
rect 141783 -3208 141835 -3156
rect 141835 -3208 141839 -3156
rect 141779 -3212 141839 -3208
rect 142776 -3210 142832 -3154
rect 134067 -4493 134133 -4425
rect 134247 -4495 134266 -4427
rect 134266 -4495 134313 -4427
rect 139082 -3541 139544 -3477
rect 135399 -4247 135872 -4178
rect 141779 -4403 141839 -4399
rect 141779 -4455 141783 -4403
rect 141783 -4455 141835 -4403
rect 141835 -4455 141839 -4403
rect 141779 -4459 141839 -4455
rect 142370 -4457 142426 -4401
rect 132467 -4676 132533 -4610
rect 139097 -4788 139559 -4724
rect 132467 -4943 132533 -4877
rect 71081 -6267 71140 -5629
rect 74345 -6267 74404 -5629
rect 77609 -6267 77668 -5629
rect 78697 -6267 78756 -5629
rect 81961 -6267 82020 -5629
rect 85225 -6267 85284 -5629
rect 67121 -6811 67249 -6683
rect 71628 -9265 71687 -8627
rect 72716 -9265 72775 -8627
rect 73804 -9265 73863 -8627
rect 74892 -9265 74951 -8627
rect 75980 -9265 76039 -8627
rect 77068 -9265 77127 -8627
rect 78156 -9265 78215 -8627
rect 79244 -9265 79303 -8627
rect 80332 -9265 80391 -8627
rect 81420 -9265 81479 -8627
rect 82508 -9265 82567 -8627
rect 83596 -9265 83655 -8627
rect 84684 -9265 84743 -8627
rect 143478 -11095 143534 -11039
rect 143168 -11353 143224 -11297
rect 144397 -11359 144463 -11293
rect 144829 -11302 144885 -11246
rect 142778 -11653 142834 -11597
rect 144399 -11657 144465 -11591
rect 142368 -11919 142424 -11863
rect 144399 -11924 144465 -11858
rect 145999 -11474 146065 -11406
rect 146179 -11476 146198 -11408
rect 146198 -11476 146245 -11408
rect 147329 -11225 147802 -11156
rect 153844 -11384 153904 -11380
rect 153844 -11436 153848 -11384
rect 153848 -11436 153900 -11384
rect 153900 -11436 153904 -11384
rect 153844 -11440 153904 -11436
rect 145705 -12250 145765 -12190
rect 151014 -11769 151476 -11705
rect 146273 -12680 146333 -12620
rect 71079 -14265 71138 -13627
rect 72167 -14265 72226 -13627
rect 73255 -14265 73314 -13627
rect 74343 -14265 74402 -13627
rect 75431 -14265 75490 -13627
rect 76519 -14265 76578 -13627
rect 77607 -14265 77666 -13627
rect 78695 -14265 78754 -13627
rect 79783 -14265 79842 -13627
rect 80871 -14265 80930 -13627
rect 81959 -14265 82018 -13627
rect 83047 -14265 83106 -13627
rect 84135 -14265 84194 -13627
rect 85223 -14265 85282 -13627
rect 71621 -17271 71685 -16617
rect 72709 -17271 72773 -16617
rect 73797 -17271 73861 -16617
rect 74885 -17271 74949 -16617
rect 75973 -17271 76037 -16617
rect 77061 -17271 77125 -16617
rect 78149 -17271 78213 -16617
rect 79237 -17271 79301 -16617
rect 80325 -17271 80389 -16617
rect 81413 -17271 81477 -16617
rect 82501 -17271 82565 -16617
rect 83589 -17271 83653 -16617
rect 84677 -17271 84741 -16617
rect 71075 -22006 71142 -21612
rect 72165 -22012 72232 -21618
rect 73253 -22012 73320 -21618
rect 74341 -22012 74408 -21618
rect 75429 -22012 75496 -21618
rect 76517 -22012 76584 -21618
rect 77605 -22012 77672 -21618
rect 81957 -22012 82024 -21618
rect 83045 -22012 83112 -21618
rect 84133 -22012 84200 -21618
rect 85221 -22012 85288 -21618
rect 77491 -23175 78491 -22175
<< metal3 >>
rect 36373 71840 37373 91353
rect 36368 71835 37378 71840
rect 36368 70835 36373 71835
rect 37373 70835 37378 71835
rect 43364 71822 44364 91353
rect 57809 71826 58809 91353
rect 36368 70830 37378 70835
rect 43359 71817 44369 71822
rect 43359 70817 43364 71817
rect 44364 70817 44369 71817
rect 43359 70812 44369 70817
rect 57804 71821 58814 71826
rect 57804 70821 57809 71821
rect 58809 70821 58814 71821
rect 64881 71776 65881 91353
rect 74883 71812 75883 91353
rect 74878 71807 75888 71812
rect 57804 70816 58814 70821
rect 64876 71771 65886 71776
rect 64876 70771 64881 71771
rect 65881 70771 65886 71771
rect 74878 70807 74883 71807
rect 75883 70807 75888 71807
rect 85758 71764 86758 91353
rect 94068 71788 95068 91353
rect 103408 71872 104408 91353
rect 103403 71867 104413 71872
rect 94063 71783 95073 71788
rect 74878 70802 75888 70807
rect 85753 71759 86763 71764
rect 64876 70766 65886 70771
rect 85753 70759 85758 71759
rect 86758 70759 86763 71759
rect 94063 70783 94068 71783
rect 95068 70783 95073 71783
rect 103403 70867 103408 71867
rect 104408 70867 104413 71867
rect 103403 70862 104413 70867
rect 94063 70778 95073 70783
rect 85753 70754 86763 70759
rect 112864 70709 113864 91353
rect 114864 70709 115864 91353
rect 116864 70709 117864 91353
rect 35275 70423 35420 70428
rect 35275 67107 35285 70423
rect 35410 67107 35420 70423
rect 45267 70421 45441 70426
rect 38284 70399 38452 70404
rect 38284 67113 38294 70399
rect 38442 67113 38452 70399
rect 38284 67108 38452 67113
rect 42285 70392 42420 70397
rect 42285 67110 42295 70392
rect 42410 67110 42420 70392
rect 35275 67102 35420 67107
rect 42285 67105 42420 67110
rect 45267 67092 45277 70421
rect 45431 67092 45441 70421
rect 87653 70406 87827 70411
rect 59702 70398 59874 70403
rect 56690 70393 56858 70398
rect 56690 67113 56700 70393
rect 56848 67113 56858 70393
rect 56690 67108 56858 67113
rect 59702 67113 59712 70398
rect 59864 67113 59874 70398
rect 59702 67108 59874 67113
rect 63778 70396 63961 70401
rect 63778 67105 63788 70396
rect 63951 67105 63961 70396
rect 66794 70395 66962 70400
rect 66794 67117 66804 70395
rect 66952 67117 66962 70395
rect 66794 67112 66962 67117
rect 73784 70398 73945 70403
rect 63778 67100 63961 67105
rect 73784 67107 73794 70398
rect 73935 67107 73945 70398
rect 76789 70396 76944 70401
rect 76789 67113 76799 70396
rect 76934 67113 76944 70396
rect 76789 67108 76944 67113
rect 84660 70393 84808 70398
rect 84660 67112 84670 70393
rect 84798 67112 84808 70393
rect 84660 67107 84808 67112
rect 87653 67108 87663 70406
rect 87817 67108 87827 70406
rect 73784 67102 73945 67107
rect 87653 67103 87827 67108
rect 92967 70406 93129 70411
rect 92967 67100 92977 70406
rect 93119 67100 93129 70406
rect 95975 70403 96123 70408
rect 95975 67112 95985 70403
rect 96113 67112 96123 70403
rect 95975 67107 96123 67112
rect 102307 70406 102469 70411
rect 92967 67095 93129 67100
rect 102307 67100 102317 70406
rect 102459 67100 102469 70406
rect 105315 70403 105463 70408
rect 105315 67112 105325 70403
rect 105453 67112 105463 70403
rect 105315 67107 105463 67112
rect 102307 67095 102469 67100
rect 45267 67087 45441 67092
rect 65048 65111 65181 65116
rect 63674 65102 63807 65107
rect 62898 65047 63143 65052
rect 62898 64980 62908 65047
rect 63133 64980 63143 65047
rect 63674 64989 63684 65102
rect 63797 64989 63807 65102
rect 63674 64984 63807 64989
rect 64222 65055 64470 65060
rect 62898 64975 63143 64980
rect 64222 64976 64232 65055
rect 64460 64976 64470 65055
rect 65048 64998 65058 65111
rect 65171 64998 65181 65111
rect 66411 65111 66544 65116
rect 65048 64993 65181 64998
rect 65606 65055 65853 65060
rect 64222 64971 64470 64976
rect 65606 64980 65616 65055
rect 65843 64980 65853 65055
rect 66411 64998 66421 65111
rect 66534 64998 66544 65111
rect 67760 65112 67893 65117
rect 66411 64993 66544 64998
rect 66987 65054 67235 65059
rect 65606 64975 65853 64980
rect 66987 64982 66997 65054
rect 67225 64982 67235 65054
rect 67760 64999 67770 65112
rect 67883 64999 67893 65112
rect 75048 65111 75181 65116
rect 73674 65102 73807 65107
rect 67760 64994 67893 64999
rect 72898 65047 73143 65052
rect 66987 64977 67235 64982
rect 72898 64980 72908 65047
rect 73133 64980 73143 65047
rect 73674 64989 73684 65102
rect 73797 64989 73807 65102
rect 73674 64984 73807 64989
rect 74222 65055 74470 65060
rect 72898 64975 73143 64980
rect 74222 64976 74232 65055
rect 74460 64976 74470 65055
rect 75048 64998 75058 65111
rect 75171 64998 75181 65111
rect 76411 65111 76544 65116
rect 75048 64993 75181 64998
rect 75606 65055 75853 65060
rect 74222 64971 74470 64976
rect 75606 64980 75616 65055
rect 75843 64980 75853 65055
rect 76411 64998 76421 65111
rect 76534 64998 76544 65111
rect 77760 65112 77893 65117
rect 76411 64993 76544 64998
rect 76987 65054 77235 65059
rect 75606 64975 75853 64980
rect 76987 64982 76997 65054
rect 77225 64982 77235 65054
rect 77760 64999 77770 65112
rect 77883 64999 77893 65112
rect 77760 64994 77893 64999
rect 76987 64977 77235 64982
rect 61519 64144 61647 64149
rect 61519 64134 61524 64144
rect 60693 64026 61524 64134
rect 61642 64134 61647 64144
rect 71632 64136 71760 64141
rect 71632 64134 71637 64136
rect 61642 64026 71637 64134
rect 60693 64018 71637 64026
rect 71755 64134 71760 64136
rect 113316 64134 113434 70709
rect 71755 64129 113434 64134
rect 71755 64021 84180 64129
rect 84288 64021 101834 64129
rect 101942 64021 113434 64129
rect 71755 64018 113434 64021
rect 60693 64016 113434 64018
rect 71632 64013 71760 64016
rect 86475 63858 86639 63863
rect 85118 63849 85328 63854
rect 85118 63757 85128 63849
rect 85318 63757 85328 63849
rect 85118 63752 85328 63757
rect 85558 63823 86012 63828
rect 85558 63736 85568 63823
rect 86002 63736 86012 63823
rect 86475 63764 86485 63858
rect 86629 63764 86639 63858
rect 104129 63858 104293 63863
rect 102772 63849 102982 63854
rect 86475 63759 86639 63764
rect 86894 63809 87338 63814
rect 85558 63731 86012 63736
rect 86894 63732 86904 63809
rect 87328 63732 87338 63809
rect 102772 63757 102782 63849
rect 102972 63757 102982 63849
rect 102772 63752 102982 63757
rect 103212 63823 103666 63828
rect 86894 63727 87338 63732
rect 103212 63736 103222 63823
rect 103656 63736 103666 63823
rect 104129 63764 104139 63858
rect 104283 63764 104293 63858
rect 104129 63759 104293 63764
rect 104548 63809 104992 63814
rect 103212 63731 103666 63736
rect 104548 63732 104558 63809
rect 104982 63732 104992 63809
rect 104548 63727 104992 63732
rect 62124 63540 62252 63545
rect 62124 63534 62129 63540
rect 60693 63422 62129 63534
rect 62247 63534 62252 63540
rect 72117 63539 72245 63544
rect 72117 63534 72122 63539
rect 62247 63422 72122 63534
rect 60693 63421 72122 63422
rect 72240 63534 72245 63539
rect 115325 63534 115443 70709
rect 72240 63421 115443 63534
rect 60693 63416 115443 63421
rect 117343 62934 117461 70709
rect 60693 62929 117461 62934
rect 60693 62821 60901 62929
rect 61009 62821 71110 62929
rect 71218 62821 88038 62929
rect 88146 62821 105692 62929
rect 105800 62821 117461 62929
rect 60693 62816 117461 62821
rect 85209 62346 85321 62351
rect 102863 62346 102975 62351
rect 85209 62237 85219 62346
rect 85311 62237 85321 62346
rect 85209 62232 85321 62237
rect 86540 62341 86652 62346
rect 86540 62232 86550 62341
rect 86642 62232 86652 62341
rect 102863 62237 102873 62346
rect 102965 62237 102975 62346
rect 102863 62232 102975 62237
rect 104194 62341 104306 62346
rect 104194 62232 104204 62341
rect 104296 62232 104306 62341
rect 86540 62227 86652 62232
rect 104194 62227 104306 62232
rect 62721 62189 62854 62194
rect 62721 62076 62731 62189
rect 62844 62076 62854 62189
rect 72721 62189 72854 62194
rect 64711 62177 64844 62182
rect 64368 62159 64501 62164
rect 62721 62071 62854 62076
rect 63419 62146 63552 62151
rect 63419 62033 63429 62146
rect 63542 62033 63552 62146
rect 64368 62045 64378 62159
rect 64491 62045 64501 62159
rect 64711 62064 64721 62177
rect 64834 62064 64844 62177
rect 64711 62059 64844 62064
rect 65446 62169 65579 62174
rect 65446 62056 65456 62169
rect 65569 62056 65579 62169
rect 65446 62051 65579 62056
rect 66165 62151 66298 62156
rect 64368 62040 64501 62045
rect 66165 62038 66175 62151
rect 66288 62038 66298 62151
rect 67533 62151 67666 62156
rect 66165 62033 66298 62038
rect 66818 62143 66951 62148
rect 63419 62028 63552 62033
rect 66818 62030 66828 62143
rect 66941 62030 66951 62143
rect 67533 62038 67543 62151
rect 67656 62038 67666 62151
rect 72721 62076 72731 62189
rect 72844 62076 72854 62189
rect 74711 62177 74844 62182
rect 74368 62159 74501 62164
rect 72721 62071 72854 62076
rect 73419 62146 73552 62151
rect 67533 62033 67666 62038
rect 73419 62033 73429 62146
rect 73542 62033 73552 62146
rect 74368 62045 74378 62159
rect 74491 62045 74501 62159
rect 74711 62064 74721 62177
rect 74834 62064 74844 62177
rect 74711 62059 74844 62064
rect 75446 62169 75579 62174
rect 75446 62056 75456 62169
rect 75569 62056 75579 62169
rect 75446 62051 75579 62056
rect 76165 62151 76298 62156
rect 74368 62040 74501 62045
rect 76165 62038 76175 62151
rect 76288 62038 76298 62151
rect 77533 62151 77666 62156
rect 76165 62033 76298 62038
rect 76818 62143 76951 62148
rect 66818 62025 66951 62030
rect 73419 62028 73552 62033
rect 76818 62030 76828 62143
rect 76941 62030 76951 62143
rect 77533 62038 77543 62151
rect 77656 62038 77666 62151
rect 77533 62033 77666 62038
rect 76818 62025 76951 62030
rect 65874 61473 65962 61478
rect 63153 61352 63244 61357
rect 63153 61245 63163 61352
rect 63234 61245 63244 61352
rect 63153 61240 63244 61245
rect 63695 61346 63786 61351
rect 63695 61242 63705 61346
rect 63776 61242 63786 61346
rect 65874 61349 65884 61473
rect 65952 61349 65962 61473
rect 75874 61473 75962 61478
rect 66961 61383 67053 61388
rect 65874 61344 65962 61349
rect 66416 61364 66504 61369
rect 63695 61237 63786 61242
rect 64241 61330 64330 61335
rect 64241 61184 64251 61330
rect 64320 61184 64330 61330
rect 64788 61321 64872 61326
rect 64788 61191 64798 61321
rect 64862 61191 64872 61321
rect 66416 61207 66426 61364
rect 66494 61207 66504 61364
rect 66961 61261 66971 61383
rect 67043 61261 67053 61383
rect 66961 61256 67053 61261
rect 67504 61356 67590 61361
rect 66416 61202 66504 61207
rect 67504 61202 67514 61356
rect 67580 61202 67590 61356
rect 73153 61352 73244 61357
rect 73153 61245 73163 61352
rect 73234 61245 73244 61352
rect 73153 61240 73244 61245
rect 73695 61346 73786 61351
rect 73695 61242 73705 61346
rect 73776 61242 73786 61346
rect 75874 61349 75884 61473
rect 75952 61349 75962 61473
rect 76961 61383 77053 61388
rect 75874 61344 75962 61349
rect 76416 61364 76504 61369
rect 73695 61237 73786 61242
rect 74241 61330 74330 61335
rect 67504 61197 67590 61202
rect 64788 61186 64872 61191
rect 64241 61179 64330 61184
rect 74241 61184 74251 61330
rect 74320 61184 74330 61330
rect 74788 61321 74872 61326
rect 74788 61191 74798 61321
rect 74862 61191 74872 61321
rect 76416 61207 76426 61364
rect 76494 61207 76504 61364
rect 76961 61261 76971 61383
rect 77043 61261 77053 61383
rect 76961 61256 77053 61261
rect 77504 61356 77590 61361
rect 76416 61202 76504 61207
rect 77504 61202 77514 61356
rect 77580 61202 77590 61356
rect 77504 61197 77590 61202
rect 74788 61186 74872 61191
rect 74241 61179 74330 61184
rect 65333 61015 65420 61020
rect 65333 60862 65343 61015
rect 65410 60862 65420 61015
rect 65333 60857 65420 60862
rect 75333 61015 75420 61020
rect 75333 60862 75343 61015
rect 75410 60862 75420 61015
rect 75333 60857 75420 60862
rect 86084 60499 86169 60504
rect 86084 60357 86094 60499
rect 86159 60357 86169 60499
rect 86084 60352 86169 60357
rect 103738 60499 103823 60504
rect 103738 60357 103748 60499
rect 103813 60357 103823 60499
rect 103738 60352 103823 60357
rect 86626 60280 86714 60285
rect 85534 60274 85625 60279
rect 85534 60170 85544 60274
rect 85615 60170 85625 60274
rect 85534 60165 85625 60170
rect 86626 60170 86636 60280
rect 86704 60170 86714 60280
rect 104280 60280 104368 60285
rect 86626 60165 86714 60170
rect 103188 60274 103279 60279
rect 103188 60170 103198 60274
rect 103269 60170 103279 60274
rect 103188 60165 103279 60170
rect 104280 60170 104290 60280
rect 104358 60170 104368 60280
rect 104280 60165 104368 60170
rect 64362 60000 64690 60005
rect 63042 59993 63315 59998
rect 63042 59916 63052 59993
rect 63305 59916 63315 59993
rect 63042 59911 63315 59916
rect 64362 59915 64372 60000
rect 64680 59915 64690 60000
rect 74362 60000 74690 60005
rect 64362 59910 64690 59915
rect 65750 59989 66052 59994
rect 65750 59918 65760 59989
rect 66042 59918 66052 59989
rect 65750 59913 66052 59918
rect 67122 59991 67424 59996
rect 67122 59920 67132 59991
rect 67414 59920 67424 59991
rect 67122 59915 67424 59920
rect 73042 59993 73315 59998
rect 73042 59916 73052 59993
rect 73305 59916 73315 59993
rect 73042 59911 73315 59916
rect 74362 59915 74372 60000
rect 74680 59915 74690 60000
rect 74362 59910 74690 59915
rect 75750 59989 76052 59994
rect 75750 59918 75760 59989
rect 76042 59918 76052 59989
rect 75750 59913 76052 59918
rect 77122 59991 77424 59996
rect 77122 59920 77132 59991
rect 77414 59920 77424 59991
rect 77122 59915 77424 59920
rect 84933 59636 85066 59641
rect 84933 59523 84943 59636
rect 85056 59523 85066 59636
rect 84933 59518 85066 59523
rect 102587 59636 102720 59641
rect 102587 59523 102597 59636
rect 102710 59523 102720 59636
rect 102587 59518 102720 59523
rect 68034 59416 68167 59421
rect 66650 59381 66783 59386
rect 65288 59363 65421 59368
rect 63927 59351 64060 59356
rect 63927 59238 63937 59351
rect 64050 59238 64060 59351
rect 65288 59250 65298 59363
rect 65411 59250 65421 59363
rect 66650 59268 66660 59381
rect 66773 59268 66783 59381
rect 68034 59303 68044 59416
rect 68157 59303 68167 59416
rect 78034 59416 78167 59421
rect 76650 59381 76783 59386
rect 75288 59363 75421 59368
rect 68034 59298 68167 59303
rect 73927 59351 74060 59356
rect 66650 59263 66783 59268
rect 65288 59245 65421 59250
rect 63927 59233 64060 59238
rect 73927 59238 73937 59351
rect 74050 59238 74060 59351
rect 75288 59250 75298 59363
rect 75411 59250 75421 59363
rect 76650 59268 76660 59381
rect 76773 59268 76783 59381
rect 78034 59303 78044 59416
rect 78157 59303 78167 59416
rect 78034 59298 78167 59303
rect 76650 59263 76783 59268
rect 75288 59245 75421 59250
rect 73927 59233 74060 59238
rect 87326 59030 87459 59035
rect 87326 58917 87336 59030
rect 87449 58917 87459 59030
rect 87326 58912 87459 58917
rect 104980 59030 105113 59035
rect 104980 58917 104990 59030
rect 105103 58917 105113 59030
rect 104980 58912 105113 58917
rect 62496 54768 62623 54773
rect 62496 54651 62501 54768
rect 62618 54763 74838 54768
rect 62618 54656 74726 54763
rect 74833 54656 74838 54763
rect 62618 54651 74838 54656
rect 62496 54646 62623 54651
rect 27435 52669 27561 52674
rect 27434 52668 48568 52669
rect 27434 52542 27435 52668
rect 27561 52636 48568 52668
rect 27561 52576 46449 52636
rect 46509 52633 48568 52636
rect 46509 52576 48449 52633
rect 27561 52573 48449 52576
rect 48509 52573 48568 52633
rect 27561 52542 48568 52573
rect 27434 52541 48568 52542
rect 27435 52536 27561 52541
rect 116728 52514 116876 52519
rect 116728 52386 116738 52514
rect 116866 52386 116876 52514
rect 116728 52381 116876 52386
rect 120652 52467 120943 52472
rect 120652 52363 120662 52467
rect 120933 52363 120943 52467
rect 120652 52358 120943 52363
rect 46143 52282 46281 52287
rect 46143 51695 46153 52282
rect 46271 51695 46281 52282
rect 48187 52230 48317 52235
rect 46143 51690 46281 51695
rect 47483 51852 47618 51857
rect 47483 51229 47493 51852
rect 47608 51229 47618 51852
rect 48187 51690 48197 52230
rect 48307 51690 48317 52230
rect 63312 52174 65303 52179
rect 58759 52159 58825 52164
rect 58759 52103 58764 52159
rect 58820 52103 58825 52159
rect 58759 52098 58825 52103
rect 48187 51685 48317 51690
rect 49501 51907 49664 51912
rect 49501 51249 49511 51907
rect 49654 51249 49664 51907
rect 49501 51244 49664 51249
rect 47483 51224 47618 51229
rect 45802 50922 49364 50923
rect 45797 50796 45803 50922
rect 45929 50892 49364 50922
rect 45929 50822 47273 50892
rect 47343 50890 49364 50892
rect 47343 50830 49271 50890
rect 49331 50830 49364 50890
rect 47343 50822 49364 50830
rect 45929 50796 49364 50822
rect 45802 50795 49364 50796
rect 24762 50635 24888 50640
rect 24761 50634 38505 50635
rect 24761 50508 24762 50634
rect 24888 50595 38505 50634
rect 24888 50593 38404 50595
rect 24888 50533 36406 50593
rect 36466 50535 38404 50593
rect 38464 50535 38505 50595
rect 36466 50533 38505 50535
rect 24888 50508 38505 50533
rect 24761 50507 38505 50508
rect 24762 50502 24888 50507
rect 39483 50313 39618 50318
rect 37437 50285 37577 50290
rect 36192 49927 36295 49932
rect 36192 49483 36202 49927
rect 36285 49483 36295 49927
rect 37437 49792 37447 50285
rect 37567 49792 37577 50285
rect 37437 49787 37577 49792
rect 38134 49857 38253 49862
rect 36192 49478 36295 49483
rect 38134 49278 38144 49857
rect 38243 49278 38253 49857
rect 39483 49780 39493 50313
rect 39608 49780 39618 50313
rect 39483 49775 39618 49780
rect 38134 49273 38253 49278
rect 25662 49058 25788 49063
rect 25661 49057 39319 49058
rect 25661 48931 25662 49057
rect 25788 49027 39319 49057
rect 25788 48967 37227 49027
rect 37287 49016 39319 49027
rect 37287 48967 39227 49016
rect 25788 48956 39227 48967
rect 39287 48956 39319 49016
rect 25788 48931 39319 48956
rect 25661 48930 39319 48931
rect 25662 48925 25788 48930
rect 26624 48330 26750 48335
rect 45802 48330 45930 48336
rect 26623 48329 45802 48330
rect 26623 48203 26624 48329
rect 26750 48203 45802 48329
rect 26623 48202 45802 48203
rect 26624 48197 26750 48202
rect 45802 48196 45930 48202
rect 56036 47379 56340 47384
rect 56036 46741 56046 47379
rect 56330 46741 56340 47379
rect 56036 46736 56340 46741
rect 58762 45847 58822 52098
rect 63312 51978 63317 52174
rect 63513 51978 65303 52174
rect 63312 51973 65303 51978
rect 119316 52130 119417 52135
rect 117719 51778 117842 51783
rect 115279 51725 115395 51730
rect 64046 51678 66239 51683
rect 62501 51663 62618 51668
rect 61618 51650 61749 51655
rect 61618 51529 61623 51650
rect 61744 51529 61749 51650
rect 61618 50392 61749 51529
rect 62501 51556 62506 51663
rect 62613 51556 62618 51663
rect 61613 50387 61754 50392
rect 61613 50256 61618 50387
rect 61749 50256 61754 50387
rect 61613 50251 61754 50256
rect 60482 47309 61506 47314
rect 60482 47109 60492 47309
rect 61496 47109 61506 47309
rect 62501 47279 62618 51556
rect 64046 51482 66038 51678
rect 66234 51482 66239 51678
rect 64046 51477 66239 51482
rect 62838 49622 63390 49627
rect 62838 49465 62848 49622
rect 63380 49465 63390 49622
rect 62838 49460 63390 49465
rect 62496 47274 62623 47279
rect 62496 47157 62501 47274
rect 62618 47157 62623 47274
rect 62496 47152 62623 47157
rect 60482 47104 61506 47109
rect 58757 45842 58827 45847
rect 58757 45782 58762 45842
rect 58822 45782 58827 45842
rect 58757 45777 58827 45782
rect 62000 42674 62290 42679
rect 33473 41686 38293 41750
rect 43345 41677 44585 41741
rect 46545 41602 47958 41666
rect 62000 41599 62010 42674
rect 62280 41599 62290 42674
rect 33296 33165 33360 41532
rect 36678 40610 36834 40618
rect 36678 40472 36688 40610
rect 36826 40472 36834 40610
rect 36678 40464 36834 40472
rect 38633 39854 38697 41321
rect 42833 39888 42897 41299
rect 44947 40533 45108 40541
rect 44947 40395 44960 40533
rect 45098 40395 45108 40533
rect 44947 40385 45108 40395
rect 42833 39435 42897 39768
rect 44984 39435 45048 39788
rect 48170 39435 48234 41599
rect 62000 41594 62290 41599
rect 62847 42671 63137 42676
rect 62847 41596 62857 42671
rect 63127 41596 63137 42671
rect 63402 42335 63627 42340
rect 63402 41747 63412 42335
rect 63617 41747 63627 42335
rect 63402 41742 63627 41747
rect 62847 41591 63137 41596
rect 56017 39355 56177 39360
rect 36482 36391 36546 38338
rect 38633 36662 38697 38130
rect 42833 35486 42897 38966
rect 44984 36102 45048 38966
rect 35195 34277 35323 34855
rect 35195 34159 35200 34277
rect 35318 34159 35323 34277
rect 35195 34154 35323 34159
rect 38633 33303 38697 34983
rect 42833 33443 42897 34962
rect 44800 34263 44918 34842
rect 44800 34155 44805 34263
rect 44913 34155 44918 34263
rect 44800 34143 44918 34155
rect 48170 33232 48234 38966
rect 56017 38731 56027 39355
rect 56167 38731 56177 39355
rect 56017 38726 56177 38731
rect 33572 33098 34985 33162
rect 36945 33023 38185 33087
rect 43237 33014 48057 33078
rect 50233 32667 50243 32672
rect 40656 32643 40666 32648
rect 40656 32525 40661 32643
rect 40656 32520 40666 32525
rect 40784 32520 40790 32648
rect 50233 32549 50238 32667
rect 50233 32544 50243 32549
rect 50361 32544 50367 32672
rect 36513 31150 36631 31797
rect 36508 31145 36636 31150
rect 36508 31027 36513 31145
rect 36631 31027 36636 31145
rect 42143 31071 42261 31802
rect 55942 31354 56309 31359
rect 36508 31022 36636 31027
rect 42138 31066 42266 31071
rect 42138 30948 42143 31066
rect 42261 30948 42266 31066
rect 42138 30943 42266 30948
rect 55942 30754 55952 31354
rect 56299 30754 56309 31354
rect 55942 30749 56309 30754
rect 60976 30188 61201 30193
rect 60976 29648 60986 30188
rect 61191 29648 61201 30188
rect 60976 29643 61201 29648
rect 64046 29335 64252 51477
rect 115279 51273 115289 51725
rect 115385 51273 115395 51725
rect 117719 51316 117729 51778
rect 117832 51316 117842 51778
rect 117719 51311 117842 51316
rect 115279 51268 115395 51273
rect 119316 51001 119326 52130
rect 119407 51001 119417 52130
rect 121699 52123 121814 52128
rect 121699 51027 121709 52123
rect 121804 51027 121814 52123
rect 121699 51022 121814 51027
rect 119316 50996 119417 51001
rect 121186 50958 121526 50963
rect 117386 50953 117563 50958
rect 115569 50928 115717 50933
rect 115569 50800 115579 50928
rect 115707 50800 115717 50928
rect 117386 50869 117396 50953
rect 117553 50869 117563 50953
rect 115569 50795 115717 50800
rect 115979 50861 116151 50866
rect 117386 50864 117563 50869
rect 119926 50944 120235 50949
rect 115979 50709 115989 50861
rect 116141 50709 116151 50861
rect 119926 50772 119936 50944
rect 120225 50772 120235 50944
rect 121186 50888 121196 50958
rect 121516 50888 121526 50958
rect 121186 50883 121526 50888
rect 119926 50767 120235 50772
rect 115979 50704 116151 50709
rect 102484 50225 102732 50230
rect 67960 50219 68208 50224
rect 66164 50207 66372 50212
rect 66164 50013 66174 50207
rect 66362 50013 66372 50207
rect 66164 50008 66372 50013
rect 67960 49987 67970 50219
rect 68198 49987 68208 50219
rect 71473 50211 71721 50216
rect 100688 50213 100896 50218
rect 67960 49982 68208 49987
rect 69654 50200 69902 50205
rect 69654 49968 69664 50200
rect 69892 49968 69902 50200
rect 71473 49979 71483 50211
rect 71711 49979 71721 50211
rect 71473 49974 71721 49979
rect 73257 50208 73505 50213
rect 73257 49976 73267 50208
rect 73495 49976 73505 50208
rect 73257 49971 73505 49976
rect 75042 50206 75290 50211
rect 75042 49974 75052 50206
rect 75280 49974 75290 50206
rect 100688 50019 100698 50213
rect 100886 50019 100896 50213
rect 100688 50014 100896 50019
rect 102484 49993 102494 50225
rect 102722 49993 102732 50225
rect 105997 50217 106245 50222
rect 102484 49988 102732 49993
rect 104178 50206 104426 50211
rect 75042 49969 75290 49974
rect 104178 49974 104188 50206
rect 104416 49974 104426 50206
rect 105997 49985 106007 50217
rect 106235 49985 106245 50217
rect 105997 49980 106245 49985
rect 107781 50214 108029 50219
rect 107781 49982 107791 50214
rect 108019 49982 108029 50214
rect 107781 49977 108029 49982
rect 109566 50212 109814 50217
rect 109566 49980 109576 50212
rect 109804 49980 109814 50212
rect 109566 49975 109814 49980
rect 104178 49969 104426 49974
rect 69654 49963 69902 49968
rect 96354 49834 97884 49839
rect 96354 49432 96364 49834
rect 97874 49432 97884 49834
rect 96354 49427 97884 49432
rect 101668 48668 101924 48673
rect 67144 48662 67400 48667
rect 65274 48632 65570 48637
rect 65274 48532 65284 48632
rect 65560 48532 65570 48632
rect 67144 48584 67154 48662
rect 67390 48584 67400 48662
rect 67144 48579 67400 48584
rect 68949 48655 69203 48660
rect 68949 48576 68959 48655
rect 69193 48576 69203 48655
rect 68949 48571 69203 48576
rect 70755 48651 70994 48656
rect 70755 48570 70765 48651
rect 70984 48570 70994 48651
rect 70755 48565 70994 48570
rect 72541 48655 72801 48660
rect 72541 48571 72551 48655
rect 72791 48571 72801 48655
rect 74342 48651 74614 48656
rect 74342 48586 74352 48651
rect 74604 48586 74614 48651
rect 74342 48581 74614 48586
rect 99798 48638 100094 48643
rect 72541 48566 72801 48571
rect 99798 48538 99808 48638
rect 100084 48538 100094 48638
rect 101668 48590 101678 48668
rect 101914 48590 101924 48668
rect 101668 48585 101924 48590
rect 103473 48661 103727 48666
rect 103473 48582 103483 48661
rect 103717 48582 103727 48661
rect 103473 48577 103727 48582
rect 105279 48657 105518 48662
rect 105279 48576 105289 48657
rect 105508 48576 105518 48657
rect 105279 48571 105518 48576
rect 107065 48661 107325 48666
rect 107065 48577 107075 48661
rect 107315 48577 107325 48661
rect 108866 48657 109138 48662
rect 108866 48592 108876 48657
rect 109128 48592 109138 48657
rect 108866 48587 109138 48592
rect 107065 48572 107325 48577
rect 99798 48533 100094 48538
rect 65274 48527 65570 48532
rect 90786 47320 91118 47325
rect 90786 46782 90796 47320
rect 91108 46782 91118 47320
rect 94977 47300 96104 47305
rect 94977 47083 94987 47300
rect 96094 47083 96104 47300
rect 94977 47078 96104 47083
rect 90786 46777 91118 46782
rect 89567 43280 89693 43285
rect 85545 43279 89694 43280
rect 85545 43237 89567 43279
rect 85545 43173 85593 43237
rect 85657 43173 87594 43237
rect 87658 43173 89567 43237
rect 85545 43153 89567 43173
rect 89693 43153 89694 43279
rect 85545 43152 89694 43153
rect 89567 43147 89693 43152
rect 96515 42681 96805 42686
rect 86519 42646 86628 42651
rect 84495 42609 84638 42614
rect 84495 42267 84505 42609
rect 84628 42267 84638 42609
rect 84495 42262 84638 42267
rect 86519 42262 86529 42646
rect 86618 42262 86628 42646
rect 86519 42257 86628 42262
rect 84739 41756 88642 41757
rect 84739 41731 88515 41756
rect 84739 41728 86765 41731
rect 84739 41664 84767 41728
rect 84831 41667 86765 41728
rect 86829 41667 88515 41731
rect 84831 41664 88515 41667
rect 84739 41630 88515 41664
rect 88641 41630 88647 41756
rect 84739 41629 88642 41630
rect 96515 41606 96525 42681
rect 96795 41606 96805 42681
rect 96515 41601 96805 41606
rect 97362 42678 97652 42683
rect 97362 41603 97372 42678
rect 97642 41603 97652 42678
rect 97962 42396 98228 42401
rect 97962 41682 97972 42396
rect 98218 41682 98228 42396
rect 97962 41677 98228 41682
rect 97362 41598 97652 41603
rect 78108 41469 83095 41470
rect 78103 41343 78109 41469
rect 78235 41440 83095 41469
rect 78235 41431 83000 41440
rect 78235 41367 81000 41431
rect 81064 41376 83000 41431
rect 83064 41376 83095 41440
rect 81064 41367 83095 41376
rect 78235 41343 83095 41367
rect 78108 41342 83095 41343
rect 85864 41241 86138 41252
rect 85864 41005 85883 41241
rect 86119 41005 86138 41241
rect 85864 40988 86138 41005
rect 87796 41223 88032 41236
rect 87796 41012 87808 41223
rect 88019 41012 88032 41223
rect 87796 41000 88032 41012
rect 79894 40739 79993 40744
rect 79894 40461 79904 40739
rect 79983 40461 79993 40739
rect 79894 40456 79993 40461
rect 81955 40703 82055 40708
rect 81955 40420 81965 40703
rect 82045 40420 82055 40703
rect 81955 40415 82055 40420
rect 79094 39950 79220 39955
rect 79093 39949 82288 39950
rect 79093 39823 79094 39949
rect 79220 39923 82288 39949
rect 79220 39921 82166 39923
rect 79220 39857 80175 39921
rect 80239 39857 82166 39921
rect 79220 39849 82166 39857
rect 82240 39849 82288 39923
rect 79220 39823 82288 39849
rect 79093 39822 82288 39823
rect 79094 39817 79220 39822
rect 83008 39719 83152 39724
rect 81151 39704 81299 39719
rect 81151 39576 81162 39704
rect 81290 39576 81299 39704
rect 83008 39595 83018 39719
rect 83142 39595 83152 39719
rect 83008 39590 83152 39595
rect 81151 39557 81299 39576
rect 114699 39378 115018 39383
rect 90773 38958 91040 38963
rect 90773 38091 90783 38958
rect 91030 38091 91040 38958
rect 114699 38737 114709 39378
rect 115008 38737 115018 39378
rect 114699 38732 115018 38737
rect 90773 38086 91040 38091
rect 123001 38345 123105 38350
rect 68823 37306 69087 37311
rect 66920 37246 67184 37251
rect 65318 37235 65582 37240
rect 65318 37035 65328 37235
rect 65572 37035 65582 37235
rect 66920 37046 66930 37246
rect 67174 37046 67184 37246
rect 68823 37106 68833 37306
rect 69077 37106 69087 37306
rect 103339 37299 103603 37304
rect 68823 37101 69087 37106
rect 70540 37290 70804 37295
rect 70540 37090 70550 37290
rect 70794 37090 70804 37290
rect 70540 37085 70804 37090
rect 72354 37285 72618 37290
rect 72354 37085 72364 37285
rect 72608 37085 72618 37285
rect 72354 37080 72618 37085
rect 74326 37279 74590 37284
rect 74326 37079 74336 37279
rect 74580 37079 74590 37279
rect 101436 37239 101700 37244
rect 74326 37074 74590 37079
rect 99834 37228 100098 37233
rect 66920 37041 67184 37046
rect 65318 37030 65582 37035
rect 99834 37028 99844 37228
rect 100088 37028 100098 37228
rect 101436 37039 101446 37239
rect 101690 37039 101700 37239
rect 103339 37099 103349 37299
rect 103593 37099 103603 37299
rect 103339 37094 103603 37099
rect 105056 37283 105320 37288
rect 105056 37083 105066 37283
rect 105310 37083 105320 37283
rect 105056 37078 105320 37083
rect 106870 37278 107134 37283
rect 106870 37078 106880 37278
rect 107124 37078 107134 37278
rect 106870 37073 107134 37078
rect 108842 37272 109106 37277
rect 108842 37072 108852 37272
rect 109096 37072 109106 37272
rect 108842 37067 109106 37072
rect 123001 37052 123011 38345
rect 123095 37052 123105 38345
rect 123001 37047 123105 37052
rect 101436 37034 101700 37039
rect 99834 37023 100098 37028
rect 123001 36885 123105 36890
rect 96839 35851 97606 35856
rect 67631 35741 68051 35746
rect 65840 35734 66244 35739
rect 65840 35656 65850 35734
rect 66234 35656 66244 35734
rect 67631 35667 67641 35741
rect 68041 35667 68051 35741
rect 67631 35662 68051 35667
rect 69437 35741 69845 35746
rect 69437 35667 69447 35741
rect 69835 35667 69845 35741
rect 96839 35740 96849 35851
rect 97596 35740 97606 35851
rect 96839 35735 97606 35740
rect 102147 35734 102567 35739
rect 100356 35727 100760 35732
rect 69437 35662 69845 35667
rect 71234 35706 71642 35711
rect 65840 35651 66244 35656
rect 71234 35632 71244 35706
rect 71632 35632 71642 35706
rect 71234 35627 71642 35632
rect 73036 35706 73443 35711
rect 73036 35628 73046 35706
rect 73433 35628 73443 35706
rect 73036 35623 73443 35628
rect 74830 35702 75245 35707
rect 74830 35625 74840 35702
rect 75235 35625 75245 35702
rect 74830 35620 75245 35625
rect 67550 35060 67668 35065
rect 67550 34952 67555 35060
rect 67663 34952 67668 35060
rect 67550 33440 67668 34952
rect 82555 34935 82619 35541
rect 83771 34895 83928 34908
rect 83771 34757 83780 34895
rect 83918 34757 83928 34895
rect 85567 34894 85631 35655
rect 100356 35649 100366 35727
rect 100750 35649 100760 35727
rect 102147 35660 102157 35734
rect 102557 35660 102567 35734
rect 102147 35655 102567 35660
rect 103953 35734 104361 35739
rect 103953 35660 103963 35734
rect 104351 35660 104361 35734
rect 103953 35655 104361 35660
rect 105750 35699 106158 35704
rect 100356 35644 100760 35649
rect 105750 35625 105760 35699
rect 106148 35625 106158 35699
rect 105750 35620 106158 35625
rect 107552 35699 107959 35704
rect 107552 35621 107562 35699
rect 107949 35621 107959 35699
rect 107552 35616 107959 35621
rect 109346 35695 109761 35700
rect 109346 35618 109356 35695
rect 109751 35618 109761 35695
rect 109346 35613 109761 35618
rect 123001 35592 123011 36885
rect 123095 35592 123105 36885
rect 123001 35587 123105 35592
rect 91354 35537 91558 35542
rect 89487 35536 91559 35537
rect 89487 35532 91354 35536
rect 86360 35330 86514 35338
rect 89487 35336 89492 35532
rect 89688 35336 91354 35532
rect 89487 35332 91354 35336
rect 91558 35332 91559 35536
rect 89487 35331 91559 35332
rect 94542 35536 94746 35542
rect 86360 35192 86368 35330
rect 86506 35192 86514 35330
rect 91354 35326 91558 35331
rect 94542 35326 94746 35332
rect 123002 35405 123105 35410
rect 86360 35183 86514 35192
rect 83771 34736 83928 34757
rect 81528 34563 83251 34627
rect 67532 33421 67681 33440
rect 67532 33303 67550 33421
rect 67668 33303 67681 33421
rect 67532 33291 67681 33303
rect 81512 30938 81576 34535
rect 82675 33515 82741 33520
rect 82675 33459 82680 33515
rect 82736 33459 82741 33515
rect 82675 33454 82741 33459
rect 82305 33160 82443 33165
rect 82305 33032 82310 33160
rect 82438 33032 82443 33160
rect 82305 33027 82443 33032
rect 82671 32063 82745 32068
rect 82671 31999 82676 32063
rect 82740 31999 82745 32063
rect 82671 31994 82745 31999
rect 81959 31877 82087 31882
rect 81959 31759 81964 31877
rect 82082 31759 82087 31877
rect 81959 31754 82087 31759
rect 82222 31334 82358 31343
rect 82222 31218 82232 31334
rect 82348 31218 82358 31334
rect 82222 31211 82358 31218
rect 83187 30938 83251 34563
rect 84505 34572 86244 34636
rect 83646 33792 83774 33797
rect 83646 33674 83651 33792
rect 83769 33674 83774 33792
rect 83646 33669 83774 33674
rect 81512 30874 83251 30938
rect 84505 30947 84569 34572
rect 85006 33512 85072 33517
rect 85006 33456 85011 33512
rect 85067 33456 85072 33512
rect 85006 33451 85072 33456
rect 85316 33167 85454 33172
rect 85316 33039 85321 33167
rect 85449 33039 85454 33167
rect 85316 33034 85454 33039
rect 85787 31835 85919 31850
rect 84966 31814 85094 31819
rect 84966 31696 84971 31814
rect 85089 31696 85094 31814
rect 85787 31719 85795 31835
rect 85911 31719 85919 31835
rect 85787 31709 85919 31719
rect 84966 31691 85094 31696
rect 86180 30975 86244 34572
rect 91312 34384 91516 34389
rect 95265 34384 95470 34389
rect 123002 34387 123012 35405
rect 123095 34387 123105 35405
rect 88556 34383 91517 34384
rect 88556 34379 91312 34383
rect 88556 34183 88561 34379
rect 88757 34183 91312 34379
rect 88556 34179 91312 34183
rect 91516 34179 91517 34383
rect 88556 34178 91517 34179
rect 95265 34383 95471 34384
rect 95470 34179 95471 34383
rect 123002 34382 123105 34387
rect 128026 34927 166970 34932
rect 95265 34178 95471 34179
rect 91312 34173 91516 34178
rect 95265 34173 95470 34178
rect 125018 34131 125358 34136
rect 119407 33914 119413 34040
rect 119539 33914 119545 34040
rect 125018 33811 125028 34131
rect 125348 33811 125358 34131
rect 128026 33937 128031 34927
rect 129021 33937 166970 34927
rect 128026 33932 166970 33937
rect 125018 33806 125358 33811
rect 127207 33739 127604 33744
rect 127207 33666 127217 33739
rect 127594 33666 127604 33739
rect 127207 33661 127604 33666
rect 123000 33617 123107 33622
rect 123000 32643 123010 33617
rect 123097 32643 123107 33617
rect 123000 32638 123107 32643
rect 127209 32617 127601 32622
rect 127209 32552 127219 32617
rect 127591 32552 127601 32617
rect 127209 32547 127601 32552
rect 122997 32470 123107 32475
rect 86661 31819 86789 31824
rect 86661 31701 86666 31819
rect 86784 31701 86789 31819
rect 86661 31696 86789 31701
rect 114706 31367 115025 31372
rect 95417 31246 95721 31251
rect 84505 30883 86228 30947
rect 95417 30789 95427 31246
rect 95711 30789 95721 31246
rect 95417 30784 95721 30789
rect 90804 30752 91066 30757
rect 82529 30047 82593 30470
rect 85524 29897 85588 30658
rect 90804 30288 90814 30752
rect 91056 30288 91066 30752
rect 114706 30726 114716 31367
rect 115015 30726 115025 31367
rect 122997 31104 123007 32470
rect 123097 31104 123107 32470
rect 122997 31099 123107 31104
rect 124319 31186 124659 31191
rect 114706 30721 115025 30726
rect 122998 30864 123109 30869
rect 90804 30283 91066 30288
rect 122998 29606 123008 30864
rect 123099 29606 123109 30864
rect 124319 30866 124329 31186
rect 124649 30866 124659 31186
rect 124319 30861 124659 30866
rect 122998 29601 123109 29606
rect 64041 29330 64257 29335
rect 64041 29124 64046 29330
rect 64252 29124 64257 29330
rect 64041 29119 64257 29124
rect 58866 27670 59072 28849
rect 59353 28687 61043 28692
rect 59353 28460 59363 28687
rect 61033 28460 61043 28687
rect 59353 28455 61043 28460
rect 45485 27628 59072 27670
rect 45485 27510 45534 27628
rect 45652 27510 59072 27628
rect 45485 27464 59072 27510
rect 93382 27680 93588 28779
rect 95193 28684 95772 28689
rect 95193 28464 95203 28684
rect 95762 28464 95772 28684
rect 95193 28459 95772 28464
rect 93382 27474 94041 27680
rect 93835 27016 94041 27474
rect 104374 27177 104528 27194
rect 104374 27049 104388 27177
rect 104516 27049 104528 27177
rect 107951 27185 107961 27190
rect 107951 27067 107956 27185
rect 107951 27062 107961 27067
rect 108079 27062 108085 27190
rect 104374 27041 104528 27049
rect 93835 26820 93840 27016
rect 94036 26820 94041 27016
rect 93835 26815 94041 26820
rect 86367 24988 86505 24993
rect 86367 24870 86377 24988
rect 86495 24870 86505 24988
rect 86367 24865 86505 24870
rect 85178 24732 85306 24759
rect 85178 24658 85207 24732
rect 85281 24658 85306 24732
rect 85178 24631 85306 24658
rect 86996 23907 87105 23928
rect 41218 23870 41366 23875
rect 41218 23742 41228 23870
rect 41356 23742 41366 23870
rect 41218 23737 41366 23742
rect 51058 23839 51196 23844
rect 51058 23721 51068 23839
rect 51186 23721 51196 23839
rect 51058 23716 51196 23721
rect 62978 23840 63116 23845
rect 62978 23722 62988 23840
rect 63106 23722 63116 23840
rect 62978 23717 63116 23722
rect 71547 23837 71685 23842
rect 71547 23719 71557 23837
rect 71675 23719 71685 23837
rect 86996 23833 87014 23907
rect 87088 23833 87105 23907
rect 86996 23809 87105 23833
rect 92580 23788 92718 23793
rect 71547 23714 71685 23719
rect 83045 23772 83183 23777
rect 83045 23654 83055 23772
rect 83173 23654 83183 23772
rect 83045 23649 83183 23654
rect 85581 23722 85719 23727
rect 41677 23590 41793 23622
rect 41677 23526 41701 23590
rect 41765 23526 41793 23590
rect 41677 23504 41793 23526
rect 52528 23580 52636 23609
rect 52528 23516 52551 23580
rect 52615 23516 52636 23580
rect 52528 23489 52636 23516
rect 64415 23588 64543 23624
rect 64415 23514 64440 23588
rect 64514 23514 64543 23588
rect 64415 23496 64543 23514
rect 72846 23592 72974 23618
rect 85581 23604 85591 23722
rect 85709 23604 85719 23722
rect 92580 23670 92590 23788
rect 92708 23670 92718 23788
rect 92580 23665 92718 23670
rect 85581 23599 85719 23604
rect 72846 23518 72870 23592
rect 72944 23518 72974 23592
rect 72846 23490 72974 23518
rect 81855 23543 81959 23568
rect 81855 23469 81872 23543
rect 81946 23469 81959 23543
rect 81855 23443 81959 23469
rect 93107 23542 93235 23569
rect 93107 23468 93131 23542
rect 93205 23468 93235 23542
rect 93107 23441 93235 23468
rect 103434 23108 103552 24172
rect 106362 23428 106510 23433
rect 106362 23300 106372 23428
rect 106500 23300 106510 23428
rect 106362 23295 106510 23300
rect 105384 23165 105512 23193
rect 105384 23091 105417 23165
rect 105491 23091 105512 23165
rect 105384 23065 105512 23091
rect 109004 23113 109122 24143
rect 103434 22984 103552 22990
rect 109004 22989 109122 22995
rect 39890 22775 40002 22808
rect 39890 22711 39914 22775
rect 39978 22711 40002 22775
rect 39890 22690 40002 22711
rect 50482 22768 50598 22793
rect 50482 22704 50506 22768
rect 50570 22704 50598 22768
rect 50482 22677 50598 22704
rect 62392 22765 62520 22784
rect 62392 22691 62415 22765
rect 62489 22691 62520 22765
rect 62392 22656 62520 22691
rect 71156 22766 71284 22796
rect 71156 22692 71181 22766
rect 71255 22692 71284 22766
rect 71156 22668 71284 22692
rect 83436 22716 83543 22732
rect 83436 22642 83454 22716
rect 83528 22642 83543 22716
rect 83436 22625 83543 22642
rect 91372 22717 91481 22738
rect 91372 22643 91387 22717
rect 91461 22643 91481 22717
rect 107980 22694 108096 22699
rect 107979 22693 108097 22694
rect 91372 22622 91481 22643
rect 104384 22674 104518 22682
rect 51930 22587 52068 22592
rect 40373 22578 40521 22583
rect 40373 22450 40383 22578
rect 40511 22450 40521 22578
rect 51930 22469 51940 22587
rect 52058 22469 52068 22587
rect 51930 22464 52068 22469
rect 63850 22582 63988 22587
rect 63850 22464 63860 22582
rect 63978 22464 63988 22582
rect 63850 22459 63988 22464
rect 72425 22578 72563 22583
rect 72425 22460 72435 22578
rect 72553 22460 72563 22578
rect 104384 22558 104394 22674
rect 104510 22558 104518 22674
rect 107979 22577 107980 22693
rect 108096 22577 108097 22693
rect 107979 22576 108097 22577
rect 107980 22571 108096 22576
rect 104384 22544 104518 22558
rect 91872 22528 92010 22533
rect 72425 22455 72563 22460
rect 82246 22522 82384 22527
rect 40373 22445 40521 22450
rect 82246 22404 82256 22522
rect 82374 22404 82384 22522
rect 91872 22410 91882 22528
rect 92000 22410 92010 22528
rect 91872 22405 92010 22410
rect 82246 22399 82384 22404
rect 107073 22355 107190 22373
rect 107073 22271 107090 22355
rect 107174 22271 107190 22355
rect 107073 22249 107190 22271
rect 105786 22156 105934 22161
rect 105786 22028 105796 22156
rect 105924 22028 105934 22156
rect 105786 22023 105934 22028
rect 36833 21883 36981 21888
rect 36833 21755 36843 21883
rect 36971 21755 36981 21883
rect 60229 21871 60367 21876
rect 36833 21750 36981 21755
rect 47785 21847 47933 21852
rect 47785 21719 47795 21847
rect 47923 21719 47933 21847
rect 60229 21753 60239 21871
rect 60357 21753 60367 21871
rect 60229 21748 60367 21753
rect 47785 21714 47933 21719
rect 43424 21662 43572 21667
rect 38290 21591 38393 21605
rect 38290 21517 38303 21591
rect 38377 21517 38393 21591
rect 43424 21534 43434 21662
rect 43562 21534 43572 21662
rect 61646 21589 61760 21607
rect 43424 21529 43572 21534
rect 48694 21584 48778 21589
rect 38290 21504 38393 21517
rect 48694 21520 48704 21584
rect 48768 21583 48778 21584
rect 48768 21520 49362 21583
rect 48694 21519 49362 21520
rect 49426 21519 49432 21583
rect 48694 21515 48778 21519
rect 61646 21515 61659 21589
rect 61733 21515 61760 21589
rect 61646 21495 61760 21515
rect 44370 21403 44436 21404
rect 44363 21399 44837 21403
rect 44363 21343 44375 21399
rect 44431 21343 44837 21399
rect 44363 21339 44837 21343
rect 44901 21339 44907 21403
rect 44370 21338 44436 21339
rect 36252 20773 36367 20795
rect 36252 20709 36278 20773
rect 36342 20709 36367 20773
rect 47727 20767 47811 20772
rect 36252 20686 36367 20709
rect 47036 20703 47042 20767
rect 47106 20703 47737 20767
rect 47801 20703 47811 20767
rect 47727 20698 47811 20703
rect 59676 20768 59788 20797
rect 59676 20694 59693 20768
rect 59767 20694 59788 20768
rect 67139 20795 67244 20815
rect 67139 20731 67161 20795
rect 67225 20731 67244 20795
rect 67139 20711 67244 20731
rect 67974 20792 68078 20808
rect 67974 20728 67989 20792
rect 68053 20728 68078 20792
rect 67974 20712 68078 20728
rect 59676 20665 59788 20694
rect 37628 20579 37776 20584
rect 37628 20451 37638 20579
rect 37766 20451 37776 20579
rect 42987 20582 43102 20610
rect 42987 20518 43010 20582
rect 43074 20518 43102 20582
rect 42987 20490 43102 20518
rect 48593 20577 48741 20582
rect 37628 20446 37776 20451
rect 48593 20449 48603 20577
rect 48731 20449 48741 20577
rect 61051 20579 61189 20584
rect 61051 20461 61061 20579
rect 61179 20461 61189 20579
rect 74007 20545 74118 20565
rect 74007 20481 74028 20545
rect 74092 20481 74118 20545
rect 74007 20463 74118 20481
rect 74825 20551 74936 20568
rect 74825 20487 74856 20551
rect 74920 20487 74936 20551
rect 74825 20469 74936 20487
rect 61051 20456 61189 20461
rect 48593 20444 48741 20449
rect 44250 20397 44398 20402
rect 44250 20269 44260 20397
rect 44388 20269 44398 20397
rect 44250 20264 44398 20269
rect 66639 20332 66777 20337
rect 66639 20214 66649 20332
rect 66767 20214 66777 20332
rect 66639 20209 66777 20214
rect 68376 20324 68514 20329
rect 68376 20206 68386 20324
rect 68504 20206 68514 20324
rect 68376 20201 68514 20206
rect 75266 20093 75404 20098
rect 73555 20070 73693 20075
rect 73555 19952 73565 20070
rect 73683 19952 73693 20070
rect 75266 19975 75276 20093
rect 75394 19975 75404 20093
rect 75266 19970 75404 19975
rect 73555 19947 73693 19952
rect 36833 19885 36981 19890
rect 36833 19757 36843 19885
rect 36971 19757 36981 19885
rect 36833 19752 36981 19757
rect 47781 19842 47929 19847
rect 47781 19714 47791 19842
rect 47919 19714 47929 19842
rect 60231 19841 60369 19846
rect 60231 19723 60241 19841
rect 60359 19723 60369 19841
rect 67140 19825 67248 19840
rect 67140 19761 67163 19825
rect 67227 19761 67248 19825
rect 67140 19744 67248 19761
rect 67972 19826 68071 19846
rect 67972 19762 67985 19826
rect 68049 19762 68071 19826
rect 67972 19745 68071 19762
rect 60231 19718 60369 19723
rect 47781 19709 47929 19714
rect 43405 19654 43553 19659
rect 38281 19592 38395 19617
rect 38281 19528 38307 19592
rect 38371 19528 38395 19592
rect 38281 19503 38395 19528
rect 43405 19526 43415 19654
rect 43543 19526 43553 19654
rect 43405 19521 43553 19526
rect 49338 19582 49447 19618
rect 49338 19518 49357 19582
rect 49421 19518 49447 19582
rect 49338 19484 49447 19518
rect 61647 19586 61757 19605
rect 61647 19512 61662 19586
rect 61736 19512 61757 19586
rect 61647 19496 61757 19512
rect 74009 19583 74122 19610
rect 74009 19519 74034 19583
rect 74098 19519 74122 19583
rect 74009 19498 74122 19519
rect 74827 19582 74938 19607
rect 74827 19518 74860 19582
rect 74924 19518 74938 19582
rect 74827 19497 74938 19518
rect 44359 19403 44443 19407
rect 44359 19402 44840 19403
rect 44359 19338 44369 19402
rect 44433 19339 44840 19402
rect 44904 19339 44910 19403
rect 44433 19338 44443 19339
rect 44359 19333 44443 19338
rect 36258 18771 36366 18796
rect 36258 18707 36280 18771
rect 36344 18707 36366 18771
rect 47725 18761 47809 18766
rect 36258 18682 36366 18707
rect 47034 18697 47040 18761
rect 47104 18697 47735 18761
rect 47799 18697 47809 18761
rect 47725 18692 47809 18697
rect 59678 18764 59793 18797
rect 59678 18700 59710 18764
rect 59774 18700 59793 18764
rect 59678 18672 59793 18700
rect 61045 18583 61183 18588
rect 37623 18578 37771 18583
rect 43408 18582 43474 18583
rect 37623 18450 37633 18578
rect 37761 18450 37771 18578
rect 43004 18518 43010 18582
rect 43074 18578 43474 18582
rect 43074 18522 43413 18578
rect 43469 18522 43474 18578
rect 43074 18518 43474 18522
rect 43408 18517 43474 18518
rect 48593 18578 48741 18583
rect 37623 18445 37771 18450
rect 48593 18450 48603 18578
rect 48731 18450 48741 18578
rect 61045 18465 61055 18583
rect 61173 18465 61183 18583
rect 61045 18460 61183 18465
rect 48593 18445 48741 18450
rect 44249 18389 44397 18394
rect 44249 18261 44259 18389
rect 44387 18261 44397 18389
rect 44249 18256 44397 18261
rect 40387 17866 40535 17871
rect 40387 17738 40397 17866
rect 40525 17738 40535 17866
rect 40387 17733 40535 17738
rect 51094 17840 51232 17845
rect 51094 17722 51104 17840
rect 51222 17722 51232 17840
rect 71574 17844 71712 17849
rect 51094 17717 51232 17722
rect 63005 17833 63143 17838
rect 63005 17715 63015 17833
rect 63133 17715 63143 17833
rect 71574 17726 71584 17844
rect 71702 17726 71712 17844
rect 92556 17819 92694 17824
rect 71574 17721 71712 17726
rect 82958 17813 83096 17818
rect 63005 17710 63143 17715
rect 82958 17695 82968 17813
rect 83086 17695 83096 17813
rect 92556 17701 92566 17819
rect 92684 17701 92694 17819
rect 92556 17696 92694 17701
rect 82958 17690 83096 17695
rect 41676 17587 41791 17615
rect 41676 17523 41702 17587
rect 41766 17523 41791 17587
rect 41676 17493 41791 17523
rect 52530 17580 52635 17605
rect 72856 17599 72969 17622
rect 52530 17516 52547 17580
rect 52611 17516 52635 17580
rect 52530 17494 52635 17516
rect 63932 17582 64016 17587
rect 63932 17518 63942 17582
rect 64006 17518 64442 17582
rect 64506 17518 64512 17582
rect 72856 17525 72877 17599
rect 72951 17525 72969 17599
rect 63932 17513 64016 17518
rect 72856 17503 72969 17525
rect 81856 17572 81959 17596
rect 81856 17498 81877 17572
rect 81951 17498 81959 17572
rect 92777 17567 92851 17572
rect 92777 17503 92782 17567
rect 92846 17503 93134 17567
rect 93198 17503 93204 17567
rect 92777 17498 92851 17503
rect 81856 17472 81959 17498
rect 86402 16962 86540 16967
rect 86402 16844 86412 16962
rect 86530 16844 86540 16962
rect 86402 16839 86540 16844
rect 39889 16765 39997 16794
rect 39889 16701 39911 16765
rect 39975 16701 39997 16765
rect 39889 16668 39997 16701
rect 50481 16762 50597 16796
rect 50481 16698 50503 16762
rect 50567 16698 50597 16762
rect 50481 16665 50597 16698
rect 62392 16768 62520 16792
rect 62392 16694 62416 16768
rect 62490 16694 62520 16768
rect 62392 16664 62520 16694
rect 71163 16779 71278 16799
rect 71163 16705 71185 16779
rect 71259 16705 71278 16779
rect 71163 16683 71278 16705
rect 83428 16752 83545 16779
rect 83428 16678 83450 16752
rect 83524 16678 83545 16752
rect 91375 16748 91489 16773
rect 83428 16655 83545 16678
rect 85186 16722 85301 16742
rect 85186 16648 85205 16722
rect 85279 16648 85301 16722
rect 85186 16630 85301 16648
rect 91375 16674 91397 16748
rect 91471 16674 91489 16748
rect 91375 16642 91489 16674
rect 51807 16582 51945 16587
rect 41201 16542 41349 16547
rect 41201 16414 41211 16542
rect 41339 16414 41349 16542
rect 51807 16464 51817 16582
rect 51935 16464 51945 16582
rect 72286 16582 72424 16587
rect 51807 16459 51945 16464
rect 63817 16573 63955 16578
rect 63817 16455 63827 16573
rect 63945 16455 63955 16573
rect 72286 16464 72296 16582
rect 72414 16464 72424 16582
rect 72286 16459 72424 16464
rect 82286 16561 82424 16566
rect 63817 16450 63955 16455
rect 82286 16443 82296 16561
rect 82414 16443 82424 16561
rect 82286 16438 82424 16443
rect 91849 16547 91987 16552
rect 91849 16429 91859 16547
rect 91977 16429 91987 16547
rect 91849 16424 91987 16429
rect 41201 16409 41349 16414
rect 86989 15897 87117 15921
rect 86989 15823 87011 15897
rect 87085 15823 87117 15897
rect 86989 15793 87117 15823
rect 85614 15695 85752 15700
rect 85614 15577 85624 15695
rect 85742 15577 85752 15695
rect 85614 15572 85752 15577
rect 42983 14533 43111 14539
rect 67124 14533 67252 14539
rect 67426 14533 67564 14538
rect 91367 14533 91495 14539
rect 105384 14533 105512 14539
rect 23789 14405 42983 14533
rect 43111 14405 67124 14533
rect 67252 14405 67431 14533
rect 67559 14405 91367 14533
rect 91495 14405 105384 14533
rect 105512 14405 125602 14533
rect 42983 14399 43111 14405
rect 67124 14399 67252 14405
rect 67426 14400 67564 14405
rect 91367 14399 91495 14405
rect 105384 14399 105512 14405
rect 44812 13991 44940 13997
rect 66749 13991 66887 13995
rect 67969 13991 68097 13997
rect 93107 13991 93235 13997
rect 107068 13991 107196 13997
rect 23789 13863 44812 13991
rect 44940 13990 67969 13991
rect 44940 13863 66754 13990
rect 44812 13857 44940 13863
rect 66749 13862 66754 13863
rect 66882 13863 67969 13990
rect 68097 13863 93107 13991
rect 93235 13863 107068 13991
rect 107196 13863 125602 13991
rect 66882 13862 66887 13863
rect 66749 13857 66887 13862
rect 67969 13857 68097 13863
rect 93107 13857 93235 13863
rect 107068 13857 107196 13863
rect 47010 12350 47138 12356
rect 71863 12350 72001 12353
rect 23789 12222 47010 12350
rect 47138 12348 120735 12350
rect 47138 12222 71868 12348
rect 47010 12216 47138 12222
rect 71863 12220 71868 12222
rect 71996 12222 120735 12348
rect 120863 12222 120869 12350
rect 71996 12220 72001 12222
rect 71863 12215 72001 12220
rect 49330 11808 49458 11814
rect 72405 11809 72543 11814
rect 72405 11808 72410 11809
rect 23789 11680 49330 11808
rect 49458 11681 72410 11808
rect 72538 11808 72543 11809
rect 72538 11681 121333 11808
rect 49458 11680 121333 11681
rect 121461 11680 121467 11808
rect 49330 11674 49458 11680
rect 72405 11676 72543 11680
rect 59672 11264 59800 11270
rect 72949 11264 73087 11265
rect 23789 11136 59672 11264
rect 59800 11260 121937 11264
rect 59800 11136 72954 11260
rect 59672 11130 59800 11136
rect 72949 11132 72954 11136
rect 73082 11136 121937 11260
rect 122065 11136 122071 11264
rect 73082 11132 73087 11136
rect 72949 11127 73087 11132
rect 73493 10738 73631 10743
rect 61642 10725 61770 10731
rect 73493 10725 73498 10738
rect 23789 10597 61642 10725
rect 61770 10610 73498 10725
rect 73626 10725 73631 10738
rect 73626 10610 122541 10725
rect 61770 10597 122541 10610
rect 122669 10597 122675 10725
rect 61642 10591 61770 10597
rect 64415 9084 64543 9090
rect 75119 9086 75257 9091
rect 75119 9084 75124 9086
rect 23789 8956 64415 9084
rect 64543 8958 75124 9084
rect 75252 9084 75257 9086
rect 75252 8958 123737 9084
rect 64543 8956 123737 8958
rect 123865 8956 123871 9084
rect 64415 8950 64543 8956
rect 75119 8953 75257 8956
rect 62392 8548 62520 8554
rect 75665 8552 75803 8557
rect 75665 8548 75670 8552
rect 23789 8420 62392 8548
rect 62520 8424 75670 8548
rect 75798 8548 75803 8552
rect 75798 8424 124335 8548
rect 62520 8420 124335 8424
rect 124463 8420 124469 8548
rect 62392 8414 62520 8420
rect 75665 8419 75803 8420
rect 76206 8003 76344 8008
rect 76206 7998 76211 8003
rect 23789 7870 52517 7998
rect 52645 7875 76211 7998
rect 76339 7998 76344 8003
rect 76339 7875 124939 7998
rect 52645 7870 124939 7875
rect 125067 7870 125073 7998
rect 50477 7462 50605 7468
rect 76754 7464 76892 7469
rect 76754 7462 76759 7464
rect 23789 7334 50477 7462
rect 50605 7336 76759 7462
rect 76887 7462 76892 7464
rect 76887 7336 125537 7462
rect 50605 7334 125537 7336
rect 125665 7334 125671 7462
rect 50477 7328 50605 7334
rect 76754 7331 76892 7334
rect 144621 7265 166969 7662
rect 141092 7205 166969 7265
rect 79471 5833 79609 5838
rect 39882 5821 40010 5827
rect 79471 5821 79476 5833
rect 23789 5693 39882 5821
rect 40010 5809 79476 5821
rect 40010 5693 76521 5809
rect 39882 5687 40010 5693
rect 76515 5685 76521 5693
rect 76645 5705 79476 5809
rect 79604 5821 79609 5833
rect 85178 5821 85306 5827
rect 79604 5705 85178 5821
rect 76645 5693 85178 5705
rect 85306 5797 126739 5821
rect 85306 5693 111040 5797
rect 76645 5685 76651 5693
rect 85178 5687 85306 5693
rect 111034 5679 111040 5693
rect 111158 5693 126739 5797
rect 126867 5693 126873 5821
rect 111158 5679 111164 5693
rect 80015 5294 80153 5299
rect 41670 5284 41798 5290
rect 80015 5284 80020 5294
rect 23789 5156 41670 5284
rect 41798 5268 80020 5284
rect 41798 5156 76910 5268
rect 41670 5150 41798 5156
rect 76904 5146 76910 5156
rect 77032 5166 80020 5268
rect 80148 5284 80153 5294
rect 86989 5284 87117 5290
rect 80148 5166 86989 5284
rect 77032 5156 86989 5166
rect 87117 5273 127339 5284
rect 87117 5157 111439 5273
rect 111555 5157 127339 5273
rect 87117 5156 127339 5157
rect 127467 5156 127473 5284
rect 77032 5146 77038 5156
rect 86989 5150 87117 5156
rect 27434 4739 27562 4745
rect 80557 4742 80695 4747
rect 80557 4739 80562 4742
rect 23789 4611 27434 4739
rect 27562 4726 80562 4739
rect 27562 4611 74000 4726
rect 27434 4605 27562 4611
rect 73994 4600 74000 4611
rect 74126 4614 80562 4726
rect 80690 4739 80695 4742
rect 89566 4739 89694 4745
rect 80690 4614 89566 4739
rect 74126 4611 89566 4614
rect 89694 4611 127933 4739
rect 128061 4611 128067 4739
rect 74126 4600 74132 4611
rect 80557 4609 80695 4611
rect 89566 4605 89694 4611
rect 26623 4191 26751 4197
rect 74813 4191 74941 4197
rect 81101 4194 81239 4199
rect 81101 4191 81106 4194
rect 23789 4063 26623 4191
rect 26751 4063 74813 4191
rect 74941 4066 81106 4191
rect 81234 4191 81239 4194
rect 88514 4191 88642 4197
rect 81234 4066 88514 4191
rect 74941 4063 88514 4066
rect 88642 4063 128545 4191
rect 128673 4063 128679 4191
rect 26623 4057 26751 4063
rect 74813 4057 74941 4063
rect 81101 4061 81239 4063
rect 88514 4057 88642 4063
rect 25661 2563 25789 2569
rect 72846 2563 72974 2569
rect 79093 2563 79221 2569
rect 82743 2566 82881 2571
rect 82743 2563 82748 2566
rect 23789 2435 25661 2563
rect 25789 2435 72846 2563
rect 72974 2435 79093 2563
rect 79221 2438 82748 2563
rect 82876 2563 82881 2566
rect 82876 2438 129748 2563
rect 79221 2435 129748 2438
rect 129876 2435 129882 2563
rect 25661 2429 25789 2435
rect 72846 2429 72974 2435
rect 79093 2429 79221 2435
rect 82743 2433 82881 2435
rect 24761 2017 24889 2023
rect 71156 2017 71284 2023
rect 78108 2017 78236 2023
rect 83284 2017 83422 2021
rect 23789 1889 24761 2017
rect 24889 1889 71156 2017
rect 71284 1889 78108 2017
rect 78236 2016 130331 2017
rect 78236 1889 83289 2016
rect 24761 1883 24889 1889
rect 71156 1883 71284 1889
rect 78108 1883 78236 1889
rect 83284 1888 83289 1889
rect 83417 1889 130331 2016
rect 130459 1889 130465 2017
rect 83417 1888 83422 1889
rect 83284 1883 83422 1888
rect 38277 1466 38405 1472
rect 83425 1466 83553 1472
rect 83825 1471 83963 1476
rect 83825 1466 83830 1471
rect 23789 1338 38277 1466
rect 38405 1459 83425 1466
rect 38405 1338 76122 1459
rect 38277 1332 38405 1338
rect 76116 1333 76122 1338
rect 76248 1338 83425 1459
rect 83553 1343 83830 1466
rect 83958 1466 83963 1471
rect 83958 1458 119412 1466
rect 83958 1343 110635 1458
rect 83553 1338 110635 1343
rect 110755 1338 119412 1458
rect 119540 1338 130936 1466
rect 131064 1338 131070 1466
rect 76248 1333 76254 1338
rect 83425 1332 83553 1338
rect 84364 948 84502 953
rect 36248 935 36376 941
rect 81845 935 81973 941
rect 84364 935 84369 948
rect 23789 807 36248 935
rect 36376 919 81845 935
rect 36376 807 75721 919
rect 36248 801 36376 807
rect 75715 793 75721 807
rect 75847 807 81845 919
rect 81973 820 84369 935
rect 84497 935 84502 948
rect 84497 931 131530 935
rect 84497 820 110236 931
rect 81973 811 110236 820
rect 110356 811 131530 931
rect 81973 807 131530 811
rect 131658 807 131670 935
rect 75847 793 75853 807
rect 81845 801 81973 807
rect 133768 687 133838 692
rect 141092 687 141152 7205
rect 144621 6662 166969 7205
rect 144621 5159 166969 5662
rect 133768 627 133773 687
rect 133833 627 141152 687
rect 142004 5099 166969 5159
rect 133768 622 133838 627
rect 134336 350 134406 355
rect 142004 350 142064 5099
rect 144621 4662 166969 5099
rect 134336 290 134341 350
rect 134401 290 142064 350
rect 134336 285 134406 290
rect 122561 158 122627 164
rect 122533 92 122561 158
rect 122627 92 132805 158
rect 122561 86 122627 92
rect 132460 -100 132536 -96
rect 128552 -166 128558 -100
rect 128624 -101 132536 -100
rect 128624 -166 132465 -101
rect 132460 -167 132465 -166
rect 132531 -167 132536 -101
rect 132460 -172 132536 -167
rect 132739 -216 132805 92
rect 135392 33 135885 38
rect 135392 -36 135402 33
rect 135875 -36 135885 33
rect 135392 -41 135885 -36
rect 132892 -54 134313 -49
rect 132892 -110 132897 -54
rect 132953 -110 134313 -54
rect 132892 -115 134313 -110
rect 134057 -214 134143 -209
rect 134247 -211 134313 -115
rect 141774 -188 141844 -183
rect 143469 -188 143535 -185
rect 133922 -216 133988 -214
rect 134057 -216 134067 -214
rect 132739 -282 134067 -216
rect 134133 -282 134143 -214
rect 134057 -287 134143 -282
rect 134237 -216 134323 -211
rect 134237 -284 134247 -216
rect 134313 -284 134323 -216
rect 141774 -248 141779 -188
rect 141839 -190 143535 -188
rect 141839 -246 143474 -190
rect 143530 -246 143535 -190
rect 141839 -248 143535 -246
rect 141774 -253 141844 -248
rect 143469 -251 143535 -248
rect 134237 -289 134323 -284
rect 132462 -399 132538 -394
rect 121973 -465 121979 -399
rect 122045 -465 132467 -399
rect 132533 -465 132538 -399
rect 132462 -470 132538 -465
rect 139072 -513 139554 -508
rect 139072 -577 139082 -513
rect 139544 -577 139554 -513
rect 139072 -582 139554 -577
rect 132462 -666 132538 -661
rect 127941 -732 127947 -666
rect 128013 -732 132467 -666
rect 132533 -732 132538 -666
rect 132462 -737 132538 -732
rect 144621 -818 166969 -338
rect 144198 -878 166969 -818
rect 123737 -1225 123743 -1159
rect 123809 -1225 132805 -1159
rect 132460 -1417 132536 -1413
rect 129760 -1483 129766 -1417
rect 129832 -1418 132536 -1417
rect 129832 -1483 132465 -1418
rect 132460 -1484 132465 -1483
rect 132531 -1484 132536 -1418
rect 132460 -1489 132536 -1484
rect 132739 -1533 132805 -1225
rect 135395 -1282 135888 -1277
rect 135395 -1351 135405 -1282
rect 135878 -1351 135888 -1282
rect 135395 -1356 135888 -1351
rect 132892 -1371 134313 -1366
rect 132892 -1427 132897 -1371
rect 132953 -1427 134313 -1371
rect 132892 -1432 134313 -1427
rect 134057 -1531 134143 -1526
rect 134247 -1528 134313 -1432
rect 141774 -1505 141844 -1500
rect 143163 -1505 143229 -1502
rect 133922 -1533 133988 -1531
rect 134057 -1533 134067 -1531
rect 132739 -1599 134067 -1533
rect 134133 -1599 134143 -1531
rect 134057 -1604 134143 -1599
rect 134237 -1533 134323 -1528
rect 134237 -1601 134247 -1533
rect 134313 -1601 134323 -1533
rect 141774 -1565 141779 -1505
rect 141839 -1507 143229 -1505
rect 141839 -1563 143168 -1507
rect 143224 -1563 143229 -1507
rect 141839 -1565 143229 -1563
rect 141774 -1570 141844 -1565
rect 143163 -1568 143229 -1565
rect 134237 -1606 134323 -1601
rect 132462 -1716 132538 -1711
rect 124347 -1782 124353 -1716
rect 124419 -1782 132467 -1716
rect 132533 -1782 132538 -1716
rect 132462 -1787 132538 -1782
rect 139082 -1827 139564 -1822
rect 139082 -1891 139092 -1827
rect 139554 -1891 139564 -1827
rect 139082 -1896 139564 -1891
rect 130362 -1983 130428 -1977
rect 132462 -1983 132538 -1978
rect 67093 -2039 67180 -2034
rect 67093 -2665 67103 -2039
rect 67170 -2665 67180 -2039
rect 130428 -2049 132467 -1983
rect 132533 -2049 132538 -1983
rect 130362 -2055 130428 -2049
rect 132462 -2054 132538 -2049
rect 133768 -2277 133838 -2272
rect 144198 -2277 144258 -878
rect 144621 -1338 166969 -878
rect 133768 -2337 133773 -2277
rect 133833 -2337 144258 -2277
rect 133768 -2342 133838 -2337
rect 67093 -2670 67180 -2665
rect 134336 -2614 134406 -2609
rect 144621 -2614 166969 -2338
rect 134336 -2674 134341 -2614
rect 134401 -2674 166969 -2614
rect 134336 -2679 134406 -2674
rect 121362 -2872 121368 -2806
rect 121434 -2872 132805 -2806
rect 132460 -3064 132536 -3060
rect 127358 -3130 127364 -3064
rect 127430 -3065 132536 -3064
rect 127430 -3130 132465 -3065
rect 132460 -3131 132465 -3130
rect 132531 -3131 132536 -3065
rect 132460 -3136 132536 -3131
rect 132739 -3180 132805 -2872
rect 135387 -2928 135880 -2923
rect 135387 -2997 135397 -2928
rect 135870 -2997 135880 -2928
rect 135387 -3002 135880 -2997
rect 132892 -3018 134313 -3013
rect 132892 -3074 132897 -3018
rect 132953 -3074 134313 -3018
rect 132892 -3079 134313 -3074
rect 134057 -3178 134143 -3173
rect 134247 -3175 134313 -3079
rect 141774 -3152 141844 -3147
rect 142771 -3152 142837 -3149
rect 133922 -3180 133988 -3178
rect 134057 -3180 134067 -3178
rect 132739 -3246 134067 -3180
rect 134133 -3246 134143 -3178
rect 134057 -3251 134143 -3246
rect 134237 -3180 134323 -3175
rect 134237 -3248 134247 -3180
rect 134313 -3248 134323 -3180
rect 141774 -3212 141779 -3152
rect 141839 -3154 142837 -3152
rect 141839 -3210 142776 -3154
rect 142832 -3210 142837 -3154
rect 141839 -3212 142837 -3210
rect 141774 -3217 141844 -3212
rect 142771 -3215 142837 -3212
rect 134237 -3253 134323 -3248
rect 144621 -3338 166969 -2674
rect 132462 -3363 132538 -3358
rect 120751 -3429 120757 -3363
rect 120823 -3429 132467 -3363
rect 132533 -3429 132538 -3363
rect 132462 -3434 132538 -3429
rect 139072 -3477 139554 -3472
rect 139072 -3541 139082 -3477
rect 139544 -3541 139554 -3477
rect 139072 -3546 139554 -3541
rect 132462 -3630 132538 -3625
rect 126757 -3696 126763 -3630
rect 126829 -3696 132467 -3630
rect 132533 -3696 132538 -3630
rect 132462 -3701 132538 -3696
rect 124952 -4119 124958 -4053
rect 125024 -4119 132805 -4053
rect 130963 -4311 131029 -4305
rect 132460 -4311 132536 -4307
rect 131029 -4312 132536 -4311
rect 131029 -4377 132465 -4312
rect 130963 -4383 131029 -4377
rect 132460 -4378 132465 -4377
rect 132531 -4378 132536 -4312
rect 132460 -4383 132536 -4378
rect 132739 -4427 132805 -4119
rect 135389 -4178 135882 -4173
rect 135389 -4247 135399 -4178
rect 135872 -4247 135882 -4178
rect 135389 -4252 135882 -4247
rect 132892 -4265 134313 -4260
rect 132892 -4321 132897 -4265
rect 132953 -4321 134313 -4265
rect 132892 -4326 134313 -4321
rect 134057 -4425 134143 -4420
rect 134247 -4422 134313 -4326
rect 141774 -4399 141844 -4394
rect 142365 -4399 142431 -4396
rect 133922 -4427 133988 -4425
rect 134057 -4427 134067 -4425
rect 132739 -4493 134067 -4427
rect 134133 -4493 134143 -4425
rect 134057 -4498 134143 -4493
rect 134237 -4427 134323 -4422
rect 134237 -4495 134247 -4427
rect 134313 -4495 134323 -4427
rect 141774 -4459 141779 -4399
rect 141839 -4401 142431 -4399
rect 141839 -4457 142370 -4401
rect 142426 -4457 142431 -4401
rect 141839 -4459 142431 -4457
rect 141774 -4464 141844 -4459
rect 142365 -4462 142431 -4459
rect 134237 -4500 134323 -4495
rect 132462 -4610 132538 -4605
rect 125562 -4676 125568 -4610
rect 125634 -4676 132467 -4610
rect 132533 -4676 132538 -4610
rect 132462 -4681 132538 -4676
rect 139087 -4724 139569 -4719
rect 139087 -4788 139097 -4724
rect 139559 -4788 139569 -4724
rect 139087 -4793 139569 -4788
rect 132462 -4877 132538 -4872
rect 131550 -4943 131556 -4877
rect 131622 -4943 132467 -4877
rect 132533 -4943 132538 -4877
rect 132462 -4948 132538 -4943
rect 66550 -5627 66637 -5622
rect 66550 -6253 66560 -5627
rect 66627 -6253 66637 -5627
rect 66550 -6258 66637 -6253
rect 71071 -5629 71150 -5624
rect 71071 -6267 71081 -5629
rect 71140 -6267 71150 -5629
rect 71071 -6272 71150 -6267
rect 74335 -5629 74414 -5624
rect 74335 -6267 74345 -5629
rect 74404 -6267 74414 -5629
rect 74335 -6272 74414 -6267
rect 77599 -5629 77678 -5624
rect 77599 -6267 77609 -5629
rect 77668 -6267 77678 -5629
rect 77599 -6272 77678 -6267
rect 78687 -5629 78766 -5624
rect 78687 -6267 78697 -5629
rect 78756 -6267 78766 -5629
rect 78687 -6272 78766 -6267
rect 81951 -5629 82030 -5624
rect 81951 -6267 81961 -5629
rect 82020 -6267 82030 -5629
rect 81951 -6272 82030 -6267
rect 85215 -5629 85294 -5624
rect 85215 -6267 85225 -5629
rect 85284 -6267 85294 -5629
rect 85215 -6272 85294 -6267
rect 67015 -6683 67352 -6678
rect 67015 -6811 67121 -6683
rect 67249 -6811 67352 -6683
rect 67015 -7736 67352 -6811
rect 66690 -40917 67690 -7736
rect 71618 -8627 71697 -8622
rect 71618 -9265 71628 -8627
rect 71687 -9265 71697 -8627
rect 71618 -9270 71697 -9265
rect 72706 -8627 72785 -8622
rect 72706 -9265 72716 -8627
rect 72775 -9265 72785 -8627
rect 72706 -9270 72785 -9265
rect 73794 -8627 73873 -8622
rect 73794 -9265 73804 -8627
rect 73863 -9265 73873 -8627
rect 73794 -9270 73873 -9265
rect 74882 -8627 74961 -8622
rect 74882 -9265 74892 -8627
rect 74951 -9265 74961 -8627
rect 74882 -9270 74961 -9265
rect 75970 -8627 76049 -8622
rect 75970 -9265 75980 -8627
rect 76039 -9265 76049 -8627
rect 75970 -9270 76049 -9265
rect 77058 -8627 77137 -8622
rect 77058 -9265 77068 -8627
rect 77127 -9265 77137 -8627
rect 77058 -9270 77137 -9265
rect 78146 -8627 78225 -8622
rect 78146 -9265 78156 -8627
rect 78215 -9265 78225 -8627
rect 78146 -9270 78225 -9265
rect 79234 -8627 79313 -8622
rect 79234 -9265 79244 -8627
rect 79303 -9265 79313 -8627
rect 79234 -9270 79313 -9265
rect 80322 -8627 80401 -8622
rect 80322 -9265 80332 -8627
rect 80391 -9265 80401 -8627
rect 80322 -9270 80401 -9265
rect 81410 -8627 81489 -8622
rect 81410 -9265 81420 -8627
rect 81479 -9265 81489 -8627
rect 81410 -9270 81489 -9265
rect 82498 -8627 82577 -8622
rect 82498 -9265 82508 -8627
rect 82567 -9265 82577 -8627
rect 82498 -9270 82577 -9265
rect 83586 -8627 83665 -8622
rect 83586 -9265 83596 -8627
rect 83655 -9265 83665 -8627
rect 83586 -9270 83665 -9265
rect 84674 -8627 84753 -8622
rect 84674 -9265 84684 -8627
rect 84743 -9265 84753 -8627
rect 84674 -9270 84753 -9265
rect 155440 -10846 166970 -10364
rect 154392 -10906 166970 -10846
rect 143473 -11039 144737 -11034
rect 143473 -11095 143478 -11039
rect 143534 -11095 144737 -11039
rect 143473 -11100 144737 -11095
rect 144392 -11292 144468 -11288
rect 143163 -11293 144468 -11292
rect 143163 -11297 144397 -11293
rect 143163 -11353 143168 -11297
rect 143224 -11353 144397 -11297
rect 143163 -11358 144397 -11353
rect 144392 -11359 144397 -11358
rect 144463 -11359 144468 -11293
rect 144392 -11364 144468 -11359
rect 144671 -11408 144737 -11100
rect 147319 -11156 147812 -11151
rect 147319 -11225 147329 -11156
rect 147802 -11225 147812 -11156
rect 147319 -11230 147812 -11225
rect 144824 -11246 146245 -11241
rect 144824 -11302 144829 -11246
rect 144885 -11302 146245 -11246
rect 144824 -11307 146245 -11302
rect 145989 -11406 146075 -11401
rect 146179 -11403 146245 -11307
rect 153839 -11380 153909 -11375
rect 154392 -11380 154452 -10906
rect 155440 -11364 166970 -10906
rect 145854 -11408 145920 -11406
rect 145989 -11408 145999 -11406
rect 144671 -11474 145999 -11408
rect 146065 -11474 146075 -11406
rect 145989 -11479 146075 -11474
rect 146169 -11408 146255 -11403
rect 146169 -11476 146179 -11408
rect 146245 -11476 146255 -11408
rect 153839 -11440 153844 -11380
rect 153904 -11440 154452 -11380
rect 153839 -11445 153909 -11440
rect 146169 -11481 146255 -11476
rect 144394 -11591 144470 -11586
rect 144358 -11592 144399 -11591
rect 142773 -11597 144399 -11592
rect 142773 -11653 142778 -11597
rect 142834 -11653 144399 -11597
rect 142773 -11657 144399 -11653
rect 144465 -11657 144470 -11591
rect 142773 -11658 144470 -11657
rect 144394 -11662 144470 -11658
rect 151004 -11705 151486 -11700
rect 151004 -11769 151014 -11705
rect 151476 -11769 151486 -11705
rect 151004 -11774 151486 -11769
rect 144394 -11858 144470 -11853
rect 142363 -11863 144399 -11858
rect 142363 -11919 142368 -11863
rect 142424 -11919 144399 -11863
rect 142363 -11924 144399 -11919
rect 144465 -11924 144470 -11858
rect 144394 -11929 144470 -11924
rect 145700 -12190 145770 -12185
rect 145700 -12250 145705 -12190
rect 145765 -12250 154910 -12190
rect 145700 -12255 145770 -12250
rect 146268 -12620 146338 -12615
rect 146268 -12680 146273 -12620
rect 146333 -12680 153882 -12620
rect 146268 -12685 146338 -12680
rect 71069 -13627 71148 -13622
rect 71069 -14265 71079 -13627
rect 71138 -14265 71148 -13627
rect 71069 -14270 71148 -14265
rect 72157 -13627 72236 -13622
rect 72157 -14265 72167 -13627
rect 72226 -14265 72236 -13627
rect 72157 -14270 72236 -14265
rect 73245 -13627 73324 -13622
rect 73245 -14265 73255 -13627
rect 73314 -14265 73324 -13627
rect 73245 -14270 73324 -14265
rect 74333 -13627 74412 -13622
rect 74333 -14265 74343 -13627
rect 74402 -14265 74412 -13627
rect 74333 -14270 74412 -14265
rect 75421 -13627 75500 -13622
rect 75421 -14265 75431 -13627
rect 75490 -14265 75500 -13627
rect 75421 -14270 75500 -14265
rect 76509 -13627 76588 -13622
rect 76509 -14265 76519 -13627
rect 76578 -14265 76588 -13627
rect 76509 -14270 76588 -14265
rect 77597 -13627 77676 -13622
rect 77597 -14265 77607 -13627
rect 77666 -14265 77676 -13627
rect 77597 -14270 77676 -14265
rect 78685 -13627 78764 -13622
rect 78685 -14265 78695 -13627
rect 78754 -14265 78764 -13627
rect 78685 -14270 78764 -14265
rect 79773 -13627 79852 -13622
rect 79773 -14265 79783 -13627
rect 79842 -14265 79852 -13627
rect 79773 -14270 79852 -14265
rect 80861 -13627 80940 -13622
rect 80861 -14265 80871 -13627
rect 80930 -14265 80940 -13627
rect 80861 -14270 80940 -14265
rect 81949 -13627 82028 -13622
rect 81949 -14265 81959 -13627
rect 82018 -14265 82028 -13627
rect 81949 -14270 82028 -14265
rect 83037 -13627 83116 -13622
rect 83037 -14265 83047 -13627
rect 83106 -14265 83116 -13627
rect 83037 -14270 83116 -14265
rect 84125 -13627 84204 -13622
rect 84125 -14265 84135 -13627
rect 84194 -14265 84204 -13627
rect 84125 -14270 84204 -14265
rect 85213 -13627 85292 -13622
rect 85213 -14265 85223 -13627
rect 85282 -14265 85292 -13627
rect 85213 -14270 85292 -14265
rect 153822 -15232 153882 -12680
rect 154850 -12954 154910 -12250
rect 155440 -12954 166970 -12484
rect 154850 -13014 166970 -12954
rect 155440 -13484 166970 -13014
rect 155440 -15232 166970 -14766
rect 153822 -15292 166970 -15232
rect 155440 -15766 166970 -15292
rect 71611 -16617 71695 -16612
rect 71611 -17271 71621 -16617
rect 71685 -17271 71695 -16617
rect 71611 -17276 71695 -17271
rect 72699 -16617 72783 -16612
rect 72699 -17271 72709 -16617
rect 72773 -17271 72783 -16617
rect 72699 -17276 72783 -17271
rect 73787 -16617 73871 -16612
rect 73787 -17271 73797 -16617
rect 73861 -17271 73871 -16617
rect 73787 -17276 73871 -17271
rect 74875 -16617 74959 -16612
rect 74875 -17271 74885 -16617
rect 74949 -17271 74959 -16617
rect 74875 -17276 74959 -17271
rect 75963 -16617 76047 -16612
rect 75963 -17271 75973 -16617
rect 76037 -17271 76047 -16617
rect 75963 -17276 76047 -17271
rect 77051 -16617 77135 -16612
rect 77051 -17271 77061 -16617
rect 77125 -17271 77135 -16617
rect 77051 -17276 77135 -17271
rect 78139 -16617 78223 -16612
rect 78139 -17271 78149 -16617
rect 78213 -17271 78223 -16617
rect 78139 -17276 78223 -17271
rect 79227 -16617 79311 -16612
rect 79227 -17271 79237 -16617
rect 79301 -17271 79311 -16617
rect 79227 -17276 79311 -17271
rect 80315 -16617 80399 -16612
rect 80315 -17271 80325 -16617
rect 80389 -17271 80399 -16617
rect 80315 -17276 80399 -17271
rect 81403 -16617 81487 -16612
rect 81403 -17271 81413 -16617
rect 81477 -17271 81487 -16617
rect 81403 -17276 81487 -17271
rect 82491 -16617 82575 -16612
rect 82491 -17271 82501 -16617
rect 82565 -17271 82575 -16617
rect 82491 -17276 82575 -17271
rect 83579 -16617 83663 -16612
rect 83579 -17271 83589 -16617
rect 83653 -17271 83663 -16617
rect 83579 -17276 83663 -17271
rect 84667 -16617 84751 -16612
rect 84667 -17271 84677 -16617
rect 84741 -17271 84751 -16617
rect 84667 -17276 84751 -17271
rect 71065 -21612 71152 -21607
rect 71065 -22006 71075 -21612
rect 71142 -22006 71152 -21612
rect 71065 -22011 71152 -22006
rect 72155 -21618 72242 -21613
rect 72155 -22012 72165 -21618
rect 72232 -22012 72242 -21618
rect 72155 -22017 72242 -22012
rect 73243 -21618 73330 -21613
rect 73243 -22012 73253 -21618
rect 73320 -22012 73330 -21618
rect 73243 -22017 73330 -22012
rect 74331 -21618 74418 -21613
rect 74331 -22012 74341 -21618
rect 74408 -22012 74418 -21618
rect 74331 -22017 74418 -22012
rect 75419 -21618 75506 -21613
rect 75419 -22012 75429 -21618
rect 75496 -22012 75506 -21618
rect 75419 -22017 75506 -22012
rect 76507 -21618 76594 -21613
rect 76507 -22012 76517 -21618
rect 76584 -22012 76594 -21618
rect 76507 -22017 76594 -22012
rect 77595 -21618 77682 -21613
rect 77595 -22012 77605 -21618
rect 77672 -22012 77682 -21618
rect 77595 -22017 77682 -22012
rect 81947 -21618 82034 -21613
rect 81947 -22012 81957 -21618
rect 82024 -22012 82034 -21618
rect 81947 -22017 82034 -22012
rect 83035 -21618 83122 -21613
rect 83035 -22012 83045 -21618
rect 83112 -22012 83122 -21618
rect 83035 -22017 83122 -22012
rect 84123 -21618 84210 -21613
rect 84123 -22012 84133 -21618
rect 84200 -22012 84210 -21618
rect 84123 -22017 84210 -22012
rect 85211 -21618 85298 -21613
rect 85211 -22012 85221 -21618
rect 85288 -22012 85298 -21618
rect 85211 -22017 85298 -22012
rect 77486 -22175 78496 -22170
rect 77486 -23175 77491 -22175
rect 78491 -23175 78496 -22175
rect 77486 -23180 78496 -23175
rect 77491 -40917 78491 -23180
<< via3 >>
rect 35285 67107 35410 70423
rect 38294 67113 38442 70399
rect 42295 67110 42410 70392
rect 45277 67092 45431 70421
rect 56700 67113 56848 70393
rect 59712 67113 59864 70398
rect 63788 67105 63951 70396
rect 66804 67117 66952 70395
rect 73794 67107 73935 70398
rect 76799 67113 76934 70396
rect 84670 67112 84798 70393
rect 87663 67108 87817 70406
rect 92977 67100 93119 70406
rect 95985 67112 96113 70403
rect 102317 67100 102459 70406
rect 105325 67112 105453 70403
rect 62908 64980 63133 65047
rect 63684 64989 63797 65102
rect 64232 64976 64460 65055
rect 65058 64998 65171 65111
rect 65616 64980 65843 65055
rect 66421 64998 66534 65111
rect 66997 64982 67225 65054
rect 67770 64999 67883 65112
rect 72908 64980 73133 65047
rect 73684 64989 73797 65102
rect 74232 64976 74460 65055
rect 75058 64998 75171 65111
rect 75616 64980 75843 65055
rect 76421 64998 76534 65111
rect 76997 64982 77225 65054
rect 77770 64999 77883 65112
rect 85128 63757 85318 63849
rect 85568 63736 86002 63823
rect 86485 63764 86629 63858
rect 86904 63732 87328 63809
rect 102782 63757 102972 63849
rect 103222 63736 103656 63823
rect 104139 63764 104283 63858
rect 104558 63732 104982 63809
rect 85219 62237 85311 62346
rect 86550 62232 86642 62341
rect 102873 62237 102965 62346
rect 104204 62232 104296 62341
rect 62731 62076 62844 62189
rect 63429 62033 63542 62146
rect 64378 62045 64491 62159
rect 64721 62064 64834 62177
rect 65456 62056 65569 62169
rect 66175 62038 66288 62151
rect 66828 62030 66941 62143
rect 67543 62038 67656 62151
rect 72731 62076 72844 62189
rect 73429 62033 73542 62146
rect 74378 62045 74491 62159
rect 74721 62064 74834 62177
rect 75456 62056 75569 62169
rect 76175 62038 76288 62151
rect 76828 62030 76941 62143
rect 77543 62038 77656 62151
rect 63163 61245 63234 61352
rect 63705 61242 63776 61346
rect 65884 61349 65952 61473
rect 64251 61184 64320 61330
rect 64798 61191 64862 61321
rect 66426 61207 66494 61364
rect 66971 61261 67043 61383
rect 67514 61202 67580 61356
rect 73163 61245 73234 61352
rect 73705 61242 73776 61346
rect 75884 61349 75952 61473
rect 74251 61184 74320 61330
rect 74798 61191 74862 61321
rect 76426 61207 76494 61364
rect 76971 61261 77043 61383
rect 77514 61202 77580 61356
rect 65343 60862 65410 61015
rect 75343 60862 75410 61015
rect 86094 60357 86159 60499
rect 103748 60357 103813 60499
rect 85544 60170 85615 60274
rect 86636 60170 86704 60280
rect 103198 60170 103269 60274
rect 104290 60170 104358 60280
rect 63052 59916 63305 59993
rect 64372 59915 64680 60000
rect 65760 59918 66042 59989
rect 67132 59920 67414 59991
rect 73052 59916 73305 59993
rect 74372 59915 74680 60000
rect 75760 59918 76042 59989
rect 77132 59920 77414 59991
rect 84943 59523 85056 59636
rect 102597 59523 102710 59636
rect 63937 59238 64050 59351
rect 65298 59250 65411 59363
rect 66660 59268 66773 59381
rect 68044 59303 68157 59416
rect 73937 59238 74050 59351
rect 75298 59250 75411 59363
rect 76660 59268 76773 59381
rect 78044 59303 78157 59416
rect 87336 58917 87449 59030
rect 104990 58917 105103 59030
rect 27435 52542 27561 52668
rect 116738 52386 116866 52514
rect 120662 52363 120933 52467
rect 46153 51695 46271 52282
rect 47493 51229 47608 51852
rect 48197 51690 48307 52230
rect 49511 51249 49654 51907
rect 45803 50796 45929 50922
rect 24762 50508 24888 50634
rect 36202 49483 36285 49927
rect 37447 49792 37567 50285
rect 38144 49278 38243 49857
rect 39493 49780 39608 50313
rect 25662 48931 25788 49057
rect 26624 48203 26750 48329
rect 45802 48202 45930 48330
rect 56046 46741 56330 47379
rect 60492 47109 61496 47309
rect 62848 49465 63380 49622
rect 62010 41599 62280 42674
rect 36688 40605 36826 40610
rect 36688 40477 36693 40605
rect 36693 40477 36821 40605
rect 36821 40477 36826 40605
rect 36688 40472 36826 40477
rect 44960 40528 45098 40533
rect 44960 40400 44965 40528
rect 44965 40400 45093 40528
rect 45093 40400 45098 40528
rect 44960 40395 45098 40400
rect 62857 41596 63127 42671
rect 63412 41747 63617 42335
rect 56027 38731 56167 39355
rect 50243 32667 50361 32672
rect 40666 32643 40784 32648
rect 40666 32525 40779 32643
rect 40779 32525 40784 32643
rect 40666 32520 40784 32525
rect 50243 32549 50356 32667
rect 50356 32549 50361 32667
rect 50243 32544 50361 32549
rect 55952 30754 56299 31354
rect 60986 29648 61191 30188
rect 115289 51273 115385 51725
rect 117729 51316 117832 51778
rect 119326 51001 119407 52130
rect 121709 51027 121804 52123
rect 115579 50800 115707 50928
rect 117396 50869 117553 50953
rect 115989 50709 116141 50861
rect 119936 50772 120225 50944
rect 121196 50888 121516 50958
rect 66174 50013 66362 50207
rect 67970 49987 68198 50219
rect 69664 49968 69892 50200
rect 71483 49979 71711 50211
rect 73267 49976 73495 50208
rect 75052 49974 75280 50206
rect 100698 50019 100886 50213
rect 102494 49993 102722 50225
rect 104188 49974 104416 50206
rect 106007 49985 106235 50217
rect 107791 49982 108019 50214
rect 109576 49980 109804 50212
rect 96364 49432 97874 49834
rect 65284 48532 65560 48632
rect 67154 48584 67390 48662
rect 68959 48576 69193 48655
rect 70765 48570 70984 48651
rect 72551 48571 72791 48655
rect 74352 48586 74604 48651
rect 99808 48538 100084 48638
rect 101678 48590 101914 48668
rect 103483 48582 103717 48661
rect 105289 48576 105508 48657
rect 107075 48577 107315 48661
rect 108876 48592 109128 48657
rect 90796 46782 91108 47320
rect 94987 47083 96094 47300
rect 89567 43153 89693 43279
rect 84505 42267 84628 42609
rect 86529 42262 86618 42646
rect 88515 41630 88641 41756
rect 96525 41606 96795 42681
rect 97372 41603 97642 42678
rect 97972 41682 98218 42396
rect 78109 41343 78235 41469
rect 85883 41236 86119 41241
rect 85883 41010 85888 41236
rect 85888 41010 86114 41236
rect 86114 41010 86119 41236
rect 85883 41005 86119 41010
rect 87808 41218 88019 41223
rect 87808 41017 87813 41218
rect 87813 41017 88014 41218
rect 88014 41017 88019 41218
rect 87808 41012 88019 41017
rect 79904 40461 79983 40739
rect 81965 40420 82045 40703
rect 79094 39823 79220 39949
rect 81162 39699 81290 39704
rect 81162 39581 81167 39699
rect 81167 39581 81285 39699
rect 81285 39581 81290 39699
rect 81162 39576 81290 39581
rect 83018 39595 83142 39719
rect 90783 38091 91030 38958
rect 114709 38737 115008 39378
rect 65328 37035 65572 37235
rect 66930 37046 67174 37246
rect 68833 37106 69077 37306
rect 70550 37090 70794 37290
rect 72364 37085 72608 37285
rect 74336 37079 74580 37279
rect 99844 37028 100088 37228
rect 101446 37039 101690 37239
rect 103349 37099 103593 37299
rect 105066 37083 105310 37283
rect 106880 37078 107124 37278
rect 108852 37072 109096 37272
rect 123011 37052 123095 38345
rect 65850 35656 66234 35734
rect 67641 35667 68041 35741
rect 69447 35667 69835 35741
rect 96849 35740 97596 35851
rect 71244 35632 71632 35706
rect 73046 35628 73433 35706
rect 74840 35625 75235 35702
rect 83780 34890 83918 34895
rect 83780 34762 83785 34890
rect 83785 34762 83913 34890
rect 83913 34762 83918 34890
rect 83780 34757 83918 34762
rect 100366 35649 100750 35727
rect 102157 35660 102557 35734
rect 103963 35660 104351 35734
rect 105760 35625 106148 35699
rect 107562 35621 107949 35699
rect 109356 35618 109751 35695
rect 123011 35592 123095 36885
rect 91354 35332 91558 35536
rect 94542 35332 94746 35536
rect 86368 35325 86506 35330
rect 86368 35197 86373 35325
rect 86373 35197 86501 35325
rect 86501 35197 86506 35325
rect 86368 35192 86506 35197
rect 82232 31330 82348 31334
rect 82232 31222 82236 31330
rect 82236 31222 82344 31330
rect 82344 31222 82348 31330
rect 82232 31218 82348 31222
rect 85795 31831 85911 31835
rect 85795 31723 85799 31831
rect 85799 31723 85907 31831
rect 85907 31723 85911 31831
rect 85795 31719 85911 31723
rect 123012 34387 123095 35405
rect 91312 34179 91516 34383
rect 95265 34379 95470 34383
rect 95265 34183 95270 34379
rect 95270 34183 95466 34379
rect 95466 34183 95470 34379
rect 95265 34179 95470 34183
rect 119413 33914 119539 34040
rect 125028 33811 125348 34131
rect 127217 33666 127594 33739
rect 123010 32643 123097 33617
rect 127219 32552 127591 32617
rect 95427 30789 95711 31246
rect 90814 30288 91056 30752
rect 114716 30726 115015 31367
rect 123007 31104 123097 32470
rect 123008 29606 123099 30864
rect 124329 30866 124649 31186
rect 59363 28460 61033 28687
rect 95203 28464 95762 28684
rect 104388 27172 104516 27177
rect 104388 27054 104393 27172
rect 104393 27054 104511 27172
rect 104511 27054 104516 27172
rect 104388 27049 104516 27054
rect 107961 27185 108079 27190
rect 107961 27067 108074 27185
rect 108074 27067 108079 27185
rect 107961 27062 108079 27067
rect 86377 24870 86495 24988
rect 85207 24727 85281 24732
rect 85207 24663 85212 24727
rect 85212 24663 85276 24727
rect 85276 24663 85281 24727
rect 85207 24658 85281 24663
rect 41228 23742 41356 23870
rect 51068 23721 51186 23839
rect 62988 23722 63106 23840
rect 71557 23719 71675 23837
rect 87014 23902 87088 23907
rect 87014 23838 87019 23902
rect 87019 23838 87083 23902
rect 87083 23838 87088 23902
rect 87014 23833 87088 23838
rect 83055 23654 83173 23772
rect 41701 23526 41765 23590
rect 52551 23516 52615 23580
rect 64440 23583 64514 23588
rect 64440 23519 64445 23583
rect 64445 23519 64509 23583
rect 64509 23519 64514 23583
rect 64440 23514 64514 23519
rect 85591 23604 85709 23722
rect 92590 23670 92708 23788
rect 72870 23587 72944 23592
rect 72870 23523 72875 23587
rect 72875 23523 72939 23587
rect 72939 23523 72944 23587
rect 72870 23518 72944 23523
rect 81872 23538 81946 23543
rect 81872 23474 81877 23538
rect 81877 23474 81941 23538
rect 81941 23474 81946 23538
rect 81872 23469 81946 23474
rect 93131 23537 93205 23542
rect 93131 23473 93136 23537
rect 93136 23473 93200 23537
rect 93200 23473 93205 23537
rect 93131 23468 93205 23473
rect 106372 23300 106500 23428
rect 103434 22990 103552 23108
rect 105417 23160 105491 23165
rect 105417 23096 105422 23160
rect 105422 23096 105486 23160
rect 105486 23096 105491 23160
rect 105417 23091 105491 23096
rect 109004 22995 109122 23113
rect 39914 22711 39978 22775
rect 50506 22704 50570 22768
rect 62415 22760 62489 22765
rect 62415 22696 62420 22760
rect 62420 22696 62484 22760
rect 62484 22696 62489 22760
rect 62415 22691 62489 22696
rect 71181 22761 71255 22766
rect 71181 22697 71186 22761
rect 71186 22697 71250 22761
rect 71250 22697 71255 22761
rect 71181 22692 71255 22697
rect 83454 22711 83528 22716
rect 83454 22647 83459 22711
rect 83459 22647 83523 22711
rect 83523 22647 83528 22711
rect 83454 22642 83528 22647
rect 91387 22712 91461 22717
rect 91387 22648 91392 22712
rect 91392 22648 91456 22712
rect 91456 22648 91461 22712
rect 91387 22643 91461 22648
rect 40383 22450 40511 22578
rect 51940 22469 52058 22587
rect 63860 22464 63978 22582
rect 72435 22460 72553 22578
rect 104394 22670 104510 22674
rect 104394 22562 104398 22670
rect 104398 22562 104506 22670
rect 104506 22562 104510 22670
rect 104394 22558 104510 22562
rect 107980 22689 108096 22693
rect 107980 22581 107984 22689
rect 107984 22581 108092 22689
rect 108092 22581 108096 22689
rect 107980 22577 108096 22581
rect 82256 22404 82374 22522
rect 91882 22410 92000 22528
rect 107090 22350 107174 22355
rect 107090 22276 107095 22350
rect 107095 22276 107169 22350
rect 107169 22276 107174 22350
rect 107090 22271 107174 22276
rect 105796 22028 105924 22156
rect 36843 21755 36971 21883
rect 47795 21719 47923 21847
rect 60239 21753 60357 21871
rect 38303 21586 38377 21591
rect 38303 21522 38308 21586
rect 38308 21522 38372 21586
rect 38372 21522 38377 21586
rect 38303 21517 38377 21522
rect 43434 21534 43562 21662
rect 49362 21519 49426 21583
rect 61659 21584 61733 21589
rect 61659 21520 61664 21584
rect 61664 21520 61728 21584
rect 61728 21520 61733 21584
rect 61659 21515 61733 21520
rect 44837 21339 44901 21403
rect 36278 20709 36342 20773
rect 47042 20703 47106 20767
rect 59693 20763 59767 20768
rect 59693 20699 59698 20763
rect 59698 20699 59762 20763
rect 59762 20699 59767 20763
rect 59693 20694 59767 20699
rect 67161 20731 67225 20795
rect 67989 20728 68053 20792
rect 37638 20451 37766 20579
rect 43010 20518 43074 20582
rect 48603 20449 48731 20577
rect 61061 20461 61179 20579
rect 74028 20481 74092 20545
rect 74856 20487 74920 20551
rect 44260 20269 44388 20397
rect 66649 20214 66767 20332
rect 68386 20206 68504 20324
rect 73565 19952 73683 20070
rect 75276 19975 75394 20093
rect 36843 19757 36971 19885
rect 47791 19714 47919 19842
rect 60241 19723 60359 19841
rect 67163 19761 67227 19825
rect 67985 19762 68049 19826
rect 38307 19528 38371 19592
rect 43415 19526 43543 19654
rect 49357 19518 49421 19582
rect 61662 19581 61736 19586
rect 61662 19517 61667 19581
rect 61667 19517 61731 19581
rect 61731 19517 61736 19581
rect 61662 19512 61736 19517
rect 74034 19519 74098 19583
rect 74860 19518 74924 19582
rect 44840 19339 44904 19403
rect 36280 18707 36344 18771
rect 47040 18697 47104 18761
rect 59710 18700 59774 18764
rect 37633 18450 37761 18578
rect 43010 18518 43074 18582
rect 48603 18450 48731 18578
rect 61055 18465 61173 18583
rect 44259 18261 44387 18389
rect 40397 17738 40525 17866
rect 51104 17722 51222 17840
rect 63015 17715 63133 17833
rect 71584 17726 71702 17844
rect 82968 17695 83086 17813
rect 92566 17701 92684 17819
rect 41702 17523 41766 17587
rect 52547 17516 52611 17580
rect 64442 17518 64506 17582
rect 72877 17594 72951 17599
rect 72877 17530 72882 17594
rect 72882 17530 72946 17594
rect 72946 17530 72951 17594
rect 72877 17525 72951 17530
rect 81877 17567 81951 17572
rect 81877 17503 81882 17567
rect 81882 17503 81946 17567
rect 81946 17503 81951 17567
rect 81877 17498 81951 17503
rect 93134 17503 93198 17567
rect 86412 16844 86530 16962
rect 39911 16701 39975 16765
rect 50503 16698 50567 16762
rect 62416 16763 62490 16768
rect 62416 16699 62421 16763
rect 62421 16699 62485 16763
rect 62485 16699 62490 16763
rect 62416 16694 62490 16699
rect 71185 16774 71259 16779
rect 71185 16710 71190 16774
rect 71190 16710 71254 16774
rect 71254 16710 71259 16774
rect 71185 16705 71259 16710
rect 83450 16747 83524 16752
rect 83450 16683 83455 16747
rect 83455 16683 83519 16747
rect 83519 16683 83524 16747
rect 83450 16678 83524 16683
rect 85205 16717 85279 16722
rect 85205 16653 85210 16717
rect 85210 16653 85274 16717
rect 85274 16653 85279 16717
rect 85205 16648 85279 16653
rect 91397 16743 91471 16748
rect 91397 16679 91402 16743
rect 91402 16679 91466 16743
rect 91466 16679 91471 16743
rect 91397 16674 91471 16679
rect 41211 16414 41339 16542
rect 51817 16464 51935 16582
rect 63827 16455 63945 16573
rect 72296 16464 72414 16582
rect 82296 16443 82414 16561
rect 91859 16429 91977 16547
rect 87011 15892 87085 15897
rect 87011 15828 87016 15892
rect 87016 15828 87080 15892
rect 87080 15828 87085 15892
rect 87011 15823 87085 15828
rect 85624 15577 85742 15695
rect 42983 14405 43111 14533
rect 67124 14405 67252 14533
rect 91367 14405 91495 14533
rect 105384 14405 105512 14533
rect 44812 13863 44940 13991
rect 67969 13863 68097 13991
rect 93107 13863 93235 13991
rect 107068 13863 107196 13991
rect 47010 12222 47138 12350
rect 120735 12222 120863 12350
rect 49330 11680 49458 11808
rect 121333 11680 121461 11808
rect 59672 11136 59800 11264
rect 121937 11136 122065 11264
rect 61642 10597 61770 10725
rect 122541 10597 122669 10725
rect 64415 8956 64543 9084
rect 123737 8956 123865 9084
rect 62392 8420 62520 8548
rect 124335 8420 124463 8548
rect 52517 7870 52645 7998
rect 124939 7870 125067 7998
rect 50477 7334 50605 7462
rect 125537 7334 125665 7462
rect 39882 5693 40010 5821
rect 76521 5685 76645 5809
rect 85178 5693 85306 5821
rect 111040 5679 111158 5797
rect 126739 5693 126867 5821
rect 41670 5156 41798 5284
rect 76910 5146 77032 5268
rect 86989 5156 87117 5284
rect 111439 5157 111555 5273
rect 127339 5156 127467 5284
rect 27434 4611 27562 4739
rect 74000 4600 74126 4726
rect 89566 4611 89694 4739
rect 127933 4611 128061 4739
rect 26623 4063 26751 4191
rect 74813 4063 74941 4191
rect 88514 4063 88642 4191
rect 128545 4063 128673 4191
rect 25661 2435 25789 2563
rect 72846 2435 72974 2563
rect 79093 2435 79221 2563
rect 129748 2435 129876 2563
rect 24761 1889 24889 2017
rect 71156 1889 71284 2017
rect 78108 1889 78236 2017
rect 130331 1889 130459 2017
rect 38277 1338 38405 1466
rect 76122 1333 76248 1459
rect 83425 1338 83553 1466
rect 110635 1338 110755 1458
rect 119412 1338 119540 1466
rect 130936 1338 131064 1466
rect 36248 807 36376 935
rect 75721 793 75847 919
rect 81845 807 81973 935
rect 110236 811 110356 931
rect 131530 807 131658 935
rect 122561 92 122627 158
rect 128558 -166 128624 -100
rect 135402 -36 135875 33
rect 121979 -465 122045 -399
rect 139082 -577 139544 -513
rect 127947 -732 128013 -666
rect 123743 -1225 123809 -1159
rect 129766 -1483 129832 -1417
rect 135405 -1351 135878 -1282
rect 124353 -1782 124419 -1716
rect 139092 -1891 139554 -1827
rect 67103 -2665 67170 -2039
rect 130362 -2049 130428 -1983
rect 121368 -2872 121434 -2806
rect 127364 -3130 127430 -3064
rect 135397 -2997 135870 -2928
rect 120757 -3429 120823 -3363
rect 139082 -3541 139544 -3477
rect 126763 -3696 126829 -3630
rect 124958 -4119 125024 -4053
rect 130963 -4377 131029 -4311
rect 135399 -4247 135872 -4178
rect 125568 -4676 125634 -4610
rect 139097 -4788 139559 -4724
rect 131556 -4943 131622 -4877
rect 66560 -6253 66627 -5627
rect 147329 -11225 147802 -11156
rect 151014 -11769 151476 -11705
rect 71621 -17271 71685 -16617
rect 72709 -17271 72773 -16617
rect 73797 -17271 73861 -16617
rect 74885 -17271 74949 -16617
rect 75973 -17271 76037 -16617
rect 77061 -17271 77125 -16617
rect 78149 -17271 78213 -16617
rect 79237 -17271 79301 -16617
rect 80325 -17271 80389 -16617
rect 81413 -17271 81477 -16617
rect 82501 -17271 82565 -16617
rect 83589 -17271 83653 -16617
rect 84677 -17271 84741 -16617
rect 71075 -22006 71142 -21612
rect 72165 -22012 72232 -21618
rect 73253 -22012 73320 -21618
rect 74341 -22012 74408 -21618
rect 75429 -22012 75496 -21618
rect 76517 -22012 76584 -21618
rect 77605 -22012 77672 -21618
rect 81957 -22012 82024 -21618
rect 83045 -22012 83112 -21618
rect 84133 -22012 84200 -21618
rect 85221 -22012 85288 -21618
<< metal4 >>
rect 9965 86397 11965 91353
rect 9965 74405 11965 84397
rect 9965 66405 11965 73705
rect 9965 58405 11965 65705
rect 9965 50405 11965 57705
rect 9965 42405 11965 49705
rect 9965 34405 11965 41705
rect 9965 26405 11965 33705
rect 9965 18405 11965 25705
rect 9965 10405 11965 17705
rect 9965 2405 11965 9705
rect 9965 -5595 11965 1705
rect 9965 -13595 11965 -6295
rect 9965 -21595 11965 -14295
rect 9965 -34385 11965 -22295
rect 9965 -40917 11965 -36385
rect 13965 82397 15965 91353
rect 155830 82397 157830 91353
rect 15965 80397 15967 82397
rect 13965 71405 15965 80397
rect 155830 71405 157830 80397
rect 38585 70751 38587 70986
rect 13965 63405 15965 70705
rect 35087 70423 35412 70499
rect 35087 67107 35285 70423
rect 35410 67107 35412 70423
rect 35087 66343 35412 67107
rect 38262 70399 38587 70751
rect 59998 70772 59999 71037
rect 38262 67113 38294 70399
rect 38442 67113 38587 70399
rect 38262 67007 38587 67113
rect 42109 70392 42434 70489
rect 45313 70422 45638 70754
rect 42109 67110 42295 70392
rect 42410 67110 42434 70392
rect 42109 66339 42434 67110
rect 45276 70421 45638 70422
rect 45276 67092 45277 70421
rect 45431 67092 45638 70421
rect 45276 67091 45638 67092
rect 45313 67051 45638 67091
rect 56491 70394 56816 70445
rect 59674 70398 59999 70772
rect 67147 70753 67150 70935
rect 56491 70393 56849 70394
rect 56491 67113 56700 70393
rect 56848 67113 56849 70393
rect 56491 67112 56849 67113
rect 59674 67113 59712 70398
rect 59864 67113 59999 70398
rect 42433 65857 42434 66339
rect 56491 66331 56816 67112
rect 59674 66985 59999 67113
rect 63595 70397 63920 70515
rect 63595 70396 63952 70397
rect 66825 70396 67150 70753
rect 88003 70747 88004 70942
rect 63595 67105 63788 70396
rect 63951 67105 63952 70396
rect 66803 70395 67150 70396
rect 66803 67117 66804 70395
rect 66952 67117 67150 70395
rect 66803 67116 67150 67117
rect 63595 67104 63952 67105
rect 63595 66343 63920 67104
rect 66825 66997 67150 67116
rect 73661 70398 73986 70528
rect 73661 67107 73794 70398
rect 73935 67107 73986 70398
rect 76822 70397 77147 70746
rect 76798 70396 77147 70397
rect 76798 67113 76799 70396
rect 76934 67113 77147 70396
rect 76798 67112 77147 67113
rect 56491 66061 56492 66331
rect 73661 66350 73986 67107
rect 76822 67093 77147 67112
rect 84508 70393 84833 70485
rect 87679 70407 88004 70747
rect 84508 67112 84670 70393
rect 84798 67112 84833 70393
rect 63595 65724 63920 65749
rect 63685 65544 63798 65724
rect 63685 65431 67884 65544
rect 63685 65103 63798 65431
rect 65058 65112 65171 65431
rect 66421 65112 66534 65431
rect 67771 65113 67884 65431
rect 68300 65408 68413 65784
rect 84508 66351 84833 67112
rect 87662 70406 88004 70407
rect 87662 67108 87663 70406
rect 87817 67108 88004 70406
rect 87662 67107 88004 67108
rect 87679 67101 88004 67107
rect 92753 70407 93078 70414
rect 92753 70406 93120 70407
rect 68292 65295 68413 65408
rect 67769 65112 67884 65113
rect 63683 65102 63798 65103
rect 62907 65047 63134 65048
rect 62907 64980 62908 65047
rect 63133 64980 63134 65047
rect 63683 64989 63684 65102
rect 63797 64989 63798 65102
rect 65057 65111 65172 65112
rect 64330 65056 64443 65068
rect 63683 64988 63798 64989
rect 62907 64979 63134 64980
rect 62967 63348 63080 64979
rect 13965 55405 15965 62705
rect 62730 62189 62845 62190
rect 62730 62076 62731 62189
rect 62844 62076 62845 62189
rect 62730 62075 62845 62076
rect 62731 61902 62844 62075
rect 62967 61902 63080 62754
rect 63685 62352 63798 64988
rect 64231 65055 64461 65056
rect 64231 64976 64232 65055
rect 64460 64976 64461 65055
rect 65057 64998 65058 65111
rect 65171 64998 65172 65111
rect 66420 65111 66535 65112
rect 65695 65056 65808 65068
rect 65057 64997 65172 64998
rect 65615 65055 65844 65056
rect 64231 64975 64461 64976
rect 63429 62239 63798 62352
rect 63429 62147 63542 62239
rect 64330 62160 64443 64975
rect 65058 62331 65171 64997
rect 65615 64980 65616 65055
rect 65843 64980 65844 65055
rect 66420 64998 66421 65111
rect 66534 64998 66535 65111
rect 67052 65055 67165 65096
rect 66420 64997 66535 64998
rect 66996 65054 67226 65055
rect 65615 64979 65844 64980
rect 64723 62218 65171 62331
rect 64723 62178 64836 62218
rect 64720 62177 64836 62178
rect 64330 62159 64492 62160
rect 63428 62146 63543 62147
rect 63428 62033 63429 62146
rect 63542 62033 63543 62146
rect 63428 62032 63543 62033
rect 64330 62045 64378 62159
rect 64491 62045 64492 62159
rect 64720 62064 64721 62177
rect 64834 62064 64836 62177
rect 64720 62063 64836 62064
rect 64723 62059 64836 62063
rect 65455 62169 65570 62170
rect 65695 62169 65808 64979
rect 66421 62323 66534 64997
rect 66996 64982 66997 65054
rect 67225 64982 67226 65054
rect 67769 64999 67770 65112
rect 67883 64999 67884 65112
rect 67769 64998 67884 64999
rect 66996 64981 67226 64982
rect 65455 62056 65456 62169
rect 65569 62056 65808 62169
rect 66175 62210 66534 62323
rect 66175 62152 66289 62210
rect 65455 62055 65570 62056
rect 64330 62044 64492 62045
rect 64330 61902 64443 62044
rect 65695 61902 65808 62056
rect 66174 62151 66289 62152
rect 66174 62038 66175 62151
rect 66288 62038 66289 62151
rect 66174 62037 66289 62038
rect 66827 62143 66942 62144
rect 67052 62143 67165 64981
rect 67771 62356 67884 64998
rect 67543 62243 67884 62356
rect 67543 62152 67656 62243
rect 66827 62030 66828 62143
rect 66941 62030 67165 62143
rect 67542 62151 67657 62152
rect 67542 62038 67543 62151
rect 67656 62038 67657 62151
rect 67542 62037 67657 62038
rect 66827 62029 66942 62030
rect 67052 61902 67165 62030
rect 62731 61790 67165 61902
rect 62731 61789 63648 61790
rect 63818 61789 67165 61790
rect 68300 61658 68413 65295
rect 73685 65544 73798 65756
rect 92753 67100 92977 70406
rect 93119 67100 93120 70406
rect 92753 67099 93120 67100
rect 95977 70403 96302 70761
rect 95977 67112 95985 70403
rect 96113 67112 96302 70403
rect 92753 66341 93078 67099
rect 95977 67083 96302 67112
rect 102093 70407 102418 70414
rect 102093 70406 102460 70407
rect 102093 67100 102317 70406
rect 102459 67100 102460 70406
rect 102093 67099 102460 67100
rect 105317 70403 105642 70761
rect 105317 67112 105325 70403
rect 105453 67112 105642 70403
rect 73685 65431 77884 65544
rect 73685 65103 73798 65431
rect 75058 65112 75171 65431
rect 76421 65112 76534 65431
rect 77771 65113 77884 65431
rect 77769 65112 77884 65113
rect 73683 65102 73798 65103
rect 72907 65047 73134 65048
rect 72907 64980 72908 65047
rect 73133 64980 73134 65047
rect 73683 64989 73684 65102
rect 73797 64989 73798 65102
rect 75057 65111 75172 65112
rect 74330 65056 74443 65068
rect 73683 64988 73798 64989
rect 72907 64979 73134 64980
rect 72967 63348 73080 64979
rect 72730 62189 72845 62190
rect 72730 62076 72731 62189
rect 72844 62076 72845 62189
rect 72730 62075 72845 62076
rect 72731 61902 72844 62075
rect 72967 61902 73080 62754
rect 73685 62352 73798 64988
rect 74231 65055 74461 65056
rect 74231 64976 74232 65055
rect 74460 64976 74461 65055
rect 75057 64998 75058 65111
rect 75171 64998 75172 65111
rect 76420 65111 76535 65112
rect 75695 65056 75808 65068
rect 75057 64997 75172 64998
rect 75615 65055 75844 65056
rect 74231 64975 74461 64976
rect 73429 62239 73798 62352
rect 73429 62147 73542 62239
rect 74330 62160 74443 64975
rect 75058 62331 75171 64997
rect 75615 64980 75616 65055
rect 75843 64980 75844 65055
rect 76420 64998 76421 65111
rect 76534 64998 76535 65111
rect 77052 65055 77165 65096
rect 76420 64997 76535 64998
rect 76996 65054 77226 65055
rect 75615 64979 75844 64980
rect 74723 62218 75171 62331
rect 74723 62178 74836 62218
rect 74720 62177 74836 62178
rect 74330 62159 74492 62160
rect 73428 62146 73543 62147
rect 73428 62033 73429 62146
rect 73542 62033 73543 62146
rect 73428 62032 73543 62033
rect 74330 62045 74378 62159
rect 74491 62045 74492 62159
rect 74720 62064 74721 62177
rect 74834 62064 74836 62177
rect 74720 62063 74836 62064
rect 74723 62059 74836 62063
rect 75455 62169 75570 62170
rect 75695 62169 75808 64979
rect 76421 62323 76534 64997
rect 76996 64982 76997 65054
rect 77225 64982 77226 65054
rect 77769 64999 77770 65112
rect 77883 64999 77884 65112
rect 77769 64998 77884 64999
rect 76996 64981 77226 64982
rect 75455 62056 75456 62169
rect 75569 62056 75808 62169
rect 76175 62210 76534 62323
rect 76175 62152 76289 62210
rect 75455 62055 75570 62056
rect 74330 62044 74492 62045
rect 74330 61902 74443 62044
rect 75695 61902 75808 62056
rect 76174 62151 76289 62152
rect 76174 62038 76175 62151
rect 76288 62038 76289 62151
rect 76174 62037 76289 62038
rect 76827 62143 76942 62144
rect 77052 62143 77165 64981
rect 77771 62356 77884 64998
rect 77543 62243 77884 62356
rect 77543 62152 77656 62243
rect 76827 62030 76828 62143
rect 76941 62030 77165 62143
rect 77542 62151 77657 62152
rect 77542 62038 77543 62151
rect 77656 62038 77657 62151
rect 77542 62037 77657 62038
rect 76827 62029 76942 62030
rect 77052 61902 77165 62030
rect 72731 61790 77165 61902
rect 72731 61789 73648 61790
rect 73818 61789 77165 61790
rect 78300 61658 78413 65751
rect 85172 64150 86615 64263
rect 85172 63850 85285 64150
rect 86502 63859 86615 64150
rect 86484 63858 86630 63859
rect 85127 63849 85319 63850
rect 85127 63757 85128 63849
rect 85318 63757 85319 63849
rect 85127 63756 85319 63757
rect 85567 63823 86003 63824
rect 85172 63217 85285 63756
rect 85567 63736 85568 63823
rect 86002 63736 86003 63823
rect 86484 63764 86485 63858
rect 86629 63764 86630 63858
rect 87108 63810 87221 65835
rect 102093 66341 102418 67099
rect 105317 67083 105642 67112
rect 102826 64150 104269 64263
rect 102826 63850 102939 64150
rect 104156 63859 104269 64150
rect 104138 63858 104284 63859
rect 102781 63849 102973 63850
rect 86484 63763 86630 63764
rect 86903 63809 87329 63810
rect 85567 63735 86003 63736
rect 85172 62347 85285 62897
rect 85172 62346 85312 62347
rect 85172 62237 85219 62346
rect 85311 62237 85312 62346
rect 85172 62236 85312 62237
rect 85172 62195 85285 62236
rect 62987 61545 68413 61658
rect 72987 61545 78413 61658
rect 63162 61352 63235 61353
rect 63162 61245 63163 61352
rect 63234 61245 63235 61352
rect 63706 61347 63777 61545
rect 63162 61244 63235 61245
rect 63704 61346 63777 61347
rect 63163 60531 63234 61244
rect 63704 61242 63705 61346
rect 63776 61242 63777 61346
rect 63704 61241 63777 61242
rect 63706 61224 63777 61241
rect 64250 61330 64321 61331
rect 64250 61184 64251 61330
rect 64320 61184 64321 61330
rect 64797 61322 64861 61545
rect 65883 61473 65953 61545
rect 65883 61349 65884 61473
rect 65952 61349 65953 61473
rect 66973 61384 67044 61545
rect 66970 61383 67044 61384
rect 65883 61347 65953 61349
rect 66425 61364 66495 61365
rect 64797 61321 64863 61322
rect 64797 61191 64798 61321
rect 64862 61191 64863 61321
rect 66425 61207 66426 61364
rect 66494 61207 66495 61364
rect 66970 61261 66971 61383
rect 67043 61261 67044 61383
rect 66970 61260 67044 61261
rect 67513 61356 67581 61357
rect 66425 61206 66495 61207
rect 64797 61190 64863 61191
rect 64250 61183 64321 61184
rect 64250 60531 64320 61183
rect 65342 61015 65411 61016
rect 65342 60862 65343 61015
rect 65410 60862 65411 61015
rect 65342 60861 65411 60862
rect 65342 60531 65409 60861
rect 66426 60531 66493 61206
rect 67513 61202 67514 61356
rect 67580 61202 67581 61356
rect 73162 61352 73235 61353
rect 73162 61245 73163 61352
rect 73234 61245 73235 61352
rect 73706 61347 73777 61545
rect 73162 61244 73235 61245
rect 73704 61346 73777 61347
rect 67513 61201 67581 61202
rect 67515 60531 67579 61201
rect 73163 60531 73234 61244
rect 73704 61242 73705 61346
rect 73776 61242 73777 61346
rect 73704 61241 73777 61242
rect 73706 61224 73777 61241
rect 74250 61330 74321 61331
rect 74250 61184 74251 61330
rect 74320 61184 74321 61330
rect 74797 61322 74861 61545
rect 75883 61473 75953 61545
rect 75883 61349 75884 61473
rect 75952 61349 75953 61473
rect 76973 61384 77044 61545
rect 76970 61383 77044 61384
rect 75883 61347 75953 61349
rect 76425 61364 76495 61365
rect 74797 61321 74863 61322
rect 74797 61191 74798 61321
rect 74862 61191 74863 61321
rect 76425 61207 76426 61364
rect 76494 61207 76495 61364
rect 76970 61261 76971 61383
rect 77043 61261 77044 61383
rect 76970 61260 77044 61261
rect 77513 61356 77581 61357
rect 76425 61206 76495 61207
rect 74797 61190 74863 61191
rect 74250 61183 74321 61184
rect 74250 60531 74320 61183
rect 75342 61015 75411 61016
rect 75342 60862 75343 61015
rect 75410 60862 75411 61015
rect 75342 60861 75411 60862
rect 75342 60531 75409 60861
rect 76426 60531 76493 61206
rect 77513 61202 77514 61356
rect 77580 61202 77581 61356
rect 77513 61201 77581 61202
rect 77515 60531 77579 61201
rect 85701 60771 85814 63735
rect 86502 63202 86615 63763
rect 86903 63732 86904 63809
rect 87328 63732 87329 63809
rect 102781 63757 102782 63849
rect 102972 63757 102973 63849
rect 102781 63756 102973 63757
rect 103221 63823 103657 63824
rect 86903 63731 87329 63732
rect 86502 62342 86615 62882
rect 86502 62341 86643 62342
rect 86502 62232 86550 62341
rect 86642 62232 86643 62341
rect 86502 62231 86643 62232
rect 86502 62198 86615 62231
rect 87108 60771 87221 63731
rect 102826 63217 102939 63756
rect 103221 63736 103222 63823
rect 103656 63736 103657 63823
rect 104138 63764 104139 63858
rect 104283 63764 104284 63858
rect 104762 63810 104875 65878
rect 104138 63763 104284 63764
rect 104557 63809 104983 63810
rect 103221 63735 103657 63736
rect 102826 62347 102939 62897
rect 102826 62346 102966 62347
rect 102826 62237 102873 62346
rect 102965 62237 102966 62346
rect 102826 62236 102966 62237
rect 102826 62195 102939 62236
rect 85701 60658 87221 60771
rect 103355 60771 103468 63735
rect 104156 63202 104269 63763
rect 104557 63732 104558 63809
rect 104982 63732 104983 63809
rect 104557 63731 104983 63732
rect 104156 62342 104269 62882
rect 104156 62341 104297 62342
rect 104156 62232 104204 62341
rect 104296 62232 104297 62341
rect 104156 62231 104297 62232
rect 104156 62198 104269 62231
rect 104762 60771 104875 63731
rect 103355 60658 104875 60771
rect 155830 63405 157830 70705
rect 62731 60418 67873 60531
rect 72746 60418 77873 60531
rect 86094 60500 86159 60658
rect 103748 60500 103813 60658
rect 63052 59994 63165 60034
rect 63051 59993 63306 59994
rect 63051 59916 63052 59993
rect 63305 59916 63306 59993
rect 63051 59915 63306 59916
rect 63052 58626 63165 59915
rect 63937 59352 64050 60418
rect 64371 60000 64681 60001
rect 64371 59915 64372 60000
rect 64680 59915 64681 60000
rect 64371 59914 64681 59915
rect 63936 59351 64051 59352
rect 63936 59238 63937 59351
rect 64050 59238 64051 59351
rect 63936 59237 64051 59238
rect 64507 58626 64620 59914
rect 65298 59364 65411 60418
rect 65863 59990 65976 60021
rect 65759 59989 66043 59990
rect 65759 59918 65760 59989
rect 66042 59918 66043 59989
rect 65759 59917 66043 59918
rect 65297 59363 65412 59364
rect 65297 59250 65298 59363
rect 65411 59250 65412 59363
rect 65297 59249 65412 59250
rect 65863 58626 65976 59917
rect 66660 59382 66773 60418
rect 67131 59991 67415 59992
rect 67131 59920 67132 59991
rect 67414 59920 67415 59991
rect 67131 59919 67415 59920
rect 66659 59381 66774 59382
rect 66659 59268 66660 59381
rect 66773 59268 66774 59381
rect 66659 59267 66774 59268
rect 67226 58626 67339 59919
rect 63052 58513 67339 58626
rect 67760 59416 67873 60418
rect 73052 59994 73165 60034
rect 73051 59993 73306 59994
rect 73051 59916 73052 59993
rect 73305 59916 73306 59993
rect 73051 59915 73306 59916
rect 68043 59416 68158 59417
rect 67760 59303 68044 59416
rect 68157 59303 68158 59416
rect 63052 58201 63165 58513
rect 67760 55213 67873 59303
rect 68043 59302 68158 59303
rect 73052 58626 73165 59915
rect 73937 59352 74050 60418
rect 74371 60000 74681 60001
rect 74371 59915 74372 60000
rect 74680 59915 74681 60000
rect 74371 59914 74681 59915
rect 73936 59351 74051 59352
rect 73936 59238 73937 59351
rect 74050 59238 74051 59351
rect 73936 59237 74051 59238
rect 74507 58626 74620 59914
rect 75298 59364 75411 60418
rect 75863 59990 75976 60021
rect 75759 59989 76043 59990
rect 75759 59918 75760 59989
rect 76042 59918 76043 59989
rect 75759 59917 76043 59918
rect 75297 59363 75412 59364
rect 75297 59250 75298 59363
rect 75411 59250 75412 59363
rect 75297 59249 75412 59250
rect 75863 58626 75976 59917
rect 76660 59382 76773 60418
rect 77131 59991 77415 59992
rect 77131 59920 77132 59991
rect 77414 59920 77415 59991
rect 77131 59919 77415 59920
rect 76659 59381 76774 59382
rect 76659 59268 76660 59381
rect 76773 59268 76774 59381
rect 76659 59267 76774 59268
rect 77226 58626 77339 59919
rect 73052 58513 77339 58626
rect 77760 59416 77873 60418
rect 86093 60499 86160 60500
rect 86093 60357 86094 60499
rect 86159 60357 86160 60499
rect 86093 60356 86160 60357
rect 103747 60499 103814 60500
rect 103747 60357 103748 60499
rect 103813 60357 103814 60499
rect 103747 60356 103814 60357
rect 86094 60344 86159 60356
rect 103748 60344 103813 60356
rect 86634 60281 86703 60283
rect 104288 60281 104357 60283
rect 86634 60280 86705 60281
rect 85543 60274 85616 60275
rect 85543 60170 85544 60274
rect 85615 60265 85616 60274
rect 85615 60170 85617 60265
rect 85543 60169 85617 60170
rect 85544 60022 85617 60169
rect 86634 60170 86636 60280
rect 86704 60170 86705 60280
rect 104288 60280 104359 60281
rect 86634 60169 86705 60170
rect 103197 60274 103270 60275
rect 103197 60170 103198 60274
rect 103269 60265 103270 60274
rect 103269 60170 103271 60265
rect 103197 60169 103271 60170
rect 86634 60022 86703 60169
rect 103198 60022 103271 60169
rect 104288 60170 104290 60280
rect 104358 60170 104359 60280
rect 104288 60169 104359 60170
rect 104288 60022 104357 60169
rect 84943 59909 87406 60022
rect 84943 59637 85056 59909
rect 84942 59636 85057 59637
rect 84942 59523 84943 59636
rect 85056 59523 85057 59636
rect 84942 59522 85057 59523
rect 78043 59416 78158 59417
rect 77760 59303 78044 59416
rect 78157 59303 78158 59416
rect 73052 58201 73165 58513
rect 77760 55217 77873 59303
rect 78043 59302 78158 59303
rect 85634 58267 85747 59687
rect 86488 58267 86601 59683
rect 85634 58218 86601 58267
rect 85851 58154 86601 58218
rect 87293 59031 87406 59909
rect 102597 59909 105060 60022
rect 102597 59637 102710 59909
rect 102596 59636 102711 59637
rect 102596 59523 102597 59636
rect 102710 59523 102711 59636
rect 102596 59522 102711 59523
rect 87293 59030 87450 59031
rect 87293 58917 87336 59030
rect 87449 58917 87450 59030
rect 87293 58916 87450 58917
rect 13965 47405 15965 54705
rect 27434 52668 27562 52669
rect 27434 52542 27435 52668
rect 27561 52542 27562 52668
rect 13965 39405 15965 46705
rect 13965 31405 15965 38705
rect 13965 23405 15965 30705
rect 13965 15405 15965 22705
rect 13965 7405 15965 14705
rect 13965 -595 15965 6705
rect 24761 50634 24889 50635
rect 24761 50508 24762 50634
rect 24888 50508 24889 50634
rect 24761 2018 24889 50508
rect 25661 49057 25789 49058
rect 25661 48931 25662 49057
rect 25788 48931 25789 49057
rect 25661 2564 25789 48931
rect 26623 48329 26751 48330
rect 26623 48203 26624 48329
rect 26750 48203 26751 48329
rect 26623 4192 26751 48203
rect 27434 4740 27562 52542
rect 46108 52283 46268 54901
rect 46108 52282 46272 52283
rect 46108 51695 46153 52282
rect 46271 51695 46272 52282
rect 48152 52230 48312 54909
rect 87293 55196 87406 58916
rect 103288 58267 103401 59687
rect 104142 58267 104255 59683
rect 103288 58218 104255 58267
rect 103505 58154 104255 58218
rect 104947 59031 105060 59909
rect 104947 59030 105104 59031
rect 104947 58917 104990 59030
rect 105103 58917 105104 59030
rect 104947 58916 105104 58917
rect 104947 55228 105060 58916
rect 155830 55405 157830 62705
rect 115496 52795 115624 54900
rect 119940 54635 120210 54888
rect 119215 54365 120931 54635
rect 46108 51694 46272 51695
rect 47476 51852 47636 51866
rect 46108 51693 46268 51694
rect 47476 51229 47493 51852
rect 47608 51229 47636 51852
rect 48152 51690 48197 52230
rect 48307 51690 48312 52230
rect 115204 52667 116866 52795
rect 49510 51907 49655 51908
rect 49510 51903 49511 51907
rect 48152 51683 48312 51690
rect 45802 50922 45930 50923
rect 45802 50796 45803 50922
rect 45929 50796 45930 50922
rect 35850 49931 36152 49935
rect 35850 49927 36290 49931
rect 35850 49483 36202 49927
rect 36285 49483 36290 49927
rect 37951 49857 38253 49894
rect 35850 49473 36290 49483
rect 35850 47283 36152 49473
rect 37951 49278 38144 49857
rect 38243 49278 38253 49857
rect 37951 47223 38253 49278
rect 45802 48331 45930 50796
rect 47476 50200 47636 51229
rect 49507 51249 49511 51903
rect 49654 51903 49655 51907
rect 49654 51249 49667 51903
rect 49507 50169 49667 51249
rect 115204 51726 115332 52667
rect 116738 52515 116866 52667
rect 116737 52514 116867 52515
rect 116737 52386 116738 52514
rect 116866 52386 116867 52514
rect 116737 52385 116867 52386
rect 116738 52345 116866 52385
rect 119215 52130 119485 54365
rect 120661 52468 120931 54365
rect 120661 52467 120934 52468
rect 120661 52363 120662 52467
rect 120933 52363 120934 52467
rect 120661 52362 120934 52363
rect 120661 52185 120931 52362
rect 117728 51778 117833 51779
rect 115204 51725 115386 51726
rect 115204 51273 115289 51725
rect 115385 51273 115386 51725
rect 117728 51316 117729 51778
rect 117832 51612 117833 51778
rect 117832 51316 117950 51612
rect 117728 51315 117950 51316
rect 115204 51272 115386 51273
rect 115204 50703 115332 51272
rect 117395 50953 117554 50954
rect 115578 50928 115708 50929
rect 115578 50800 115579 50928
rect 115707 50800 115708 50928
rect 117395 50869 117396 50953
rect 117553 50869 117554 50953
rect 117395 50868 117554 50869
rect 116124 50862 116204 50864
rect 115578 50799 115708 50800
rect 115988 50861 116204 50862
rect 115579 50703 115707 50799
rect 115988 50709 115989 50861
rect 116141 50709 116204 50861
rect 115988 50708 116204 50709
rect 115204 50575 115707 50703
rect 115989 50700 116204 50708
rect 117398 50700 117550 50868
rect 117798 50700 117950 51315
rect 119215 51001 119326 52130
rect 119407 51001 119485 52130
rect 121708 52123 121805 52124
rect 121708 51731 121709 52123
rect 121653 51411 121709 51731
rect 121708 51027 121709 51411
rect 121804 51731 121805 52123
rect 121804 51411 122409 51731
rect 121804 51027 121805 51411
rect 121708 51026 121805 51027
rect 119215 50968 119485 51001
rect 115989 50548 117950 50700
rect 119718 50944 120241 51000
rect 119718 50772 119936 50944
rect 120225 50772 120241 50944
rect 119718 50680 120241 50772
rect 121195 50958 121517 50959
rect 121195 50888 121196 50958
rect 121516 50888 121517 50958
rect 121195 50887 121517 50888
rect 63349 49801 63357 50255
rect 62822 49623 63357 49801
rect 62822 49622 63381 49623
rect 62822 49465 62848 49622
rect 63380 49465 63381 49622
rect 62822 49464 63381 49465
rect 62822 49450 63357 49464
rect 67147 48662 67404 48678
rect 65246 48632 65588 48650
rect 65246 48532 65284 48632
rect 65560 48532 65588 48632
rect 65246 48450 65588 48532
rect 67147 48584 67154 48662
rect 67390 48584 67404 48662
rect 67147 48450 67404 48584
rect 68945 48655 69202 48663
rect 68945 48576 68959 48655
rect 69193 48576 69202 48655
rect 68945 48450 69202 48576
rect 70741 48651 70996 48659
rect 70741 48570 70765 48651
rect 70984 48570 70996 48651
rect 70741 48450 70996 48570
rect 72544 48655 72799 48662
rect 72544 48571 72551 48655
rect 72791 48571 72799 48655
rect 72544 48450 72799 48571
rect 74331 48651 74622 48652
rect 74331 48586 74352 48651
rect 74604 48586 74622 48651
rect 74331 48450 74622 48586
rect 45801 48330 45931 48331
rect 45801 48202 45802 48330
rect 45930 48202 45931 48330
rect 45801 48201 45931 48202
rect 64066 48130 75300 48450
rect 56045 47379 56331 47380
rect 56045 46741 56046 47379
rect 56330 46741 56331 47379
rect 64066 47220 64386 48130
rect 95481 47377 95601 50324
rect 117398 50228 117550 50548
rect 119718 50212 120038 50680
rect 120037 49921 120038 50212
rect 96363 49432 96364 49764
rect 97874 49432 97875 49764
rect 96363 49431 97875 49432
rect 101671 48668 101928 48684
rect 99770 48638 100112 48656
rect 99770 48538 99808 48638
rect 100084 48538 100112 48638
rect 99770 48456 100112 48538
rect 101671 48590 101678 48668
rect 101914 48590 101928 48668
rect 101671 48456 101928 48590
rect 103469 48661 103726 48669
rect 103469 48582 103483 48661
rect 103717 48582 103726 48661
rect 103469 48456 103726 48582
rect 105265 48657 105520 48665
rect 105265 48576 105289 48657
rect 105508 48576 105520 48657
rect 105265 48456 105520 48576
rect 107068 48661 107323 48668
rect 107068 48577 107075 48661
rect 107315 48577 107323 48661
rect 107068 48456 107323 48577
rect 108855 48657 109146 48658
rect 108855 48592 108876 48657
rect 109128 48592 109146 48657
rect 108855 48456 109146 48592
rect 98590 48136 109824 48456
rect 90872 47321 90992 47358
rect 64384 47078 64386 47220
rect 90795 47320 91109 47321
rect 90795 46782 90796 47320
rect 91108 46782 91109 47320
rect 98590 47226 98910 48136
rect 98908 47084 98910 47226
rect 121195 47216 121515 50887
rect 122089 50227 122409 51411
rect 122089 50022 122091 50227
rect 121514 47189 121515 47216
rect 155830 47405 157830 54705
rect 90795 46781 91109 46782
rect 56045 46740 56331 46741
rect 89566 43279 89694 43280
rect 89566 43153 89567 43279
rect 89693 43153 89694 43279
rect 43141 42670 44785 42734
rect 46323 42666 47956 42730
rect 61879 42674 63777 42709
rect 33426 42574 38481 42638
rect 61879 42335 62010 42674
rect 62280 42671 63777 42674
rect 62280 42335 62857 42671
rect 63127 42335 63777 42671
rect 86528 42646 86619 42647
rect 84504 42609 84629 42610
rect 84504 42520 84505 42609
rect 61879 41731 61951 42335
rect 63172 41747 63412 42335
rect 63617 41747 63777 42335
rect 84216 42377 84505 42520
rect 84216 42237 84359 42377
rect 84504 42267 84505 42377
rect 84628 42267 84629 42609
rect 86528 42511 86529 42646
rect 84504 42266 84629 42267
rect 86349 42262 86529 42511
rect 86618 42511 86619 42646
rect 86618 42368 86625 42511
rect 86618 42262 86623 42368
rect 86349 42229 86623 42262
rect 86590 41944 86623 42229
rect 63172 41731 63777 41747
rect 61879 41599 62010 41731
rect 62280 41599 62857 41731
rect 61879 41596 62857 41599
rect 63127 41596 63777 41731
rect 61879 41565 63777 41596
rect 78108 41469 78236 41470
rect 32097 33415 32161 41442
rect 36687 40610 36827 40611
rect 36687 40472 36688 40610
rect 36826 40472 36827 40610
rect 36687 40471 36827 40472
rect 36693 39678 36821 40471
rect 39642 39823 39706 41431
rect 41824 39823 41888 41341
rect 44959 40533 45099 40534
rect 44959 40395 44960 40533
rect 45098 40395 45099 40533
rect 44959 40394 45099 40395
rect 44965 39609 45093 40394
rect 49369 39435 49433 41349
rect 78108 41343 78109 41469
rect 78235 41343 78236 41469
rect 56026 39355 56168 39356
rect 35459 36623 35523 38141
rect 39642 36623 39706 38141
rect 41824 36623 41888 38141
rect 46007 36623 46071 38141
rect 49369 35888 49433 38966
rect 56026 38731 56027 39355
rect 56167 39337 56168 39355
rect 56167 38731 56168 38752
rect 56026 38730 56168 38731
rect 64123 37306 75204 37559
rect 64123 37246 68833 37306
rect 64123 37239 66930 37246
rect 49315 35813 49570 35888
rect 49315 35682 49606 35813
rect 49369 35607 49606 35682
rect 39642 33423 39706 34941
rect 41824 33333 41888 34941
rect 49369 33322 49433 35607
rect 50242 32672 50362 32673
rect 50242 32667 50243 32672
rect 40665 32648 40785 32649
rect 40665 32643 40666 32648
rect 39809 32525 40666 32643
rect 40665 32520 40666 32525
rect 40784 32520 40785 32648
rect 49436 32549 50243 32667
rect 50242 32544 50243 32549
rect 50361 32544 50362 32672
rect 50242 32543 50362 32544
rect 40665 32519 40785 32520
rect 43049 32126 48104 32190
rect 33529 32030 38556 32098
rect 55951 31354 56300 31355
rect 55951 30754 55952 31354
rect 56299 30754 56300 31354
rect 55951 30753 56300 30754
rect 64123 31125 64374 37239
rect 65294 37235 65614 37239
rect 65294 37035 65328 37235
rect 65572 37035 65614 37235
rect 66929 37046 66930 37239
rect 67174 37239 68833 37246
rect 67174 37046 67175 37239
rect 68832 37106 68833 37239
rect 69077 37290 75204 37306
rect 69077 37239 70550 37290
rect 69077 37106 69078 37239
rect 68832 37105 69078 37106
rect 70549 37090 70550 37239
rect 70794 37285 75204 37290
rect 70794 37239 72364 37285
rect 70794 37090 70795 37239
rect 70549 37089 70795 37090
rect 72363 37085 72364 37239
rect 72608 37279 75204 37285
rect 72608 37239 74336 37279
rect 72608 37085 72609 37239
rect 72363 37084 72609 37085
rect 74335 37079 74336 37239
rect 74580 37239 75204 37279
rect 74580 37079 74581 37239
rect 74335 37078 74581 37079
rect 66929 37045 67175 37046
rect 65294 37028 65614 37035
rect 67642 35742 68044 35743
rect 67640 35741 68044 35742
rect 65840 35734 66241 35740
rect 65840 35656 65850 35734
rect 66234 35656 66241 35734
rect 67640 35667 67641 35741
rect 68041 35667 68044 35741
rect 67640 35666 68044 35667
rect 69446 35741 69836 35742
rect 69446 35667 69447 35741
rect 69835 35667 69836 35741
rect 69446 35666 69836 35667
rect 71243 35706 71633 35707
rect 65840 35546 66241 35656
rect 67642 35546 68044 35666
rect 69513 35546 69781 35666
rect 71243 35632 71244 35706
rect 71632 35632 71633 35706
rect 71243 35631 71633 35632
rect 73044 35706 73435 35711
rect 71244 35546 71632 35631
rect 73044 35628 73046 35706
rect 73433 35628 73435 35706
rect 73044 35546 73435 35628
rect 74836 35702 75237 35705
rect 74836 35625 74840 35702
rect 75235 35625 75237 35702
rect 74836 35546 75237 35625
rect 65176 35226 75256 35546
rect 70278 34224 70598 35226
rect 60380 30104 60700 30856
rect 60985 30188 61192 30189
rect 60985 30104 60986 30188
rect 60380 29784 60986 30104
rect 60380 28688 60700 29784
rect 60985 29648 60986 29784
rect 61191 30104 61192 30188
rect 61191 29784 61197 30104
rect 61191 29648 61192 29784
rect 60985 29647 61192 29648
rect 59362 28687 61034 28688
rect 59362 28460 59363 28687
rect 61033 28460 61034 28687
rect 59362 28459 61034 28460
rect 41220 23871 41348 25829
rect 41220 23870 41357 23871
rect 41220 23755 41228 23870
rect 41227 23742 41228 23755
rect 41356 23742 41357 23870
rect 51066 23840 51184 25870
rect 62990 23841 63108 25942
rect 62987 23840 63108 23841
rect 51066 23839 51187 23840
rect 51066 23796 51068 23839
rect 41227 23741 41357 23742
rect 51067 23721 51068 23796
rect 51186 23721 51187 23839
rect 62987 23722 62988 23840
rect 63106 23767 63108 23840
rect 71554 23838 71672 25841
rect 71554 23837 71676 23838
rect 71554 23786 71557 23837
rect 63106 23722 63107 23767
rect 62987 23721 63107 23722
rect 51067 23720 51187 23721
rect 71556 23719 71557 23786
rect 71675 23719 71676 23837
rect 71556 23718 71676 23719
rect 41670 23590 41798 23634
rect 41670 23526 41701 23590
rect 41765 23526 41798 23590
rect 36826 21884 36954 21921
rect 36826 21883 36972 21884
rect 36826 21755 36843 21883
rect 36971 21755 36972 21883
rect 36826 21754 36972 21755
rect 36248 20773 36376 20804
rect 36248 20709 36278 20773
rect 36342 20709 36376 20773
rect 36248 18771 36376 20709
rect 36248 18707 36280 18771
rect 36344 18707 36376 18771
rect 27433 4739 27563 4740
rect 27433 4611 27434 4739
rect 27562 4611 27563 4739
rect 27433 4610 27563 4611
rect 26622 4191 26752 4192
rect 26622 4063 26623 4191
rect 26751 4063 26752 4191
rect 26622 4062 26752 4063
rect 25660 2563 25790 2564
rect 25660 2435 25661 2563
rect 25789 2435 25790 2563
rect 25660 2434 25790 2435
rect 24760 2017 24890 2018
rect 24760 1889 24761 2017
rect 24889 1889 24890 2017
rect 24760 1888 24890 1889
rect 36248 936 36376 18707
rect 36826 19886 36954 21754
rect 37633 20580 37761 22884
rect 39882 22775 40010 22802
rect 39882 22711 39914 22775
rect 39978 22711 40010 22775
rect 38277 21591 38405 21615
rect 38277 21517 38303 21591
rect 38377 21517 38405 21591
rect 37633 20579 37767 20580
rect 37633 20451 37638 20579
rect 37766 20451 37767 20579
rect 37633 20450 37767 20451
rect 36826 19885 36972 19886
rect 36826 19757 36843 19885
rect 36971 19757 36972 19885
rect 36826 19756 36972 19757
rect 36826 18194 36954 19756
rect 37633 18579 37761 20450
rect 38277 19592 38405 21517
rect 38277 19528 38307 19592
rect 38371 19528 38405 19592
rect 37632 18578 37762 18579
rect 37632 18450 37633 18578
rect 37761 18450 37762 18578
rect 37632 18449 37762 18450
rect 37633 18425 37761 18449
rect 38277 1467 38405 19528
rect 39882 16765 40010 22711
rect 40392 22579 40520 22881
rect 40382 22578 40520 22579
rect 40382 22450 40383 22578
rect 40511 22455 40520 22578
rect 40511 22450 40512 22455
rect 40382 22449 40512 22450
rect 40292 18197 40633 18243
rect 40292 17877 40301 18197
rect 40621 17877 40633 18197
rect 40292 17866 40633 17877
rect 40292 17835 40397 17866
rect 40396 17738 40397 17835
rect 40525 17835 40633 17866
rect 40525 17738 40526 17835
rect 40396 17737 40526 17738
rect 39882 16701 39911 16765
rect 39975 16701 40010 16765
rect 39882 5822 40010 16701
rect 41670 17587 41798 23526
rect 52517 23580 52645 23641
rect 52517 23516 52551 23580
rect 52615 23516 52645 23580
rect 43431 21663 43559 22933
rect 50477 22768 50605 22798
rect 50477 22704 50506 22768
rect 50570 22704 50605 22768
rect 47795 21848 47923 21888
rect 47794 21847 47924 21848
rect 47794 21719 47795 21847
rect 47923 21719 47924 21847
rect 47794 21718 47924 21719
rect 43431 21662 43563 21663
rect 43431 21534 43434 21662
rect 43562 21534 43563 21662
rect 43431 21533 43563 21534
rect 41670 17523 41702 17587
rect 41766 17523 41798 17587
rect 41211 16543 41339 16550
rect 41210 16542 41340 16543
rect 41210 16414 41211 16542
rect 41339 16414 41340 16542
rect 41210 16413 41340 16414
rect 41211 15209 41339 16413
rect 39881 5821 40011 5822
rect 39881 5693 39882 5821
rect 40010 5693 40011 5821
rect 39881 5692 40011 5693
rect 41670 5285 41798 17523
rect 42983 20582 43111 20631
rect 42983 20518 43010 20582
rect 43074 20518 43111 20582
rect 42983 18582 43111 20518
rect 43431 19655 43559 21533
rect 44812 21403 44940 21433
rect 44812 21339 44837 21403
rect 44901 21339 44940 21403
rect 44259 20397 44389 20398
rect 44259 20269 44260 20397
rect 44388 20269 44389 20397
rect 44259 20268 44389 20269
rect 43414 19654 43559 19655
rect 43414 19526 43415 19654
rect 43543 19544 43559 19654
rect 43543 19526 43544 19544
rect 43414 19525 43544 19526
rect 42983 18518 43010 18582
rect 43074 18518 43111 18582
rect 42983 14534 43111 18518
rect 44261 18390 44389 20268
rect 44258 18389 44389 18390
rect 44258 18344 44259 18389
rect 44166 18261 44259 18344
rect 44387 18344 44389 18389
rect 44812 19403 44940 21339
rect 44812 19339 44840 19403
rect 44904 19339 44940 19403
rect 44387 18261 44486 18344
rect 44166 18205 44486 18261
rect 44485 18123 44486 18205
rect 42982 14533 43112 14534
rect 42982 14405 42983 14533
rect 43111 14405 43112 14533
rect 42982 14404 43112 14405
rect 44812 13992 44940 19339
rect 47010 20767 47138 20788
rect 47010 20703 47042 20767
rect 47106 20703 47138 20767
rect 47010 18761 47138 20703
rect 47795 19843 47923 21718
rect 49330 21583 49458 21608
rect 49330 21519 49362 21583
rect 49426 21519 49458 21583
rect 48602 20577 48732 20578
rect 48602 20449 48603 20577
rect 48731 20449 48732 20577
rect 48602 20448 48732 20449
rect 47790 19842 47923 19843
rect 47790 19714 47791 19842
rect 47919 19714 47923 19842
rect 47790 19713 47923 19714
rect 47010 18697 47040 18761
rect 47104 18697 47138 18761
rect 44811 13991 44941 13992
rect 44811 13863 44812 13991
rect 44940 13863 44941 13991
rect 44811 13862 44941 13863
rect 47010 12351 47138 18697
rect 47795 18146 47923 19713
rect 48603 18579 48731 20448
rect 49330 19582 49458 21519
rect 49330 19518 49357 19582
rect 49421 19518 49458 19582
rect 48602 18578 48732 18579
rect 48602 18450 48603 18578
rect 48731 18450 48732 18578
rect 48602 18449 48732 18450
rect 48603 15172 48731 18449
rect 47009 12350 47139 12351
rect 47009 12222 47010 12350
rect 47138 12222 47139 12350
rect 47009 12221 47139 12222
rect 49330 11809 49458 19518
rect 50477 16762 50605 22704
rect 51944 22588 52062 22877
rect 51939 22587 52062 22588
rect 51939 22469 51940 22587
rect 52058 22482 52062 22587
rect 52058 22469 52059 22482
rect 51939 22468 52059 22469
rect 51103 17840 51223 17841
rect 51103 17722 51104 17840
rect 51222 17722 51223 17840
rect 51103 17721 51223 17722
rect 50477 16698 50503 16762
rect 50567 16698 50605 16762
rect 49329 11808 49459 11809
rect 49329 11680 49330 11808
rect 49458 11680 49459 11808
rect 49329 11679 49459 11680
rect 50477 7463 50605 16698
rect 52517 17580 52645 23516
rect 64415 23588 64543 23640
rect 64415 23514 64440 23588
rect 64514 23514 64543 23588
rect 60238 21871 60358 21872
rect 60238 21753 60239 21871
rect 60357 21753 60358 21871
rect 60238 21752 60358 21753
rect 52517 17516 52547 17580
rect 52611 17516 52645 17580
rect 51816 16582 51936 16583
rect 51816 16464 51817 16582
rect 51935 16563 51936 16582
rect 51935 16464 51939 16563
rect 51816 16463 51939 16464
rect 51821 15195 51939 16463
rect 52517 7999 52645 17516
rect 59672 20768 59800 20940
rect 59672 20694 59693 20768
rect 59767 20694 59800 20768
rect 59672 18764 59800 20694
rect 59672 18700 59710 18764
rect 59774 18700 59800 18764
rect 59672 11265 59800 18700
rect 60239 19842 60357 21752
rect 61061 20580 61179 22953
rect 62392 22765 62520 22793
rect 62392 22691 62415 22765
rect 62489 22691 62520 22765
rect 61642 21589 61770 21617
rect 61642 21515 61659 21589
rect 61733 21515 61770 21589
rect 61060 20579 61180 20580
rect 61060 20461 61061 20579
rect 61179 20461 61180 20579
rect 61060 20460 61180 20461
rect 60239 19841 60360 19842
rect 60239 19723 60241 19841
rect 60359 19723 60360 19841
rect 60239 19722 60360 19723
rect 60239 18233 60357 19722
rect 61061 18584 61179 20460
rect 61054 18583 61179 18584
rect 61054 18465 61055 18583
rect 61173 18485 61179 18583
rect 61642 19586 61770 21515
rect 61642 19512 61662 19586
rect 61736 19512 61770 19586
rect 61173 18465 61174 18485
rect 61054 18464 61174 18465
rect 59671 11264 59801 11265
rect 59671 11136 59672 11264
rect 59800 11136 59801 11264
rect 59671 11135 59801 11136
rect 61642 10726 61770 19512
rect 62392 16768 62520 22691
rect 63864 22583 63982 22857
rect 63859 22582 63982 22583
rect 63859 22464 63860 22582
rect 63978 22525 63982 22582
rect 63978 22464 63979 22525
rect 63859 22463 63979 22464
rect 63016 17834 63134 17895
rect 63014 17833 63134 17834
rect 63014 17715 63015 17833
rect 63133 17715 63134 17833
rect 63014 17714 63134 17715
rect 62392 16694 62416 16768
rect 62490 16694 62520 16768
rect 61641 10725 61771 10726
rect 61641 10597 61642 10725
rect 61770 10597 61771 10725
rect 61641 10596 61771 10597
rect 62392 8549 62520 16694
rect 64415 17582 64543 23514
rect 72846 23592 72974 23618
rect 72846 23518 72870 23592
rect 72944 23518 72974 23592
rect 67124 20795 67252 20819
rect 67124 20731 67161 20795
rect 67225 20731 67252 20795
rect 66647 20333 66765 20338
rect 66647 20332 66768 20333
rect 66647 20214 66649 20332
rect 66767 20214 66768 20332
rect 66647 20213 66768 20214
rect 66647 18200 66765 20213
rect 67124 19825 67252 20731
rect 67124 19761 67163 19825
rect 67227 19761 67252 19825
rect 64415 17518 64442 17582
rect 64506 17518 64543 17582
rect 63826 16573 63946 16574
rect 63826 16455 63827 16573
rect 63945 16455 63946 16573
rect 63826 16454 63946 16455
rect 63826 15246 63944 16454
rect 64415 9085 64543 17518
rect 67124 14534 67252 19761
rect 67969 20792 68097 20816
rect 67969 20728 67989 20792
rect 68053 20728 68097 20792
rect 67969 19826 68097 20728
rect 68386 20325 68504 22911
rect 71156 22766 71284 22799
rect 71156 22692 71181 22766
rect 71255 22692 71284 22766
rect 68385 20324 68505 20325
rect 68385 20206 68386 20324
rect 68504 20206 68505 20324
rect 68385 20205 68505 20206
rect 67969 19762 67985 19826
rect 68049 19762 68097 19826
rect 67123 14533 67253 14534
rect 67123 14405 67124 14533
rect 67252 14405 67253 14533
rect 67123 14404 67253 14405
rect 67969 13992 68097 19762
rect 71156 16779 71284 22692
rect 72435 22579 72553 22901
rect 72434 22578 72554 22579
rect 72434 22460 72435 22578
rect 72553 22460 72554 22578
rect 72434 22459 72554 22460
rect 71483 18190 71823 18203
rect 71483 17870 71485 18190
rect 71805 17870 71823 18190
rect 71483 17844 71823 17870
rect 71483 17797 71584 17844
rect 71583 17726 71584 17797
rect 71702 17797 71823 17844
rect 71702 17777 71704 17797
rect 71702 17726 71703 17777
rect 71583 17725 71703 17726
rect 71156 16705 71185 16779
rect 71259 16705 71284 16779
rect 67968 13991 68098 13992
rect 67968 13863 67969 13991
rect 68097 13863 68098 13991
rect 67968 13862 68098 13863
rect 64414 9084 64544 9085
rect 64414 8956 64415 9084
rect 64543 8956 64544 9084
rect 64414 8955 64544 8956
rect 62391 8548 62521 8549
rect 62391 8420 62392 8548
rect 62520 8420 62521 8548
rect 62391 8419 62521 8420
rect 52516 7998 52646 7999
rect 52516 7870 52517 7998
rect 52645 7870 52646 7998
rect 52516 7869 52646 7870
rect 50476 7462 50606 7463
rect 50476 7334 50477 7462
rect 50605 7334 50606 7462
rect 50476 7333 50606 7334
rect 41669 5284 41799 5285
rect 41669 5156 41670 5284
rect 41798 5156 41799 5284
rect 41669 5155 41799 5156
rect 71156 2018 71284 16705
rect 72846 17599 72974 23518
rect 73566 20071 73684 22875
rect 73564 20070 73684 20071
rect 73564 19952 73565 20070
rect 73683 19952 73684 20070
rect 73564 19951 73684 19952
rect 73999 20545 74127 20574
rect 73999 20481 74028 20545
rect 74092 20481 74127 20545
rect 72846 17525 72877 17599
rect 72951 17525 72974 17599
rect 72295 16582 72415 16583
rect 72295 16464 72296 16582
rect 72414 16464 72415 16582
rect 72295 16463 72415 16464
rect 72295 15191 72413 16463
rect 72846 2564 72974 17525
rect 73999 19583 74127 20481
rect 73999 19519 74034 19583
rect 74098 19519 74127 19583
rect 73999 4726 74127 19519
rect 73999 4600 74000 4726
rect 74126 4600 74127 4726
rect 73999 4599 74127 4600
rect 74813 20551 74941 20572
rect 74813 20487 74856 20551
rect 74920 20487 74941 20551
rect 74813 19582 74941 20487
rect 74813 19518 74860 19582
rect 74924 19518 74941 19582
rect 74813 4192 74941 19518
rect 75275 20093 75395 20094
rect 75275 19975 75276 20093
rect 75394 19975 75395 20093
rect 75275 19974 75395 19975
rect 75275 18144 75393 19974
rect 74812 4191 74942 4192
rect 74812 4063 74813 4191
rect 74941 4063 74942 4191
rect 74812 4062 74942 4063
rect 72845 2563 72975 2564
rect 72845 2435 72846 2563
rect 72974 2435 72975 2563
rect 72845 2434 72975 2435
rect 71155 2017 71285 2018
rect 71155 1889 71156 2017
rect 71284 1889 71285 2017
rect 71155 1888 71285 1889
rect 38276 1466 38406 1467
rect 38276 1338 38277 1466
rect 38405 1338 38406 1466
rect 38276 1337 38406 1338
rect 36247 935 36377 936
rect 36247 807 36248 935
rect 36376 807 36377 935
rect 36247 806 36377 807
rect 75720 919 75848 36965
rect 76121 1459 76249 36964
rect 76520 5809 76646 36991
rect 76520 5685 76521 5809
rect 76645 5685 76646 5809
rect 76520 5684 76646 5685
rect 76909 5268 77033 36983
rect 76909 5146 76910 5268
rect 77032 5146 77033 5268
rect 76909 5145 77033 5146
rect 78108 2018 78236 41343
rect 79804 40740 79965 41893
rect 81823 40750 81962 41893
rect 88514 41756 88642 41757
rect 88514 41630 88515 41756
rect 88641 41630 88642 41756
rect 85864 41241 86138 41252
rect 85864 41005 85883 41241
rect 86119 41005 86138 41241
rect 85864 40988 86138 41005
rect 87796 41223 88032 41236
rect 87796 41012 87808 41223
rect 88019 41012 88032 41223
rect 87796 41000 88032 41012
rect 79804 40739 79984 40740
rect 79804 40499 79904 40739
rect 79903 40461 79904 40499
rect 79983 40461 79984 40739
rect 79903 40460 79984 40461
rect 81822 40703 82060 40750
rect 81822 40420 81965 40703
rect 82045 40420 82060 40703
rect 81822 40393 82060 40420
rect 79093 39949 79221 39950
rect 79093 39823 79094 39949
rect 79220 39823 79221 39949
rect 79093 2564 79221 39823
rect 80840 39719 83228 39798
rect 80840 39704 83018 39719
rect 80840 39576 81162 39704
rect 81290 39595 83018 39704
rect 83142 39595 83228 39719
rect 81290 39576 83228 39595
rect 80840 39478 83228 39576
rect 81530 39193 81850 39478
rect 85888 39205 86114 40988
rect 87813 39207 88014 41000
rect 82211 34922 82275 35607
rect 81216 34918 83541 34922
rect 85220 34920 85284 35655
rect 86360 35330 86514 35338
rect 86360 35192 86368 35330
rect 86506 35192 86514 35330
rect 86360 35183 86514 35192
rect 86373 34920 86501 35183
rect 81216 34890 83557 34918
rect 83771 34895 83928 34908
rect 83771 34890 83780 34895
rect 81216 34858 83780 34890
rect 81216 30850 81280 34858
rect 83471 34762 83780 34858
rect 83477 34712 83557 34762
rect 83771 34757 83780 34762
rect 83918 34757 83928 34895
rect 83771 34736 83928 34757
rect 84215 34856 86534 34920
rect 82259 31894 82323 33614
rect 82231 31334 82349 31636
rect 82231 31218 82232 31334
rect 82348 31218 82349 31334
rect 82231 31217 82349 31218
rect 83477 30654 83541 34712
rect 81222 30590 83541 30654
rect 84215 30652 84279 34856
rect 85433 31896 85497 33616
rect 85519 31835 85912 31836
rect 85519 31719 85795 31835
rect 85911 31719 85912 31835
rect 85519 31718 85912 31719
rect 86476 30652 86540 34660
rect 82216 29893 82280 30590
rect 84215 30588 86540 30652
rect 85218 29886 85282 30588
rect 81845 23543 81973 23613
rect 81845 23469 81872 23543
rect 81946 23469 81973 23543
rect 81845 17572 81973 23469
rect 82259 22523 82377 25916
rect 85178 24732 85306 24759
rect 85178 24658 85207 24732
rect 85281 24658 85306 24732
rect 83057 23773 83175 23782
rect 83054 23772 83175 23773
rect 83054 23654 83055 23772
rect 83173 23654 83175 23772
rect 83054 23653 83175 23654
rect 83057 23225 83175 23653
rect 82255 22522 82377 22523
rect 82255 22404 82256 22522
rect 82374 22414 82377 22522
rect 83425 22716 83553 23515
rect 83425 22642 83454 22716
rect 83528 22642 83553 22716
rect 82374 22404 82375 22414
rect 82255 22403 82375 22404
rect 81845 17498 81877 17572
rect 81951 17498 81973 17572
rect 79092 2563 79222 2564
rect 79092 2435 79093 2563
rect 79221 2435 79222 2563
rect 79092 2434 79222 2435
rect 78107 2017 78237 2018
rect 78107 1889 78108 2017
rect 78236 1889 78237 2017
rect 78107 1888 78237 1889
rect 76121 1333 76122 1459
rect 76248 1333 76249 1459
rect 76121 1332 76249 1333
rect 81845 936 81973 17498
rect 82303 16562 82421 17851
rect 82967 17813 83089 17814
rect 82967 17695 82968 17813
rect 83086 17695 83089 17813
rect 82967 17694 83089 17695
rect 82295 16561 82421 16562
rect 82295 16443 82296 16561
rect 82414 16483 82421 16561
rect 82414 16443 82415 16483
rect 82295 16442 82415 16443
rect 82971 15215 83089 17694
rect 83425 16752 83553 22642
rect 83425 16678 83450 16752
rect 83524 16678 83553 16752
rect 83425 1467 83553 16678
rect 85178 16722 85306 24658
rect 85591 23723 85709 25883
rect 86377 24989 86495 24993
rect 86376 24988 86496 24989
rect 86376 24870 86377 24988
rect 86495 24870 86496 24988
rect 86376 24869 86496 24870
rect 85590 23722 85710 23723
rect 85590 23604 85591 23722
rect 85709 23604 85710 23722
rect 85590 23603 85710 23604
rect 85591 23599 85709 23603
rect 86377 23220 86495 24869
rect 86989 23907 87117 23967
rect 86989 23833 87014 23907
rect 87088 23833 87117 23907
rect 85178 16648 85205 16722
rect 85279 16648 85306 16722
rect 85178 5822 85306 16648
rect 85631 15696 85749 17918
rect 86413 16963 86531 16990
rect 86411 16962 86531 16963
rect 86411 16844 86412 16962
rect 86530 16844 86531 16962
rect 86411 16843 86531 16844
rect 85623 15695 85749 15696
rect 85623 15577 85624 15695
rect 85742 15595 85749 15695
rect 85742 15577 85743 15595
rect 85623 15576 85743 15577
rect 86413 15188 86531 16843
rect 86989 15897 87117 23833
rect 86989 15823 87011 15897
rect 87085 15823 87117 15897
rect 85177 5821 85307 5822
rect 85177 5693 85178 5821
rect 85306 5693 85307 5821
rect 85177 5692 85307 5693
rect 86989 5285 87117 15823
rect 86988 5284 87118 5285
rect 86988 5156 86989 5284
rect 87117 5156 87118 5284
rect 86988 5155 87118 5156
rect 88514 4192 88642 41630
rect 89566 4740 89694 43153
rect 96365 42681 98263 42719
rect 96365 42342 96525 42681
rect 96795 42678 98263 42681
rect 96795 42342 97372 42678
rect 97642 42396 98263 42678
rect 97642 42342 97972 42396
rect 96365 41738 96466 42342
rect 97687 41738 97972 42342
rect 96365 41606 96525 41738
rect 96795 41606 97372 41738
rect 96365 41603 97372 41606
rect 97642 41682 97972 41738
rect 98218 41682 98263 42396
rect 97642 41603 98263 41682
rect 96365 41575 98263 41603
rect 155830 39405 157830 46705
rect 114708 39378 115009 39379
rect 90782 38958 90794 38959
rect 90782 38091 90783 38958
rect 91030 38091 91031 38748
rect 114708 38737 114709 39378
rect 115008 38737 115009 39378
rect 114708 38736 115009 38737
rect 90782 38090 91031 38091
rect 122924 38345 123200 38372
rect 98570 37299 109720 37552
rect 98570 37239 103349 37299
rect 98570 37232 101446 37239
rect 96848 35851 97597 35852
rect 96848 35836 96849 35851
rect 96846 35740 96849 35836
rect 97596 35836 97597 35851
rect 97596 35740 97601 35836
rect 91353 35536 94747 35537
rect 91353 35332 91354 35536
rect 91558 35332 94542 35536
rect 94746 35332 94747 35536
rect 91353 35331 94747 35332
rect 91311 34383 95471 34384
rect 91311 34179 91312 34383
rect 91516 34179 95265 34383
rect 95470 34179 95471 34383
rect 91311 34178 95471 34179
rect 96846 34291 97601 35740
rect 90787 30813 90805 30935
rect 95426 31246 95712 31247
rect 95426 31243 95427 31246
rect 90787 30752 91087 30813
rect 90787 30288 90814 30752
rect 91056 30288 91087 30752
rect 90787 30268 91087 30288
rect 95424 30789 95427 31243
rect 95711 30789 95712 31246
rect 98570 31241 98890 37232
rect 99810 37228 100130 37232
rect 99810 37028 99844 37228
rect 100088 37028 100130 37228
rect 101445 37039 101446 37232
rect 101690 37232 103349 37239
rect 101690 37039 101691 37232
rect 103348 37099 103349 37232
rect 103593 37283 109720 37299
rect 103593 37232 105066 37283
rect 103593 37099 103594 37232
rect 103348 37098 103594 37099
rect 105065 37083 105066 37232
rect 105310 37278 109720 37283
rect 105310 37232 106880 37278
rect 105310 37083 105311 37232
rect 105065 37082 105311 37083
rect 106879 37078 106880 37232
rect 107124 37272 109720 37278
rect 107124 37232 108852 37272
rect 107124 37078 107125 37232
rect 106879 37077 107125 37078
rect 108851 37072 108852 37232
rect 109096 37232 109720 37272
rect 109096 37072 109097 37232
rect 108851 37071 109097 37072
rect 101445 37038 101691 37039
rect 122924 37052 123011 38345
rect 123095 38339 123200 38345
rect 123095 37052 123201 38339
rect 99810 37021 100130 37028
rect 122924 36885 123201 37052
rect 102158 35735 102560 35736
rect 102156 35734 102560 35735
rect 100356 35727 100757 35733
rect 100356 35649 100366 35727
rect 100750 35649 100757 35727
rect 102156 35660 102157 35734
rect 102557 35660 102560 35734
rect 102156 35659 102560 35660
rect 103962 35734 104352 35735
rect 103962 35660 103963 35734
rect 104351 35660 104352 35734
rect 103962 35659 104352 35660
rect 105759 35699 106149 35700
rect 100356 35539 100757 35649
rect 102158 35539 102560 35659
rect 104029 35539 104297 35659
rect 105759 35625 105760 35699
rect 106148 35625 106149 35699
rect 105759 35624 106149 35625
rect 107560 35699 107951 35704
rect 105760 35539 106148 35624
rect 107560 35621 107562 35699
rect 107949 35621 107951 35699
rect 107560 35539 107951 35621
rect 109352 35695 109753 35698
rect 109352 35618 109356 35695
rect 109751 35618 109753 35695
rect 109352 35539 109753 35618
rect 99692 35219 109772 35539
rect 104794 34198 105114 35219
rect 95424 30788 95712 30789
rect 95424 28685 95704 30788
rect 95202 28684 95763 28685
rect 95202 28464 95203 28684
rect 95762 28464 95763 28684
rect 95202 28463 95763 28464
rect 107960 27190 108080 27191
rect 104387 27177 104517 27178
rect 104387 27049 104388 27177
rect 104516 27049 104517 27177
rect 107960 27062 107961 27190
rect 108079 27062 108080 27190
rect 107960 27061 108080 27062
rect 104387 27048 104517 27049
rect 91367 22717 91495 22767
rect 91367 22643 91387 22717
rect 91461 22643 91495 22717
rect 91367 16748 91495 22643
rect 91882 22529 92000 25860
rect 92589 23788 92709 23789
rect 92589 23670 92590 23788
rect 92708 23670 92709 23788
rect 92589 23669 92709 23670
rect 92589 23205 92707 23669
rect 93107 23542 93235 23569
rect 93107 23468 93131 23542
rect 93205 23468 93235 23542
rect 91881 22528 92001 22529
rect 91881 22410 91882 22528
rect 92000 22410 92001 22528
rect 91881 22409 92001 22410
rect 91367 16674 91397 16748
rect 91471 16674 91495 16748
rect 91367 14534 91495 16674
rect 91859 16548 91977 17843
rect 92565 17819 92685 17820
rect 92565 17701 92566 17819
rect 92684 17701 92685 17819
rect 92565 17700 92685 17701
rect 91858 16547 91978 16548
rect 91858 16429 91859 16547
rect 91977 16429 91978 16547
rect 91858 16428 91978 16429
rect 92566 15235 92684 17700
rect 93107 17567 93235 23468
rect 104393 22682 104511 27048
rect 107961 26657 108079 27061
rect 107961 26386 108097 26657
rect 106334 25920 106501 26144
rect 106268 25918 106501 25920
rect 106373 23429 106501 25918
rect 106371 23428 106501 23429
rect 106371 23300 106372 23428
rect 106500 23300 106501 23428
rect 106371 23299 106501 23300
rect 105384 23165 105512 23193
rect 105384 23091 105417 23165
rect 105491 23091 105512 23165
rect 104384 22674 104518 22682
rect 104384 22558 104394 22674
rect 104510 22558 104518 22674
rect 104384 22544 104518 22558
rect 93107 17503 93134 17567
rect 93198 17503 93235 17567
rect 91366 14533 91496 14534
rect 91366 14405 91367 14533
rect 91495 14405 91496 14533
rect 91366 14404 91496 14405
rect 93107 13992 93235 17503
rect 105384 14534 105512 23091
rect 105806 22157 105934 22857
rect 105795 22156 105934 22157
rect 105795 22028 105796 22156
rect 105924 22057 105934 22156
rect 107068 22355 107196 23242
rect 107979 22693 108097 26386
rect 107979 22577 107980 22693
rect 108096 22577 108097 22693
rect 107979 22576 108097 22577
rect 107068 22271 107090 22355
rect 107174 22271 107196 22355
rect 105924 22028 105925 22057
rect 105795 22027 105925 22028
rect 105383 14533 105513 14534
rect 105383 14405 105384 14533
rect 105512 14405 105513 14533
rect 105383 14404 105513 14405
rect 107068 13992 107196 22271
rect 93106 13991 93236 13992
rect 93106 13863 93107 13991
rect 93235 13863 93236 13991
rect 93106 13862 93236 13863
rect 107067 13991 107197 13992
rect 107067 13863 107068 13991
rect 107196 13863 107197 13991
rect 107067 13862 107197 13863
rect 89565 4739 89695 4740
rect 89565 4611 89566 4739
rect 89694 4611 89695 4739
rect 89565 4610 89695 4611
rect 88513 4191 88643 4192
rect 88513 4063 88514 4191
rect 88642 4063 88643 4191
rect 88513 4062 88643 4063
rect 83424 1466 83554 1467
rect 83424 1338 83425 1466
rect 83553 1338 83554 1466
rect 83424 1337 83554 1338
rect 75720 793 75721 919
rect 75847 793 75848 919
rect 81844 935 81974 936
rect 81844 807 81845 935
rect 81973 807 81974 935
rect 110235 931 110357 36787
rect 110634 1458 110756 36784
rect 111039 5797 111159 36786
rect 111039 5679 111040 5797
rect 111158 5679 111159 5797
rect 111039 5678 111159 5679
rect 111438 5273 111556 36790
rect 122924 35592 123011 36885
rect 123095 35592 123201 36885
rect 122924 35432 123201 35592
rect 122910 35405 123201 35432
rect 122910 34622 123012 35405
rect 122924 34387 123012 34622
rect 123095 34387 123201 35405
rect 122924 34384 123201 34387
rect 119412 34040 119540 34041
rect 119412 33914 119413 34040
rect 119539 33914 119540 34040
rect 114715 31367 115016 31368
rect 114715 30726 114716 31367
rect 115015 30726 115016 31367
rect 114715 30725 115016 30726
rect 111438 5157 111439 5273
rect 111555 5157 111556 5273
rect 111438 5156 111556 5157
rect 119412 1467 119540 33914
rect 122924 33723 122951 34384
rect 125027 34131 125349 34132
rect 125027 33811 125028 34131
rect 125348 33811 125349 34131
rect 125027 33810 125349 33811
rect 127171 33739 127633 33771
rect 122924 33617 123201 33723
rect 127171 33666 127217 33739
rect 127594 33666 127633 33739
rect 127171 33665 127633 33666
rect 122924 32643 123010 33617
rect 123097 32643 123201 33617
rect 122924 32470 123201 32643
rect 127218 32617 127592 32618
rect 127218 32552 127219 32617
rect 127591 32552 127592 32617
rect 127218 32551 127592 32552
rect 122924 31104 123007 32470
rect 123097 31104 123201 32470
rect 127347 31321 127475 32551
rect 155830 31405 157830 38705
rect 122924 30864 123201 31104
rect 124328 31186 124650 31187
rect 124328 30866 124329 31186
rect 124649 30866 124650 31186
rect 124328 30865 124650 30866
rect 122924 29606 123008 30864
rect 123099 29606 123201 30864
rect 122924 29575 123201 29606
rect 122924 29570 123200 29575
rect 155830 23405 157830 30705
rect 155830 15405 157830 22705
rect 120733 12351 120861 12826
rect 120733 12350 120864 12351
rect 120733 12222 120735 12350
rect 120863 12222 120864 12350
rect 120733 12221 120864 12222
rect 110634 1338 110635 1458
rect 110755 1338 110756 1458
rect 110634 1337 110756 1338
rect 119411 1466 119541 1467
rect 119411 1338 119412 1466
rect 119540 1338 119541 1466
rect 119411 1337 119541 1338
rect 110235 811 110236 931
rect 110356 811 110357 931
rect 110235 810 110357 811
rect 81844 806 81974 807
rect 75720 792 75848 793
rect 13965 -8595 15965 -1295
rect 67103 -2038 67170 -1266
rect 67102 -2039 67171 -2038
rect 67102 -2665 67103 -2039
rect 67170 -2665 67171 -2039
rect 67102 -2666 67171 -2665
rect 120733 -3363 120861 12221
rect 121333 11809 121461 12826
rect 121332 11808 121462 11809
rect 121332 11680 121333 11808
rect 121461 11680 121462 11808
rect 121332 11679 121462 11680
rect 120733 -3429 120757 -3363
rect 120823 -3429 120861 -3363
rect 120733 -5121 120861 -3429
rect 121333 -2806 121461 11679
rect 121333 -2872 121368 -2806
rect 121434 -2872 121461 -2806
rect 121333 -5121 121461 -2872
rect 121933 11265 122061 12826
rect 121933 11264 122066 11265
rect 121933 11136 121937 11264
rect 122065 11136 122066 11264
rect 121933 11135 122066 11136
rect 121933 -399 122061 11135
rect 121933 -465 121979 -399
rect 122045 -465 122061 -399
rect 121933 -5121 122061 -465
rect 122533 10726 122661 12826
rect 122533 10725 122670 10726
rect 122533 10597 122541 10725
rect 122669 10597 122670 10725
rect 122533 10596 122670 10597
rect 122533 158 122661 10596
rect 122533 92 122561 158
rect 122627 92 122661 158
rect 122533 -5121 122661 92
rect 123733 9085 123861 12826
rect 123733 9084 123866 9085
rect 123733 8956 123737 9084
rect 123865 8956 123866 9084
rect 123733 8955 123866 8956
rect 123733 -1159 123861 8955
rect 123733 -1225 123743 -1159
rect 123809 -1225 123861 -1159
rect 123733 -5121 123861 -1225
rect 124333 8549 124461 12826
rect 124333 8548 124464 8549
rect 124333 8420 124335 8548
rect 124463 8420 124464 8548
rect 124333 8419 124464 8420
rect 124333 -1716 124461 8419
rect 124333 -1782 124353 -1716
rect 124419 -1782 124461 -1716
rect 124333 -5121 124461 -1782
rect 124933 7999 125061 12826
rect 124933 7998 125068 7999
rect 124933 7870 124939 7998
rect 125067 7870 125068 7998
rect 124933 7869 125068 7870
rect 124933 -4053 125061 7869
rect 124933 -4119 124958 -4053
rect 125024 -4119 125061 -4053
rect 124933 -5121 125061 -4119
rect 125533 7463 125661 12826
rect 125533 7462 125666 7463
rect 125533 7334 125537 7462
rect 125665 7334 125666 7462
rect 125533 7333 125666 7334
rect 125533 -4610 125661 7333
rect 125533 -4676 125568 -4610
rect 125634 -4676 125661 -4610
rect 125533 -5121 125661 -4676
rect 126733 5822 126861 12826
rect 126733 5821 126868 5822
rect 126733 5693 126739 5821
rect 126867 5693 126868 5821
rect 126733 5692 126868 5693
rect 126733 -3630 126861 5692
rect 126733 -3696 126763 -3630
rect 126829 -3696 126861 -3630
rect 126733 -5121 126861 -3696
rect 127333 5285 127461 12826
rect 127333 5284 127468 5285
rect 127333 5156 127339 5284
rect 127467 5156 127468 5284
rect 127333 5155 127468 5156
rect 127333 -3064 127461 5155
rect 127933 4740 128061 12826
rect 127932 4739 128062 4740
rect 127932 4611 127933 4739
rect 128061 4611 128062 4739
rect 127932 4610 128062 4611
rect 127333 -3130 127364 -3064
rect 127430 -3130 127461 -3064
rect 127333 -5121 127461 -3130
rect 127933 -666 128061 4610
rect 127933 -732 127947 -666
rect 128013 -732 128061 -666
rect 127933 -5121 128061 -732
rect 128533 4192 128661 12826
rect 128533 4191 128674 4192
rect 128533 4063 128545 4191
rect 128673 4063 128674 4191
rect 128533 4062 128674 4063
rect 128533 -100 128661 4062
rect 128533 -166 128558 -100
rect 128624 -166 128661 -100
rect 128533 -5121 128661 -166
rect 129733 2564 129861 12826
rect 129733 2563 129877 2564
rect 129733 2435 129748 2563
rect 129876 2435 129877 2563
rect 129733 2434 129877 2435
rect 129733 -1417 129861 2434
rect 130333 2018 130461 12826
rect 130330 2017 130461 2018
rect 130330 1889 130331 2017
rect 130459 1889 130461 2017
rect 130330 1888 130461 1889
rect 129733 -1483 129766 -1417
rect 129832 -1483 129861 -1417
rect 129733 -5121 129861 -1483
rect 130333 -1983 130461 1888
rect 130333 -2049 130362 -1983
rect 130428 -2049 130461 -1983
rect 130333 -5121 130461 -2049
rect 130933 1467 131061 12826
rect 130933 1466 131065 1467
rect 130933 1338 130936 1466
rect 131064 1338 131065 1466
rect 130933 1337 131065 1338
rect 130933 -4311 131061 1337
rect 131533 936 131661 12826
rect 155830 7405 157830 14705
rect 131529 935 131661 936
rect 131529 807 131530 935
rect 131658 807 131661 935
rect 131529 806 131661 807
rect 130933 -4377 130963 -4311
rect 131029 -4377 131061 -4311
rect 130933 -5121 131061 -4377
rect 131533 -4877 131661 806
rect 131533 -4943 131556 -4877
rect 131622 -4943 131661 -4877
rect 131533 -5121 131661 -4943
rect 135364 33 135912 1776
rect 135364 -36 135402 33
rect 135875 -36 135912 33
rect 135364 -1282 135912 -36
rect 139037 -513 139585 448
rect 139037 -577 139082 -513
rect 139544 -577 139585 -513
rect 139037 -651 139585 -577
rect 139584 -1210 139585 -651
rect 135364 -1351 135405 -1282
rect 135878 -1351 135912 -1282
rect 135364 -2928 135912 -1351
rect 135364 -2997 135397 -2928
rect 135870 -2997 135912 -2928
rect 135364 -4178 135912 -2997
rect 135364 -4247 135399 -4178
rect 135872 -4247 135912 -4178
rect 66559 -5627 66628 -5626
rect 66559 -5628 66560 -5627
rect 66627 -5628 66628 -5627
rect 135364 -5686 135912 -4247
rect 139037 -1827 139585 -1210
rect 139037 -1891 139092 -1827
rect 139554 -1891 139585 -1827
rect 139037 -3477 139585 -1891
rect 139037 -3541 139082 -3477
rect 139544 -3541 139585 -3477
rect 139037 -4724 139585 -3541
rect 139037 -4788 139097 -4724
rect 139559 -4788 139585 -4724
rect 139037 -5091 139585 -4788
rect 155830 -595 157830 6705
rect 13965 -16595 15965 -9295
rect 147296 -11156 147844 -6226
rect 155830 -8595 157830 -1295
rect 147296 -11225 147329 -11156
rect 147802 -11225 147844 -11156
rect 147296 -11260 147844 -11225
rect 150970 -11705 151518 -9216
rect 150970 -11769 151014 -11705
rect 151476 -11769 151518 -11705
rect 150970 -11804 151518 -11769
rect 155830 -16595 157830 -9295
rect 71620 -16617 71686 -16616
rect 71620 -16625 71621 -16617
rect 71685 -16625 71686 -16617
rect 72708 -16617 72774 -16616
rect 72708 -16625 72709 -16617
rect 72773 -16625 72774 -16617
rect 73796 -16617 73862 -16616
rect 73796 -16625 73797 -16617
rect 73861 -16625 73862 -16617
rect 74884 -16617 74950 -16616
rect 74884 -16625 74885 -16617
rect 74949 -16625 74950 -16617
rect 75972 -16617 76038 -16616
rect 75972 -16625 75973 -16617
rect 76037 -16625 76038 -16617
rect 77060 -16617 77126 -16616
rect 77060 -16625 77061 -16617
rect 77125 -16625 77126 -16617
rect 78148 -16617 78214 -16616
rect 78148 -16625 78149 -16617
rect 78213 -16625 78214 -16617
rect 79236 -16617 79302 -16616
rect 79236 -16625 79237 -16617
rect 79301 -16625 79302 -16617
rect 80324 -16617 80390 -16616
rect 80324 -16625 80325 -16617
rect 80389 -16625 80390 -16617
rect 81412 -16617 81478 -16616
rect 81412 -16625 81413 -16617
rect 81477 -16625 81478 -16617
rect 82500 -16617 82566 -16616
rect 82500 -16625 82501 -16617
rect 82565 -16625 82566 -16617
rect 83588 -16617 83654 -16616
rect 83588 -16625 83589 -16617
rect 83653 -16625 83654 -16617
rect 84676 -16617 84742 -16616
rect 84676 -16625 84677 -16617
rect 84741 -16625 84742 -16617
rect 71620 -17271 71621 -17264
rect 71685 -17271 71686 -17264
rect 71620 -17272 71686 -17271
rect 72708 -17271 72709 -17264
rect 72773 -17271 72774 -17264
rect 72708 -17272 72774 -17271
rect 73796 -17271 73797 -17264
rect 73861 -17271 73862 -17264
rect 73796 -17272 73862 -17271
rect 74884 -17271 74885 -17264
rect 74949 -17271 74950 -17264
rect 74884 -17272 74950 -17271
rect 75972 -17271 75973 -17264
rect 76037 -17271 76038 -17264
rect 75972 -17272 76038 -17271
rect 77060 -17271 77061 -17264
rect 77125 -17271 77126 -17264
rect 77060 -17272 77126 -17271
rect 78148 -17271 78149 -17264
rect 78213 -17271 78214 -17264
rect 78148 -17272 78214 -17271
rect 79236 -17271 79237 -17264
rect 79301 -17271 79302 -17264
rect 79236 -17272 79302 -17271
rect 80324 -17271 80325 -17264
rect 80389 -17271 80390 -17264
rect 80324 -17272 80390 -17271
rect 81412 -17271 81413 -17264
rect 81477 -17271 81478 -17264
rect 81412 -17272 81478 -17271
rect 82500 -17271 82501 -17264
rect 82565 -17271 82566 -17264
rect 82500 -17272 82566 -17271
rect 83588 -17271 83589 -17264
rect 83653 -17271 83654 -17264
rect 83588 -17272 83654 -17271
rect 84676 -17271 84677 -17264
rect 84741 -17271 84742 -17264
rect 84676 -17272 84742 -17271
rect 13965 -24595 15965 -17295
rect 71074 -21612 71143 -21611
rect 71074 -21630 71075 -21612
rect 71142 -21630 71143 -21612
rect 72164 -21618 72233 -21617
rect 72164 -21646 72165 -21618
rect 72232 -21646 72233 -21618
rect 73252 -21618 73321 -21617
rect 73252 -21646 73253 -21618
rect 73320 -21646 73321 -21618
rect 74340 -21618 74409 -21617
rect 74340 -21646 74341 -21618
rect 74408 -21646 74409 -21618
rect 75428 -21618 75497 -21617
rect 75428 -21646 75429 -21618
rect 75496 -21646 75497 -21618
rect 76516 -21618 76585 -21617
rect 76516 -21646 76517 -21618
rect 76584 -21646 76585 -21618
rect 77604 -21618 77673 -21617
rect 77604 -21646 77605 -21618
rect 77672 -21646 77673 -21618
rect 81956 -21618 82025 -21617
rect 81956 -21646 81957 -21618
rect 82024 -21646 82025 -21618
rect 83044 -21618 83113 -21617
rect 83044 -21646 83045 -21618
rect 83112 -21646 83113 -21618
rect 84132 -21618 84201 -21617
rect 84132 -21646 84133 -21618
rect 84200 -21646 84201 -21618
rect 85220 -21618 85289 -21617
rect 85220 -21646 85221 -21618
rect 85288 -21646 85289 -21618
rect 13965 -30385 15965 -25295
rect 13965 -40917 15965 -32385
rect 155830 -24595 157830 -17295
rect 155830 -30385 157830 -25295
rect 155830 -40917 157830 -32385
rect 159830 86397 161830 91353
rect 159830 74405 161830 84397
rect 159830 66405 161830 73705
rect 159830 58405 161830 65705
rect 159830 50405 161830 57705
rect 159830 42405 161830 49705
rect 159830 34405 161830 41705
rect 159830 26405 161830 33705
rect 159830 18405 161830 25705
rect 159830 10405 161830 17705
rect 159830 2405 161830 9705
rect 159830 -5595 161830 1705
rect 159830 -13595 161830 -6295
rect 159830 -21595 161830 -14295
rect 159830 -34385 161830 -22295
rect 159830 -40917 161830 -36385
<< via4 >>
rect 9965 84397 11965 86397
rect 9965 73705 11965 74405
rect 9965 65705 11965 66405
rect 9965 57705 11965 58405
rect 9965 49705 11965 50405
rect 9965 41705 11965 42405
rect 9965 33705 11965 34405
rect 9965 25705 11965 26405
rect 9965 17705 11965 18405
rect 9965 9705 11965 10405
rect 9965 1705 11965 2405
rect 9965 -6295 11965 -5595
rect 9965 -14295 11965 -13595
rect 9965 -22295 11965 -21595
rect 9965 -36385 11965 -34385
rect 13965 80397 15965 82397
rect 155830 80397 157830 82397
rect 13965 70705 15965 71405
rect 38260 70751 38585 71345
rect 45313 70754 45638 71348
rect 59673 70772 59998 71366
rect 35087 65749 35412 66343
rect 66822 70753 67147 71347
rect 42108 65745 42433 66339
rect 76822 70746 77147 71340
rect 87678 70747 88003 71341
rect 56492 65737 56817 66331
rect 63595 65749 63920 66343
rect 68212 65784 68537 66378
rect 95977 70761 96302 71355
rect 73661 65756 73986 66350
rect 13965 62705 15965 63405
rect 62881 62754 63206 63348
rect 78180 65751 78505 66345
rect 84508 65757 84833 66351
rect 105317 70761 105642 71355
rect 86984 65835 87304 66155
rect 72881 62754 73206 63348
rect 92753 65747 93078 66341
rect 155830 70705 157830 71405
rect 102093 65747 102418 66341
rect 104659 65878 104979 66198
rect 85069 62897 85389 63217
rect 86409 62882 86729 63202
rect 102723 62897 103043 63217
rect 104063 62882 104383 63202
rect 155830 62705 157830 63405
rect 62949 57881 63269 58201
rect 13965 54705 15965 55405
rect 46028 54901 46348 55221
rect 48072 54909 48392 55229
rect 72949 57881 73269 58201
rect 85531 57898 85851 58218
rect 13965 46705 15965 47405
rect 13965 38705 15965 39405
rect 13965 30705 15965 31405
rect 13965 22705 15965 23405
rect 13965 14705 15965 15405
rect 13965 6705 15965 7405
rect 67678 54893 67998 55213
rect 77657 54897 77977 55217
rect 103185 57898 103505 58218
rect 87209 54876 87529 55196
rect 104844 54908 105164 55228
rect 115401 54900 115721 55220
rect 119915 54888 120235 55208
rect 155830 54705 157830 55405
rect 37392 50285 37636 50368
rect 37392 49792 37447 50285
rect 37447 49792 37567 50285
rect 37567 49792 37636 50285
rect 39437 50313 39681 50370
rect 37392 49739 37636 49792
rect 39437 49780 39493 50313
rect 39493 49780 39608 50313
rect 39608 49780 39681 50313
rect 39437 49741 39681 49780
rect 35841 46963 36161 47283
rect 47393 49880 47713 50200
rect 49430 49849 49750 50169
rect 62820 49801 63349 50269
rect 66106 50207 66426 50266
rect 66106 50013 66174 50207
rect 66174 50013 66362 50207
rect 66362 50013 66426 50207
rect 66106 49946 66426 50013
rect 67927 50219 68247 50265
rect 67927 49987 67970 50219
rect 67970 49987 68198 50219
rect 68198 49987 68247 50219
rect 67927 49945 68247 49987
rect 69624 50200 69944 50250
rect 69624 49968 69664 50200
rect 69664 49968 69892 50200
rect 69892 49968 69944 50200
rect 69624 49930 69944 49968
rect 71438 50211 71758 50252
rect 71438 49979 71483 50211
rect 71483 49979 71711 50211
rect 71711 49979 71758 50211
rect 71438 49932 71758 49979
rect 73214 50208 73534 50254
rect 73214 49976 73267 50208
rect 73267 49976 73495 50208
rect 73495 49976 73534 50208
rect 73214 49934 73534 49976
rect 74999 50206 75319 50250
rect 74999 49974 75052 50206
rect 75052 49974 75280 50206
rect 75280 49974 75319 50206
rect 74999 49930 75319 49974
rect 37944 46903 38264 47223
rect 56046 46741 56330 47379
rect 60427 47309 61558 47368
rect 60427 47109 60492 47309
rect 60492 47109 61496 47309
rect 61496 47109 61558 47309
rect 96360 49834 97880 50310
rect 100630 50213 100950 50272
rect 100630 50019 100698 50213
rect 100698 50019 100886 50213
rect 100886 50019 100950 50213
rect 100630 49952 100950 50019
rect 102451 50225 102771 50271
rect 102451 49993 102494 50225
rect 102494 49993 102722 50225
rect 102722 49993 102771 50225
rect 102451 49951 102771 49993
rect 104148 50206 104468 50256
rect 104148 49974 104188 50206
rect 104188 49974 104416 50206
rect 104416 49974 104468 50206
rect 104148 49936 104468 49974
rect 105962 50217 106282 50258
rect 105962 49985 106007 50217
rect 106007 49985 106235 50217
rect 106235 49985 106282 50217
rect 105962 49938 106282 49985
rect 107738 50214 108058 50260
rect 107738 49982 107791 50214
rect 107791 49982 108019 50214
rect 108019 49982 108058 50214
rect 107738 49940 108058 49982
rect 109523 50212 109843 50256
rect 109523 49980 109576 50212
rect 109576 49980 109804 50212
rect 109804 49980 109843 50212
rect 109523 49936 109843 49980
rect 117310 49908 117630 50228
rect 119717 49892 120037 50212
rect 96360 49764 96364 49834
rect 96364 49764 97874 49834
rect 97874 49764 97880 49834
rect 60427 46779 61558 47109
rect 64064 46900 64384 47220
rect 90796 46782 91108 47320
rect 94914 47300 96166 47377
rect 94914 47083 94987 47300
rect 94987 47083 96094 47300
rect 96094 47083 96166 47300
rect 94914 46794 96166 47083
rect 98588 46906 98908 47226
rect 122091 49907 122411 50227
rect 121194 46896 121514 47216
rect 155830 46705 157830 47405
rect 61951 41731 62010 42335
rect 62010 41731 62280 42335
rect 62280 41731 62857 42335
rect 62857 41731 63127 42335
rect 63127 41731 63172 42335
rect 79732 41893 80052 42213
rect 81727 41893 82047 42213
rect 84128 41917 84448 42237
rect 86270 41909 86590 42229
rect 56068 38752 56167 39337
rect 56167 38752 56350 39337
rect 55952 30754 56299 31354
rect 60380 30856 60700 31176
rect 70278 33904 70598 34224
rect 64089 30805 64409 31125
rect 41124 25829 41444 26149
rect 50965 25870 51285 26190
rect 62889 25942 63209 26262
rect 71453 25841 71773 26161
rect 37537 22884 37857 23204
rect 40296 22881 40616 23201
rect 36730 17874 37050 18194
rect 40301 17877 40621 18197
rect 43335 22933 43655 23253
rect 51843 22877 52163 23197
rect 41115 14889 41435 15209
rect 44165 17885 44485 18205
rect 47699 17826 48019 18146
rect 48507 14852 48827 15172
rect 51003 17841 51323 18161
rect 60960 22953 61280 23273
rect 51720 14875 52040 15195
rect 63763 22857 64083 23177
rect 60138 17913 60458 18233
rect 62915 17895 63235 18215
rect 68285 22911 68605 23231
rect 66546 17880 66866 18200
rect 63725 14926 64045 15246
rect 72334 22901 72654 23221
rect 71485 17870 71805 18190
rect 73465 22875 73785 23195
rect 72194 14871 72514 15191
rect 75174 17824 75494 18144
rect 81530 38873 81850 39193
rect 85841 38885 86161 39205
rect 87754 38887 88074 39207
rect 82158 25916 82478 26236
rect 85490 25883 85810 26203
rect 82956 22905 83276 23225
rect 82202 17851 82522 18171
rect 82870 14895 83190 15215
rect 86276 22900 86596 23220
rect 85530 17918 85850 18238
rect 86312 14868 86632 15188
rect 96466 41738 96525 42342
rect 96525 41738 96795 42342
rect 96795 41738 97372 42342
rect 97372 41738 97642 42342
rect 97642 41738 97687 42342
rect 90794 38958 91103 39357
rect 90794 38748 91030 38958
rect 91030 38748 91103 38958
rect 114709 38737 115008 39378
rect 155830 38705 157830 39405
rect 96846 33763 97601 34291
rect 90805 30813 91089 31270
rect 95427 30789 95711 31246
rect 104794 33878 105114 34198
rect 98570 30921 98890 31241
rect 91781 25860 92101 26180
rect 92488 22885 92808 23205
rect 91758 17843 92078 18163
rect 103333 23108 103653 23209
rect 103333 22990 103434 23108
rect 103434 22990 103552 23108
rect 103552 22990 103653 23108
rect 103333 22889 103653 22990
rect 106014 25920 106334 26240
rect 92465 14915 92785 15235
rect 105710 22857 106030 23177
rect 108903 23113 109223 23214
rect 108903 22995 109004 23113
rect 109004 22995 109122 23113
rect 109122 22995 109223 23113
rect 108903 22894 109223 22995
rect 114716 30726 115015 31367
rect 122951 33723 123238 34384
rect 125028 33811 125348 34131
rect 127109 33771 127757 34341
rect 124329 30866 124649 31186
rect 127085 30751 127733 31321
rect 155830 30705 157830 31405
rect 155830 22705 157830 23405
rect 155830 14705 157830 15405
rect 13965 -1295 15965 -595
rect 67007 -1266 67285 -627
rect 155830 6705 157830 7405
rect 135364 1776 135912 2335
rect 139036 -1210 139584 -651
rect 66477 -6253 66560 -5628
rect 66560 -6253 66627 -5628
rect 66627 -6253 66755 -5628
rect 66477 -6267 66755 -6253
rect 70975 -6283 71253 -5644
rect 74239 -6283 74517 -5644
rect 77503 -6283 77781 -5644
rect 78591 -6283 78869 -5644
rect 81855 -6283 82133 -5644
rect 85119 -6283 85397 -5644
rect 155830 -1295 157830 -595
rect 135364 -6234 135912 -5686
rect 147296 -6226 147844 -5678
rect 13965 -9295 15965 -8595
rect 71521 -9269 71799 -8630
rect 72609 -9269 72887 -8630
rect 73697 -9269 73975 -8630
rect 74785 -9269 75063 -8630
rect 75873 -9269 76151 -8630
rect 76961 -9269 77239 -8630
rect 78049 -9269 78327 -8630
rect 79137 -9269 79415 -8630
rect 80225 -9269 80503 -8630
rect 81313 -9269 81591 -8630
rect 82401 -9269 82679 -8630
rect 83489 -9269 83767 -8630
rect 84577 -9269 84855 -8630
rect 150970 -9216 151518 -8668
rect 155830 -9295 157830 -8595
rect 70961 -14268 71239 -13629
rect 72064 -14268 72342 -13629
rect 73137 -14268 73415 -13629
rect 74225 -14268 74503 -13629
rect 75313 -14268 75591 -13629
rect 76401 -14268 76679 -13629
rect 77489 -14268 77767 -13629
rect 78577 -14268 78855 -13629
rect 79665 -14268 79943 -13629
rect 80753 -14268 81031 -13629
rect 81841 -14268 82119 -13629
rect 82929 -14268 83207 -13629
rect 84017 -14268 84295 -13629
rect 85105 -14268 85383 -13629
rect 13965 -17295 15965 -16595
rect 71519 -17264 71621 -16625
rect 71621 -17264 71685 -16625
rect 71685 -17264 71797 -16625
rect 72607 -17264 72709 -16625
rect 72709 -17264 72773 -16625
rect 72773 -17264 72885 -16625
rect 73695 -17264 73797 -16625
rect 73797 -17264 73861 -16625
rect 73861 -17264 73973 -16625
rect 74783 -17264 74885 -16625
rect 74885 -17264 74949 -16625
rect 74949 -17264 75061 -16625
rect 75871 -17264 75973 -16625
rect 75973 -17264 76037 -16625
rect 76037 -17264 76149 -16625
rect 76959 -17264 77061 -16625
rect 77061 -17264 77125 -16625
rect 77125 -17264 77237 -16625
rect 78047 -17264 78149 -16625
rect 78149 -17264 78213 -16625
rect 78213 -17264 78325 -16625
rect 79135 -17264 79237 -16625
rect 79237 -17264 79301 -16625
rect 79301 -17264 79413 -16625
rect 80223 -17264 80325 -16625
rect 80325 -17264 80389 -16625
rect 80389 -17264 80501 -16625
rect 81311 -17264 81413 -16625
rect 81413 -17264 81477 -16625
rect 81477 -17264 81589 -16625
rect 82399 -17264 82501 -16625
rect 82501 -17264 82565 -16625
rect 82565 -17264 82677 -16625
rect 83487 -17264 83589 -16625
rect 83589 -17264 83653 -16625
rect 83653 -17264 83765 -16625
rect 84575 -17264 84677 -16625
rect 84677 -17264 84741 -16625
rect 84741 -17264 84853 -16625
rect 155830 -17295 157830 -16595
rect 70977 -22006 71075 -21630
rect 71075 -22006 71142 -21630
rect 71142 -22006 71255 -21630
rect 70977 -22269 71255 -22006
rect 72072 -22012 72165 -21646
rect 72165 -22012 72232 -21646
rect 72232 -22012 72350 -21646
rect 72072 -22285 72350 -22012
rect 73160 -22012 73253 -21646
rect 73253 -22012 73320 -21646
rect 73320 -22012 73438 -21646
rect 73160 -22285 73438 -22012
rect 74248 -22012 74341 -21646
rect 74341 -22012 74408 -21646
rect 74408 -22012 74526 -21646
rect 74248 -22285 74526 -22012
rect 75336 -22012 75429 -21646
rect 75429 -22012 75496 -21646
rect 75496 -22012 75614 -21646
rect 75336 -22285 75614 -22012
rect 76424 -22012 76517 -21646
rect 76517 -22012 76584 -21646
rect 76584 -22012 76702 -21646
rect 76424 -22285 76702 -22012
rect 77512 -22012 77605 -21646
rect 77605 -22012 77672 -21646
rect 77672 -22012 77790 -21646
rect 77512 -22285 77790 -22012
rect 81864 -22012 81957 -21646
rect 81957 -22012 82024 -21646
rect 82024 -22012 82142 -21646
rect 81864 -22285 82142 -22012
rect 82952 -22012 83045 -21646
rect 83045 -22012 83112 -21646
rect 83112 -22012 83230 -21646
rect 82952 -22285 83230 -22012
rect 84040 -22012 84133 -21646
rect 84133 -22012 84200 -21646
rect 84200 -22012 84318 -21646
rect 84040 -22285 84318 -22012
rect 85128 -22012 85221 -21646
rect 85221 -22012 85288 -21646
rect 85288 -22012 85406 -21646
rect 85128 -22285 85406 -22012
rect 13965 -25295 15965 -24595
rect 13965 -32385 15965 -30385
rect 155830 -25295 157830 -24595
rect 155830 -32385 157830 -30385
rect 159830 84397 161830 86397
rect 159830 73705 161830 74405
rect 159830 65705 161830 66405
rect 159830 57705 161830 58405
rect 159830 49705 161830 50405
rect 159830 41705 161830 42405
rect 159830 33705 161830 34405
rect 159830 25705 161830 26405
rect 159830 17705 161830 18405
rect 159830 9705 161830 10405
rect 159830 1705 161830 2405
rect 159830 -6295 161830 -5595
rect 159830 -14295 161830 -13595
rect 159830 -22295 161830 -21595
rect 159830 -36385 161830 -34385
<< metal5 >>
rect 9941 86397 11989 86421
rect 159806 86397 161854 86421
rect 4703 84397 9965 86397
rect 11965 84397 159830 86397
rect 161830 84397 166970 86397
rect 9941 84373 11989 84397
rect 159806 84373 161854 84397
rect 13941 82397 15989 82421
rect 155806 82397 157854 82421
rect 4703 80397 13965 82397
rect 15965 80397 155830 82397
rect 157830 80397 166970 82397
rect 13941 80373 15989 80397
rect 155806 80373 157854 80397
rect 9941 74405 11989 74429
rect 159806 74405 161854 74429
rect 9941 73705 9965 74405
rect 11965 73705 159830 74405
rect 161830 73705 161854 74405
rect 9941 73681 11989 73705
rect 159806 73681 161854 73705
rect 13941 71405 15989 71429
rect 155806 71405 157854 71429
rect 9941 70705 13965 71405
rect 15965 71366 155830 71405
rect 15965 71348 59673 71366
rect 15965 71345 45313 71348
rect 15965 70751 38260 71345
rect 38585 70754 45313 71345
rect 45638 70772 59673 71348
rect 59998 71355 155830 71366
rect 59998 71347 95977 71355
rect 59998 70772 66822 71347
rect 45638 70754 66822 70772
rect 38585 70753 66822 70754
rect 67147 71341 95977 71347
rect 67147 71340 87678 71341
rect 67147 70753 76822 71340
rect 38585 70751 76822 70753
rect 15965 70746 76822 70751
rect 77147 70747 87678 71340
rect 88003 70761 95977 71341
rect 96302 70761 105317 71355
rect 105642 70761 155830 71355
rect 88003 70747 155830 70761
rect 77147 70746 155830 70747
rect 15965 70705 155830 70746
rect 157830 70705 161854 71405
rect 13941 70681 15989 70705
rect 155806 70681 157854 70705
rect 9941 66405 11989 66429
rect 159806 66405 161854 66429
rect 9941 65705 9965 66405
rect 11965 66378 159830 66405
rect 11965 66343 68212 66378
rect 11965 65749 35087 66343
rect 35412 66339 63595 66343
rect 35412 65749 42108 66339
rect 11965 65745 42108 65749
rect 42433 66331 63595 66339
rect 42433 65745 56492 66331
rect 11965 65737 56492 65745
rect 56817 65749 63595 66331
rect 63920 65784 68212 66343
rect 68537 66351 159830 66378
rect 68537 66350 84508 66351
rect 68537 65784 73661 66350
rect 63920 65756 73661 65784
rect 73986 66345 84508 66350
rect 73986 65756 78180 66345
rect 63920 65751 78180 65756
rect 78505 65757 84508 66345
rect 84833 66341 159830 66351
rect 84833 66155 92753 66341
rect 84833 65835 86984 66155
rect 87304 65835 92753 66155
rect 84833 65757 92753 65835
rect 78505 65751 92753 65757
rect 63920 65749 92753 65751
rect 56817 65747 92753 65749
rect 93078 65747 102093 66341
rect 102418 66198 159830 66341
rect 102418 65878 104659 66198
rect 104979 65878 159830 66198
rect 102418 65747 159830 65878
rect 56817 65737 159830 65747
rect 11965 65705 159830 65737
rect 161830 65705 161854 66405
rect 9941 65681 11989 65705
rect 159806 65681 161854 65705
rect 13941 63405 15989 63429
rect 155806 63405 157854 63429
rect 9941 62705 13965 63405
rect 15965 63348 155830 63405
rect 15965 62754 62881 63348
rect 63206 62754 72881 63348
rect 73206 63217 155830 63348
rect 73206 62897 85069 63217
rect 85389 63202 102723 63217
rect 85389 62897 86409 63202
rect 73206 62882 86409 62897
rect 86729 62897 102723 63202
rect 103043 63202 155830 63217
rect 103043 62897 104063 63202
rect 86729 62882 104063 62897
rect 104383 62882 155830 63202
rect 73206 62754 155830 62882
rect 15965 62705 155830 62754
rect 157830 62705 161854 63405
rect 13941 62681 15989 62705
rect 155806 62681 157854 62705
rect 9941 58405 11989 58429
rect 159806 58405 161854 58429
rect 9941 57705 9965 58405
rect 11965 58218 159830 58405
rect 11965 58201 85531 58218
rect 11965 57881 62949 58201
rect 63269 57881 72949 58201
rect 73269 57898 85531 58201
rect 85851 57898 103185 58218
rect 103505 57898 159830 58218
rect 73269 57881 159830 57898
rect 11965 57705 159830 57881
rect 161830 57705 161854 58405
rect 9941 57681 11989 57705
rect 159806 57681 161854 57705
rect 13941 55405 15989 55429
rect 155806 55405 157854 55429
rect 9941 54705 13965 55405
rect 15965 55229 155830 55405
rect 15965 55221 48072 55229
rect 15965 54901 46028 55221
rect 46348 54909 48072 55221
rect 48392 55228 155830 55229
rect 48392 55217 104844 55228
rect 48392 55213 77657 55217
rect 48392 54909 67678 55213
rect 46348 54901 67678 54909
rect 15965 54893 67678 54901
rect 67998 54897 77657 55213
rect 77977 55196 104844 55217
rect 77977 54897 87209 55196
rect 67998 54893 87209 54897
rect 15965 54876 87209 54893
rect 87529 54908 104844 55196
rect 105164 55220 155830 55228
rect 105164 54908 115401 55220
rect 87529 54900 115401 54908
rect 115721 55208 155830 55220
rect 115721 54900 119915 55208
rect 87529 54888 119915 54900
rect 120235 54888 155830 55208
rect 87529 54876 155830 54888
rect 15965 54705 155830 54876
rect 157830 54705 161854 55405
rect 13941 54681 15989 54705
rect 155806 54681 157854 54705
rect 9941 50405 11989 50429
rect 159806 50405 161854 50429
rect 9941 49705 9965 50405
rect 11965 50370 159830 50405
rect 11965 50368 39437 50370
rect 11965 49739 37392 50368
rect 37636 49741 39437 50368
rect 39681 50310 159830 50370
rect 39681 50269 96360 50310
rect 39681 50200 62820 50269
rect 39681 49880 47393 50200
rect 47713 50169 62820 50200
rect 47713 49880 49430 50169
rect 39681 49849 49430 49880
rect 49750 49849 62820 50169
rect 39681 49801 62820 49849
rect 63349 50266 96360 50269
rect 63349 49946 66106 50266
rect 66426 50265 96360 50266
rect 66426 49946 67927 50265
rect 63349 49945 67927 49946
rect 68247 50254 96360 50265
rect 68247 50252 73214 50254
rect 68247 50250 71438 50252
rect 68247 49945 69624 50250
rect 63349 49930 69624 49945
rect 69944 49932 71438 50250
rect 71758 49934 73214 50252
rect 73534 50250 96360 50254
rect 73534 49934 74999 50250
rect 71758 49932 74999 49934
rect 69944 49930 74999 49932
rect 75319 49930 96360 50250
rect 63349 49801 96360 49930
rect 39681 49764 96360 49801
rect 97880 50272 159830 50310
rect 97880 49952 100630 50272
rect 100950 50271 159830 50272
rect 100950 49952 102451 50271
rect 97880 49951 102451 49952
rect 102771 50260 159830 50271
rect 102771 50258 107738 50260
rect 102771 50256 105962 50258
rect 102771 49951 104148 50256
rect 97880 49936 104148 49951
rect 104468 49938 105962 50256
rect 106282 49940 107738 50258
rect 108058 50256 159830 50260
rect 108058 49940 109523 50256
rect 106282 49938 109523 49940
rect 104468 49936 109523 49938
rect 109843 50228 159830 50256
rect 109843 49936 117310 50228
rect 97880 49908 117310 49936
rect 117630 50227 159830 50228
rect 117630 50212 122091 50227
rect 117630 49908 119717 50212
rect 97880 49892 119717 49908
rect 120037 49907 122091 50212
rect 122411 49907 159830 50227
rect 120037 49892 159830 49907
rect 97880 49764 159830 49892
rect 39681 49741 159830 49764
rect 37636 49739 159830 49741
rect 11965 49705 159830 49739
rect 161830 49705 161854 50405
rect 9941 49681 11989 49705
rect 63915 49699 75867 49705
rect 159806 49681 161854 49705
rect 13941 47405 15989 47429
rect 155806 47405 157854 47429
rect 9941 46705 13965 47405
rect 15965 47379 90710 47405
rect 15965 47283 56046 47379
rect 15965 46963 35841 47283
rect 36161 47223 56046 47283
rect 36161 46963 37944 47223
rect 15965 46903 37944 46963
rect 38264 46903 56046 47223
rect 15965 46741 56046 46903
rect 56330 47368 90710 47379
rect 56330 46779 60427 47368
rect 61558 47358 90710 47368
rect 91072 47377 155830 47405
rect 91072 47358 94914 47377
rect 61558 47320 94914 47358
rect 61558 47220 90796 47320
rect 61558 46900 64064 47220
rect 64384 46900 90796 47220
rect 61558 46782 90796 46900
rect 91108 46794 94914 47320
rect 96166 47226 155830 47377
rect 96166 46906 98588 47226
rect 98908 47216 155830 47226
rect 98908 46906 121194 47216
rect 96166 46896 121194 46906
rect 121514 46896 155830 47216
rect 96166 46794 155830 46896
rect 91108 46782 155830 46794
rect 61558 46779 155830 46782
rect 56330 46741 155830 46779
rect 15965 46705 155830 46741
rect 157830 46705 161854 47405
rect 13941 46681 15989 46705
rect 63915 46699 75867 46705
rect 155806 46681 157854 46705
rect 9941 42405 11989 42429
rect 159806 42405 161854 42429
rect 9941 41705 9965 42405
rect 11965 42342 159830 42405
rect 11965 42335 96466 42342
rect 11965 41731 61951 42335
rect 63172 42237 96466 42335
rect 63172 42213 84128 42237
rect 63172 41893 79732 42213
rect 80052 41893 81727 42213
rect 82047 41917 84128 42213
rect 84448 42229 96466 42237
rect 84448 41917 86270 42229
rect 82047 41909 86270 41917
rect 86590 41909 96466 42229
rect 82047 41893 96466 41909
rect 63172 41738 96466 41893
rect 97687 41738 159830 42342
rect 63172 41731 159830 41738
rect 11965 41705 159830 41731
rect 161830 41705 161854 42405
rect 9941 41681 11989 41705
rect 61878 41698 63242 41705
rect 159806 41681 161854 41705
rect 13941 39405 15989 39429
rect 155806 39405 157854 39429
rect 9941 38705 13965 39405
rect 15965 39378 155830 39405
rect 15965 39357 114709 39378
rect 15965 39337 90794 39357
rect 15965 38752 56068 39337
rect 56350 39207 90794 39337
rect 56350 39205 87754 39207
rect 56350 39193 85841 39205
rect 56350 38873 81530 39193
rect 81850 38885 85841 39193
rect 86161 38887 87754 39205
rect 88074 38887 90794 39207
rect 86161 38885 90794 38887
rect 81850 38873 90794 38885
rect 56350 38752 90794 38873
rect 15965 38748 90794 38752
rect 91103 38748 114709 39357
rect 15965 38737 114709 38748
rect 115008 38737 155830 39378
rect 15965 38705 155830 38737
rect 157830 38705 161854 39405
rect 13941 38681 15989 38705
rect 155806 38681 157854 38705
rect 9941 34405 11989 34429
rect 122927 34405 123262 34408
rect 159806 34405 161854 34429
rect 9941 33705 9965 34405
rect 11965 34384 159830 34405
rect 11965 34291 122951 34384
rect 11965 34224 96846 34291
rect 11965 33904 70278 34224
rect 70598 33904 96846 34224
rect 11965 33763 96846 33904
rect 97601 34198 122951 34291
rect 97601 33878 104794 34198
rect 105114 33878 122951 34198
rect 97601 33763 122951 33878
rect 11965 33723 122951 33763
rect 123238 34341 159830 34384
rect 123238 34131 127109 34341
rect 123238 33811 125028 34131
rect 125348 33811 127109 34131
rect 123238 33771 127109 33811
rect 127757 33771 159830 34341
rect 123238 33723 159830 33771
rect 11965 33705 159830 33723
rect 161830 33705 161854 34405
rect 9941 33681 11989 33705
rect 122927 33699 123262 33705
rect 159806 33681 161854 33705
rect 13941 31405 15989 31429
rect 155806 31405 157854 31429
rect 9941 30705 13965 31405
rect 15965 31367 155830 31405
rect 15965 31354 114716 31367
rect 15965 30754 55952 31354
rect 56299 31270 114716 31354
rect 56299 31176 90805 31270
rect 56299 30856 60380 31176
rect 60700 31125 90805 31176
rect 60700 30856 64089 31125
rect 56299 30805 64089 30856
rect 64409 30813 90805 31125
rect 91089 31246 114716 31270
rect 91089 30813 95427 31246
rect 64409 30805 95427 30813
rect 56299 30789 95427 30805
rect 95711 31241 114716 31246
rect 95711 30921 98570 31241
rect 98890 30921 114716 31241
rect 95711 30789 114716 30921
rect 56299 30754 114716 30789
rect 15965 30726 114716 30754
rect 115015 31321 155830 31367
rect 115015 31186 127085 31321
rect 115015 30866 124329 31186
rect 124649 30866 127085 31186
rect 115015 30751 127085 30866
rect 127733 30751 155830 31321
rect 115015 30726 155830 30751
rect 15965 30705 155830 30726
rect 157830 30705 161854 31405
rect 13941 30681 15989 30705
rect 114692 30702 115039 30705
rect 155806 30681 157854 30705
rect 9941 26405 11989 26429
rect 159806 26405 161854 26429
rect 9941 25705 9965 26405
rect 11965 26382 49228 26405
rect 50458 26382 159830 26405
rect 11965 26262 159830 26382
rect 11965 26190 62889 26262
rect 11965 26149 50965 26190
rect 11965 25829 41124 26149
rect 41444 25870 50965 26149
rect 51285 25942 62889 26190
rect 63209 26240 159830 26262
rect 63209 26236 106014 26240
rect 63209 26161 82158 26236
rect 63209 25942 71453 26161
rect 51285 25870 71453 25942
rect 41444 25841 71453 25870
rect 71773 25916 82158 26161
rect 82478 26203 106014 26236
rect 82478 25916 85490 26203
rect 71773 25883 85490 25916
rect 85810 26180 106014 26203
rect 85810 25883 91781 26180
rect 71773 25860 91781 25883
rect 92101 25920 106014 26180
rect 106334 25920 159830 26240
rect 92101 25860 159830 25920
rect 71773 25841 159830 25860
rect 41444 25829 159830 25841
rect 11965 25705 159830 25829
rect 161830 25705 161854 26405
rect 9941 25681 11989 25705
rect 159806 25681 161854 25705
rect 13941 23405 15989 23429
rect 155806 23405 157854 23429
rect 9941 22705 13965 23405
rect 15965 23273 155830 23405
rect 15965 23253 60960 23273
rect 15965 23204 43335 23253
rect 15965 22884 37537 23204
rect 37857 23201 43335 23204
rect 37857 22884 40296 23201
rect 15965 22881 40296 22884
rect 40616 22933 43335 23201
rect 43655 23197 60960 23253
rect 43655 22933 51843 23197
rect 40616 22881 51843 22933
rect 15965 22877 51843 22881
rect 52163 22953 60960 23197
rect 61280 23231 155830 23273
rect 61280 23177 68285 23231
rect 61280 22953 63763 23177
rect 52163 22877 63763 22953
rect 15965 22857 63763 22877
rect 64083 22911 68285 23177
rect 68605 23225 155830 23231
rect 68605 23221 82956 23225
rect 68605 22911 72334 23221
rect 64083 22901 72334 22911
rect 72654 23195 82956 23221
rect 72654 22901 73465 23195
rect 64083 22875 73465 22901
rect 73785 22905 82956 23195
rect 83276 23220 155830 23225
rect 83276 22905 86276 23220
rect 73785 22900 86276 22905
rect 86596 23214 155830 23220
rect 86596 23209 108903 23214
rect 86596 23205 103333 23209
rect 86596 22900 92488 23205
rect 73785 22885 92488 22900
rect 92808 22889 103333 23205
rect 103653 23177 108903 23209
rect 103653 22889 105710 23177
rect 92808 22885 105710 22889
rect 73785 22875 105710 22885
rect 64083 22857 105710 22875
rect 106030 22894 108903 23177
rect 109223 22894 155830 23214
rect 106030 22857 155830 22894
rect 15965 22705 155830 22857
rect 157830 22705 161854 23405
rect 13941 22681 15989 22705
rect 155806 22681 157854 22705
rect 9941 18405 11989 18429
rect 159806 18405 161854 18429
rect 9941 17705 9965 18405
rect 11965 18238 159830 18405
rect 11965 18233 85530 18238
rect 11965 18205 60138 18233
rect 11965 18197 44165 18205
rect 11965 18194 40301 18197
rect 11965 17874 36730 18194
rect 37050 17877 40301 18194
rect 40621 17885 44165 18197
rect 44485 18161 60138 18205
rect 44485 18146 51003 18161
rect 44485 17885 47699 18146
rect 40621 17877 47699 17885
rect 37050 17874 47699 17877
rect 11965 17826 47699 17874
rect 48019 17841 51003 18146
rect 51323 17913 60138 18161
rect 60458 18215 85530 18233
rect 60458 17913 62915 18215
rect 51323 17895 62915 17913
rect 63235 18200 85530 18215
rect 63235 17895 66546 18200
rect 51323 17880 66546 17895
rect 66866 18190 85530 18200
rect 66866 17880 71485 18190
rect 51323 17870 71485 17880
rect 71805 18171 85530 18190
rect 71805 18144 82202 18171
rect 71805 17870 75174 18144
rect 51323 17841 75174 17870
rect 48019 17826 75174 17841
rect 11965 17824 75174 17826
rect 75494 17851 82202 18144
rect 82522 17918 85530 18171
rect 85850 18163 159830 18238
rect 85850 17918 91758 18163
rect 82522 17851 91758 17918
rect 75494 17843 91758 17851
rect 92078 17843 159830 18163
rect 75494 17824 159830 17843
rect 11965 17705 159830 17824
rect 161830 17705 161854 18405
rect 9941 17681 11989 17705
rect 159806 17681 161854 17705
rect 13941 15405 15989 15429
rect 155806 15405 157854 15429
rect 9941 14705 13965 15405
rect 15965 15246 155830 15405
rect 15965 15209 63725 15246
rect 15965 14889 41115 15209
rect 41435 15195 63725 15209
rect 41435 15172 51720 15195
rect 41435 14889 48507 15172
rect 15965 14852 48507 14889
rect 48827 14875 51720 15172
rect 52040 14926 63725 15195
rect 64045 15235 155830 15246
rect 64045 15215 92465 15235
rect 64045 15191 82870 15215
rect 64045 14926 72194 15191
rect 52040 14875 72194 14926
rect 48827 14871 72194 14875
rect 72514 14895 82870 15191
rect 83190 15188 92465 15215
rect 83190 14895 86312 15188
rect 72514 14871 86312 14895
rect 48827 14868 86312 14871
rect 86632 14915 92465 15188
rect 92785 14915 155830 15235
rect 86632 14868 155830 14915
rect 48827 14852 155830 14868
rect 15965 14705 155830 14852
rect 157830 14705 161854 15405
rect 13941 14681 15989 14705
rect 155806 14681 157854 14705
rect 9941 10405 11989 10429
rect 159806 10405 161854 10429
rect 9941 9705 9965 10405
rect 11965 9705 159830 10405
rect 161830 9705 161854 10405
rect 9941 9681 11989 9705
rect 159806 9681 161854 9705
rect 13941 7405 15989 7429
rect 155806 7405 157854 7429
rect 9941 6705 13965 7405
rect 15965 6705 155830 7405
rect 157830 6705 161854 7405
rect 13941 6681 15989 6705
rect 155806 6681 157854 6705
rect 9941 2405 11989 2429
rect 159806 2405 161854 2429
rect 9941 1705 9965 2405
rect 11965 2335 159830 2405
rect 11965 1776 135364 2335
rect 135912 1776 159830 2335
rect 11965 1705 159830 1776
rect 161830 1705 161854 2405
rect 9941 1681 11989 1705
rect 159806 1681 161854 1705
rect 13941 -595 15989 -571
rect 155806 -595 157854 -571
rect 9941 -1295 13965 -595
rect 15965 -627 155830 -595
rect 15965 -1266 67007 -627
rect 67285 -651 155830 -627
rect 67285 -1210 139036 -651
rect 139584 -1210 155830 -651
rect 67285 -1266 155830 -1210
rect 15965 -1295 155830 -1266
rect 157830 -1295 161854 -595
rect 13941 -1319 15989 -1295
rect 155806 -1319 157854 -1295
rect 9941 -5595 11989 -5571
rect 159806 -5595 161854 -5571
rect 9941 -6295 9965 -5595
rect 11965 -5628 159830 -5595
rect 11965 -6267 66477 -5628
rect 66755 -5644 159830 -5628
rect 66755 -6267 70975 -5644
rect 11965 -6283 70975 -6267
rect 71253 -6283 74239 -5644
rect 74517 -6283 77503 -5644
rect 77781 -6283 78591 -5644
rect 78869 -6283 81855 -5644
rect 82133 -6283 85119 -5644
rect 85397 -5678 159830 -5644
rect 85397 -5686 147296 -5678
rect 85397 -6234 135364 -5686
rect 135912 -6226 147296 -5686
rect 147844 -6226 159830 -5678
rect 135912 -6234 159830 -6226
rect 85397 -6283 159830 -6234
rect 11965 -6295 159830 -6283
rect 161830 -6295 161854 -5595
rect 9941 -6319 11989 -6295
rect 70951 -6307 71277 -6295
rect 74215 -6307 74541 -6295
rect 77479 -6307 77805 -6295
rect 78567 -6307 78893 -6295
rect 81831 -6307 82157 -6295
rect 85095 -6307 85421 -6295
rect 159806 -6319 161854 -6295
rect 13941 -8595 15989 -8571
rect 155806 -8595 157854 -8571
rect 9941 -9295 13965 -8595
rect 15965 -8630 155830 -8595
rect 15965 -9269 71521 -8630
rect 71799 -9269 72609 -8630
rect 72887 -9269 73697 -8630
rect 73975 -9269 74785 -8630
rect 75063 -9269 75873 -8630
rect 76151 -9269 76961 -8630
rect 77239 -9269 78049 -8630
rect 78327 -9269 79137 -8630
rect 79415 -9269 80225 -8630
rect 80503 -9269 81313 -8630
rect 81591 -9269 82401 -8630
rect 82679 -9269 83489 -8630
rect 83767 -9269 84577 -8630
rect 84855 -8668 155830 -8630
rect 84855 -9216 150970 -8668
rect 151518 -9216 155830 -8668
rect 84855 -9269 155830 -9216
rect 15965 -9295 155830 -9269
rect 157830 -9295 161854 -8595
rect 13941 -9319 15989 -9295
rect 155806 -9319 157854 -9295
rect 9941 -13595 11989 -13571
rect 159806 -13595 161854 -13571
rect 9941 -14295 9965 -13595
rect 11965 -13629 159830 -13595
rect 11965 -14268 70961 -13629
rect 71239 -14268 72064 -13629
rect 72342 -14268 73137 -13629
rect 73415 -14268 74225 -13629
rect 74503 -14268 75313 -13629
rect 75591 -14268 76401 -13629
rect 76679 -14268 77489 -13629
rect 77767 -14268 78577 -13629
rect 78855 -14268 79665 -13629
rect 79943 -14268 80753 -13629
rect 81031 -14268 81841 -13629
rect 82119 -14268 82929 -13629
rect 83207 -14268 84017 -13629
rect 84295 -14268 85105 -13629
rect 85383 -14268 159830 -13629
rect 11965 -14295 159830 -14268
rect 161830 -14295 161854 -13595
rect 9941 -14319 11989 -14295
rect 159806 -14319 161854 -14295
rect 13941 -16595 15989 -16571
rect 155806 -16595 157854 -16571
rect 9941 -17295 13965 -16595
rect 15965 -16625 155830 -16595
rect 15965 -17264 71519 -16625
rect 71797 -17264 72607 -16625
rect 72885 -17264 73695 -16625
rect 73973 -17264 74783 -16625
rect 75061 -17264 75871 -16625
rect 76149 -17264 76959 -16625
rect 77237 -17264 78047 -16625
rect 78325 -17264 79135 -16625
rect 79413 -17264 80223 -16625
rect 80501 -17264 81311 -16625
rect 81589 -17264 82399 -16625
rect 82677 -17264 83487 -16625
rect 83765 -17264 84575 -16625
rect 84853 -17264 155830 -16625
rect 15965 -17295 155830 -17264
rect 157830 -17295 161854 -16595
rect 13941 -17319 15989 -17295
rect 155806 -17319 157854 -17295
rect 9941 -21595 11989 -21571
rect 159806 -21595 161854 -21571
rect 9941 -22295 9965 -21595
rect 11965 -21630 159830 -21595
rect 11965 -22269 70977 -21630
rect 71255 -21646 159830 -21630
rect 71255 -22269 72072 -21646
rect 11965 -22285 72072 -22269
rect 72350 -22285 73160 -21646
rect 73438 -22285 74248 -21646
rect 74526 -22285 75336 -21646
rect 75614 -22285 76424 -21646
rect 76702 -22285 77512 -21646
rect 77790 -22285 81864 -21646
rect 82142 -22285 82952 -21646
rect 83230 -22285 84040 -21646
rect 84318 -22285 85128 -21646
rect 85406 -22285 159830 -21646
rect 11965 -22295 159830 -22285
rect 161830 -22295 161854 -21595
rect 9941 -22319 11989 -22295
rect 72048 -22309 72374 -22295
rect 73136 -22309 73462 -22295
rect 74224 -22309 74550 -22295
rect 75312 -22309 75638 -22295
rect 76400 -22309 76726 -22295
rect 77488 -22309 77814 -22295
rect 81840 -22309 82166 -22295
rect 82928 -22309 83254 -22295
rect 84016 -22309 84342 -22295
rect 85104 -22309 85430 -22295
rect 159806 -22319 161854 -22295
rect 13941 -24595 15989 -24571
rect 155806 -24595 157854 -24571
rect 9941 -25295 13965 -24595
rect 15965 -25295 155830 -24595
rect 157830 -25295 161854 -24595
rect 13941 -25319 15989 -25295
rect 155806 -25319 157854 -25295
rect 13941 -30385 15989 -30361
rect 155806 -30385 157854 -30361
rect 4703 -32385 13965 -30385
rect 15965 -32385 155830 -30385
rect 157830 -32385 166970 -30385
rect 13941 -32409 15989 -32385
rect 155806 -32409 157854 -32385
rect 9941 -34385 11989 -34361
rect 159806 -34385 161854 -34361
rect 4703 -36385 9965 -34385
rect 11965 -36385 159830 -34385
rect 161830 -36385 166970 -34385
rect 9941 -36409 11989 -36385
rect 159806 -36409 161854 -36385
use a_mux2_en  a_mux2_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/a_mux2_en
timestamp 1655484843
transform 0 -1 84928 1 0 60716
box -2638 -2806 3466 243
use a_mux2_en  a_mux2_en_1
timestamp 1655484843
transform 0 -1 102582 1 0 60716
box -2638 -2806 3466 243
use a_mux4_en  a_mux4_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/a_mux4_en
timestamp 1655484843
transform 0 -1 62720 1 0 61957
box -3843 -5692 3675 352
use a_mux4_en  a_mux4_en_1
timestamp 1655484843
transform 0 -1 72720 1 0 61957
box -3843 -5692 3675 352
use clock_v2  clock_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/clock_v2
timestamp 1655484843
transform 0 -1 71097 1 0 -19032
box -3377 -14204 17044 36
use comparator_v2  comparator_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/comparator_v2
timestamp 1655484843
transform 0 1 115004 1 0 32246
box -3788 -193 7250 10729
use esd_cell  esd_cell_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/esd_cell
timestamp 1655484843
transform 0 -1 66871 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_1
timestamp 1655484843
transform 0 -1 76871 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_2
timestamp 1655484843
transform 0 -1 87741 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_3
timestamp 1655484843
transform 0 -1 105391 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_4
timestamp 1655484843
transform 0 -1 59771 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_5
timestamp 1655484843
transform 0 -1 96051 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_6
timestamp 1655484843
transform 0 -1 45351 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_7
timestamp 1655484843
transform 0 -1 38351 1 0 67009
box -64 -64 3554 3096
use onebit_dac  onebit_dac_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/onebit_dac
timestamp 1655484843
transform 0 1 116581 1 0 50758
box -6 -1274 1554 1238
use onebit_dac  onebit_dac_1
timestamp 1655484843
transform 0 1 120581 1 0 50758
box -6 -1274 1554 1238
use ota_v2  ota_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/ota_v2
timestamp 1655484843
transform 0 1 90907 1 0 28504
box -170 1 23753 20628
use ota_w_test_v2  ota_w_test_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/ota_w_test_v2
timestamp 1655484843
transform 0 1 56391 1 0 28511
box -170 1 23753 20628
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/analog_top_v2
timestamp 1655484843
transform 1 0 80428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_1
timestamp 1655484843
transform 1 0 82428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_2
timestamp 1655484843
transform 1 0 81428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_3
timestamp 1655484843
transform 1 0 83428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_4
timestamp 1655484843
transform -1 0 87328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_5
timestamp 1655484843
transform -1 0 87328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_6
timestamp 1655484843
transform -1 0 86328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_7
timestamp 1655484843
transform -1 0 86328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_8
timestamp 1655484843
transform -1 0 85328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_9
timestamp 1655484843
transform 1 0 81428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_10
timestamp 1655484843
transform 1 0 82428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_11
timestamp 1655484843
transform 1 0 83428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_12
timestamp 1655484843
transform -1 0 85328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_13
timestamp 1655484843
transform -1 0 84328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_14
timestamp 1655484843
transform -1 0 84328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_15
timestamp 1655484843
transform 1 0 80428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_16
timestamp 1655484843
transform 1 0 80428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_17
timestamp 1655484843
transform 1 0 81428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_18
timestamp 1655484843
transform 1 0 82428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_19
timestamp 1655484843
transform 1 0 83428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_20
timestamp 1655484843
transform -1 0 87328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_21
timestamp 1655484843
transform -1 0 87328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_22
timestamp 1655484843
transform -1 0 86328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_23
timestamp 1655484843
transform -1 0 86328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_24
timestamp 1655484843
transform 1 0 80428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_25
timestamp 1655484843
transform 1 0 81428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_26
timestamp 1655484843
transform 1 0 82428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_27
timestamp 1655484843
transform 1 0 83428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_28
timestamp 1655484843
transform -1 0 85328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_29
timestamp 1655484843
transform -1 0 85328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_30
timestamp 1655484843
transform -1 0 84328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_31
timestamp 1655484843
transform -1 0 84328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_32
timestamp 1655484843
transform 1 0 80428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_33
timestamp 1655484843
transform 1 0 81428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_34
timestamp 1655484843
transform 1 0 82428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_35
timestamp 1655484843
transform 1 0 83428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_36
timestamp 1655484843
transform -1 0 87328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_37
timestamp 1655484843
transform -1 0 86328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_38
timestamp 1655484843
transform -1 0 85328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_39
timestamp 1655484843
transform -1 0 84328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_40
timestamp 1655484843
transform 1 0 80428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_41
timestamp 1655484843
transform 1 0 81428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_42
timestamp 1655484843
transform 1 0 82428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_43
timestamp 1655484843
transform 1 0 83428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_44
timestamp 1655484843
transform -1 0 87328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_45
timestamp 1655484843
transform -1 0 87328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_46
timestamp 1655484843
transform -1 0 86328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_47
timestamp 1655484843
transform -1 0 86328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_48
timestamp 1655484843
transform 1 0 80428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_49
timestamp 1655484843
transform 1 0 81428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_50
timestamp 1655484843
transform 1 0 82428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_51
timestamp 1655484843
transform 1 0 83428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_52
timestamp 1655484843
transform -1 0 85328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_53
timestamp 1655484843
transform -1 0 85328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_54
timestamp 1655484843
transform -1 0 84328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_55
timestamp 1655484843
transform -1 0 84328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_56
timestamp 1655484843
transform 1 0 80428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_57
timestamp 1655484843
transform 1 0 81428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_58
timestamp 1655484843
transform 1 0 82428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_59
timestamp 1655484843
transform 1 0 83428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_60
timestamp 1655484843
transform -1 0 87328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_61
timestamp 1655484843
transform -1 0 87328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_62
timestamp 1655484843
transform -1 0 86328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_63
timestamp 1655484843
transform -1 0 86328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_64
timestamp 1655484843
transform 1 0 80428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_65
timestamp 1655484843
transform 1 0 81428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_66
timestamp 1655484843
transform 1 0 82428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_67
timestamp 1655484843
transform 1 0 83428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_68
timestamp 1655484843
transform -1 0 85328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_69
timestamp 1655484843
transform -1 0 85328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_70
timestamp 1655484843
transform -1 0 84328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_71
timestamp 1655484843
transform -1 0 84328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/analog_top_v2
timestamp 1655484843
transform 0 -1 39165 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_1
timestamp 1655484843
transform 0 -1 39165 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_2
timestamp 1655484843
transform 0 -1 39165 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_3
timestamp 1655484843
transform 0 -1 39165 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_4
timestamp 1655484843
transform 0 -1 39165 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_5
timestamp 1655484843
transform 0 -1 39165 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_6
timestamp 1655484843
transform 0 -1 35965 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_7
timestamp 1655484843
transform 0 -1 35965 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_8
timestamp 1655484843
transform 0 -1 35965 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_9
timestamp 1655484843
transform 0 -1 35965 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_10
timestamp 1655484843
transform 0 -1 35965 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_11
timestamp 1655484843
transform 0 -1 35965 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_12
timestamp 1655484843
transform 0 -1 32765 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_13
timestamp 1655484843
transform 0 -1 32765 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_14
timestamp 1655484843
transform 0 -1 32765 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_15
timestamp 1655484843
transform 0 -1 32765 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_16
timestamp 1655484843
transform 0 -1 32765 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_17
timestamp 1655484843
transform 0 -1 32765 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_18
timestamp 1655484843
transform 0 -1 29565 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_19
timestamp 1655484843
transform 0 -1 29565 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_20
timestamp 1655484843
transform 0 -1 29565 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_21
timestamp 1655484843
transform 0 -1 29565 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_22
timestamp 1655484843
transform 0 -1 29565 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_23
timestamp 1655484843
transform 0 -1 29565 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_24
timestamp 1655484843
transform 0 1 42365 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_25
timestamp 1655484843
transform 0 1 42365 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_26
timestamp 1655484843
transform 0 1 42365 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_27
timestamp 1655484843
transform 0 1 42365 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_28
timestamp 1655484843
transform 0 1 42365 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_29
timestamp 1655484843
transform 0 1 42365 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_30
timestamp 1655484843
transform 0 1 45565 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_31
timestamp 1655484843
transform 0 1 45565 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_32
timestamp 1655484843
transform 0 1 45565 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_33
timestamp 1655484843
transform 0 1 45565 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_34
timestamp 1655484843
transform 0 1 45565 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_35
timestamp 1655484843
transform 0 1 45565 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_36
timestamp 1655484843
transform 0 1 48765 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_37
timestamp 1655484843
transform 0 1 48765 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_38
timestamp 1655484843
transform 0 1 48765 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_39
timestamp 1655484843
transform 0 1 48765 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_40
timestamp 1655484843
transform 0 1 48765 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_41
timestamp 1655484843
transform 0 1 48765 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_42
timestamp 1655484843
transform 0 1 51965 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_43
timestamp 1655484843
transform 0 1 51965 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_44
timestamp 1655484843
transform 0 1 51965 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_45
timestamp 1655484843
transform 0 1 51965 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_46
timestamp 1655484843
transform 0 1 51965 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_47
timestamp 1655484843
transform 0 1 51965 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/analog_top_v2
timestamp 1655484843
transform 0 1 108064 -1 0 25313
box -1310 -1260 1210 1260
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_1
timestamp 1655484843
transform 0 1 104396 -1 0 25315
box -1310 -1260 1210 1260
use sky130_fd_pr__nfet_01v8_CFEPS5  sky130_fd_pr__nfet_01v8_CFEPS5_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/analog_top_v2
timestamp 1655484843
transform 1 0 127406 0 -1 32821
box -311 -274 311 276
use sky130_fd_pr__pfet_01v8_hvt_XAYTAL  sky130_fd_pr__pfet_01v8_hvt_XAYTAL_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/analog_top_v2
timestamp 1655484843
transform 1 0 127406 0 -1 33415
box -311 -319 311 319
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 136247 0 1 -3507
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1655484843
transform 1 0 136247 0 1 -1860
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_2
timestamp 1655484843
transform 1 0 136247 0 1 -543
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_3
timestamp 1655484843
transform 1 0 136247 0 1 -4754
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_4
timestamp 1655484843
transform 1 0 148179 0 1 -11735
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 0 -1 67137 1 0 -5429
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1655484843
transform 1 0 138179 0 1 -3507
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_2
timestamp 1655484843
transform 1 0 138179 0 1 -1860
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_3
timestamp 1655484843
transform 1 0 138179 0 1 -543
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_4
timestamp 1655484843
transform 1 0 138179 0 1 -4754
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_5
timestamp 1655484843
transform 1 0 150111 0 1 -11735
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 0 -1 67137 1 0 -6625
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1655484843
transform 0 -1 67137 1 0 -3129
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_2
timestamp 1655484843
transform 1 0 136983 0 1 -3507
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_3
timestamp 1655484843
transform 1 0 135051 0 1 -3507
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_4
timestamp 1655484843
transform 1 0 140479 0 1 -3507
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_5
timestamp 1655484843
transform 1 0 140479 0 1 -1860
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_6
timestamp 1655484843
transform 1 0 136983 0 1 -1860
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_7
timestamp 1655484843
transform 1 0 135051 0 1 -1860
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_8
timestamp 1655484843
transform 1 0 140479 0 1 -543
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_9
timestamp 1655484843
transform 1 0 136983 0 1 -543
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_10
timestamp 1655484843
transform 1 0 135051 0 1 -543
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_11
timestamp 1655484843
transform 1 0 135051 0 1 -4754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_12
timestamp 1655484843
transform 1 0 136983 0 1 -4754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_13
timestamp 1655484843
transform 1 0 140479 0 1 -4754
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_14
timestamp 1655484843
transform 1 0 152411 0 1 -11735
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_15
timestamp 1655484843
transform 1 0 148915 0 1 -11735
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_16
timestamp 1655484843
transform 1 0 146983 0 1 -11735
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 133119 0 1 -3507
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_1
timestamp 1655484843
transform 1 0 133119 0 1 -1860
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_2
timestamp 1655484843
transform 1 0 133119 0 1 -543
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_3
timestamp 1655484843
transform 1 0 133119 0 1 -4754
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_4
timestamp 1655484843
transform 1 0 145051 0 1 -11735
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 0 -1 67137 1 0 -5521
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1655484843
transform 0 -1 67137 1 0 -3221
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1655484843
transform 1 0 136891 0 1 -3507
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1655484843
transform 1 0 136155 0 1 -3507
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1655484843
transform 1 0 133027 0 1 -3507
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1655484843
transform 1 0 140387 0 1 -3507
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1655484843
transform 1 0 138087 0 1 -3507
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1655484843
transform 1 0 140387 0 1 -1860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1655484843
transform 1 0 138087 0 1 -1860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1655484843
transform 1 0 136891 0 1 -1860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1655484843
transform 1 0 136155 0 1 -1860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1655484843
transform 1 0 133027 0 1 -1860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1655484843
transform 1 0 140387 0 1 -543
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1655484843
transform 1 0 138087 0 1 -543
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1655484843
transform 1 0 136891 0 1 -543
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1655484843
transform 1 0 136155 0 1 -543
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1655484843
transform 1 0 133027 0 1 -543
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1655484843
transform 1 0 133027 0 1 -4754
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1655484843
transform 1 0 136155 0 1 -4754
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1655484843
transform 1 0 136891 0 1 -4754
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1655484843
transform 1 0 138087 0 1 -4754
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1655484843
transform 1 0 140387 0 1 -4754
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1655484843
transform 1 0 152319 0 1 -11735
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1655484843
transform 1 0 150019 0 1 -11735
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1655484843
transform 1 0 148823 0 1 -11735
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1655484843
transform 1 0 148087 0 1 -11735
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1655484843
transform 1 0 144959 0 1 -11735
box -38 -48 130 592
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/transmission_gate
timestamp 1655484843
transform 1 0 50965 0 1 22637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_1
timestamp 1655484843
transform 1 0 47655 0 1 20637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_2
timestamp 1655484843
transform 1 0 47655 0 1 18637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_3
timestamp 1655484843
transform 1 0 50965 0 1 16637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_4
timestamp 1655484843
transform 1 0 40287 0 1 22642
box -53 -49 1241 1063
use transmission_gate  transmission_gate_5
timestamp 1655484843
transform 1 0 40287 0 1 16642
box -53 -49 1241 1063
use transmission_gate  transmission_gate_6
timestamp 1655484843
transform -1 0 44518 0 -1 21462
box -53 -49 1241 1063
use transmission_gate  transmission_gate_7
timestamp 1655484843
transform -1 0 44518 0 -1 19462
box -53 -49 1241 1063
use transmission_gate  transmission_gate_8
timestamp 1655484843
transform 1 0 36712 0 1 20644
box -53 -49 1241 1063
use transmission_gate  transmission_gate_9
timestamp 1655484843
transform 1 0 36712 0 1 18644
box -53 -49 1241 1063
use transmission_gate  transmission_gate_10
timestamp 1655484843
transform 0 1 36343 -1 0 50351
box -53 -49 1241 1063
use transmission_gate  transmission_gate_11
timestamp 1655484843
transform 0 1 38343 -1 0 50351
box -53 -49 1241 1063
use transmission_gate  transmission_gate_12
timestamp 1655484843
transform 1 0 60175 0 1 18637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_13
timestamp 1655484843
transform 1 0 62895 0 1 16637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_14
timestamp 1655484843
transform 1 0 62895 0 1 22637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_15
timestamp 1655484843
transform 1 0 60175 0 1 20637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_16
timestamp 1655484843
transform 0 -1 68108 1 0 19681
box -53 -49 1241 1063
use transmission_gate  transmission_gate_17
timestamp 1655484843
transform 0 -1 85714 -1 0 43032
box -53 -49 1241 1063
use transmission_gate  transmission_gate_18
timestamp 1655484843
transform 0 -1 87714 -1 0 43032
box -53 -49 1241 1063
use transmission_gate  transmission_gate_19
timestamp 1655484843
transform 1 0 71459 0 1 22638
box -53 -49 1241 1063
use transmission_gate  transmission_gate_20
timestamp 1655484843
transform 1 0 71459 0 1 16648
box -53 -49 1241 1063
use transmission_gate  transmission_gate_21
timestamp 1655484843
transform 0 1 73976 1 0 19436
box -53 -49 1241 1063
use transmission_gate  transmission_gate_22
timestamp 1655484843
transform 1 0 85498 0 -1 16775
box -53 -49 1241 1063
use transmission_gate  transmission_gate_23
timestamp 1655484843
transform 1 0 82138 0 -1 17625
box -53 -49 1241 1063
use transmission_gate  transmission_gate_24
timestamp 1655484843
transform 1 0 82138 0 -1 23595
box -53 -49 1241 1063
use transmission_gate  transmission_gate_25
timestamp 1655484843
transform 1 0 85498 0 -1 24785
box -53 -49 1241 1063
use transmission_gate  transmission_gate_26
timestamp 1655484843
transform -1 0 92927 0 -1 23595
box -53 -49 1241 1063
use transmission_gate  transmission_gate_27
timestamp 1655484843
transform -1 0 92927 0 -1 17625
box -53 -49 1241 1063
use transmission_gate  transmission_gate_28
timestamp 1655484843
transform -1 0 106850 0 1 22217
box -53 -49 1241 1063
use transmission_gate  transmission_gate_29
timestamp 1655484843
transform 0 -1 83121 -1 0 41228
box -53 -49 1241 1063
use transmission_gate  transmission_gate_30
timestamp 1655484843
transform 0 -1 81121 -1 0 41228
box -53 -49 1241 1063
use transmission_gate  transmission_gate_31
timestamp 1655484843
transform 0 1 48389 -1 0 52358
box -53 -49 1241 1063
use transmission_gate  transmission_gate_32
timestamp 1655484843
transform 0 1 46389 -1 0 52348
box -53 -49 1241 1063
<< labels >>
flabel metal3 166522 7170 166522 7170 1 FreeSans 8000 0 0 0 d_clk_grp_2_ctrl_0
port 21 n
flabel metal3 166482 5138 166482 5138 1 FreeSans 8000 0 0 0 d_clk_grp_2_ctrl_1
port 22 n
flabel metal3 166471 -867 166471 -867 1 FreeSans 8000 0 0 0 d_clk_grp_1_ctrl_0
port 19 n
flabel metal3 166471 -2775 166471 -2775 1 FreeSans 8000 0 0 0 d_clk_grp_1_ctrl_1
port 20 n
flabel metal3 67147 -40491 67147 -40491 1 FreeSans 8000 0 0 0 rst_n
port 3 n
flabel metal3 77988 -40479 77988 -40479 1 FreeSans 8000 0 0 0 clk
port 14 n
flabel metal3 117368 90901 117368 90901 1 FreeSans 8000 0 0 0 debug
port 8 n
flabel metal3 115397 89837 115397 89837 1 FreeSans 8000 0 0 0 a_mod_grp_ctrl_1
port 7 n
flabel metal3 113347 88615 113347 88615 1 FreeSans 8000 0 0 0 a_mod_grp_ctrl_0
port 6 n
flabel metal3 103942 90507 103942 90507 1 FreeSans 8000 0 0 0 a_probe_1
port 11 n
flabel metal3 86275 90560 86275 90560 1 FreeSans 8000 0 0 0 a_probe_0
port 10 n
flabel metal3 94580 90666 94580 90666 1 FreeSans 8000 0 0 0 i_bias_2
port 5 n
flabel metal3 75485 90718 75485 90718 1 FreeSans 8000 0 0 0 a_probe_3
port 13 n
flabel metal3 65329 90613 65329 90613 1 FreeSans 8000 0 0 0 a_probe_2
port 12 n
flabel metal3 58241 90613 58241 90613 1 FreeSans 8000 0 0 0 i_bias_1
port 4 n
flabel metal3 36925 90771 36925 90771 1 FreeSans 8000 0 0 0 ip
port 1 n
flabel metal3 43854 90771 43854 90771 1 FreeSans 8000 0 0 0 in
port 2 n
flabel metal5 5498 85359 5498 85359 1 FreeSans 8000 0 0 0 VDD
port 23 n power bidirectional
flabel metal5 5307 81285 5307 81285 1 FreeSans 8000 0 0 0 VSS
port 24 n power bidirectional
flabel metal3 166446 34396 166446 34396 1 FreeSans 8000 0 0 0 op
port 9 n
flabel metal3 166538 -10922 166538 -10922 1 FreeSans 8000 0 0 0 d_probe
port 25 n
flabel metal3 166388 -12956 166388 -12956 1 FreeSans 8000 0 0 0 d_probe_ctrl_0
port 26 n
flabel metal3 166388 -15258 166388 -15258 1 FreeSans 8000 0 0 0 d_probe_ctrl_1
port 27 n
<< end >>
