magic
tech sky130A
timestamp 1654711401
<< error_p >>
rect -38 90 -9 93
rect 9 90 38 93
rect -38 73 -32 90
rect 9 73 15 90
rect -38 70 -9 73
rect 9 70 38 73
rect -38 -73 -9 -70
rect 9 -73 38 -70
rect -38 -90 -32 -73
rect 9 -90 15 -73
rect -38 -93 -9 -90
rect 9 -93 38 -90
<< nwell >>
rect -155 -159 155 159
<< pmoshvt >>
rect -55 -50 -40 50
rect -7 -50 7 50
rect 40 -50 55 50
<< pdiff >>
rect -86 44 -55 50
rect -86 -44 -80 44
rect -63 -44 -55 44
rect -86 -50 -55 -44
rect -40 44 -7 50
rect -40 -44 -32 44
rect -15 -44 -7 44
rect -40 -50 -7 -44
rect 7 44 40 50
rect 7 -44 15 44
rect 32 -44 40 44
rect 7 -50 40 -44
rect 55 44 86 50
rect 55 -44 63 44
rect 80 -44 86 44
rect 55 -50 86 -44
<< pdiffc >>
rect -80 -44 -63 44
rect -32 -44 -15 44
rect 15 -44 32 44
rect 63 -44 80 44
<< nsubdiff >>
rect -137 124 -89 141
rect 89 124 137 141
rect -137 93 -120 124
rect 120 93 137 124
rect -137 -124 -120 -93
rect 120 -124 137 -93
rect -137 -141 -89 -124
rect 89 -141 137 -124
<< nsubdiffcont >>
rect -89 124 89 141
rect -137 -93 -120 93
rect 120 -93 137 93
rect -89 -141 89 -124
<< poly >>
rect -64 90 64 98
rect -64 73 -32 90
rect -15 73 15 90
rect 32 73 64 90
rect -64 63 64 73
rect -55 50 -40 63
rect -7 50 7 63
rect 40 50 55 63
rect -55 -65 -40 -50
rect -7 -65 7 -50
rect 40 -65 55 -50
rect -64 -73 64 -65
rect -64 -90 -32 -73
rect -15 -90 15 -73
rect 32 -90 64 -73
rect -64 -101 64 -90
<< polycont >>
rect -32 73 -15 90
rect 15 73 32 90
rect -32 -90 -15 -73
rect 15 -90 32 -73
<< locali >>
rect -137 124 -89 141
rect 89 124 137 141
rect -137 93 -120 124
rect 120 93 137 124
rect -40 73 -32 90
rect -15 73 15 90
rect 32 73 40 90
rect -80 44 -63 52
rect -80 -52 -63 -44
rect -32 44 -15 52
rect -32 -52 -15 -44
rect 15 44 32 52
rect 15 -52 32 -44
rect 63 44 80 52
rect 63 -52 80 -44
rect -40 -90 -32 -73
rect -15 -90 15 -73
rect 32 -90 40 -73
rect -137 -124 -120 -93
rect 120 -124 137 -93
rect -137 -141 -89 -124
rect 89 -141 137 -124
<< viali >>
rect -32 73 -15 90
rect 15 73 32 90
rect -80 -44 -63 44
rect -32 -44 -15 44
rect 15 -44 32 44
rect 63 -44 80 44
rect -32 -90 -15 -73
rect 15 -90 32 -73
<< metal1 >>
rect -38 90 -9 93
rect -38 73 -32 90
rect -15 73 -9 90
rect -38 70 -9 73
rect 9 90 38 93
rect 9 73 15 90
rect 32 73 38 90
rect 9 70 38 73
rect -83 44 -60 50
rect -83 8 -80 44
rect -137 -8 -80 8
rect -83 -44 -80 -8
rect -63 8 -60 44
rect -35 44 -12 50
rect -35 8 -32 44
rect -63 -8 -32 8
rect -63 -44 -60 -8
rect -83 -50 -60 -44
rect -35 -44 -32 -8
rect -15 8 -12 44
rect 12 44 35 50
rect 12 8 15 44
rect -15 -8 15 8
rect -15 -44 -12 -8
rect -35 -50 -12 -44
rect 12 -44 15 -8
rect 32 8 35 44
rect 60 44 83 50
rect 60 8 63 44
rect 32 -8 63 8
rect 32 -44 35 -8
rect 12 -50 35 -44
rect 60 -44 63 -8
rect 80 -44 83 44
rect 60 -50 83 -44
rect -38 -73 -9 -70
rect -38 -90 -32 -73
rect -15 -90 -9 -73
rect -38 -93 -9 -90
rect 9 -73 38 -70
rect 9 -90 15 -73
rect 32 -90 38 -73
rect 9 -93 38 -90
<< properties >>
string FIXED_BBOX -129 -133 129 133
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 1 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
