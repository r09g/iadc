* NGSPICE file created from a_mux4_en_flat.ext - technology: sky130A

.subckt a_mux4_en_flat en s1 s0 in0 in1 in2 in3 out VDD VSS
X0 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=1.05536e+13p pd=8.08e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X1 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X2 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X3 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X4 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X5 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X6 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X7 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X8 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=0p ps=0u w=1.36e+06u l=150000u
X9 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=4.0352e+12p ps=4.048e+07u w=520000u l=150000u
X10 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X11 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X12 a_n499_n2830# sky130_fd_sc_hd__nand2_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=2.439e+12p ps=2.634e+07u w=650000u l=150000u
X13 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X14 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X15 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X16 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X17 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X18 a_n499_n1742# sky130_fd_sc_hd__nand2_1_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X19 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X20 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X21 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X22 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X23 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X24 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X25 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X26 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X27 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X28 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X29 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X30 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X31 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X32 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X33 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X34 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X35 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X36 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X37 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X38 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X39 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X40 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X41 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X42 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X43 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X44 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X45 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X46 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X47 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X48 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X49 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X50 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X51 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X52 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X53 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X54 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X55 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X56 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__nand2_1_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=3.9e+12p ps=3.78e+07u w=1e+06u l=150000u
X57 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X58 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X59 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X60 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X61 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X62 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X63 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/en_b VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X64 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X65 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X66 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X67 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X68 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X69 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X70 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X71 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X72 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X73 switch_5t_3/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X74 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X75 VDD s0 switch_5t_2/transmission_gate_0/en_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X76 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X77 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X78 switch_5t_3/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X79 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X80 VDD sky130_fd_sc_hd__nand2_1_3/A switch_5t_1/transmission_gate_0/en_b VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X81 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X82 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X83 sky130_fd_sc_hd__nand2_1_0/Y s0 a_n499_n3694# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X84 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X85 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X86 VDD s0 sky130_fd_sc_hd__nand2_1_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X87 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X88 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X89 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X90 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X91 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X92 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X93 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X94 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X95 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X96 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X97 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X98 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X99 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X100 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X101 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X102 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X103 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X104 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X105 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X106 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X107 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X108 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X109 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X110 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X111 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X112 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X113 switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X114 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X115 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X116 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X117 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X118 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X119 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X120 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X121 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X122 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X123 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X124 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X125 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X127 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X129 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X130 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X131 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X132 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X133 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X134 a_n499_n3694# s1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X135 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X136 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X137 sky130_fd_sc_hd__nand2_1_3/B s0 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X138 sky130_fd_sc_hd__nand2_1_0/Y s1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X140 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X141 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X142 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X143 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X144 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X145 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X146 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X147 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X148 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X149 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X150 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X151 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X152 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X153 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X154 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X155 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X156 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X157 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X158 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X159 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X160 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X161 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X162 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X163 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X164 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X165 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X166 transmission_gate_0/en_b en VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X167 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X168 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X169 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X170 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X171 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X172 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X173 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X174 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X175 sky130_fd_sc_hd__nand2_1_3/A s1 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X176 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X177 switch_5t_3/transmission_gate_0/in transmission_gate_0/en_b in3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X178 switch_5t_3/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X179 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X180 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X181 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X182 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X183 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X184 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X185 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X186 in0 transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X187 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X188 out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X189 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X190 switch_5t_0/transmission_gate_0/in en in1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X191 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X192 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X193 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X194 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X195 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X196 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X197 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X198 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X199 in3 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X200 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X201 switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/en_b VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X202 sky130_fd_sc_hd__nand2_1_3/B s0 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X203 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X204 sky130_fd_sc_hd__inv_1_3/A s1 a_n499_n2606# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X205 out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X206 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X207 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X208 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b in0 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X209 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X210 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X211 out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X212 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X213 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X214 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X215 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X216 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X217 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X218 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X219 in1 en switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X220 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X221 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X222 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X223 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X224 out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X225 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X226 out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X227 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X228 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/en_b VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X229 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X230 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X231 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X232 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X233 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X234 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X235 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X236 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X237 in2 transmission_gate_0/en_b switch_5t_2/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X238 switch_5t_2/transmission_gate_0/en_b s0 a_n499_n2830# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X239 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X240 out switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X241 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A a_n499_n1742# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X242 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X243 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X244 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X245 transmission_gate_0/en_b en VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X246 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X247 in3 en switch_5t_3/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X248 switch_5t_1/transmission_gate_0/in en in0 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X249 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X250 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X251 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X252 a_n499_n2606# sky130_fd_sc_hd__nand2_1_3/B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X253 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b in2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X254 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X255 switch_5t_3/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X256 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X257 in1 transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X258 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X259 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/A out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X260 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X261 sky130_fd_sc_hd__nand2_1_3/A s1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X262 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X263 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b in1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X264 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y switch_5t_0/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X265 switch_5t_3/transmission_gate_0/in en in3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X266 switch_5t_2/transmission_gate_0/in en in2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X267 in0 en switch_5t_1/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X268 VDD s1 sky130_fd_sc_hd__inv_1_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X269 out switch_5t_2/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X270 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X271 switch_5t_3/transmission_gate_0/in switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X272 in2 en switch_5t_2/transmission_gate_0/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X273 out switch_5t_1/transmission_gate_0/en switch_5t_1/transmission_gate_0/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 switch_5t_2/transmission_gate_0/in switch_5t_3/transmission_gate_0/out 0.07fF
C1 switch_5t_0/transmission_gate_0/in switch_5t_1/transmission_gate_0/in 0.45fF
C2 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en 1.51fF
C3 s0 en 0.55fF
C4 sky130_fd_sc_hd__inv_1_3/Y switch_5t_1/transmission_gate_0/out 0.09fF
C5 VDD switch_5t_0/transmission_gate_0/in 2.86fF
C6 sky130_fd_sc_hd__inv_1_3/Y switch_5t_1/transmission_gate_0/in 0.12fF
C7 VDD sky130_fd_sc_hd__inv_1_3/Y 0.57fF
C8 switch_5t_0/transmission_gate_0/out switch_5t_0/transmission_gate_0/in 7.36fF
C9 s1 switch_5t_1/transmission_gate_0/en 0.03fF
C10 switch_5t_2/transmission_gate_0/out switch_5t_0/transmission_gate_0/in 0.07fF
C11 sky130_fd_sc_hd__nand2_1_3/B sky130_fd_sc_hd__nand2_1_3/A 0.49fF
C12 transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in 0.49fF
C13 switch_5t_2/transmission_gate_0/in en 0.66fF
C14 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y 1.95fF
C15 switch_5t_2/transmission_gate_0/out sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C16 switch_5t_1/transmission_gate_0/out transmission_gate_0/en_b 0.02fF
C17 switch_5t_1/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in 0.13fF
C18 switch_5t_1/transmission_gate_0/in transmission_gate_0/en_b 0.73fF
C19 sky130_fd_sc_hd__nand2_1_0/Y s0 0.21fF
C20 s0 switch_5t_2/transmission_gate_0/en_b 0.45fF
C21 switch_5t_2/transmission_gate_0/en switch_5t_0/transmission_gate_0/in 0.05fF
C22 VDD transmission_gate_0/en_b 5.66fF
C23 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__inv_1_3/Y 0.67fF
C24 switch_5t_3/transmission_gate_0/en transmission_gate_0/en_b 0.00fF
C25 switch_5t_2/transmission_gate_0/en sky130_fd_sc_hd__inv_1_3/Y 0.16fF
C26 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/en_b 1.46fF
C27 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/in 0.09fF
C28 en switch_5t_0/transmission_gate_0/in 0.68fF
C29 sky130_fd_sc_hd__nand2_1_0/Y a_n499_n3694# 0.02fF
C30 switch_5t_1/transmission_gate_0/en_b transmission_gate_0/en_b 0.06fF
C31 s1 switch_5t_3/transmission_gate_0/in 0.02fF
C32 s0 sky130_fd_sc_hd__nand2_1_3/B 0.34fF
C33 switch_5t_2/transmission_gate_0/en transmission_gate_0/en_b 0.04fF
C34 switch_5t_2/transmission_gate_0/in out 0.43fF
C35 s1 switch_5t_1/transmission_gate_0/in 0.06fF
C36 VDD s1 1.02fF
C37 switch_5t_1/transmission_gate_0/out switch_5t_1/transmission_gate_0/en 2.01fF
C38 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/en 1.53fF
C39 a_n499_n2606# s1 0.00fF
C40 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/B 0.02fF
C41 switch_5t_2/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/in 0.02fF
C42 en transmission_gate_0/en_b 3.34fF
C43 VDD switch_5t_1/transmission_gate_0/en 0.44fF
C44 switch_5t_2/transmission_gate_0/out s1 0.01fF
C45 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C46 switch_5t_0/transmission_gate_0/out switch_5t_1/transmission_gate_0/en 0.03fF
C47 s0 in1 0.00fF
C48 switch_5t_1/transmission_gate_0/en_b s1 0.07fF
C49 out switch_5t_0/transmission_gate_0/in 0.43fF
C50 in2 sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C51 switch_5t_2/transmission_gate_0/en s1 0.03fF
C52 in2 in3 0.23fF
C53 out sky130_fd_sc_hd__inv_1_3/Y 0.64fF
C54 switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/en 0.54fF
C55 sky130_fd_sc_hd__nand2_1_0/Y transmission_gate_0/en_b 0.04fF
C56 switch_5t_2/transmission_gate_0/en_b transmission_gate_0/en_b 0.04fF
C57 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/B 0.07fF
C58 switch_5t_2/transmission_gate_0/in in1 0.06fF
C59 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nand2_1_3/B 0.00fF
C60 en s1 0.66fF
C61 VDD switch_5t_3/transmission_gate_0/in 2.44fF
C62 switch_5t_3/transmission_gate_0/en switch_5t_3/transmission_gate_0/in 1.57fF
C63 switch_5t_1/transmission_gate_0/in switch_5t_1/transmission_gate_0/out 7.39fF
C64 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__nand2_1_3/A 0.19fF
C65 en switch_5t_1/transmission_gate_0/en 0.07fF
C66 VDD switch_5t_1/transmission_gate_0/out 2.93fF
C67 VDD switch_5t_1/transmission_gate_0/in 3.13fF
C68 switch_5t_2/transmission_gate_0/out switch_5t_3/transmission_gate_0/in 0.06fF
C69 transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B 0.04fF
C70 VDD switch_5t_3/transmission_gate_0/en 0.58fF
C71 s0 in2 0.00fF
C72 switch_5t_0/transmission_gate_0/out switch_5t_1/transmission_gate_0/out 0.33fF
C73 in1 switch_5t_0/transmission_gate_0/in 6.76fF
C74 switch_5t_0/transmission_gate_0/out switch_5t_1/transmission_gate_0/in 0.07fF
C75 VDD switch_5t_0/transmission_gate_0/out 3.04fF
C76 sky130_fd_sc_hd__nand2_1_0/Y s1 0.08fF
C77 switch_5t_2/transmission_gate_0/en_b s1 0.07fF
C78 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/in 7.32fF
C79 switch_5t_2/transmission_gate_0/out VDD 3.01fF
C80 switch_5t_2/transmission_gate_0/en switch_5t_3/transmission_gate_0/in 0.04fF
C81 switch_5t_2/transmission_gate_0/out switch_5t_3/transmission_gate_0/en 0.09fF
C82 switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/out 1.88fF
C83 switch_5t_1/transmission_gate_0/en_b switch_5t_1/transmission_gate_0/in 1.39fF
C84 switch_5t_1/transmission_gate_0/en_b VDD 3.71fF
C85 switch_5t_2/transmission_gate_0/in in2 6.62fF
C86 switch_5t_0/transmission_gate_0/in in0 0.06fF
C87 switch_5t_2/transmission_gate_0/out switch_5t_0/transmission_gate_0/out 0.30fF
C88 VDD switch_5t_3/transmission_gate_0/out 2.72fF
C89 switch_5t_2/transmission_gate_0/en VDD 0.57fF
C90 switch_5t_3/transmission_gate_0/out switch_5t_3/transmission_gate_0/en 1.97fF
C91 switch_5t_2/transmission_gate_0/en switch_5t_3/transmission_gate_0/en 0.25fF
C92 s0 sky130_fd_sc_hd__inv_1_3/A 0.10fF
C93 en switch_5t_3/transmission_gate_0/in 0.63fF
C94 switch_5t_1/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/out 0.12fF
C95 in1 transmission_gate_0/en_b 1.29fF
C96 out switch_5t_1/transmission_gate_0/en 0.58fF
C97 a_n499_n2830# switch_5t_2/transmission_gate_0/en_b 0.01fF
C98 switch_5t_2/transmission_gate_0/out switch_5t_3/transmission_gate_0/out 0.30fF
C99 switch_5t_2/transmission_gate_0/en switch_5t_0/transmission_gate_0/out 0.09fF
C100 en switch_5t_1/transmission_gate_0/out 0.00fF
C101 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/out 1.96fF
C102 s1 sky130_fd_sc_hd__nand2_1_3/B 0.36fF
C103 en switch_5t_1/transmission_gate_0/in 0.70fF
C104 en VDD 0.48fF
C105 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/A 0.06fF
C106 in0 transmission_gate_0/en_b 1.33fF
C107 switch_5t_2/transmission_gate_0/en switch_5t_3/transmission_gate_0/out 0.02fF
C108 in2 switch_5t_0/transmission_gate_0/in 0.07fF
C109 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/in 1.40fF
C110 switch_5t_2/transmission_gate_0/en_b switch_5t_3/transmission_gate_0/in 0.09fF
C111 switch_5t_1/transmission_gate_0/en_b a_n499_n1742# 0.01fF
C112 s0 sky130_fd_sc_hd__nand2_1_3/A 1.04fF
C113 en switch_5t_1/transmission_gate_0/en_b 0.07fF
C114 switch_5t_2/transmission_gate_0/en en 0.03fF
C115 sky130_fd_sc_hd__nand2_1_0/Y VDD 3.70fF
C116 switch_5t_2/transmission_gate_0/en_b VDD 3.75fF
C117 out switch_5t_3/transmission_gate_0/in 0.43fF
C118 switch_5t_2/transmission_gate_0/en_b switch_5t_3/transmission_gate_0/en 0.46fF
C119 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/en 0.55fF
C120 sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/in 1.59fF
C121 in2 transmission_gate_0/en_b 1.30fF
C122 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/A 0.08fF
C123 out switch_5t_1/transmission_gate_0/out 7.54fF
C124 switch_5t_2/transmission_gate_0/in in3 0.07fF
C125 switch_5t_2/transmission_gate_0/en_b switch_5t_0/transmission_gate_0/out 0.02fF
C126 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_3/Y 0.62fF
C127 out switch_5t_1/transmission_gate_0/in 0.43fF
C128 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/out 0.06fF
C129 switch_5t_2/transmission_gate_0/out switch_5t_2/transmission_gate_0/en_b 1.89fF
C130 out VDD 6.03fF
C131 out switch_5t_3/transmission_gate_0/en 0.63fF
C132 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_1/transmission_gate_0/en_b 0.00fF
C133 switch_5t_1/transmission_gate_0/en_b switch_5t_2/transmission_gate_0/en_b 0.01fF
C134 switch_5t_1/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/B 0.02fF
C135 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_3/transmission_gate_0/out 1.85fF
C136 switch_5t_2/transmission_gate_0/en_b switch_5t_3/transmission_gate_0/out 0.09fF
C137 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/en 0.19fF
C138 switch_5t_2/transmission_gate_0/en switch_5t_2/transmission_gate_0/en_b 1.01fF
C139 out switch_5t_0/transmission_gate_0/out 7.67fF
C140 VDD sky130_fd_sc_hd__nand2_1_3/B 1.22fF
C141 out switch_5t_2/transmission_gate_0/out 7.67fF
C142 sky130_fd_sc_hd__inv_1_3/A transmission_gate_0/en_b 0.04fF
C143 out switch_5t_1/transmission_gate_0/en_b 0.50fF
C144 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/A 0.08fF
C145 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_3/B 0.02fF
C146 out switch_5t_3/transmission_gate_0/out 7.47fF
C147 switch_5t_2/transmission_gate_0/en out 0.64fF
C148 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C149 en switch_5t_2/transmission_gate_0/en_b 0.03fF
C150 sky130_fd_sc_hd__nand2_1_0/Y en 0.06fF
C151 in2 s1 0.00fF
C152 switch_5t_2/transmission_gate_0/in s0 0.46fF
C153 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B 0.06fF
C154 in1 switch_5t_1/transmission_gate_0/in 0.07fF
C155 VDD in1 1.23fF
C156 transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A 0.10fF
C157 in3 transmission_gate_0/en_b 1.23fF
C158 sky130_fd_sc_hd__inv_1_3/A s1 0.39fF
C159 sky130_fd_sc_hd__nand2_1_0/Y switch_5t_2/transmission_gate_0/en_b 0.39fF
C160 en sky130_fd_sc_hd__nand2_1_3/B 0.03fF
C161 switch_5t_1/transmission_gate_0/in in0 6.63fF
C162 VDD in0 1.35fF
C163 s0 switch_5t_0/transmission_gate_0/in 0.07fF
C164 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/en 0.02fF
C165 s0 sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C166 out switch_5t_2/transmission_gate_0/en_b 0.51fF
C167 sky130_fd_sc_hd__nand2_1_0/Y out 0.45fF
C168 in2 switch_5t_3/transmission_gate_0/in 0.06fF
C169 switch_5t_2/transmission_gate_0/in switch_5t_0/transmission_gate_0/in 0.30fF
C170 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/B 0.00fF
C171 switch_5t_2/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C172 s1 sky130_fd_sc_hd__nand2_1_3/A 0.51fF
C173 s0 transmission_gate_0/en_b 0.47fF
C174 in2 VDD 1.28fF
C175 en in1 1.35fF
C176 switch_5t_1/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C177 en in0 1.35fF
C178 switch_5t_2/transmission_gate_0/in transmission_gate_0/en_b 0.58fF
C179 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/out 0.03fF
C180 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/in 0.05fF
C181 switch_5t_0/transmission_gate_0/in sky130_fd_sc_hd__inv_1_3/Y 1.57fF
C182 sky130_fd_sc_hd__inv_1_3/A VDD 3.71fF
C183 sky130_fd_sc_hd__inv_1_3/A a_n499_n2606# 0.02fF
C184 s0 s1 2.22fF
C185 sky130_fd_sc_hd__inv_1_3/A switch_5t_0/transmission_gate_0/out 1.89fF
C186 sky130_fd_sc_hd__inv_1_3/A switch_5t_2/transmission_gate_0/out 0.09fF
C187 in2 en 1.37fF
C188 s0 switch_5t_1/transmission_gate_0/en 0.03fF
C189 switch_5t_0/transmission_gate_0/in transmission_gate_0/en_b 0.82fF
C190 in3 switch_5t_3/transmission_gate_0/in 6.62fF
C191 sky130_fd_sc_hd__inv_1_3/A switch_5t_1/transmission_gate_0/en_b 0.47fF
C192 sky130_fd_sc_hd__inv_1_3/Y transmission_gate_0/en_b 0.01fF
C193 switch_5t_2/transmission_gate_0/en sky130_fd_sc_hd__inv_1_3/A 0.42fF
C194 switch_5t_2/transmission_gate_0/in s1 0.30fF
C195 switch_5t_1/transmission_gate_0/in sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C196 in1 sky130_fd_sc_hd__nand2_1_3/B 0.01fF
C197 VDD sky130_fd_sc_hd__nand2_1_3/A 1.38fF
C198 VDD in3 1.13fF
C199 a_n499_n2830# s0 0.00fF
C200 switch_5t_0/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C201 switch_5t_2/transmission_gate_0/out sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C202 sky130_fd_sc_hd__inv_1_3/A en 0.03fF
C203 switch_5t_1/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A 0.21fF
C204 s1 switch_5t_0/transmission_gate_0/in 0.08fF
C205 switch_5t_2/transmission_gate_0/en sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C206 s0 switch_5t_3/transmission_gate_0/in 0.01fF
C207 s1 sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C208 switch_5t_0/transmission_gate_0/in switch_5t_1/transmission_gate_0/en 0.01fF
C209 s0 switch_5t_1/transmission_gate_0/in 0.04fF
C210 s0 VDD 1.24fF
C211 sky130_fd_sc_hd__inv_1_3/Y switch_5t_1/transmission_gate_0/en 0.20fF
C212 sky130_fd_sc_hd__inv_1_3/A switch_5t_2/transmission_gate_0/en_b 0.23fF
C213 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_3/A 0.01fF
C214 s0 switch_5t_3/transmission_gate_0/en 0.01fF
C215 en sky130_fd_sc_hd__nand2_1_3/A 0.07fF
C216 switch_5t_2/transmission_gate_0/in switch_5t_3/transmission_gate_0/in 0.35fF
C217 in1 in0 0.25fF
C218 en in3 1.34fF
C219 s0 switch_5t_2/transmission_gate_0/out 0.02fF
C220 s1 transmission_gate_0/en_b 1.15fF
C221 sky130_fd_sc_hd__inv_1_3/A out 0.51fF
C222 switch_5t_2/transmission_gate_0/in VDD 3.32fF
C223 switch_5t_2/transmission_gate_0/in switch_5t_3/transmission_gate_0/en 0.07fF
C224 s0 switch_5t_1/transmission_gate_0/en_b 0.08fF
C225 switch_5t_1/transmission_gate_0/en transmission_gate_0/en_b 0.07fF
C226 switch_5t_2/transmission_gate_0/en s0 0.09fF
C227 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__nand2_1_3/B 0.20fF
C228 switch_5t_2/transmission_gate_0/in switch_5t_0/transmission_gate_0/out 0.06fF
C229 switch_5t_2/transmission_gate_0/in switch_5t_2/transmission_gate_0/out 7.32fF
C230 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C231 switch_5t_2/transmission_gate_0/en_b sky130_fd_sc_hd__nand2_1_3/A 0.09fF
C232 in2 in1 0.23fF
C233 switch_5t_2/transmission_gate_0/in switch_5t_1/transmission_gate_0/en_b 0.00fF
C234 switch_5t_0/transmission_gate_0/in switch_5t_1/transmission_gate_0/out 0.06fF
C235 switch_5t_3/transmission_gate_0/out VSS 2.21fF
C236 switch_5t_3/transmission_gate_0/en VSS 3.37fF
C237 in3 VSS 1.22fF
C238 switch_5t_3/transmission_gate_0/in VSS 2.54fF
C239 a_n499_n3694# VSS 0.00fF
C240 sky130_fd_sc_hd__nand2_1_0/Y VSS 1.45fF
C241 switch_5t_2/transmission_gate_0/out VSS 2.35fF
C242 switch_5t_2/transmission_gate_0/en VSS 3.94fF
C243 in2 VSS 1.28fF
C244 switch_5t_2/transmission_gate_0/in VSS 2.87fF
C245 switch_5t_2/transmission_gate_0/en_b VSS 1.41fF
C246 a_n499_n2830# VSS 0.01fF
C247 a_n499_n2606# VSS 0.00fF
C248 s1 VSS 2.28fF
C249 s0 VSS 1.60fF
C250 switch_5t_0/transmission_gate_0/out VSS 2.34fF
C251 a_n499_n1742# VSS 0.01fF
C252 sky130_fd_sc_hd__nand2_1_3/A VSS 0.97fF
C253 sky130_fd_sc_hd__nand2_1_3/B VSS 0.70fF
C254 in1 VSS 1.30fF
C255 switch_5t_0/transmission_gate_0/in VSS 3.43fF
C256 sky130_fd_sc_hd__inv_1_3/Y VSS 3.75fF
C257 sky130_fd_sc_hd__inv_1_3/A VSS 1.52fF
C258 en VSS 9.89fF
C259 out VSS 5.26fF
C260 switch_5t_1/transmission_gate_0/en_b VSS 1.23fF
C261 switch_5t_1/transmission_gate_0/out VSS 2.45fF
C262 switch_5t_1/transmission_gate_0/en VSS 4.40fF
C263 in0 VSS 1.28fF
C264 switch_5t_1/transmission_gate_0/in VSS 3.06fF
C265 transmission_gate_0/en_b VSS 3.07fF
C266 VDD VSS 47.88fF
.ends

