magic
tech sky130A
magscale 1 2
timestamp 1654675174
<< metal1 >>
rect 103391 71867 104426 71889
rect 36352 71835 37396 71862
rect 36352 70835 36373 71835
rect 37373 70835 37396 71835
rect 36352 70810 37396 70835
rect 43351 71817 44375 71828
rect 43351 70817 43364 71817
rect 44364 70817 44375 71817
rect 36795 70435 36923 70810
rect 43351 70806 44375 70817
rect 57794 71821 58825 71840
rect 57794 70821 57809 71821
rect 58809 70821 58825 71821
rect 74871 71807 75895 71820
rect 43795 70435 43923 70806
rect 57794 70802 58825 70821
rect 64867 71771 65896 71786
rect 58215 70435 58343 70802
rect 64867 70771 64881 71771
rect 65881 70771 65896 71771
rect 74871 70807 74883 71807
rect 75883 70807 75895 71807
rect 94051 71783 95086 71805
rect 74871 70796 75895 70807
rect 85821 71759 86856 71781
rect 64867 70758 65896 70771
rect 65315 70435 65443 70758
rect 75315 70435 75443 70796
rect 85821 70759 85838 71759
rect 86838 70759 86856 71759
rect 94051 70783 94068 71783
rect 95068 70783 95086 71783
rect 103391 70867 103408 71867
rect 104408 70867 104426 71867
rect 103391 70852 104426 70867
rect 94051 70768 95086 70783
rect 85821 70744 86856 70759
rect 86265 70435 86393 70744
rect 94495 70563 94623 70768
rect 103835 70435 103963 70852
rect 36795 66876 36923 67015
rect 36795 66742 36923 66748
rect 43795 66816 43923 67196
rect 43795 66682 43923 66688
rect 38709 57231 38837 57237
rect 43795 57231 43923 57237
rect 82647 57231 82775 57237
rect 38837 57103 43795 57231
rect 43923 57103 82647 57231
rect 38709 57097 38837 57103
rect 43795 57097 43923 57103
rect 82647 57097 82775 57103
rect 36795 55845 36923 55851
rect 80625 55845 80753 55851
rect 36923 55717 80625 55845
rect 36795 55711 36923 55717
rect 80625 55711 80753 55717
rect 48941 54451 49059 54457
rect 48934 54333 48941 54451
rect 49059 54450 120608 54451
rect 49059 54333 87250 54450
rect 48941 54327 49059 54333
rect 87244 54332 87250 54333
rect 87368 54333 120608 54450
rect 87368 54332 87374 54333
rect 85345 53410 85463 53416
rect 46935 53292 85345 53410
rect 85463 53292 116623 53410
rect 46935 52387 47053 53292
rect 85345 53286 85463 53292
rect 48935 52399 48941 52517
rect 49059 52399 49065 52517
rect 116505 52230 116623 53292
rect 120490 52241 120608 54333
rect 48730 51289 48873 51297
rect 46745 51153 46751 51281
rect 46879 51153 46885 51281
rect 48730 51161 48737 51289
rect 48865 51161 48873 51289
rect 48730 51154 48873 51161
rect 36789 50498 36795 50626
rect 36923 50498 36929 50626
rect 38703 50500 38709 50628
rect 38837 50500 38843 50628
rect 36795 50381 36923 50498
rect 38709 50376 38837 50500
rect 116873 50236 116991 50242
rect 120884 50236 121002 50242
rect 126619 50236 126751 50243
rect 116991 50118 120884 50236
rect 121002 50118 126626 50236
rect 126744 50118 126751 50236
rect 116873 50112 116991 50118
rect 120884 50112 121002 50118
rect 126619 50111 126751 50118
rect 116334 49381 116452 49387
rect 120328 49381 120460 49387
rect 125957 49381 126075 49387
rect 36683 49210 36693 49338
rect 36821 49210 36831 49338
rect 38682 49225 38692 49353
rect 38820 49225 38830 49353
rect 116452 49263 120335 49381
rect 120453 49263 125957 49381
rect 116334 49257 116452 49263
rect 120328 49256 120460 49263
rect 125957 49257 126075 49263
rect 36693 48424 36821 48430
rect 46751 48424 46879 48430
rect 36821 48296 46751 48424
rect 36693 48290 36821 48296
rect 46751 48290 46879 48296
rect 48737 47288 48865 47294
rect 38674 47160 38680 47288
rect 38808 47160 48737 47288
rect 48737 47154 48865 47160
rect 38686 45429 38692 45557
rect 38820 45429 44965 45557
rect 45093 45429 45099 45557
rect 85345 43190 85463 43196
rect 85345 43066 85463 43072
rect 87250 43186 87368 43192
rect 87250 43062 87368 43068
rect 85234 41840 85240 41968
rect 85368 41840 85374 41968
rect 87241 41829 87247 41957
rect 87375 41829 87381 41957
rect 80619 41245 80625 41373
rect 80753 41245 80759 41373
rect 82641 41261 82647 41389
rect 82775 41261 82781 41389
rect 80633 40168 80780 40176
rect 80633 40040 80643 40168
rect 80771 40040 80780 40168
rect 80633 40033 80780 40040
rect 82645 40162 82773 40168
rect 82645 40028 82773 40034
rect 86311 39407 86317 39417
rect 82639 39279 82645 39407
rect 82773 39289 86317 39407
rect 86445 39407 86451 39417
rect 87247 39407 87375 39413
rect 86445 39289 87247 39407
rect 82773 39279 87247 39289
rect 87247 39273 87375 39279
rect 40699 39232 40931 39246
rect 51833 39232 52039 39238
rect 40699 39026 40712 39232
rect 40918 39026 51833 39232
rect 40699 39012 40931 39026
rect 51833 39020 52039 39026
rect 82310 38567 82438 38573
rect 85240 38567 85368 38573
rect 80637 38439 80643 38567
rect 80771 38439 82310 38567
rect 82438 38439 85240 38567
rect 82310 38433 82438 38439
rect 85240 38433 85368 38439
rect 85321 37663 85449 37669
rect 85449 37535 86317 37663
rect 86445 37535 86451 37663
rect 85321 37529 85449 37535
rect 89487 36058 89693 36064
rect 86373 36022 86501 36028
rect 86501 35894 89487 36022
rect 86373 35888 86501 35894
rect 89487 35846 89693 35852
rect 50201 35813 50433 35828
rect 50201 35607 50215 35813
rect 50421 35607 54340 35813
rect 54546 35607 54552 35813
rect 50201 35594 50433 35607
rect 86360 35183 86514 35338
rect 83771 34890 83928 34908
rect 88533 34890 88556 34918
rect 83771 34762 83785 34890
rect 83913 34762 88556 34890
rect 83771 34736 83928 34762
rect 88533 34712 88556 34762
rect 88762 34712 88768 34918
rect 107424 34896 108254 35014
rect 108372 34896 108378 35014
rect 110860 34896 110866 35014
rect 110984 34896 110990 35014
rect 67544 33674 67550 33792
rect 67668 33674 67674 33792
rect 60673 33204 63007 33322
rect 60702 33185 60712 33204
rect 60676 31414 61695 31532
rect 60699 31382 60712 31414
rect 61569 28056 61687 31414
rect 61568 27997 61687 28056
rect 38285 27752 38403 27758
rect 42065 27752 42183 27758
rect 38403 27634 42065 27752
rect 42183 27634 44800 27752
rect 44918 27634 44924 27752
rect 38285 27628 38403 27634
rect 42065 27628 42183 27634
rect 61568 26993 61686 27997
rect 55807 26875 55813 26993
rect 55931 26875 61686 26993
rect 45223 26341 45341 26347
rect 45341 26223 46166 26341
rect 46284 26223 46290 26341
rect 45223 26217 45341 26223
rect 56821 26199 56939 26205
rect 62889 26200 63007 33204
rect 67550 27921 67668 33674
rect 67544 27803 67550 27921
rect 67668 27803 67674 27921
rect 69183 27908 69301 34332
rect 83813 33792 83961 33810
rect 83813 33674 83827 33792
rect 83945 33674 88643 33792
rect 88761 33674 88767 33792
rect 83813 33655 83961 33674
rect 107303 33517 107421 34312
rect 107297 33399 107303 33517
rect 107421 33399 107427 33517
rect 95208 33207 97247 33325
rect 95223 33112 95228 33207
rect 77070 31877 77188 31883
rect 81834 31877 81976 31890
rect 77188 31759 81847 31877
rect 81965 31759 81976 31877
rect 77070 31753 77188 31759
rect 81834 31746 81976 31759
rect 86778 31819 86965 31853
rect 86778 31701 86818 31819
rect 86936 31701 87767 31819
rect 87885 31701 87891 31819
rect 86778 31671 86965 31701
rect 95177 31414 96047 31532
rect 95219 31382 95228 31414
rect 78343 29370 78461 29376
rect 84866 29370 84984 29376
rect 78340 29252 78343 29370
rect 78461 29252 84866 29370
rect 78343 29246 78461 29252
rect 84866 29246 84984 29252
rect 82222 28351 82355 28361
rect 80004 28233 80010 28351
rect 80128 28233 82231 28351
rect 82349 28233 82355 28351
rect 82222 28226 82355 28233
rect 92040 28019 92246 28025
rect 93382 28019 93588 28025
rect 69177 27790 69183 27908
rect 69301 27790 69307 27908
rect 92246 27813 93382 28019
rect 92040 27807 92246 27813
rect 93382 27807 93588 27813
rect 80943 27024 80949 27142
rect 81067 27024 85794 27142
rect 85912 27024 85918 27142
rect 88643 26607 88761 26613
rect 95929 26607 96047 31414
rect 88761 26489 96047 26607
rect 88643 26483 88761 26489
rect 61176 26199 63007 26200
rect 56939 26082 63007 26199
rect 56939 26081 61191 26082
rect 56821 26075 56939 26081
rect 58184 25335 58302 25341
rect 67550 25335 67668 25341
rect 58302 25217 67550 25335
rect 58184 25211 58302 25217
rect 67550 25211 67668 25217
rect 97129 25170 97247 33207
rect 107303 32812 107421 33399
rect 110866 32825 110984 34896
rect 125957 34488 126075 34494
rect 125632 34370 125957 34382
rect 127075 34382 127203 34425
rect 126075 34370 127203 34382
rect 125632 34348 127203 34370
rect 127075 34297 127203 34348
rect 126626 33700 126744 33706
rect 125624 33582 126626 33597
rect 126744 33582 127505 33597
rect 125624 33563 127505 33582
rect 126900 33268 126934 33563
rect 126900 33234 127488 33268
rect 126900 32957 126934 33234
rect 126900 32923 127487 32957
rect 110860 32707 110866 32825
rect 110984 32707 110990 32825
rect 126900 32717 126934 32923
rect 107303 32688 107421 32694
rect 126900 32683 127487 32717
rect 110889 28334 111007 28340
rect 107294 28315 107428 28322
rect 107294 28197 107303 28315
rect 107421 28197 108683 28315
rect 109786 28216 110889 28334
rect 110889 28210 111007 28216
rect 107294 28184 107428 28197
rect 93204 25052 93210 25170
rect 93328 25052 97247 25170
rect 39593 24596 39711 24602
rect 39711 24478 45918 24596
rect 46036 24478 46042 24596
rect 39593 24472 39711 24478
rect 88643 24435 88761 24441
rect 82029 24422 82147 24428
rect 69183 24414 69301 24420
rect 59549 24296 59555 24414
rect 59673 24296 69183 24414
rect 82147 24304 85449 24422
rect 86555 24317 88643 24435
rect 88643 24311 88761 24317
rect 82029 24298 82147 24304
rect 69183 24290 69301 24296
rect 88643 23243 88761 23249
rect 36559 23142 36699 23148
rect 36559 23014 36565 23142
rect 36693 23014 43321 23142
rect 44435 23112 49046 23116
rect 36559 23008 36699 23014
rect 44435 22998 45918 23112
rect 45912 22994 45918 22998
rect 46036 22998 49046 23112
rect 49164 22998 53351 23116
rect 55813 23110 55931 23116
rect 46036 22994 46042 22998
rect 54451 22992 55813 23110
rect 59549 23015 59555 23133
rect 59673 23015 62367 23133
rect 83734 23123 84288 23241
rect 84406 23123 84412 23241
rect 88761 23125 89438 23243
rect 90859 23241 90977 23247
rect 63471 23105 67640 23110
rect 63471 22992 65692 23105
rect 55813 22986 55931 22992
rect 65686 22987 65692 22992
rect 65810 22992 67640 23105
rect 67758 22992 71434 23110
rect 77064 23108 77070 23123
rect 65810 22987 65816 22992
rect 72533 22990 74332 23108
rect 74450 23005 77070 23108
rect 77188 23108 77194 23123
rect 80010 23117 80128 23123
rect 88643 23119 88761 23125
rect 90536 23123 90859 23241
rect 90859 23117 90977 23123
rect 77188 23005 80010 23108
rect 74450 22999 80010 23005
rect 82029 23108 82147 23114
rect 80128 22999 82029 23108
rect 74450 22990 82029 22999
rect 82147 22990 82621 23108
rect 82029 22984 82147 22990
rect 36554 21115 36700 21124
rect 36554 20987 36565 21115
rect 36693 20987 39756 21115
rect 41572 21108 41690 21114
rect 47715 21109 47833 21115
rect 40858 20990 41572 21108
rect 45912 20990 45918 21108
rect 46036 20990 46337 21108
rect 47449 20991 47715 21109
rect 49564 21009 49570 21127
rect 49688 21009 50149 21127
rect 55813 21113 55931 21119
rect 51245 20995 55813 21113
rect 59549 20996 59555 21114
rect 59673 20996 60152 21114
rect 64422 21111 64540 21117
rect 36554 20977 36700 20987
rect 41572 20984 41690 20990
rect 47715 20985 47833 20991
rect 55813 20989 55931 20995
rect 61241 20993 64422 21111
rect 64422 20987 64540 20993
rect 67630 20753 67640 20871
rect 67758 20753 67768 20871
rect 74322 20507 74332 20625
rect 74450 20507 74460 20625
rect 92040 20242 92246 20248
rect 84278 20208 84416 20218
rect 90811 20208 92040 20242
rect 47715 20171 47833 20172
rect 48344 20171 48462 20177
rect 47648 20166 48344 20171
rect 41566 20048 41572 20166
rect 41690 20048 47715 20166
rect 47833 20053 48344 20166
rect 84278 20090 84288 20208
rect 84406 20090 90859 20208
rect 90977 20090 92040 20208
rect 84278 20084 84416 20090
rect 47833 20048 47842 20053
rect 47715 20042 47833 20048
rect 48344 20047 48462 20053
rect 90811 20036 92040 20090
rect 92040 20030 92246 20036
rect 67627 19527 67637 19645
rect 67755 19527 67765 19645
rect 74330 19411 74448 19417
rect 74330 19287 74448 19293
rect 49046 19143 49164 19149
rect 38285 19128 38403 19134
rect 38403 19010 39763 19128
rect 41572 19118 41690 19124
rect 38285 19004 38403 19010
rect 40869 19000 41572 19118
rect 41572 18994 41690 19000
rect 45223 19116 45341 19122
rect 45341 18998 45909 19116
rect 46027 18998 46338 19116
rect 47715 19109 47833 19115
rect 45223 18992 45341 18998
rect 47439 18991 47715 19109
rect 49164 19025 50128 19143
rect 55826 19112 55944 19118
rect 49046 19019 49164 19025
rect 51249 18994 55826 19112
rect 58178 18995 58184 19113
rect 58302 18995 60137 19113
rect 61249 18994 65692 19112
rect 65810 18994 65816 19112
rect 47715 18985 47833 18991
rect 55826 18988 55944 18994
rect 93210 18837 93328 18843
rect 87761 18719 87767 18837
rect 87885 18719 88626 18837
rect 88744 18719 93210 18837
rect 93210 18713 93328 18719
rect 56821 18089 56939 18095
rect 55820 17971 55826 18089
rect 55944 17971 56821 18089
rect 56821 17965 56939 17971
rect 58184 17157 58302 17163
rect 83725 17161 84288 17279
rect 84406 17161 84412 17279
rect 90859 17274 90977 17280
rect 45903 17115 45909 17127
rect 38285 17093 38403 17099
rect 38403 16975 43332 17093
rect 44439 17009 45909 17115
rect 46027 17115 46033 17127
rect 46027 17009 49570 17115
rect 44439 16997 49570 17009
rect 49688 16997 53335 17115
rect 55826 17109 55944 17115
rect 54444 16991 55826 17109
rect 58302 17039 62353 17157
rect 88620 17155 88626 17273
rect 88744 17155 89431 17273
rect 90533 17156 90859 17274
rect 90859 17150 90977 17156
rect 80943 17123 80949 17124
rect 67628 17112 67638 17113
rect 58184 17033 58302 17039
rect 63464 16994 64422 17112
rect 64540 16995 67638 17112
rect 67756 17112 67766 17113
rect 67756 16995 71417 17112
rect 72540 17005 74330 17123
rect 74448 17121 80949 17123
rect 74448 17005 78343 17121
rect 78337 17003 78343 17005
rect 78461 17006 80949 17121
rect 81067 17123 81073 17124
rect 82020 17123 82160 17137
rect 81067 17006 82030 17123
rect 78461 17005 82030 17006
rect 82148 17005 82613 17123
rect 78461 17003 78467 17005
rect 64540 16994 71417 16995
rect 82020 16993 82160 17005
rect 55826 16985 55944 16991
rect 38285 16969 38403 16975
rect 88626 16423 88744 16429
rect 82030 16379 82148 16385
rect 82148 16261 85434 16379
rect 86554 16305 88626 16423
rect 88626 16299 88744 16305
rect 82030 16255 82148 16261
rect 71861 -2025 71989 -2015
rect 71861 -2163 71989 -2153
rect 72403 -2026 72531 -2016
rect 72403 -2164 72531 -2154
rect 72947 -2025 73075 -2015
rect 72947 -2163 73075 -2153
rect 73486 -2026 73614 -2016
rect 73486 -2164 73614 -2154
rect 75127 -2025 75255 -2015
rect 75127 -2163 75255 -2153
rect 75663 -2026 75791 -2016
rect 75663 -2164 75791 -2154
rect 76213 -2025 76341 -2015
rect 76213 -2163 76341 -2153
rect 76749 -2026 76877 -2016
rect 76749 -2164 76877 -2154
rect 79480 -2026 79608 -2016
rect 79480 -2164 79608 -2154
rect 80017 -2025 80145 -2015
rect 80017 -2163 80145 -2153
rect 80562 -2027 80690 -2017
rect 80562 -2165 80690 -2155
rect 81110 -2026 81238 -2016
rect 81110 -2164 81238 -2154
rect 82738 -2026 82866 -2016
rect 82738 -2164 82866 -2154
rect 83284 -2026 83412 -2016
rect 83284 -2164 83412 -2154
rect 83835 -2025 83963 -2015
rect 83835 -2163 83963 -2153
rect 84366 -2026 84494 -2016
rect 84366 -2164 84494 -2154
<< via1 >>
rect 36373 70835 37373 71835
rect 43364 70817 44364 71817
rect 57809 70821 58809 71821
rect 64881 70771 65881 71771
rect 74883 70807 75883 71807
rect 85838 70759 86838 71759
rect 94068 70783 95068 71783
rect 103408 70867 104408 71867
rect 36795 66748 36923 66876
rect 43795 66688 43923 66816
rect 38709 57103 38837 57231
rect 43795 57103 43923 57231
rect 82647 57103 82775 57231
rect 36795 55717 36923 55845
rect 80625 55717 80753 55845
rect 48941 54333 49059 54451
rect 87250 54332 87368 54450
rect 85345 53292 85463 53410
rect 48941 52399 49059 52517
rect 46751 51153 46879 51281
rect 48737 51161 48865 51289
rect 36795 50498 36923 50626
rect 38709 50500 38837 50628
rect 116873 50118 116991 50236
rect 120884 50118 121002 50236
rect 126626 50118 126744 50236
rect 36693 49210 36821 49338
rect 38692 49225 38820 49353
rect 116334 49263 116452 49381
rect 120335 49263 120453 49381
rect 125957 49263 126075 49381
rect 36693 48296 36821 48424
rect 46751 48296 46879 48424
rect 38680 47160 38808 47288
rect 48737 47160 48865 47288
rect 38692 45429 38820 45557
rect 44965 45429 45093 45557
rect 85345 43072 85463 43190
rect 87250 43068 87368 43186
rect 85240 41840 85368 41968
rect 87247 41829 87375 41957
rect 80625 41245 80753 41373
rect 82647 41261 82775 41389
rect 80643 40040 80771 40168
rect 82645 40034 82773 40162
rect 82645 39279 82773 39407
rect 86317 39289 86445 39417
rect 87247 39279 87375 39407
rect 40712 39026 40918 39232
rect 51833 39026 52039 39232
rect 80643 38439 80771 38567
rect 82310 38439 82438 38567
rect 85240 38439 85368 38567
rect 85321 37535 85449 37663
rect 86317 37535 86445 37663
rect 86373 35894 86501 36022
rect 89487 35852 89693 36058
rect 50215 35607 50421 35813
rect 54340 35607 54546 35813
rect 83785 34762 83913 34890
rect 88556 34712 88762 34918
rect 108254 34896 108372 35014
rect 110866 34896 110984 35014
rect 67550 33674 67668 33792
rect 38285 27634 38403 27752
rect 42065 27634 42183 27752
rect 44800 27634 44918 27752
rect 55813 26875 55931 26993
rect 45223 26223 45341 26341
rect 46166 26223 46284 26341
rect 67550 27803 67668 27921
rect 83827 33674 83945 33792
rect 88643 33674 88761 33792
rect 107303 33399 107421 33517
rect 77070 31759 77188 31877
rect 81847 31759 81965 31877
rect 86818 31701 86936 31819
rect 87767 31701 87885 31819
rect 78343 29252 78461 29370
rect 84866 29252 84984 29370
rect 80010 28233 80128 28351
rect 82231 28233 82349 28351
rect 69183 27790 69301 27908
rect 92040 27813 92246 28019
rect 93382 27813 93588 28019
rect 80949 27024 81067 27142
rect 85794 27024 85912 27142
rect 88643 26489 88761 26607
rect 56821 26081 56939 26199
rect 58184 25217 58302 25335
rect 67550 25217 67668 25335
rect 125957 34370 126075 34488
rect 126626 33582 126744 33700
rect 107303 32694 107421 32812
rect 110866 32707 110984 32825
rect 107303 28197 107421 28315
rect 110889 28216 111007 28334
rect 93210 25052 93328 25170
rect 39593 24478 39711 24596
rect 45918 24478 46036 24596
rect 59555 24296 59673 24414
rect 69183 24296 69301 24414
rect 82029 24304 82147 24422
rect 88643 24317 88761 24435
rect 36565 23014 36693 23142
rect 45918 22994 46036 23112
rect 49046 22998 49164 23116
rect 55813 22992 55931 23110
rect 59555 23015 59673 23133
rect 84288 23123 84406 23241
rect 88643 23125 88761 23243
rect 65692 22987 65810 23105
rect 67640 22992 67758 23110
rect 74332 22990 74450 23108
rect 77070 23005 77188 23123
rect 90859 23123 90977 23241
rect 80010 22999 80128 23117
rect 82029 22990 82147 23108
rect 36565 20987 36693 21115
rect 41572 20990 41690 21108
rect 45918 20990 46036 21108
rect 47715 20991 47833 21109
rect 49570 21009 49688 21127
rect 55813 20995 55931 21113
rect 59555 20996 59673 21114
rect 64422 20993 64540 21111
rect 67640 20753 67758 20871
rect 74332 20507 74450 20625
rect 41572 20048 41690 20166
rect 47715 20048 47833 20166
rect 48344 20053 48462 20171
rect 84288 20090 84406 20208
rect 90859 20090 90977 20208
rect 92040 20036 92246 20242
rect 67637 19527 67755 19645
rect 74330 19293 74448 19411
rect 38285 19010 38403 19128
rect 41572 19000 41690 19118
rect 45223 18998 45341 19116
rect 45909 18998 46027 19116
rect 47715 18991 47833 19109
rect 49046 19025 49164 19143
rect 55826 18994 55944 19112
rect 58184 18995 58302 19113
rect 65692 18994 65810 19112
rect 87767 18719 87885 18837
rect 88626 18719 88744 18837
rect 93210 18719 93328 18837
rect 55826 17971 55944 18089
rect 56821 17971 56939 18089
rect 84288 17161 84406 17279
rect 38285 16975 38403 17093
rect 45909 17009 46027 17127
rect 49570 16997 49688 17115
rect 55826 16991 55944 17109
rect 58184 17039 58302 17157
rect 88626 17155 88744 17273
rect 90859 17156 90977 17274
rect 64422 16994 64540 17112
rect 67638 16995 67756 17113
rect 74330 17005 74448 17123
rect 78343 17003 78461 17121
rect 80949 17006 81067 17124
rect 82030 17005 82148 17123
rect 82030 16261 82148 16379
rect 88626 16305 88744 16423
rect 71861 -2153 71989 -2025
rect 72403 -2154 72531 -2026
rect 72947 -2153 73075 -2025
rect 73486 -2154 73614 -2026
rect 75127 -2153 75255 -2025
rect 75663 -2154 75791 -2026
rect 76213 -2153 76341 -2025
rect 76749 -2154 76877 -2026
rect 79480 -2154 79608 -2026
rect 80017 -2153 80145 -2025
rect 80562 -2155 80690 -2027
rect 81110 -2154 81238 -2026
rect 82738 -2154 82866 -2026
rect 83284 -2154 83412 -2026
rect 83835 -2153 83963 -2025
rect 84366 -2154 84494 -2026
<< metal2 >>
rect 103391 71867 104426 71889
rect 36373 71835 37373 71844
rect 36373 70826 37373 70835
rect 43351 71817 44375 71828
rect 43351 70817 43364 71817
rect 44364 70817 44375 71817
rect 43351 70806 44375 70817
rect 57794 71821 58825 71840
rect 57794 70821 57809 71821
rect 58809 70821 58825 71821
rect 74871 71807 75895 71820
rect 57794 70802 58825 70821
rect 64867 71771 65896 71786
rect 64867 70771 64881 71771
rect 65881 70771 65896 71771
rect 74871 70807 74883 71807
rect 75883 70807 75895 71807
rect 94051 71783 95086 71805
rect 74871 70796 75895 70807
rect 85821 71759 86856 71781
rect 64867 70758 65896 70771
rect 85821 70759 85838 71759
rect 86838 70759 86856 71759
rect 94051 70783 94068 71783
rect 95068 70783 95086 71783
rect 103391 70867 103408 71867
rect 104408 70867 104426 71867
rect 103391 70852 104426 70867
rect 94051 70768 95086 70783
rect 85821 70744 86856 70759
rect 36789 66748 36795 66876
rect 36923 66748 36929 66876
rect 36795 55845 36923 66748
rect 43789 66688 43795 66816
rect 43923 66688 43929 66816
rect 43795 57231 43923 66688
rect 38703 57103 38709 57231
rect 38837 57103 38843 57231
rect 43789 57103 43795 57231
rect 43923 57103 43929 57231
rect 82641 57103 82647 57231
rect 82775 57103 82781 57231
rect 36789 55717 36795 55845
rect 36923 55717 36929 55845
rect 36795 50626 36923 55717
rect 36795 50492 36923 50498
rect 38709 50628 38837 57103
rect 80619 55717 80625 55845
rect 80753 55717 80759 55845
rect 48935 54333 48941 54451
rect 49059 54333 49065 54451
rect 48941 52517 49059 54333
rect 48941 52393 49059 52399
rect 48730 51289 48873 51297
rect 38709 50494 38837 50500
rect 46751 51281 46879 51287
rect 48730 51161 48737 51289
rect 48865 51161 48873 51289
rect 48730 51154 48873 51161
rect 38692 49353 38820 49363
rect 36693 49338 36821 49348
rect 36693 48424 36821 49210
rect 36687 48296 36693 48424
rect 36821 48296 36827 48424
rect 36693 40605 36821 48296
rect 38692 47294 38820 49225
rect 46751 48424 46879 51153
rect 46745 48296 46751 48424
rect 46879 48296 46885 48424
rect 38680 47288 38820 47294
rect 48737 47288 48865 51154
rect 38808 47160 38820 47288
rect 48731 47160 48737 47288
rect 48865 47160 48871 47288
rect 38680 47154 38820 47160
rect 38692 45557 38820 47154
rect 38692 45423 38820 45429
rect 44965 45557 45093 45563
rect 44965 40528 45093 45429
rect 80625 41373 80753 55717
rect 82647 41389 82775 57103
rect 87250 54450 87368 54456
rect 85339 53292 85345 53410
rect 85463 53292 85469 53410
rect 85345 43190 85463 53292
rect 85339 43072 85345 43190
rect 85463 43072 85469 43190
rect 87250 43186 87368 54332
rect 116367 50862 116419 50910
rect 116334 49381 116452 50862
rect 116911 50850 116963 50914
rect 116873 50236 116991 50850
rect 116867 50118 116873 50236
rect 116991 50118 116997 50236
rect 120335 49387 120453 50858
rect 120884 50236 121002 50864
rect 126619 50236 126751 50243
rect 120878 50118 120884 50236
rect 121002 50118 121008 50236
rect 126619 50118 126626 50236
rect 126744 50118 126751 50236
rect 126619 50111 126751 50118
rect 120328 49381 120460 49387
rect 116328 49263 116334 49381
rect 116452 49263 116458 49381
rect 120328 49263 120335 49381
rect 120453 49263 120460 49381
rect 125951 49263 125957 49381
rect 126075 49263 126081 49381
rect 120328 49256 120460 49263
rect 87244 43068 87250 43186
rect 87368 43068 87374 43186
rect 82647 41255 82775 41261
rect 85240 41968 85368 41974
rect 80625 41239 80753 41245
rect 36693 40468 36821 40477
rect 44956 40400 44965 40528
rect 45093 40400 45102 40528
rect 80633 40168 80780 40176
rect 80633 40040 80643 40168
rect 80771 40040 80780 40168
rect 80633 40033 80780 40040
rect 82639 40034 82645 40162
rect 82773 40034 82779 40162
rect 40699 39232 40931 39246
rect 40699 39026 40712 39232
rect 40918 39026 40931 39232
rect 51827 39026 51833 39232
rect 52039 39026 52045 39232
rect 40699 39012 40931 39026
rect 50201 35813 50433 35828
rect 50201 35607 50215 35813
rect 50421 35607 50433 35813
rect 50201 35594 50433 35607
rect 51833 34367 52039 39026
rect 80643 38567 80771 40033
rect 82645 39407 82773 40034
rect 82645 39273 82773 39279
rect 85240 38567 85368 41840
rect 87247 41957 87375 41963
rect 86317 39417 86445 39423
rect 87247 39407 87375 41829
rect 113191 39618 117167 39736
rect 82304 38439 82310 38567
rect 82438 38439 82444 38567
rect 85234 38439 85240 38567
rect 85368 38439 85374 38567
rect 80643 38433 80771 38439
rect 54340 35813 54546 35819
rect 54340 35601 54546 35607
rect 67224 34846 68039 35053
rect 36565 34277 36693 34282
rect 36561 34159 36570 34277
rect 36688 34159 36697 34277
rect 44800 34263 44918 34268
rect 36565 23148 36693 34159
rect 44796 34155 44805 34263
rect 44913 34155 44922 34263
rect 51833 34171 51838 34367
rect 52034 34171 52039 34367
rect 51833 34166 52039 34171
rect 51838 34162 52034 34166
rect 39593 31145 39711 31154
rect 38279 27634 38285 27752
rect 38403 27634 38409 27752
rect 36559 23142 36699 23148
rect 36559 23014 36565 23142
rect 36693 23014 36699 23142
rect 36559 23008 36699 23014
rect 36565 21124 36693 23008
rect 36554 21115 36700 21124
rect 36554 20987 36565 21115
rect 36693 20987 36700 21115
rect 36554 20977 36700 20987
rect 38285 19128 38403 27634
rect 39593 24596 39711 31027
rect 44800 27752 44918 34155
rect 67550 33792 67668 34846
rect 67550 33668 67668 33674
rect 82310 33331 82438 38439
rect 86317 37663 86445 39289
rect 87241 39279 87247 39407
rect 87375 39279 87381 39407
rect 85315 37535 85321 37663
rect 85449 37535 85455 37663
rect 83771 34890 83928 34908
rect 83771 34762 83785 34890
rect 83913 34762 83928 34890
rect 83771 34736 83928 34762
rect 83813 33792 83961 33810
rect 83813 33674 83827 33792
rect 83945 33674 83961 33792
rect 83813 33655 83961 33674
rect 82310 33194 82438 33203
rect 85321 33320 85449 37535
rect 86317 37529 86445 37535
rect 86367 35894 86373 36022
rect 86501 35894 86507 36022
rect 86373 35338 86501 35894
rect 89481 35852 89487 36058
rect 89693 35852 89699 36058
rect 89487 35532 89693 35852
rect 86360 35325 86514 35338
rect 89483 35336 89492 35532
rect 89688 35336 89697 35532
rect 89487 35331 89693 35336
rect 86360 35197 86373 35325
rect 86501 35197 86514 35325
rect 86360 35183 86514 35197
rect 108254 35014 108372 35020
rect 110866 35014 110984 35020
rect 113191 35014 113309 39618
rect 117049 38289 117167 39618
rect 88556 34918 88762 34924
rect 108372 34896 110866 35014
rect 110984 34896 113309 35014
rect 108254 34890 108372 34896
rect 110866 34890 110984 34896
rect 88556 34379 88762 34712
rect 125957 34488 126075 49263
rect 88552 34183 88561 34379
rect 88757 34183 88766 34379
rect 125951 34370 125957 34488
rect 126075 34370 126081 34488
rect 88556 34178 88762 34183
rect 85321 33183 85449 33192
rect 88643 33792 88761 33798
rect 126626 33700 126744 50111
rect 81834 31877 81976 31890
rect 77064 31759 77070 31877
rect 77188 31759 77194 31877
rect 81834 31759 81847 31877
rect 81965 31759 81976 31877
rect 84866 31850 84984 31879
rect 42059 27634 42065 27752
rect 42183 27634 42189 27752
rect 44800 27628 44918 27634
rect 46166 31025 46284 31034
rect 46166 26341 46284 30907
rect 67550 27921 67668 27927
rect 45217 26223 45223 26341
rect 45341 26223 45347 26341
rect 39587 24478 39593 24596
rect 39711 24478 39717 24596
rect 41566 20990 41572 21108
rect 41690 20990 41696 21108
rect 41572 20166 41690 20990
rect 38279 19010 38285 19128
rect 38403 19010 38409 19128
rect 41572 19118 41690 20048
rect 38285 17093 38403 19010
rect 41566 19000 41572 19118
rect 41690 19000 41696 19118
rect 45223 19116 45341 26223
rect 46166 26217 46284 26223
rect 48344 27628 48462 27638
rect 45918 24596 46036 24602
rect 45918 23112 46036 24478
rect 45918 21108 46036 22994
rect 47709 20991 47715 21109
rect 47833 20991 47839 21109
rect 45918 20984 46036 20990
rect 47715 20166 47833 20991
rect 48344 20171 48462 27510
rect 55813 26993 55931 26999
rect 49046 23116 49164 23122
rect 55813 23110 55931 26875
rect 56815 26081 56821 26199
rect 56939 26081 56945 26199
rect 47709 20048 47715 20166
rect 47833 20048 47839 20166
rect 48338 20053 48344 20171
rect 48462 20053 48468 20171
rect 45909 19116 46027 19122
rect 45217 18998 45223 19116
rect 45341 18998 45347 19116
rect 47715 19109 47833 20048
rect 49046 19143 49164 22998
rect 55807 22992 55813 23110
rect 55931 22992 55937 23110
rect 49570 21127 49688 21133
rect 55813 21113 55931 22992
rect 45909 17127 46027 18998
rect 47709 18991 47715 19109
rect 47833 18991 47839 19109
rect 49040 19025 49046 19143
rect 49164 19025 49170 19143
rect 38279 16975 38285 17093
rect 38403 16975 38409 17093
rect 45909 17003 46027 17009
rect 49570 17115 49688 21009
rect 55807 20995 55813 21113
rect 55931 20995 55937 21113
rect 55820 18994 55826 19112
rect 55944 18994 55950 19112
rect 55826 18089 55944 18994
rect 56821 18089 56939 26081
rect 67550 25335 67668 27803
rect 69183 27908 69301 27914
rect 58178 25217 58184 25335
rect 58302 25217 58308 25335
rect 67544 25217 67550 25335
rect 67668 25217 67674 25335
rect 58184 19113 58302 25217
rect 59555 24414 59673 24420
rect 69183 24414 69301 27790
rect 69177 24296 69183 24414
rect 69301 24296 69307 24414
rect 59555 23133 59673 24296
rect 77070 23123 77188 31759
rect 81834 31746 81976 31759
rect 84836 31840 84984 31850
rect 84954 31722 84984 31840
rect 84836 31712 84984 31722
rect 82222 31330 82358 31343
rect 82222 31222 82236 31330
rect 82344 31222 82358 31330
rect 82222 31211 82358 31222
rect 78337 29252 78343 29370
rect 78461 29252 78467 29370
rect 59555 21114 59673 23015
rect 65692 23105 65810 23111
rect 59555 20990 59673 20996
rect 64416 20993 64422 21111
rect 64540 20993 64546 21111
rect 56815 17971 56821 18089
rect 56939 17971 56945 18089
rect 55826 17109 55944 17971
rect 58184 17157 58302 18995
rect 49570 16991 49688 16997
rect 55820 16991 55826 17109
rect 55944 16991 55950 17109
rect 58178 17039 58184 17157
rect 58302 17039 58308 17157
rect 64422 17112 64540 20993
rect 65692 19112 65810 22987
rect 67640 23110 67758 23120
rect 67640 20871 67758 22992
rect 67640 20743 67758 20753
rect 74332 23108 74450 23118
rect 77070 22999 77188 23005
rect 74332 20625 74450 22990
rect 74332 20497 74450 20507
rect 65692 18988 65810 18994
rect 67637 19645 67755 19655
rect 64422 16988 64540 16994
rect 67637 17123 67755 19527
rect 74324 19293 74330 19411
rect 74448 19293 74454 19411
rect 74330 17123 74448 19293
rect 67637 17113 67756 17123
rect 67637 16995 67638 17113
rect 74330 16999 74448 17005
rect 78343 17121 78461 29252
rect 82231 28361 82349 31211
rect 84866 29370 84984 31712
rect 85787 31831 85919 31850
rect 85787 31723 85799 31831
rect 85907 31723 85919 31831
rect 85787 31709 85919 31723
rect 86778 31819 86965 31853
rect 84860 29252 84866 29370
rect 84984 29252 84990 29370
rect 80010 28351 80128 28357
rect 80010 23117 80128 28233
rect 82222 28351 82355 28361
rect 82222 28233 82231 28351
rect 82349 28233 82355 28351
rect 82222 28226 82355 28233
rect 82231 28220 82349 28226
rect 80949 27142 81067 27148
rect 80004 22999 80010 23117
rect 80128 22999 80134 23117
rect 78343 16997 78461 17003
rect 80949 17124 81067 27024
rect 85794 27142 85912 31709
rect 86778 31701 86818 31819
rect 86936 31701 86965 31819
rect 86778 31671 86965 31701
rect 87767 31819 87885 31825
rect 85794 27018 85912 27024
rect 82023 24304 82029 24422
rect 82147 24304 82153 24422
rect 82029 23108 82147 24304
rect 84288 23241 84406 23247
rect 82023 22990 82029 23108
rect 82147 22990 82153 23108
rect 84288 20218 84406 23123
rect 84278 20208 84416 20218
rect 84278 20090 84288 20208
rect 84406 20090 84416 20208
rect 84278 20084 84416 20090
rect 84288 17279 84406 20084
rect 87767 18837 87885 31701
rect 88643 26607 88761 33674
rect 126620 33582 126626 33700
rect 126744 33582 126750 33700
rect 107303 33517 107421 33523
rect 107421 33399 113269 33517
rect 107303 33393 107421 33399
rect 110866 32825 110984 32831
rect 107303 32812 107421 32821
rect 107297 32694 107303 32812
rect 107421 32694 107427 32812
rect 110857 32707 110866 32825
rect 110984 32707 110993 32825
rect 110866 32701 110984 32707
rect 107303 32685 107421 32694
rect 113151 28435 113269 33399
rect 117180 28437 117298 29684
rect 113620 28435 117298 28437
rect 110894 28334 111002 28338
rect 107294 28315 107428 28322
rect 107294 28197 107303 28315
rect 107421 28197 107428 28315
rect 110883 28216 110889 28334
rect 111007 28216 111013 28334
rect 113151 28319 117298 28435
rect 113151 28317 113697 28319
rect 110894 28212 111002 28216
rect 107294 28184 107428 28197
rect 92034 27813 92040 28019
rect 92246 27813 92252 28019
rect 93376 27813 93382 28019
rect 93588 27813 93594 28019
rect 88637 26489 88643 26607
rect 88761 26489 88767 26607
rect 88643 24435 88761 26489
rect 88637 24317 88643 24435
rect 88761 24317 88767 24435
rect 88643 23243 88761 24317
rect 88637 23125 88643 23243
rect 88761 23125 88767 23243
rect 90853 23123 90859 23241
rect 90977 23123 90983 23241
rect 90859 20208 90977 23123
rect 92040 20242 92246 27813
rect 93210 25170 93328 25176
rect 90853 20090 90859 20208
rect 90977 20090 90983 20208
rect 87767 18713 87885 18719
rect 88626 18837 88744 18843
rect 84288 17155 84406 17161
rect 88626 17273 88744 18719
rect 90859 17274 90977 20090
rect 92034 20036 92040 20242
rect 92246 20036 92252 20242
rect 93210 18837 93328 25052
rect 93204 18719 93210 18837
rect 93328 18719 93334 18837
rect 90853 17156 90859 17274
rect 90977 17156 90983 17274
rect 80949 17000 81067 17006
rect 82020 17123 82160 17137
rect 82020 17005 82030 17123
rect 82148 17005 82160 17123
rect 67637 16990 67756 16995
rect 82020 16993 82160 17005
rect 67638 16985 67756 16990
rect 82030 16379 82148 16993
rect 88626 16423 88744 17155
rect 82024 16261 82030 16379
rect 82148 16261 82154 16379
rect 88620 16305 88626 16423
rect 88744 16305 88750 16423
rect 71851 -2153 71861 -2025
rect 71989 -2153 71999 -2025
rect 72393 -2154 72403 -2026
rect 72531 -2154 72541 -2026
rect 72937 -2153 72947 -2025
rect 73075 -2153 73085 -2025
rect 73476 -2154 73486 -2026
rect 73614 -2154 73624 -2026
rect 75117 -2153 75127 -2025
rect 75255 -2153 75265 -2025
rect 75653 -2154 75663 -2026
rect 75791 -2154 75801 -2026
rect 76203 -2153 76213 -2025
rect 76341 -2153 76351 -2025
rect 76739 -2154 76749 -2026
rect 76877 -2154 76887 -2026
rect 79470 -2154 79480 -2026
rect 79608 -2154 79618 -2026
rect 80007 -2153 80017 -2025
rect 80145 -2153 80155 -2025
rect 80552 -2155 80562 -2027
rect 80690 -2155 80700 -2027
rect 81100 -2154 81110 -2026
rect 81238 -2154 81248 -2026
rect 82728 -2154 82738 -2026
rect 82866 -2154 82876 -2026
rect 83274 -2154 83284 -2026
rect 83412 -2154 83422 -2026
rect 83825 -2153 83835 -2025
rect 83963 -2153 83973 -2025
rect 84356 -2154 84366 -2026
rect 84494 -2154 84504 -2026
<< via2 >>
rect 36373 70835 37373 71835
rect 43364 70817 44364 71817
rect 57809 70821 58809 71821
rect 64881 70771 65881 71771
rect 74883 70807 75883 71807
rect 85838 70759 86838 71759
rect 94068 70783 95068 71783
rect 103408 70867 104408 71867
rect 36693 40477 36821 40605
rect 44965 40400 45093 40528
rect 40712 39026 40918 39232
rect 50215 35607 50421 35813
rect 54345 35612 54541 35808
rect 36570 34159 36688 34277
rect 44805 34155 44913 34263
rect 51838 34171 52034 34367
rect 39593 31027 39711 31145
rect 83785 34762 83913 34890
rect 83827 33674 83945 33792
rect 82310 33203 82438 33331
rect 89492 35336 89688 35532
rect 86373 35197 86501 35325
rect 88561 34183 88757 34379
rect 85321 33192 85449 33320
rect 81847 31759 81965 31877
rect 46166 30907 46284 31025
rect 48344 27510 48462 27628
rect 84836 31722 84954 31840
rect 82236 31222 82344 31330
rect 85799 31723 85907 31831
rect 86818 31701 86936 31819
rect 107303 32694 107421 32812
rect 110866 32707 110984 32825
rect 107308 28202 107416 28310
rect 110894 28221 111002 28329
rect 93387 27818 93583 28014
rect 71861 -2153 71989 -2025
rect 72403 -2154 72531 -2026
rect 72947 -2153 73075 -2025
rect 73486 -2154 73614 -2026
rect 75127 -2153 75255 -2025
rect 75663 -2154 75791 -2026
rect 76213 -2153 76341 -2025
rect 76749 -2154 76877 -2026
rect 79480 -2154 79608 -2026
rect 80017 -2153 80145 -2025
rect 80562 -2155 80690 -2027
rect 81110 -2154 81238 -2026
rect 82738 -2154 82866 -2026
rect 83284 -2154 83412 -2026
rect 83835 -2153 83963 -2025
rect 84366 -2154 84494 -2026
<< metal3 >>
rect 36373 71840 37373 87729
rect 36368 71835 37378 71840
rect 36368 70835 36373 71835
rect 37373 70835 37378 71835
rect 43364 71822 44364 87636
rect 57809 71826 58809 75167
rect 36368 70830 37378 70835
rect 43359 71817 44369 71822
rect 43359 70817 43364 71817
rect 44364 70817 44369 71817
rect 43359 70812 44369 70817
rect 57804 71821 58814 71826
rect 57804 70821 57809 71821
rect 58809 70821 58814 71821
rect 64881 71776 65881 75198
rect 74883 71812 75883 74992
rect 74878 71807 75888 71812
rect 57804 70816 58814 70821
rect 64876 71771 65886 71776
rect 64876 70771 64881 71771
rect 65881 70771 65886 71771
rect 74878 70807 74883 71807
rect 75883 70807 75888 71807
rect 85838 71764 86838 74971
rect 94068 71788 95068 74995
rect 103408 71872 104408 75079
rect 103403 71867 104413 71872
rect 94063 71783 95073 71788
rect 74878 70802 75888 70807
rect 85833 71759 86843 71764
rect 64876 70766 65886 70771
rect 85833 70759 85838 71759
rect 86838 70759 86843 71759
rect 94063 70783 94068 71783
rect 95068 70783 95073 71783
rect 103403 70867 103408 71867
rect 104408 70867 104413 71867
rect 103403 70862 104413 70867
rect 94063 70778 95073 70783
rect 85833 70754 86843 70759
rect 33473 41686 38293 41750
rect 43345 41677 44585 41741
rect 46545 41602 47958 41666
rect 33296 33165 33360 41532
rect 36678 40610 36834 40618
rect 36678 40472 36688 40610
rect 36826 40472 36834 40610
rect 36678 40464 36834 40472
rect 38633 39962 38697 41321
rect 42833 39962 42897 41202
rect 44947 40533 45108 40541
rect 44947 40395 44960 40533
rect 45098 40395 45108 40533
rect 44947 40385 45108 40395
rect 40699 39237 40931 39246
rect 40699 39021 40707 39237
rect 40923 39021 40931 39237
rect 40699 39012 40931 39021
rect 36482 36762 36546 38002
rect 38633 36762 38697 38002
rect 42833 36762 42897 38002
rect 44984 36762 45048 38002
rect 36565 34277 36693 34855
rect 36565 34159 36570 34277
rect 36688 34159 36693 34277
rect 36565 34154 36693 34159
rect 38633 33562 38697 34802
rect 42833 33443 42897 34802
rect 44800 34263 44918 34842
rect 44800 34155 44805 34263
rect 44913 34155 44918 34263
rect 44800 34143 44918 34155
rect 48170 33232 48234 41599
rect 50201 35818 50433 35828
rect 50201 35602 50210 35818
rect 50426 35602 50433 35818
rect 56624 35813 56828 35818
rect 54340 35812 56829 35813
rect 54340 35808 56624 35812
rect 54340 35612 54345 35808
rect 54541 35612 56624 35808
rect 54340 35608 56624 35612
rect 56828 35608 56829 35812
rect 54340 35607 56829 35608
rect 56624 35602 56828 35607
rect 50201 35594 50433 35602
rect 82555 34935 82619 35541
rect 83771 34895 83928 34908
rect 83771 34757 83780 34895
rect 83918 34757 83928 34895
rect 85567 34894 85631 35655
rect 91354 35537 91558 35542
rect 94546 35537 94752 35543
rect 89487 35536 91559 35537
rect 89487 35532 91354 35536
rect 86360 35330 86514 35338
rect 89487 35336 89492 35532
rect 89688 35336 91354 35532
rect 89487 35332 91354 35336
rect 91558 35332 91559 35536
rect 89487 35331 91559 35332
rect 86360 35192 86368 35330
rect 86506 35192 86514 35330
rect 91354 35326 91558 35331
rect 94546 35325 94752 35331
rect 86360 35183 86514 35192
rect 83771 34736 83928 34757
rect 56642 34372 56846 34377
rect 60430 34372 60636 34682
rect 81528 34563 83251 34627
rect 51833 34371 56847 34372
rect 51833 34367 56642 34371
rect 51833 34171 51838 34367
rect 52034 34171 56642 34367
rect 51833 34167 56642 34171
rect 56846 34167 56847 34371
rect 51833 34166 56847 34167
rect 56642 34161 56846 34166
rect 60430 34160 60636 34166
rect 33572 33098 34985 33162
rect 36945 33023 38185 33087
rect 43237 33014 48057 33078
rect 39593 31150 39711 31797
rect 39588 31145 39716 31150
rect 39588 31027 39593 31145
rect 39711 31027 39716 31145
rect 46166 31030 46284 31861
rect 39588 31022 39716 31027
rect 46161 31025 46289 31030
rect 46161 30907 46166 31025
rect 46284 30907 46289 31025
rect 46161 30902 46289 30907
rect 81512 30938 81576 34535
rect 82649 33707 82859 33771
rect 82305 33331 82443 33336
rect 82305 33203 82310 33331
rect 82438 33203 82443 33331
rect 82305 33198 82443 33203
rect 82310 32974 82438 33198
rect 81834 31877 81976 31890
rect 81834 31759 81847 31877
rect 81965 31759 82184 31877
rect 82790 31796 82854 33707
rect 81834 31746 81976 31759
rect 82619 31732 82854 31796
rect 82222 31334 82358 31343
rect 82222 31218 82232 31334
rect 82348 31218 82358 31334
rect 82222 31211 82358 31218
rect 83187 30938 83251 34563
rect 84505 34572 86244 34636
rect 83813 33792 83961 33810
rect 83598 33674 83827 33792
rect 83945 33674 83961 33792
rect 83813 33655 83961 33674
rect 81512 30874 83251 30938
rect 84505 30947 84569 34572
rect 84862 33707 85097 33771
rect 84862 31845 84926 33707
rect 85316 33320 85454 33325
rect 85316 33192 85321 33320
rect 85449 33192 85454 33320
rect 85316 33187 85454 33192
rect 85321 32989 85449 33187
rect 84826 31840 84964 31845
rect 84826 31722 84836 31840
rect 84954 31804 84964 31840
rect 85787 31835 85919 31850
rect 84954 31740 85090 31804
rect 84954 31722 84964 31740
rect 84826 31717 84964 31722
rect 85787 31719 85795 31835
rect 85911 31719 85919 31835
rect 85787 31709 85919 31719
rect 86180 30975 86244 34572
rect 91312 34384 91516 34389
rect 94946 34384 95152 34765
rect 88556 34383 91517 34384
rect 88556 34379 91312 34383
rect 88556 34183 88561 34379
rect 88757 34183 91312 34379
rect 88556 34179 91312 34183
rect 91516 34179 91517 34383
rect 88556 34178 91517 34179
rect 91312 34173 91516 34178
rect 94946 34172 95152 34178
rect 107284 32817 107438 32834
rect 107284 32689 107298 32817
rect 107426 32689 107438 32817
rect 110861 32825 110871 32830
rect 110861 32707 110866 32825
rect 110861 32702 110871 32707
rect 110989 32702 110995 32830
rect 107284 32681 107438 32689
rect 86778 31819 86965 31853
rect 86610 31701 86818 31819
rect 86936 31701 86965 31819
rect 86778 31671 86965 31701
rect 84505 30883 86228 30947
rect 82529 30047 82593 30470
rect 85524 29897 85588 30658
rect 58866 27670 59072 28849
rect 93382 28014 93588 28779
rect 110890 28334 111006 28339
rect 110889 28333 111007 28334
rect 107294 28314 107428 28322
rect 107294 28198 107304 28314
rect 107420 28198 107428 28314
rect 110889 28217 110890 28333
rect 111006 28217 111007 28333
rect 110889 28216 111007 28217
rect 110890 28211 111006 28216
rect 107294 28184 107428 28198
rect 93382 27818 93387 28014
rect 93583 27818 93588 28014
rect 93382 27813 93588 27818
rect 48295 27628 59072 27670
rect 48295 27510 48344 27628
rect 48462 27510 59072 27628
rect 48295 27464 59072 27510
rect 24674 13863 132085 13991
rect 71856 12350 71862 12351
rect 24674 12225 71862 12350
rect 71988 12350 71994 12351
rect 71988 12225 132085 12350
rect 24674 12222 132085 12225
rect 24674 11682 72404 11808
rect 72530 11682 132085 11808
rect 24674 11680 132085 11682
rect 24674 11136 72947 11264
rect 73075 11136 132085 11264
rect 24674 10720 132085 10725
rect 24674 10597 73487 10720
rect 73481 10594 73487 10597
rect 73613 10597 132085 10720
rect 73613 10594 73619 10597
rect 24674 9083 132085 9084
rect 24674 8957 75128 9083
rect 75254 8957 132085 9083
rect 24674 8956 132085 8957
rect 75658 8548 75664 8549
rect 24674 8423 75664 8548
rect 75790 8548 75796 8549
rect 75790 8423 132085 8548
rect 24674 8420 132085 8423
rect 76208 7998 76214 8001
rect 24674 7875 76214 7998
rect 76340 7998 76346 8001
rect 76340 7875 132085 7998
rect 24674 7870 132085 7875
rect 24674 7459 132085 7462
rect 24674 7334 76750 7459
rect 76744 7333 76750 7334
rect 76876 7334 132085 7459
rect 76876 7333 76882 7334
rect 24674 5820 132085 5821
rect 24674 5694 79481 5820
rect 79607 5694 132085 5820
rect 24674 5693 132085 5694
rect 24674 5158 80018 5284
rect 80144 5158 132085 5284
rect 24674 5156 132085 5158
rect 80557 4739 80563 4749
rect 24674 4623 80563 4739
rect 80689 4739 80695 4749
rect 80689 4623 132085 4739
rect 24674 4611 132085 4623
rect 24674 4185 132085 4191
rect 24674 4063 81111 4185
rect 81105 4059 81111 4063
rect 81237 4063 132085 4185
rect 81237 4059 81243 4063
rect 24674 2562 132085 2563
rect 24674 2436 82739 2562
rect 82865 2436 132085 2562
rect 24674 2435 132085 2436
rect 83279 2017 83285 2019
rect 24674 1893 83285 2017
rect 83411 2017 83417 2019
rect 83411 1893 132085 2017
rect 24674 1889 132085 1893
rect 83830 1466 83836 1471
rect 24674 1345 83836 1466
rect 83962 1466 83968 1471
rect 83962 1345 132085 1466
rect 24674 1338 132085 1345
rect 24674 929 132085 935
rect 24674 807 84367 929
rect 84361 803 84367 807
rect 84493 807 132085 929
rect 84493 803 84499 807
rect 71861 -2015 71989 -2011
rect 71856 -2024 71994 -2015
rect 72403 -2016 72531 -2011
rect 72947 -2015 73075 -2011
rect 71856 -2153 71861 -2024
rect 71989 -2153 71994 -2024
rect 71856 -2163 71994 -2153
rect 72398 -2026 72536 -2016
rect 72398 -2158 72403 -2026
rect 72531 -2158 72536 -2026
rect 72398 -2164 72536 -2158
rect 72942 -2025 73080 -2015
rect 73486 -2016 73614 -2011
rect 75127 -2015 75255 -2011
rect 72942 -2155 72947 -2025
rect 73075 -2155 73080 -2025
rect 72942 -2163 73080 -2155
rect 73481 -2026 73619 -2016
rect 73481 -2158 73486 -2026
rect 73614 -2158 73619 -2026
rect 73481 -2164 73619 -2158
rect 75122 -2025 75260 -2015
rect 75663 -2016 75791 -2011
rect 76213 -2015 76341 -2011
rect 75122 -2155 75127 -2025
rect 75255 -2155 75260 -2025
rect 75122 -2163 75260 -2155
rect 75658 -2024 75796 -2016
rect 75658 -2154 75663 -2024
rect 75791 -2154 75796 -2024
rect 75658 -2164 75796 -2154
rect 76208 -2024 76346 -2015
rect 76749 -2016 76877 -2011
rect 79480 -2016 79608 -2011
rect 80017 -2015 80145 -2011
rect 76208 -2153 76213 -2024
rect 76341 -2153 76346 -2024
rect 76208 -2163 76346 -2153
rect 76744 -2024 76882 -2016
rect 76744 -2154 76749 -2024
rect 76877 -2154 76882 -2024
rect 76744 -2164 76882 -2154
rect 79475 -2023 79613 -2016
rect 79475 -2154 79480 -2023
rect 79608 -2154 79613 -2023
rect 79475 -2164 79613 -2154
rect 80012 -2023 80150 -2015
rect 80562 -2017 80690 -2011
rect 81110 -2016 81238 -2011
rect 82738 -2016 82866 -2011
rect 83284 -2016 83412 -2011
rect 83835 -2015 83963 -2011
rect 80012 -2153 80017 -2023
rect 80145 -2153 80150 -2023
rect 80012 -2163 80150 -2153
rect 80557 -2027 80695 -2017
rect 80557 -2155 80562 -2027
rect 80690 -2155 80695 -2027
rect 80557 -2165 80695 -2155
rect 81105 -2026 81243 -2016
rect 81105 -2160 81110 -2026
rect 81238 -2160 81243 -2026
rect 81105 -2164 81243 -2160
rect 82733 -2026 82871 -2016
rect 82733 -2155 82738 -2026
rect 82866 -2155 82871 -2026
rect 82733 -2164 82871 -2155
rect 83279 -2026 83417 -2016
rect 83279 -2155 83284 -2026
rect 83412 -2155 83417 -2026
rect 83279 -2164 83417 -2155
rect 83830 -2025 83968 -2015
rect 84366 -2016 84494 -2011
rect 83830 -2155 83835 -2025
rect 83963 -2155 83968 -2025
rect 83830 -2163 83968 -2155
rect 84361 -2023 84499 -2016
rect 84361 -2154 84366 -2023
rect 84494 -2154 84499 -2023
rect 84361 -2164 84499 -2154
rect 81110 -2166 81238 -2164
<< via3 >>
rect 36688 40605 36826 40610
rect 36688 40477 36693 40605
rect 36693 40477 36821 40605
rect 36821 40477 36826 40605
rect 36688 40472 36826 40477
rect 44960 40528 45098 40533
rect 44960 40400 44965 40528
rect 44965 40400 45093 40528
rect 45093 40400 45098 40528
rect 44960 40395 45098 40400
rect 40707 39232 40923 39237
rect 40707 39026 40712 39232
rect 40712 39026 40918 39232
rect 40918 39026 40923 39232
rect 40707 39021 40923 39026
rect 50210 35813 50426 35818
rect 50210 35607 50215 35813
rect 50215 35607 50421 35813
rect 50421 35607 50426 35813
rect 50210 35602 50426 35607
rect 56624 35608 56828 35812
rect 60030 35607 60236 35813
rect 83780 34890 83918 34895
rect 83780 34762 83785 34890
rect 83785 34762 83913 34890
rect 83913 34762 83918 34890
rect 83780 34757 83918 34762
rect 91354 35332 91558 35536
rect 94546 35331 94752 35537
rect 86368 35325 86506 35330
rect 86368 35197 86373 35325
rect 86373 35197 86501 35325
rect 86501 35197 86506 35325
rect 86368 35192 86506 35197
rect 56642 34167 56846 34371
rect 60430 34166 60636 34372
rect 82232 31330 82348 31334
rect 82232 31222 82236 31330
rect 82236 31222 82344 31330
rect 82344 31222 82348 31330
rect 82232 31218 82348 31222
rect 85795 31831 85911 31835
rect 85795 31723 85799 31831
rect 85799 31723 85907 31831
rect 85907 31723 85911 31831
rect 85795 31719 85911 31723
rect 91312 34179 91516 34383
rect 94946 34178 95152 34384
rect 107298 32812 107426 32817
rect 107298 32694 107303 32812
rect 107303 32694 107421 32812
rect 107421 32694 107426 32812
rect 107298 32689 107426 32694
rect 110871 32825 110989 32830
rect 110871 32707 110984 32825
rect 110984 32707 110989 32825
rect 110871 32702 110989 32707
rect 107304 28310 107420 28314
rect 107304 28202 107308 28310
rect 107308 28202 107416 28310
rect 107416 28202 107420 28310
rect 107304 28198 107420 28202
rect 110890 28329 111006 28333
rect 110890 28221 110894 28329
rect 110894 28221 111002 28329
rect 111002 28221 111006 28329
rect 110890 28217 111006 28221
rect 71862 12225 71988 12351
rect 72404 11682 72530 11808
rect 72947 11136 73075 11264
rect 73487 10594 73613 10720
rect 75128 8957 75254 9083
rect 75664 8423 75790 8549
rect 76214 7875 76340 8001
rect 76750 7333 76876 7459
rect 79481 5694 79607 5820
rect 80018 5158 80144 5284
rect 80563 4623 80689 4749
rect 81111 4059 81237 4185
rect 82739 2436 82865 2562
rect 83285 1893 83411 2019
rect 83836 1345 83962 1471
rect 84367 803 84493 929
rect 71861 -2025 71989 -2024
rect 71861 -2152 71989 -2025
rect 72403 -2154 72531 -2030
rect 72403 -2158 72531 -2154
rect 72947 -2153 73075 -2027
rect 72947 -2155 73075 -2153
rect 73486 -2154 73614 -2030
rect 73486 -2158 73614 -2154
rect 75127 -2153 75255 -2027
rect 75127 -2155 75255 -2153
rect 75663 -2026 75791 -2024
rect 75663 -2152 75791 -2026
rect 76213 -2025 76341 -2024
rect 76213 -2152 76341 -2025
rect 76749 -2026 76877 -2024
rect 76749 -2152 76877 -2026
rect 79480 -2026 79608 -2023
rect 79480 -2151 79608 -2026
rect 80017 -2025 80145 -2023
rect 80017 -2151 80145 -2025
rect 80562 -2155 80690 -2027
rect 81110 -2154 81238 -2032
rect 81110 -2160 81238 -2154
rect 82738 -2154 82866 -2027
rect 82738 -2155 82866 -2154
rect 83284 -2154 83412 -2027
rect 83284 -2155 83412 -2154
rect 83835 -2153 83963 -2027
rect 83835 -2155 83963 -2153
rect 84366 -2026 84494 -2023
rect 84366 -2151 84494 -2026
<< metal4 >>
rect 43206 42670 44724 42734
rect 46406 42666 47956 42730
rect 33426 42574 38481 42638
rect 32097 33415 32161 41442
rect 36687 40610 36827 40611
rect 36687 40472 36688 40610
rect 36826 40472 36827 40610
rect 36687 40471 36827 40472
rect 36693 39678 36821 40471
rect 39642 39823 39706 41431
rect 41824 39823 41888 41341
rect 44959 40533 45099 40534
rect 44959 40395 44960 40533
rect 45098 40395 45099 40533
rect 44959 40394 45099 40395
rect 44965 39609 45093 40394
rect 40699 39237 40931 39246
rect 40699 39232 40707 39237
rect 39968 39026 40707 39232
rect 40699 39021 40707 39026
rect 40923 39021 40931 39237
rect 40699 39012 40931 39021
rect 35459 36623 35523 38141
rect 39642 36623 39706 38141
rect 41824 36623 41888 38141
rect 46007 36623 46071 38141
rect 49369 35888 49433 41349
rect 49315 35813 49570 35888
rect 50201 35818 50433 35828
rect 50201 35813 50210 35818
rect 49315 35682 50210 35813
rect 49369 35607 50210 35682
rect 39642 33423 39706 34941
rect 41824 33333 41888 34941
rect 49369 33322 49433 35607
rect 50201 35602 50210 35607
rect 50426 35602 50433 35818
rect 60029 35813 60237 35814
rect 56623 35812 60030 35813
rect 56623 35608 56624 35812
rect 56828 35608 60030 35812
rect 56623 35607 60030 35608
rect 60236 35607 60237 35813
rect 60029 35606 60237 35607
rect 50201 35594 50433 35602
rect 82211 34922 82275 35607
rect 81216 34918 83541 34922
rect 85220 34920 85284 35655
rect 94545 35537 94753 35538
rect 91353 35536 94546 35537
rect 86360 35330 86514 35338
rect 91353 35332 91354 35536
rect 91558 35332 94546 35536
rect 91353 35331 94546 35332
rect 94752 35331 94753 35537
rect 94545 35330 94753 35331
rect 86360 35192 86368 35330
rect 86506 35192 86514 35330
rect 86360 35183 86514 35192
rect 86373 34920 86501 35183
rect 81216 34890 83557 34918
rect 83771 34895 83928 34908
rect 83771 34890 83780 34895
rect 81216 34858 83780 34890
rect 60429 34372 60637 34373
rect 56641 34371 60430 34372
rect 56641 34167 56642 34371
rect 56846 34167 60430 34371
rect 56641 34166 60430 34167
rect 60636 34166 60637 34372
rect 60429 34165 60637 34166
rect 43049 32126 48104 32190
rect 33574 32034 35124 32098
rect 36806 32030 38324 32094
rect 81216 30850 81280 34858
rect 83471 34762 83780 34858
rect 83477 34712 83557 34762
rect 83771 34757 83780 34762
rect 83918 34757 83928 34895
rect 83771 34736 83928 34757
rect 84215 34856 86534 34920
rect 82259 31894 82323 33614
rect 82231 31334 82349 31636
rect 82231 31218 82232 31334
rect 82348 31218 82349 31334
rect 82231 31217 82349 31218
rect 83477 30654 83541 34712
rect 81222 30590 83541 30654
rect 84215 30652 84279 34856
rect 85433 31896 85497 33616
rect 85519 31835 85912 31836
rect 85519 31719 85795 31835
rect 85911 31719 85912 31835
rect 85519 31718 85912 31719
rect 86476 30652 86540 34660
rect 94945 34384 95153 34385
rect 91311 34383 94946 34384
rect 91311 34179 91312 34383
rect 91516 34179 94946 34383
rect 91311 34178 94946 34179
rect 95152 34178 95153 34384
rect 94945 34177 95153 34178
rect 110870 32830 110990 32831
rect 107297 32817 107427 32818
rect 107297 32689 107298 32817
rect 107426 32689 107427 32817
rect 110870 32702 110871 32830
rect 110989 32702 110990 32830
rect 110870 32701 110990 32702
rect 107297 32688 107427 32689
rect 82216 29893 82280 30590
rect 84215 30588 86540 30652
rect 85218 29886 85282 30588
rect 107303 28322 107421 32688
rect 110871 32026 110989 32701
rect 110889 28333 111007 29930
rect 107294 28314 107428 28322
rect 107294 28198 107304 28314
rect 107420 28198 107428 28314
rect 110889 28217 110890 28333
rect 111006 28217 111007 28333
rect 110889 28216 111007 28217
rect 107294 28184 107428 28198
rect 71861 12351 71989 12352
rect 71861 12225 71862 12351
rect 71988 12225 71989 12351
rect 71861 -2023 71989 12225
rect 72403 11808 72531 11809
rect 72403 11682 72404 11808
rect 72530 11682 72531 11808
rect 71860 -2024 71990 -2023
rect 71860 -2152 71861 -2024
rect 71989 -2152 71990 -2024
rect 72403 -2029 72531 11682
rect 72947 11265 73075 11266
rect 72946 11264 73076 11265
rect 72946 11136 72947 11264
rect 73075 11136 73076 11264
rect 72946 11135 73076 11136
rect 72947 -2026 73075 11135
rect 73486 10720 73614 10721
rect 73486 10594 73487 10720
rect 73613 10594 73614 10720
rect 72946 -2027 73076 -2026
rect 71860 -2153 71990 -2152
rect 72402 -2030 72532 -2029
rect 72402 -2158 72403 -2030
rect 72531 -2158 72532 -2030
rect 72946 -2155 72947 -2027
rect 73075 -2155 73076 -2027
rect 73486 -2029 73614 10594
rect 75127 9083 75255 9084
rect 75127 8957 75128 9083
rect 75254 8957 75255 9083
rect 75127 -2026 75255 8957
rect 75663 8549 75791 8550
rect 75663 8423 75664 8549
rect 75790 8423 75791 8549
rect 75663 -2023 75791 8423
rect 76213 8001 76341 8002
rect 76213 7875 76214 8001
rect 76340 7875 76341 8001
rect 76213 -2023 76341 7875
rect 76749 7459 76877 7460
rect 76749 7333 76750 7459
rect 76876 7333 76877 7459
rect 76749 -2023 76877 7333
rect 79480 5820 79608 5821
rect 79480 5694 79481 5820
rect 79607 5694 79608 5820
rect 79480 -2022 79608 5694
rect 80017 5284 80145 5285
rect 80017 5158 80018 5284
rect 80144 5158 80145 5284
rect 80017 -2022 80145 5158
rect 80562 4749 80690 4750
rect 80562 4623 80563 4749
rect 80689 4623 80690 4749
rect 79479 -2023 79609 -2022
rect 75662 -2024 75792 -2023
rect 75126 -2027 75256 -2026
rect 72946 -2156 73076 -2155
rect 73485 -2030 73615 -2029
rect 72402 -2159 72532 -2158
rect 73485 -2158 73486 -2030
rect 73614 -2158 73615 -2030
rect 75126 -2155 75127 -2027
rect 75255 -2155 75256 -2027
rect 75662 -2152 75663 -2024
rect 75791 -2152 75792 -2024
rect 75662 -2153 75792 -2152
rect 76212 -2024 76342 -2023
rect 76212 -2152 76213 -2024
rect 76341 -2152 76342 -2024
rect 76212 -2153 76342 -2152
rect 76748 -2024 76878 -2023
rect 76748 -2152 76749 -2024
rect 76877 -2152 76878 -2024
rect 79479 -2151 79480 -2023
rect 79608 -2151 79609 -2023
rect 79479 -2152 79609 -2151
rect 80016 -2023 80146 -2022
rect 80016 -2151 80017 -2023
rect 80145 -2151 80146 -2023
rect 80562 -2026 80690 4623
rect 81110 4185 81238 4186
rect 81110 4059 81111 4185
rect 81237 4059 81238 4185
rect 80016 -2152 80146 -2151
rect 80561 -2027 80691 -2026
rect 76748 -2153 76878 -2152
rect 75126 -2156 75256 -2155
rect 80561 -2155 80562 -2027
rect 80690 -2155 80691 -2027
rect 81110 -2031 81238 4059
rect 82738 2562 82866 2563
rect 82738 2436 82739 2562
rect 82865 2436 82866 2562
rect 82738 -2026 82866 2436
rect 83284 2019 83412 2020
rect 83284 1893 83285 2019
rect 83411 1893 83412 2019
rect 83284 -2026 83412 1893
rect 83835 1471 83963 1472
rect 83835 1345 83836 1471
rect 83962 1345 83963 1471
rect 83835 -2026 83963 1345
rect 84366 929 84494 930
rect 84366 803 84367 929
rect 84493 803 84494 929
rect 84366 -2022 84494 803
rect 84365 -2023 84495 -2022
rect 82737 -2027 82867 -2026
rect 80561 -2156 80691 -2155
rect 81109 -2032 81239 -2031
rect 73485 -2159 73615 -2158
rect 81109 -2160 81110 -2032
rect 81238 -2160 81239 -2032
rect 82737 -2155 82738 -2027
rect 82866 -2155 82867 -2027
rect 82737 -2156 82867 -2155
rect 83283 -2027 83413 -2026
rect 83283 -2155 83284 -2027
rect 83412 -2155 83413 -2027
rect 83283 -2156 83413 -2155
rect 83834 -2027 83964 -2026
rect 83834 -2155 83835 -2027
rect 83963 -2155 83964 -2027
rect 84365 -2151 84366 -2023
rect 84494 -2151 84495 -2023
rect 84365 -2152 84495 -2151
rect 83834 -2156 83964 -2155
rect 81109 -2161 81239 -2160
use a_mux2_en  a_mux2_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/a_mux2_en
timestamp 1654674840
transform 0 -1 84928 1 0 60716
box -2638 -2806 3466 243
use a_mux2_en  a_mux2_en_1
timestamp 1654674840
transform 0 -1 102578 1 0 60716
box -2638 -2806 3466 243
use a_mux4_en  a_mux4_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/a_mux4_en
timestamp 1654674840
transform 0 -1 62720 1 0 61957
box -3843 -5692 3675 352
use a_mux4_en  a_mux4_en_1
timestamp 1654674840
transform 0 -1 72720 1 0 61957
box -3843 -5692 3675 352
use clock_v2  clock_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/clock_v2
timestamp 1654674840
transform 0 -1 71097 1 0 -19032
box -3377 -14204 17044 36
use comparator_v2  comparator_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/comparator_v2
timestamp 1654674840
transform 0 1 115004 1 0 32246
box -3788 -193 7250 10729
use esd_cell  esd_cell_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/esd_cell
timestamp 1654674269
transform 0 -1 66871 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_1
timestamp 1654674269
transform 0 -1 76871 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_2
timestamp 1654674269
transform 0 -1 87821 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_3
timestamp 1654674269
transform 0 -1 105391 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_4
timestamp 1654674269
transform 0 -1 59771 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_5
timestamp 1654674269
transform 0 -1 96051 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_6
timestamp 1654674269
transform 0 -1 45351 1 0 67009
box -64 -64 3554 3096
use esd_cell  esd_cell_7
timestamp 1654674269
transform 0 -1 38351 1 0 67009
box -64 -64 3554 3096
use onebit_dac  onebit_dac_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/onebit_dac
timestamp 1654674269
transform 0 1 116581 1 0 50758
box -6 -1274 1554 1238
use onebit_dac  onebit_dac_1
timestamp 1654674269
transform 0 1 120581 1 0 50758
box -6 -1274 1554 1238
use ota_w_test_v2  ota_w_test_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/ota_w_test_v2
timestamp 1654674269
transform 0 1 56391 1 0 28511
box -170 1 23753 20628
use ota_w_test_v2  ota_w_test_v2_1
timestamp 1654674269
transform 0 1 90907 1 0 28504
box -170 1 23753 20628
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_0
timestamp 1654674269
transform 1 0 80428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_1
timestamp 1654674269
transform 1 0 82428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_2
timestamp 1654674269
transform 1 0 81428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_3
timestamp 1654674269
transform 1 0 83428 0 -1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_4
timestamp 1654674269
transform -1 0 87328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_5
timestamp 1654674269
transform -1 0 87328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_6
timestamp 1654674269
transform -1 0 86328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_7
timestamp 1654674269
transform -1 0 86328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_8
timestamp 1654674269
transform -1 0 85328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_9
timestamp 1654674269
transform 1 0 81428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_10
timestamp 1654674269
transform 1 0 82428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_11
timestamp 1654674269
transform 1 0 83428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_12
timestamp 1654674269
transform -1 0 85328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_13
timestamp 1654674269
transform -1 0 84328 0 1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_14
timestamp 1654674269
transform -1 0 84328 0 1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_15
timestamp 1654674269
transform 1 0 80428 0 -1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_16
timestamp 1654674269
transform 1 0 80428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_17
timestamp 1654674269
transform 1 0 81428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_18
timestamp 1654674269
transform 1 0 82428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_19
timestamp 1654674269
transform 1 0 83428 0 -1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_20
timestamp 1654674269
transform -1 0 87328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_21
timestamp 1654674269
transform -1 0 87328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_22
timestamp 1654674269
transform -1 0 86328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_23
timestamp 1654674269
transform -1 0 86328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_24
timestamp 1654674269
transform 1 0 80428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_25
timestamp 1654674269
transform 1 0 81428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_26
timestamp 1654674269
transform 1 0 82428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_27
timestamp 1654674269
transform 1 0 83428 0 -1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_28
timestamp 1654674269
transform -1 0 85328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_29
timestamp 1654674269
transform -1 0 85328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_30
timestamp 1654674269
transform -1 0 84328 0 1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_31
timestamp 1654674269
transform -1 0 84328 0 1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_32
timestamp 1654674269
transform 1 0 80428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_33
timestamp 1654674269
transform 1 0 81428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_34
timestamp 1654674269
transform 1 0 82428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_35
timestamp 1654674269
transform 1 0 83428 0 -1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_36
timestamp 1654674269
transform -1 0 87328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_37
timestamp 1654674269
transform -1 0 86328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_38
timestamp 1654674269
transform -1 0 85328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_39
timestamp 1654674269
transform -1 0 84328 0 1 32755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_40
timestamp 1654674269
transform 1 0 80428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_41
timestamp 1654674269
transform 1 0 81428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_42
timestamp 1654674269
transform 1 0 82428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_43
timestamp 1654674269
transform 1 0 83428 0 -1 31755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_44
timestamp 1654674269
transform -1 0 87328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_45
timestamp 1654674269
transform -1 0 87328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_46
timestamp 1654674269
transform -1 0 86328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_47
timestamp 1654674269
transform -1 0 86328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_48
timestamp 1654674269
transform 1 0 80428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_49
timestamp 1654674269
transform 1 0 81428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_50
timestamp 1654674269
transform 1 0 82428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_51
timestamp 1654674269
transform 1 0 83428 0 -1 30755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_52
timestamp 1654674269
transform -1 0 85328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_53
timestamp 1654674269
transform -1 0 85328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_54
timestamp 1654674269
transform -1 0 84328 0 1 33755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_55
timestamp 1654674269
transform -1 0 84328 0 1 34755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_56
timestamp 1654674269
transform 1 0 80428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_57
timestamp 1654674269
transform 1 0 81428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_58
timestamp 1654674269
transform 1 0 82428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_59
timestamp 1654674269
transform 1 0 83428 0 -1 29755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_60
timestamp 1654674269
transform -1 0 87328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_61
timestamp 1654674269
transform -1 0 87328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_62
timestamp 1654674269
transform -1 0 86328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_63
timestamp 1654674269
transform -1 0 86328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_64
timestamp 1654674269
transform 1 0 80428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_65
timestamp 1654674269
transform 1 0 81428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_66
timestamp 1654674269
transform 1 0 82428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_67
timestamp 1654674269
transform 1 0 83428 0 -1 28755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_68
timestamp 1654674269
transform -1 0 85328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_69
timestamp 1654674269
transform -1 0 85328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_70
timestamp 1654674269
transform -1 0 84328 0 1 35755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_71
timestamp 1654674269
transform -1 0 84328 0 1 36755
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_0
timestamp 1654674269
transform 0 -1 39165 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_1
timestamp 1654674269
transform 0 -1 39165 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_2
timestamp 1654674269
transform 0 -1 39165 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_3
timestamp 1654674269
transform 0 -1 39165 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_4
timestamp 1654674269
transform 0 -1 39165 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_5
timestamp 1654674269
transform 0 -1 39165 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_6
timestamp 1654674269
transform 0 -1 35965 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_7
timestamp 1654674269
transform 0 -1 35965 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_8
timestamp 1654674269
transform 0 -1 35965 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_9
timestamp 1654674269
transform 0 -1 35965 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_10
timestamp 1654674269
transform 0 -1 35965 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_11
timestamp 1654674269
transform 0 -1 35965 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_12
timestamp 1654674269
transform 0 -1 32765 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_13
timestamp 1654674269
transform 0 -1 32765 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_14
timestamp 1654674269
transform 0 -1 32765 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_15
timestamp 1654674269
transform 0 -1 32765 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_16
timestamp 1654674269
transform 0 -1 32765 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_17
timestamp 1654674269
transform 0 -1 32765 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_18
timestamp 1654674269
transform 0 -1 29565 1 0 29433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_19
timestamp 1654674269
transform 0 -1 29565 1 0 32633
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_20
timestamp 1654674269
transform 0 -1 29565 1 0 35833
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_21
timestamp 1654674269
transform 0 -1 29565 1 0 39033
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_22
timestamp 1654674269
transform 0 -1 29565 1 0 42233
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_23
timestamp 1654674269
transform 0 -1 29565 1 0 45433
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_24
timestamp 1654674269
transform 0 1 42365 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_25
timestamp 1654674269
transform 0 1 42365 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_26
timestamp 1654674269
transform 0 1 42365 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_27
timestamp 1654674269
transform 0 1 42365 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_28
timestamp 1654674269
transform 0 1 42365 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_29
timestamp 1654674269
transform 0 1 42365 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_30
timestamp 1654674269
transform 0 1 45565 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_31
timestamp 1654674269
transform 0 1 45565 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_32
timestamp 1654674269
transform 0 1 45565 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_33
timestamp 1654674269
transform 0 1 45565 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_34
timestamp 1654674269
transform 0 1 45565 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_35
timestamp 1654674269
transform 0 1 45565 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_36
timestamp 1654674269
transform 0 1 48765 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_37
timestamp 1654674269
transform 0 1 48765 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_38
timestamp 1654674269
transform 0 1 48765 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_39
timestamp 1654674269
transform 0 1 48765 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_40
timestamp 1654674269
transform 0 1 48765 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_41
timestamp 1654674269
transform 0 1 48765 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_42
timestamp 1654674269
transform 0 1 51965 -1 0 45331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_43
timestamp 1654674269
transform 0 1 51965 -1 0 42131
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_44
timestamp 1654674269
transform 0 1 51965 -1 0 38931
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_45
timestamp 1654674269
transform 0 1 51965 -1 0 35731
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_46
timestamp 1654674269
transform 0 1 51965 -1 0 32531
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_47
timestamp 1654674269
transform 0 1 51965 -1 0 29331
box -1031 -980 929 980
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_0
timestamp 1654674269
transform 0 1 110974 -1 0 30953
box -1310 -1260 1210 1260
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_1
timestamp 1654674269
transform 0 1 107306 -1 0 30955
box -1310 -1260 1210 1260
use sky130_fd_pr__nfet_01v8_CFEPS5  sky130_fd_pr__nfet_01v8_CFEPS5_0
timestamp 1654674269
transform 1 0 127406 0 -1 32821
box -311 -274 311 276
use sky130_fd_pr__pfet_01v8_hvt_XAYTAL  sky130_fd_pr__pfet_01v8_hvt_XAYTAL_0
timestamp 1654674269
transform 1 0 127406 0 -1 33415
box -311 -319 311 319
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 137539 0 1 11212
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1650294714
transform 1 0 137547 0 1 7951
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_2
timestamp 1650294714
transform 1 0 137547 0 1 4723
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_3
timestamp 1650294714
transform 1 0 137547 0 1 1356
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 -1 67137 1 0 -5429
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1650294714
transform 1 0 139471 0 1 11212
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_2
timestamp 1650294714
transform 1 0 139479 0 1 7951
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_3
timestamp 1650294714
transform 1 0 139479 0 1 4723
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_4
timestamp 1650294714
transform 1 0 139479 0 1 1356
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 -1 67137 1 0 -6625
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1650294714
transform 0 -1 67137 1 0 -3129
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_2
timestamp 1650294714
transform 1 0 136343 0 1 11212
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_3
timestamp 1650294714
transform 1 0 138275 0 1 11212
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_4
timestamp 1650294714
transform 1 0 141771 0 1 11212
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_5
timestamp 1650294714
transform 1 0 136351 0 1 7951
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_6
timestamp 1650294714
transform 1 0 138283 0 1 7951
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_7
timestamp 1650294714
transform 1 0 141779 0 1 7951
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_8
timestamp 1650294714
transform 1 0 136351 0 1 4723
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_9
timestamp 1650294714
transform 1 0 138283 0 1 4723
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_10
timestamp 1650294714
transform 1 0 141779 0 1 4723
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_11
timestamp 1650294714
transform 1 0 136351 0 1 1356
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_12
timestamp 1650294714
transform 1 0 138283 0 1 1356
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_13
timestamp 1650294714
transform 1 0 141779 0 1 1356
box -38 -48 1142 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 134411 0 1 11212
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_1
timestamp 1650294714
transform 1 0 134419 0 1 7951
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_2
timestamp 1650294714
transform 1 0 134419 0 1 4723
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_3
timestamp 1650294714
transform 1 0 134419 0 1 1356
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 -1 67137 1 0 -5521
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1650294714
transform 0 -1 67137 1 0 -3221
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1650294714
transform 1 0 134319 0 1 11212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1650294714
transform 1 0 137447 0 1 11212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1650294714
transform 1 0 138183 0 1 11212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1650294714
transform 1 0 139379 0 1 11212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1650294714
transform 1 0 141679 0 1 11212
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1650294714
transform 1 0 134327 0 1 7951
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1650294714
transform 1 0 137455 0 1 7951
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1650294714
transform 1 0 138191 0 1 7951
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1650294714
transform 1 0 139387 0 1 7951
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1650294714
transform 1 0 141687 0 1 7951
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1650294714
transform 1 0 134327 0 1 4723
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1650294714
transform 1 0 137455 0 1 4723
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1650294714
transform 1 0 138191 0 1 4723
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1650294714
transform 1 0 139387 0 1 4723
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1650294714
transform 1 0 141687 0 1 4723
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1650294714
transform 1 0 134327 0 1 1356
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1650294714
transform 1 0 137455 0 1 1356
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1650294714
transform 1 0 138191 0 1 1356
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1650294714
transform 1 0 139387 0 1 1356
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1650294714
transform 1 0 141687 0 1 1356
box -38 -48 130 592
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/transmission_gate
timestamp 1654674269
transform 1 0 53375 0 1 22637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_1
timestamp 1654674269
transform 1 0 50175 0 1 20637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_2
timestamp 1654674269
transform 1 0 50175 0 1 18637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_3
timestamp 1654674269
transform 1 0 53375 0 1 16637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_4
timestamp 1654674269
transform 1 0 43367 0 1 22642
box -53 -49 1241 1063
use transmission_gate  transmission_gate_5
timestamp 1654674269
transform 1 0 43367 0 1 16642
box -53 -49 1241 1063
use transmission_gate  transmission_gate_6
timestamp 1654674269
transform -1 0 47418 0 -1 21462
box -53 -49 1241 1063
use transmission_gate  transmission_gate_7
timestamp 1654674269
transform -1 0 47418 0 -1 19462
box -53 -49 1241 1063
use transmission_gate  transmission_gate_8
timestamp 1654674269
transform 1 0 39792 0 1 20644
box -53 -49 1241 1063
use transmission_gate  transmission_gate_9
timestamp 1654674269
transform 1 0 39792 0 1 18644
box -53 -49 1241 1063
use transmission_gate  transmission_gate_10
timestamp 1654674269
transform 0 1 36343 -1 0 50351
box -53 -49 1241 1063
use transmission_gate  transmission_gate_11
timestamp 1654674269
transform 0 1 38343 -1 0 50351
box -53 -49 1241 1063
use transmission_gate  transmission_gate_12
timestamp 1654674269
transform 1 0 60175 0 1 18637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_13
timestamp 1654674269
transform 1 0 62395 0 1 16637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_14
timestamp 1654674269
transform 1 0 62395 0 1 22637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_15
timestamp 1654674269
transform 1 0 60175 0 1 20637
box -53 -49 1241 1063
use transmission_gate  transmission_gate_16
timestamp 1654674269
transform 0 -1 68108 1 0 19681
box -53 -49 1241 1063
use transmission_gate  transmission_gate_17
timestamp 1654674269
transform 0 -1 85714 -1 0 43032
box -53 -49 1241 1063
use transmission_gate  transmission_gate_18
timestamp 1654674269
transform 0 -1 87714 -1 0 43032
box -53 -49 1241 1063
use transmission_gate  transmission_gate_19
timestamp 1654674269
transform 1 0 71459 0 1 22638
box -53 -49 1241 1063
use transmission_gate  transmission_gate_20
timestamp 1654674269
transform 1 0 71459 0 1 16648
box -53 -49 1241 1063
use transmission_gate  transmission_gate_21
timestamp 1654674269
transform 0 1 73976 1 0 19436
box -53 -49 1241 1063
use transmission_gate  transmission_gate_22
timestamp 1654674269
transform 1 0 85478 0 -1 16775
box -53 -49 1241 1063
use transmission_gate  transmission_gate_23
timestamp 1654674269
transform 1 0 82658 0 -1 17625
box -53 -49 1241 1063
use transmission_gate  transmission_gate_24
timestamp 1654674269
transform 1 0 82658 0 -1 23595
box -53 -49 1241 1063
use transmission_gate  transmission_gate_25
timestamp 1654674269
transform 1 0 85478 0 -1 24785
box -53 -49 1241 1063
use transmission_gate  transmission_gate_26
timestamp 1654674269
transform -1 0 90507 0 -1 23595
box -53 -49 1241 1063
use transmission_gate  transmission_gate_27
timestamp 1654674269
transform -1 0 90507 0 -1 17625
box -53 -49 1241 1063
use transmission_gate  transmission_gate_28
timestamp 1654674269
transform -1 0 109760 0 1 27857
box -53 -49 1241 1063
use transmission_gate  transmission_gate_29
timestamp 1654674269
transform 0 -1 83121 -1 0 41228
box -53 -49 1241 1063
use transmission_gate  transmission_gate_30
timestamp 1654674269
transform 0 -1 81121 -1 0 41228
box -53 -49 1241 1063
use transmission_gate  transmission_gate_31
timestamp 1654674269
transform 0 1 48389 -1 0 52358
box -53 -49 1241 1063
use transmission_gate  transmission_gate_32
timestamp 1654674269
transform 0 1 46389 -1 0 52348
box -53 -49 1241 1063
<< end >>
