magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< metal3 >>
rect -360 -310 260 310
<< mimcap >>
rect -260 152 160 210
rect -260 -152 -202 152
rect 102 -152 160 152
rect -260 -210 160 -152
<< mimcapcontact >>
rect -202 -152 102 152
<< metal4 >>
rect -221 152 121 171
rect -221 -152 -202 152
rect 102 -152 121 152
rect -221 -171 121 -152
<< properties >>
string FIXED_BBOX -360 -310 260 310
<< end >>
