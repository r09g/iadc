magic
tech sky130A
timestamp 1654894986
<< end >>
