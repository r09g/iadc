magic
tech sky130A
magscale 1 2
timestamp 1654526415
<< nwell >>
rect -1129 -2208 -869 -2205
rect -599 -2208 -428 -2205
rect -592 -2332 -540 -2280
rect -434 -2290 -428 -2208
<< pwell >>
rect -934 -525 -635 -498
rect -934 -680 -384 -525
rect -701 -1768 -384 -1362
rect -1253 -2605 -337 -2450
rect -1241 -2632 -337 -2605
rect -1253 -2856 -340 -2701
rect -701 -3693 -337 -3538
rect -702 -3944 -338 -3789
rect -701 -4781 -337 -4626
<< locali >>
rect -3843 224 3659 352
rect -1670 -118 -1542 224
rect -2022 -182 -1542 -118
rect -1670 -989 -1542 -182
rect -165 -133 1647 -5
rect -165 -444 -37 -133
rect -355 -508 -37 -444
rect -3564 -1088 -3222 -1024
rect -1670 -1053 -891 -989
rect -3564 -2383 -3500 -1088
rect -1670 -1443 -1542 -1053
rect -165 -1334 -37 -508
rect 3329 -1069 3457 224
rect 3042 -1121 3457 -1069
rect 1677 -1249 3457 -1121
rect -2030 -1507 -1542 -1443
rect -1670 -2082 -1542 -1507
rect -165 -1462 1650 -1334
rect -165 -1503 327 -1462
rect -165 -1548 -37 -1503
rect -358 -1581 -37 -1548
rect -345 -1582 -37 -1581
rect -1670 -2146 -1220 -2082
rect -3564 -2447 -3210 -2383
rect -3564 -3782 -3500 -2447
rect -1670 -2841 -1542 -2146
rect -592 -2332 -540 -2280
rect -165 -2636 -37 -1582
rect 3329 -2396 3457 -1249
rect 3042 -2447 3457 -2396
rect 1686 -2575 3457 -2447
rect -343 -2670 -37 -2636
rect -2031 -2905 -1542 -2841
rect -165 -2713 -37 -2670
rect -165 -2841 1647 -2713
rect -1670 -3164 -1542 -2905
rect -165 -2882 340 -2841
rect -1670 -3228 -1203 -3164
rect -3564 -3846 -3211 -3782
rect -3564 -5168 -3500 -3846
rect -1670 -4239 -1542 -3228
rect -165 -3724 -37 -2882
rect -349 -3758 -37 -3724
rect -165 -4083 -37 -3758
rect 3329 -3779 3457 -2575
rect 3039 -3831 3457 -3779
rect 1686 -3959 3457 -3831
rect -2023 -4258 -1542 -4239
rect -165 -4211 1661 -4083
rect -2023 -4303 -649 -4258
rect -1670 -4322 -649 -4303
rect -165 -4264 340 -4211
rect -1670 -4324 -1542 -4322
rect -165 -4812 -37 -4264
rect -348 -4846 -37 -4812
rect -3564 -5232 -3216 -5168
rect -3564 -5564 -3500 -5232
rect -165 -5564 -37 -4846
rect 3329 -5227 3457 -3959
rect 1661 -5355 3457 -5227
rect -3827 -5692 3675 -5564
<< viali >>
rect -822 -637 -788 -603
rect -452 -628 -418 -594
rect -905 -732 -871 -698
rect -538 -734 -504 -700
rect -453 -1231 -419 -1197
rect -534 -1346 -500 -1312
rect -469 -1710 -435 -1676
rect -582 -1818 -548 -1784
rect -408 -1819 -374 -1785
rect -1004 -2270 -970 -2236
rect -489 -2304 -455 -2270
rect -1091 -2432 -1057 -2398
rect -583 -2432 -549 -2398
rect -402 -2429 -368 -2395
rect -1089 -2908 -1055 -2874
rect -994 -2908 -960 -2874
rect -574 -2908 -540 -2874
rect -401 -2909 -367 -2875
rect -490 -3070 -456 -3036
rect -576 -3526 -542 -3492
rect -405 -3521 -371 -3487
rect -492 -3624 -458 -3590
rect -539 -3995 -505 -3961
rect -453 -4154 -419 -4120
rect -452 -4452 -418 -4418
rect -540 -4608 -506 -4574
<< metal1 >>
rect -1597 -121 -1587 -69
rect -1535 -121 -914 -69
rect -862 -121 -852 -69
rect -1952 -246 -1942 -194
rect -1890 -246 -1416 -194
rect -1364 -246 -1354 -194
rect -80 -547 124 -513
rect -1426 -645 -1416 -593
rect -1364 -597 -1354 -593
rect -1364 -603 -776 -597
rect -1364 -637 -822 -603
rect -788 -637 -776 -603
rect -471 -636 -461 -584
rect -409 -636 -399 -584
rect -1364 -643 -776 -637
rect -1364 -645 -1354 -643
rect -3461 -742 -3272 -690
rect -1984 -733 -1797 -699
rect -1831 -870 -1797 -733
rect -924 -742 -914 -690
rect -862 -742 -852 -690
rect -559 -746 -549 -694
rect -497 -746 -487 -694
rect -80 -870 -46 -547
rect 3080 -556 3317 -504
rect -1831 -904 -46 -870
rect 88 -1191 98 -1188
rect -465 -1197 98 -1191
rect -465 -1231 -453 -1197
rect -419 -1231 98 -1197
rect -465 -1237 98 -1231
rect 88 -1240 98 -1237
rect 150 -1240 160 -1188
rect -549 -1312 -287 -1303
rect -549 -1346 -534 -1312
rect -500 -1346 -287 -1312
rect -549 -1355 -287 -1346
rect -235 -1355 -225 -1303
rect -1852 -1446 -50 -1412
rect -3461 -2075 -3274 -2023
rect -1852 -2033 -1818 -1446
rect -1734 -1580 -1724 -1528
rect -1672 -1580 -1416 -1528
rect -1364 -1580 -1354 -1528
rect -488 -1721 -478 -1669
rect -426 -1721 -416 -1669
rect -602 -1828 -592 -1776
rect -540 -1828 -530 -1776
rect -426 -1831 -416 -1779
rect -364 -1831 -354 -1779
rect -84 -1847 -50 -1446
rect 3265 -1839 3317 -556
rect -84 -1881 122 -1847
rect 3075 -1891 3317 -1839
rect -882 -1971 -872 -1919
rect -820 -1971 -416 -1919
rect -364 -1971 -354 -1919
rect -1976 -2067 -1818 -2033
rect -602 -2230 -592 -2225
rect -1016 -2236 -592 -2230
rect -1016 -2270 -1004 -2236
rect -970 -2270 -592 -2236
rect -1016 -2276 -592 -2270
rect -602 -2277 -592 -2276
rect -540 -2277 -530 -2225
rect -297 -2264 -287 -2261
rect -501 -2270 -287 -2264
rect -501 -2304 -489 -2270
rect -455 -2304 -287 -2270
rect -501 -2310 -287 -2304
rect -297 -2313 -287 -2310
rect -235 -2313 -225 -2261
rect -1111 -2440 -1101 -2388
rect -1049 -2440 -762 -2388
rect -710 -2440 -700 -2388
rect -602 -2442 -592 -2390
rect -540 -2442 -530 -2390
rect -422 -2437 -412 -2385
rect -360 -2437 -350 -2385
rect 87 -2386 179 -2334
rect -1250 -2543 -1240 -2491
rect -1188 -2543 -412 -2491
rect -360 -2543 -350 -2491
rect 3265 -2617 3317 -1891
rect 3265 -2626 3454 -2617
rect 3265 -2660 3456 -2626
rect 3265 -2669 3454 -2660
rect -772 -2827 -762 -2775
rect -710 -2827 -412 -2775
rect -360 -2827 -350 -2775
rect -1936 -2958 -1926 -2906
rect -1874 -2958 -1416 -2906
rect -1364 -2958 -1354 -2906
rect -1108 -2917 -1098 -2865
rect -1046 -2917 -1036 -2865
rect -1002 -2868 -872 -2864
rect -1006 -2874 -872 -2868
rect -1006 -2908 -994 -2874
rect -960 -2908 -872 -2874
rect -1006 -2914 -872 -2908
rect -1002 -2916 -872 -2914
rect -820 -2874 -527 -2864
rect -820 -2908 -574 -2874
rect -540 -2908 -527 -2874
rect -820 -2916 -527 -2908
rect -1002 -2918 -527 -2916
rect -422 -2918 -412 -2866
rect -360 -2918 -350 -2866
rect -246 -3030 -236 -3026
rect -502 -3036 -236 -3030
rect -502 -3070 -490 -3036
rect -456 -3070 -236 -3036
rect -502 -3076 -236 -3070
rect -246 -3078 -236 -3076
rect -184 -3078 -174 -3026
rect 3265 -3216 3317 -2669
rect -44 -3259 140 -3225
rect -44 -3308 -10 -3259
rect 3077 -3268 3317 -3216
rect -1812 -3342 -10 -3308
rect -3461 -3455 -3271 -3403
rect -1812 -3411 -1778 -3342
rect -1982 -3445 -1778 -3411
rect -773 -3445 -762 -3393
rect -710 -3445 -414 -3393
rect -362 -3445 -352 -3393
rect -1251 -3539 -1241 -3485
rect -1187 -3492 -528 -3485
rect -1187 -3526 -576 -3492
rect -542 -3526 -528 -3492
rect -424 -3526 -414 -3474
rect -362 -3526 -352 -3474
rect -1187 -3539 -528 -3526
rect -417 -3527 -359 -3526
rect -510 -3632 -500 -3580
rect -448 -3632 -438 -3580
rect -245 -3764 -235 -3712
rect -183 -3764 122 -3712
rect -579 -3961 -236 -3951
rect -579 -3995 -539 -3961
rect -505 -3995 -236 -3961
rect -579 -4003 -236 -3995
rect -184 -4003 -173 -3951
rect -91 -4114 -81 -4111
rect -465 -4120 -81 -4114
rect -465 -4154 -453 -4120
rect -419 -4154 -81 -4120
rect -465 -4160 -81 -4154
rect -91 -4163 -81 -4160
rect -29 -4163 -19 -4111
rect -1953 -4336 -1943 -4284
rect -1891 -4336 -1416 -4284
rect -1364 -4336 -1354 -4284
rect 82 -4412 92 -4409
rect -464 -4418 92 -4412
rect -464 -4452 -452 -4418
rect -418 -4452 92 -4418
rect -464 -4458 92 -4452
rect 82 -4461 92 -4458
rect 144 -4461 154 -4409
rect -558 -4617 -548 -4565
rect -496 -4617 -486 -4565
rect 3265 -4595 3317 -3268
rect -48 -4637 104 -4603
rect -48 -4674 -14 -4637
rect 3075 -4647 3317 -4595
rect -1808 -4708 -14 -4674
rect -3461 -4832 -3278 -4780
rect -1808 -4789 -1774 -4708
rect -1975 -4823 -1774 -4789
<< via1 >>
rect -1587 -121 -1535 -69
rect -914 -121 -862 -69
rect -1942 -246 -1890 -194
rect -1416 -246 -1364 -194
rect -1416 -645 -1364 -593
rect -461 -594 -409 -584
rect -461 -628 -452 -594
rect -452 -628 -418 -594
rect -418 -628 -409 -594
rect -461 -636 -409 -628
rect -914 -698 -862 -690
rect -914 -732 -905 -698
rect -905 -732 -871 -698
rect -871 -732 -862 -698
rect -914 -742 -862 -732
rect -549 -700 -497 -694
rect -549 -734 -538 -700
rect -538 -734 -504 -700
rect -504 -734 -497 -700
rect -549 -746 -497 -734
rect 98 -1240 150 -1188
rect -287 -1355 -235 -1303
rect -1724 -1580 -1672 -1528
rect -1416 -1580 -1364 -1528
rect -478 -1676 -426 -1669
rect -478 -1710 -469 -1676
rect -469 -1710 -435 -1676
rect -435 -1710 -426 -1676
rect -478 -1721 -426 -1710
rect -592 -1784 -540 -1776
rect -592 -1818 -582 -1784
rect -582 -1818 -548 -1784
rect -548 -1818 -540 -1784
rect -592 -1828 -540 -1818
rect -416 -1785 -364 -1779
rect -416 -1819 -408 -1785
rect -408 -1819 -374 -1785
rect -374 -1819 -364 -1785
rect -416 -1831 -364 -1819
rect -872 -1971 -820 -1919
rect -416 -1971 -364 -1919
rect -592 -2277 -540 -2225
rect -287 -2313 -235 -2261
rect -1101 -2398 -1049 -2388
rect -1101 -2432 -1091 -2398
rect -1091 -2432 -1057 -2398
rect -1057 -2432 -1049 -2398
rect -1101 -2440 -1049 -2432
rect -762 -2440 -710 -2388
rect -592 -2398 -540 -2390
rect -592 -2432 -583 -2398
rect -583 -2432 -549 -2398
rect -549 -2432 -540 -2398
rect -592 -2442 -540 -2432
rect -412 -2395 -360 -2385
rect -412 -2429 -402 -2395
rect -402 -2429 -368 -2395
rect -368 -2429 -360 -2395
rect -412 -2437 -360 -2429
rect -1240 -2543 -1188 -2491
rect -412 -2543 -360 -2491
rect -762 -2827 -710 -2775
rect -412 -2827 -360 -2775
rect -1926 -2958 -1874 -2906
rect -1416 -2958 -1364 -2906
rect -1098 -2874 -1046 -2865
rect -1098 -2908 -1089 -2874
rect -1089 -2908 -1055 -2874
rect -1055 -2908 -1046 -2874
rect -1098 -2917 -1046 -2908
rect -872 -2916 -820 -2864
rect -412 -2875 -360 -2866
rect -412 -2909 -401 -2875
rect -401 -2909 -367 -2875
rect -367 -2909 -360 -2875
rect -412 -2918 -360 -2909
rect -236 -3078 -184 -3026
rect -762 -3445 -710 -3393
rect -414 -3445 -362 -3393
rect -1241 -3539 -1187 -3485
rect -414 -3487 -362 -3474
rect -414 -3521 -405 -3487
rect -405 -3521 -371 -3487
rect -371 -3521 -362 -3487
rect -414 -3526 -362 -3521
rect -500 -3590 -448 -3580
rect -500 -3624 -492 -3590
rect -492 -3624 -458 -3590
rect -458 -3624 -448 -3590
rect -500 -3632 -448 -3624
rect -235 -3764 -183 -3712
rect -236 -4003 -184 -3951
rect -81 -4163 -29 -4111
rect -1943 -4336 -1891 -4284
rect -1416 -4336 -1364 -4284
rect 92 -4461 144 -4409
rect -548 -4574 -496 -4565
rect -548 -4608 -540 -4574
rect -540 -4608 -506 -4574
rect -506 -4608 -496 -4574
rect -548 -4617 -496 -4608
<< metal2 >>
rect -1587 -69 -1535 148
rect -1942 -194 -1890 -184
rect -2217 -246 -1942 -194
rect -1942 -256 -1890 -246
rect -1587 -1001 -1535 -121
rect -2241 -1053 -1535 -1001
rect -1724 -1528 -1672 -1518
rect -2238 -1580 -1724 -1528
rect -1724 -1590 -1672 -1580
rect -1587 -2335 -1535 -1053
rect -2224 -2387 -1535 -2335
rect -1926 -2906 -1874 -2896
rect -2222 -2958 -1926 -2906
rect -1926 -2968 -1874 -2958
rect -1587 -3713 -1535 -2387
rect -1416 -194 -1364 -184
rect -1416 -593 -1364 -246
rect -1416 -1528 -1364 -645
rect -1416 -2906 -1364 -1580
rect -2217 -3765 -1532 -3713
rect -1943 -4284 -1891 -4274
rect -2222 -4336 -1943 -4284
rect -1943 -4346 -1891 -4336
rect -1587 -5091 -1535 -3765
rect -1416 -4284 -1364 -2958
rect -1241 -2491 -1187 148
rect -1101 -2388 -1049 148
rect -914 -69 -862 -60
rect -914 -690 -862 -121
rect -461 -245 227 -193
rect -461 -584 -409 -245
rect -461 -646 -409 -636
rect -914 -752 -862 -742
rect -549 -694 -497 -684
rect -497 -746 -426 -694
rect -549 -756 -426 -746
rect -478 -1000 -426 -756
rect -478 -1052 255 -1000
rect -478 -1669 -426 -1052
rect 98 -1188 150 -1178
rect -478 -1731 -426 -1721
rect -287 -1303 -235 -1293
rect -592 -1776 -540 -1766
rect -1101 -2450 -1049 -2440
rect -872 -1919 -820 -1909
rect -1241 -2543 -1240 -2491
rect -1188 -2543 -1187 -2491
rect -1241 -2864 -1187 -2543
rect -1098 -2864 -1046 -2855
rect -872 -2864 -820 -1971
rect -592 -2225 -540 -1828
rect -416 -1779 -364 -1769
rect -416 -1919 -364 -1831
rect -416 -1981 -364 -1971
rect -1241 -2865 -1045 -2864
rect -1241 -2917 -1098 -2865
rect -1046 -2917 -1045 -2865
rect -1241 -2918 -1045 -2917
rect -1241 -3485 -1187 -2918
rect -1098 -2927 -1046 -2918
rect -872 -2926 -820 -2916
rect -762 -2388 -710 -2378
rect -762 -2775 -710 -2440
rect -592 -2390 -540 -2277
rect -287 -2261 -235 -1355
rect 98 -1589 150 -1240
rect -235 -2313 148 -2261
rect -287 -2323 -235 -2313
rect 96 -2324 148 -2313
rect 96 -2334 201 -2324
rect -592 -2450 -540 -2442
rect -412 -2385 -360 -2375
rect 96 -2386 253 -2334
rect 96 -2389 196 -2386
rect 96 -2397 201 -2389
rect -412 -2491 -360 -2437
rect -412 -2553 -360 -2543
rect -762 -3393 -710 -2827
rect -412 -2775 -360 -2765
rect -412 -2866 -360 -2827
rect -412 -2928 -360 -2918
rect -81 -2957 201 -2905
rect -236 -3026 -184 -3016
rect -762 -3475 -710 -3445
rect -414 -3393 -362 -3383
rect -414 -3474 -362 -3445
rect -414 -3536 -362 -3526
rect -1241 -3549 -1187 -3539
rect -1416 -4346 -1364 -4336
rect -500 -3580 -448 -3570
rect -500 -4555 -448 -3632
rect -236 -3702 -184 -3078
rect -236 -3712 -183 -3702
rect -236 -3764 -235 -3712
rect -236 -3774 -183 -3764
rect -236 -3951 -184 -3774
rect -236 -4013 -184 -4003
rect -81 -4111 -29 -2957
rect -81 -4173 -29 -4163
rect 92 -4325 189 -4273
rect 92 -4345 164 -4325
rect 92 -4409 144 -4345
rect 92 -4471 144 -4461
rect -548 -4565 -448 -4555
rect -496 -4617 -448 -4565
rect -548 -4627 -448 -4617
rect -2223 -5143 -1535 -5091
rect -500 -5089 -448 -4627
rect -500 -5141 203 -5089
rect -1587 -5148 -1535 -5143
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform -1 0 -704 0 -1 -2653
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_1
timestamp 1650294714
transform 1 0 -888 0 1 -2653
box -38 -48 222 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654309566
transform 1 0 -1164 0 -1 -2653
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1654309566
transform 1 0 -1164 0 1 -2653
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1654309566
transform 1 0 -612 0 1 -1565
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1654309566
transform 1 0 -612 0 -1 -477
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1654309566
transform 1 0 -612 0 -1 -3741
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1654309566
transform 1 0 -612 0 1 -4829
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1654309566
transform 1 0 -980 0 -1 -477
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 -612 0 1 -3741
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1650294714
transform 1 0 -612 0 -1 -2653
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2
timestamp 1650294714
transform 1 0 -612 0 1 -2653
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_3
timestamp 1650294714
transform 1 0 -612 0 -1 -1565
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform -1 0 -1164 0 -1 -2653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1650294714
transform 1 0 -1256 0 1 -2653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1650294714
transform -1 0 -612 0 -1 -1565
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1650294714
transform 1 0 -704 0 1 -3741
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1650294714
transform 1 0 -704 0 1 -1565
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1650294714
transform -1 0 -612 0 -1 -477
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1650294714
transform -1 0 -612 0 -1 -3741
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1650294714
transform 1 0 -704 0 1 -4829
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1650294714
transform -1 0 -612 0 -1 -2653
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1650294714
transform 1 0 -704 0 1 -2653
box -38 -48 130 592
use switch_5t  switch_5t_0
timestamp 1654526415
transform 1 0 123 0 -1 -62
box -53 4 3056 1118
use switch_5t  switch_5t_1
timestamp 1654526415
transform 1 0 123 0 -1 -1396
box -53 4 3056 1118
use switch_5t  switch_5t_2
timestamp 1654526415
transform 1 0 123 0 -1 -2774
box -53 4 3056 1118
use switch_5t  switch_5t_3
timestamp 1654526415
transform 1 0 123 0 -1 -4152
box -53 4 3056 1118
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/transmission_gate
timestamp 1654522530
transform 1 0 -3213 0 1 -1129
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1654522530
transform 1 0 -3213 0 1 -2463
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1654522530
transform 1 0 -3213 0 1 -3841
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1654522530
transform 1 0 -3213 0 1 -5219
box -216 -51 1283 1063
<< labels >>
flabel metal1 3438 -2641 3438 -2641 1 FreeSans 400 0 0 0 out
flabel metal2 -1562 128 -1562 128 1 FreeSans 400 0 0 0 en
flabel metal2 -1216 128 -1216 128 1 FreeSans 400 0 0 0 s1
flabel metal2 -1073 128 -1073 128 1 FreeSans 400 0 0 0 s0
flabel metal1 -3454 -717 -3454 -717 1 FreeSans 400 0 0 0 in0
flabel metal1 -3454 -2051 -3454 -2051 1 FreeSans 400 0 0 0 in1
flabel metal1 -3455 -3430 -3455 -3430 1 FreeSans 400 0 0 0 in2
flabel metal1 -3453 -4807 -3453 -4807 1 FreeSans 400 0 0 0 in3
flabel locali -3783 -5630 -3783 -5630 1 FreeSans 400 0 0 0 VSS
flabel locali -3801 286 -3801 286 1 FreeSans 400 0 0 0 VDD
<< end >>
