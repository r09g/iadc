magic
tech sky130A
magscale 1 2
timestamp 1654717932
<< nwell >>
rect 7153 18323 8447 18973
rect 20083 18323 21377 18973
rect 7153 16523 8447 17173
rect 20083 16523 21377 17173
rect 7153 14723 8447 15373
rect 20083 14723 21377 15373
rect 7153 12923 8447 13573
rect 20083 12923 21377 13573
rect 7153 11123 8447 11773
rect 20083 11123 21377 11773
rect 7153 9323 8447 9973
rect 20083 9323 21377 9973
rect 14291 7047 21042 7048
rect 7215 5341 21042 7047
rect 7215 4020 13093 5341
<< pwell >>
rect 7153 17861 8447 18323
rect 20083 17861 21377 18323
rect 7153 16061 8447 16523
rect 20083 16061 21377 16523
rect 7153 14261 8447 14723
rect 20083 14261 21377 14723
rect 7153 12461 8447 12923
rect 20083 12461 21377 12923
rect 7153 10661 8447 11123
rect 20083 10661 21377 11123
rect 7153 8861 8447 9323
rect 20083 8861 21377 9323
rect -116 3990 7122 4864
rect 13288 3990 22069 5305
rect -116 3 22069 3990
rect 13288 1 22069 3
<< nmos >>
rect 7353 18071 7383 18175
rect 7449 18071 7479 18175
rect 7545 18071 7575 18175
rect 7641 18071 7671 18175
rect 7737 18071 7767 18175
rect 7833 18071 7863 18175
rect 7929 18071 7959 18175
rect 8025 18071 8055 18175
rect 8121 18071 8151 18175
rect 8217 18071 8247 18175
rect 20283 18071 20313 18175
rect 20379 18071 20409 18175
rect 20475 18071 20505 18175
rect 20571 18071 20601 18175
rect 20667 18071 20697 18175
rect 20763 18071 20793 18175
rect 20859 18071 20889 18175
rect 20955 18071 20985 18175
rect 21051 18071 21081 18175
rect 21147 18071 21177 18175
rect 7353 16271 7383 16375
rect 7449 16271 7479 16375
rect 7545 16271 7575 16375
rect 7641 16271 7671 16375
rect 7737 16271 7767 16375
rect 7833 16271 7863 16375
rect 7929 16271 7959 16375
rect 8025 16271 8055 16375
rect 8121 16271 8151 16375
rect 8217 16271 8247 16375
rect 20283 16271 20313 16375
rect 20379 16271 20409 16375
rect 20475 16271 20505 16375
rect 20571 16271 20601 16375
rect 20667 16271 20697 16375
rect 20763 16271 20793 16375
rect 20859 16271 20889 16375
rect 20955 16271 20985 16375
rect 21051 16271 21081 16375
rect 21147 16271 21177 16375
rect 7353 14471 7383 14575
rect 7449 14471 7479 14575
rect 7545 14471 7575 14575
rect 7641 14471 7671 14575
rect 7737 14471 7767 14575
rect 7833 14471 7863 14575
rect 7929 14471 7959 14575
rect 8025 14471 8055 14575
rect 8121 14471 8151 14575
rect 8217 14471 8247 14575
rect 20283 14471 20313 14575
rect 20379 14471 20409 14575
rect 20475 14471 20505 14575
rect 20571 14471 20601 14575
rect 20667 14471 20697 14575
rect 20763 14471 20793 14575
rect 20859 14471 20889 14575
rect 20955 14471 20985 14575
rect 21051 14471 21081 14575
rect 21147 14471 21177 14575
rect 7353 12671 7383 12775
rect 7449 12671 7479 12775
rect 7545 12671 7575 12775
rect 7641 12671 7671 12775
rect 7737 12671 7767 12775
rect 7833 12671 7863 12775
rect 7929 12671 7959 12775
rect 8025 12671 8055 12775
rect 8121 12671 8151 12775
rect 8217 12671 8247 12775
rect 20283 12671 20313 12775
rect 20379 12671 20409 12775
rect 20475 12671 20505 12775
rect 20571 12671 20601 12775
rect 20667 12671 20697 12775
rect 20763 12671 20793 12775
rect 20859 12671 20889 12775
rect 20955 12671 20985 12775
rect 21051 12671 21081 12775
rect 21147 12671 21177 12775
rect 7353 10871 7383 10975
rect 7449 10871 7479 10975
rect 7545 10871 7575 10975
rect 7641 10871 7671 10975
rect 7737 10871 7767 10975
rect 7833 10871 7863 10975
rect 7929 10871 7959 10975
rect 8025 10871 8055 10975
rect 8121 10871 8151 10975
rect 8217 10871 8247 10975
rect 20283 10871 20313 10975
rect 20379 10871 20409 10975
rect 20475 10871 20505 10975
rect 20571 10871 20601 10975
rect 20667 10871 20697 10975
rect 20763 10871 20793 10975
rect 20859 10871 20889 10975
rect 20955 10871 20985 10975
rect 21051 10871 21081 10975
rect 21147 10871 21177 10975
rect 7353 9071 7383 9175
rect 7449 9071 7479 9175
rect 7545 9071 7575 9175
rect 7641 9071 7671 9175
rect 7737 9071 7767 9175
rect 7833 9071 7863 9175
rect 7929 9071 7959 9175
rect 8025 9071 8055 9175
rect 8121 9071 8151 9175
rect 8217 9071 8247 9175
rect 20283 9071 20313 9175
rect 20379 9071 20409 9175
rect 20475 9071 20505 9175
rect 20571 9071 20601 9175
rect 20667 9071 20697 9175
rect 20763 9071 20793 9175
rect 20859 9071 20889 9175
rect 20955 9071 20985 9175
rect 21051 9071 21081 9175
rect 21147 9071 21177 9175
rect 474 3171 594 3451
rect 652 3171 772 3451
rect 830 3171 950 3451
rect 1008 3171 1128 3451
rect 1186 3171 1306 3451
rect 1364 3171 1484 3451
rect 1542 3171 1662 3451
rect 1720 3171 1840 3451
rect 1898 3171 2018 3451
rect 2076 3171 2196 3451
rect 2254 3171 2374 3451
rect 2432 3171 2552 3451
rect 2610 3171 2730 3451
rect 2788 3171 2908 3451
rect 2966 3171 3086 3451
rect 3144 3171 3264 3451
rect 3322 3171 3442 3451
rect 3500 3171 3620 3451
rect 3874 3171 3994 3451
rect 4052 3171 4172 3451
rect 4230 3171 4350 3451
rect 4408 3171 4528 3451
rect 4586 3171 4706 3451
rect 4764 3171 4884 3451
rect 4942 3171 5062 3451
rect 5120 3171 5240 3451
rect 5298 3171 5418 3451
rect 5476 3171 5596 3451
rect 5654 3171 5774 3451
rect 5832 3171 5952 3451
rect 6010 3171 6130 3451
rect 6188 3171 6308 3451
rect 6366 3171 6486 3451
rect 6544 3171 6664 3451
rect 6722 3171 6842 3451
rect 6900 3171 7020 3451
rect 7603 3371 7723 3651
rect 7781 3371 7901 3651
rect 7959 3371 8079 3651
rect 8137 3371 8257 3651
rect 8315 3371 8435 3651
rect 8493 3371 8613 3651
rect 8671 3371 8791 3651
rect 8849 3371 8969 3651
rect 9027 3371 9147 3651
rect 9205 3371 9325 3651
rect 9383 3371 9503 3651
rect 9561 3371 9681 3651
rect 9739 3371 9859 3651
rect 9917 3371 10037 3651
rect 10290 3371 10410 3651
rect 10468 3371 10588 3651
rect 10646 3371 10766 3651
rect 10824 3371 10944 3651
rect 11002 3371 11122 3651
rect 11180 3371 11300 3651
rect 11358 3371 11478 3651
rect 11536 3371 11656 3651
rect 11714 3371 11834 3651
rect 11892 3371 12012 3651
rect 12070 3371 12190 3651
rect 12248 3371 12368 3651
rect 12426 3371 12546 3651
rect 12604 3371 12724 3651
rect 474 2671 594 2951
rect 652 2671 772 2951
rect 830 2671 950 2951
rect 1008 2671 1128 2951
rect 1186 2671 1306 2951
rect 1364 2671 1484 2951
rect 1542 2671 1662 2951
rect 1720 2671 1840 2951
rect 1898 2671 2018 2951
rect 2076 2671 2196 2951
rect 2254 2671 2374 2951
rect 2432 2671 2552 2951
rect 2610 2671 2730 2951
rect 2788 2671 2908 2951
rect 2966 2671 3086 2951
rect 3144 2671 3264 2951
rect 3322 2671 3442 2951
rect 3500 2671 3620 2951
rect 3874 2671 3994 2951
rect 4052 2671 4172 2951
rect 4230 2671 4350 2951
rect 4408 2671 4528 2951
rect 4586 2671 4706 2951
rect 4764 2671 4884 2951
rect 4942 2671 5062 2951
rect 5120 2671 5240 2951
rect 5298 2671 5418 2951
rect 5476 2671 5596 2951
rect 5654 2671 5774 2951
rect 5832 2671 5952 2951
rect 6010 2671 6130 2951
rect 6188 2671 6308 2951
rect 6366 2671 6486 2951
rect 6544 2671 6664 2951
rect 6722 2671 6842 2951
rect 6900 2671 7020 2951
rect 7603 2871 7723 3151
rect 7781 2871 7901 3151
rect 7959 2871 8079 3151
rect 8137 2871 8257 3151
rect 8315 2871 8435 3151
rect 8493 2871 8613 3151
rect 8671 2871 8791 3151
rect 8849 2871 8969 3151
rect 9027 2871 9147 3151
rect 9205 2871 9325 3151
rect 9383 2871 9503 3151
rect 9561 2871 9681 3151
rect 9739 2871 9859 3151
rect 9917 2871 10037 3151
rect 10290 2871 10410 3151
rect 10468 2871 10588 3151
rect 10646 2871 10766 3151
rect 10824 2871 10944 3151
rect 11002 2871 11122 3151
rect 11180 2871 11300 3151
rect 11358 2871 11478 3151
rect 11536 2871 11656 3151
rect 11714 2871 11834 3151
rect 11892 2871 12012 3151
rect 12070 2871 12190 3151
rect 12248 2871 12368 3151
rect 12426 2871 12546 3151
rect 12604 2871 12724 3151
rect 474 2171 594 2451
rect 652 2171 772 2451
rect 830 2171 950 2451
rect 1008 2171 1128 2451
rect 1186 2171 1306 2451
rect 1364 2171 1484 2451
rect 1542 2171 1662 2451
rect 1720 2171 1840 2451
rect 1898 2171 2018 2451
rect 2076 2171 2196 2451
rect 2254 2171 2374 2451
rect 2432 2171 2552 2451
rect 2610 2171 2730 2451
rect 2788 2171 2908 2451
rect 2966 2171 3086 2451
rect 3144 2171 3264 2451
rect 3322 2171 3442 2451
rect 3500 2171 3620 2451
rect 3874 2171 3994 2451
rect 4052 2171 4172 2451
rect 4230 2171 4350 2451
rect 4408 2171 4528 2451
rect 4586 2171 4706 2451
rect 4764 2171 4884 2451
rect 4942 2171 5062 2451
rect 5120 2171 5240 2451
rect 5298 2171 5418 2451
rect 5476 2171 5596 2451
rect 5654 2171 5774 2451
rect 5832 2171 5952 2451
rect 6010 2171 6130 2451
rect 6188 2171 6308 2451
rect 6366 2171 6486 2451
rect 6544 2171 6664 2451
rect 6722 2171 6842 2451
rect 6900 2171 7020 2451
rect 7603 2371 7723 2651
rect 7781 2371 7901 2651
rect 7959 2371 8079 2651
rect 8137 2371 8257 2651
rect 8315 2371 8435 2651
rect 8493 2371 8613 2651
rect 8671 2371 8791 2651
rect 8849 2371 8969 2651
rect 9027 2371 9147 2651
rect 9205 2371 9325 2651
rect 9383 2371 9503 2651
rect 9561 2371 9681 2651
rect 9739 2371 9859 2651
rect 9917 2371 10037 2651
rect 10290 2371 10410 2651
rect 10468 2371 10588 2651
rect 10646 2371 10766 2651
rect 10824 2371 10944 2651
rect 11002 2371 11122 2651
rect 11180 2371 11300 2651
rect 11358 2371 11478 2651
rect 11536 2371 11656 2651
rect 11714 2371 11834 2651
rect 11892 2371 12012 2651
rect 12070 2371 12190 2651
rect 12248 2371 12368 2651
rect 12426 2371 12546 2651
rect 12604 2371 12724 2651
rect 474 1671 594 1951
rect 652 1671 772 1951
rect 830 1671 950 1951
rect 1008 1671 1128 1951
rect 1186 1671 1306 1951
rect 1364 1671 1484 1951
rect 1542 1671 1662 1951
rect 1720 1671 1840 1951
rect 1898 1671 2018 1951
rect 2076 1671 2196 1951
rect 2254 1671 2374 1951
rect 2432 1671 2552 1951
rect 2610 1671 2730 1951
rect 2788 1671 2908 1951
rect 2966 1671 3086 1951
rect 3144 1671 3264 1951
rect 3322 1671 3442 1951
rect 3500 1671 3620 1951
rect 3874 1671 3994 1951
rect 4052 1671 4172 1951
rect 4230 1671 4350 1951
rect 4408 1671 4528 1951
rect 4586 1671 4706 1951
rect 4764 1671 4884 1951
rect 4942 1671 5062 1951
rect 5120 1671 5240 1951
rect 5298 1671 5418 1951
rect 5476 1671 5596 1951
rect 5654 1671 5774 1951
rect 5832 1671 5952 1951
rect 6010 1671 6130 1951
rect 6188 1671 6308 1951
rect 6366 1671 6486 1951
rect 6544 1671 6664 1951
rect 6722 1671 6842 1951
rect 6900 1671 7020 1951
rect 7603 1671 7723 1951
rect 7781 1671 7901 1951
rect 7959 1671 8079 1951
rect 8137 1671 8257 1951
rect 8315 1671 8435 1951
rect 8493 1671 8613 1951
rect 8671 1671 8791 1951
rect 8849 1671 8969 1951
rect 9027 1671 9147 1951
rect 9205 1671 9325 1951
rect 9383 1671 9503 1951
rect 9561 1671 9681 1951
rect 9739 1671 9859 1951
rect 9917 1671 10037 1951
rect 10290 1671 10410 1951
rect 10468 1671 10588 1951
rect 10646 1671 10766 1951
rect 10824 1671 10944 1951
rect 11002 1671 11122 1951
rect 11180 1671 11300 1951
rect 11358 1671 11478 1951
rect 11536 1671 11656 1951
rect 11714 1671 11834 1951
rect 11892 1671 12012 1951
rect 12070 1671 12190 1951
rect 12248 1671 12368 1951
rect 12426 1671 12546 1951
rect 12604 1671 12724 1951
rect 474 1171 594 1451
rect 652 1171 772 1451
rect 830 1171 950 1451
rect 1008 1171 1128 1451
rect 1186 1171 1306 1451
rect 1364 1171 1484 1451
rect 1542 1171 1662 1451
rect 1720 1171 1840 1451
rect 1898 1171 2018 1451
rect 2076 1171 2196 1451
rect 2254 1171 2374 1451
rect 2432 1171 2552 1451
rect 2610 1171 2730 1451
rect 2788 1171 2908 1451
rect 2966 1171 3086 1451
rect 3144 1171 3264 1451
rect 3322 1171 3442 1451
rect 3500 1171 3620 1451
rect 3874 1171 3994 1451
rect 4052 1171 4172 1451
rect 4230 1171 4350 1451
rect 4408 1171 4528 1451
rect 4586 1171 4706 1451
rect 4764 1171 4884 1451
rect 4942 1171 5062 1451
rect 5120 1171 5240 1451
rect 5298 1171 5418 1451
rect 5476 1171 5596 1451
rect 5654 1171 5774 1451
rect 5832 1171 5952 1451
rect 6010 1171 6130 1451
rect 6188 1171 6308 1451
rect 6366 1171 6486 1451
rect 6544 1171 6664 1451
rect 6722 1171 6842 1451
rect 6900 1171 7020 1451
rect 7603 1171 7723 1451
rect 7781 1171 7901 1451
rect 7959 1171 8079 1451
rect 8137 1171 8257 1451
rect 8315 1171 8435 1451
rect 8493 1171 8613 1451
rect 8671 1171 8791 1451
rect 8849 1171 8969 1451
rect 9027 1171 9147 1451
rect 9205 1171 9325 1451
rect 9383 1171 9503 1451
rect 9561 1171 9681 1451
rect 9739 1171 9859 1451
rect 9917 1171 10037 1451
rect 10290 1171 10410 1451
rect 10468 1171 10588 1451
rect 10646 1171 10766 1451
rect 10824 1171 10944 1451
rect 11002 1171 11122 1451
rect 11180 1171 11300 1451
rect 11358 1171 11478 1451
rect 11536 1171 11656 1451
rect 11714 1171 11834 1451
rect 11892 1171 12012 1451
rect 12070 1171 12190 1451
rect 12248 1171 12368 1451
rect 12426 1171 12546 1451
rect 12604 1171 12724 1451
rect 474 671 594 951
rect 652 671 772 951
rect 830 671 950 951
rect 1008 671 1128 951
rect 1186 671 1306 951
rect 1364 671 1484 951
rect 1542 671 1662 951
rect 1720 671 1840 951
rect 1898 671 2018 951
rect 2076 671 2196 951
rect 2254 671 2374 951
rect 2432 671 2552 951
rect 2610 671 2730 951
rect 2788 671 2908 951
rect 2966 671 3086 951
rect 3144 671 3264 951
rect 3322 671 3442 951
rect 3500 671 3620 951
rect 3874 671 3994 951
rect 4052 671 4172 951
rect 4230 671 4350 951
rect 4408 671 4528 951
rect 4586 671 4706 951
rect 4764 671 4884 951
rect 4942 671 5062 951
rect 5120 671 5240 951
rect 5298 671 5418 951
rect 5476 671 5596 951
rect 5654 671 5774 951
rect 5832 671 5952 951
rect 6010 671 6130 951
rect 6188 671 6308 951
rect 6366 671 6486 951
rect 6544 671 6664 951
rect 6722 671 6842 951
rect 6900 671 7020 951
rect 7603 671 7723 951
rect 7781 671 7901 951
rect 7959 671 8079 951
rect 8137 671 8257 951
rect 8315 671 8435 951
rect 8493 671 8613 951
rect 8671 671 8791 951
rect 8849 671 8969 951
rect 9027 671 9147 951
rect 9205 671 9325 951
rect 9383 671 9503 951
rect 9561 671 9681 951
rect 9739 671 9859 951
rect 9917 671 10037 951
rect 10290 671 10410 951
rect 10468 671 10588 951
rect 10646 671 10766 951
rect 10824 671 10944 951
rect 11002 671 11122 951
rect 11180 671 11300 951
rect 11358 671 11478 951
rect 11536 671 11656 951
rect 11714 671 11834 951
rect 11892 671 12012 951
rect 12070 671 12190 951
rect 12248 671 12368 951
rect 12426 671 12546 951
rect 12604 671 12724 951
rect 13596 4779 13716 5059
rect 13774 4779 13894 5059
rect 13952 4779 14072 5059
rect 14130 4779 14250 5059
rect 14308 4779 14428 5059
rect 14486 4779 14606 5059
rect 14664 4779 14784 5059
rect 14842 4779 14962 5059
rect 15020 4779 15140 5059
rect 15198 4779 15318 5059
rect 15376 4779 15496 5059
rect 15554 4779 15674 5059
rect 15732 4779 15852 5059
rect 15910 4779 16030 5059
rect 16088 4779 16208 5059
rect 16266 4779 16386 5059
rect 16444 4779 16564 5059
rect 16622 4779 16742 5059
rect 16800 4779 16920 5059
rect 16978 4779 17098 5059
rect 17156 4779 17276 5059
rect 17334 4779 17454 5059
rect 17512 4779 17632 5059
rect 17690 4779 17810 5059
rect 17868 4779 17988 5059
rect 18046 4779 18166 5059
rect 18224 4779 18344 5059
rect 13596 4279 13716 4559
rect 13774 4279 13894 4559
rect 13952 4279 14072 4559
rect 14130 4279 14250 4559
rect 14308 4279 14428 4559
rect 14486 4279 14606 4559
rect 14664 4279 14784 4559
rect 14842 4279 14962 4559
rect 15020 4279 15140 4559
rect 15198 4279 15318 4559
rect 15376 4279 15496 4559
rect 15554 4279 15674 4559
rect 15732 4279 15852 4559
rect 15910 4279 16030 4559
rect 16088 4279 16208 4559
rect 16266 4279 16386 4559
rect 16444 4279 16564 4559
rect 16622 4279 16742 4559
rect 16800 4279 16920 4559
rect 16978 4279 17098 4559
rect 17156 4279 17276 4559
rect 17334 4279 17454 4559
rect 17512 4279 17632 4559
rect 17690 4279 17810 4559
rect 17868 4279 17988 4559
rect 18046 4279 18166 4559
rect 18224 4279 18344 4559
rect 17154 3275 17274 3555
rect 17332 3275 17452 3555
rect 17510 3275 17630 3555
rect 17688 3275 17808 3555
rect 13722 2270 13842 2550
rect 14014 2270 14134 2550
rect 14306 2270 14426 2550
rect 14598 2270 14718 2550
rect 14890 2270 15010 2550
rect 15182 2270 15302 2550
rect 15474 2270 15594 2550
rect 16440 2336 16560 2616
rect 16618 2336 16738 2616
rect 16796 2336 16916 2616
rect 16974 2336 17094 2616
rect 17152 2336 17272 2616
rect 17330 2336 17450 2616
rect 17508 2336 17628 2616
rect 17686 2336 17806 2616
rect 17864 2336 17984 2616
rect 18042 2336 18162 2616
rect 18220 2336 18340 2616
rect 13722 1772 13842 2052
rect 14014 1772 14134 2052
rect 14306 1772 14426 2052
rect 14598 1772 14718 2052
rect 14890 1772 15010 2052
rect 15182 1772 15302 2052
rect 15474 1772 15594 2052
rect 16440 1836 16560 2116
rect 16618 1836 16738 2116
rect 16796 1836 16916 2116
rect 16974 1836 17094 2116
rect 17152 1836 17272 2116
rect 17330 1836 17450 2116
rect 17508 1836 17628 2116
rect 17686 1836 17806 2116
rect 17864 1836 17984 2116
rect 18042 1836 18162 2116
rect 18220 1836 18340 2116
rect 13722 1274 13842 1554
rect 14014 1274 14134 1554
rect 14306 1274 14426 1554
rect 14598 1274 14718 1554
rect 14890 1274 15010 1554
rect 15182 1274 15302 1554
rect 15474 1274 15594 1554
rect 16440 1276 16560 1556
rect 16618 1276 16738 1556
rect 16796 1276 16916 1556
rect 16974 1276 17094 1556
rect 17152 1276 17272 1556
rect 17330 1276 17450 1556
rect 17508 1276 17628 1556
rect 17686 1276 17806 1556
rect 17864 1276 17984 1556
rect 18042 1276 18162 1556
rect 18220 1276 18340 1556
rect 13722 776 13842 1056
rect 14014 776 14134 1056
rect 14306 776 14426 1056
rect 14598 776 14718 1056
rect 14890 776 15010 1056
rect 15182 776 15302 1056
rect 15474 776 15594 1056
rect 16440 776 16560 1056
rect 16618 776 16738 1056
rect 16796 776 16916 1056
rect 16974 776 17094 1056
rect 17152 776 17272 1056
rect 17330 776 17450 1056
rect 17508 776 17628 1056
rect 17686 776 17806 1056
rect 17864 776 17984 1056
rect 18042 776 18162 1056
rect 18220 776 18340 1056
rect 19413 2262 19533 2542
rect 19591 2262 19711 2542
rect 19769 2262 19889 2542
rect 19947 2262 20067 2542
rect 20125 2262 20245 2542
rect 20303 2262 20423 2542
rect 20481 2262 20601 2542
rect 20659 2262 20779 2542
rect 20837 2262 20957 2542
rect 21015 2262 21135 2542
rect 21193 2262 21313 2542
rect 19413 1764 19533 2044
rect 19591 1764 19711 2044
rect 19769 1764 19889 2044
rect 19947 1764 20067 2044
rect 20125 1764 20245 2044
rect 20303 1764 20423 2044
rect 20481 1764 20601 2044
rect 20659 1764 20779 2044
rect 20837 1764 20957 2044
rect 21015 1764 21135 2044
rect 21193 1764 21313 2044
rect 19413 1266 19533 1546
rect 19591 1266 19711 1546
rect 19769 1266 19889 1546
rect 19947 1266 20067 1546
rect 20125 1266 20245 1546
rect 20303 1266 20423 1546
rect 20481 1266 20601 1546
rect 20659 1266 20779 1546
rect 20837 1266 20957 1546
rect 21015 1266 21135 1546
rect 21193 1266 21313 1546
rect 19413 768 19533 1048
rect 19591 768 19711 1048
rect 19769 768 19889 1048
rect 19947 768 20067 1048
rect 20125 768 20245 1048
rect 20303 768 20423 1048
rect 20481 768 20601 1048
rect 20659 768 20779 1048
rect 20837 768 20957 1048
rect 21015 768 21135 1048
rect 21193 768 21313 1048
<< pmos >>
rect 7353 18481 7383 18753
rect 7449 18481 7479 18753
rect 7545 18481 7575 18753
rect 7641 18481 7671 18753
rect 7737 18481 7767 18753
rect 7833 18481 7863 18753
rect 7929 18481 7959 18753
rect 8025 18481 8055 18753
rect 8121 18481 8151 18753
rect 8217 18481 8247 18753
rect 20283 18481 20313 18753
rect 20379 18481 20409 18753
rect 20475 18481 20505 18753
rect 20571 18481 20601 18753
rect 20667 18481 20697 18753
rect 20763 18481 20793 18753
rect 20859 18481 20889 18753
rect 20955 18481 20985 18753
rect 21051 18481 21081 18753
rect 21147 18481 21177 18753
rect 7353 16681 7383 16953
rect 7449 16681 7479 16953
rect 7545 16681 7575 16953
rect 7641 16681 7671 16953
rect 7737 16681 7767 16953
rect 7833 16681 7863 16953
rect 7929 16681 7959 16953
rect 8025 16681 8055 16953
rect 8121 16681 8151 16953
rect 8217 16681 8247 16953
rect 20283 16681 20313 16953
rect 20379 16681 20409 16953
rect 20475 16681 20505 16953
rect 20571 16681 20601 16953
rect 20667 16681 20697 16953
rect 20763 16681 20793 16953
rect 20859 16681 20889 16953
rect 20955 16681 20985 16953
rect 21051 16681 21081 16953
rect 21147 16681 21177 16953
rect 7353 14881 7383 15153
rect 7449 14881 7479 15153
rect 7545 14881 7575 15153
rect 7641 14881 7671 15153
rect 7737 14881 7767 15153
rect 7833 14881 7863 15153
rect 7929 14881 7959 15153
rect 8025 14881 8055 15153
rect 8121 14881 8151 15153
rect 8217 14881 8247 15153
rect 20283 14881 20313 15153
rect 20379 14881 20409 15153
rect 20475 14881 20505 15153
rect 20571 14881 20601 15153
rect 20667 14881 20697 15153
rect 20763 14881 20793 15153
rect 20859 14881 20889 15153
rect 20955 14881 20985 15153
rect 21051 14881 21081 15153
rect 21147 14881 21177 15153
rect 7353 13081 7383 13353
rect 7449 13081 7479 13353
rect 7545 13081 7575 13353
rect 7641 13081 7671 13353
rect 7737 13081 7767 13353
rect 7833 13081 7863 13353
rect 7929 13081 7959 13353
rect 8025 13081 8055 13353
rect 8121 13081 8151 13353
rect 8217 13081 8247 13353
rect 20283 13081 20313 13353
rect 20379 13081 20409 13353
rect 20475 13081 20505 13353
rect 20571 13081 20601 13353
rect 20667 13081 20697 13353
rect 20763 13081 20793 13353
rect 20859 13081 20889 13353
rect 20955 13081 20985 13353
rect 21051 13081 21081 13353
rect 21147 13081 21177 13353
rect 7353 11281 7383 11553
rect 7449 11281 7479 11553
rect 7545 11281 7575 11553
rect 7641 11281 7671 11553
rect 7737 11281 7767 11553
rect 7833 11281 7863 11553
rect 7929 11281 7959 11553
rect 8025 11281 8055 11553
rect 8121 11281 8151 11553
rect 8217 11281 8247 11553
rect 20283 11281 20313 11553
rect 20379 11281 20409 11553
rect 20475 11281 20505 11553
rect 20571 11281 20601 11553
rect 20667 11281 20697 11553
rect 20763 11281 20793 11553
rect 20859 11281 20889 11553
rect 20955 11281 20985 11553
rect 21051 11281 21081 11553
rect 21147 11281 21177 11553
rect 7353 9481 7383 9753
rect 7449 9481 7479 9753
rect 7545 9481 7575 9753
rect 7641 9481 7671 9753
rect 7737 9481 7767 9753
rect 7833 9481 7863 9753
rect 7929 9481 7959 9753
rect 8025 9481 8055 9753
rect 8121 9481 8151 9753
rect 8217 9481 8247 9753
rect 20283 9481 20313 9753
rect 20379 9481 20409 9753
rect 20475 9481 20505 9753
rect 20571 9481 20601 9753
rect 20667 9481 20697 9753
rect 20763 9481 20793 9753
rect 20859 9481 20889 9753
rect 20955 9481 20985 9753
rect 21051 9481 21081 9753
rect 21147 9481 21177 9753
rect 14743 5631 14863 5911
rect 14921 5631 15041 5911
rect 15099 5631 15219 5911
rect 15277 5631 15397 5911
rect 15455 5631 15575 5911
rect 15633 5631 15753 5911
rect 15811 5631 15931 5911
rect 15989 5631 16109 5911
rect 16943 5631 17063 5911
rect 17121 5631 17241 5911
rect 17299 5631 17419 5911
rect 17477 5631 17597 5911
rect 17655 5631 17775 5911
rect 17833 5631 17953 5911
rect 18011 5631 18131 5911
rect 18189 5631 18309 5911
rect 19143 5631 19263 5911
rect 19321 5631 19441 5911
rect 19499 5631 19619 5911
rect 19677 5631 19797 5911
rect 19855 5631 19975 5911
rect 20033 5631 20153 5911
rect 20211 5631 20331 5911
rect 20389 5631 20509 5911
rect 7958 4871 8078 5151
rect 8136 4871 8256 5151
rect 8314 4871 8434 5151
rect 8492 4871 8612 5151
rect 8670 4871 8790 5151
rect 8848 4871 8968 5151
rect 9026 4871 9146 5151
rect 9204 4871 9324 5151
rect 9382 4871 9502 5151
rect 9560 4871 9680 5151
rect 9738 4871 9858 5151
rect 9916 4871 10036 5151
rect 10288 4871 10408 5151
rect 10466 4871 10586 5151
rect 10644 4871 10764 5151
rect 10822 4871 10942 5151
rect 11000 4871 11120 5151
rect 11178 4871 11298 5151
rect 11356 4871 11476 5151
rect 11534 4871 11654 5151
rect 11712 4871 11832 5151
rect 11890 4871 12010 5151
rect 12068 4871 12188 5151
rect 12246 4871 12366 5151
rect 7958 4301 8078 4581
rect 8136 4301 8256 4581
rect 8314 4301 8434 4581
rect 8492 4301 8612 4581
rect 8670 4301 8790 4581
rect 8848 4301 8968 4581
rect 9026 4301 9146 4581
rect 9204 4301 9324 4581
rect 9382 4301 9502 4581
rect 9560 4301 9680 4581
rect 9738 4301 9858 4581
rect 9916 4301 10036 4581
rect 10288 4301 10408 4581
rect 10466 4301 10586 4581
rect 10644 4301 10764 4581
rect 10822 4301 10942 4581
rect 11000 4301 11120 4581
rect 11178 4301 11298 4581
rect 11356 4301 11476 4581
rect 11534 4301 11654 4581
rect 11712 4301 11832 4581
rect 11890 4301 12010 4581
rect 12068 4301 12188 4581
rect 12246 4301 12366 4581
<< pmoslvt >>
rect 7602 6329 7722 6609
rect 7780 6329 7900 6609
rect 7958 6329 8078 6609
rect 8136 6329 8256 6609
rect 8314 6329 8434 6609
rect 8492 6329 8612 6609
rect 8670 6329 8790 6609
rect 8848 6329 8968 6609
rect 9026 6329 9146 6609
rect 9204 6329 9324 6609
rect 9382 6329 9502 6609
rect 9560 6329 9680 6609
rect 9738 6329 9858 6609
rect 9916 6329 10036 6609
rect 10288 6329 10408 6609
rect 10466 6329 10586 6609
rect 10644 6329 10764 6609
rect 10822 6329 10942 6609
rect 11000 6329 11120 6609
rect 11178 6329 11298 6609
rect 11356 6329 11476 6609
rect 11534 6329 11654 6609
rect 11712 6329 11832 6609
rect 11890 6329 12010 6609
rect 12068 6329 12188 6609
rect 12246 6329 12366 6609
rect 12424 6329 12544 6609
rect 12602 6329 12722 6609
rect 7602 5751 7722 6031
rect 7780 5751 7900 6031
rect 7958 5751 8078 6031
rect 8136 5751 8256 6031
rect 8314 5751 8434 6031
rect 8492 5751 8612 6031
rect 8670 5751 8790 6031
rect 8848 5751 8968 6031
rect 9026 5751 9146 6031
rect 9204 5751 9324 6031
rect 9382 5751 9502 6031
rect 9560 5751 9680 6031
rect 9738 5751 9858 6031
rect 9916 5751 10036 6031
rect 10288 5752 10408 6032
rect 10466 5752 10586 6032
rect 10644 5752 10764 6032
rect 10822 5752 10942 6032
rect 11000 5752 11120 6032
rect 11178 5752 11298 6032
rect 11356 5752 11476 6032
rect 11534 5752 11654 6032
rect 11712 5752 11832 6032
rect 11890 5752 12010 6032
rect 12068 5752 12188 6032
rect 12246 5752 12366 6032
rect 12424 5752 12544 6032
rect 12602 5752 12722 6032
rect 14742 6398 14862 6678
rect 14920 6398 15040 6678
rect 15098 6398 15218 6678
rect 15276 6398 15396 6678
rect 15454 6398 15574 6678
rect 15632 6398 15752 6678
rect 15810 6398 15930 6678
rect 15988 6398 16108 6678
rect 16942 6398 17062 6678
rect 17120 6398 17240 6678
rect 17298 6398 17418 6678
rect 17476 6398 17596 6678
rect 17654 6398 17774 6678
rect 17832 6398 17952 6678
rect 18010 6398 18130 6678
rect 18188 6398 18308 6678
rect 19142 6398 19262 6678
rect 19320 6398 19440 6678
rect 19498 6398 19618 6678
rect 19676 6398 19796 6678
rect 19854 6398 19974 6678
rect 20032 6398 20152 6678
rect 20210 6398 20330 6678
rect 20388 6398 20508 6678
<< nmoslvt >>
rect 2096 3991 2136 4231
rect 2308 3991 2348 4231
rect 2520 3991 2560 4231
rect 2732 3991 2772 4231
rect 2944 3991 2984 4231
rect 3156 3991 3196 4231
rect 3368 3991 3408 4231
rect 3580 3991 3620 4231
rect 3876 3991 3916 4231
rect 4088 3991 4128 4231
rect 4300 3991 4340 4231
rect 4512 3991 4552 4231
rect 4724 3991 4764 4231
rect 4936 3991 4976 4231
rect 5148 3991 5188 4231
rect 5360 3991 5400 4231
rect 19055 4770 19175 5050
rect 19233 4770 19353 5050
rect 19411 4770 19531 5050
rect 19589 4770 19709 5050
rect 19767 4770 19887 5050
rect 19945 4770 20065 5050
rect 20123 4770 20243 5050
rect 20301 4770 20421 5050
rect 20479 4770 20599 5050
rect 20657 4770 20777 5050
rect 20835 4770 20955 5050
rect 21013 4770 21133 5050
rect 21191 4770 21311 5050
rect 21369 4770 21489 5050
rect 21547 4770 21667 5050
rect 21725 4770 21845 5050
rect 19055 4272 19175 4552
rect 19233 4272 19353 4552
rect 19411 4272 19531 4552
rect 19589 4272 19709 4552
rect 19767 4272 19887 4552
rect 19945 4272 20065 4552
rect 20123 4272 20243 4552
rect 20301 4272 20421 4552
rect 20479 4272 20599 4552
rect 20657 4272 20777 4552
rect 20835 4272 20955 4552
rect 21013 4272 21133 4552
rect 21191 4272 21311 4552
rect 21369 4272 21489 4552
rect 21547 4272 21667 4552
rect 21725 4272 21845 4552
rect 19055 3774 19175 4054
rect 19233 3774 19353 4054
rect 19411 3774 19531 4054
rect 19589 3774 19709 4054
rect 19767 3774 19887 4054
rect 19945 3774 20065 4054
rect 20123 3774 20243 4054
rect 20301 3774 20421 4054
rect 20479 3774 20599 4054
rect 20657 3774 20777 4054
rect 20835 3774 20955 4054
rect 21013 3774 21133 4054
rect 21191 3774 21311 4054
rect 21369 3774 21489 4054
rect 21547 3774 21667 4054
rect 21725 3774 21845 4054
rect 19055 3276 19175 3556
rect 19233 3276 19353 3556
rect 19411 3276 19531 3556
rect 19589 3276 19709 3556
rect 19767 3276 19887 3556
rect 19945 3276 20065 3556
rect 20123 3276 20243 3556
rect 20301 3276 20421 3556
rect 20479 3276 20599 3556
rect 20657 3276 20777 3556
rect 20835 3276 20955 3556
rect 21013 3276 21133 3556
rect 21191 3276 21311 3556
rect 21369 3276 21489 3556
rect 21547 3276 21667 3556
rect 21725 3276 21845 3556
<< ndiff >>
rect 7291 18163 7353 18175
rect 7291 18083 7303 18163
rect 7337 18083 7353 18163
rect 7291 18071 7353 18083
rect 7383 18163 7449 18175
rect 7383 18083 7399 18163
rect 7433 18083 7449 18163
rect 7383 18071 7449 18083
rect 7479 18163 7545 18175
rect 7479 18083 7495 18163
rect 7529 18083 7545 18163
rect 7479 18071 7545 18083
rect 7575 18163 7641 18175
rect 7575 18083 7591 18163
rect 7625 18083 7641 18163
rect 7575 18071 7641 18083
rect 7671 18163 7737 18175
rect 7671 18083 7687 18163
rect 7721 18083 7737 18163
rect 7671 18071 7737 18083
rect 7767 18163 7833 18175
rect 7767 18083 7783 18163
rect 7817 18083 7833 18163
rect 7767 18071 7833 18083
rect 7863 18163 7929 18175
rect 7863 18083 7879 18163
rect 7913 18083 7929 18163
rect 7863 18071 7929 18083
rect 7959 18163 8025 18175
rect 7959 18083 7975 18163
rect 8009 18083 8025 18163
rect 7959 18071 8025 18083
rect 8055 18163 8121 18175
rect 8055 18083 8071 18163
rect 8105 18083 8121 18163
rect 8055 18071 8121 18083
rect 8151 18163 8217 18175
rect 8151 18083 8167 18163
rect 8201 18083 8217 18163
rect 8151 18071 8217 18083
rect 8247 18163 8309 18175
rect 8247 18083 8263 18163
rect 8297 18083 8309 18163
rect 8247 18071 8309 18083
rect 20221 18163 20283 18175
rect 20221 18083 20233 18163
rect 20267 18083 20283 18163
rect 20221 18071 20283 18083
rect 20313 18163 20379 18175
rect 20313 18083 20329 18163
rect 20363 18083 20379 18163
rect 20313 18071 20379 18083
rect 20409 18163 20475 18175
rect 20409 18083 20425 18163
rect 20459 18083 20475 18163
rect 20409 18071 20475 18083
rect 20505 18163 20571 18175
rect 20505 18083 20521 18163
rect 20555 18083 20571 18163
rect 20505 18071 20571 18083
rect 20601 18163 20667 18175
rect 20601 18083 20617 18163
rect 20651 18083 20667 18163
rect 20601 18071 20667 18083
rect 20697 18163 20763 18175
rect 20697 18083 20713 18163
rect 20747 18083 20763 18163
rect 20697 18071 20763 18083
rect 20793 18163 20859 18175
rect 20793 18083 20809 18163
rect 20843 18083 20859 18163
rect 20793 18071 20859 18083
rect 20889 18163 20955 18175
rect 20889 18083 20905 18163
rect 20939 18083 20955 18163
rect 20889 18071 20955 18083
rect 20985 18163 21051 18175
rect 20985 18083 21001 18163
rect 21035 18083 21051 18163
rect 20985 18071 21051 18083
rect 21081 18163 21147 18175
rect 21081 18083 21097 18163
rect 21131 18083 21147 18163
rect 21081 18071 21147 18083
rect 21177 18163 21239 18175
rect 21177 18083 21193 18163
rect 21227 18083 21239 18163
rect 21177 18071 21239 18083
rect 7291 16363 7353 16375
rect 7291 16283 7303 16363
rect 7337 16283 7353 16363
rect 7291 16271 7353 16283
rect 7383 16363 7449 16375
rect 7383 16283 7399 16363
rect 7433 16283 7449 16363
rect 7383 16271 7449 16283
rect 7479 16363 7545 16375
rect 7479 16283 7495 16363
rect 7529 16283 7545 16363
rect 7479 16271 7545 16283
rect 7575 16363 7641 16375
rect 7575 16283 7591 16363
rect 7625 16283 7641 16363
rect 7575 16271 7641 16283
rect 7671 16363 7737 16375
rect 7671 16283 7687 16363
rect 7721 16283 7737 16363
rect 7671 16271 7737 16283
rect 7767 16363 7833 16375
rect 7767 16283 7783 16363
rect 7817 16283 7833 16363
rect 7767 16271 7833 16283
rect 7863 16363 7929 16375
rect 7863 16283 7879 16363
rect 7913 16283 7929 16363
rect 7863 16271 7929 16283
rect 7959 16363 8025 16375
rect 7959 16283 7975 16363
rect 8009 16283 8025 16363
rect 7959 16271 8025 16283
rect 8055 16363 8121 16375
rect 8055 16283 8071 16363
rect 8105 16283 8121 16363
rect 8055 16271 8121 16283
rect 8151 16363 8217 16375
rect 8151 16283 8167 16363
rect 8201 16283 8217 16363
rect 8151 16271 8217 16283
rect 8247 16363 8309 16375
rect 8247 16283 8263 16363
rect 8297 16283 8309 16363
rect 8247 16271 8309 16283
rect 20221 16363 20283 16375
rect 20221 16283 20233 16363
rect 20267 16283 20283 16363
rect 20221 16271 20283 16283
rect 20313 16363 20379 16375
rect 20313 16283 20329 16363
rect 20363 16283 20379 16363
rect 20313 16271 20379 16283
rect 20409 16363 20475 16375
rect 20409 16283 20425 16363
rect 20459 16283 20475 16363
rect 20409 16271 20475 16283
rect 20505 16363 20571 16375
rect 20505 16283 20521 16363
rect 20555 16283 20571 16363
rect 20505 16271 20571 16283
rect 20601 16363 20667 16375
rect 20601 16283 20617 16363
rect 20651 16283 20667 16363
rect 20601 16271 20667 16283
rect 20697 16363 20763 16375
rect 20697 16283 20713 16363
rect 20747 16283 20763 16363
rect 20697 16271 20763 16283
rect 20793 16363 20859 16375
rect 20793 16283 20809 16363
rect 20843 16283 20859 16363
rect 20793 16271 20859 16283
rect 20889 16363 20955 16375
rect 20889 16283 20905 16363
rect 20939 16283 20955 16363
rect 20889 16271 20955 16283
rect 20985 16363 21051 16375
rect 20985 16283 21001 16363
rect 21035 16283 21051 16363
rect 20985 16271 21051 16283
rect 21081 16363 21147 16375
rect 21081 16283 21097 16363
rect 21131 16283 21147 16363
rect 21081 16271 21147 16283
rect 21177 16363 21239 16375
rect 21177 16283 21193 16363
rect 21227 16283 21239 16363
rect 21177 16271 21239 16283
rect 7291 14563 7353 14575
rect 7291 14483 7303 14563
rect 7337 14483 7353 14563
rect 7291 14471 7353 14483
rect 7383 14563 7449 14575
rect 7383 14483 7399 14563
rect 7433 14483 7449 14563
rect 7383 14471 7449 14483
rect 7479 14563 7545 14575
rect 7479 14483 7495 14563
rect 7529 14483 7545 14563
rect 7479 14471 7545 14483
rect 7575 14563 7641 14575
rect 7575 14483 7591 14563
rect 7625 14483 7641 14563
rect 7575 14471 7641 14483
rect 7671 14563 7737 14575
rect 7671 14483 7687 14563
rect 7721 14483 7737 14563
rect 7671 14471 7737 14483
rect 7767 14563 7833 14575
rect 7767 14483 7783 14563
rect 7817 14483 7833 14563
rect 7767 14471 7833 14483
rect 7863 14563 7929 14575
rect 7863 14483 7879 14563
rect 7913 14483 7929 14563
rect 7863 14471 7929 14483
rect 7959 14563 8025 14575
rect 7959 14483 7975 14563
rect 8009 14483 8025 14563
rect 7959 14471 8025 14483
rect 8055 14563 8121 14575
rect 8055 14483 8071 14563
rect 8105 14483 8121 14563
rect 8055 14471 8121 14483
rect 8151 14563 8217 14575
rect 8151 14483 8167 14563
rect 8201 14483 8217 14563
rect 8151 14471 8217 14483
rect 8247 14563 8309 14575
rect 8247 14483 8263 14563
rect 8297 14483 8309 14563
rect 8247 14471 8309 14483
rect 20221 14563 20283 14575
rect 20221 14483 20233 14563
rect 20267 14483 20283 14563
rect 20221 14471 20283 14483
rect 20313 14563 20379 14575
rect 20313 14483 20329 14563
rect 20363 14483 20379 14563
rect 20313 14471 20379 14483
rect 20409 14563 20475 14575
rect 20409 14483 20425 14563
rect 20459 14483 20475 14563
rect 20409 14471 20475 14483
rect 20505 14563 20571 14575
rect 20505 14483 20521 14563
rect 20555 14483 20571 14563
rect 20505 14471 20571 14483
rect 20601 14563 20667 14575
rect 20601 14483 20617 14563
rect 20651 14483 20667 14563
rect 20601 14471 20667 14483
rect 20697 14563 20763 14575
rect 20697 14483 20713 14563
rect 20747 14483 20763 14563
rect 20697 14471 20763 14483
rect 20793 14563 20859 14575
rect 20793 14483 20809 14563
rect 20843 14483 20859 14563
rect 20793 14471 20859 14483
rect 20889 14563 20955 14575
rect 20889 14483 20905 14563
rect 20939 14483 20955 14563
rect 20889 14471 20955 14483
rect 20985 14563 21051 14575
rect 20985 14483 21001 14563
rect 21035 14483 21051 14563
rect 20985 14471 21051 14483
rect 21081 14563 21147 14575
rect 21081 14483 21097 14563
rect 21131 14483 21147 14563
rect 21081 14471 21147 14483
rect 21177 14563 21239 14575
rect 21177 14483 21193 14563
rect 21227 14483 21239 14563
rect 21177 14471 21239 14483
rect 7291 12763 7353 12775
rect 7291 12683 7303 12763
rect 7337 12683 7353 12763
rect 7291 12671 7353 12683
rect 7383 12763 7449 12775
rect 7383 12683 7399 12763
rect 7433 12683 7449 12763
rect 7383 12671 7449 12683
rect 7479 12763 7545 12775
rect 7479 12683 7495 12763
rect 7529 12683 7545 12763
rect 7479 12671 7545 12683
rect 7575 12763 7641 12775
rect 7575 12683 7591 12763
rect 7625 12683 7641 12763
rect 7575 12671 7641 12683
rect 7671 12763 7737 12775
rect 7671 12683 7687 12763
rect 7721 12683 7737 12763
rect 7671 12671 7737 12683
rect 7767 12763 7833 12775
rect 7767 12683 7783 12763
rect 7817 12683 7833 12763
rect 7767 12671 7833 12683
rect 7863 12763 7929 12775
rect 7863 12683 7879 12763
rect 7913 12683 7929 12763
rect 7863 12671 7929 12683
rect 7959 12763 8025 12775
rect 7959 12683 7975 12763
rect 8009 12683 8025 12763
rect 7959 12671 8025 12683
rect 8055 12763 8121 12775
rect 8055 12683 8071 12763
rect 8105 12683 8121 12763
rect 8055 12671 8121 12683
rect 8151 12763 8217 12775
rect 8151 12683 8167 12763
rect 8201 12683 8217 12763
rect 8151 12671 8217 12683
rect 8247 12763 8309 12775
rect 8247 12683 8263 12763
rect 8297 12683 8309 12763
rect 8247 12671 8309 12683
rect 20221 12763 20283 12775
rect 20221 12683 20233 12763
rect 20267 12683 20283 12763
rect 20221 12671 20283 12683
rect 20313 12763 20379 12775
rect 20313 12683 20329 12763
rect 20363 12683 20379 12763
rect 20313 12671 20379 12683
rect 20409 12763 20475 12775
rect 20409 12683 20425 12763
rect 20459 12683 20475 12763
rect 20409 12671 20475 12683
rect 20505 12763 20571 12775
rect 20505 12683 20521 12763
rect 20555 12683 20571 12763
rect 20505 12671 20571 12683
rect 20601 12763 20667 12775
rect 20601 12683 20617 12763
rect 20651 12683 20667 12763
rect 20601 12671 20667 12683
rect 20697 12763 20763 12775
rect 20697 12683 20713 12763
rect 20747 12683 20763 12763
rect 20697 12671 20763 12683
rect 20793 12763 20859 12775
rect 20793 12683 20809 12763
rect 20843 12683 20859 12763
rect 20793 12671 20859 12683
rect 20889 12763 20955 12775
rect 20889 12683 20905 12763
rect 20939 12683 20955 12763
rect 20889 12671 20955 12683
rect 20985 12763 21051 12775
rect 20985 12683 21001 12763
rect 21035 12683 21051 12763
rect 20985 12671 21051 12683
rect 21081 12763 21147 12775
rect 21081 12683 21097 12763
rect 21131 12683 21147 12763
rect 21081 12671 21147 12683
rect 21177 12763 21239 12775
rect 21177 12683 21193 12763
rect 21227 12683 21239 12763
rect 21177 12671 21239 12683
rect 7291 10963 7353 10975
rect 7291 10883 7303 10963
rect 7337 10883 7353 10963
rect 7291 10871 7353 10883
rect 7383 10963 7449 10975
rect 7383 10883 7399 10963
rect 7433 10883 7449 10963
rect 7383 10871 7449 10883
rect 7479 10963 7545 10975
rect 7479 10883 7495 10963
rect 7529 10883 7545 10963
rect 7479 10871 7545 10883
rect 7575 10963 7641 10975
rect 7575 10883 7591 10963
rect 7625 10883 7641 10963
rect 7575 10871 7641 10883
rect 7671 10963 7737 10975
rect 7671 10883 7687 10963
rect 7721 10883 7737 10963
rect 7671 10871 7737 10883
rect 7767 10963 7833 10975
rect 7767 10883 7783 10963
rect 7817 10883 7833 10963
rect 7767 10871 7833 10883
rect 7863 10963 7929 10975
rect 7863 10883 7879 10963
rect 7913 10883 7929 10963
rect 7863 10871 7929 10883
rect 7959 10963 8025 10975
rect 7959 10883 7975 10963
rect 8009 10883 8025 10963
rect 7959 10871 8025 10883
rect 8055 10963 8121 10975
rect 8055 10883 8071 10963
rect 8105 10883 8121 10963
rect 8055 10871 8121 10883
rect 8151 10963 8217 10975
rect 8151 10883 8167 10963
rect 8201 10883 8217 10963
rect 8151 10871 8217 10883
rect 8247 10963 8309 10975
rect 8247 10883 8263 10963
rect 8297 10883 8309 10963
rect 8247 10871 8309 10883
rect 20221 10963 20283 10975
rect 20221 10883 20233 10963
rect 20267 10883 20283 10963
rect 20221 10871 20283 10883
rect 20313 10963 20379 10975
rect 20313 10883 20329 10963
rect 20363 10883 20379 10963
rect 20313 10871 20379 10883
rect 20409 10963 20475 10975
rect 20409 10883 20425 10963
rect 20459 10883 20475 10963
rect 20409 10871 20475 10883
rect 20505 10963 20571 10975
rect 20505 10883 20521 10963
rect 20555 10883 20571 10963
rect 20505 10871 20571 10883
rect 20601 10963 20667 10975
rect 20601 10883 20617 10963
rect 20651 10883 20667 10963
rect 20601 10871 20667 10883
rect 20697 10963 20763 10975
rect 20697 10883 20713 10963
rect 20747 10883 20763 10963
rect 20697 10871 20763 10883
rect 20793 10963 20859 10975
rect 20793 10883 20809 10963
rect 20843 10883 20859 10963
rect 20793 10871 20859 10883
rect 20889 10963 20955 10975
rect 20889 10883 20905 10963
rect 20939 10883 20955 10963
rect 20889 10871 20955 10883
rect 20985 10963 21051 10975
rect 20985 10883 21001 10963
rect 21035 10883 21051 10963
rect 20985 10871 21051 10883
rect 21081 10963 21147 10975
rect 21081 10883 21097 10963
rect 21131 10883 21147 10963
rect 21081 10871 21147 10883
rect 21177 10963 21239 10975
rect 21177 10883 21193 10963
rect 21227 10883 21239 10963
rect 21177 10871 21239 10883
rect 7291 9163 7353 9175
rect 7291 9083 7303 9163
rect 7337 9083 7353 9163
rect 7291 9071 7353 9083
rect 7383 9163 7449 9175
rect 7383 9083 7399 9163
rect 7433 9083 7449 9163
rect 7383 9071 7449 9083
rect 7479 9163 7545 9175
rect 7479 9083 7495 9163
rect 7529 9083 7545 9163
rect 7479 9071 7545 9083
rect 7575 9163 7641 9175
rect 7575 9083 7591 9163
rect 7625 9083 7641 9163
rect 7575 9071 7641 9083
rect 7671 9163 7737 9175
rect 7671 9083 7687 9163
rect 7721 9083 7737 9163
rect 7671 9071 7737 9083
rect 7767 9163 7833 9175
rect 7767 9083 7783 9163
rect 7817 9083 7833 9163
rect 7767 9071 7833 9083
rect 7863 9163 7929 9175
rect 7863 9083 7879 9163
rect 7913 9083 7929 9163
rect 7863 9071 7929 9083
rect 7959 9163 8025 9175
rect 7959 9083 7975 9163
rect 8009 9083 8025 9163
rect 7959 9071 8025 9083
rect 8055 9163 8121 9175
rect 8055 9083 8071 9163
rect 8105 9083 8121 9163
rect 8055 9071 8121 9083
rect 8151 9163 8217 9175
rect 8151 9083 8167 9163
rect 8201 9083 8217 9163
rect 8151 9071 8217 9083
rect 8247 9163 8309 9175
rect 8247 9083 8263 9163
rect 8297 9083 8309 9163
rect 8247 9071 8309 9083
rect 20221 9163 20283 9175
rect 20221 9083 20233 9163
rect 20267 9083 20283 9163
rect 20221 9071 20283 9083
rect 20313 9163 20379 9175
rect 20313 9083 20329 9163
rect 20363 9083 20379 9163
rect 20313 9071 20379 9083
rect 20409 9163 20475 9175
rect 20409 9083 20425 9163
rect 20459 9083 20475 9163
rect 20409 9071 20475 9083
rect 20505 9163 20571 9175
rect 20505 9083 20521 9163
rect 20555 9083 20571 9163
rect 20505 9071 20571 9083
rect 20601 9163 20667 9175
rect 20601 9083 20617 9163
rect 20651 9083 20667 9163
rect 20601 9071 20667 9083
rect 20697 9163 20763 9175
rect 20697 9083 20713 9163
rect 20747 9083 20763 9163
rect 20697 9071 20763 9083
rect 20793 9163 20859 9175
rect 20793 9083 20809 9163
rect 20843 9083 20859 9163
rect 20793 9071 20859 9083
rect 20889 9163 20955 9175
rect 20889 9083 20905 9163
rect 20939 9083 20955 9163
rect 20889 9071 20955 9083
rect 20985 9163 21051 9175
rect 20985 9083 21001 9163
rect 21035 9083 21051 9163
rect 20985 9071 21051 9083
rect 21081 9163 21147 9175
rect 21081 9083 21097 9163
rect 21131 9083 21147 9163
rect 21081 9071 21147 9083
rect 21177 9163 21239 9175
rect 21177 9083 21193 9163
rect 21227 9083 21239 9163
rect 21177 9071 21239 9083
rect 2038 4219 2096 4231
rect 2038 4003 2050 4219
rect 2084 4003 2096 4219
rect 2038 3991 2096 4003
rect 2136 4219 2194 4231
rect 2136 4003 2148 4219
rect 2182 4003 2194 4219
rect 2136 3991 2194 4003
rect 2250 4219 2308 4231
rect 2250 4003 2262 4219
rect 2296 4003 2308 4219
rect 2250 3991 2308 4003
rect 2348 4219 2406 4231
rect 2348 4003 2360 4219
rect 2394 4003 2406 4219
rect 2348 3991 2406 4003
rect 2462 4219 2520 4231
rect 2462 4003 2474 4219
rect 2508 4003 2520 4219
rect 2462 3991 2520 4003
rect 2560 4219 2618 4231
rect 2560 4003 2572 4219
rect 2606 4003 2618 4219
rect 2560 3991 2618 4003
rect 2674 4219 2732 4231
rect 2674 4003 2686 4219
rect 2720 4003 2732 4219
rect 2674 3991 2732 4003
rect 2772 4219 2830 4231
rect 2772 4003 2784 4219
rect 2818 4003 2830 4219
rect 2772 3991 2830 4003
rect 2886 4219 2944 4231
rect 2886 4003 2898 4219
rect 2932 4003 2944 4219
rect 2886 3991 2944 4003
rect 2984 4219 3042 4231
rect 2984 4003 2996 4219
rect 3030 4003 3042 4219
rect 2984 3991 3042 4003
rect 3098 4219 3156 4231
rect 3098 4003 3110 4219
rect 3144 4003 3156 4219
rect 3098 3991 3156 4003
rect 3196 4219 3254 4231
rect 3196 4003 3208 4219
rect 3242 4003 3254 4219
rect 3196 3991 3254 4003
rect 3310 4219 3368 4231
rect 3310 4003 3322 4219
rect 3356 4003 3368 4219
rect 3310 3991 3368 4003
rect 3408 4219 3466 4231
rect 3408 4003 3420 4219
rect 3454 4003 3466 4219
rect 3408 3991 3466 4003
rect 3522 4219 3580 4231
rect 3522 4003 3534 4219
rect 3568 4003 3580 4219
rect 3522 3991 3580 4003
rect 3620 4219 3678 4231
rect 3620 4003 3632 4219
rect 3666 4003 3678 4219
rect 3620 3991 3678 4003
rect 3818 4219 3876 4231
rect 3818 4003 3830 4219
rect 3864 4003 3876 4219
rect 3818 3991 3876 4003
rect 3916 4219 3974 4231
rect 3916 4003 3928 4219
rect 3962 4003 3974 4219
rect 3916 3991 3974 4003
rect 4030 4219 4088 4231
rect 4030 4003 4042 4219
rect 4076 4003 4088 4219
rect 4030 3991 4088 4003
rect 4128 4219 4186 4231
rect 4128 4003 4140 4219
rect 4174 4003 4186 4219
rect 4128 3991 4186 4003
rect 4242 4219 4300 4231
rect 4242 4003 4254 4219
rect 4288 4003 4300 4219
rect 4242 3991 4300 4003
rect 4340 4219 4398 4231
rect 4340 4003 4352 4219
rect 4386 4003 4398 4219
rect 4340 3991 4398 4003
rect 4454 4219 4512 4231
rect 4454 4003 4466 4219
rect 4500 4003 4512 4219
rect 4454 3991 4512 4003
rect 4552 4219 4610 4231
rect 4552 4003 4564 4219
rect 4598 4003 4610 4219
rect 4552 3991 4610 4003
rect 4666 4219 4724 4231
rect 4666 4003 4678 4219
rect 4712 4003 4724 4219
rect 4666 3991 4724 4003
rect 4764 4219 4822 4231
rect 4764 4003 4776 4219
rect 4810 4003 4822 4219
rect 4764 3991 4822 4003
rect 4878 4219 4936 4231
rect 4878 4003 4890 4219
rect 4924 4003 4936 4219
rect 4878 3991 4936 4003
rect 4976 4219 5034 4231
rect 4976 4003 4988 4219
rect 5022 4003 5034 4219
rect 4976 3991 5034 4003
rect 5090 4219 5148 4231
rect 5090 4003 5102 4219
rect 5136 4003 5148 4219
rect 5090 3991 5148 4003
rect 5188 4219 5246 4231
rect 5188 4003 5200 4219
rect 5234 4003 5246 4219
rect 5188 3991 5246 4003
rect 5302 4219 5360 4231
rect 5302 4003 5314 4219
rect 5348 4003 5360 4219
rect 5302 3991 5360 4003
rect 5400 4219 5458 4231
rect 5400 4003 5412 4219
rect 5446 4003 5458 4219
rect 5400 3991 5458 4003
rect 7545 3639 7603 3651
rect 416 3439 474 3451
rect 416 3183 428 3439
rect 462 3183 474 3439
rect 416 3171 474 3183
rect 594 3439 652 3451
rect 594 3183 606 3439
rect 640 3183 652 3439
rect 594 3171 652 3183
rect 772 3439 830 3451
rect 772 3183 784 3439
rect 818 3183 830 3439
rect 772 3171 830 3183
rect 950 3439 1008 3451
rect 950 3183 962 3439
rect 996 3183 1008 3439
rect 950 3171 1008 3183
rect 1128 3439 1186 3451
rect 1128 3183 1140 3439
rect 1174 3183 1186 3439
rect 1128 3171 1186 3183
rect 1306 3439 1364 3451
rect 1306 3183 1318 3439
rect 1352 3183 1364 3439
rect 1306 3171 1364 3183
rect 1484 3439 1542 3451
rect 1484 3183 1496 3439
rect 1530 3183 1542 3439
rect 1484 3171 1542 3183
rect 1662 3439 1720 3451
rect 1662 3183 1674 3439
rect 1708 3183 1720 3439
rect 1662 3171 1720 3183
rect 1840 3439 1898 3451
rect 1840 3183 1852 3439
rect 1886 3183 1898 3439
rect 1840 3171 1898 3183
rect 2018 3439 2076 3451
rect 2018 3183 2030 3439
rect 2064 3183 2076 3439
rect 2018 3171 2076 3183
rect 2196 3439 2254 3451
rect 2196 3183 2208 3439
rect 2242 3183 2254 3439
rect 2196 3171 2254 3183
rect 2374 3439 2432 3451
rect 2374 3183 2386 3439
rect 2420 3183 2432 3439
rect 2374 3171 2432 3183
rect 2552 3439 2610 3451
rect 2552 3183 2564 3439
rect 2598 3183 2610 3439
rect 2552 3171 2610 3183
rect 2730 3439 2788 3451
rect 2730 3183 2742 3439
rect 2776 3183 2788 3439
rect 2730 3171 2788 3183
rect 2908 3439 2966 3451
rect 2908 3183 2920 3439
rect 2954 3183 2966 3439
rect 2908 3171 2966 3183
rect 3086 3439 3144 3451
rect 3086 3183 3098 3439
rect 3132 3183 3144 3439
rect 3086 3171 3144 3183
rect 3264 3439 3322 3451
rect 3264 3183 3276 3439
rect 3310 3183 3322 3439
rect 3264 3171 3322 3183
rect 3442 3439 3500 3451
rect 3442 3183 3454 3439
rect 3488 3183 3500 3439
rect 3442 3171 3500 3183
rect 3620 3439 3678 3451
rect 3620 3183 3632 3439
rect 3666 3183 3678 3439
rect 3620 3171 3678 3183
rect 3816 3439 3874 3451
rect 3816 3183 3828 3439
rect 3862 3183 3874 3439
rect 3816 3171 3874 3183
rect 3994 3439 4052 3451
rect 3994 3183 4006 3439
rect 4040 3183 4052 3439
rect 3994 3171 4052 3183
rect 4172 3439 4230 3451
rect 4172 3183 4184 3439
rect 4218 3183 4230 3439
rect 4172 3171 4230 3183
rect 4350 3439 4408 3451
rect 4350 3183 4362 3439
rect 4396 3183 4408 3439
rect 4350 3171 4408 3183
rect 4528 3439 4586 3451
rect 4528 3183 4540 3439
rect 4574 3183 4586 3439
rect 4528 3171 4586 3183
rect 4706 3439 4764 3451
rect 4706 3183 4718 3439
rect 4752 3183 4764 3439
rect 4706 3171 4764 3183
rect 4884 3439 4942 3451
rect 4884 3183 4896 3439
rect 4930 3183 4942 3439
rect 4884 3171 4942 3183
rect 5062 3439 5120 3451
rect 5062 3183 5074 3439
rect 5108 3183 5120 3439
rect 5062 3171 5120 3183
rect 5240 3439 5298 3451
rect 5240 3183 5252 3439
rect 5286 3183 5298 3439
rect 5240 3171 5298 3183
rect 5418 3439 5476 3451
rect 5418 3183 5430 3439
rect 5464 3183 5476 3439
rect 5418 3171 5476 3183
rect 5596 3439 5654 3451
rect 5596 3183 5608 3439
rect 5642 3183 5654 3439
rect 5596 3171 5654 3183
rect 5774 3439 5832 3451
rect 5774 3183 5786 3439
rect 5820 3183 5832 3439
rect 5774 3171 5832 3183
rect 5952 3439 6010 3451
rect 5952 3183 5964 3439
rect 5998 3183 6010 3439
rect 5952 3171 6010 3183
rect 6130 3439 6188 3451
rect 6130 3183 6142 3439
rect 6176 3183 6188 3439
rect 6130 3171 6188 3183
rect 6308 3439 6366 3451
rect 6308 3183 6320 3439
rect 6354 3183 6366 3439
rect 6308 3171 6366 3183
rect 6486 3439 6544 3451
rect 6486 3183 6498 3439
rect 6532 3183 6544 3439
rect 6486 3171 6544 3183
rect 6664 3439 6722 3451
rect 6664 3183 6676 3439
rect 6710 3183 6722 3439
rect 6664 3171 6722 3183
rect 6842 3439 6900 3451
rect 6842 3183 6854 3439
rect 6888 3183 6900 3439
rect 6842 3171 6900 3183
rect 7020 3439 7078 3451
rect 7020 3183 7032 3439
rect 7066 3183 7078 3439
rect 7545 3383 7557 3639
rect 7591 3383 7603 3639
rect 7545 3371 7603 3383
rect 7723 3639 7781 3651
rect 7723 3383 7735 3639
rect 7769 3383 7781 3639
rect 7723 3371 7781 3383
rect 7901 3639 7959 3651
rect 7901 3383 7913 3639
rect 7947 3383 7959 3639
rect 7901 3371 7959 3383
rect 8079 3639 8137 3651
rect 8079 3383 8091 3639
rect 8125 3383 8137 3639
rect 8079 3371 8137 3383
rect 8257 3639 8315 3651
rect 8257 3383 8269 3639
rect 8303 3383 8315 3639
rect 8257 3371 8315 3383
rect 8435 3639 8493 3651
rect 8435 3383 8447 3639
rect 8481 3383 8493 3639
rect 8435 3371 8493 3383
rect 8613 3639 8671 3651
rect 8613 3383 8625 3639
rect 8659 3383 8671 3639
rect 8613 3371 8671 3383
rect 8791 3639 8849 3651
rect 8791 3383 8803 3639
rect 8837 3383 8849 3639
rect 8791 3371 8849 3383
rect 8969 3639 9027 3651
rect 8969 3383 8981 3639
rect 9015 3383 9027 3639
rect 8969 3371 9027 3383
rect 9147 3639 9205 3651
rect 9147 3383 9159 3639
rect 9193 3383 9205 3639
rect 9147 3371 9205 3383
rect 9325 3639 9383 3651
rect 9325 3383 9337 3639
rect 9371 3383 9383 3639
rect 9325 3371 9383 3383
rect 9503 3639 9561 3651
rect 9503 3383 9515 3639
rect 9549 3383 9561 3639
rect 9503 3371 9561 3383
rect 9681 3639 9739 3651
rect 9681 3383 9693 3639
rect 9727 3383 9739 3639
rect 9681 3371 9739 3383
rect 9859 3639 9917 3651
rect 9859 3383 9871 3639
rect 9905 3383 9917 3639
rect 9859 3371 9917 3383
rect 10037 3639 10095 3651
rect 10037 3383 10049 3639
rect 10083 3383 10095 3639
rect 10037 3371 10095 3383
rect 10232 3639 10290 3651
rect 10232 3383 10244 3639
rect 10278 3383 10290 3639
rect 10232 3371 10290 3383
rect 10410 3639 10468 3651
rect 10410 3383 10422 3639
rect 10456 3383 10468 3639
rect 10410 3371 10468 3383
rect 10588 3639 10646 3651
rect 10588 3383 10600 3639
rect 10634 3383 10646 3639
rect 10588 3371 10646 3383
rect 10766 3639 10824 3651
rect 10766 3383 10778 3639
rect 10812 3383 10824 3639
rect 10766 3371 10824 3383
rect 10944 3639 11002 3651
rect 10944 3383 10956 3639
rect 10990 3383 11002 3639
rect 10944 3371 11002 3383
rect 11122 3639 11180 3651
rect 11122 3383 11134 3639
rect 11168 3383 11180 3639
rect 11122 3371 11180 3383
rect 11300 3639 11358 3651
rect 11300 3383 11312 3639
rect 11346 3383 11358 3639
rect 11300 3371 11358 3383
rect 11478 3639 11536 3651
rect 11478 3383 11490 3639
rect 11524 3383 11536 3639
rect 11478 3371 11536 3383
rect 11656 3639 11714 3651
rect 11656 3383 11668 3639
rect 11702 3383 11714 3639
rect 11656 3371 11714 3383
rect 11834 3639 11892 3651
rect 11834 3383 11846 3639
rect 11880 3383 11892 3639
rect 11834 3371 11892 3383
rect 12012 3639 12070 3651
rect 12012 3383 12024 3639
rect 12058 3383 12070 3639
rect 12012 3371 12070 3383
rect 12190 3639 12248 3651
rect 12190 3383 12202 3639
rect 12236 3383 12248 3639
rect 12190 3371 12248 3383
rect 12368 3639 12426 3651
rect 12368 3383 12380 3639
rect 12414 3383 12426 3639
rect 12368 3371 12426 3383
rect 12546 3639 12604 3651
rect 12546 3383 12558 3639
rect 12592 3383 12604 3639
rect 12546 3371 12604 3383
rect 12724 3639 12782 3651
rect 12724 3383 12736 3639
rect 12770 3383 12782 3639
rect 12724 3371 12782 3383
rect 7020 3171 7078 3183
rect 7545 3139 7603 3151
rect 416 2939 474 2951
rect 416 2683 428 2939
rect 462 2683 474 2939
rect 416 2671 474 2683
rect 594 2939 652 2951
rect 594 2683 606 2939
rect 640 2683 652 2939
rect 594 2671 652 2683
rect 772 2939 830 2951
rect 772 2683 784 2939
rect 818 2683 830 2939
rect 772 2671 830 2683
rect 950 2939 1008 2951
rect 950 2683 962 2939
rect 996 2683 1008 2939
rect 950 2671 1008 2683
rect 1128 2939 1186 2951
rect 1128 2683 1140 2939
rect 1174 2683 1186 2939
rect 1128 2671 1186 2683
rect 1306 2939 1364 2951
rect 1306 2683 1318 2939
rect 1352 2683 1364 2939
rect 1306 2671 1364 2683
rect 1484 2939 1542 2951
rect 1484 2683 1496 2939
rect 1530 2683 1542 2939
rect 1484 2671 1542 2683
rect 1662 2939 1720 2951
rect 1662 2683 1674 2939
rect 1708 2683 1720 2939
rect 1662 2671 1720 2683
rect 1840 2939 1898 2951
rect 1840 2683 1852 2939
rect 1886 2683 1898 2939
rect 1840 2671 1898 2683
rect 2018 2939 2076 2951
rect 2018 2683 2030 2939
rect 2064 2683 2076 2939
rect 2018 2671 2076 2683
rect 2196 2939 2254 2951
rect 2196 2683 2208 2939
rect 2242 2683 2254 2939
rect 2196 2671 2254 2683
rect 2374 2939 2432 2951
rect 2374 2683 2386 2939
rect 2420 2683 2432 2939
rect 2374 2671 2432 2683
rect 2552 2939 2610 2951
rect 2552 2683 2564 2939
rect 2598 2683 2610 2939
rect 2552 2671 2610 2683
rect 2730 2939 2788 2951
rect 2730 2683 2742 2939
rect 2776 2683 2788 2939
rect 2730 2671 2788 2683
rect 2908 2939 2966 2951
rect 2908 2683 2920 2939
rect 2954 2683 2966 2939
rect 2908 2671 2966 2683
rect 3086 2939 3144 2951
rect 3086 2683 3098 2939
rect 3132 2683 3144 2939
rect 3086 2671 3144 2683
rect 3264 2939 3322 2951
rect 3264 2683 3276 2939
rect 3310 2683 3322 2939
rect 3264 2671 3322 2683
rect 3442 2939 3500 2951
rect 3442 2683 3454 2939
rect 3488 2683 3500 2939
rect 3442 2671 3500 2683
rect 3620 2939 3678 2951
rect 3620 2683 3632 2939
rect 3666 2683 3678 2939
rect 3620 2671 3678 2683
rect 3816 2939 3874 2951
rect 3816 2683 3828 2939
rect 3862 2683 3874 2939
rect 3816 2671 3874 2683
rect 3994 2939 4052 2951
rect 3994 2683 4006 2939
rect 4040 2683 4052 2939
rect 3994 2671 4052 2683
rect 4172 2939 4230 2951
rect 4172 2683 4184 2939
rect 4218 2683 4230 2939
rect 4172 2671 4230 2683
rect 4350 2939 4408 2951
rect 4350 2683 4362 2939
rect 4396 2683 4408 2939
rect 4350 2671 4408 2683
rect 4528 2939 4586 2951
rect 4528 2683 4540 2939
rect 4574 2683 4586 2939
rect 4528 2671 4586 2683
rect 4706 2939 4764 2951
rect 4706 2683 4718 2939
rect 4752 2683 4764 2939
rect 4706 2671 4764 2683
rect 4884 2939 4942 2951
rect 4884 2683 4896 2939
rect 4930 2683 4942 2939
rect 4884 2671 4942 2683
rect 5062 2939 5120 2951
rect 5062 2683 5074 2939
rect 5108 2683 5120 2939
rect 5062 2671 5120 2683
rect 5240 2939 5298 2951
rect 5240 2683 5252 2939
rect 5286 2683 5298 2939
rect 5240 2671 5298 2683
rect 5418 2939 5476 2951
rect 5418 2683 5430 2939
rect 5464 2683 5476 2939
rect 5418 2671 5476 2683
rect 5596 2939 5654 2951
rect 5596 2683 5608 2939
rect 5642 2683 5654 2939
rect 5596 2671 5654 2683
rect 5774 2939 5832 2951
rect 5774 2683 5786 2939
rect 5820 2683 5832 2939
rect 5774 2671 5832 2683
rect 5952 2939 6010 2951
rect 5952 2683 5964 2939
rect 5998 2683 6010 2939
rect 5952 2671 6010 2683
rect 6130 2939 6188 2951
rect 6130 2683 6142 2939
rect 6176 2683 6188 2939
rect 6130 2671 6188 2683
rect 6308 2939 6366 2951
rect 6308 2683 6320 2939
rect 6354 2683 6366 2939
rect 6308 2671 6366 2683
rect 6486 2939 6544 2951
rect 6486 2683 6498 2939
rect 6532 2683 6544 2939
rect 6486 2671 6544 2683
rect 6664 2939 6722 2951
rect 6664 2683 6676 2939
rect 6710 2683 6722 2939
rect 6664 2671 6722 2683
rect 6842 2939 6900 2951
rect 6842 2683 6854 2939
rect 6888 2683 6900 2939
rect 6842 2671 6900 2683
rect 7020 2939 7078 2951
rect 7020 2683 7032 2939
rect 7066 2683 7078 2939
rect 7545 2883 7557 3139
rect 7591 2883 7603 3139
rect 7545 2871 7603 2883
rect 7723 3139 7781 3151
rect 7723 2883 7735 3139
rect 7769 2883 7781 3139
rect 7723 2871 7781 2883
rect 7901 3139 7959 3151
rect 7901 2883 7913 3139
rect 7947 2883 7959 3139
rect 7901 2871 7959 2883
rect 8079 3139 8137 3151
rect 8079 2883 8091 3139
rect 8125 2883 8137 3139
rect 8079 2871 8137 2883
rect 8257 3139 8315 3151
rect 8257 2883 8269 3139
rect 8303 2883 8315 3139
rect 8257 2871 8315 2883
rect 8435 3139 8493 3151
rect 8435 2883 8447 3139
rect 8481 2883 8493 3139
rect 8435 2871 8493 2883
rect 8613 3139 8671 3151
rect 8613 2883 8625 3139
rect 8659 2883 8671 3139
rect 8613 2871 8671 2883
rect 8791 3139 8849 3151
rect 8791 2883 8803 3139
rect 8837 2883 8849 3139
rect 8791 2871 8849 2883
rect 8969 3139 9027 3151
rect 8969 2883 8981 3139
rect 9015 2883 9027 3139
rect 8969 2871 9027 2883
rect 9147 3139 9205 3151
rect 9147 2883 9159 3139
rect 9193 2883 9205 3139
rect 9147 2871 9205 2883
rect 9325 3139 9383 3151
rect 9325 2883 9337 3139
rect 9371 2883 9383 3139
rect 9325 2871 9383 2883
rect 9503 3139 9561 3151
rect 9503 2883 9515 3139
rect 9549 2883 9561 3139
rect 9503 2871 9561 2883
rect 9681 3139 9739 3151
rect 9681 2883 9693 3139
rect 9727 2883 9739 3139
rect 9681 2871 9739 2883
rect 9859 3139 9917 3151
rect 9859 2883 9871 3139
rect 9905 2883 9917 3139
rect 9859 2871 9917 2883
rect 10037 3139 10095 3151
rect 10037 2883 10049 3139
rect 10083 2883 10095 3139
rect 10037 2871 10095 2883
rect 10232 3139 10290 3151
rect 10232 2883 10244 3139
rect 10278 2883 10290 3139
rect 10232 2871 10290 2883
rect 10410 3139 10468 3151
rect 10410 2883 10422 3139
rect 10456 2883 10468 3139
rect 10410 2871 10468 2883
rect 10588 3139 10646 3151
rect 10588 2883 10600 3139
rect 10634 2883 10646 3139
rect 10588 2871 10646 2883
rect 10766 3139 10824 3151
rect 10766 2883 10778 3139
rect 10812 2883 10824 3139
rect 10766 2871 10824 2883
rect 10944 3139 11002 3151
rect 10944 2883 10956 3139
rect 10990 2883 11002 3139
rect 10944 2871 11002 2883
rect 11122 3139 11180 3151
rect 11122 2883 11134 3139
rect 11168 2883 11180 3139
rect 11122 2871 11180 2883
rect 11300 3139 11358 3151
rect 11300 2883 11312 3139
rect 11346 2883 11358 3139
rect 11300 2871 11358 2883
rect 11478 3139 11536 3151
rect 11478 2883 11490 3139
rect 11524 2883 11536 3139
rect 11478 2871 11536 2883
rect 11656 3139 11714 3151
rect 11656 2883 11668 3139
rect 11702 2883 11714 3139
rect 11656 2871 11714 2883
rect 11834 3139 11892 3151
rect 11834 2883 11846 3139
rect 11880 2883 11892 3139
rect 11834 2871 11892 2883
rect 12012 3139 12070 3151
rect 12012 2883 12024 3139
rect 12058 2883 12070 3139
rect 12012 2871 12070 2883
rect 12190 3139 12248 3151
rect 12190 2883 12202 3139
rect 12236 2883 12248 3139
rect 12190 2871 12248 2883
rect 12368 3139 12426 3151
rect 12368 2883 12380 3139
rect 12414 2883 12426 3139
rect 12368 2871 12426 2883
rect 12546 3139 12604 3151
rect 12546 2883 12558 3139
rect 12592 2883 12604 3139
rect 12546 2871 12604 2883
rect 12724 3139 12782 3151
rect 12724 2883 12736 3139
rect 12770 2883 12782 3139
rect 12724 2871 12782 2883
rect 7020 2671 7078 2683
rect 7545 2639 7603 2651
rect 416 2439 474 2451
rect 416 2183 428 2439
rect 462 2183 474 2439
rect 416 2171 474 2183
rect 594 2439 652 2451
rect 594 2183 606 2439
rect 640 2183 652 2439
rect 594 2171 652 2183
rect 772 2439 830 2451
rect 772 2183 784 2439
rect 818 2183 830 2439
rect 772 2171 830 2183
rect 950 2439 1008 2451
rect 950 2183 962 2439
rect 996 2183 1008 2439
rect 950 2171 1008 2183
rect 1128 2439 1186 2451
rect 1128 2183 1140 2439
rect 1174 2183 1186 2439
rect 1128 2171 1186 2183
rect 1306 2439 1364 2451
rect 1306 2183 1318 2439
rect 1352 2183 1364 2439
rect 1306 2171 1364 2183
rect 1484 2439 1542 2451
rect 1484 2183 1496 2439
rect 1530 2183 1542 2439
rect 1484 2171 1542 2183
rect 1662 2439 1720 2451
rect 1662 2183 1674 2439
rect 1708 2183 1720 2439
rect 1662 2171 1720 2183
rect 1840 2439 1898 2451
rect 1840 2183 1852 2439
rect 1886 2183 1898 2439
rect 1840 2171 1898 2183
rect 2018 2439 2076 2451
rect 2018 2183 2030 2439
rect 2064 2183 2076 2439
rect 2018 2171 2076 2183
rect 2196 2439 2254 2451
rect 2196 2183 2208 2439
rect 2242 2183 2254 2439
rect 2196 2171 2254 2183
rect 2374 2439 2432 2451
rect 2374 2183 2386 2439
rect 2420 2183 2432 2439
rect 2374 2171 2432 2183
rect 2552 2439 2610 2451
rect 2552 2183 2564 2439
rect 2598 2183 2610 2439
rect 2552 2171 2610 2183
rect 2730 2439 2788 2451
rect 2730 2183 2742 2439
rect 2776 2183 2788 2439
rect 2730 2171 2788 2183
rect 2908 2439 2966 2451
rect 2908 2183 2920 2439
rect 2954 2183 2966 2439
rect 2908 2171 2966 2183
rect 3086 2439 3144 2451
rect 3086 2183 3098 2439
rect 3132 2183 3144 2439
rect 3086 2171 3144 2183
rect 3264 2439 3322 2451
rect 3264 2183 3276 2439
rect 3310 2183 3322 2439
rect 3264 2171 3322 2183
rect 3442 2439 3500 2451
rect 3442 2183 3454 2439
rect 3488 2183 3500 2439
rect 3442 2171 3500 2183
rect 3620 2439 3678 2451
rect 3620 2183 3632 2439
rect 3666 2183 3678 2439
rect 3620 2171 3678 2183
rect 3816 2439 3874 2451
rect 3816 2183 3828 2439
rect 3862 2183 3874 2439
rect 3816 2171 3874 2183
rect 3994 2439 4052 2451
rect 3994 2183 4006 2439
rect 4040 2183 4052 2439
rect 3994 2171 4052 2183
rect 4172 2439 4230 2451
rect 4172 2183 4184 2439
rect 4218 2183 4230 2439
rect 4172 2171 4230 2183
rect 4350 2439 4408 2451
rect 4350 2183 4362 2439
rect 4396 2183 4408 2439
rect 4350 2171 4408 2183
rect 4528 2439 4586 2451
rect 4528 2183 4540 2439
rect 4574 2183 4586 2439
rect 4528 2171 4586 2183
rect 4706 2439 4764 2451
rect 4706 2183 4718 2439
rect 4752 2183 4764 2439
rect 4706 2171 4764 2183
rect 4884 2439 4942 2451
rect 4884 2183 4896 2439
rect 4930 2183 4942 2439
rect 4884 2171 4942 2183
rect 5062 2439 5120 2451
rect 5062 2183 5074 2439
rect 5108 2183 5120 2439
rect 5062 2171 5120 2183
rect 5240 2439 5298 2451
rect 5240 2183 5252 2439
rect 5286 2183 5298 2439
rect 5240 2171 5298 2183
rect 5418 2439 5476 2451
rect 5418 2183 5430 2439
rect 5464 2183 5476 2439
rect 5418 2171 5476 2183
rect 5596 2439 5654 2451
rect 5596 2183 5608 2439
rect 5642 2183 5654 2439
rect 5596 2171 5654 2183
rect 5774 2439 5832 2451
rect 5774 2183 5786 2439
rect 5820 2183 5832 2439
rect 5774 2171 5832 2183
rect 5952 2439 6010 2451
rect 5952 2183 5964 2439
rect 5998 2183 6010 2439
rect 5952 2171 6010 2183
rect 6130 2439 6188 2451
rect 6130 2183 6142 2439
rect 6176 2183 6188 2439
rect 6130 2171 6188 2183
rect 6308 2439 6366 2451
rect 6308 2183 6320 2439
rect 6354 2183 6366 2439
rect 6308 2171 6366 2183
rect 6486 2439 6544 2451
rect 6486 2183 6498 2439
rect 6532 2183 6544 2439
rect 6486 2171 6544 2183
rect 6664 2439 6722 2451
rect 6664 2183 6676 2439
rect 6710 2183 6722 2439
rect 6664 2171 6722 2183
rect 6842 2439 6900 2451
rect 6842 2183 6854 2439
rect 6888 2183 6900 2439
rect 6842 2171 6900 2183
rect 7020 2439 7078 2451
rect 7020 2183 7032 2439
rect 7066 2183 7078 2439
rect 7545 2383 7557 2639
rect 7591 2383 7603 2639
rect 7545 2371 7603 2383
rect 7723 2639 7781 2651
rect 7723 2383 7735 2639
rect 7769 2383 7781 2639
rect 7723 2371 7781 2383
rect 7901 2639 7959 2651
rect 7901 2383 7913 2639
rect 7947 2383 7959 2639
rect 7901 2371 7959 2383
rect 8079 2639 8137 2651
rect 8079 2383 8091 2639
rect 8125 2383 8137 2639
rect 8079 2371 8137 2383
rect 8257 2639 8315 2651
rect 8257 2383 8269 2639
rect 8303 2383 8315 2639
rect 8257 2371 8315 2383
rect 8435 2639 8493 2651
rect 8435 2383 8447 2639
rect 8481 2383 8493 2639
rect 8435 2371 8493 2383
rect 8613 2639 8671 2651
rect 8613 2383 8625 2639
rect 8659 2383 8671 2639
rect 8613 2371 8671 2383
rect 8791 2639 8849 2651
rect 8791 2383 8803 2639
rect 8837 2383 8849 2639
rect 8791 2371 8849 2383
rect 8969 2639 9027 2651
rect 8969 2383 8981 2639
rect 9015 2383 9027 2639
rect 8969 2371 9027 2383
rect 9147 2639 9205 2651
rect 9147 2383 9159 2639
rect 9193 2383 9205 2639
rect 9147 2371 9205 2383
rect 9325 2639 9383 2651
rect 9325 2383 9337 2639
rect 9371 2383 9383 2639
rect 9325 2371 9383 2383
rect 9503 2639 9561 2651
rect 9503 2383 9515 2639
rect 9549 2383 9561 2639
rect 9503 2371 9561 2383
rect 9681 2639 9739 2651
rect 9681 2383 9693 2639
rect 9727 2383 9739 2639
rect 9681 2371 9739 2383
rect 9859 2639 9917 2651
rect 9859 2383 9871 2639
rect 9905 2383 9917 2639
rect 9859 2371 9917 2383
rect 10037 2639 10095 2651
rect 10037 2383 10049 2639
rect 10083 2383 10095 2639
rect 10037 2371 10095 2383
rect 10232 2639 10290 2651
rect 10232 2383 10244 2639
rect 10278 2383 10290 2639
rect 10232 2371 10290 2383
rect 10410 2639 10468 2651
rect 10410 2383 10422 2639
rect 10456 2383 10468 2639
rect 10410 2371 10468 2383
rect 10588 2639 10646 2651
rect 10588 2383 10600 2639
rect 10634 2383 10646 2639
rect 10588 2371 10646 2383
rect 10766 2639 10824 2651
rect 10766 2383 10778 2639
rect 10812 2383 10824 2639
rect 10766 2371 10824 2383
rect 10944 2639 11002 2651
rect 10944 2383 10956 2639
rect 10990 2383 11002 2639
rect 10944 2371 11002 2383
rect 11122 2639 11180 2651
rect 11122 2383 11134 2639
rect 11168 2383 11180 2639
rect 11122 2371 11180 2383
rect 11300 2639 11358 2651
rect 11300 2383 11312 2639
rect 11346 2383 11358 2639
rect 11300 2371 11358 2383
rect 11478 2639 11536 2651
rect 11478 2383 11490 2639
rect 11524 2383 11536 2639
rect 11478 2371 11536 2383
rect 11656 2639 11714 2651
rect 11656 2383 11668 2639
rect 11702 2383 11714 2639
rect 11656 2371 11714 2383
rect 11834 2639 11892 2651
rect 11834 2383 11846 2639
rect 11880 2383 11892 2639
rect 11834 2371 11892 2383
rect 12012 2639 12070 2651
rect 12012 2383 12024 2639
rect 12058 2383 12070 2639
rect 12012 2371 12070 2383
rect 12190 2639 12248 2651
rect 12190 2383 12202 2639
rect 12236 2383 12248 2639
rect 12190 2371 12248 2383
rect 12368 2639 12426 2651
rect 12368 2383 12380 2639
rect 12414 2383 12426 2639
rect 12368 2371 12426 2383
rect 12546 2639 12604 2651
rect 12546 2383 12558 2639
rect 12592 2383 12604 2639
rect 12546 2371 12604 2383
rect 12724 2639 12782 2651
rect 12724 2383 12736 2639
rect 12770 2383 12782 2639
rect 12724 2371 12782 2383
rect 7020 2171 7078 2183
rect 416 1939 474 1951
rect 416 1683 428 1939
rect 462 1683 474 1939
rect 416 1671 474 1683
rect 594 1939 652 1951
rect 594 1683 606 1939
rect 640 1683 652 1939
rect 594 1671 652 1683
rect 772 1939 830 1951
rect 772 1683 784 1939
rect 818 1683 830 1939
rect 772 1671 830 1683
rect 950 1939 1008 1951
rect 950 1683 962 1939
rect 996 1683 1008 1939
rect 950 1671 1008 1683
rect 1128 1939 1186 1951
rect 1128 1683 1140 1939
rect 1174 1683 1186 1939
rect 1128 1671 1186 1683
rect 1306 1939 1364 1951
rect 1306 1683 1318 1939
rect 1352 1683 1364 1939
rect 1306 1671 1364 1683
rect 1484 1939 1542 1951
rect 1484 1683 1496 1939
rect 1530 1683 1542 1939
rect 1484 1671 1542 1683
rect 1662 1939 1720 1951
rect 1662 1683 1674 1939
rect 1708 1683 1720 1939
rect 1662 1671 1720 1683
rect 1840 1939 1898 1951
rect 1840 1683 1852 1939
rect 1886 1683 1898 1939
rect 1840 1671 1898 1683
rect 2018 1939 2076 1951
rect 2018 1683 2030 1939
rect 2064 1683 2076 1939
rect 2018 1671 2076 1683
rect 2196 1939 2254 1951
rect 2196 1683 2208 1939
rect 2242 1683 2254 1939
rect 2196 1671 2254 1683
rect 2374 1939 2432 1951
rect 2374 1683 2386 1939
rect 2420 1683 2432 1939
rect 2374 1671 2432 1683
rect 2552 1939 2610 1951
rect 2552 1683 2564 1939
rect 2598 1683 2610 1939
rect 2552 1671 2610 1683
rect 2730 1939 2788 1951
rect 2730 1683 2742 1939
rect 2776 1683 2788 1939
rect 2730 1671 2788 1683
rect 2908 1939 2966 1951
rect 2908 1683 2920 1939
rect 2954 1683 2966 1939
rect 2908 1671 2966 1683
rect 3086 1939 3144 1951
rect 3086 1683 3098 1939
rect 3132 1683 3144 1939
rect 3086 1671 3144 1683
rect 3264 1939 3322 1951
rect 3264 1683 3276 1939
rect 3310 1683 3322 1939
rect 3264 1671 3322 1683
rect 3442 1939 3500 1951
rect 3442 1683 3454 1939
rect 3488 1683 3500 1939
rect 3442 1671 3500 1683
rect 3620 1939 3678 1951
rect 3620 1683 3632 1939
rect 3666 1683 3678 1939
rect 3620 1671 3678 1683
rect 3816 1939 3874 1951
rect 3816 1683 3828 1939
rect 3862 1683 3874 1939
rect 3816 1671 3874 1683
rect 3994 1939 4052 1951
rect 3994 1683 4006 1939
rect 4040 1683 4052 1939
rect 3994 1671 4052 1683
rect 4172 1939 4230 1951
rect 4172 1683 4184 1939
rect 4218 1683 4230 1939
rect 4172 1671 4230 1683
rect 4350 1939 4408 1951
rect 4350 1683 4362 1939
rect 4396 1683 4408 1939
rect 4350 1671 4408 1683
rect 4528 1939 4586 1951
rect 4528 1683 4540 1939
rect 4574 1683 4586 1939
rect 4528 1671 4586 1683
rect 4706 1939 4764 1951
rect 4706 1683 4718 1939
rect 4752 1683 4764 1939
rect 4706 1671 4764 1683
rect 4884 1939 4942 1951
rect 4884 1683 4896 1939
rect 4930 1683 4942 1939
rect 4884 1671 4942 1683
rect 5062 1939 5120 1951
rect 5062 1683 5074 1939
rect 5108 1683 5120 1939
rect 5062 1671 5120 1683
rect 5240 1939 5298 1951
rect 5240 1683 5252 1939
rect 5286 1683 5298 1939
rect 5240 1671 5298 1683
rect 5418 1939 5476 1951
rect 5418 1683 5430 1939
rect 5464 1683 5476 1939
rect 5418 1671 5476 1683
rect 5596 1939 5654 1951
rect 5596 1683 5608 1939
rect 5642 1683 5654 1939
rect 5596 1671 5654 1683
rect 5774 1939 5832 1951
rect 5774 1683 5786 1939
rect 5820 1683 5832 1939
rect 5774 1671 5832 1683
rect 5952 1939 6010 1951
rect 5952 1683 5964 1939
rect 5998 1683 6010 1939
rect 5952 1671 6010 1683
rect 6130 1939 6188 1951
rect 6130 1683 6142 1939
rect 6176 1683 6188 1939
rect 6130 1671 6188 1683
rect 6308 1939 6366 1951
rect 6308 1683 6320 1939
rect 6354 1683 6366 1939
rect 6308 1671 6366 1683
rect 6486 1939 6544 1951
rect 6486 1683 6498 1939
rect 6532 1683 6544 1939
rect 6486 1671 6544 1683
rect 6664 1939 6722 1951
rect 6664 1683 6676 1939
rect 6710 1683 6722 1939
rect 6664 1671 6722 1683
rect 6842 1939 6900 1951
rect 6842 1683 6854 1939
rect 6888 1683 6900 1939
rect 6842 1671 6900 1683
rect 7020 1939 7078 1951
rect 7020 1683 7032 1939
rect 7066 1683 7078 1939
rect 7020 1671 7078 1683
rect 7545 1939 7603 1951
rect 7545 1683 7557 1939
rect 7591 1683 7603 1939
rect 7545 1671 7603 1683
rect 7723 1939 7781 1951
rect 7723 1683 7735 1939
rect 7769 1683 7781 1939
rect 7723 1671 7781 1683
rect 7901 1939 7959 1951
rect 7901 1683 7913 1939
rect 7947 1683 7959 1939
rect 7901 1671 7959 1683
rect 8079 1939 8137 1951
rect 8079 1683 8091 1939
rect 8125 1683 8137 1939
rect 8079 1671 8137 1683
rect 8257 1939 8315 1951
rect 8257 1683 8269 1939
rect 8303 1683 8315 1939
rect 8257 1671 8315 1683
rect 8435 1939 8493 1951
rect 8435 1683 8447 1939
rect 8481 1683 8493 1939
rect 8435 1671 8493 1683
rect 8613 1939 8671 1951
rect 8613 1683 8625 1939
rect 8659 1683 8671 1939
rect 8613 1671 8671 1683
rect 8791 1939 8849 1951
rect 8791 1683 8803 1939
rect 8837 1683 8849 1939
rect 8791 1671 8849 1683
rect 8969 1939 9027 1951
rect 8969 1683 8981 1939
rect 9015 1683 9027 1939
rect 8969 1671 9027 1683
rect 9147 1939 9205 1951
rect 9147 1683 9159 1939
rect 9193 1683 9205 1939
rect 9147 1671 9205 1683
rect 9325 1939 9383 1951
rect 9325 1683 9337 1939
rect 9371 1683 9383 1939
rect 9325 1671 9383 1683
rect 9503 1939 9561 1951
rect 9503 1683 9515 1939
rect 9549 1683 9561 1939
rect 9503 1671 9561 1683
rect 9681 1939 9739 1951
rect 9681 1683 9693 1939
rect 9727 1683 9739 1939
rect 9681 1671 9739 1683
rect 9859 1939 9917 1951
rect 9859 1683 9871 1939
rect 9905 1683 9917 1939
rect 9859 1671 9917 1683
rect 10037 1939 10095 1951
rect 10037 1683 10049 1939
rect 10083 1683 10095 1939
rect 10037 1671 10095 1683
rect 10232 1939 10290 1951
rect 10232 1683 10244 1939
rect 10278 1683 10290 1939
rect 10232 1671 10290 1683
rect 10410 1939 10468 1951
rect 10410 1683 10422 1939
rect 10456 1683 10468 1939
rect 10410 1671 10468 1683
rect 10588 1939 10646 1951
rect 10588 1683 10600 1939
rect 10634 1683 10646 1939
rect 10588 1671 10646 1683
rect 10766 1939 10824 1951
rect 10766 1683 10778 1939
rect 10812 1683 10824 1939
rect 10766 1671 10824 1683
rect 10944 1939 11002 1951
rect 10944 1683 10956 1939
rect 10990 1683 11002 1939
rect 10944 1671 11002 1683
rect 11122 1939 11180 1951
rect 11122 1683 11134 1939
rect 11168 1683 11180 1939
rect 11122 1671 11180 1683
rect 11300 1939 11358 1951
rect 11300 1683 11312 1939
rect 11346 1683 11358 1939
rect 11300 1671 11358 1683
rect 11478 1939 11536 1951
rect 11478 1683 11490 1939
rect 11524 1683 11536 1939
rect 11478 1671 11536 1683
rect 11656 1939 11714 1951
rect 11656 1683 11668 1939
rect 11702 1683 11714 1939
rect 11656 1671 11714 1683
rect 11834 1939 11892 1951
rect 11834 1683 11846 1939
rect 11880 1683 11892 1939
rect 11834 1671 11892 1683
rect 12012 1939 12070 1951
rect 12012 1683 12024 1939
rect 12058 1683 12070 1939
rect 12012 1671 12070 1683
rect 12190 1939 12248 1951
rect 12190 1683 12202 1939
rect 12236 1683 12248 1939
rect 12190 1671 12248 1683
rect 12368 1939 12426 1951
rect 12368 1683 12380 1939
rect 12414 1683 12426 1939
rect 12368 1671 12426 1683
rect 12546 1939 12604 1951
rect 12546 1683 12558 1939
rect 12592 1683 12604 1939
rect 12546 1671 12604 1683
rect 12724 1939 12782 1951
rect 12724 1683 12736 1939
rect 12770 1683 12782 1939
rect 12724 1671 12782 1683
rect 416 1439 474 1451
rect 416 1183 428 1439
rect 462 1183 474 1439
rect 416 1171 474 1183
rect 594 1439 652 1451
rect 594 1183 606 1439
rect 640 1183 652 1439
rect 594 1171 652 1183
rect 772 1439 830 1451
rect 772 1183 784 1439
rect 818 1183 830 1439
rect 772 1171 830 1183
rect 950 1439 1008 1451
rect 950 1183 962 1439
rect 996 1183 1008 1439
rect 950 1171 1008 1183
rect 1128 1439 1186 1451
rect 1128 1183 1140 1439
rect 1174 1183 1186 1439
rect 1128 1171 1186 1183
rect 1306 1439 1364 1451
rect 1306 1183 1318 1439
rect 1352 1183 1364 1439
rect 1306 1171 1364 1183
rect 1484 1439 1542 1451
rect 1484 1183 1496 1439
rect 1530 1183 1542 1439
rect 1484 1171 1542 1183
rect 1662 1439 1720 1451
rect 1662 1183 1674 1439
rect 1708 1183 1720 1439
rect 1662 1171 1720 1183
rect 1840 1439 1898 1451
rect 1840 1183 1852 1439
rect 1886 1183 1898 1439
rect 1840 1171 1898 1183
rect 2018 1439 2076 1451
rect 2018 1183 2030 1439
rect 2064 1183 2076 1439
rect 2018 1171 2076 1183
rect 2196 1439 2254 1451
rect 2196 1183 2208 1439
rect 2242 1183 2254 1439
rect 2196 1171 2254 1183
rect 2374 1439 2432 1451
rect 2374 1183 2386 1439
rect 2420 1183 2432 1439
rect 2374 1171 2432 1183
rect 2552 1439 2610 1451
rect 2552 1183 2564 1439
rect 2598 1183 2610 1439
rect 2552 1171 2610 1183
rect 2730 1439 2788 1451
rect 2730 1183 2742 1439
rect 2776 1183 2788 1439
rect 2730 1171 2788 1183
rect 2908 1439 2966 1451
rect 2908 1183 2920 1439
rect 2954 1183 2966 1439
rect 2908 1171 2966 1183
rect 3086 1439 3144 1451
rect 3086 1183 3098 1439
rect 3132 1183 3144 1439
rect 3086 1171 3144 1183
rect 3264 1439 3322 1451
rect 3264 1183 3276 1439
rect 3310 1183 3322 1439
rect 3264 1171 3322 1183
rect 3442 1439 3500 1451
rect 3442 1183 3454 1439
rect 3488 1183 3500 1439
rect 3442 1171 3500 1183
rect 3620 1439 3678 1451
rect 3620 1183 3632 1439
rect 3666 1183 3678 1439
rect 3620 1171 3678 1183
rect 3816 1439 3874 1451
rect 3816 1183 3828 1439
rect 3862 1183 3874 1439
rect 3816 1171 3874 1183
rect 3994 1439 4052 1451
rect 3994 1183 4006 1439
rect 4040 1183 4052 1439
rect 3994 1171 4052 1183
rect 4172 1439 4230 1451
rect 4172 1183 4184 1439
rect 4218 1183 4230 1439
rect 4172 1171 4230 1183
rect 4350 1439 4408 1451
rect 4350 1183 4362 1439
rect 4396 1183 4408 1439
rect 4350 1171 4408 1183
rect 4528 1439 4586 1451
rect 4528 1183 4540 1439
rect 4574 1183 4586 1439
rect 4528 1171 4586 1183
rect 4706 1439 4764 1451
rect 4706 1183 4718 1439
rect 4752 1183 4764 1439
rect 4706 1171 4764 1183
rect 4884 1439 4942 1451
rect 4884 1183 4896 1439
rect 4930 1183 4942 1439
rect 4884 1171 4942 1183
rect 5062 1439 5120 1451
rect 5062 1183 5074 1439
rect 5108 1183 5120 1439
rect 5062 1171 5120 1183
rect 5240 1439 5298 1451
rect 5240 1183 5252 1439
rect 5286 1183 5298 1439
rect 5240 1171 5298 1183
rect 5418 1439 5476 1451
rect 5418 1183 5430 1439
rect 5464 1183 5476 1439
rect 5418 1171 5476 1183
rect 5596 1439 5654 1451
rect 5596 1183 5608 1439
rect 5642 1183 5654 1439
rect 5596 1171 5654 1183
rect 5774 1439 5832 1451
rect 5774 1183 5786 1439
rect 5820 1183 5832 1439
rect 5774 1171 5832 1183
rect 5952 1439 6010 1451
rect 5952 1183 5964 1439
rect 5998 1183 6010 1439
rect 5952 1171 6010 1183
rect 6130 1439 6188 1451
rect 6130 1183 6142 1439
rect 6176 1183 6188 1439
rect 6130 1171 6188 1183
rect 6308 1439 6366 1451
rect 6308 1183 6320 1439
rect 6354 1183 6366 1439
rect 6308 1171 6366 1183
rect 6486 1439 6544 1451
rect 6486 1183 6498 1439
rect 6532 1183 6544 1439
rect 6486 1171 6544 1183
rect 6664 1439 6722 1451
rect 6664 1183 6676 1439
rect 6710 1183 6722 1439
rect 6664 1171 6722 1183
rect 6842 1439 6900 1451
rect 6842 1183 6854 1439
rect 6888 1183 6900 1439
rect 6842 1171 6900 1183
rect 7020 1439 7078 1451
rect 7020 1183 7032 1439
rect 7066 1183 7078 1439
rect 7020 1171 7078 1183
rect 7545 1439 7603 1451
rect 7545 1183 7557 1439
rect 7591 1183 7603 1439
rect 7545 1171 7603 1183
rect 7723 1439 7781 1451
rect 7723 1183 7735 1439
rect 7769 1183 7781 1439
rect 7723 1171 7781 1183
rect 7901 1439 7959 1451
rect 7901 1183 7913 1439
rect 7947 1183 7959 1439
rect 7901 1171 7959 1183
rect 8079 1439 8137 1451
rect 8079 1183 8091 1439
rect 8125 1183 8137 1439
rect 8079 1171 8137 1183
rect 8257 1439 8315 1451
rect 8257 1183 8269 1439
rect 8303 1183 8315 1439
rect 8257 1171 8315 1183
rect 8435 1439 8493 1451
rect 8435 1183 8447 1439
rect 8481 1183 8493 1439
rect 8435 1171 8493 1183
rect 8613 1439 8671 1451
rect 8613 1183 8625 1439
rect 8659 1183 8671 1439
rect 8613 1171 8671 1183
rect 8791 1439 8849 1451
rect 8791 1183 8803 1439
rect 8837 1183 8849 1439
rect 8791 1171 8849 1183
rect 8969 1439 9027 1451
rect 8969 1183 8981 1439
rect 9015 1183 9027 1439
rect 8969 1171 9027 1183
rect 9147 1439 9205 1451
rect 9147 1183 9159 1439
rect 9193 1183 9205 1439
rect 9147 1171 9205 1183
rect 9325 1439 9383 1451
rect 9325 1183 9337 1439
rect 9371 1183 9383 1439
rect 9325 1171 9383 1183
rect 9503 1439 9561 1451
rect 9503 1183 9515 1439
rect 9549 1183 9561 1439
rect 9503 1171 9561 1183
rect 9681 1439 9739 1451
rect 9681 1183 9693 1439
rect 9727 1183 9739 1439
rect 9681 1171 9739 1183
rect 9859 1439 9917 1451
rect 9859 1183 9871 1439
rect 9905 1183 9917 1439
rect 9859 1171 9917 1183
rect 10037 1439 10095 1451
rect 10037 1183 10049 1439
rect 10083 1183 10095 1439
rect 10037 1171 10095 1183
rect 10232 1439 10290 1451
rect 10232 1183 10244 1439
rect 10278 1183 10290 1439
rect 10232 1171 10290 1183
rect 10410 1439 10468 1451
rect 10410 1183 10422 1439
rect 10456 1183 10468 1439
rect 10410 1171 10468 1183
rect 10588 1439 10646 1451
rect 10588 1183 10600 1439
rect 10634 1183 10646 1439
rect 10588 1171 10646 1183
rect 10766 1439 10824 1451
rect 10766 1183 10778 1439
rect 10812 1183 10824 1439
rect 10766 1171 10824 1183
rect 10944 1439 11002 1451
rect 10944 1183 10956 1439
rect 10990 1183 11002 1439
rect 10944 1171 11002 1183
rect 11122 1439 11180 1451
rect 11122 1183 11134 1439
rect 11168 1183 11180 1439
rect 11122 1171 11180 1183
rect 11300 1439 11358 1451
rect 11300 1183 11312 1439
rect 11346 1183 11358 1439
rect 11300 1171 11358 1183
rect 11478 1439 11536 1451
rect 11478 1183 11490 1439
rect 11524 1183 11536 1439
rect 11478 1171 11536 1183
rect 11656 1439 11714 1451
rect 11656 1183 11668 1439
rect 11702 1183 11714 1439
rect 11656 1171 11714 1183
rect 11834 1439 11892 1451
rect 11834 1183 11846 1439
rect 11880 1183 11892 1439
rect 11834 1171 11892 1183
rect 12012 1439 12070 1451
rect 12012 1183 12024 1439
rect 12058 1183 12070 1439
rect 12012 1171 12070 1183
rect 12190 1439 12248 1451
rect 12190 1183 12202 1439
rect 12236 1183 12248 1439
rect 12190 1171 12248 1183
rect 12368 1439 12426 1451
rect 12368 1183 12380 1439
rect 12414 1183 12426 1439
rect 12368 1171 12426 1183
rect 12546 1439 12604 1451
rect 12546 1183 12558 1439
rect 12592 1183 12604 1439
rect 12546 1171 12604 1183
rect 12724 1439 12782 1451
rect 12724 1183 12736 1439
rect 12770 1183 12782 1439
rect 12724 1171 12782 1183
rect 416 939 474 951
rect 416 683 428 939
rect 462 683 474 939
rect 416 671 474 683
rect 594 939 652 951
rect 594 683 606 939
rect 640 683 652 939
rect 594 671 652 683
rect 772 939 830 951
rect 772 683 784 939
rect 818 683 830 939
rect 772 671 830 683
rect 950 939 1008 951
rect 950 683 962 939
rect 996 683 1008 939
rect 950 671 1008 683
rect 1128 939 1186 951
rect 1128 683 1140 939
rect 1174 683 1186 939
rect 1128 671 1186 683
rect 1306 939 1364 951
rect 1306 683 1318 939
rect 1352 683 1364 939
rect 1306 671 1364 683
rect 1484 939 1542 951
rect 1484 683 1496 939
rect 1530 683 1542 939
rect 1484 671 1542 683
rect 1662 939 1720 951
rect 1662 683 1674 939
rect 1708 683 1720 939
rect 1662 671 1720 683
rect 1840 939 1898 951
rect 1840 683 1852 939
rect 1886 683 1898 939
rect 1840 671 1898 683
rect 2018 939 2076 951
rect 2018 683 2030 939
rect 2064 683 2076 939
rect 2018 671 2076 683
rect 2196 939 2254 951
rect 2196 683 2208 939
rect 2242 683 2254 939
rect 2196 671 2254 683
rect 2374 939 2432 951
rect 2374 683 2386 939
rect 2420 683 2432 939
rect 2374 671 2432 683
rect 2552 939 2610 951
rect 2552 683 2564 939
rect 2598 683 2610 939
rect 2552 671 2610 683
rect 2730 939 2788 951
rect 2730 683 2742 939
rect 2776 683 2788 939
rect 2730 671 2788 683
rect 2908 939 2966 951
rect 2908 683 2920 939
rect 2954 683 2966 939
rect 2908 671 2966 683
rect 3086 939 3144 951
rect 3086 683 3098 939
rect 3132 683 3144 939
rect 3086 671 3144 683
rect 3264 939 3322 951
rect 3264 683 3276 939
rect 3310 683 3322 939
rect 3264 671 3322 683
rect 3442 939 3500 951
rect 3442 683 3454 939
rect 3488 683 3500 939
rect 3442 671 3500 683
rect 3620 939 3678 951
rect 3620 683 3632 939
rect 3666 683 3678 939
rect 3620 671 3678 683
rect 3816 939 3874 951
rect 3816 683 3828 939
rect 3862 683 3874 939
rect 3816 671 3874 683
rect 3994 939 4052 951
rect 3994 683 4006 939
rect 4040 683 4052 939
rect 3994 671 4052 683
rect 4172 939 4230 951
rect 4172 683 4184 939
rect 4218 683 4230 939
rect 4172 671 4230 683
rect 4350 939 4408 951
rect 4350 683 4362 939
rect 4396 683 4408 939
rect 4350 671 4408 683
rect 4528 939 4586 951
rect 4528 683 4540 939
rect 4574 683 4586 939
rect 4528 671 4586 683
rect 4706 939 4764 951
rect 4706 683 4718 939
rect 4752 683 4764 939
rect 4706 671 4764 683
rect 4884 939 4942 951
rect 4884 683 4896 939
rect 4930 683 4942 939
rect 4884 671 4942 683
rect 5062 939 5120 951
rect 5062 683 5074 939
rect 5108 683 5120 939
rect 5062 671 5120 683
rect 5240 939 5298 951
rect 5240 683 5252 939
rect 5286 683 5298 939
rect 5240 671 5298 683
rect 5418 939 5476 951
rect 5418 683 5430 939
rect 5464 683 5476 939
rect 5418 671 5476 683
rect 5596 939 5654 951
rect 5596 683 5608 939
rect 5642 683 5654 939
rect 5596 671 5654 683
rect 5774 939 5832 951
rect 5774 683 5786 939
rect 5820 683 5832 939
rect 5774 671 5832 683
rect 5952 939 6010 951
rect 5952 683 5964 939
rect 5998 683 6010 939
rect 5952 671 6010 683
rect 6130 939 6188 951
rect 6130 683 6142 939
rect 6176 683 6188 939
rect 6130 671 6188 683
rect 6308 939 6366 951
rect 6308 683 6320 939
rect 6354 683 6366 939
rect 6308 671 6366 683
rect 6486 939 6544 951
rect 6486 683 6498 939
rect 6532 683 6544 939
rect 6486 671 6544 683
rect 6664 939 6722 951
rect 6664 683 6676 939
rect 6710 683 6722 939
rect 6664 671 6722 683
rect 6842 939 6900 951
rect 6842 683 6854 939
rect 6888 683 6900 939
rect 6842 671 6900 683
rect 7020 939 7078 951
rect 7020 683 7032 939
rect 7066 683 7078 939
rect 7020 671 7078 683
rect 7545 939 7603 951
rect 7545 683 7557 939
rect 7591 683 7603 939
rect 7545 671 7603 683
rect 7723 939 7781 951
rect 7723 683 7735 939
rect 7769 683 7781 939
rect 7723 671 7781 683
rect 7901 939 7959 951
rect 7901 683 7913 939
rect 7947 683 7959 939
rect 7901 671 7959 683
rect 8079 939 8137 951
rect 8079 683 8091 939
rect 8125 683 8137 939
rect 8079 671 8137 683
rect 8257 939 8315 951
rect 8257 683 8269 939
rect 8303 683 8315 939
rect 8257 671 8315 683
rect 8435 939 8493 951
rect 8435 683 8447 939
rect 8481 683 8493 939
rect 8435 671 8493 683
rect 8613 939 8671 951
rect 8613 683 8625 939
rect 8659 683 8671 939
rect 8613 671 8671 683
rect 8791 939 8849 951
rect 8791 683 8803 939
rect 8837 683 8849 939
rect 8791 671 8849 683
rect 8969 939 9027 951
rect 8969 683 8981 939
rect 9015 683 9027 939
rect 8969 671 9027 683
rect 9147 939 9205 951
rect 9147 683 9159 939
rect 9193 683 9205 939
rect 9147 671 9205 683
rect 9325 939 9383 951
rect 9325 683 9337 939
rect 9371 683 9383 939
rect 9325 671 9383 683
rect 9503 939 9561 951
rect 9503 683 9515 939
rect 9549 683 9561 939
rect 9503 671 9561 683
rect 9681 939 9739 951
rect 9681 683 9693 939
rect 9727 683 9739 939
rect 9681 671 9739 683
rect 9859 939 9917 951
rect 9859 683 9871 939
rect 9905 683 9917 939
rect 9859 671 9917 683
rect 10037 939 10095 951
rect 10037 683 10049 939
rect 10083 683 10095 939
rect 10037 671 10095 683
rect 10232 939 10290 951
rect 10232 683 10244 939
rect 10278 683 10290 939
rect 10232 671 10290 683
rect 10410 939 10468 951
rect 10410 683 10422 939
rect 10456 683 10468 939
rect 10410 671 10468 683
rect 10588 939 10646 951
rect 10588 683 10600 939
rect 10634 683 10646 939
rect 10588 671 10646 683
rect 10766 939 10824 951
rect 10766 683 10778 939
rect 10812 683 10824 939
rect 10766 671 10824 683
rect 10944 939 11002 951
rect 10944 683 10956 939
rect 10990 683 11002 939
rect 10944 671 11002 683
rect 11122 939 11180 951
rect 11122 683 11134 939
rect 11168 683 11180 939
rect 11122 671 11180 683
rect 11300 939 11358 951
rect 11300 683 11312 939
rect 11346 683 11358 939
rect 11300 671 11358 683
rect 11478 939 11536 951
rect 11478 683 11490 939
rect 11524 683 11536 939
rect 11478 671 11536 683
rect 11656 939 11714 951
rect 11656 683 11668 939
rect 11702 683 11714 939
rect 11656 671 11714 683
rect 11834 939 11892 951
rect 11834 683 11846 939
rect 11880 683 11892 939
rect 11834 671 11892 683
rect 12012 939 12070 951
rect 12012 683 12024 939
rect 12058 683 12070 939
rect 12012 671 12070 683
rect 12190 939 12248 951
rect 12190 683 12202 939
rect 12236 683 12248 939
rect 12190 671 12248 683
rect 12368 939 12426 951
rect 12368 683 12380 939
rect 12414 683 12426 939
rect 12368 671 12426 683
rect 12546 939 12604 951
rect 12546 683 12558 939
rect 12592 683 12604 939
rect 12546 671 12604 683
rect 12724 939 12782 951
rect 12724 683 12736 939
rect 12770 683 12782 939
rect 12724 671 12782 683
rect 13538 5047 13596 5059
rect 13538 4791 13550 5047
rect 13584 4791 13596 5047
rect 13538 4779 13596 4791
rect 13716 5047 13774 5059
rect 13716 4791 13728 5047
rect 13762 4791 13774 5047
rect 13716 4779 13774 4791
rect 13894 5047 13952 5059
rect 13894 4791 13906 5047
rect 13940 4791 13952 5047
rect 13894 4779 13952 4791
rect 14072 5047 14130 5059
rect 14072 4791 14084 5047
rect 14118 4791 14130 5047
rect 14072 4779 14130 4791
rect 14250 5047 14308 5059
rect 14250 4791 14262 5047
rect 14296 4791 14308 5047
rect 14250 4779 14308 4791
rect 14428 5047 14486 5059
rect 14428 4791 14440 5047
rect 14474 4791 14486 5047
rect 14428 4779 14486 4791
rect 14606 5047 14664 5059
rect 14606 4791 14618 5047
rect 14652 4791 14664 5047
rect 14606 4779 14664 4791
rect 14784 5047 14842 5059
rect 14784 4791 14796 5047
rect 14830 4791 14842 5047
rect 14784 4779 14842 4791
rect 14962 5047 15020 5059
rect 14962 4791 14974 5047
rect 15008 4791 15020 5047
rect 14962 4779 15020 4791
rect 15140 5047 15198 5059
rect 15140 4791 15152 5047
rect 15186 4791 15198 5047
rect 15140 4779 15198 4791
rect 15318 5047 15376 5059
rect 15318 4791 15330 5047
rect 15364 4791 15376 5047
rect 15318 4779 15376 4791
rect 15496 5047 15554 5059
rect 15496 4791 15508 5047
rect 15542 4791 15554 5047
rect 15496 4779 15554 4791
rect 15674 5047 15732 5059
rect 15674 4791 15686 5047
rect 15720 4791 15732 5047
rect 15674 4779 15732 4791
rect 15852 5047 15910 5059
rect 15852 4791 15864 5047
rect 15898 4791 15910 5047
rect 15852 4779 15910 4791
rect 16030 5047 16088 5059
rect 16030 4791 16042 5047
rect 16076 4791 16088 5047
rect 16030 4779 16088 4791
rect 16208 5047 16266 5059
rect 16208 4791 16220 5047
rect 16254 4791 16266 5047
rect 16208 4779 16266 4791
rect 16386 5047 16444 5059
rect 16386 4791 16398 5047
rect 16432 4791 16444 5047
rect 16386 4779 16444 4791
rect 16564 5047 16622 5059
rect 16564 4791 16576 5047
rect 16610 4791 16622 5047
rect 16564 4779 16622 4791
rect 16742 5047 16800 5059
rect 16742 4791 16754 5047
rect 16788 4791 16800 5047
rect 16742 4779 16800 4791
rect 16920 5047 16978 5059
rect 16920 4791 16932 5047
rect 16966 4791 16978 5047
rect 16920 4779 16978 4791
rect 17098 5047 17156 5059
rect 17098 4791 17110 5047
rect 17144 4791 17156 5047
rect 17098 4779 17156 4791
rect 17276 5047 17334 5059
rect 17276 4791 17288 5047
rect 17322 4791 17334 5047
rect 17276 4779 17334 4791
rect 17454 5047 17512 5059
rect 17454 4791 17466 5047
rect 17500 4791 17512 5047
rect 17454 4779 17512 4791
rect 17632 5047 17690 5059
rect 17632 4791 17644 5047
rect 17678 4791 17690 5047
rect 17632 4779 17690 4791
rect 17810 5047 17868 5059
rect 17810 4791 17822 5047
rect 17856 4791 17868 5047
rect 17810 4779 17868 4791
rect 17988 5047 18046 5059
rect 17988 4791 18000 5047
rect 18034 4791 18046 5047
rect 17988 4779 18046 4791
rect 18166 5047 18224 5059
rect 18166 4791 18178 5047
rect 18212 4791 18224 5047
rect 18166 4779 18224 4791
rect 18344 5047 18402 5059
rect 18344 4791 18356 5047
rect 18390 4791 18402 5047
rect 18344 4779 18402 4791
rect 13538 4547 13596 4559
rect 13538 4291 13550 4547
rect 13584 4291 13596 4547
rect 13538 4279 13596 4291
rect 13716 4547 13774 4559
rect 13716 4291 13728 4547
rect 13762 4291 13774 4547
rect 13716 4279 13774 4291
rect 13894 4547 13952 4559
rect 13894 4291 13906 4547
rect 13940 4291 13952 4547
rect 13894 4279 13952 4291
rect 14072 4547 14130 4559
rect 14072 4291 14084 4547
rect 14118 4291 14130 4547
rect 14072 4279 14130 4291
rect 14250 4547 14308 4559
rect 14250 4291 14262 4547
rect 14296 4291 14308 4547
rect 14250 4279 14308 4291
rect 14428 4547 14486 4559
rect 14428 4291 14440 4547
rect 14474 4291 14486 4547
rect 14428 4279 14486 4291
rect 14606 4547 14664 4559
rect 14606 4291 14618 4547
rect 14652 4291 14664 4547
rect 14606 4279 14664 4291
rect 14784 4547 14842 4559
rect 14784 4291 14796 4547
rect 14830 4291 14842 4547
rect 14784 4279 14842 4291
rect 14962 4547 15020 4559
rect 14962 4291 14974 4547
rect 15008 4291 15020 4547
rect 14962 4279 15020 4291
rect 15140 4547 15198 4559
rect 15140 4291 15152 4547
rect 15186 4291 15198 4547
rect 15140 4279 15198 4291
rect 15318 4547 15376 4559
rect 15318 4291 15330 4547
rect 15364 4291 15376 4547
rect 15318 4279 15376 4291
rect 15496 4547 15554 4559
rect 15496 4291 15508 4547
rect 15542 4291 15554 4547
rect 15496 4279 15554 4291
rect 15674 4547 15732 4559
rect 15674 4291 15686 4547
rect 15720 4291 15732 4547
rect 15674 4279 15732 4291
rect 15852 4547 15910 4559
rect 15852 4291 15864 4547
rect 15898 4291 15910 4547
rect 15852 4279 15910 4291
rect 16030 4547 16088 4559
rect 16030 4291 16042 4547
rect 16076 4291 16088 4547
rect 16030 4279 16088 4291
rect 16208 4547 16266 4559
rect 16208 4291 16220 4547
rect 16254 4291 16266 4547
rect 16208 4279 16266 4291
rect 16386 4547 16444 4559
rect 16386 4291 16398 4547
rect 16432 4291 16444 4547
rect 16386 4279 16444 4291
rect 16564 4547 16622 4559
rect 16564 4291 16576 4547
rect 16610 4291 16622 4547
rect 16564 4279 16622 4291
rect 16742 4547 16800 4559
rect 16742 4291 16754 4547
rect 16788 4291 16800 4547
rect 16742 4279 16800 4291
rect 16920 4547 16978 4559
rect 16920 4291 16932 4547
rect 16966 4291 16978 4547
rect 16920 4279 16978 4291
rect 17098 4547 17156 4559
rect 17098 4291 17110 4547
rect 17144 4291 17156 4547
rect 17098 4279 17156 4291
rect 17276 4547 17334 4559
rect 17276 4291 17288 4547
rect 17322 4291 17334 4547
rect 17276 4279 17334 4291
rect 17454 4547 17512 4559
rect 17454 4291 17466 4547
rect 17500 4291 17512 4547
rect 17454 4279 17512 4291
rect 17632 4547 17690 4559
rect 17632 4291 17644 4547
rect 17678 4291 17690 4547
rect 17632 4279 17690 4291
rect 17810 4547 17868 4559
rect 17810 4291 17822 4547
rect 17856 4291 17868 4547
rect 17810 4279 17868 4291
rect 17988 4547 18046 4559
rect 17988 4291 18000 4547
rect 18034 4291 18046 4547
rect 17988 4279 18046 4291
rect 18166 4547 18224 4559
rect 18166 4291 18178 4547
rect 18212 4291 18224 4547
rect 18166 4279 18224 4291
rect 18344 4547 18402 4559
rect 18344 4291 18356 4547
rect 18390 4291 18402 4547
rect 18344 4279 18402 4291
rect 17096 3543 17154 3555
rect 17096 3287 17108 3543
rect 17142 3287 17154 3543
rect 17096 3275 17154 3287
rect 17274 3543 17332 3555
rect 17274 3287 17286 3543
rect 17320 3287 17332 3543
rect 17274 3275 17332 3287
rect 17452 3543 17510 3555
rect 17452 3287 17464 3543
rect 17498 3287 17510 3543
rect 17452 3275 17510 3287
rect 17630 3543 17688 3555
rect 17630 3287 17642 3543
rect 17676 3287 17688 3543
rect 17630 3275 17688 3287
rect 17808 3543 17866 3555
rect 17808 3287 17820 3543
rect 17854 3287 17866 3543
rect 17808 3275 17866 3287
rect 16382 2604 16440 2616
rect 13664 2538 13722 2550
rect 13664 2282 13676 2538
rect 13710 2282 13722 2538
rect 13664 2270 13722 2282
rect 13842 2538 13900 2550
rect 13842 2282 13854 2538
rect 13888 2282 13900 2538
rect 13842 2270 13900 2282
rect 13956 2538 14014 2550
rect 13956 2282 13968 2538
rect 14002 2282 14014 2538
rect 13956 2270 14014 2282
rect 14134 2538 14192 2550
rect 14134 2282 14146 2538
rect 14180 2282 14192 2538
rect 14134 2270 14192 2282
rect 14248 2538 14306 2550
rect 14248 2282 14260 2538
rect 14294 2282 14306 2538
rect 14248 2270 14306 2282
rect 14426 2538 14484 2550
rect 14426 2282 14438 2538
rect 14472 2282 14484 2538
rect 14426 2270 14484 2282
rect 14540 2538 14598 2550
rect 14540 2282 14552 2538
rect 14586 2282 14598 2538
rect 14540 2270 14598 2282
rect 14718 2538 14776 2550
rect 14718 2282 14730 2538
rect 14764 2282 14776 2538
rect 14718 2270 14776 2282
rect 14832 2538 14890 2550
rect 14832 2282 14844 2538
rect 14878 2282 14890 2538
rect 14832 2270 14890 2282
rect 15010 2538 15068 2550
rect 15010 2282 15022 2538
rect 15056 2282 15068 2538
rect 15010 2270 15068 2282
rect 15124 2538 15182 2550
rect 15124 2282 15136 2538
rect 15170 2282 15182 2538
rect 15124 2270 15182 2282
rect 15302 2538 15360 2550
rect 15302 2282 15314 2538
rect 15348 2282 15360 2538
rect 15302 2270 15360 2282
rect 15416 2538 15474 2550
rect 15416 2282 15428 2538
rect 15462 2282 15474 2538
rect 15416 2270 15474 2282
rect 15594 2538 15652 2550
rect 15594 2282 15606 2538
rect 15640 2282 15652 2538
rect 16382 2348 16394 2604
rect 16428 2348 16440 2604
rect 16382 2336 16440 2348
rect 16560 2604 16618 2616
rect 16560 2348 16572 2604
rect 16606 2348 16618 2604
rect 16560 2336 16618 2348
rect 16738 2604 16796 2616
rect 16738 2348 16750 2604
rect 16784 2348 16796 2604
rect 16738 2336 16796 2348
rect 16916 2604 16974 2616
rect 16916 2348 16928 2604
rect 16962 2348 16974 2604
rect 16916 2336 16974 2348
rect 17094 2604 17152 2616
rect 17094 2348 17106 2604
rect 17140 2348 17152 2604
rect 17094 2336 17152 2348
rect 17272 2604 17330 2616
rect 17272 2348 17284 2604
rect 17318 2348 17330 2604
rect 17272 2336 17330 2348
rect 17450 2604 17508 2616
rect 17450 2348 17462 2604
rect 17496 2348 17508 2604
rect 17450 2336 17508 2348
rect 17628 2604 17686 2616
rect 17628 2348 17640 2604
rect 17674 2348 17686 2604
rect 17628 2336 17686 2348
rect 17806 2604 17864 2616
rect 17806 2348 17818 2604
rect 17852 2348 17864 2604
rect 17806 2336 17864 2348
rect 17984 2604 18042 2616
rect 17984 2348 17996 2604
rect 18030 2348 18042 2604
rect 17984 2336 18042 2348
rect 18162 2604 18220 2616
rect 18162 2348 18174 2604
rect 18208 2348 18220 2604
rect 18162 2336 18220 2348
rect 18340 2604 18398 2616
rect 18340 2348 18352 2604
rect 18386 2348 18398 2604
rect 18340 2336 18398 2348
rect 15594 2270 15652 2282
rect 16382 2104 16440 2116
rect 13664 2040 13722 2052
rect 13664 1784 13676 2040
rect 13710 1784 13722 2040
rect 13664 1772 13722 1784
rect 13842 2040 13900 2052
rect 13842 1784 13854 2040
rect 13888 1784 13900 2040
rect 13842 1772 13900 1784
rect 13956 2040 14014 2052
rect 13956 1784 13968 2040
rect 14002 1784 14014 2040
rect 13956 1772 14014 1784
rect 14134 2040 14192 2052
rect 14134 1784 14146 2040
rect 14180 1784 14192 2040
rect 14134 1772 14192 1784
rect 14248 2040 14306 2052
rect 14248 1784 14260 2040
rect 14294 1784 14306 2040
rect 14248 1772 14306 1784
rect 14426 2040 14484 2052
rect 14426 1784 14438 2040
rect 14472 1784 14484 2040
rect 14426 1772 14484 1784
rect 14540 2040 14598 2052
rect 14540 1784 14552 2040
rect 14586 1784 14598 2040
rect 14540 1772 14598 1784
rect 14718 2040 14776 2052
rect 14718 1784 14730 2040
rect 14764 1784 14776 2040
rect 14718 1772 14776 1784
rect 14832 2040 14890 2052
rect 14832 1784 14844 2040
rect 14878 1784 14890 2040
rect 14832 1772 14890 1784
rect 15010 2040 15068 2052
rect 15010 1784 15022 2040
rect 15056 1784 15068 2040
rect 15010 1772 15068 1784
rect 15124 2040 15182 2052
rect 15124 1784 15136 2040
rect 15170 1784 15182 2040
rect 15124 1772 15182 1784
rect 15302 2040 15360 2052
rect 15302 1784 15314 2040
rect 15348 1784 15360 2040
rect 15302 1772 15360 1784
rect 15416 2040 15474 2052
rect 15416 1784 15428 2040
rect 15462 1784 15474 2040
rect 15416 1772 15474 1784
rect 15594 2040 15652 2052
rect 15594 1784 15606 2040
rect 15640 1784 15652 2040
rect 16382 1848 16394 2104
rect 16428 1848 16440 2104
rect 16382 1836 16440 1848
rect 16560 2104 16618 2116
rect 16560 1848 16572 2104
rect 16606 1848 16618 2104
rect 16560 1836 16618 1848
rect 16738 2104 16796 2116
rect 16738 1848 16750 2104
rect 16784 1848 16796 2104
rect 16738 1836 16796 1848
rect 16916 2104 16974 2116
rect 16916 1848 16928 2104
rect 16962 1848 16974 2104
rect 16916 1836 16974 1848
rect 17094 2104 17152 2116
rect 17094 1848 17106 2104
rect 17140 1848 17152 2104
rect 17094 1836 17152 1848
rect 17272 2104 17330 2116
rect 17272 1848 17284 2104
rect 17318 1848 17330 2104
rect 17272 1836 17330 1848
rect 17450 2104 17508 2116
rect 17450 1848 17462 2104
rect 17496 1848 17508 2104
rect 17450 1836 17508 1848
rect 17628 2104 17686 2116
rect 17628 1848 17640 2104
rect 17674 1848 17686 2104
rect 17628 1836 17686 1848
rect 17806 2104 17864 2116
rect 17806 1848 17818 2104
rect 17852 1848 17864 2104
rect 17806 1836 17864 1848
rect 17984 2104 18042 2116
rect 17984 1848 17996 2104
rect 18030 1848 18042 2104
rect 17984 1836 18042 1848
rect 18162 2104 18220 2116
rect 18162 1848 18174 2104
rect 18208 1848 18220 2104
rect 18162 1836 18220 1848
rect 18340 2104 18398 2116
rect 18340 1848 18352 2104
rect 18386 1848 18398 2104
rect 18340 1836 18398 1848
rect 15594 1772 15652 1784
rect 13664 1542 13722 1554
rect 13664 1286 13676 1542
rect 13710 1286 13722 1542
rect 13664 1274 13722 1286
rect 13842 1542 13900 1554
rect 13842 1286 13854 1542
rect 13888 1286 13900 1542
rect 13842 1274 13900 1286
rect 13956 1542 14014 1554
rect 13956 1286 13968 1542
rect 14002 1286 14014 1542
rect 13956 1274 14014 1286
rect 14134 1542 14192 1554
rect 14134 1286 14146 1542
rect 14180 1286 14192 1542
rect 14134 1274 14192 1286
rect 14248 1542 14306 1554
rect 14248 1286 14260 1542
rect 14294 1286 14306 1542
rect 14248 1274 14306 1286
rect 14426 1542 14484 1554
rect 14426 1286 14438 1542
rect 14472 1286 14484 1542
rect 14426 1274 14484 1286
rect 14540 1542 14598 1554
rect 14540 1286 14552 1542
rect 14586 1286 14598 1542
rect 14540 1274 14598 1286
rect 14718 1542 14776 1554
rect 14718 1286 14730 1542
rect 14764 1286 14776 1542
rect 14718 1274 14776 1286
rect 14832 1542 14890 1554
rect 14832 1286 14844 1542
rect 14878 1286 14890 1542
rect 14832 1274 14890 1286
rect 15010 1542 15068 1554
rect 15010 1286 15022 1542
rect 15056 1286 15068 1542
rect 15010 1274 15068 1286
rect 15124 1542 15182 1554
rect 15124 1286 15136 1542
rect 15170 1286 15182 1542
rect 15124 1274 15182 1286
rect 15302 1542 15360 1554
rect 15302 1286 15314 1542
rect 15348 1286 15360 1542
rect 15302 1274 15360 1286
rect 15416 1542 15474 1554
rect 15416 1286 15428 1542
rect 15462 1286 15474 1542
rect 15416 1274 15474 1286
rect 15594 1542 15652 1554
rect 15594 1286 15606 1542
rect 15640 1286 15652 1542
rect 15594 1274 15652 1286
rect 16382 1544 16440 1556
rect 16382 1288 16394 1544
rect 16428 1288 16440 1544
rect 16382 1276 16440 1288
rect 16560 1544 16618 1556
rect 16560 1288 16572 1544
rect 16606 1288 16618 1544
rect 16560 1276 16618 1288
rect 16738 1544 16796 1556
rect 16738 1288 16750 1544
rect 16784 1288 16796 1544
rect 16738 1276 16796 1288
rect 16916 1544 16974 1556
rect 16916 1288 16928 1544
rect 16962 1288 16974 1544
rect 16916 1276 16974 1288
rect 17094 1544 17152 1556
rect 17094 1288 17106 1544
rect 17140 1288 17152 1544
rect 17094 1276 17152 1288
rect 17272 1544 17330 1556
rect 17272 1288 17284 1544
rect 17318 1288 17330 1544
rect 17272 1276 17330 1288
rect 17450 1544 17508 1556
rect 17450 1288 17462 1544
rect 17496 1288 17508 1544
rect 17450 1276 17508 1288
rect 17628 1544 17686 1556
rect 17628 1288 17640 1544
rect 17674 1288 17686 1544
rect 17628 1276 17686 1288
rect 17806 1544 17864 1556
rect 17806 1288 17818 1544
rect 17852 1288 17864 1544
rect 17806 1276 17864 1288
rect 17984 1544 18042 1556
rect 17984 1288 17996 1544
rect 18030 1288 18042 1544
rect 17984 1276 18042 1288
rect 18162 1544 18220 1556
rect 18162 1288 18174 1544
rect 18208 1288 18220 1544
rect 18162 1276 18220 1288
rect 18340 1544 18398 1556
rect 18340 1288 18352 1544
rect 18386 1288 18398 1544
rect 18340 1276 18398 1288
rect 13664 1044 13722 1056
rect 13664 788 13676 1044
rect 13710 788 13722 1044
rect 13664 776 13722 788
rect 13842 1044 13900 1056
rect 13842 788 13854 1044
rect 13888 788 13900 1044
rect 13842 776 13900 788
rect 13956 1044 14014 1056
rect 13956 788 13968 1044
rect 14002 788 14014 1044
rect 13956 776 14014 788
rect 14134 1044 14192 1056
rect 14134 788 14146 1044
rect 14180 788 14192 1044
rect 14134 776 14192 788
rect 14248 1044 14306 1056
rect 14248 788 14260 1044
rect 14294 788 14306 1044
rect 14248 776 14306 788
rect 14426 1044 14484 1056
rect 14426 788 14438 1044
rect 14472 788 14484 1044
rect 14426 776 14484 788
rect 14540 1044 14598 1056
rect 14540 788 14552 1044
rect 14586 788 14598 1044
rect 14540 776 14598 788
rect 14718 1044 14776 1056
rect 14718 788 14730 1044
rect 14764 788 14776 1044
rect 14718 776 14776 788
rect 14832 1044 14890 1056
rect 14832 788 14844 1044
rect 14878 788 14890 1044
rect 14832 776 14890 788
rect 15010 1044 15068 1056
rect 15010 788 15022 1044
rect 15056 788 15068 1044
rect 15010 776 15068 788
rect 15124 1044 15182 1056
rect 15124 788 15136 1044
rect 15170 788 15182 1044
rect 15124 776 15182 788
rect 15302 1044 15360 1056
rect 15302 788 15314 1044
rect 15348 788 15360 1044
rect 15302 776 15360 788
rect 15416 1044 15474 1056
rect 15416 788 15428 1044
rect 15462 788 15474 1044
rect 15416 776 15474 788
rect 15594 1044 15652 1056
rect 15594 788 15606 1044
rect 15640 788 15652 1044
rect 15594 776 15652 788
rect 16382 1044 16440 1056
rect 16382 788 16394 1044
rect 16428 788 16440 1044
rect 16382 776 16440 788
rect 16560 1044 16618 1056
rect 16560 788 16572 1044
rect 16606 788 16618 1044
rect 16560 776 16618 788
rect 16738 1044 16796 1056
rect 16738 788 16750 1044
rect 16784 788 16796 1044
rect 16738 776 16796 788
rect 16916 1044 16974 1056
rect 16916 788 16928 1044
rect 16962 788 16974 1044
rect 16916 776 16974 788
rect 17094 1044 17152 1056
rect 17094 788 17106 1044
rect 17140 788 17152 1044
rect 17094 776 17152 788
rect 17272 1044 17330 1056
rect 17272 788 17284 1044
rect 17318 788 17330 1044
rect 17272 776 17330 788
rect 17450 1044 17508 1056
rect 17450 788 17462 1044
rect 17496 788 17508 1044
rect 17450 776 17508 788
rect 17628 1044 17686 1056
rect 17628 788 17640 1044
rect 17674 788 17686 1044
rect 17628 776 17686 788
rect 17806 1044 17864 1056
rect 17806 788 17818 1044
rect 17852 788 17864 1044
rect 17806 776 17864 788
rect 17984 1044 18042 1056
rect 17984 788 17996 1044
rect 18030 788 18042 1044
rect 17984 776 18042 788
rect 18162 1044 18220 1056
rect 18162 788 18174 1044
rect 18208 788 18220 1044
rect 18162 776 18220 788
rect 18340 1044 18398 1056
rect 18340 788 18352 1044
rect 18386 788 18398 1044
rect 18340 776 18398 788
rect 18997 5038 19055 5050
rect 18997 4782 19009 5038
rect 19043 4782 19055 5038
rect 18997 4770 19055 4782
rect 19175 5038 19233 5050
rect 19175 4782 19187 5038
rect 19221 4782 19233 5038
rect 19175 4770 19233 4782
rect 19353 5038 19411 5050
rect 19353 4782 19365 5038
rect 19399 4782 19411 5038
rect 19353 4770 19411 4782
rect 19531 5038 19589 5050
rect 19531 4782 19543 5038
rect 19577 4782 19589 5038
rect 19531 4770 19589 4782
rect 19709 5038 19767 5050
rect 19709 4782 19721 5038
rect 19755 4782 19767 5038
rect 19709 4770 19767 4782
rect 19887 5038 19945 5050
rect 19887 4782 19899 5038
rect 19933 4782 19945 5038
rect 19887 4770 19945 4782
rect 20065 5038 20123 5050
rect 20065 4782 20077 5038
rect 20111 4782 20123 5038
rect 20065 4770 20123 4782
rect 20243 5038 20301 5050
rect 20243 4782 20255 5038
rect 20289 4782 20301 5038
rect 20243 4770 20301 4782
rect 20421 5038 20479 5050
rect 20421 4782 20433 5038
rect 20467 4782 20479 5038
rect 20421 4770 20479 4782
rect 20599 5038 20657 5050
rect 20599 4782 20611 5038
rect 20645 4782 20657 5038
rect 20599 4770 20657 4782
rect 20777 5038 20835 5050
rect 20777 4782 20789 5038
rect 20823 4782 20835 5038
rect 20777 4770 20835 4782
rect 20955 5038 21013 5050
rect 20955 4782 20967 5038
rect 21001 4782 21013 5038
rect 20955 4770 21013 4782
rect 21133 5038 21191 5050
rect 21133 4782 21145 5038
rect 21179 4782 21191 5038
rect 21133 4770 21191 4782
rect 21311 5038 21369 5050
rect 21311 4782 21323 5038
rect 21357 4782 21369 5038
rect 21311 4770 21369 4782
rect 21489 5038 21547 5050
rect 21489 4782 21501 5038
rect 21535 4782 21547 5038
rect 21489 4770 21547 4782
rect 21667 5038 21725 5050
rect 21667 4782 21679 5038
rect 21713 4782 21725 5038
rect 21667 4770 21725 4782
rect 21845 5038 21903 5050
rect 21845 4782 21857 5038
rect 21891 4782 21903 5038
rect 21845 4770 21903 4782
rect 18997 4540 19055 4552
rect 18997 4284 19009 4540
rect 19043 4284 19055 4540
rect 18997 4272 19055 4284
rect 19175 4540 19233 4552
rect 19175 4284 19187 4540
rect 19221 4284 19233 4540
rect 19175 4272 19233 4284
rect 19353 4540 19411 4552
rect 19353 4284 19365 4540
rect 19399 4284 19411 4540
rect 19353 4272 19411 4284
rect 19531 4540 19589 4552
rect 19531 4284 19543 4540
rect 19577 4284 19589 4540
rect 19531 4272 19589 4284
rect 19709 4540 19767 4552
rect 19709 4284 19721 4540
rect 19755 4284 19767 4540
rect 19709 4272 19767 4284
rect 19887 4540 19945 4552
rect 19887 4284 19899 4540
rect 19933 4284 19945 4540
rect 19887 4272 19945 4284
rect 20065 4540 20123 4552
rect 20065 4284 20077 4540
rect 20111 4284 20123 4540
rect 20065 4272 20123 4284
rect 20243 4540 20301 4552
rect 20243 4284 20255 4540
rect 20289 4284 20301 4540
rect 20243 4272 20301 4284
rect 20421 4540 20479 4552
rect 20421 4284 20433 4540
rect 20467 4284 20479 4540
rect 20421 4272 20479 4284
rect 20599 4540 20657 4552
rect 20599 4284 20611 4540
rect 20645 4284 20657 4540
rect 20599 4272 20657 4284
rect 20777 4540 20835 4552
rect 20777 4284 20789 4540
rect 20823 4284 20835 4540
rect 20777 4272 20835 4284
rect 20955 4540 21013 4552
rect 20955 4284 20967 4540
rect 21001 4284 21013 4540
rect 20955 4272 21013 4284
rect 21133 4540 21191 4552
rect 21133 4284 21145 4540
rect 21179 4284 21191 4540
rect 21133 4272 21191 4284
rect 21311 4540 21369 4552
rect 21311 4284 21323 4540
rect 21357 4284 21369 4540
rect 21311 4272 21369 4284
rect 21489 4540 21547 4552
rect 21489 4284 21501 4540
rect 21535 4284 21547 4540
rect 21489 4272 21547 4284
rect 21667 4540 21725 4552
rect 21667 4284 21679 4540
rect 21713 4284 21725 4540
rect 21667 4272 21725 4284
rect 21845 4540 21903 4552
rect 21845 4284 21857 4540
rect 21891 4284 21903 4540
rect 21845 4272 21903 4284
rect 18997 4042 19055 4054
rect 18997 3786 19009 4042
rect 19043 3786 19055 4042
rect 18997 3774 19055 3786
rect 19175 4042 19233 4054
rect 19175 3786 19187 4042
rect 19221 3786 19233 4042
rect 19175 3774 19233 3786
rect 19353 4042 19411 4054
rect 19353 3786 19365 4042
rect 19399 3786 19411 4042
rect 19353 3774 19411 3786
rect 19531 4042 19589 4054
rect 19531 3786 19543 4042
rect 19577 3786 19589 4042
rect 19531 3774 19589 3786
rect 19709 4042 19767 4054
rect 19709 3786 19721 4042
rect 19755 3786 19767 4042
rect 19709 3774 19767 3786
rect 19887 4042 19945 4054
rect 19887 3786 19899 4042
rect 19933 3786 19945 4042
rect 19887 3774 19945 3786
rect 20065 4042 20123 4054
rect 20065 3786 20077 4042
rect 20111 3786 20123 4042
rect 20065 3774 20123 3786
rect 20243 4042 20301 4054
rect 20243 3786 20255 4042
rect 20289 3786 20301 4042
rect 20243 3774 20301 3786
rect 20421 4042 20479 4054
rect 20421 3786 20433 4042
rect 20467 3786 20479 4042
rect 20421 3774 20479 3786
rect 20599 4042 20657 4054
rect 20599 3786 20611 4042
rect 20645 3786 20657 4042
rect 20599 3774 20657 3786
rect 20777 4042 20835 4054
rect 20777 3786 20789 4042
rect 20823 3786 20835 4042
rect 20777 3774 20835 3786
rect 20955 4042 21013 4054
rect 20955 3786 20967 4042
rect 21001 3786 21013 4042
rect 20955 3774 21013 3786
rect 21133 4042 21191 4054
rect 21133 3786 21145 4042
rect 21179 3786 21191 4042
rect 21133 3774 21191 3786
rect 21311 4042 21369 4054
rect 21311 3786 21323 4042
rect 21357 3786 21369 4042
rect 21311 3774 21369 3786
rect 21489 4042 21547 4054
rect 21489 3786 21501 4042
rect 21535 3786 21547 4042
rect 21489 3774 21547 3786
rect 21667 4042 21725 4054
rect 21667 3786 21679 4042
rect 21713 3786 21725 4042
rect 21667 3774 21725 3786
rect 21845 4042 21903 4054
rect 21845 3786 21857 4042
rect 21891 3786 21903 4042
rect 21845 3774 21903 3786
rect 18997 3544 19055 3556
rect 18997 3288 19009 3544
rect 19043 3288 19055 3544
rect 18997 3276 19055 3288
rect 19175 3544 19233 3556
rect 19175 3288 19187 3544
rect 19221 3288 19233 3544
rect 19175 3276 19233 3288
rect 19353 3544 19411 3556
rect 19353 3288 19365 3544
rect 19399 3288 19411 3544
rect 19353 3276 19411 3288
rect 19531 3544 19589 3556
rect 19531 3288 19543 3544
rect 19577 3288 19589 3544
rect 19531 3276 19589 3288
rect 19709 3544 19767 3556
rect 19709 3288 19721 3544
rect 19755 3288 19767 3544
rect 19709 3276 19767 3288
rect 19887 3544 19945 3556
rect 19887 3288 19899 3544
rect 19933 3288 19945 3544
rect 19887 3276 19945 3288
rect 20065 3544 20123 3556
rect 20065 3288 20077 3544
rect 20111 3288 20123 3544
rect 20065 3276 20123 3288
rect 20243 3544 20301 3556
rect 20243 3288 20255 3544
rect 20289 3288 20301 3544
rect 20243 3276 20301 3288
rect 20421 3544 20479 3556
rect 20421 3288 20433 3544
rect 20467 3288 20479 3544
rect 20421 3276 20479 3288
rect 20599 3544 20657 3556
rect 20599 3288 20611 3544
rect 20645 3288 20657 3544
rect 20599 3276 20657 3288
rect 20777 3544 20835 3556
rect 20777 3288 20789 3544
rect 20823 3288 20835 3544
rect 20777 3276 20835 3288
rect 20955 3544 21013 3556
rect 20955 3288 20967 3544
rect 21001 3288 21013 3544
rect 20955 3276 21013 3288
rect 21133 3544 21191 3556
rect 21133 3288 21145 3544
rect 21179 3288 21191 3544
rect 21133 3276 21191 3288
rect 21311 3544 21369 3556
rect 21311 3288 21323 3544
rect 21357 3288 21369 3544
rect 21311 3276 21369 3288
rect 21489 3544 21547 3556
rect 21489 3288 21501 3544
rect 21535 3288 21547 3544
rect 21489 3276 21547 3288
rect 21667 3544 21725 3556
rect 21667 3288 21679 3544
rect 21713 3288 21725 3544
rect 21667 3276 21725 3288
rect 21845 3544 21903 3556
rect 21845 3288 21857 3544
rect 21891 3288 21903 3544
rect 21845 3276 21903 3288
rect 19355 2530 19413 2542
rect 19355 2274 19367 2530
rect 19401 2274 19413 2530
rect 19355 2262 19413 2274
rect 19533 2530 19591 2542
rect 19533 2274 19545 2530
rect 19579 2274 19591 2530
rect 19533 2262 19591 2274
rect 19711 2530 19769 2542
rect 19711 2274 19723 2530
rect 19757 2274 19769 2530
rect 19711 2262 19769 2274
rect 19889 2530 19947 2542
rect 19889 2274 19901 2530
rect 19935 2274 19947 2530
rect 19889 2262 19947 2274
rect 20067 2530 20125 2542
rect 20067 2274 20079 2530
rect 20113 2274 20125 2530
rect 20067 2262 20125 2274
rect 20245 2530 20303 2542
rect 20245 2274 20257 2530
rect 20291 2274 20303 2530
rect 20245 2262 20303 2274
rect 20423 2530 20481 2542
rect 20423 2274 20435 2530
rect 20469 2274 20481 2530
rect 20423 2262 20481 2274
rect 20601 2530 20659 2542
rect 20601 2274 20613 2530
rect 20647 2274 20659 2530
rect 20601 2262 20659 2274
rect 20779 2530 20837 2542
rect 20779 2274 20791 2530
rect 20825 2274 20837 2530
rect 20779 2262 20837 2274
rect 20957 2530 21015 2542
rect 20957 2274 20969 2530
rect 21003 2274 21015 2530
rect 20957 2262 21015 2274
rect 21135 2530 21193 2542
rect 21135 2274 21147 2530
rect 21181 2274 21193 2530
rect 21135 2262 21193 2274
rect 21313 2530 21371 2542
rect 21313 2274 21325 2530
rect 21359 2274 21371 2530
rect 21313 2262 21371 2274
rect 19355 2032 19413 2044
rect 19355 1776 19367 2032
rect 19401 1776 19413 2032
rect 19355 1764 19413 1776
rect 19533 2032 19591 2044
rect 19533 1776 19545 2032
rect 19579 1776 19591 2032
rect 19533 1764 19591 1776
rect 19711 2032 19769 2044
rect 19711 1776 19723 2032
rect 19757 1776 19769 2032
rect 19711 1764 19769 1776
rect 19889 2032 19947 2044
rect 19889 1776 19901 2032
rect 19935 1776 19947 2032
rect 19889 1764 19947 1776
rect 20067 2032 20125 2044
rect 20067 1776 20079 2032
rect 20113 1776 20125 2032
rect 20067 1764 20125 1776
rect 20245 2032 20303 2044
rect 20245 1776 20257 2032
rect 20291 1776 20303 2032
rect 20245 1764 20303 1776
rect 20423 2032 20481 2044
rect 20423 1776 20435 2032
rect 20469 1776 20481 2032
rect 20423 1764 20481 1776
rect 20601 2032 20659 2044
rect 20601 1776 20613 2032
rect 20647 1776 20659 2032
rect 20601 1764 20659 1776
rect 20779 2032 20837 2044
rect 20779 1776 20791 2032
rect 20825 1776 20837 2032
rect 20779 1764 20837 1776
rect 20957 2032 21015 2044
rect 20957 1776 20969 2032
rect 21003 1776 21015 2032
rect 20957 1764 21015 1776
rect 21135 2032 21193 2044
rect 21135 1776 21147 2032
rect 21181 1776 21193 2032
rect 21135 1764 21193 1776
rect 21313 2032 21371 2044
rect 21313 1776 21325 2032
rect 21359 1776 21371 2032
rect 21313 1764 21371 1776
rect 19355 1534 19413 1546
rect 19355 1278 19367 1534
rect 19401 1278 19413 1534
rect 19355 1266 19413 1278
rect 19533 1534 19591 1546
rect 19533 1278 19545 1534
rect 19579 1278 19591 1534
rect 19533 1266 19591 1278
rect 19711 1534 19769 1546
rect 19711 1278 19723 1534
rect 19757 1278 19769 1534
rect 19711 1266 19769 1278
rect 19889 1534 19947 1546
rect 19889 1278 19901 1534
rect 19935 1278 19947 1534
rect 19889 1266 19947 1278
rect 20067 1534 20125 1546
rect 20067 1278 20079 1534
rect 20113 1278 20125 1534
rect 20067 1266 20125 1278
rect 20245 1534 20303 1546
rect 20245 1278 20257 1534
rect 20291 1278 20303 1534
rect 20245 1266 20303 1278
rect 20423 1534 20481 1546
rect 20423 1278 20435 1534
rect 20469 1278 20481 1534
rect 20423 1266 20481 1278
rect 20601 1534 20659 1546
rect 20601 1278 20613 1534
rect 20647 1278 20659 1534
rect 20601 1266 20659 1278
rect 20779 1534 20837 1546
rect 20779 1278 20791 1534
rect 20825 1278 20837 1534
rect 20779 1266 20837 1278
rect 20957 1534 21015 1546
rect 20957 1278 20969 1534
rect 21003 1278 21015 1534
rect 20957 1266 21015 1278
rect 21135 1534 21193 1546
rect 21135 1278 21147 1534
rect 21181 1278 21193 1534
rect 21135 1266 21193 1278
rect 21313 1534 21371 1546
rect 21313 1278 21325 1534
rect 21359 1278 21371 1534
rect 21313 1266 21371 1278
rect 19355 1036 19413 1048
rect 19355 780 19367 1036
rect 19401 780 19413 1036
rect 19355 768 19413 780
rect 19533 1036 19591 1048
rect 19533 780 19545 1036
rect 19579 780 19591 1036
rect 19533 768 19591 780
rect 19711 1036 19769 1048
rect 19711 780 19723 1036
rect 19757 780 19769 1036
rect 19711 768 19769 780
rect 19889 1036 19947 1048
rect 19889 780 19901 1036
rect 19935 780 19947 1036
rect 19889 768 19947 780
rect 20067 1036 20125 1048
rect 20067 780 20079 1036
rect 20113 780 20125 1036
rect 20067 768 20125 780
rect 20245 1036 20303 1048
rect 20245 780 20257 1036
rect 20291 780 20303 1036
rect 20245 768 20303 780
rect 20423 1036 20481 1048
rect 20423 780 20435 1036
rect 20469 780 20481 1036
rect 20423 768 20481 780
rect 20601 1036 20659 1048
rect 20601 780 20613 1036
rect 20647 780 20659 1036
rect 20601 768 20659 780
rect 20779 1036 20837 1048
rect 20779 780 20791 1036
rect 20825 780 20837 1036
rect 20779 768 20837 780
rect 20957 1036 21015 1048
rect 20957 780 20969 1036
rect 21003 780 21015 1036
rect 20957 768 21015 780
rect 21135 1036 21193 1048
rect 21135 780 21147 1036
rect 21181 780 21193 1036
rect 21135 768 21193 780
rect 21313 1036 21371 1048
rect 21313 780 21325 1036
rect 21359 780 21371 1036
rect 21313 768 21371 780
<< pdiff >>
rect 7291 18741 7353 18753
rect 7291 18493 7303 18741
rect 7337 18493 7353 18741
rect 7291 18481 7353 18493
rect 7383 18741 7449 18753
rect 7383 18493 7399 18741
rect 7433 18493 7449 18741
rect 7383 18481 7449 18493
rect 7479 18741 7545 18753
rect 7479 18493 7495 18741
rect 7529 18493 7545 18741
rect 7479 18481 7545 18493
rect 7575 18741 7641 18753
rect 7575 18493 7591 18741
rect 7625 18493 7641 18741
rect 7575 18481 7641 18493
rect 7671 18741 7737 18753
rect 7671 18493 7687 18741
rect 7721 18493 7737 18741
rect 7671 18481 7737 18493
rect 7767 18741 7833 18753
rect 7767 18493 7783 18741
rect 7817 18493 7833 18741
rect 7767 18481 7833 18493
rect 7863 18741 7929 18753
rect 7863 18493 7879 18741
rect 7913 18493 7929 18741
rect 7863 18481 7929 18493
rect 7959 18741 8025 18753
rect 7959 18493 7975 18741
rect 8009 18493 8025 18741
rect 7959 18481 8025 18493
rect 8055 18741 8121 18753
rect 8055 18493 8071 18741
rect 8105 18493 8121 18741
rect 8055 18481 8121 18493
rect 8151 18741 8217 18753
rect 8151 18493 8167 18741
rect 8201 18493 8217 18741
rect 8151 18481 8217 18493
rect 8247 18741 8309 18753
rect 8247 18493 8263 18741
rect 8297 18493 8309 18741
rect 8247 18481 8309 18493
rect 20221 18741 20283 18753
rect 20221 18493 20233 18741
rect 20267 18493 20283 18741
rect 20221 18481 20283 18493
rect 20313 18741 20379 18753
rect 20313 18493 20329 18741
rect 20363 18493 20379 18741
rect 20313 18481 20379 18493
rect 20409 18741 20475 18753
rect 20409 18493 20425 18741
rect 20459 18493 20475 18741
rect 20409 18481 20475 18493
rect 20505 18741 20571 18753
rect 20505 18493 20521 18741
rect 20555 18493 20571 18741
rect 20505 18481 20571 18493
rect 20601 18741 20667 18753
rect 20601 18493 20617 18741
rect 20651 18493 20667 18741
rect 20601 18481 20667 18493
rect 20697 18741 20763 18753
rect 20697 18493 20713 18741
rect 20747 18493 20763 18741
rect 20697 18481 20763 18493
rect 20793 18741 20859 18753
rect 20793 18493 20809 18741
rect 20843 18493 20859 18741
rect 20793 18481 20859 18493
rect 20889 18741 20955 18753
rect 20889 18493 20905 18741
rect 20939 18493 20955 18741
rect 20889 18481 20955 18493
rect 20985 18741 21051 18753
rect 20985 18493 21001 18741
rect 21035 18493 21051 18741
rect 20985 18481 21051 18493
rect 21081 18741 21147 18753
rect 21081 18493 21097 18741
rect 21131 18493 21147 18741
rect 21081 18481 21147 18493
rect 21177 18741 21239 18753
rect 21177 18493 21193 18741
rect 21227 18493 21239 18741
rect 21177 18481 21239 18493
rect 7291 16941 7353 16953
rect 7291 16693 7303 16941
rect 7337 16693 7353 16941
rect 7291 16681 7353 16693
rect 7383 16941 7449 16953
rect 7383 16693 7399 16941
rect 7433 16693 7449 16941
rect 7383 16681 7449 16693
rect 7479 16941 7545 16953
rect 7479 16693 7495 16941
rect 7529 16693 7545 16941
rect 7479 16681 7545 16693
rect 7575 16941 7641 16953
rect 7575 16693 7591 16941
rect 7625 16693 7641 16941
rect 7575 16681 7641 16693
rect 7671 16941 7737 16953
rect 7671 16693 7687 16941
rect 7721 16693 7737 16941
rect 7671 16681 7737 16693
rect 7767 16941 7833 16953
rect 7767 16693 7783 16941
rect 7817 16693 7833 16941
rect 7767 16681 7833 16693
rect 7863 16941 7929 16953
rect 7863 16693 7879 16941
rect 7913 16693 7929 16941
rect 7863 16681 7929 16693
rect 7959 16941 8025 16953
rect 7959 16693 7975 16941
rect 8009 16693 8025 16941
rect 7959 16681 8025 16693
rect 8055 16941 8121 16953
rect 8055 16693 8071 16941
rect 8105 16693 8121 16941
rect 8055 16681 8121 16693
rect 8151 16941 8217 16953
rect 8151 16693 8167 16941
rect 8201 16693 8217 16941
rect 8151 16681 8217 16693
rect 8247 16941 8309 16953
rect 8247 16693 8263 16941
rect 8297 16693 8309 16941
rect 8247 16681 8309 16693
rect 20221 16941 20283 16953
rect 20221 16693 20233 16941
rect 20267 16693 20283 16941
rect 20221 16681 20283 16693
rect 20313 16941 20379 16953
rect 20313 16693 20329 16941
rect 20363 16693 20379 16941
rect 20313 16681 20379 16693
rect 20409 16941 20475 16953
rect 20409 16693 20425 16941
rect 20459 16693 20475 16941
rect 20409 16681 20475 16693
rect 20505 16941 20571 16953
rect 20505 16693 20521 16941
rect 20555 16693 20571 16941
rect 20505 16681 20571 16693
rect 20601 16941 20667 16953
rect 20601 16693 20617 16941
rect 20651 16693 20667 16941
rect 20601 16681 20667 16693
rect 20697 16941 20763 16953
rect 20697 16693 20713 16941
rect 20747 16693 20763 16941
rect 20697 16681 20763 16693
rect 20793 16941 20859 16953
rect 20793 16693 20809 16941
rect 20843 16693 20859 16941
rect 20793 16681 20859 16693
rect 20889 16941 20955 16953
rect 20889 16693 20905 16941
rect 20939 16693 20955 16941
rect 20889 16681 20955 16693
rect 20985 16941 21051 16953
rect 20985 16693 21001 16941
rect 21035 16693 21051 16941
rect 20985 16681 21051 16693
rect 21081 16941 21147 16953
rect 21081 16693 21097 16941
rect 21131 16693 21147 16941
rect 21081 16681 21147 16693
rect 21177 16941 21239 16953
rect 21177 16693 21193 16941
rect 21227 16693 21239 16941
rect 21177 16681 21239 16693
rect 7291 15141 7353 15153
rect 7291 14893 7303 15141
rect 7337 14893 7353 15141
rect 7291 14881 7353 14893
rect 7383 15141 7449 15153
rect 7383 14893 7399 15141
rect 7433 14893 7449 15141
rect 7383 14881 7449 14893
rect 7479 15141 7545 15153
rect 7479 14893 7495 15141
rect 7529 14893 7545 15141
rect 7479 14881 7545 14893
rect 7575 15141 7641 15153
rect 7575 14893 7591 15141
rect 7625 14893 7641 15141
rect 7575 14881 7641 14893
rect 7671 15141 7737 15153
rect 7671 14893 7687 15141
rect 7721 14893 7737 15141
rect 7671 14881 7737 14893
rect 7767 15141 7833 15153
rect 7767 14893 7783 15141
rect 7817 14893 7833 15141
rect 7767 14881 7833 14893
rect 7863 15141 7929 15153
rect 7863 14893 7879 15141
rect 7913 14893 7929 15141
rect 7863 14881 7929 14893
rect 7959 15141 8025 15153
rect 7959 14893 7975 15141
rect 8009 14893 8025 15141
rect 7959 14881 8025 14893
rect 8055 15141 8121 15153
rect 8055 14893 8071 15141
rect 8105 14893 8121 15141
rect 8055 14881 8121 14893
rect 8151 15141 8217 15153
rect 8151 14893 8167 15141
rect 8201 14893 8217 15141
rect 8151 14881 8217 14893
rect 8247 15141 8309 15153
rect 8247 14893 8263 15141
rect 8297 14893 8309 15141
rect 8247 14881 8309 14893
rect 20221 15141 20283 15153
rect 20221 14893 20233 15141
rect 20267 14893 20283 15141
rect 20221 14881 20283 14893
rect 20313 15141 20379 15153
rect 20313 14893 20329 15141
rect 20363 14893 20379 15141
rect 20313 14881 20379 14893
rect 20409 15141 20475 15153
rect 20409 14893 20425 15141
rect 20459 14893 20475 15141
rect 20409 14881 20475 14893
rect 20505 15141 20571 15153
rect 20505 14893 20521 15141
rect 20555 14893 20571 15141
rect 20505 14881 20571 14893
rect 20601 15141 20667 15153
rect 20601 14893 20617 15141
rect 20651 14893 20667 15141
rect 20601 14881 20667 14893
rect 20697 15141 20763 15153
rect 20697 14893 20713 15141
rect 20747 14893 20763 15141
rect 20697 14881 20763 14893
rect 20793 15141 20859 15153
rect 20793 14893 20809 15141
rect 20843 14893 20859 15141
rect 20793 14881 20859 14893
rect 20889 15141 20955 15153
rect 20889 14893 20905 15141
rect 20939 14893 20955 15141
rect 20889 14881 20955 14893
rect 20985 15141 21051 15153
rect 20985 14893 21001 15141
rect 21035 14893 21051 15141
rect 20985 14881 21051 14893
rect 21081 15141 21147 15153
rect 21081 14893 21097 15141
rect 21131 14893 21147 15141
rect 21081 14881 21147 14893
rect 21177 15141 21239 15153
rect 21177 14893 21193 15141
rect 21227 14893 21239 15141
rect 21177 14881 21239 14893
rect 7291 13341 7353 13353
rect 7291 13093 7303 13341
rect 7337 13093 7353 13341
rect 7291 13081 7353 13093
rect 7383 13341 7449 13353
rect 7383 13093 7399 13341
rect 7433 13093 7449 13341
rect 7383 13081 7449 13093
rect 7479 13341 7545 13353
rect 7479 13093 7495 13341
rect 7529 13093 7545 13341
rect 7479 13081 7545 13093
rect 7575 13341 7641 13353
rect 7575 13093 7591 13341
rect 7625 13093 7641 13341
rect 7575 13081 7641 13093
rect 7671 13341 7737 13353
rect 7671 13093 7687 13341
rect 7721 13093 7737 13341
rect 7671 13081 7737 13093
rect 7767 13341 7833 13353
rect 7767 13093 7783 13341
rect 7817 13093 7833 13341
rect 7767 13081 7833 13093
rect 7863 13341 7929 13353
rect 7863 13093 7879 13341
rect 7913 13093 7929 13341
rect 7863 13081 7929 13093
rect 7959 13341 8025 13353
rect 7959 13093 7975 13341
rect 8009 13093 8025 13341
rect 7959 13081 8025 13093
rect 8055 13341 8121 13353
rect 8055 13093 8071 13341
rect 8105 13093 8121 13341
rect 8055 13081 8121 13093
rect 8151 13341 8217 13353
rect 8151 13093 8167 13341
rect 8201 13093 8217 13341
rect 8151 13081 8217 13093
rect 8247 13341 8309 13353
rect 8247 13093 8263 13341
rect 8297 13093 8309 13341
rect 8247 13081 8309 13093
rect 20221 13341 20283 13353
rect 20221 13093 20233 13341
rect 20267 13093 20283 13341
rect 20221 13081 20283 13093
rect 20313 13341 20379 13353
rect 20313 13093 20329 13341
rect 20363 13093 20379 13341
rect 20313 13081 20379 13093
rect 20409 13341 20475 13353
rect 20409 13093 20425 13341
rect 20459 13093 20475 13341
rect 20409 13081 20475 13093
rect 20505 13341 20571 13353
rect 20505 13093 20521 13341
rect 20555 13093 20571 13341
rect 20505 13081 20571 13093
rect 20601 13341 20667 13353
rect 20601 13093 20617 13341
rect 20651 13093 20667 13341
rect 20601 13081 20667 13093
rect 20697 13341 20763 13353
rect 20697 13093 20713 13341
rect 20747 13093 20763 13341
rect 20697 13081 20763 13093
rect 20793 13341 20859 13353
rect 20793 13093 20809 13341
rect 20843 13093 20859 13341
rect 20793 13081 20859 13093
rect 20889 13341 20955 13353
rect 20889 13093 20905 13341
rect 20939 13093 20955 13341
rect 20889 13081 20955 13093
rect 20985 13341 21051 13353
rect 20985 13093 21001 13341
rect 21035 13093 21051 13341
rect 20985 13081 21051 13093
rect 21081 13341 21147 13353
rect 21081 13093 21097 13341
rect 21131 13093 21147 13341
rect 21081 13081 21147 13093
rect 21177 13341 21239 13353
rect 21177 13093 21193 13341
rect 21227 13093 21239 13341
rect 21177 13081 21239 13093
rect 7291 11541 7353 11553
rect 7291 11293 7303 11541
rect 7337 11293 7353 11541
rect 7291 11281 7353 11293
rect 7383 11541 7449 11553
rect 7383 11293 7399 11541
rect 7433 11293 7449 11541
rect 7383 11281 7449 11293
rect 7479 11541 7545 11553
rect 7479 11293 7495 11541
rect 7529 11293 7545 11541
rect 7479 11281 7545 11293
rect 7575 11541 7641 11553
rect 7575 11293 7591 11541
rect 7625 11293 7641 11541
rect 7575 11281 7641 11293
rect 7671 11541 7737 11553
rect 7671 11293 7687 11541
rect 7721 11293 7737 11541
rect 7671 11281 7737 11293
rect 7767 11541 7833 11553
rect 7767 11293 7783 11541
rect 7817 11293 7833 11541
rect 7767 11281 7833 11293
rect 7863 11541 7929 11553
rect 7863 11293 7879 11541
rect 7913 11293 7929 11541
rect 7863 11281 7929 11293
rect 7959 11541 8025 11553
rect 7959 11293 7975 11541
rect 8009 11293 8025 11541
rect 7959 11281 8025 11293
rect 8055 11541 8121 11553
rect 8055 11293 8071 11541
rect 8105 11293 8121 11541
rect 8055 11281 8121 11293
rect 8151 11541 8217 11553
rect 8151 11293 8167 11541
rect 8201 11293 8217 11541
rect 8151 11281 8217 11293
rect 8247 11541 8309 11553
rect 8247 11293 8263 11541
rect 8297 11293 8309 11541
rect 8247 11281 8309 11293
rect 20221 11541 20283 11553
rect 20221 11293 20233 11541
rect 20267 11293 20283 11541
rect 20221 11281 20283 11293
rect 20313 11541 20379 11553
rect 20313 11293 20329 11541
rect 20363 11293 20379 11541
rect 20313 11281 20379 11293
rect 20409 11541 20475 11553
rect 20409 11293 20425 11541
rect 20459 11293 20475 11541
rect 20409 11281 20475 11293
rect 20505 11541 20571 11553
rect 20505 11293 20521 11541
rect 20555 11293 20571 11541
rect 20505 11281 20571 11293
rect 20601 11541 20667 11553
rect 20601 11293 20617 11541
rect 20651 11293 20667 11541
rect 20601 11281 20667 11293
rect 20697 11541 20763 11553
rect 20697 11293 20713 11541
rect 20747 11293 20763 11541
rect 20697 11281 20763 11293
rect 20793 11541 20859 11553
rect 20793 11293 20809 11541
rect 20843 11293 20859 11541
rect 20793 11281 20859 11293
rect 20889 11541 20955 11553
rect 20889 11293 20905 11541
rect 20939 11293 20955 11541
rect 20889 11281 20955 11293
rect 20985 11541 21051 11553
rect 20985 11293 21001 11541
rect 21035 11293 21051 11541
rect 20985 11281 21051 11293
rect 21081 11541 21147 11553
rect 21081 11293 21097 11541
rect 21131 11293 21147 11541
rect 21081 11281 21147 11293
rect 21177 11541 21239 11553
rect 21177 11293 21193 11541
rect 21227 11293 21239 11541
rect 21177 11281 21239 11293
rect 7291 9741 7353 9753
rect 7291 9493 7303 9741
rect 7337 9493 7353 9741
rect 7291 9481 7353 9493
rect 7383 9741 7449 9753
rect 7383 9493 7399 9741
rect 7433 9493 7449 9741
rect 7383 9481 7449 9493
rect 7479 9741 7545 9753
rect 7479 9493 7495 9741
rect 7529 9493 7545 9741
rect 7479 9481 7545 9493
rect 7575 9741 7641 9753
rect 7575 9493 7591 9741
rect 7625 9493 7641 9741
rect 7575 9481 7641 9493
rect 7671 9741 7737 9753
rect 7671 9493 7687 9741
rect 7721 9493 7737 9741
rect 7671 9481 7737 9493
rect 7767 9741 7833 9753
rect 7767 9493 7783 9741
rect 7817 9493 7833 9741
rect 7767 9481 7833 9493
rect 7863 9741 7929 9753
rect 7863 9493 7879 9741
rect 7913 9493 7929 9741
rect 7863 9481 7929 9493
rect 7959 9741 8025 9753
rect 7959 9493 7975 9741
rect 8009 9493 8025 9741
rect 7959 9481 8025 9493
rect 8055 9741 8121 9753
rect 8055 9493 8071 9741
rect 8105 9493 8121 9741
rect 8055 9481 8121 9493
rect 8151 9741 8217 9753
rect 8151 9493 8167 9741
rect 8201 9493 8217 9741
rect 8151 9481 8217 9493
rect 8247 9741 8309 9753
rect 8247 9493 8263 9741
rect 8297 9493 8309 9741
rect 8247 9481 8309 9493
rect 20221 9741 20283 9753
rect 20221 9493 20233 9741
rect 20267 9493 20283 9741
rect 20221 9481 20283 9493
rect 20313 9741 20379 9753
rect 20313 9493 20329 9741
rect 20363 9493 20379 9741
rect 20313 9481 20379 9493
rect 20409 9741 20475 9753
rect 20409 9493 20425 9741
rect 20459 9493 20475 9741
rect 20409 9481 20475 9493
rect 20505 9741 20571 9753
rect 20505 9493 20521 9741
rect 20555 9493 20571 9741
rect 20505 9481 20571 9493
rect 20601 9741 20667 9753
rect 20601 9493 20617 9741
rect 20651 9493 20667 9741
rect 20601 9481 20667 9493
rect 20697 9741 20763 9753
rect 20697 9493 20713 9741
rect 20747 9493 20763 9741
rect 20697 9481 20763 9493
rect 20793 9741 20859 9753
rect 20793 9493 20809 9741
rect 20843 9493 20859 9741
rect 20793 9481 20859 9493
rect 20889 9741 20955 9753
rect 20889 9493 20905 9741
rect 20939 9493 20955 9741
rect 20889 9481 20955 9493
rect 20985 9741 21051 9753
rect 20985 9493 21001 9741
rect 21035 9493 21051 9741
rect 20985 9481 21051 9493
rect 21081 9741 21147 9753
rect 21081 9493 21097 9741
rect 21131 9493 21147 9741
rect 21081 9481 21147 9493
rect 21177 9741 21239 9753
rect 21177 9493 21193 9741
rect 21227 9493 21239 9741
rect 21177 9481 21239 9493
rect 7544 6597 7602 6609
rect 7544 6341 7556 6597
rect 7590 6341 7602 6597
rect 7544 6329 7602 6341
rect 7722 6597 7780 6609
rect 7722 6341 7734 6597
rect 7768 6341 7780 6597
rect 7722 6329 7780 6341
rect 7900 6597 7958 6609
rect 7900 6341 7912 6597
rect 7946 6341 7958 6597
rect 7900 6329 7958 6341
rect 8078 6597 8136 6609
rect 8078 6341 8090 6597
rect 8124 6341 8136 6597
rect 8078 6329 8136 6341
rect 8256 6597 8314 6609
rect 8256 6341 8268 6597
rect 8302 6341 8314 6597
rect 8256 6329 8314 6341
rect 8434 6597 8492 6609
rect 8434 6341 8446 6597
rect 8480 6341 8492 6597
rect 8434 6329 8492 6341
rect 8612 6597 8670 6609
rect 8612 6341 8624 6597
rect 8658 6341 8670 6597
rect 8612 6329 8670 6341
rect 8790 6597 8848 6609
rect 8790 6341 8802 6597
rect 8836 6341 8848 6597
rect 8790 6329 8848 6341
rect 8968 6597 9026 6609
rect 8968 6341 8980 6597
rect 9014 6341 9026 6597
rect 8968 6329 9026 6341
rect 9146 6597 9204 6609
rect 9146 6341 9158 6597
rect 9192 6341 9204 6597
rect 9146 6329 9204 6341
rect 9324 6597 9382 6609
rect 9324 6341 9336 6597
rect 9370 6341 9382 6597
rect 9324 6329 9382 6341
rect 9502 6597 9560 6609
rect 9502 6341 9514 6597
rect 9548 6341 9560 6597
rect 9502 6329 9560 6341
rect 9680 6597 9738 6609
rect 9680 6341 9692 6597
rect 9726 6341 9738 6597
rect 9680 6329 9738 6341
rect 9858 6597 9916 6609
rect 9858 6341 9870 6597
rect 9904 6341 9916 6597
rect 9858 6329 9916 6341
rect 10036 6597 10094 6609
rect 10036 6341 10048 6597
rect 10082 6341 10094 6597
rect 10036 6329 10094 6341
rect 10230 6597 10288 6609
rect 10230 6341 10242 6597
rect 10276 6341 10288 6597
rect 10230 6329 10288 6341
rect 10408 6597 10466 6609
rect 10408 6341 10420 6597
rect 10454 6341 10466 6597
rect 10408 6329 10466 6341
rect 10586 6597 10644 6609
rect 10586 6341 10598 6597
rect 10632 6341 10644 6597
rect 10586 6329 10644 6341
rect 10764 6597 10822 6609
rect 10764 6341 10776 6597
rect 10810 6341 10822 6597
rect 10764 6329 10822 6341
rect 10942 6597 11000 6609
rect 10942 6341 10954 6597
rect 10988 6341 11000 6597
rect 10942 6329 11000 6341
rect 11120 6597 11178 6609
rect 11120 6341 11132 6597
rect 11166 6341 11178 6597
rect 11120 6329 11178 6341
rect 11298 6597 11356 6609
rect 11298 6341 11310 6597
rect 11344 6341 11356 6597
rect 11298 6329 11356 6341
rect 11476 6597 11534 6609
rect 11476 6341 11488 6597
rect 11522 6341 11534 6597
rect 11476 6329 11534 6341
rect 11654 6597 11712 6609
rect 11654 6341 11666 6597
rect 11700 6341 11712 6597
rect 11654 6329 11712 6341
rect 11832 6597 11890 6609
rect 11832 6341 11844 6597
rect 11878 6341 11890 6597
rect 11832 6329 11890 6341
rect 12010 6597 12068 6609
rect 12010 6341 12022 6597
rect 12056 6341 12068 6597
rect 12010 6329 12068 6341
rect 12188 6597 12246 6609
rect 12188 6341 12200 6597
rect 12234 6341 12246 6597
rect 12188 6329 12246 6341
rect 12366 6597 12424 6609
rect 12366 6341 12378 6597
rect 12412 6341 12424 6597
rect 12366 6329 12424 6341
rect 12544 6597 12602 6609
rect 12544 6341 12556 6597
rect 12590 6341 12602 6597
rect 12544 6329 12602 6341
rect 12722 6597 12780 6609
rect 12722 6341 12734 6597
rect 12768 6341 12780 6597
rect 12722 6329 12780 6341
rect 7544 6019 7602 6031
rect 7544 5763 7556 6019
rect 7590 5763 7602 6019
rect 7544 5751 7602 5763
rect 7722 6019 7780 6031
rect 7722 5763 7734 6019
rect 7768 5763 7780 6019
rect 7722 5751 7780 5763
rect 7900 6019 7958 6031
rect 7900 5763 7912 6019
rect 7946 5763 7958 6019
rect 7900 5751 7958 5763
rect 8078 6019 8136 6031
rect 8078 5763 8090 6019
rect 8124 5763 8136 6019
rect 8078 5751 8136 5763
rect 8256 6019 8314 6031
rect 8256 5763 8268 6019
rect 8302 5763 8314 6019
rect 8256 5751 8314 5763
rect 8434 6019 8492 6031
rect 8434 5763 8446 6019
rect 8480 5763 8492 6019
rect 8434 5751 8492 5763
rect 8612 6019 8670 6031
rect 8612 5763 8624 6019
rect 8658 5763 8670 6019
rect 8612 5751 8670 5763
rect 8790 6019 8848 6031
rect 8790 5763 8802 6019
rect 8836 5763 8848 6019
rect 8790 5751 8848 5763
rect 8968 6019 9026 6031
rect 8968 5763 8980 6019
rect 9014 5763 9026 6019
rect 8968 5751 9026 5763
rect 9146 6019 9204 6031
rect 9146 5763 9158 6019
rect 9192 5763 9204 6019
rect 9146 5751 9204 5763
rect 9324 6019 9382 6031
rect 9324 5763 9336 6019
rect 9370 5763 9382 6019
rect 9324 5751 9382 5763
rect 9502 6019 9560 6031
rect 9502 5763 9514 6019
rect 9548 5763 9560 6019
rect 9502 5751 9560 5763
rect 9680 6019 9738 6031
rect 9680 5763 9692 6019
rect 9726 5763 9738 6019
rect 9680 5751 9738 5763
rect 9858 6019 9916 6031
rect 9858 5763 9870 6019
rect 9904 5763 9916 6019
rect 9858 5751 9916 5763
rect 10036 6019 10094 6031
rect 10036 5763 10048 6019
rect 10082 5763 10094 6019
rect 10036 5751 10094 5763
rect 10230 6020 10288 6032
rect 10230 5764 10242 6020
rect 10276 5764 10288 6020
rect 10230 5752 10288 5764
rect 10408 6020 10466 6032
rect 10408 5764 10420 6020
rect 10454 5764 10466 6020
rect 10408 5752 10466 5764
rect 10586 6020 10644 6032
rect 10586 5764 10598 6020
rect 10632 5764 10644 6020
rect 10586 5752 10644 5764
rect 10764 6020 10822 6032
rect 10764 5764 10776 6020
rect 10810 5764 10822 6020
rect 10764 5752 10822 5764
rect 10942 6020 11000 6032
rect 10942 5764 10954 6020
rect 10988 5764 11000 6020
rect 10942 5752 11000 5764
rect 11120 6020 11178 6032
rect 11120 5764 11132 6020
rect 11166 5764 11178 6020
rect 11120 5752 11178 5764
rect 11298 6020 11356 6032
rect 11298 5764 11310 6020
rect 11344 5764 11356 6020
rect 11298 5752 11356 5764
rect 11476 6020 11534 6032
rect 11476 5764 11488 6020
rect 11522 5764 11534 6020
rect 11476 5752 11534 5764
rect 11654 6020 11712 6032
rect 11654 5764 11666 6020
rect 11700 5764 11712 6020
rect 11654 5752 11712 5764
rect 11832 6020 11890 6032
rect 11832 5764 11844 6020
rect 11878 5764 11890 6020
rect 11832 5752 11890 5764
rect 12010 6020 12068 6032
rect 12010 5764 12022 6020
rect 12056 5764 12068 6020
rect 12010 5752 12068 5764
rect 12188 6020 12246 6032
rect 12188 5764 12200 6020
rect 12234 5764 12246 6020
rect 12188 5752 12246 5764
rect 12366 6020 12424 6032
rect 12366 5764 12378 6020
rect 12412 5764 12424 6020
rect 12366 5752 12424 5764
rect 12544 6020 12602 6032
rect 12544 5764 12556 6020
rect 12590 5764 12602 6020
rect 12544 5752 12602 5764
rect 12722 6020 12780 6032
rect 12722 5764 12734 6020
rect 12768 5764 12780 6020
rect 12722 5752 12780 5764
rect 14684 6666 14742 6678
rect 14684 6410 14696 6666
rect 14730 6410 14742 6666
rect 14684 6398 14742 6410
rect 14862 6666 14920 6678
rect 14862 6410 14874 6666
rect 14908 6410 14920 6666
rect 14862 6398 14920 6410
rect 15040 6666 15098 6678
rect 15040 6410 15052 6666
rect 15086 6410 15098 6666
rect 15040 6398 15098 6410
rect 15218 6666 15276 6678
rect 15218 6410 15230 6666
rect 15264 6410 15276 6666
rect 15218 6398 15276 6410
rect 15396 6666 15454 6678
rect 15396 6410 15408 6666
rect 15442 6410 15454 6666
rect 15396 6398 15454 6410
rect 15574 6666 15632 6678
rect 15574 6410 15586 6666
rect 15620 6410 15632 6666
rect 15574 6398 15632 6410
rect 15752 6666 15810 6678
rect 15752 6410 15764 6666
rect 15798 6410 15810 6666
rect 15752 6398 15810 6410
rect 15930 6666 15988 6678
rect 15930 6410 15942 6666
rect 15976 6410 15988 6666
rect 15930 6398 15988 6410
rect 16108 6666 16166 6678
rect 16108 6410 16120 6666
rect 16154 6410 16166 6666
rect 16108 6398 16166 6410
rect 16884 6666 16942 6678
rect 16884 6410 16896 6666
rect 16930 6410 16942 6666
rect 16884 6398 16942 6410
rect 17062 6666 17120 6678
rect 17062 6410 17074 6666
rect 17108 6410 17120 6666
rect 17062 6398 17120 6410
rect 17240 6666 17298 6678
rect 17240 6410 17252 6666
rect 17286 6410 17298 6666
rect 17240 6398 17298 6410
rect 17418 6666 17476 6678
rect 17418 6410 17430 6666
rect 17464 6410 17476 6666
rect 17418 6398 17476 6410
rect 17596 6666 17654 6678
rect 17596 6410 17608 6666
rect 17642 6410 17654 6666
rect 17596 6398 17654 6410
rect 17774 6666 17832 6678
rect 17774 6410 17786 6666
rect 17820 6410 17832 6666
rect 17774 6398 17832 6410
rect 17952 6666 18010 6678
rect 17952 6410 17964 6666
rect 17998 6410 18010 6666
rect 17952 6398 18010 6410
rect 18130 6666 18188 6678
rect 18130 6410 18142 6666
rect 18176 6410 18188 6666
rect 18130 6398 18188 6410
rect 18308 6666 18366 6678
rect 18308 6410 18320 6666
rect 18354 6410 18366 6666
rect 18308 6398 18366 6410
rect 19084 6666 19142 6678
rect 19084 6410 19096 6666
rect 19130 6410 19142 6666
rect 19084 6398 19142 6410
rect 19262 6666 19320 6678
rect 19262 6410 19274 6666
rect 19308 6410 19320 6666
rect 19262 6398 19320 6410
rect 19440 6666 19498 6678
rect 19440 6410 19452 6666
rect 19486 6410 19498 6666
rect 19440 6398 19498 6410
rect 19618 6666 19676 6678
rect 19618 6410 19630 6666
rect 19664 6410 19676 6666
rect 19618 6398 19676 6410
rect 19796 6666 19854 6678
rect 19796 6410 19808 6666
rect 19842 6410 19854 6666
rect 19796 6398 19854 6410
rect 19974 6666 20032 6678
rect 19974 6410 19986 6666
rect 20020 6410 20032 6666
rect 19974 6398 20032 6410
rect 20152 6666 20210 6678
rect 20152 6410 20164 6666
rect 20198 6410 20210 6666
rect 20152 6398 20210 6410
rect 20330 6666 20388 6678
rect 20330 6410 20342 6666
rect 20376 6410 20388 6666
rect 20330 6398 20388 6410
rect 20508 6666 20566 6678
rect 20508 6410 20520 6666
rect 20554 6410 20566 6666
rect 20508 6398 20566 6410
rect 14685 5899 14743 5911
rect 14685 5643 14697 5899
rect 14731 5643 14743 5899
rect 14685 5631 14743 5643
rect 14863 5899 14921 5911
rect 14863 5643 14875 5899
rect 14909 5643 14921 5899
rect 14863 5631 14921 5643
rect 15041 5899 15099 5911
rect 15041 5643 15053 5899
rect 15087 5643 15099 5899
rect 15041 5631 15099 5643
rect 15219 5899 15277 5911
rect 15219 5643 15231 5899
rect 15265 5643 15277 5899
rect 15219 5631 15277 5643
rect 15397 5899 15455 5911
rect 15397 5643 15409 5899
rect 15443 5643 15455 5899
rect 15397 5631 15455 5643
rect 15575 5899 15633 5911
rect 15575 5643 15587 5899
rect 15621 5643 15633 5899
rect 15575 5631 15633 5643
rect 15753 5899 15811 5911
rect 15753 5643 15765 5899
rect 15799 5643 15811 5899
rect 15753 5631 15811 5643
rect 15931 5899 15989 5911
rect 15931 5643 15943 5899
rect 15977 5643 15989 5899
rect 15931 5631 15989 5643
rect 16109 5899 16167 5911
rect 16109 5643 16121 5899
rect 16155 5643 16167 5899
rect 16109 5631 16167 5643
rect 16885 5899 16943 5911
rect 16885 5643 16897 5899
rect 16931 5643 16943 5899
rect 16885 5631 16943 5643
rect 17063 5899 17121 5911
rect 17063 5643 17075 5899
rect 17109 5643 17121 5899
rect 17063 5631 17121 5643
rect 17241 5899 17299 5911
rect 17241 5643 17253 5899
rect 17287 5643 17299 5899
rect 17241 5631 17299 5643
rect 17419 5899 17477 5911
rect 17419 5643 17431 5899
rect 17465 5643 17477 5899
rect 17419 5631 17477 5643
rect 17597 5899 17655 5911
rect 17597 5643 17609 5899
rect 17643 5643 17655 5899
rect 17597 5631 17655 5643
rect 17775 5899 17833 5911
rect 17775 5643 17787 5899
rect 17821 5643 17833 5899
rect 17775 5631 17833 5643
rect 17953 5899 18011 5911
rect 17953 5643 17965 5899
rect 17999 5643 18011 5899
rect 17953 5631 18011 5643
rect 18131 5899 18189 5911
rect 18131 5643 18143 5899
rect 18177 5643 18189 5899
rect 18131 5631 18189 5643
rect 18309 5899 18367 5911
rect 18309 5643 18321 5899
rect 18355 5643 18367 5899
rect 18309 5631 18367 5643
rect 19085 5899 19143 5911
rect 19085 5643 19097 5899
rect 19131 5643 19143 5899
rect 19085 5631 19143 5643
rect 19263 5899 19321 5911
rect 19263 5643 19275 5899
rect 19309 5643 19321 5899
rect 19263 5631 19321 5643
rect 19441 5899 19499 5911
rect 19441 5643 19453 5899
rect 19487 5643 19499 5899
rect 19441 5631 19499 5643
rect 19619 5899 19677 5911
rect 19619 5643 19631 5899
rect 19665 5643 19677 5899
rect 19619 5631 19677 5643
rect 19797 5899 19855 5911
rect 19797 5643 19809 5899
rect 19843 5643 19855 5899
rect 19797 5631 19855 5643
rect 19975 5899 20033 5911
rect 19975 5643 19987 5899
rect 20021 5643 20033 5899
rect 19975 5631 20033 5643
rect 20153 5899 20211 5911
rect 20153 5643 20165 5899
rect 20199 5643 20211 5899
rect 20153 5631 20211 5643
rect 20331 5899 20389 5911
rect 20331 5643 20343 5899
rect 20377 5643 20389 5899
rect 20331 5631 20389 5643
rect 20509 5899 20567 5911
rect 20509 5643 20521 5899
rect 20555 5643 20567 5899
rect 20509 5631 20567 5643
rect 7900 5139 7958 5151
rect 7900 4883 7912 5139
rect 7946 4883 7958 5139
rect 7900 4871 7958 4883
rect 8078 5139 8136 5151
rect 8078 4883 8090 5139
rect 8124 4883 8136 5139
rect 8078 4871 8136 4883
rect 8256 5139 8314 5151
rect 8256 4883 8268 5139
rect 8302 4883 8314 5139
rect 8256 4871 8314 4883
rect 8434 5139 8492 5151
rect 8434 4883 8446 5139
rect 8480 4883 8492 5139
rect 8434 4871 8492 4883
rect 8612 5139 8670 5151
rect 8612 4883 8624 5139
rect 8658 4883 8670 5139
rect 8612 4871 8670 4883
rect 8790 5139 8848 5151
rect 8790 4883 8802 5139
rect 8836 4883 8848 5139
rect 8790 4871 8848 4883
rect 8968 5139 9026 5151
rect 8968 4883 8980 5139
rect 9014 4883 9026 5139
rect 8968 4871 9026 4883
rect 9146 5139 9204 5151
rect 9146 4883 9158 5139
rect 9192 4883 9204 5139
rect 9146 4871 9204 4883
rect 9324 5139 9382 5151
rect 9324 4883 9336 5139
rect 9370 4883 9382 5139
rect 9324 4871 9382 4883
rect 9502 5139 9560 5151
rect 9502 4883 9514 5139
rect 9548 4883 9560 5139
rect 9502 4871 9560 4883
rect 9680 5139 9738 5151
rect 9680 4883 9692 5139
rect 9726 4883 9738 5139
rect 9680 4871 9738 4883
rect 9858 5139 9916 5151
rect 9858 4883 9870 5139
rect 9904 4883 9916 5139
rect 9858 4871 9916 4883
rect 10036 5139 10094 5151
rect 10036 4883 10048 5139
rect 10082 4883 10094 5139
rect 10036 4871 10094 4883
rect 10230 5139 10288 5151
rect 10230 4883 10242 5139
rect 10276 4883 10288 5139
rect 10230 4871 10288 4883
rect 10408 5139 10466 5151
rect 10408 4883 10420 5139
rect 10454 4883 10466 5139
rect 10408 4871 10466 4883
rect 10586 5139 10644 5151
rect 10586 4883 10598 5139
rect 10632 4883 10644 5139
rect 10586 4871 10644 4883
rect 10764 5139 10822 5151
rect 10764 4883 10776 5139
rect 10810 4883 10822 5139
rect 10764 4871 10822 4883
rect 10942 5139 11000 5151
rect 10942 4883 10954 5139
rect 10988 4883 11000 5139
rect 10942 4871 11000 4883
rect 11120 5139 11178 5151
rect 11120 4883 11132 5139
rect 11166 4883 11178 5139
rect 11120 4871 11178 4883
rect 11298 5139 11356 5151
rect 11298 4883 11310 5139
rect 11344 4883 11356 5139
rect 11298 4871 11356 4883
rect 11476 5139 11534 5151
rect 11476 4883 11488 5139
rect 11522 4883 11534 5139
rect 11476 4871 11534 4883
rect 11654 5139 11712 5151
rect 11654 4883 11666 5139
rect 11700 4883 11712 5139
rect 11654 4871 11712 4883
rect 11832 5139 11890 5151
rect 11832 4883 11844 5139
rect 11878 4883 11890 5139
rect 11832 4871 11890 4883
rect 12010 5139 12068 5151
rect 12010 4883 12022 5139
rect 12056 4883 12068 5139
rect 12010 4871 12068 4883
rect 12188 5139 12246 5151
rect 12188 4883 12200 5139
rect 12234 4883 12246 5139
rect 12188 4871 12246 4883
rect 12366 5139 12424 5151
rect 12366 4883 12378 5139
rect 12412 4883 12424 5139
rect 12366 4871 12424 4883
rect 7900 4569 7958 4581
rect 7900 4313 7912 4569
rect 7946 4313 7958 4569
rect 7900 4301 7958 4313
rect 8078 4569 8136 4581
rect 8078 4313 8090 4569
rect 8124 4313 8136 4569
rect 8078 4301 8136 4313
rect 8256 4569 8314 4581
rect 8256 4313 8268 4569
rect 8302 4313 8314 4569
rect 8256 4301 8314 4313
rect 8434 4569 8492 4581
rect 8434 4313 8446 4569
rect 8480 4313 8492 4569
rect 8434 4301 8492 4313
rect 8612 4569 8670 4581
rect 8612 4313 8624 4569
rect 8658 4313 8670 4569
rect 8612 4301 8670 4313
rect 8790 4569 8848 4581
rect 8790 4313 8802 4569
rect 8836 4313 8848 4569
rect 8790 4301 8848 4313
rect 8968 4569 9026 4581
rect 8968 4313 8980 4569
rect 9014 4313 9026 4569
rect 8968 4301 9026 4313
rect 9146 4569 9204 4581
rect 9146 4313 9158 4569
rect 9192 4313 9204 4569
rect 9146 4301 9204 4313
rect 9324 4569 9382 4581
rect 9324 4313 9336 4569
rect 9370 4313 9382 4569
rect 9324 4301 9382 4313
rect 9502 4569 9560 4581
rect 9502 4313 9514 4569
rect 9548 4313 9560 4569
rect 9502 4301 9560 4313
rect 9680 4569 9738 4581
rect 9680 4313 9692 4569
rect 9726 4313 9738 4569
rect 9680 4301 9738 4313
rect 9858 4569 9916 4581
rect 9858 4313 9870 4569
rect 9904 4313 9916 4569
rect 9858 4301 9916 4313
rect 10036 4569 10094 4581
rect 10036 4313 10048 4569
rect 10082 4313 10094 4569
rect 10036 4301 10094 4313
rect 10230 4569 10288 4581
rect 10230 4313 10242 4569
rect 10276 4313 10288 4569
rect 10230 4301 10288 4313
rect 10408 4569 10466 4581
rect 10408 4313 10420 4569
rect 10454 4313 10466 4569
rect 10408 4301 10466 4313
rect 10586 4569 10644 4581
rect 10586 4313 10598 4569
rect 10632 4313 10644 4569
rect 10586 4301 10644 4313
rect 10764 4569 10822 4581
rect 10764 4313 10776 4569
rect 10810 4313 10822 4569
rect 10764 4301 10822 4313
rect 10942 4569 11000 4581
rect 10942 4313 10954 4569
rect 10988 4313 11000 4569
rect 10942 4301 11000 4313
rect 11120 4569 11178 4581
rect 11120 4313 11132 4569
rect 11166 4313 11178 4569
rect 11120 4301 11178 4313
rect 11298 4569 11356 4581
rect 11298 4313 11310 4569
rect 11344 4313 11356 4569
rect 11298 4301 11356 4313
rect 11476 4569 11534 4581
rect 11476 4313 11488 4569
rect 11522 4313 11534 4569
rect 11476 4301 11534 4313
rect 11654 4569 11712 4581
rect 11654 4313 11666 4569
rect 11700 4313 11712 4569
rect 11654 4301 11712 4313
rect 11832 4569 11890 4581
rect 11832 4313 11844 4569
rect 11878 4313 11890 4569
rect 11832 4301 11890 4313
rect 12010 4569 12068 4581
rect 12010 4313 12022 4569
rect 12056 4313 12068 4569
rect 12010 4301 12068 4313
rect 12188 4569 12246 4581
rect 12188 4313 12200 4569
rect 12234 4313 12246 4569
rect 12188 4301 12246 4313
rect 12366 4569 12424 4581
rect 12366 4313 12378 4569
rect 12412 4313 12424 4569
rect 12366 4301 12424 4313
<< ndiffc >>
rect 7303 18083 7337 18163
rect 7399 18083 7433 18163
rect 7495 18083 7529 18163
rect 7591 18083 7625 18163
rect 7687 18083 7721 18163
rect 7783 18083 7817 18163
rect 7879 18083 7913 18163
rect 7975 18083 8009 18163
rect 8071 18083 8105 18163
rect 8167 18083 8201 18163
rect 8263 18083 8297 18163
rect 20233 18083 20267 18163
rect 20329 18083 20363 18163
rect 20425 18083 20459 18163
rect 20521 18083 20555 18163
rect 20617 18083 20651 18163
rect 20713 18083 20747 18163
rect 20809 18083 20843 18163
rect 20905 18083 20939 18163
rect 21001 18083 21035 18163
rect 21097 18083 21131 18163
rect 21193 18083 21227 18163
rect 7303 16283 7337 16363
rect 7399 16283 7433 16363
rect 7495 16283 7529 16363
rect 7591 16283 7625 16363
rect 7687 16283 7721 16363
rect 7783 16283 7817 16363
rect 7879 16283 7913 16363
rect 7975 16283 8009 16363
rect 8071 16283 8105 16363
rect 8167 16283 8201 16363
rect 8263 16283 8297 16363
rect 20233 16283 20267 16363
rect 20329 16283 20363 16363
rect 20425 16283 20459 16363
rect 20521 16283 20555 16363
rect 20617 16283 20651 16363
rect 20713 16283 20747 16363
rect 20809 16283 20843 16363
rect 20905 16283 20939 16363
rect 21001 16283 21035 16363
rect 21097 16283 21131 16363
rect 21193 16283 21227 16363
rect 7303 14483 7337 14563
rect 7399 14483 7433 14563
rect 7495 14483 7529 14563
rect 7591 14483 7625 14563
rect 7687 14483 7721 14563
rect 7783 14483 7817 14563
rect 7879 14483 7913 14563
rect 7975 14483 8009 14563
rect 8071 14483 8105 14563
rect 8167 14483 8201 14563
rect 8263 14483 8297 14563
rect 20233 14483 20267 14563
rect 20329 14483 20363 14563
rect 20425 14483 20459 14563
rect 20521 14483 20555 14563
rect 20617 14483 20651 14563
rect 20713 14483 20747 14563
rect 20809 14483 20843 14563
rect 20905 14483 20939 14563
rect 21001 14483 21035 14563
rect 21097 14483 21131 14563
rect 21193 14483 21227 14563
rect 7303 12683 7337 12763
rect 7399 12683 7433 12763
rect 7495 12683 7529 12763
rect 7591 12683 7625 12763
rect 7687 12683 7721 12763
rect 7783 12683 7817 12763
rect 7879 12683 7913 12763
rect 7975 12683 8009 12763
rect 8071 12683 8105 12763
rect 8167 12683 8201 12763
rect 8263 12683 8297 12763
rect 20233 12683 20267 12763
rect 20329 12683 20363 12763
rect 20425 12683 20459 12763
rect 20521 12683 20555 12763
rect 20617 12683 20651 12763
rect 20713 12683 20747 12763
rect 20809 12683 20843 12763
rect 20905 12683 20939 12763
rect 21001 12683 21035 12763
rect 21097 12683 21131 12763
rect 21193 12683 21227 12763
rect 7303 10883 7337 10963
rect 7399 10883 7433 10963
rect 7495 10883 7529 10963
rect 7591 10883 7625 10963
rect 7687 10883 7721 10963
rect 7783 10883 7817 10963
rect 7879 10883 7913 10963
rect 7975 10883 8009 10963
rect 8071 10883 8105 10963
rect 8167 10883 8201 10963
rect 8263 10883 8297 10963
rect 20233 10883 20267 10963
rect 20329 10883 20363 10963
rect 20425 10883 20459 10963
rect 20521 10883 20555 10963
rect 20617 10883 20651 10963
rect 20713 10883 20747 10963
rect 20809 10883 20843 10963
rect 20905 10883 20939 10963
rect 21001 10883 21035 10963
rect 21097 10883 21131 10963
rect 21193 10883 21227 10963
rect 7303 9083 7337 9163
rect 7399 9083 7433 9163
rect 7495 9083 7529 9163
rect 7591 9083 7625 9163
rect 7687 9083 7721 9163
rect 7783 9083 7817 9163
rect 7879 9083 7913 9163
rect 7975 9083 8009 9163
rect 8071 9083 8105 9163
rect 8167 9083 8201 9163
rect 8263 9083 8297 9163
rect 20233 9083 20267 9163
rect 20329 9083 20363 9163
rect 20425 9083 20459 9163
rect 20521 9083 20555 9163
rect 20617 9083 20651 9163
rect 20713 9083 20747 9163
rect 20809 9083 20843 9163
rect 20905 9083 20939 9163
rect 21001 9083 21035 9163
rect 21097 9083 21131 9163
rect 21193 9083 21227 9163
rect 2050 4003 2084 4219
rect 2148 4003 2182 4219
rect 2262 4003 2296 4219
rect 2360 4003 2394 4219
rect 2474 4003 2508 4219
rect 2572 4003 2606 4219
rect 2686 4003 2720 4219
rect 2784 4003 2818 4219
rect 2898 4003 2932 4219
rect 2996 4003 3030 4219
rect 3110 4003 3144 4219
rect 3208 4003 3242 4219
rect 3322 4003 3356 4219
rect 3420 4003 3454 4219
rect 3534 4003 3568 4219
rect 3632 4003 3666 4219
rect 3830 4003 3864 4219
rect 3928 4003 3962 4219
rect 4042 4003 4076 4219
rect 4140 4003 4174 4219
rect 4254 4003 4288 4219
rect 4352 4003 4386 4219
rect 4466 4003 4500 4219
rect 4564 4003 4598 4219
rect 4678 4003 4712 4219
rect 4776 4003 4810 4219
rect 4890 4003 4924 4219
rect 4988 4003 5022 4219
rect 5102 4003 5136 4219
rect 5200 4003 5234 4219
rect 5314 4003 5348 4219
rect 5412 4003 5446 4219
rect 428 3183 462 3439
rect 606 3183 640 3439
rect 784 3183 818 3439
rect 962 3183 996 3439
rect 1140 3183 1174 3439
rect 1318 3183 1352 3439
rect 1496 3183 1530 3439
rect 1674 3183 1708 3439
rect 1852 3183 1886 3439
rect 2030 3183 2064 3439
rect 2208 3183 2242 3439
rect 2386 3183 2420 3439
rect 2564 3183 2598 3439
rect 2742 3183 2776 3439
rect 2920 3183 2954 3439
rect 3098 3183 3132 3439
rect 3276 3183 3310 3439
rect 3454 3183 3488 3439
rect 3632 3183 3666 3439
rect 3828 3183 3862 3439
rect 4006 3183 4040 3439
rect 4184 3183 4218 3439
rect 4362 3183 4396 3439
rect 4540 3183 4574 3439
rect 4718 3183 4752 3439
rect 4896 3183 4930 3439
rect 5074 3183 5108 3439
rect 5252 3183 5286 3439
rect 5430 3183 5464 3439
rect 5608 3183 5642 3439
rect 5786 3183 5820 3439
rect 5964 3183 5998 3439
rect 6142 3183 6176 3439
rect 6320 3183 6354 3439
rect 6498 3183 6532 3439
rect 6676 3183 6710 3439
rect 6854 3183 6888 3439
rect 7032 3183 7066 3439
rect 7557 3383 7591 3639
rect 7735 3383 7769 3639
rect 7913 3383 7947 3639
rect 8091 3383 8125 3639
rect 8269 3383 8303 3639
rect 8447 3383 8481 3639
rect 8625 3383 8659 3639
rect 8803 3383 8837 3639
rect 8981 3383 9015 3639
rect 9159 3383 9193 3639
rect 9337 3383 9371 3639
rect 9515 3383 9549 3639
rect 9693 3383 9727 3639
rect 9871 3383 9905 3639
rect 10049 3383 10083 3639
rect 10244 3383 10278 3639
rect 10422 3383 10456 3639
rect 10600 3383 10634 3639
rect 10778 3383 10812 3639
rect 10956 3383 10990 3639
rect 11134 3383 11168 3639
rect 11312 3383 11346 3639
rect 11490 3383 11524 3639
rect 11668 3383 11702 3639
rect 11846 3383 11880 3639
rect 12024 3383 12058 3639
rect 12202 3383 12236 3639
rect 12380 3383 12414 3639
rect 12558 3383 12592 3639
rect 12736 3383 12770 3639
rect 428 2683 462 2939
rect 606 2683 640 2939
rect 784 2683 818 2939
rect 962 2683 996 2939
rect 1140 2683 1174 2939
rect 1318 2683 1352 2939
rect 1496 2683 1530 2939
rect 1674 2683 1708 2939
rect 1852 2683 1886 2939
rect 2030 2683 2064 2939
rect 2208 2683 2242 2939
rect 2386 2683 2420 2939
rect 2564 2683 2598 2939
rect 2742 2683 2776 2939
rect 2920 2683 2954 2939
rect 3098 2683 3132 2939
rect 3276 2683 3310 2939
rect 3454 2683 3488 2939
rect 3632 2683 3666 2939
rect 3828 2683 3862 2939
rect 4006 2683 4040 2939
rect 4184 2683 4218 2939
rect 4362 2683 4396 2939
rect 4540 2683 4574 2939
rect 4718 2683 4752 2939
rect 4896 2683 4930 2939
rect 5074 2683 5108 2939
rect 5252 2683 5286 2939
rect 5430 2683 5464 2939
rect 5608 2683 5642 2939
rect 5786 2683 5820 2939
rect 5964 2683 5998 2939
rect 6142 2683 6176 2939
rect 6320 2683 6354 2939
rect 6498 2683 6532 2939
rect 6676 2683 6710 2939
rect 6854 2683 6888 2939
rect 7032 2683 7066 2939
rect 7557 2883 7591 3139
rect 7735 2883 7769 3139
rect 7913 2883 7947 3139
rect 8091 2883 8125 3139
rect 8269 2883 8303 3139
rect 8447 2883 8481 3139
rect 8625 2883 8659 3139
rect 8803 2883 8837 3139
rect 8981 2883 9015 3139
rect 9159 2883 9193 3139
rect 9337 2883 9371 3139
rect 9515 2883 9549 3139
rect 9693 2883 9727 3139
rect 9871 2883 9905 3139
rect 10049 2883 10083 3139
rect 10244 2883 10278 3139
rect 10422 2883 10456 3139
rect 10600 2883 10634 3139
rect 10778 2883 10812 3139
rect 10956 2883 10990 3139
rect 11134 2883 11168 3139
rect 11312 2883 11346 3139
rect 11490 2883 11524 3139
rect 11668 2883 11702 3139
rect 11846 2883 11880 3139
rect 12024 2883 12058 3139
rect 12202 2883 12236 3139
rect 12380 2883 12414 3139
rect 12558 2883 12592 3139
rect 12736 2883 12770 3139
rect 428 2183 462 2439
rect 606 2183 640 2439
rect 784 2183 818 2439
rect 962 2183 996 2439
rect 1140 2183 1174 2439
rect 1318 2183 1352 2439
rect 1496 2183 1530 2439
rect 1674 2183 1708 2439
rect 1852 2183 1886 2439
rect 2030 2183 2064 2439
rect 2208 2183 2242 2439
rect 2386 2183 2420 2439
rect 2564 2183 2598 2439
rect 2742 2183 2776 2439
rect 2920 2183 2954 2439
rect 3098 2183 3132 2439
rect 3276 2183 3310 2439
rect 3454 2183 3488 2439
rect 3632 2183 3666 2439
rect 3828 2183 3862 2439
rect 4006 2183 4040 2439
rect 4184 2183 4218 2439
rect 4362 2183 4396 2439
rect 4540 2183 4574 2439
rect 4718 2183 4752 2439
rect 4896 2183 4930 2439
rect 5074 2183 5108 2439
rect 5252 2183 5286 2439
rect 5430 2183 5464 2439
rect 5608 2183 5642 2439
rect 5786 2183 5820 2439
rect 5964 2183 5998 2439
rect 6142 2183 6176 2439
rect 6320 2183 6354 2439
rect 6498 2183 6532 2439
rect 6676 2183 6710 2439
rect 6854 2183 6888 2439
rect 7032 2183 7066 2439
rect 7557 2383 7591 2639
rect 7735 2383 7769 2639
rect 7913 2383 7947 2639
rect 8091 2383 8125 2639
rect 8269 2383 8303 2639
rect 8447 2383 8481 2639
rect 8625 2383 8659 2639
rect 8803 2383 8837 2639
rect 8981 2383 9015 2639
rect 9159 2383 9193 2639
rect 9337 2383 9371 2639
rect 9515 2383 9549 2639
rect 9693 2383 9727 2639
rect 9871 2383 9905 2639
rect 10049 2383 10083 2639
rect 10244 2383 10278 2639
rect 10422 2383 10456 2639
rect 10600 2383 10634 2639
rect 10778 2383 10812 2639
rect 10956 2383 10990 2639
rect 11134 2383 11168 2639
rect 11312 2383 11346 2639
rect 11490 2383 11524 2639
rect 11668 2383 11702 2639
rect 11846 2383 11880 2639
rect 12024 2383 12058 2639
rect 12202 2383 12236 2639
rect 12380 2383 12414 2639
rect 12558 2383 12592 2639
rect 12736 2383 12770 2639
rect 428 1683 462 1939
rect 606 1683 640 1939
rect 784 1683 818 1939
rect 962 1683 996 1939
rect 1140 1683 1174 1939
rect 1318 1683 1352 1939
rect 1496 1683 1530 1939
rect 1674 1683 1708 1939
rect 1852 1683 1886 1939
rect 2030 1683 2064 1939
rect 2208 1683 2242 1939
rect 2386 1683 2420 1939
rect 2564 1683 2598 1939
rect 2742 1683 2776 1939
rect 2920 1683 2954 1939
rect 3098 1683 3132 1939
rect 3276 1683 3310 1939
rect 3454 1683 3488 1939
rect 3632 1683 3666 1939
rect 3828 1683 3862 1939
rect 4006 1683 4040 1939
rect 4184 1683 4218 1939
rect 4362 1683 4396 1939
rect 4540 1683 4574 1939
rect 4718 1683 4752 1939
rect 4896 1683 4930 1939
rect 5074 1683 5108 1939
rect 5252 1683 5286 1939
rect 5430 1683 5464 1939
rect 5608 1683 5642 1939
rect 5786 1683 5820 1939
rect 5964 1683 5998 1939
rect 6142 1683 6176 1939
rect 6320 1683 6354 1939
rect 6498 1683 6532 1939
rect 6676 1683 6710 1939
rect 6854 1683 6888 1939
rect 7032 1683 7066 1939
rect 7557 1683 7591 1939
rect 7735 1683 7769 1939
rect 7913 1683 7947 1939
rect 8091 1683 8125 1939
rect 8269 1683 8303 1939
rect 8447 1683 8481 1939
rect 8625 1683 8659 1939
rect 8803 1683 8837 1939
rect 8981 1683 9015 1939
rect 9159 1683 9193 1939
rect 9337 1683 9371 1939
rect 9515 1683 9549 1939
rect 9693 1683 9727 1939
rect 9871 1683 9905 1939
rect 10049 1683 10083 1939
rect 10244 1683 10278 1939
rect 10422 1683 10456 1939
rect 10600 1683 10634 1939
rect 10778 1683 10812 1939
rect 10956 1683 10990 1939
rect 11134 1683 11168 1939
rect 11312 1683 11346 1939
rect 11490 1683 11524 1939
rect 11668 1683 11702 1939
rect 11846 1683 11880 1939
rect 12024 1683 12058 1939
rect 12202 1683 12236 1939
rect 12380 1683 12414 1939
rect 12558 1683 12592 1939
rect 12736 1683 12770 1939
rect 428 1183 462 1439
rect 606 1183 640 1439
rect 784 1183 818 1439
rect 962 1183 996 1439
rect 1140 1183 1174 1439
rect 1318 1183 1352 1439
rect 1496 1183 1530 1439
rect 1674 1183 1708 1439
rect 1852 1183 1886 1439
rect 2030 1183 2064 1439
rect 2208 1183 2242 1439
rect 2386 1183 2420 1439
rect 2564 1183 2598 1439
rect 2742 1183 2776 1439
rect 2920 1183 2954 1439
rect 3098 1183 3132 1439
rect 3276 1183 3310 1439
rect 3454 1183 3488 1439
rect 3632 1183 3666 1439
rect 3828 1183 3862 1439
rect 4006 1183 4040 1439
rect 4184 1183 4218 1439
rect 4362 1183 4396 1439
rect 4540 1183 4574 1439
rect 4718 1183 4752 1439
rect 4896 1183 4930 1439
rect 5074 1183 5108 1439
rect 5252 1183 5286 1439
rect 5430 1183 5464 1439
rect 5608 1183 5642 1439
rect 5786 1183 5820 1439
rect 5964 1183 5998 1439
rect 6142 1183 6176 1439
rect 6320 1183 6354 1439
rect 6498 1183 6532 1439
rect 6676 1183 6710 1439
rect 6854 1183 6888 1439
rect 7032 1183 7066 1439
rect 7557 1183 7591 1439
rect 7735 1183 7769 1439
rect 7913 1183 7947 1439
rect 8091 1183 8125 1439
rect 8269 1183 8303 1439
rect 8447 1183 8481 1439
rect 8625 1183 8659 1439
rect 8803 1183 8837 1439
rect 8981 1183 9015 1439
rect 9159 1183 9193 1439
rect 9337 1183 9371 1439
rect 9515 1183 9549 1439
rect 9693 1183 9727 1439
rect 9871 1183 9905 1439
rect 10049 1183 10083 1439
rect 10244 1183 10278 1439
rect 10422 1183 10456 1439
rect 10600 1183 10634 1439
rect 10778 1183 10812 1439
rect 10956 1183 10990 1439
rect 11134 1183 11168 1439
rect 11312 1183 11346 1439
rect 11490 1183 11524 1439
rect 11668 1183 11702 1439
rect 11846 1183 11880 1439
rect 12024 1183 12058 1439
rect 12202 1183 12236 1439
rect 12380 1183 12414 1439
rect 12558 1183 12592 1439
rect 12736 1183 12770 1439
rect 428 683 462 939
rect 606 683 640 939
rect 784 683 818 939
rect 962 683 996 939
rect 1140 683 1174 939
rect 1318 683 1352 939
rect 1496 683 1530 939
rect 1674 683 1708 939
rect 1852 683 1886 939
rect 2030 683 2064 939
rect 2208 683 2242 939
rect 2386 683 2420 939
rect 2564 683 2598 939
rect 2742 683 2776 939
rect 2920 683 2954 939
rect 3098 683 3132 939
rect 3276 683 3310 939
rect 3454 683 3488 939
rect 3632 683 3666 939
rect 3828 683 3862 939
rect 4006 683 4040 939
rect 4184 683 4218 939
rect 4362 683 4396 939
rect 4540 683 4574 939
rect 4718 683 4752 939
rect 4896 683 4930 939
rect 5074 683 5108 939
rect 5252 683 5286 939
rect 5430 683 5464 939
rect 5608 683 5642 939
rect 5786 683 5820 939
rect 5964 683 5998 939
rect 6142 683 6176 939
rect 6320 683 6354 939
rect 6498 683 6532 939
rect 6676 683 6710 939
rect 6854 683 6888 939
rect 7032 683 7066 939
rect 7557 683 7591 939
rect 7735 683 7769 939
rect 7913 683 7947 939
rect 8091 683 8125 939
rect 8269 683 8303 939
rect 8447 683 8481 939
rect 8625 683 8659 939
rect 8803 683 8837 939
rect 8981 683 9015 939
rect 9159 683 9193 939
rect 9337 683 9371 939
rect 9515 683 9549 939
rect 9693 683 9727 939
rect 9871 683 9905 939
rect 10049 683 10083 939
rect 10244 683 10278 939
rect 10422 683 10456 939
rect 10600 683 10634 939
rect 10778 683 10812 939
rect 10956 683 10990 939
rect 11134 683 11168 939
rect 11312 683 11346 939
rect 11490 683 11524 939
rect 11668 683 11702 939
rect 11846 683 11880 939
rect 12024 683 12058 939
rect 12202 683 12236 939
rect 12380 683 12414 939
rect 12558 683 12592 939
rect 12736 683 12770 939
rect 13550 4791 13584 5047
rect 13728 4791 13762 5047
rect 13906 4791 13940 5047
rect 14084 4791 14118 5047
rect 14262 4791 14296 5047
rect 14440 4791 14474 5047
rect 14618 4791 14652 5047
rect 14796 4791 14830 5047
rect 14974 4791 15008 5047
rect 15152 4791 15186 5047
rect 15330 4791 15364 5047
rect 15508 4791 15542 5047
rect 15686 4791 15720 5047
rect 15864 4791 15898 5047
rect 16042 4791 16076 5047
rect 16220 4791 16254 5047
rect 16398 4791 16432 5047
rect 16576 4791 16610 5047
rect 16754 4791 16788 5047
rect 16932 4791 16966 5047
rect 17110 4791 17144 5047
rect 17288 4791 17322 5047
rect 17466 4791 17500 5047
rect 17644 4791 17678 5047
rect 17822 4791 17856 5047
rect 18000 4791 18034 5047
rect 18178 4791 18212 5047
rect 18356 4791 18390 5047
rect 13550 4291 13584 4547
rect 13728 4291 13762 4547
rect 13906 4291 13940 4547
rect 14084 4291 14118 4547
rect 14262 4291 14296 4547
rect 14440 4291 14474 4547
rect 14618 4291 14652 4547
rect 14796 4291 14830 4547
rect 14974 4291 15008 4547
rect 15152 4291 15186 4547
rect 15330 4291 15364 4547
rect 15508 4291 15542 4547
rect 15686 4291 15720 4547
rect 15864 4291 15898 4547
rect 16042 4291 16076 4547
rect 16220 4291 16254 4547
rect 16398 4291 16432 4547
rect 16576 4291 16610 4547
rect 16754 4291 16788 4547
rect 16932 4291 16966 4547
rect 17110 4291 17144 4547
rect 17288 4291 17322 4547
rect 17466 4291 17500 4547
rect 17644 4291 17678 4547
rect 17822 4291 17856 4547
rect 18000 4291 18034 4547
rect 18178 4291 18212 4547
rect 18356 4291 18390 4547
rect 17108 3287 17142 3543
rect 17286 3287 17320 3543
rect 17464 3287 17498 3543
rect 17642 3287 17676 3543
rect 17820 3287 17854 3543
rect 13676 2282 13710 2538
rect 13854 2282 13888 2538
rect 13968 2282 14002 2538
rect 14146 2282 14180 2538
rect 14260 2282 14294 2538
rect 14438 2282 14472 2538
rect 14552 2282 14586 2538
rect 14730 2282 14764 2538
rect 14844 2282 14878 2538
rect 15022 2282 15056 2538
rect 15136 2282 15170 2538
rect 15314 2282 15348 2538
rect 15428 2282 15462 2538
rect 15606 2282 15640 2538
rect 16394 2348 16428 2604
rect 16572 2348 16606 2604
rect 16750 2348 16784 2604
rect 16928 2348 16962 2604
rect 17106 2348 17140 2604
rect 17284 2348 17318 2604
rect 17462 2348 17496 2604
rect 17640 2348 17674 2604
rect 17818 2348 17852 2604
rect 17996 2348 18030 2604
rect 18174 2348 18208 2604
rect 18352 2348 18386 2604
rect 13676 1784 13710 2040
rect 13854 1784 13888 2040
rect 13968 1784 14002 2040
rect 14146 1784 14180 2040
rect 14260 1784 14294 2040
rect 14438 1784 14472 2040
rect 14552 1784 14586 2040
rect 14730 1784 14764 2040
rect 14844 1784 14878 2040
rect 15022 1784 15056 2040
rect 15136 1784 15170 2040
rect 15314 1784 15348 2040
rect 15428 1784 15462 2040
rect 15606 1784 15640 2040
rect 16394 1848 16428 2104
rect 16572 1848 16606 2104
rect 16750 1848 16784 2104
rect 16928 1848 16962 2104
rect 17106 1848 17140 2104
rect 17284 1848 17318 2104
rect 17462 1848 17496 2104
rect 17640 1848 17674 2104
rect 17818 1848 17852 2104
rect 17996 1848 18030 2104
rect 18174 1848 18208 2104
rect 18352 1848 18386 2104
rect 13676 1286 13710 1542
rect 13854 1286 13888 1542
rect 13968 1286 14002 1542
rect 14146 1286 14180 1542
rect 14260 1286 14294 1542
rect 14438 1286 14472 1542
rect 14552 1286 14586 1542
rect 14730 1286 14764 1542
rect 14844 1286 14878 1542
rect 15022 1286 15056 1542
rect 15136 1286 15170 1542
rect 15314 1286 15348 1542
rect 15428 1286 15462 1542
rect 15606 1286 15640 1542
rect 16394 1288 16428 1544
rect 16572 1288 16606 1544
rect 16750 1288 16784 1544
rect 16928 1288 16962 1544
rect 17106 1288 17140 1544
rect 17284 1288 17318 1544
rect 17462 1288 17496 1544
rect 17640 1288 17674 1544
rect 17818 1288 17852 1544
rect 17996 1288 18030 1544
rect 18174 1288 18208 1544
rect 18352 1288 18386 1544
rect 13676 788 13710 1044
rect 13854 788 13888 1044
rect 13968 788 14002 1044
rect 14146 788 14180 1044
rect 14260 788 14294 1044
rect 14438 788 14472 1044
rect 14552 788 14586 1044
rect 14730 788 14764 1044
rect 14844 788 14878 1044
rect 15022 788 15056 1044
rect 15136 788 15170 1044
rect 15314 788 15348 1044
rect 15428 788 15462 1044
rect 15606 788 15640 1044
rect 16394 788 16428 1044
rect 16572 788 16606 1044
rect 16750 788 16784 1044
rect 16928 788 16962 1044
rect 17106 788 17140 1044
rect 17284 788 17318 1044
rect 17462 788 17496 1044
rect 17640 788 17674 1044
rect 17818 788 17852 1044
rect 17996 788 18030 1044
rect 18174 788 18208 1044
rect 18352 788 18386 1044
rect 19009 4782 19043 5038
rect 19187 4782 19221 5038
rect 19365 4782 19399 5038
rect 19543 4782 19577 5038
rect 19721 4782 19755 5038
rect 19899 4782 19933 5038
rect 20077 4782 20111 5038
rect 20255 4782 20289 5038
rect 20433 4782 20467 5038
rect 20611 4782 20645 5038
rect 20789 4782 20823 5038
rect 20967 4782 21001 5038
rect 21145 4782 21179 5038
rect 21323 4782 21357 5038
rect 21501 4782 21535 5038
rect 21679 4782 21713 5038
rect 21857 4782 21891 5038
rect 19009 4284 19043 4540
rect 19187 4284 19221 4540
rect 19365 4284 19399 4540
rect 19543 4284 19577 4540
rect 19721 4284 19755 4540
rect 19899 4284 19933 4540
rect 20077 4284 20111 4540
rect 20255 4284 20289 4540
rect 20433 4284 20467 4540
rect 20611 4284 20645 4540
rect 20789 4284 20823 4540
rect 20967 4284 21001 4540
rect 21145 4284 21179 4540
rect 21323 4284 21357 4540
rect 21501 4284 21535 4540
rect 21679 4284 21713 4540
rect 21857 4284 21891 4540
rect 19009 3786 19043 4042
rect 19187 3786 19221 4042
rect 19365 3786 19399 4042
rect 19543 3786 19577 4042
rect 19721 3786 19755 4042
rect 19899 3786 19933 4042
rect 20077 3786 20111 4042
rect 20255 3786 20289 4042
rect 20433 3786 20467 4042
rect 20611 3786 20645 4042
rect 20789 3786 20823 4042
rect 20967 3786 21001 4042
rect 21145 3786 21179 4042
rect 21323 3786 21357 4042
rect 21501 3786 21535 4042
rect 21679 3786 21713 4042
rect 21857 3786 21891 4042
rect 19009 3288 19043 3544
rect 19187 3288 19221 3544
rect 19365 3288 19399 3544
rect 19543 3288 19577 3544
rect 19721 3288 19755 3544
rect 19899 3288 19933 3544
rect 20077 3288 20111 3544
rect 20255 3288 20289 3544
rect 20433 3288 20467 3544
rect 20611 3288 20645 3544
rect 20789 3288 20823 3544
rect 20967 3288 21001 3544
rect 21145 3288 21179 3544
rect 21323 3288 21357 3544
rect 21501 3288 21535 3544
rect 21679 3288 21713 3544
rect 21857 3288 21891 3544
rect 19367 2274 19401 2530
rect 19545 2274 19579 2530
rect 19723 2274 19757 2530
rect 19901 2274 19935 2530
rect 20079 2274 20113 2530
rect 20257 2274 20291 2530
rect 20435 2274 20469 2530
rect 20613 2274 20647 2530
rect 20791 2274 20825 2530
rect 20969 2274 21003 2530
rect 21147 2274 21181 2530
rect 21325 2274 21359 2530
rect 19367 1776 19401 2032
rect 19545 1776 19579 2032
rect 19723 1776 19757 2032
rect 19901 1776 19935 2032
rect 20079 1776 20113 2032
rect 20257 1776 20291 2032
rect 20435 1776 20469 2032
rect 20613 1776 20647 2032
rect 20791 1776 20825 2032
rect 20969 1776 21003 2032
rect 21147 1776 21181 2032
rect 21325 1776 21359 2032
rect 19367 1278 19401 1534
rect 19545 1278 19579 1534
rect 19723 1278 19757 1534
rect 19901 1278 19935 1534
rect 20079 1278 20113 1534
rect 20257 1278 20291 1534
rect 20435 1278 20469 1534
rect 20613 1278 20647 1534
rect 20791 1278 20825 1534
rect 20969 1278 21003 1534
rect 21147 1278 21181 1534
rect 21325 1278 21359 1534
rect 19367 780 19401 1036
rect 19545 780 19579 1036
rect 19723 780 19757 1036
rect 19901 780 19935 1036
rect 20079 780 20113 1036
rect 20257 780 20291 1036
rect 20435 780 20469 1036
rect 20613 780 20647 1036
rect 20791 780 20825 1036
rect 20969 780 21003 1036
rect 21147 780 21181 1036
rect 21325 780 21359 1036
<< pdiffc >>
rect 7303 18493 7337 18741
rect 7399 18493 7433 18741
rect 7495 18493 7529 18741
rect 7591 18493 7625 18741
rect 7687 18493 7721 18741
rect 7783 18493 7817 18741
rect 7879 18493 7913 18741
rect 7975 18493 8009 18741
rect 8071 18493 8105 18741
rect 8167 18493 8201 18741
rect 8263 18493 8297 18741
rect 20233 18493 20267 18741
rect 20329 18493 20363 18741
rect 20425 18493 20459 18741
rect 20521 18493 20555 18741
rect 20617 18493 20651 18741
rect 20713 18493 20747 18741
rect 20809 18493 20843 18741
rect 20905 18493 20939 18741
rect 21001 18493 21035 18741
rect 21097 18493 21131 18741
rect 21193 18493 21227 18741
rect 7303 16693 7337 16941
rect 7399 16693 7433 16941
rect 7495 16693 7529 16941
rect 7591 16693 7625 16941
rect 7687 16693 7721 16941
rect 7783 16693 7817 16941
rect 7879 16693 7913 16941
rect 7975 16693 8009 16941
rect 8071 16693 8105 16941
rect 8167 16693 8201 16941
rect 8263 16693 8297 16941
rect 20233 16693 20267 16941
rect 20329 16693 20363 16941
rect 20425 16693 20459 16941
rect 20521 16693 20555 16941
rect 20617 16693 20651 16941
rect 20713 16693 20747 16941
rect 20809 16693 20843 16941
rect 20905 16693 20939 16941
rect 21001 16693 21035 16941
rect 21097 16693 21131 16941
rect 21193 16693 21227 16941
rect 7303 14893 7337 15141
rect 7399 14893 7433 15141
rect 7495 14893 7529 15141
rect 7591 14893 7625 15141
rect 7687 14893 7721 15141
rect 7783 14893 7817 15141
rect 7879 14893 7913 15141
rect 7975 14893 8009 15141
rect 8071 14893 8105 15141
rect 8167 14893 8201 15141
rect 8263 14893 8297 15141
rect 20233 14893 20267 15141
rect 20329 14893 20363 15141
rect 20425 14893 20459 15141
rect 20521 14893 20555 15141
rect 20617 14893 20651 15141
rect 20713 14893 20747 15141
rect 20809 14893 20843 15141
rect 20905 14893 20939 15141
rect 21001 14893 21035 15141
rect 21097 14893 21131 15141
rect 21193 14893 21227 15141
rect 7303 13093 7337 13341
rect 7399 13093 7433 13341
rect 7495 13093 7529 13341
rect 7591 13093 7625 13341
rect 7687 13093 7721 13341
rect 7783 13093 7817 13341
rect 7879 13093 7913 13341
rect 7975 13093 8009 13341
rect 8071 13093 8105 13341
rect 8167 13093 8201 13341
rect 8263 13093 8297 13341
rect 20233 13093 20267 13341
rect 20329 13093 20363 13341
rect 20425 13093 20459 13341
rect 20521 13093 20555 13341
rect 20617 13093 20651 13341
rect 20713 13093 20747 13341
rect 20809 13093 20843 13341
rect 20905 13093 20939 13341
rect 21001 13093 21035 13341
rect 21097 13093 21131 13341
rect 21193 13093 21227 13341
rect 7303 11293 7337 11541
rect 7399 11293 7433 11541
rect 7495 11293 7529 11541
rect 7591 11293 7625 11541
rect 7687 11293 7721 11541
rect 7783 11293 7817 11541
rect 7879 11293 7913 11541
rect 7975 11293 8009 11541
rect 8071 11293 8105 11541
rect 8167 11293 8201 11541
rect 8263 11293 8297 11541
rect 20233 11293 20267 11541
rect 20329 11293 20363 11541
rect 20425 11293 20459 11541
rect 20521 11293 20555 11541
rect 20617 11293 20651 11541
rect 20713 11293 20747 11541
rect 20809 11293 20843 11541
rect 20905 11293 20939 11541
rect 21001 11293 21035 11541
rect 21097 11293 21131 11541
rect 21193 11293 21227 11541
rect 7303 9493 7337 9741
rect 7399 9493 7433 9741
rect 7495 9493 7529 9741
rect 7591 9493 7625 9741
rect 7687 9493 7721 9741
rect 7783 9493 7817 9741
rect 7879 9493 7913 9741
rect 7975 9493 8009 9741
rect 8071 9493 8105 9741
rect 8167 9493 8201 9741
rect 8263 9493 8297 9741
rect 20233 9493 20267 9741
rect 20329 9493 20363 9741
rect 20425 9493 20459 9741
rect 20521 9493 20555 9741
rect 20617 9493 20651 9741
rect 20713 9493 20747 9741
rect 20809 9493 20843 9741
rect 20905 9493 20939 9741
rect 21001 9493 21035 9741
rect 21097 9493 21131 9741
rect 21193 9493 21227 9741
rect 7556 6341 7590 6597
rect 7734 6341 7768 6597
rect 7912 6341 7946 6597
rect 8090 6341 8124 6597
rect 8268 6341 8302 6597
rect 8446 6341 8480 6597
rect 8624 6341 8658 6597
rect 8802 6341 8836 6597
rect 8980 6341 9014 6597
rect 9158 6341 9192 6597
rect 9336 6341 9370 6597
rect 9514 6341 9548 6597
rect 9692 6341 9726 6597
rect 9870 6341 9904 6597
rect 10048 6341 10082 6597
rect 10242 6341 10276 6597
rect 10420 6341 10454 6597
rect 10598 6341 10632 6597
rect 10776 6341 10810 6597
rect 10954 6341 10988 6597
rect 11132 6341 11166 6597
rect 11310 6341 11344 6597
rect 11488 6341 11522 6597
rect 11666 6341 11700 6597
rect 11844 6341 11878 6597
rect 12022 6341 12056 6597
rect 12200 6341 12234 6597
rect 12378 6341 12412 6597
rect 12556 6341 12590 6597
rect 12734 6341 12768 6597
rect 7556 5763 7590 6019
rect 7734 5763 7768 6019
rect 7912 5763 7946 6019
rect 8090 5763 8124 6019
rect 8268 5763 8302 6019
rect 8446 5763 8480 6019
rect 8624 5763 8658 6019
rect 8802 5763 8836 6019
rect 8980 5763 9014 6019
rect 9158 5763 9192 6019
rect 9336 5763 9370 6019
rect 9514 5763 9548 6019
rect 9692 5763 9726 6019
rect 9870 5763 9904 6019
rect 10048 5763 10082 6019
rect 10242 5764 10276 6020
rect 10420 5764 10454 6020
rect 10598 5764 10632 6020
rect 10776 5764 10810 6020
rect 10954 5764 10988 6020
rect 11132 5764 11166 6020
rect 11310 5764 11344 6020
rect 11488 5764 11522 6020
rect 11666 5764 11700 6020
rect 11844 5764 11878 6020
rect 12022 5764 12056 6020
rect 12200 5764 12234 6020
rect 12378 5764 12412 6020
rect 12556 5764 12590 6020
rect 12734 5764 12768 6020
rect 14696 6410 14730 6666
rect 14874 6410 14908 6666
rect 15052 6410 15086 6666
rect 15230 6410 15264 6666
rect 15408 6410 15442 6666
rect 15586 6410 15620 6666
rect 15764 6410 15798 6666
rect 15942 6410 15976 6666
rect 16120 6410 16154 6666
rect 16896 6410 16930 6666
rect 17074 6410 17108 6666
rect 17252 6410 17286 6666
rect 17430 6410 17464 6666
rect 17608 6410 17642 6666
rect 17786 6410 17820 6666
rect 17964 6410 17998 6666
rect 18142 6410 18176 6666
rect 18320 6410 18354 6666
rect 19096 6410 19130 6666
rect 19274 6410 19308 6666
rect 19452 6410 19486 6666
rect 19630 6410 19664 6666
rect 19808 6410 19842 6666
rect 19986 6410 20020 6666
rect 20164 6410 20198 6666
rect 20342 6410 20376 6666
rect 20520 6410 20554 6666
rect 14697 5643 14731 5899
rect 14875 5643 14909 5899
rect 15053 5643 15087 5899
rect 15231 5643 15265 5899
rect 15409 5643 15443 5899
rect 15587 5643 15621 5899
rect 15765 5643 15799 5899
rect 15943 5643 15977 5899
rect 16121 5643 16155 5899
rect 16897 5643 16931 5899
rect 17075 5643 17109 5899
rect 17253 5643 17287 5899
rect 17431 5643 17465 5899
rect 17609 5643 17643 5899
rect 17787 5643 17821 5899
rect 17965 5643 17999 5899
rect 18143 5643 18177 5899
rect 18321 5643 18355 5899
rect 19097 5643 19131 5899
rect 19275 5643 19309 5899
rect 19453 5643 19487 5899
rect 19631 5643 19665 5899
rect 19809 5643 19843 5899
rect 19987 5643 20021 5899
rect 20165 5643 20199 5899
rect 20343 5643 20377 5899
rect 20521 5643 20555 5899
rect 7912 4883 7946 5139
rect 8090 4883 8124 5139
rect 8268 4883 8302 5139
rect 8446 4883 8480 5139
rect 8624 4883 8658 5139
rect 8802 4883 8836 5139
rect 8980 4883 9014 5139
rect 9158 4883 9192 5139
rect 9336 4883 9370 5139
rect 9514 4883 9548 5139
rect 9692 4883 9726 5139
rect 9870 4883 9904 5139
rect 10048 4883 10082 5139
rect 10242 4883 10276 5139
rect 10420 4883 10454 5139
rect 10598 4883 10632 5139
rect 10776 4883 10810 5139
rect 10954 4883 10988 5139
rect 11132 4883 11166 5139
rect 11310 4883 11344 5139
rect 11488 4883 11522 5139
rect 11666 4883 11700 5139
rect 11844 4883 11878 5139
rect 12022 4883 12056 5139
rect 12200 4883 12234 5139
rect 12378 4883 12412 5139
rect 7912 4313 7946 4569
rect 8090 4313 8124 4569
rect 8268 4313 8302 4569
rect 8446 4313 8480 4569
rect 8624 4313 8658 4569
rect 8802 4313 8836 4569
rect 8980 4313 9014 4569
rect 9158 4313 9192 4569
rect 9336 4313 9370 4569
rect 9514 4313 9548 4569
rect 9692 4313 9726 4569
rect 9870 4313 9904 4569
rect 10048 4313 10082 4569
rect 10242 4313 10276 4569
rect 10420 4313 10454 4569
rect 10598 4313 10632 4569
rect 10776 4313 10810 4569
rect 10954 4313 10988 4569
rect 11132 4313 11166 4569
rect 11310 4313 11344 4569
rect 11488 4313 11522 4569
rect 11666 4313 11700 4569
rect 11844 4313 11878 4569
rect 12022 4313 12056 4569
rect 12200 4313 12234 4569
rect 12378 4313 12412 4569
<< psubdiff >>
rect 7189 18253 7285 18287
rect 8315 18253 8411 18287
rect 7189 18191 7223 18253
rect 8377 18191 8411 18253
rect 7189 17931 7223 17993
rect 8377 17931 8411 17993
rect 7189 17897 7285 17931
rect 8315 17897 8411 17931
rect 20119 18253 20215 18287
rect 21245 18253 21341 18287
rect 20119 18191 20153 18253
rect 21307 18191 21341 18253
rect 20119 17931 20153 17993
rect 21307 17931 21341 17993
rect 20119 17897 20215 17931
rect 21245 17897 21341 17931
rect 7189 16453 7285 16487
rect 8315 16453 8411 16487
rect 7189 16391 7223 16453
rect 8377 16391 8411 16453
rect 7189 16131 7223 16193
rect 8377 16131 8411 16193
rect 7189 16097 7285 16131
rect 8315 16097 8411 16131
rect 20119 16453 20215 16487
rect 21245 16453 21341 16487
rect 20119 16391 20153 16453
rect 21307 16391 21341 16453
rect 20119 16131 20153 16193
rect 21307 16131 21341 16193
rect 20119 16097 20215 16131
rect 21245 16097 21341 16131
rect 7189 14653 7285 14687
rect 8315 14653 8411 14687
rect 7189 14591 7223 14653
rect 8377 14591 8411 14653
rect 7189 14331 7223 14393
rect 8377 14331 8411 14393
rect 7189 14297 7285 14331
rect 8315 14297 8411 14331
rect 20119 14653 20215 14687
rect 21245 14653 21341 14687
rect 20119 14591 20153 14653
rect 21307 14591 21341 14653
rect 20119 14331 20153 14393
rect 21307 14331 21341 14393
rect 20119 14297 20215 14331
rect 21245 14297 21341 14331
rect 7189 12853 7285 12887
rect 8315 12853 8411 12887
rect 7189 12791 7223 12853
rect 8377 12791 8411 12853
rect 7189 12531 7223 12593
rect 8377 12531 8411 12593
rect 7189 12497 7285 12531
rect 8315 12497 8411 12531
rect 20119 12853 20215 12887
rect 21245 12853 21341 12887
rect 20119 12791 20153 12853
rect 21307 12791 21341 12853
rect 20119 12531 20153 12593
rect 21307 12531 21341 12593
rect 20119 12497 20215 12531
rect 21245 12497 21341 12531
rect 7189 11053 7285 11087
rect 8315 11053 8411 11087
rect 7189 10991 7223 11053
rect 8377 10991 8411 11053
rect 7189 10731 7223 10793
rect 8377 10731 8411 10793
rect 7189 10697 7285 10731
rect 8315 10697 8411 10731
rect 20119 11053 20215 11087
rect 21245 11053 21341 11087
rect 20119 10991 20153 11053
rect 21307 10991 21341 11053
rect 20119 10731 20153 10793
rect 21307 10731 21341 10793
rect 20119 10697 20215 10731
rect 21245 10697 21341 10731
rect 7189 9253 7285 9287
rect 8315 9253 8411 9287
rect 7189 9191 7223 9253
rect 8377 9191 8411 9253
rect 7189 8931 7223 8993
rect 8377 8931 8411 8993
rect 7189 8897 7285 8931
rect 8315 8897 8411 8931
rect 20119 9253 20215 9287
rect 21245 9253 21341 9287
rect 20119 9191 20153 9253
rect 21307 9191 21341 9253
rect 20119 8931 20153 8993
rect 21307 8931 21341 8993
rect 20119 8897 20215 8931
rect 21245 8897 21341 8931
rect 161 4600 272 4649
rect 6855 4600 6973 4649
rect 161 4548 210 4600
rect 6924 4564 6973 4600
rect 13318 5260 13367 5261
rect 13318 5211 13584 5260
rect 18360 5211 18506 5260
rect 13318 5128 13367 5211
rect 6924 3934 6973 3960
rect 6924 3885 7001 3934
rect 13229 3885 13318 3934
rect 161 71 210 149
rect 18457 5145 18506 5211
rect 13318 71 13367 113
rect 18895 5190 18991 5224
rect 21909 5190 22005 5224
rect 18895 5128 18929 5190
rect 21971 5128 22005 5190
rect 18895 3136 18929 3198
rect 21971 3136 22005 3198
rect 18895 3102 18991 3136
rect 21909 3102 22005 3136
rect 19253 2682 19349 2716
rect 21377 2682 21473 2716
rect 19253 2620 19287 2682
rect 21439 2620 21473 2682
rect 19253 628 19287 690
rect 21439 628 21473 690
rect 19253 594 19349 628
rect 21377 594 21473 628
rect 161 22 304 71
rect 13205 70 13460 71
rect 18457 70 18506 149
rect 13205 22 13476 70
rect 13318 21 13476 22
rect 18366 21 18506 70
<< nsubdiff >>
rect 7189 18903 7285 18937
rect 8315 18903 8411 18937
rect 7189 18841 7223 18903
rect 8377 18841 8411 18903
rect 7189 18393 7223 18455
rect 8377 18393 8411 18455
rect 7189 18359 7285 18393
rect 8315 18359 8411 18393
rect 20119 18903 20215 18937
rect 21245 18903 21341 18937
rect 20119 18841 20153 18903
rect 21307 18841 21341 18903
rect 20119 18393 20153 18455
rect 21307 18393 21341 18455
rect 20119 18359 20215 18393
rect 21245 18359 21341 18393
rect 7189 17103 7285 17137
rect 8315 17103 8411 17137
rect 7189 17041 7223 17103
rect 8377 17041 8411 17103
rect 7189 16593 7223 16655
rect 8377 16593 8411 16655
rect 7189 16559 7285 16593
rect 8315 16559 8411 16593
rect 20119 17103 20215 17137
rect 21245 17103 21341 17137
rect 20119 17041 20153 17103
rect 21307 17041 21341 17103
rect 20119 16593 20153 16655
rect 21307 16593 21341 16655
rect 20119 16559 20215 16593
rect 21245 16559 21341 16593
rect 7189 15303 7285 15337
rect 8315 15303 8411 15337
rect 7189 15241 7223 15303
rect 8377 15241 8411 15303
rect 7189 14793 7223 14855
rect 8377 14793 8411 14855
rect 7189 14759 7285 14793
rect 8315 14759 8411 14793
rect 20119 15303 20215 15337
rect 21245 15303 21341 15337
rect 20119 15241 20153 15303
rect 21307 15241 21341 15303
rect 20119 14793 20153 14855
rect 21307 14793 21341 14855
rect 20119 14759 20215 14793
rect 21245 14759 21341 14793
rect 7189 13503 7285 13537
rect 8315 13503 8411 13537
rect 7189 13441 7223 13503
rect 8377 13441 8411 13503
rect 7189 12993 7223 13055
rect 8377 12993 8411 13055
rect 7189 12959 7285 12993
rect 8315 12959 8411 12993
rect 20119 13503 20215 13537
rect 21245 13503 21341 13537
rect 20119 13441 20153 13503
rect 21307 13441 21341 13503
rect 20119 12993 20153 13055
rect 21307 12993 21341 13055
rect 20119 12959 20215 12993
rect 21245 12959 21341 12993
rect 7189 11703 7285 11737
rect 8315 11703 8411 11737
rect 7189 11641 7223 11703
rect 8377 11641 8411 11703
rect 7189 11193 7223 11255
rect 8377 11193 8411 11255
rect 7189 11159 7285 11193
rect 8315 11159 8411 11193
rect 20119 11703 20215 11737
rect 21245 11703 21341 11737
rect 20119 11641 20153 11703
rect 21307 11641 21341 11703
rect 20119 11193 20153 11255
rect 21307 11193 21341 11255
rect 20119 11159 20215 11193
rect 21245 11159 21341 11193
rect 7189 9903 7285 9937
rect 8315 9903 8411 9937
rect 7189 9841 7223 9903
rect 8377 9841 8411 9903
rect 7189 9393 7223 9455
rect 8377 9393 8411 9455
rect 7189 9359 7285 9393
rect 8315 9359 8411 9393
rect 20119 9903 20215 9937
rect 21245 9903 21341 9937
rect 20119 9841 20153 9903
rect 21307 9841 21341 9903
rect 20119 9393 20153 9455
rect 21307 9393 21341 9455
rect 20119 9359 20215 9393
rect 21245 9359 21341 9393
rect 7310 6957 7445 6991
rect 14299 6957 14467 6991
rect 20872 6957 20977 6991
rect 7310 6852 7344 6957
rect 14358 6892 14392 6957
rect 20943 6919 20977 6957
rect 14358 5413 14392 5525
rect 20943 5413 20977 5483
rect 12999 5379 13108 5413
rect 14264 5379 14464 5413
rect 20857 5379 20977 5413
rect 12999 5315 13033 5379
rect 7310 4124 7344 4198
rect 12999 4124 13033 4221
rect 7310 4090 7453 4124
rect 12924 4090 13033 4124
<< psubdiffcont >>
rect 7285 18253 8315 18287
rect 7189 17993 7223 18191
rect 8377 17993 8411 18191
rect 7285 17897 8315 17931
rect 20215 18253 21245 18287
rect 20119 17993 20153 18191
rect 21307 17993 21341 18191
rect 20215 17897 21245 17931
rect 7285 16453 8315 16487
rect 7189 16193 7223 16391
rect 8377 16193 8411 16391
rect 7285 16097 8315 16131
rect 20215 16453 21245 16487
rect 20119 16193 20153 16391
rect 21307 16193 21341 16391
rect 20215 16097 21245 16131
rect 7285 14653 8315 14687
rect 7189 14393 7223 14591
rect 8377 14393 8411 14591
rect 7285 14297 8315 14331
rect 20215 14653 21245 14687
rect 20119 14393 20153 14591
rect 21307 14393 21341 14591
rect 20215 14297 21245 14331
rect 7285 12853 8315 12887
rect 7189 12593 7223 12791
rect 8377 12593 8411 12791
rect 7285 12497 8315 12531
rect 20215 12853 21245 12887
rect 20119 12593 20153 12791
rect 21307 12593 21341 12791
rect 20215 12497 21245 12531
rect 7285 11053 8315 11087
rect 7189 10793 7223 10991
rect 8377 10793 8411 10991
rect 7285 10697 8315 10731
rect 20215 11053 21245 11087
rect 20119 10793 20153 10991
rect 21307 10793 21341 10991
rect 20215 10697 21245 10731
rect 7285 9253 8315 9287
rect 7189 8993 7223 9191
rect 8377 8993 8411 9191
rect 7285 8897 8315 8931
rect 20215 9253 21245 9287
rect 20119 8993 20153 9191
rect 21307 8993 21341 9191
rect 20215 8897 21245 8931
rect 272 4600 6855 4649
rect 161 149 210 4548
rect 6924 3960 6973 4564
rect 13584 5211 18360 5260
rect 7001 3885 13229 3934
rect 13318 113 13367 5128
rect 18457 149 18506 5145
rect 18991 5190 21909 5224
rect 18895 3198 18929 5128
rect 21971 3198 22005 5128
rect 18991 3102 21909 3136
rect 19349 2682 21377 2716
rect 19253 690 19287 2620
rect 21439 690 21473 2620
rect 19349 594 21377 628
rect 304 22 13205 71
rect 13476 21 18366 70
<< nsubdiffcont >>
rect 7285 18903 8315 18937
rect 7189 18455 7223 18841
rect 8377 18455 8411 18841
rect 7285 18359 8315 18393
rect 20215 18903 21245 18937
rect 20119 18455 20153 18841
rect 21307 18455 21341 18841
rect 20215 18359 21245 18393
rect 7285 17103 8315 17137
rect 7189 16655 7223 17041
rect 8377 16655 8411 17041
rect 7285 16559 8315 16593
rect 20215 17103 21245 17137
rect 20119 16655 20153 17041
rect 21307 16655 21341 17041
rect 20215 16559 21245 16593
rect 7285 15303 8315 15337
rect 7189 14855 7223 15241
rect 8377 14855 8411 15241
rect 7285 14759 8315 14793
rect 20215 15303 21245 15337
rect 20119 14855 20153 15241
rect 21307 14855 21341 15241
rect 20215 14759 21245 14793
rect 7285 13503 8315 13537
rect 7189 13055 7223 13441
rect 8377 13055 8411 13441
rect 7285 12959 8315 12993
rect 20215 13503 21245 13537
rect 20119 13055 20153 13441
rect 21307 13055 21341 13441
rect 20215 12959 21245 12993
rect 7285 11703 8315 11737
rect 7189 11255 7223 11641
rect 8377 11255 8411 11641
rect 7285 11159 8315 11193
rect 20215 11703 21245 11737
rect 20119 11255 20153 11641
rect 21307 11255 21341 11641
rect 20215 11159 21245 11193
rect 7285 9903 8315 9937
rect 7189 9455 7223 9841
rect 8377 9455 8411 9841
rect 7285 9359 8315 9393
rect 20215 9903 21245 9937
rect 20119 9455 20153 9841
rect 21307 9455 21341 9841
rect 20215 9359 21245 9393
rect 7445 6957 14299 6991
rect 14467 6957 20872 6991
rect 7310 4198 7344 6852
rect 14358 5525 14392 6892
rect 20943 5483 20977 6919
rect 13108 5379 14264 5413
rect 14464 5379 20857 5413
rect 12999 4221 13033 5315
rect 7453 4090 12924 4124
<< poly >>
rect 7287 18835 8313 18851
rect 7287 18801 7303 18835
rect 7337 18801 7495 18835
rect 7529 18801 7687 18835
rect 7721 18801 7879 18835
rect 7913 18801 8071 18835
rect 8105 18801 8263 18835
rect 8297 18801 8313 18835
rect 7287 18785 8313 18801
rect 7353 18753 7383 18785
rect 7449 18753 7479 18785
rect 7545 18753 7575 18785
rect 7641 18753 7671 18785
rect 7737 18753 7767 18785
rect 7833 18753 7863 18785
rect 7929 18753 7959 18785
rect 8025 18753 8055 18785
rect 8121 18753 8151 18785
rect 8217 18753 8247 18785
rect 7353 18455 7383 18481
rect 7449 18455 7479 18481
rect 7545 18455 7575 18481
rect 7641 18455 7671 18481
rect 7737 18455 7767 18481
rect 7833 18455 7863 18481
rect 7929 18455 7959 18481
rect 8025 18455 8055 18481
rect 8121 18455 8151 18481
rect 8217 18455 8247 18481
rect 20217 18835 21243 18851
rect 20217 18801 20233 18835
rect 20267 18801 20425 18835
rect 20459 18801 20617 18835
rect 20651 18801 20809 18835
rect 20843 18801 21001 18835
rect 21035 18801 21193 18835
rect 21227 18801 21243 18835
rect 20217 18785 21243 18801
rect 20283 18753 20313 18785
rect 20379 18753 20409 18785
rect 20475 18753 20505 18785
rect 20571 18753 20601 18785
rect 20667 18753 20697 18785
rect 20763 18753 20793 18785
rect 20859 18753 20889 18785
rect 20955 18753 20985 18785
rect 21051 18753 21081 18785
rect 21147 18753 21177 18785
rect 20283 18455 20313 18481
rect 20379 18455 20409 18481
rect 20475 18455 20505 18481
rect 20571 18455 20601 18481
rect 20667 18455 20697 18481
rect 20763 18455 20793 18481
rect 20859 18455 20889 18481
rect 20955 18455 20985 18481
rect 21051 18455 21081 18481
rect 21147 18455 21177 18481
rect 7353 18175 7383 18201
rect 7449 18175 7479 18201
rect 7545 18175 7575 18201
rect 7641 18175 7671 18201
rect 7737 18175 7767 18201
rect 7833 18175 7863 18201
rect 7929 18175 7959 18201
rect 8025 18175 8055 18201
rect 8121 18175 8151 18201
rect 8217 18175 8247 18201
rect 7353 18040 7383 18071
rect 7449 18040 7479 18071
rect 7545 18040 7575 18071
rect 7641 18040 7671 18071
rect 7737 18040 7767 18071
rect 7833 18040 7863 18071
rect 7929 18040 7959 18071
rect 8025 18040 8055 18071
rect 8121 18040 8151 18071
rect 8217 18040 8247 18071
rect 7287 18024 8313 18040
rect 7287 17990 7303 18024
rect 7337 17990 7495 18024
rect 7529 17990 7687 18024
rect 7721 17990 7879 18024
rect 7913 17990 8071 18024
rect 8105 17990 8263 18024
rect 8297 17990 8313 18024
rect 7287 17974 8313 17990
rect 20283 18175 20313 18201
rect 20379 18175 20409 18201
rect 20475 18175 20505 18201
rect 20571 18175 20601 18201
rect 20667 18175 20697 18201
rect 20763 18175 20793 18201
rect 20859 18175 20889 18201
rect 20955 18175 20985 18201
rect 21051 18175 21081 18201
rect 21147 18175 21177 18201
rect 20283 18040 20313 18071
rect 20379 18040 20409 18071
rect 20475 18040 20505 18071
rect 20571 18040 20601 18071
rect 20667 18040 20697 18071
rect 20763 18040 20793 18071
rect 20859 18040 20889 18071
rect 20955 18040 20985 18071
rect 21051 18040 21081 18071
rect 21147 18040 21177 18071
rect 20217 18024 21243 18040
rect 20217 17990 20233 18024
rect 20267 17990 20425 18024
rect 20459 17990 20617 18024
rect 20651 17990 20809 18024
rect 20843 17990 21001 18024
rect 21035 17990 21193 18024
rect 21227 17990 21243 18024
rect 20217 17974 21243 17990
rect 7287 17035 8313 17051
rect 7287 17001 7303 17035
rect 7337 17001 7495 17035
rect 7529 17001 7687 17035
rect 7721 17001 7879 17035
rect 7913 17001 8071 17035
rect 8105 17001 8263 17035
rect 8297 17001 8313 17035
rect 7287 16985 8313 17001
rect 7353 16953 7383 16985
rect 7449 16953 7479 16985
rect 7545 16953 7575 16985
rect 7641 16953 7671 16985
rect 7737 16953 7767 16985
rect 7833 16953 7863 16985
rect 7929 16953 7959 16985
rect 8025 16953 8055 16985
rect 8121 16953 8151 16985
rect 8217 16953 8247 16985
rect 7353 16655 7383 16681
rect 7449 16655 7479 16681
rect 7545 16655 7575 16681
rect 7641 16655 7671 16681
rect 7737 16655 7767 16681
rect 7833 16655 7863 16681
rect 7929 16655 7959 16681
rect 8025 16655 8055 16681
rect 8121 16655 8151 16681
rect 8217 16655 8247 16681
rect 20217 17035 21243 17051
rect 20217 17001 20233 17035
rect 20267 17001 20425 17035
rect 20459 17001 20617 17035
rect 20651 17001 20809 17035
rect 20843 17001 21001 17035
rect 21035 17001 21193 17035
rect 21227 17001 21243 17035
rect 20217 16985 21243 17001
rect 20283 16953 20313 16985
rect 20379 16953 20409 16985
rect 20475 16953 20505 16985
rect 20571 16953 20601 16985
rect 20667 16953 20697 16985
rect 20763 16953 20793 16985
rect 20859 16953 20889 16985
rect 20955 16953 20985 16985
rect 21051 16953 21081 16985
rect 21147 16953 21177 16985
rect 20283 16655 20313 16681
rect 20379 16655 20409 16681
rect 20475 16655 20505 16681
rect 20571 16655 20601 16681
rect 20667 16655 20697 16681
rect 20763 16655 20793 16681
rect 20859 16655 20889 16681
rect 20955 16655 20985 16681
rect 21051 16655 21081 16681
rect 21147 16655 21177 16681
rect 7353 16375 7383 16401
rect 7449 16375 7479 16401
rect 7545 16375 7575 16401
rect 7641 16375 7671 16401
rect 7737 16375 7767 16401
rect 7833 16375 7863 16401
rect 7929 16375 7959 16401
rect 8025 16375 8055 16401
rect 8121 16375 8151 16401
rect 8217 16375 8247 16401
rect 7353 16240 7383 16271
rect 7449 16240 7479 16271
rect 7545 16240 7575 16271
rect 7641 16240 7671 16271
rect 7737 16240 7767 16271
rect 7833 16240 7863 16271
rect 7929 16240 7959 16271
rect 8025 16240 8055 16271
rect 8121 16240 8151 16271
rect 8217 16240 8247 16271
rect 7287 16224 8313 16240
rect 7287 16190 7303 16224
rect 7337 16190 7495 16224
rect 7529 16190 7687 16224
rect 7721 16190 7879 16224
rect 7913 16190 8071 16224
rect 8105 16190 8263 16224
rect 8297 16190 8313 16224
rect 7287 16174 8313 16190
rect 20283 16375 20313 16401
rect 20379 16375 20409 16401
rect 20475 16375 20505 16401
rect 20571 16375 20601 16401
rect 20667 16375 20697 16401
rect 20763 16375 20793 16401
rect 20859 16375 20889 16401
rect 20955 16375 20985 16401
rect 21051 16375 21081 16401
rect 21147 16375 21177 16401
rect 20283 16240 20313 16271
rect 20379 16240 20409 16271
rect 20475 16240 20505 16271
rect 20571 16240 20601 16271
rect 20667 16240 20697 16271
rect 20763 16240 20793 16271
rect 20859 16240 20889 16271
rect 20955 16240 20985 16271
rect 21051 16240 21081 16271
rect 21147 16240 21177 16271
rect 20217 16224 21243 16240
rect 20217 16190 20233 16224
rect 20267 16190 20425 16224
rect 20459 16190 20617 16224
rect 20651 16190 20809 16224
rect 20843 16190 21001 16224
rect 21035 16190 21193 16224
rect 21227 16190 21243 16224
rect 20217 16174 21243 16190
rect 7287 15235 8313 15251
rect 7287 15201 7303 15235
rect 7337 15201 7495 15235
rect 7529 15201 7687 15235
rect 7721 15201 7879 15235
rect 7913 15201 8071 15235
rect 8105 15201 8263 15235
rect 8297 15201 8313 15235
rect 7287 15185 8313 15201
rect 7353 15153 7383 15185
rect 7449 15153 7479 15185
rect 7545 15153 7575 15185
rect 7641 15153 7671 15185
rect 7737 15153 7767 15185
rect 7833 15153 7863 15185
rect 7929 15153 7959 15185
rect 8025 15153 8055 15185
rect 8121 15153 8151 15185
rect 8217 15153 8247 15185
rect 7353 14855 7383 14881
rect 7449 14855 7479 14881
rect 7545 14855 7575 14881
rect 7641 14855 7671 14881
rect 7737 14855 7767 14881
rect 7833 14855 7863 14881
rect 7929 14855 7959 14881
rect 8025 14855 8055 14881
rect 8121 14855 8151 14881
rect 8217 14855 8247 14881
rect 20217 15235 21243 15251
rect 20217 15201 20233 15235
rect 20267 15201 20425 15235
rect 20459 15201 20617 15235
rect 20651 15201 20809 15235
rect 20843 15201 21001 15235
rect 21035 15201 21193 15235
rect 21227 15201 21243 15235
rect 20217 15185 21243 15201
rect 20283 15153 20313 15185
rect 20379 15153 20409 15185
rect 20475 15153 20505 15185
rect 20571 15153 20601 15185
rect 20667 15153 20697 15185
rect 20763 15153 20793 15185
rect 20859 15153 20889 15185
rect 20955 15153 20985 15185
rect 21051 15153 21081 15185
rect 21147 15153 21177 15185
rect 20283 14855 20313 14881
rect 20379 14855 20409 14881
rect 20475 14855 20505 14881
rect 20571 14855 20601 14881
rect 20667 14855 20697 14881
rect 20763 14855 20793 14881
rect 20859 14855 20889 14881
rect 20955 14855 20985 14881
rect 21051 14855 21081 14881
rect 21147 14855 21177 14881
rect 7353 14575 7383 14601
rect 7449 14575 7479 14601
rect 7545 14575 7575 14601
rect 7641 14575 7671 14601
rect 7737 14575 7767 14601
rect 7833 14575 7863 14601
rect 7929 14575 7959 14601
rect 8025 14575 8055 14601
rect 8121 14575 8151 14601
rect 8217 14575 8247 14601
rect 7353 14440 7383 14471
rect 7449 14440 7479 14471
rect 7545 14440 7575 14471
rect 7641 14440 7671 14471
rect 7737 14440 7767 14471
rect 7833 14440 7863 14471
rect 7929 14440 7959 14471
rect 8025 14440 8055 14471
rect 8121 14440 8151 14471
rect 8217 14440 8247 14471
rect 7287 14424 8313 14440
rect 7287 14390 7303 14424
rect 7337 14390 7495 14424
rect 7529 14390 7687 14424
rect 7721 14390 7879 14424
rect 7913 14390 8071 14424
rect 8105 14390 8263 14424
rect 8297 14390 8313 14424
rect 7287 14374 8313 14390
rect 20283 14575 20313 14601
rect 20379 14575 20409 14601
rect 20475 14575 20505 14601
rect 20571 14575 20601 14601
rect 20667 14575 20697 14601
rect 20763 14575 20793 14601
rect 20859 14575 20889 14601
rect 20955 14575 20985 14601
rect 21051 14575 21081 14601
rect 21147 14575 21177 14601
rect 20283 14440 20313 14471
rect 20379 14440 20409 14471
rect 20475 14440 20505 14471
rect 20571 14440 20601 14471
rect 20667 14440 20697 14471
rect 20763 14440 20793 14471
rect 20859 14440 20889 14471
rect 20955 14440 20985 14471
rect 21051 14440 21081 14471
rect 21147 14440 21177 14471
rect 20217 14424 21243 14440
rect 20217 14390 20233 14424
rect 20267 14390 20425 14424
rect 20459 14390 20617 14424
rect 20651 14390 20809 14424
rect 20843 14390 21001 14424
rect 21035 14390 21193 14424
rect 21227 14390 21243 14424
rect 20217 14374 21243 14390
rect 7287 13435 8313 13451
rect 7287 13401 7303 13435
rect 7337 13401 7495 13435
rect 7529 13401 7687 13435
rect 7721 13401 7879 13435
rect 7913 13401 8071 13435
rect 8105 13401 8263 13435
rect 8297 13401 8313 13435
rect 7287 13385 8313 13401
rect 7353 13353 7383 13385
rect 7449 13353 7479 13385
rect 7545 13353 7575 13385
rect 7641 13353 7671 13385
rect 7737 13353 7767 13385
rect 7833 13353 7863 13385
rect 7929 13353 7959 13385
rect 8025 13353 8055 13385
rect 8121 13353 8151 13385
rect 8217 13353 8247 13385
rect 7353 13055 7383 13081
rect 7449 13055 7479 13081
rect 7545 13055 7575 13081
rect 7641 13055 7671 13081
rect 7737 13055 7767 13081
rect 7833 13055 7863 13081
rect 7929 13055 7959 13081
rect 8025 13055 8055 13081
rect 8121 13055 8151 13081
rect 8217 13055 8247 13081
rect 20217 13435 21243 13451
rect 20217 13401 20233 13435
rect 20267 13401 20425 13435
rect 20459 13401 20617 13435
rect 20651 13401 20809 13435
rect 20843 13401 21001 13435
rect 21035 13401 21193 13435
rect 21227 13401 21243 13435
rect 20217 13385 21243 13401
rect 20283 13353 20313 13385
rect 20379 13353 20409 13385
rect 20475 13353 20505 13385
rect 20571 13353 20601 13385
rect 20667 13353 20697 13385
rect 20763 13353 20793 13385
rect 20859 13353 20889 13385
rect 20955 13353 20985 13385
rect 21051 13353 21081 13385
rect 21147 13353 21177 13385
rect 20283 13055 20313 13081
rect 20379 13055 20409 13081
rect 20475 13055 20505 13081
rect 20571 13055 20601 13081
rect 20667 13055 20697 13081
rect 20763 13055 20793 13081
rect 20859 13055 20889 13081
rect 20955 13055 20985 13081
rect 21051 13055 21081 13081
rect 21147 13055 21177 13081
rect 7353 12775 7383 12801
rect 7449 12775 7479 12801
rect 7545 12775 7575 12801
rect 7641 12775 7671 12801
rect 7737 12775 7767 12801
rect 7833 12775 7863 12801
rect 7929 12775 7959 12801
rect 8025 12775 8055 12801
rect 8121 12775 8151 12801
rect 8217 12775 8247 12801
rect 7353 12640 7383 12671
rect 7449 12640 7479 12671
rect 7545 12640 7575 12671
rect 7641 12640 7671 12671
rect 7737 12640 7767 12671
rect 7833 12640 7863 12671
rect 7929 12640 7959 12671
rect 8025 12640 8055 12671
rect 8121 12640 8151 12671
rect 8217 12640 8247 12671
rect 7287 12624 8313 12640
rect 7287 12590 7303 12624
rect 7337 12590 7495 12624
rect 7529 12590 7687 12624
rect 7721 12590 7879 12624
rect 7913 12590 8071 12624
rect 8105 12590 8263 12624
rect 8297 12590 8313 12624
rect 7287 12574 8313 12590
rect 20283 12775 20313 12801
rect 20379 12775 20409 12801
rect 20475 12775 20505 12801
rect 20571 12775 20601 12801
rect 20667 12775 20697 12801
rect 20763 12775 20793 12801
rect 20859 12775 20889 12801
rect 20955 12775 20985 12801
rect 21051 12775 21081 12801
rect 21147 12775 21177 12801
rect 20283 12640 20313 12671
rect 20379 12640 20409 12671
rect 20475 12640 20505 12671
rect 20571 12640 20601 12671
rect 20667 12640 20697 12671
rect 20763 12640 20793 12671
rect 20859 12640 20889 12671
rect 20955 12640 20985 12671
rect 21051 12640 21081 12671
rect 21147 12640 21177 12671
rect 20217 12624 21243 12640
rect 20217 12590 20233 12624
rect 20267 12590 20425 12624
rect 20459 12590 20617 12624
rect 20651 12590 20809 12624
rect 20843 12590 21001 12624
rect 21035 12590 21193 12624
rect 21227 12590 21243 12624
rect 20217 12574 21243 12590
rect 7287 11635 8313 11651
rect 7287 11601 7303 11635
rect 7337 11601 7495 11635
rect 7529 11601 7687 11635
rect 7721 11601 7879 11635
rect 7913 11601 8071 11635
rect 8105 11601 8263 11635
rect 8297 11601 8313 11635
rect 7287 11585 8313 11601
rect 7353 11553 7383 11585
rect 7449 11553 7479 11585
rect 7545 11553 7575 11585
rect 7641 11553 7671 11585
rect 7737 11553 7767 11585
rect 7833 11553 7863 11585
rect 7929 11553 7959 11585
rect 8025 11553 8055 11585
rect 8121 11553 8151 11585
rect 8217 11553 8247 11585
rect 7353 11255 7383 11281
rect 7449 11255 7479 11281
rect 7545 11255 7575 11281
rect 7641 11255 7671 11281
rect 7737 11255 7767 11281
rect 7833 11255 7863 11281
rect 7929 11255 7959 11281
rect 8025 11255 8055 11281
rect 8121 11255 8151 11281
rect 8217 11255 8247 11281
rect 20217 11635 21243 11651
rect 20217 11601 20233 11635
rect 20267 11601 20425 11635
rect 20459 11601 20617 11635
rect 20651 11601 20809 11635
rect 20843 11601 21001 11635
rect 21035 11601 21193 11635
rect 21227 11601 21243 11635
rect 20217 11585 21243 11601
rect 20283 11553 20313 11585
rect 20379 11553 20409 11585
rect 20475 11553 20505 11585
rect 20571 11553 20601 11585
rect 20667 11553 20697 11585
rect 20763 11553 20793 11585
rect 20859 11553 20889 11585
rect 20955 11553 20985 11585
rect 21051 11553 21081 11585
rect 21147 11553 21177 11585
rect 20283 11255 20313 11281
rect 20379 11255 20409 11281
rect 20475 11255 20505 11281
rect 20571 11255 20601 11281
rect 20667 11255 20697 11281
rect 20763 11255 20793 11281
rect 20859 11255 20889 11281
rect 20955 11255 20985 11281
rect 21051 11255 21081 11281
rect 21147 11255 21177 11281
rect 7353 10975 7383 11001
rect 7449 10975 7479 11001
rect 7545 10975 7575 11001
rect 7641 10975 7671 11001
rect 7737 10975 7767 11001
rect 7833 10975 7863 11001
rect 7929 10975 7959 11001
rect 8025 10975 8055 11001
rect 8121 10975 8151 11001
rect 8217 10975 8247 11001
rect 7353 10840 7383 10871
rect 7449 10840 7479 10871
rect 7545 10840 7575 10871
rect 7641 10840 7671 10871
rect 7737 10840 7767 10871
rect 7833 10840 7863 10871
rect 7929 10840 7959 10871
rect 8025 10840 8055 10871
rect 8121 10840 8151 10871
rect 8217 10840 8247 10871
rect 7287 10824 8313 10840
rect 7287 10790 7303 10824
rect 7337 10790 7495 10824
rect 7529 10790 7687 10824
rect 7721 10790 7879 10824
rect 7913 10790 8071 10824
rect 8105 10790 8263 10824
rect 8297 10790 8313 10824
rect 7287 10774 8313 10790
rect 20283 10975 20313 11001
rect 20379 10975 20409 11001
rect 20475 10975 20505 11001
rect 20571 10975 20601 11001
rect 20667 10975 20697 11001
rect 20763 10975 20793 11001
rect 20859 10975 20889 11001
rect 20955 10975 20985 11001
rect 21051 10975 21081 11001
rect 21147 10975 21177 11001
rect 20283 10840 20313 10871
rect 20379 10840 20409 10871
rect 20475 10840 20505 10871
rect 20571 10840 20601 10871
rect 20667 10840 20697 10871
rect 20763 10840 20793 10871
rect 20859 10840 20889 10871
rect 20955 10840 20985 10871
rect 21051 10840 21081 10871
rect 21147 10840 21177 10871
rect 20217 10824 21243 10840
rect 20217 10790 20233 10824
rect 20267 10790 20425 10824
rect 20459 10790 20617 10824
rect 20651 10790 20809 10824
rect 20843 10790 21001 10824
rect 21035 10790 21193 10824
rect 21227 10790 21243 10824
rect 20217 10774 21243 10790
rect 7287 9835 8313 9851
rect 7287 9801 7303 9835
rect 7337 9801 7495 9835
rect 7529 9801 7687 9835
rect 7721 9801 7879 9835
rect 7913 9801 8071 9835
rect 8105 9801 8263 9835
rect 8297 9801 8313 9835
rect 7287 9785 8313 9801
rect 7353 9753 7383 9785
rect 7449 9753 7479 9785
rect 7545 9753 7575 9785
rect 7641 9753 7671 9785
rect 7737 9753 7767 9785
rect 7833 9753 7863 9785
rect 7929 9753 7959 9785
rect 8025 9753 8055 9785
rect 8121 9753 8151 9785
rect 8217 9753 8247 9785
rect 7353 9455 7383 9481
rect 7449 9455 7479 9481
rect 7545 9455 7575 9481
rect 7641 9455 7671 9481
rect 7737 9455 7767 9481
rect 7833 9455 7863 9481
rect 7929 9455 7959 9481
rect 8025 9455 8055 9481
rect 8121 9455 8151 9481
rect 8217 9455 8247 9481
rect 20217 9835 21243 9851
rect 20217 9801 20233 9835
rect 20267 9801 20425 9835
rect 20459 9801 20617 9835
rect 20651 9801 20809 9835
rect 20843 9801 21001 9835
rect 21035 9801 21193 9835
rect 21227 9801 21243 9835
rect 20217 9785 21243 9801
rect 20283 9753 20313 9785
rect 20379 9753 20409 9785
rect 20475 9753 20505 9785
rect 20571 9753 20601 9785
rect 20667 9753 20697 9785
rect 20763 9753 20793 9785
rect 20859 9753 20889 9785
rect 20955 9753 20985 9785
rect 21051 9753 21081 9785
rect 21147 9753 21177 9785
rect 20283 9455 20313 9481
rect 20379 9455 20409 9481
rect 20475 9455 20505 9481
rect 20571 9455 20601 9481
rect 20667 9455 20697 9481
rect 20763 9455 20793 9481
rect 20859 9455 20889 9481
rect 20955 9455 20985 9481
rect 21051 9455 21081 9481
rect 21147 9455 21177 9481
rect 7353 9175 7383 9201
rect 7449 9175 7479 9201
rect 7545 9175 7575 9201
rect 7641 9175 7671 9201
rect 7737 9175 7767 9201
rect 7833 9175 7863 9201
rect 7929 9175 7959 9201
rect 8025 9175 8055 9201
rect 8121 9175 8151 9201
rect 8217 9175 8247 9201
rect 7353 9040 7383 9071
rect 7449 9040 7479 9071
rect 7545 9040 7575 9071
rect 7641 9040 7671 9071
rect 7737 9040 7767 9071
rect 7833 9040 7863 9071
rect 7929 9040 7959 9071
rect 8025 9040 8055 9071
rect 8121 9040 8151 9071
rect 8217 9040 8247 9071
rect 7287 9024 8313 9040
rect 7287 8990 7303 9024
rect 7337 8990 7495 9024
rect 7529 8990 7687 9024
rect 7721 8990 7879 9024
rect 7913 8990 8071 9024
rect 8105 8990 8263 9024
rect 8297 8990 8313 9024
rect 7287 8974 8313 8990
rect 20283 9175 20313 9201
rect 20379 9175 20409 9201
rect 20475 9175 20505 9201
rect 20571 9175 20601 9201
rect 20667 9175 20697 9201
rect 20763 9175 20793 9201
rect 20859 9175 20889 9201
rect 20955 9175 20985 9201
rect 21051 9175 21081 9201
rect 21147 9175 21177 9201
rect 20283 9040 20313 9071
rect 20379 9040 20409 9071
rect 20475 9040 20505 9071
rect 20571 9040 20601 9071
rect 20667 9040 20697 9071
rect 20763 9040 20793 9071
rect 20859 9040 20889 9071
rect 20955 9040 20985 9071
rect 21051 9040 21081 9071
rect 21147 9040 21177 9071
rect 20217 9024 21243 9040
rect 20217 8990 20233 9024
rect 20267 8990 20425 9024
rect 20459 8990 20617 9024
rect 20651 8990 20809 9024
rect 20843 8990 21001 9024
rect 21035 8990 21193 9024
rect 21227 8990 21243 9024
rect 20217 8974 21243 8990
rect 2084 4303 2150 4319
rect 2084 4269 2100 4303
rect 2134 4269 2150 4303
rect 2084 4253 2150 4269
rect 2508 4303 2574 4319
rect 2508 4269 2524 4303
rect 2558 4269 2574 4303
rect 2096 4231 2136 4253
rect 2308 4231 2348 4257
rect 2508 4253 2574 4269
rect 2930 4303 2996 4319
rect 2930 4269 2946 4303
rect 2980 4269 2996 4303
rect 2520 4231 2560 4253
rect 2732 4231 2772 4257
rect 2930 4253 2996 4269
rect 3354 4303 3420 4319
rect 3354 4269 3370 4303
rect 3404 4269 3420 4303
rect 2944 4231 2984 4253
rect 3156 4231 3196 4257
rect 3354 4253 3420 4269
rect 3864 4303 3930 4319
rect 3864 4269 3880 4303
rect 3914 4269 3930 4303
rect 3368 4231 3408 4253
rect 3580 4231 3620 4257
rect 3864 4253 3930 4269
rect 4288 4303 4354 4319
rect 4288 4269 4304 4303
rect 4338 4269 4354 4303
rect 3876 4231 3916 4253
rect 4088 4231 4128 4257
rect 4288 4253 4354 4269
rect 4710 4303 4776 4319
rect 4710 4269 4726 4303
rect 4760 4269 4776 4303
rect 4300 4231 4340 4253
rect 4512 4231 4552 4257
rect 4710 4253 4776 4269
rect 5134 4303 5200 4319
rect 5134 4269 5150 4303
rect 5184 4269 5200 4303
rect 4724 4231 4764 4253
rect 4936 4231 4976 4257
rect 5134 4253 5200 4269
rect 5148 4231 5188 4253
rect 5360 4231 5400 4257
rect 2096 3965 2136 3991
rect 2308 3969 2348 3991
rect 2296 3953 2362 3969
rect 2520 3965 2560 3991
rect 2732 3969 2772 3991
rect 2296 3919 2312 3953
rect 2346 3919 2362 3953
rect 2296 3903 2362 3919
rect 2720 3953 2786 3969
rect 2944 3965 2984 3991
rect 3156 3969 3196 3991
rect 2720 3919 2736 3953
rect 2770 3919 2786 3953
rect 2720 3903 2786 3919
rect 3142 3953 3208 3969
rect 3368 3965 3408 3991
rect 3580 3969 3620 3991
rect 3142 3919 3158 3953
rect 3192 3919 3208 3953
rect 3142 3903 3208 3919
rect 3566 3953 3632 3969
rect 3876 3965 3916 3991
rect 4088 3969 4128 3991
rect 3566 3919 3582 3953
rect 3616 3919 3632 3953
rect 3566 3903 3632 3919
rect 4076 3953 4142 3969
rect 4300 3965 4340 3991
rect 4512 3969 4552 3991
rect 4076 3919 4092 3953
rect 4126 3919 4142 3953
rect 4076 3903 4142 3919
rect 4500 3953 4566 3969
rect 4724 3965 4764 3991
rect 4936 3969 4976 3991
rect 4500 3919 4516 3953
rect 4550 3919 4566 3953
rect 4500 3903 4566 3919
rect 4922 3953 4988 3969
rect 5148 3965 5188 3991
rect 5360 3969 5400 3991
rect 4922 3919 4938 3953
rect 4972 3919 4988 3953
rect 4922 3903 4988 3919
rect 5346 3953 5412 3969
rect 5346 3919 5362 3953
rect 5396 3919 5412 3953
rect 5346 3903 5412 3919
rect 7620 6690 7704 6706
rect 7620 6674 7636 6690
rect 7602 6656 7636 6674
rect 7688 6674 7704 6690
rect 7798 6690 7882 6706
rect 7798 6674 7814 6690
rect 7688 6656 7722 6674
rect 7602 6609 7722 6656
rect 7780 6656 7814 6674
rect 7866 6674 7882 6690
rect 7976 6690 8060 6706
rect 7976 6674 7992 6690
rect 7866 6656 7900 6674
rect 7780 6609 7900 6656
rect 7958 6656 7992 6674
rect 8044 6674 8060 6690
rect 8154 6690 8238 6706
rect 8154 6674 8170 6690
rect 8044 6656 8078 6674
rect 7958 6609 8078 6656
rect 8136 6656 8170 6674
rect 8222 6674 8238 6690
rect 8332 6690 8416 6706
rect 8332 6674 8348 6690
rect 8222 6656 8256 6674
rect 8136 6609 8256 6656
rect 8314 6656 8348 6674
rect 8400 6674 8416 6690
rect 8510 6690 8594 6706
rect 8510 6674 8526 6690
rect 8400 6656 8434 6674
rect 8314 6609 8434 6656
rect 8492 6656 8526 6674
rect 8578 6674 8594 6690
rect 8688 6690 8772 6706
rect 8688 6674 8704 6690
rect 8578 6656 8612 6674
rect 8492 6609 8612 6656
rect 8670 6656 8704 6674
rect 8756 6674 8772 6690
rect 8866 6690 8950 6706
rect 8866 6674 8882 6690
rect 8756 6656 8790 6674
rect 8670 6609 8790 6656
rect 8848 6656 8882 6674
rect 8934 6674 8950 6690
rect 9044 6690 9128 6706
rect 9044 6674 9060 6690
rect 8934 6656 8968 6674
rect 8848 6609 8968 6656
rect 9026 6656 9060 6674
rect 9112 6674 9128 6690
rect 9222 6690 9306 6706
rect 9222 6674 9238 6690
rect 9112 6656 9146 6674
rect 9026 6609 9146 6656
rect 9204 6656 9238 6674
rect 9290 6674 9306 6690
rect 9400 6690 9484 6706
rect 9400 6674 9416 6690
rect 9290 6656 9324 6674
rect 9204 6609 9324 6656
rect 9382 6656 9416 6674
rect 9468 6674 9484 6690
rect 9578 6690 9662 6706
rect 9578 6674 9594 6690
rect 9468 6656 9502 6674
rect 9382 6609 9502 6656
rect 9560 6656 9594 6674
rect 9646 6674 9662 6690
rect 9756 6690 9840 6706
rect 9756 6674 9772 6690
rect 9646 6656 9680 6674
rect 9560 6609 9680 6656
rect 9738 6656 9772 6674
rect 9824 6674 9840 6690
rect 9934 6690 10018 6706
rect 9934 6674 9950 6690
rect 9824 6656 9858 6674
rect 9738 6609 9858 6656
rect 9916 6656 9950 6674
rect 10002 6674 10018 6690
rect 10306 6690 10390 6706
rect 10306 6674 10322 6690
rect 10002 6656 10036 6674
rect 9916 6609 10036 6656
rect 10288 6656 10322 6674
rect 10374 6674 10390 6690
rect 10484 6690 10568 6706
rect 10484 6674 10500 6690
rect 10374 6656 10408 6674
rect 10288 6609 10408 6656
rect 10466 6656 10500 6674
rect 10552 6674 10568 6690
rect 10662 6690 10746 6706
rect 10662 6674 10678 6690
rect 10552 6656 10586 6674
rect 10466 6609 10586 6656
rect 10644 6656 10678 6674
rect 10730 6674 10746 6690
rect 10840 6690 10924 6706
rect 10840 6674 10856 6690
rect 10730 6656 10764 6674
rect 10644 6609 10764 6656
rect 10822 6656 10856 6674
rect 10908 6674 10924 6690
rect 11018 6690 11102 6706
rect 11018 6674 11034 6690
rect 10908 6656 10942 6674
rect 10822 6609 10942 6656
rect 11000 6656 11034 6674
rect 11086 6674 11102 6690
rect 11196 6690 11280 6706
rect 11196 6674 11212 6690
rect 11086 6656 11120 6674
rect 11000 6609 11120 6656
rect 11178 6656 11212 6674
rect 11264 6674 11280 6690
rect 11374 6690 11458 6706
rect 11374 6674 11390 6690
rect 11264 6656 11298 6674
rect 11178 6609 11298 6656
rect 11356 6656 11390 6674
rect 11442 6674 11458 6690
rect 11552 6690 11636 6706
rect 11552 6674 11568 6690
rect 11442 6656 11476 6674
rect 11356 6609 11476 6656
rect 11534 6656 11568 6674
rect 11620 6674 11636 6690
rect 11730 6690 11814 6706
rect 11730 6674 11746 6690
rect 11620 6656 11654 6674
rect 11534 6609 11654 6656
rect 11712 6656 11746 6674
rect 11798 6674 11814 6690
rect 11908 6690 11992 6706
rect 11908 6674 11924 6690
rect 11798 6656 11832 6674
rect 11712 6609 11832 6656
rect 11890 6656 11924 6674
rect 11976 6674 11992 6690
rect 12086 6690 12170 6706
rect 12086 6674 12102 6690
rect 11976 6656 12010 6674
rect 11890 6609 12010 6656
rect 12068 6656 12102 6674
rect 12154 6674 12170 6690
rect 12264 6690 12348 6706
rect 12264 6674 12280 6690
rect 12154 6656 12188 6674
rect 12068 6609 12188 6656
rect 12246 6656 12280 6674
rect 12332 6674 12348 6690
rect 12442 6690 12526 6706
rect 12442 6674 12458 6690
rect 12332 6656 12366 6674
rect 12246 6609 12366 6656
rect 12424 6656 12458 6674
rect 12510 6674 12526 6690
rect 12620 6690 12704 6706
rect 12620 6674 12636 6690
rect 12510 6656 12544 6674
rect 12424 6609 12544 6656
rect 12602 6656 12636 6674
rect 12688 6674 12704 6690
rect 12688 6656 12722 6674
rect 12602 6609 12722 6656
rect 7602 6282 7722 6329
rect 7602 6264 7636 6282
rect 7620 6248 7636 6264
rect 7688 6264 7722 6282
rect 7780 6282 7900 6329
rect 7780 6264 7814 6282
rect 7688 6248 7704 6264
rect 7620 6232 7704 6248
rect 7798 6248 7814 6264
rect 7866 6264 7900 6282
rect 7958 6282 8078 6329
rect 7958 6264 7992 6282
rect 7866 6248 7882 6264
rect 7798 6232 7882 6248
rect 7976 6248 7992 6264
rect 8044 6264 8078 6282
rect 8136 6282 8256 6329
rect 8136 6264 8170 6282
rect 8044 6248 8060 6264
rect 7976 6232 8060 6248
rect 8154 6248 8170 6264
rect 8222 6264 8256 6282
rect 8314 6282 8434 6329
rect 8314 6264 8348 6282
rect 8222 6248 8238 6264
rect 8154 6232 8238 6248
rect 8332 6248 8348 6264
rect 8400 6264 8434 6282
rect 8492 6282 8612 6329
rect 8492 6264 8526 6282
rect 8400 6248 8416 6264
rect 8332 6232 8416 6248
rect 8510 6248 8526 6264
rect 8578 6264 8612 6282
rect 8670 6282 8790 6329
rect 8670 6264 8704 6282
rect 8578 6248 8594 6264
rect 8510 6232 8594 6248
rect 8688 6248 8704 6264
rect 8756 6264 8790 6282
rect 8848 6282 8968 6329
rect 8848 6264 8882 6282
rect 8756 6248 8772 6264
rect 8688 6232 8772 6248
rect 8866 6248 8882 6264
rect 8934 6264 8968 6282
rect 9026 6282 9146 6329
rect 9026 6264 9060 6282
rect 8934 6248 8950 6264
rect 8866 6232 8950 6248
rect 9044 6248 9060 6264
rect 9112 6264 9146 6282
rect 9204 6282 9324 6329
rect 9204 6264 9238 6282
rect 9112 6248 9128 6264
rect 9044 6232 9128 6248
rect 9222 6248 9238 6264
rect 9290 6264 9324 6282
rect 9382 6282 9502 6329
rect 9382 6264 9416 6282
rect 9290 6248 9306 6264
rect 9222 6232 9306 6248
rect 9400 6248 9416 6264
rect 9468 6264 9502 6282
rect 9560 6282 9680 6329
rect 9560 6264 9594 6282
rect 9468 6248 9484 6264
rect 9400 6232 9484 6248
rect 9578 6248 9594 6264
rect 9646 6264 9680 6282
rect 9738 6282 9858 6329
rect 9738 6264 9772 6282
rect 9646 6248 9662 6264
rect 9578 6232 9662 6248
rect 9756 6248 9772 6264
rect 9824 6264 9858 6282
rect 9916 6282 10036 6329
rect 9916 6264 9950 6282
rect 9824 6248 9840 6264
rect 9756 6232 9840 6248
rect 9934 6248 9950 6264
rect 10002 6264 10036 6282
rect 10288 6282 10408 6329
rect 10288 6264 10322 6282
rect 10002 6248 10018 6264
rect 9934 6232 10018 6248
rect 10306 6248 10322 6264
rect 10374 6264 10408 6282
rect 10466 6282 10586 6329
rect 10466 6264 10500 6282
rect 10374 6248 10390 6264
rect 10306 6232 10390 6248
rect 10484 6248 10500 6264
rect 10552 6264 10586 6282
rect 10644 6282 10764 6329
rect 10644 6264 10678 6282
rect 10552 6248 10568 6264
rect 10484 6232 10568 6248
rect 10662 6248 10678 6264
rect 10730 6264 10764 6282
rect 10822 6282 10942 6329
rect 10822 6264 10856 6282
rect 10730 6248 10746 6264
rect 10662 6232 10746 6248
rect 10840 6248 10856 6264
rect 10908 6264 10942 6282
rect 11000 6282 11120 6329
rect 11000 6264 11034 6282
rect 10908 6248 10924 6264
rect 10840 6232 10924 6248
rect 11018 6248 11034 6264
rect 11086 6264 11120 6282
rect 11178 6282 11298 6329
rect 11178 6264 11212 6282
rect 11086 6248 11102 6264
rect 11018 6232 11102 6248
rect 11196 6248 11212 6264
rect 11264 6264 11298 6282
rect 11356 6282 11476 6329
rect 11356 6264 11390 6282
rect 11264 6248 11280 6264
rect 11196 6232 11280 6248
rect 11374 6248 11390 6264
rect 11442 6264 11476 6282
rect 11534 6282 11654 6329
rect 11534 6264 11568 6282
rect 11442 6248 11458 6264
rect 11374 6232 11458 6248
rect 11552 6248 11568 6264
rect 11620 6264 11654 6282
rect 11712 6282 11832 6329
rect 11712 6264 11746 6282
rect 11620 6248 11636 6264
rect 11552 6232 11636 6248
rect 11730 6248 11746 6264
rect 11798 6264 11832 6282
rect 11890 6282 12010 6329
rect 11890 6264 11924 6282
rect 11798 6248 11814 6264
rect 11730 6232 11814 6248
rect 11908 6248 11924 6264
rect 11976 6264 12010 6282
rect 12068 6282 12188 6329
rect 12068 6264 12102 6282
rect 11976 6248 11992 6264
rect 11908 6232 11992 6248
rect 12086 6248 12102 6264
rect 12154 6264 12188 6282
rect 12246 6282 12366 6329
rect 12246 6264 12280 6282
rect 12154 6248 12170 6264
rect 12086 6232 12170 6248
rect 12264 6248 12280 6264
rect 12332 6264 12366 6282
rect 12424 6282 12544 6329
rect 12424 6264 12458 6282
rect 12332 6248 12348 6264
rect 12264 6232 12348 6248
rect 12442 6248 12458 6264
rect 12510 6264 12544 6282
rect 12602 6282 12722 6329
rect 12602 6264 12636 6282
rect 12510 6248 12526 6264
rect 12442 6232 12526 6248
rect 12620 6248 12636 6264
rect 12688 6264 12722 6282
rect 12688 6248 12704 6264
rect 12620 6232 12704 6248
rect 7620 6112 7704 6128
rect 7620 6096 7636 6112
rect 7602 6078 7636 6096
rect 7688 6096 7704 6112
rect 7798 6112 7882 6128
rect 7798 6096 7814 6112
rect 7688 6078 7722 6096
rect 7602 6031 7722 6078
rect 7780 6078 7814 6096
rect 7866 6096 7882 6112
rect 7976 6112 8060 6128
rect 7976 6096 7992 6112
rect 7866 6078 7900 6096
rect 7780 6031 7900 6078
rect 7958 6078 7992 6096
rect 8044 6096 8060 6112
rect 8154 6112 8238 6128
rect 8154 6096 8170 6112
rect 8044 6078 8078 6096
rect 7958 6031 8078 6078
rect 8136 6078 8170 6096
rect 8222 6096 8238 6112
rect 8332 6112 8416 6128
rect 8332 6096 8348 6112
rect 8222 6078 8256 6096
rect 8136 6031 8256 6078
rect 8314 6078 8348 6096
rect 8400 6096 8416 6112
rect 8510 6112 8594 6128
rect 8510 6096 8526 6112
rect 8400 6078 8434 6096
rect 8314 6031 8434 6078
rect 8492 6078 8526 6096
rect 8578 6096 8594 6112
rect 8688 6112 8772 6128
rect 8688 6096 8704 6112
rect 8578 6078 8612 6096
rect 8492 6031 8612 6078
rect 8670 6078 8704 6096
rect 8756 6096 8772 6112
rect 8866 6112 8950 6128
rect 8866 6096 8882 6112
rect 8756 6078 8790 6096
rect 8670 6031 8790 6078
rect 8848 6078 8882 6096
rect 8934 6096 8950 6112
rect 9044 6112 9128 6128
rect 9044 6096 9060 6112
rect 8934 6078 8968 6096
rect 8848 6031 8968 6078
rect 9026 6078 9060 6096
rect 9112 6096 9128 6112
rect 9222 6112 9306 6128
rect 9222 6096 9238 6112
rect 9112 6078 9146 6096
rect 9026 6031 9146 6078
rect 9204 6078 9238 6096
rect 9290 6096 9306 6112
rect 9400 6112 9484 6128
rect 9400 6096 9416 6112
rect 9290 6078 9324 6096
rect 9204 6031 9324 6078
rect 9382 6078 9416 6096
rect 9468 6096 9484 6112
rect 9578 6112 9662 6128
rect 9578 6096 9594 6112
rect 9468 6078 9502 6096
rect 9382 6031 9502 6078
rect 9560 6078 9594 6096
rect 9646 6096 9662 6112
rect 9756 6112 9840 6128
rect 9756 6096 9772 6112
rect 9646 6078 9680 6096
rect 9560 6031 9680 6078
rect 9738 6078 9772 6096
rect 9824 6096 9840 6112
rect 9934 6112 10018 6128
rect 9934 6096 9950 6112
rect 9824 6078 9858 6096
rect 9738 6031 9858 6078
rect 9916 6078 9950 6096
rect 10002 6096 10018 6112
rect 10306 6113 10390 6129
rect 10306 6097 10322 6113
rect 10002 6078 10036 6096
rect 9916 6031 10036 6078
rect 10288 6079 10322 6097
rect 10374 6097 10390 6113
rect 10484 6113 10568 6129
rect 10484 6097 10500 6113
rect 10374 6079 10408 6097
rect 10288 6032 10408 6079
rect 10466 6079 10500 6097
rect 10552 6097 10568 6113
rect 10662 6113 10746 6129
rect 10662 6097 10678 6113
rect 10552 6079 10586 6097
rect 10466 6032 10586 6079
rect 10644 6079 10678 6097
rect 10730 6097 10746 6113
rect 10840 6113 10924 6129
rect 10840 6097 10856 6113
rect 10730 6079 10764 6097
rect 10644 6032 10764 6079
rect 10822 6079 10856 6097
rect 10908 6097 10924 6113
rect 11018 6113 11102 6129
rect 11018 6097 11034 6113
rect 10908 6079 10942 6097
rect 10822 6032 10942 6079
rect 11000 6079 11034 6097
rect 11086 6097 11102 6113
rect 11196 6113 11280 6129
rect 11196 6097 11212 6113
rect 11086 6079 11120 6097
rect 11000 6032 11120 6079
rect 11178 6079 11212 6097
rect 11264 6097 11280 6113
rect 11374 6113 11458 6129
rect 11374 6097 11390 6113
rect 11264 6079 11298 6097
rect 11178 6032 11298 6079
rect 11356 6079 11390 6097
rect 11442 6097 11458 6113
rect 11552 6113 11636 6129
rect 11552 6097 11568 6113
rect 11442 6079 11476 6097
rect 11356 6032 11476 6079
rect 11534 6079 11568 6097
rect 11620 6097 11636 6113
rect 11730 6113 11814 6129
rect 11730 6097 11746 6113
rect 11620 6079 11654 6097
rect 11534 6032 11654 6079
rect 11712 6079 11746 6097
rect 11798 6097 11814 6113
rect 11908 6113 11992 6129
rect 11908 6097 11924 6113
rect 11798 6079 11832 6097
rect 11712 6032 11832 6079
rect 11890 6079 11924 6097
rect 11976 6097 11992 6113
rect 12086 6113 12170 6129
rect 12086 6097 12102 6113
rect 11976 6079 12010 6097
rect 11890 6032 12010 6079
rect 12068 6079 12102 6097
rect 12154 6097 12170 6113
rect 12264 6113 12348 6129
rect 12264 6097 12280 6113
rect 12154 6079 12188 6097
rect 12068 6032 12188 6079
rect 12246 6079 12280 6097
rect 12332 6097 12348 6113
rect 12442 6113 12526 6129
rect 12442 6097 12458 6113
rect 12332 6079 12366 6097
rect 12246 6032 12366 6079
rect 12424 6079 12458 6097
rect 12510 6097 12526 6113
rect 12620 6113 12704 6129
rect 12620 6097 12636 6113
rect 12510 6079 12544 6097
rect 12424 6032 12544 6079
rect 12602 6079 12636 6097
rect 12688 6097 12704 6113
rect 12688 6079 12722 6097
rect 12602 6032 12722 6079
rect 7602 5704 7722 5751
rect 7602 5686 7636 5704
rect 7620 5670 7636 5686
rect 7688 5686 7722 5704
rect 7780 5704 7900 5751
rect 7780 5686 7814 5704
rect 7688 5670 7704 5686
rect 7620 5654 7704 5670
rect 7798 5670 7814 5686
rect 7866 5686 7900 5704
rect 7958 5704 8078 5751
rect 7958 5686 7992 5704
rect 7866 5670 7882 5686
rect 7798 5654 7882 5670
rect 7976 5670 7992 5686
rect 8044 5686 8078 5704
rect 8136 5704 8256 5751
rect 8136 5686 8170 5704
rect 8044 5670 8060 5686
rect 7976 5654 8060 5670
rect 8154 5670 8170 5686
rect 8222 5686 8256 5704
rect 8314 5704 8434 5751
rect 8314 5686 8348 5704
rect 8222 5670 8238 5686
rect 8154 5654 8238 5670
rect 8332 5670 8348 5686
rect 8400 5686 8434 5704
rect 8492 5704 8612 5751
rect 8492 5686 8526 5704
rect 8400 5670 8416 5686
rect 8332 5654 8416 5670
rect 8510 5670 8526 5686
rect 8578 5686 8612 5704
rect 8670 5704 8790 5751
rect 8670 5686 8704 5704
rect 8578 5670 8594 5686
rect 8510 5654 8594 5670
rect 8688 5670 8704 5686
rect 8756 5686 8790 5704
rect 8848 5704 8968 5751
rect 8848 5686 8882 5704
rect 8756 5670 8772 5686
rect 8688 5654 8772 5670
rect 8866 5670 8882 5686
rect 8934 5686 8968 5704
rect 9026 5704 9146 5751
rect 9026 5686 9060 5704
rect 8934 5670 8950 5686
rect 8866 5654 8950 5670
rect 9044 5670 9060 5686
rect 9112 5686 9146 5704
rect 9204 5704 9324 5751
rect 9204 5686 9238 5704
rect 9112 5670 9128 5686
rect 9044 5654 9128 5670
rect 9222 5670 9238 5686
rect 9290 5686 9324 5704
rect 9382 5704 9502 5751
rect 9382 5686 9416 5704
rect 9290 5670 9306 5686
rect 9222 5654 9306 5670
rect 9400 5670 9416 5686
rect 9468 5686 9502 5704
rect 9560 5704 9680 5751
rect 9560 5686 9594 5704
rect 9468 5670 9484 5686
rect 9400 5654 9484 5670
rect 9578 5670 9594 5686
rect 9646 5686 9680 5704
rect 9738 5704 9858 5751
rect 9738 5686 9772 5704
rect 9646 5670 9662 5686
rect 9578 5654 9662 5670
rect 9756 5670 9772 5686
rect 9824 5686 9858 5704
rect 9916 5704 10036 5751
rect 9916 5686 9950 5704
rect 9824 5670 9840 5686
rect 9756 5654 9840 5670
rect 9934 5670 9950 5686
rect 10002 5686 10036 5704
rect 10288 5705 10408 5752
rect 10288 5687 10322 5705
rect 10002 5670 10018 5686
rect 9934 5654 10018 5670
rect 10306 5671 10322 5687
rect 10374 5687 10408 5705
rect 10466 5705 10586 5752
rect 10466 5687 10500 5705
rect 10374 5671 10390 5687
rect 10306 5655 10390 5671
rect 10484 5671 10500 5687
rect 10552 5687 10586 5705
rect 10644 5705 10764 5752
rect 10644 5687 10678 5705
rect 10552 5671 10568 5687
rect 10484 5655 10568 5671
rect 10662 5671 10678 5687
rect 10730 5687 10764 5705
rect 10822 5705 10942 5752
rect 10822 5687 10856 5705
rect 10730 5671 10746 5687
rect 10662 5655 10746 5671
rect 10840 5671 10856 5687
rect 10908 5687 10942 5705
rect 11000 5705 11120 5752
rect 11000 5687 11034 5705
rect 10908 5671 10924 5687
rect 10840 5655 10924 5671
rect 11018 5671 11034 5687
rect 11086 5687 11120 5705
rect 11178 5705 11298 5752
rect 11178 5687 11212 5705
rect 11086 5671 11102 5687
rect 11018 5655 11102 5671
rect 11196 5671 11212 5687
rect 11264 5687 11298 5705
rect 11356 5705 11476 5752
rect 11356 5687 11390 5705
rect 11264 5671 11280 5687
rect 11196 5655 11280 5671
rect 11374 5671 11390 5687
rect 11442 5687 11476 5705
rect 11534 5705 11654 5752
rect 11534 5687 11568 5705
rect 11442 5671 11458 5687
rect 11374 5655 11458 5671
rect 11552 5671 11568 5687
rect 11620 5687 11654 5705
rect 11712 5705 11832 5752
rect 11712 5687 11746 5705
rect 11620 5671 11636 5687
rect 11552 5655 11636 5671
rect 11730 5671 11746 5687
rect 11798 5687 11832 5705
rect 11890 5705 12010 5752
rect 11890 5687 11924 5705
rect 11798 5671 11814 5687
rect 11730 5655 11814 5671
rect 11908 5671 11924 5687
rect 11976 5687 12010 5705
rect 12068 5705 12188 5752
rect 12068 5687 12102 5705
rect 11976 5671 11992 5687
rect 11908 5655 11992 5671
rect 12086 5671 12102 5687
rect 12154 5687 12188 5705
rect 12246 5705 12366 5752
rect 12246 5687 12280 5705
rect 12154 5671 12170 5687
rect 12086 5655 12170 5671
rect 12264 5671 12280 5687
rect 12332 5687 12366 5705
rect 12424 5705 12544 5752
rect 12424 5687 12458 5705
rect 12332 5671 12348 5687
rect 12264 5655 12348 5671
rect 12442 5671 12458 5687
rect 12510 5687 12544 5705
rect 12602 5705 12722 5752
rect 12602 5687 12636 5705
rect 12510 5671 12526 5687
rect 12442 5655 12526 5671
rect 12620 5671 12636 5687
rect 12688 5687 12722 5705
rect 12688 5671 12704 5687
rect 12620 5655 12704 5671
rect 14760 6759 14844 6775
rect 14760 6742 14776 6759
rect 14742 6725 14776 6742
rect 14828 6742 14844 6759
rect 14938 6759 15022 6775
rect 14938 6742 14954 6759
rect 14828 6725 14862 6742
rect 14742 6678 14862 6725
rect 14920 6725 14954 6742
rect 15006 6742 15022 6759
rect 15116 6759 15200 6775
rect 15116 6742 15132 6759
rect 15006 6725 15040 6742
rect 14920 6678 15040 6725
rect 15098 6725 15132 6742
rect 15184 6742 15200 6759
rect 15294 6759 15378 6775
rect 15294 6742 15310 6759
rect 15184 6725 15218 6742
rect 15098 6678 15218 6725
rect 15276 6725 15310 6742
rect 15362 6742 15378 6759
rect 15472 6759 15556 6775
rect 15472 6742 15488 6759
rect 15362 6725 15396 6742
rect 15276 6678 15396 6725
rect 15454 6725 15488 6742
rect 15540 6742 15556 6759
rect 15650 6759 15734 6775
rect 15650 6742 15666 6759
rect 15540 6725 15574 6742
rect 15454 6678 15574 6725
rect 15632 6725 15666 6742
rect 15718 6742 15734 6759
rect 15828 6759 15912 6775
rect 15828 6742 15844 6759
rect 15718 6725 15752 6742
rect 15632 6678 15752 6725
rect 15810 6725 15844 6742
rect 15896 6742 15912 6759
rect 16006 6759 16090 6775
rect 16006 6742 16022 6759
rect 15896 6725 15930 6742
rect 15810 6678 15930 6725
rect 15988 6725 16022 6742
rect 16074 6742 16090 6759
rect 16960 6759 17044 6775
rect 16960 6742 16976 6759
rect 16074 6725 16108 6742
rect 15988 6678 16108 6725
rect 16942 6725 16976 6742
rect 17028 6742 17044 6759
rect 17138 6759 17222 6775
rect 17138 6742 17154 6759
rect 17028 6725 17062 6742
rect 16942 6678 17062 6725
rect 17120 6725 17154 6742
rect 17206 6742 17222 6759
rect 17316 6759 17400 6775
rect 17316 6742 17332 6759
rect 17206 6725 17240 6742
rect 17120 6678 17240 6725
rect 17298 6725 17332 6742
rect 17384 6742 17400 6759
rect 17494 6759 17578 6775
rect 17494 6742 17510 6759
rect 17384 6725 17418 6742
rect 17298 6678 17418 6725
rect 17476 6725 17510 6742
rect 17562 6742 17578 6759
rect 17672 6759 17756 6775
rect 17672 6742 17688 6759
rect 17562 6725 17596 6742
rect 17476 6678 17596 6725
rect 17654 6725 17688 6742
rect 17740 6742 17756 6759
rect 17850 6759 17934 6775
rect 17850 6742 17866 6759
rect 17740 6725 17774 6742
rect 17654 6678 17774 6725
rect 17832 6725 17866 6742
rect 17918 6742 17934 6759
rect 18028 6759 18112 6775
rect 18028 6742 18044 6759
rect 17918 6725 17952 6742
rect 17832 6678 17952 6725
rect 18010 6725 18044 6742
rect 18096 6742 18112 6759
rect 18206 6759 18290 6775
rect 18206 6742 18222 6759
rect 18096 6725 18130 6742
rect 18010 6678 18130 6725
rect 18188 6725 18222 6742
rect 18274 6742 18290 6759
rect 19160 6759 19244 6775
rect 19160 6742 19176 6759
rect 18274 6725 18308 6742
rect 18188 6678 18308 6725
rect 19142 6725 19176 6742
rect 19228 6742 19244 6759
rect 19338 6759 19422 6775
rect 19338 6742 19354 6759
rect 19228 6725 19262 6742
rect 19142 6678 19262 6725
rect 19320 6725 19354 6742
rect 19406 6742 19422 6759
rect 19516 6759 19600 6775
rect 19516 6742 19532 6759
rect 19406 6725 19440 6742
rect 19320 6678 19440 6725
rect 19498 6725 19532 6742
rect 19584 6742 19600 6759
rect 19694 6759 19778 6775
rect 19694 6742 19710 6759
rect 19584 6725 19618 6742
rect 19498 6678 19618 6725
rect 19676 6725 19710 6742
rect 19762 6742 19778 6759
rect 19872 6759 19956 6775
rect 19872 6742 19888 6759
rect 19762 6725 19796 6742
rect 19676 6678 19796 6725
rect 19854 6725 19888 6742
rect 19940 6742 19956 6759
rect 20050 6759 20134 6775
rect 20050 6742 20066 6759
rect 19940 6725 19974 6742
rect 19854 6678 19974 6725
rect 20032 6725 20066 6742
rect 20118 6742 20134 6759
rect 20228 6759 20312 6775
rect 20228 6742 20244 6759
rect 20118 6725 20152 6742
rect 20032 6678 20152 6725
rect 20210 6725 20244 6742
rect 20296 6742 20312 6759
rect 20406 6759 20490 6775
rect 20406 6742 20422 6759
rect 20296 6725 20330 6742
rect 20210 6678 20330 6725
rect 20388 6725 20422 6742
rect 20474 6742 20490 6759
rect 20474 6725 20508 6742
rect 20388 6678 20508 6725
rect 14742 6351 14862 6398
rect 14742 6334 14776 6351
rect 14760 6317 14776 6334
rect 14828 6334 14862 6351
rect 14920 6351 15040 6398
rect 14920 6334 14954 6351
rect 14828 6317 14844 6334
rect 14760 6301 14844 6317
rect 14938 6317 14954 6334
rect 15006 6334 15040 6351
rect 15098 6351 15218 6398
rect 15098 6334 15132 6351
rect 15006 6317 15022 6334
rect 14938 6301 15022 6317
rect 15116 6317 15132 6334
rect 15184 6334 15218 6351
rect 15276 6351 15396 6398
rect 15276 6334 15310 6351
rect 15184 6317 15200 6334
rect 15116 6301 15200 6317
rect 15294 6317 15310 6334
rect 15362 6334 15396 6351
rect 15454 6351 15574 6398
rect 15454 6334 15488 6351
rect 15362 6317 15378 6334
rect 15294 6301 15378 6317
rect 15472 6317 15488 6334
rect 15540 6334 15574 6351
rect 15632 6351 15752 6398
rect 15632 6334 15666 6351
rect 15540 6317 15556 6334
rect 15472 6301 15556 6317
rect 15650 6317 15666 6334
rect 15718 6334 15752 6351
rect 15810 6351 15930 6398
rect 15810 6334 15844 6351
rect 15718 6317 15734 6334
rect 15650 6301 15734 6317
rect 15828 6317 15844 6334
rect 15896 6334 15930 6351
rect 15988 6351 16108 6398
rect 15988 6334 16022 6351
rect 15896 6317 15912 6334
rect 15828 6301 15912 6317
rect 16006 6317 16022 6334
rect 16074 6334 16108 6351
rect 16942 6351 17062 6398
rect 16942 6334 16976 6351
rect 16074 6317 16090 6334
rect 16006 6301 16090 6317
rect 16960 6317 16976 6334
rect 17028 6334 17062 6351
rect 17120 6351 17240 6398
rect 17120 6334 17154 6351
rect 17028 6317 17044 6334
rect 16960 6301 17044 6317
rect 17138 6317 17154 6334
rect 17206 6334 17240 6351
rect 17298 6351 17418 6398
rect 17298 6334 17332 6351
rect 17206 6317 17222 6334
rect 17138 6301 17222 6317
rect 17316 6317 17332 6334
rect 17384 6334 17418 6351
rect 17476 6351 17596 6398
rect 17476 6334 17510 6351
rect 17384 6317 17400 6334
rect 17316 6301 17400 6317
rect 17494 6317 17510 6334
rect 17562 6334 17596 6351
rect 17654 6351 17774 6398
rect 17654 6334 17688 6351
rect 17562 6317 17578 6334
rect 17494 6301 17578 6317
rect 17672 6317 17688 6334
rect 17740 6334 17774 6351
rect 17832 6351 17952 6398
rect 17832 6334 17866 6351
rect 17740 6317 17756 6334
rect 17672 6301 17756 6317
rect 17850 6317 17866 6334
rect 17918 6334 17952 6351
rect 18010 6351 18130 6398
rect 18010 6334 18044 6351
rect 17918 6317 17934 6334
rect 17850 6301 17934 6317
rect 18028 6317 18044 6334
rect 18096 6334 18130 6351
rect 18188 6351 18308 6398
rect 18188 6334 18222 6351
rect 18096 6317 18112 6334
rect 18028 6301 18112 6317
rect 18206 6317 18222 6334
rect 18274 6334 18308 6351
rect 19142 6351 19262 6398
rect 19142 6334 19176 6351
rect 18274 6317 18290 6334
rect 18206 6301 18290 6317
rect 19160 6317 19176 6334
rect 19228 6334 19262 6351
rect 19320 6351 19440 6398
rect 19320 6334 19354 6351
rect 19228 6317 19244 6334
rect 19160 6301 19244 6317
rect 19338 6317 19354 6334
rect 19406 6334 19440 6351
rect 19498 6351 19618 6398
rect 19498 6334 19532 6351
rect 19406 6317 19422 6334
rect 19338 6301 19422 6317
rect 19516 6317 19532 6334
rect 19584 6334 19618 6351
rect 19676 6351 19796 6398
rect 19676 6334 19710 6351
rect 19584 6317 19600 6334
rect 19516 6301 19600 6317
rect 19694 6317 19710 6334
rect 19762 6334 19796 6351
rect 19854 6351 19974 6398
rect 19854 6334 19888 6351
rect 19762 6317 19778 6334
rect 19694 6301 19778 6317
rect 19872 6317 19888 6334
rect 19940 6334 19974 6351
rect 20032 6351 20152 6398
rect 20032 6334 20066 6351
rect 19940 6317 19956 6334
rect 19872 6301 19956 6317
rect 20050 6317 20066 6334
rect 20118 6334 20152 6351
rect 20210 6351 20330 6398
rect 20210 6334 20244 6351
rect 20118 6317 20134 6334
rect 20050 6301 20134 6317
rect 20228 6317 20244 6334
rect 20296 6334 20330 6351
rect 20388 6351 20508 6398
rect 20388 6334 20422 6351
rect 20296 6317 20312 6334
rect 20228 6301 20312 6317
rect 20406 6317 20422 6334
rect 20474 6334 20508 6351
rect 20474 6317 20490 6334
rect 20406 6301 20490 6317
rect 14761 5992 14845 6008
rect 14761 5976 14777 5992
rect 14743 5958 14777 5976
rect 14829 5976 14845 5992
rect 14939 5992 15023 6008
rect 14939 5976 14955 5992
rect 14829 5958 14863 5976
rect 14743 5911 14863 5958
rect 14921 5958 14955 5976
rect 15007 5976 15023 5992
rect 15117 5992 15201 6008
rect 15117 5976 15133 5992
rect 15007 5958 15041 5976
rect 14921 5911 15041 5958
rect 15099 5958 15133 5976
rect 15185 5976 15201 5992
rect 15295 5992 15379 6008
rect 15295 5976 15311 5992
rect 15185 5958 15219 5976
rect 15099 5911 15219 5958
rect 15277 5958 15311 5976
rect 15363 5976 15379 5992
rect 15473 5992 15557 6008
rect 15473 5976 15489 5992
rect 15363 5958 15397 5976
rect 15277 5911 15397 5958
rect 15455 5958 15489 5976
rect 15541 5976 15557 5992
rect 15651 5992 15735 6008
rect 15651 5976 15667 5992
rect 15541 5958 15575 5976
rect 15455 5911 15575 5958
rect 15633 5958 15667 5976
rect 15719 5976 15735 5992
rect 15829 5992 15913 6008
rect 15829 5976 15845 5992
rect 15719 5958 15753 5976
rect 15633 5911 15753 5958
rect 15811 5958 15845 5976
rect 15897 5976 15913 5992
rect 16007 5992 16091 6008
rect 16007 5976 16023 5992
rect 15897 5958 15931 5976
rect 15811 5911 15931 5958
rect 15989 5958 16023 5976
rect 16075 5976 16091 5992
rect 16961 5992 17045 6008
rect 16961 5976 16977 5992
rect 16075 5958 16109 5976
rect 15989 5911 16109 5958
rect 16943 5958 16977 5976
rect 17029 5976 17045 5992
rect 17139 5992 17223 6008
rect 17139 5976 17155 5992
rect 17029 5958 17063 5976
rect 16943 5911 17063 5958
rect 17121 5958 17155 5976
rect 17207 5976 17223 5992
rect 17317 5992 17401 6008
rect 17317 5976 17333 5992
rect 17207 5958 17241 5976
rect 17121 5911 17241 5958
rect 17299 5958 17333 5976
rect 17385 5976 17401 5992
rect 17495 5992 17579 6008
rect 17495 5976 17511 5992
rect 17385 5958 17419 5976
rect 17299 5911 17419 5958
rect 17477 5958 17511 5976
rect 17563 5976 17579 5992
rect 17673 5992 17757 6008
rect 17673 5976 17689 5992
rect 17563 5958 17597 5976
rect 17477 5911 17597 5958
rect 17655 5958 17689 5976
rect 17741 5976 17757 5992
rect 17851 5992 17935 6008
rect 17851 5976 17867 5992
rect 17741 5958 17775 5976
rect 17655 5911 17775 5958
rect 17833 5958 17867 5976
rect 17919 5976 17935 5992
rect 18029 5992 18113 6008
rect 18029 5976 18045 5992
rect 17919 5958 17953 5976
rect 17833 5911 17953 5958
rect 18011 5958 18045 5976
rect 18097 5976 18113 5992
rect 18207 5992 18291 6008
rect 18207 5976 18223 5992
rect 18097 5958 18131 5976
rect 18011 5911 18131 5958
rect 18189 5958 18223 5976
rect 18275 5976 18291 5992
rect 19161 5992 19245 6008
rect 19161 5976 19177 5992
rect 18275 5958 18309 5976
rect 18189 5911 18309 5958
rect 19143 5958 19177 5976
rect 19229 5976 19245 5992
rect 19339 5992 19423 6008
rect 19339 5976 19355 5992
rect 19229 5958 19263 5976
rect 19143 5911 19263 5958
rect 19321 5958 19355 5976
rect 19407 5976 19423 5992
rect 19517 5992 19601 6008
rect 19517 5976 19533 5992
rect 19407 5958 19441 5976
rect 19321 5911 19441 5958
rect 19499 5958 19533 5976
rect 19585 5976 19601 5992
rect 19695 5992 19779 6008
rect 19695 5976 19711 5992
rect 19585 5958 19619 5976
rect 19499 5911 19619 5958
rect 19677 5958 19711 5976
rect 19763 5976 19779 5992
rect 19873 5992 19957 6008
rect 19873 5976 19889 5992
rect 19763 5958 19797 5976
rect 19677 5911 19797 5958
rect 19855 5958 19889 5976
rect 19941 5976 19957 5992
rect 20051 5992 20135 6008
rect 20051 5976 20067 5992
rect 19941 5958 19975 5976
rect 19855 5911 19975 5958
rect 20033 5958 20067 5976
rect 20119 5976 20135 5992
rect 20229 5992 20313 6008
rect 20229 5976 20245 5992
rect 20119 5958 20153 5976
rect 20033 5911 20153 5958
rect 20211 5958 20245 5976
rect 20297 5976 20313 5992
rect 20407 5992 20491 6008
rect 20407 5976 20423 5992
rect 20297 5958 20331 5976
rect 20211 5911 20331 5958
rect 20389 5958 20423 5976
rect 20475 5976 20491 5992
rect 20475 5958 20509 5976
rect 20389 5911 20509 5958
rect 14743 5584 14863 5631
rect 14743 5566 14777 5584
rect 14761 5550 14777 5566
rect 14829 5566 14863 5584
rect 14921 5584 15041 5631
rect 14921 5566 14955 5584
rect 14829 5550 14845 5566
rect 14761 5534 14845 5550
rect 14939 5550 14955 5566
rect 15007 5566 15041 5584
rect 15099 5584 15219 5631
rect 15099 5566 15133 5584
rect 15007 5550 15023 5566
rect 14939 5534 15023 5550
rect 15117 5550 15133 5566
rect 15185 5566 15219 5584
rect 15277 5584 15397 5631
rect 15277 5566 15311 5584
rect 15185 5550 15201 5566
rect 15117 5534 15201 5550
rect 15295 5550 15311 5566
rect 15363 5566 15397 5584
rect 15455 5584 15575 5631
rect 15455 5566 15489 5584
rect 15363 5550 15379 5566
rect 15295 5534 15379 5550
rect 15473 5550 15489 5566
rect 15541 5566 15575 5584
rect 15633 5584 15753 5631
rect 15633 5566 15667 5584
rect 15541 5550 15557 5566
rect 15473 5534 15557 5550
rect 15651 5550 15667 5566
rect 15719 5566 15753 5584
rect 15811 5584 15931 5631
rect 15811 5566 15845 5584
rect 15719 5550 15735 5566
rect 15651 5534 15735 5550
rect 15829 5550 15845 5566
rect 15897 5566 15931 5584
rect 15989 5584 16109 5631
rect 15989 5566 16023 5584
rect 15897 5550 15913 5566
rect 15829 5534 15913 5550
rect 16007 5550 16023 5566
rect 16075 5566 16109 5584
rect 16943 5584 17063 5631
rect 16943 5566 16977 5584
rect 16075 5550 16091 5566
rect 16007 5534 16091 5550
rect 16961 5550 16977 5566
rect 17029 5566 17063 5584
rect 17121 5584 17241 5631
rect 17121 5566 17155 5584
rect 17029 5550 17045 5566
rect 16961 5534 17045 5550
rect 17139 5550 17155 5566
rect 17207 5566 17241 5584
rect 17299 5584 17419 5631
rect 17299 5566 17333 5584
rect 17207 5550 17223 5566
rect 17139 5534 17223 5550
rect 17317 5550 17333 5566
rect 17385 5566 17419 5584
rect 17477 5584 17597 5631
rect 17477 5566 17511 5584
rect 17385 5550 17401 5566
rect 17317 5534 17401 5550
rect 17495 5550 17511 5566
rect 17563 5566 17597 5584
rect 17655 5584 17775 5631
rect 17655 5566 17689 5584
rect 17563 5550 17579 5566
rect 17495 5534 17579 5550
rect 17673 5550 17689 5566
rect 17741 5566 17775 5584
rect 17833 5584 17953 5631
rect 17833 5566 17867 5584
rect 17741 5550 17757 5566
rect 17673 5534 17757 5550
rect 17851 5550 17867 5566
rect 17919 5566 17953 5584
rect 18011 5584 18131 5631
rect 18011 5566 18045 5584
rect 17919 5550 17935 5566
rect 17851 5534 17935 5550
rect 18029 5550 18045 5566
rect 18097 5566 18131 5584
rect 18189 5584 18309 5631
rect 18189 5566 18223 5584
rect 18097 5550 18113 5566
rect 18029 5534 18113 5550
rect 18207 5550 18223 5566
rect 18275 5566 18309 5584
rect 19143 5584 19263 5631
rect 19143 5566 19177 5584
rect 18275 5550 18291 5566
rect 18207 5534 18291 5550
rect 19161 5550 19177 5566
rect 19229 5566 19263 5584
rect 19321 5584 19441 5631
rect 19321 5566 19355 5584
rect 19229 5550 19245 5566
rect 19161 5534 19245 5550
rect 19339 5550 19355 5566
rect 19407 5566 19441 5584
rect 19499 5584 19619 5631
rect 19499 5566 19533 5584
rect 19407 5550 19423 5566
rect 19339 5534 19423 5550
rect 19517 5550 19533 5566
rect 19585 5566 19619 5584
rect 19677 5584 19797 5631
rect 19677 5566 19711 5584
rect 19585 5550 19601 5566
rect 19517 5534 19601 5550
rect 19695 5550 19711 5566
rect 19763 5566 19797 5584
rect 19855 5584 19975 5631
rect 19855 5566 19889 5584
rect 19763 5550 19779 5566
rect 19695 5534 19779 5550
rect 19873 5550 19889 5566
rect 19941 5566 19975 5584
rect 20033 5584 20153 5631
rect 20033 5566 20067 5584
rect 19941 5550 19957 5566
rect 19873 5534 19957 5550
rect 20051 5550 20067 5566
rect 20119 5566 20153 5584
rect 20211 5584 20331 5631
rect 20211 5566 20245 5584
rect 20119 5550 20135 5566
rect 20051 5534 20135 5550
rect 20229 5550 20245 5566
rect 20297 5566 20331 5584
rect 20389 5584 20509 5631
rect 20389 5566 20423 5584
rect 20297 5550 20313 5566
rect 20229 5534 20313 5550
rect 20407 5550 20423 5566
rect 20475 5566 20509 5584
rect 20475 5550 20491 5566
rect 20407 5534 20491 5550
rect 7976 5232 8060 5248
rect 7976 5216 7992 5232
rect 7958 5198 7992 5216
rect 8044 5216 8060 5232
rect 8154 5232 8238 5248
rect 8154 5216 8170 5232
rect 8044 5198 8078 5216
rect 7958 5151 8078 5198
rect 8136 5198 8170 5216
rect 8222 5216 8238 5232
rect 8332 5232 8416 5248
rect 8332 5216 8348 5232
rect 8222 5198 8256 5216
rect 8136 5151 8256 5198
rect 8314 5198 8348 5216
rect 8400 5216 8416 5232
rect 8510 5232 8594 5248
rect 8510 5216 8526 5232
rect 8400 5198 8434 5216
rect 8314 5151 8434 5198
rect 8492 5198 8526 5216
rect 8578 5216 8594 5232
rect 8688 5232 8772 5248
rect 8688 5216 8704 5232
rect 8578 5198 8612 5216
rect 8492 5151 8612 5198
rect 8670 5198 8704 5216
rect 8756 5216 8772 5232
rect 8866 5232 8950 5248
rect 8866 5216 8882 5232
rect 8756 5198 8790 5216
rect 8670 5151 8790 5198
rect 8848 5198 8882 5216
rect 8934 5216 8950 5232
rect 9044 5232 9128 5248
rect 9044 5216 9060 5232
rect 8934 5198 8968 5216
rect 8848 5151 8968 5198
rect 9026 5198 9060 5216
rect 9112 5216 9128 5232
rect 9222 5232 9306 5248
rect 9222 5216 9238 5232
rect 9112 5198 9146 5216
rect 9026 5151 9146 5198
rect 9204 5198 9238 5216
rect 9290 5216 9306 5232
rect 9400 5232 9484 5248
rect 9400 5216 9416 5232
rect 9290 5198 9324 5216
rect 9204 5151 9324 5198
rect 9382 5198 9416 5216
rect 9468 5216 9484 5232
rect 9578 5232 9662 5248
rect 9578 5216 9594 5232
rect 9468 5198 9502 5216
rect 9382 5151 9502 5198
rect 9560 5198 9594 5216
rect 9646 5216 9662 5232
rect 9756 5232 9840 5248
rect 9756 5216 9772 5232
rect 9646 5198 9680 5216
rect 9560 5151 9680 5198
rect 9738 5198 9772 5216
rect 9824 5216 9840 5232
rect 9934 5232 10018 5248
rect 9934 5216 9950 5232
rect 9824 5198 9858 5216
rect 9738 5151 9858 5198
rect 9916 5198 9950 5216
rect 10002 5216 10018 5232
rect 10306 5232 10390 5248
rect 10306 5216 10322 5232
rect 10002 5198 10036 5216
rect 9916 5151 10036 5198
rect 10288 5198 10322 5216
rect 10374 5216 10390 5232
rect 10484 5232 10568 5248
rect 10484 5216 10500 5232
rect 10374 5198 10408 5216
rect 10288 5151 10408 5198
rect 10466 5198 10500 5216
rect 10552 5216 10568 5232
rect 10662 5232 10746 5248
rect 10662 5216 10678 5232
rect 10552 5198 10586 5216
rect 10466 5151 10586 5198
rect 10644 5198 10678 5216
rect 10730 5216 10746 5232
rect 10840 5232 10924 5248
rect 10840 5216 10856 5232
rect 10730 5198 10764 5216
rect 10644 5151 10764 5198
rect 10822 5198 10856 5216
rect 10908 5216 10924 5232
rect 11018 5232 11102 5248
rect 11018 5216 11034 5232
rect 10908 5198 10942 5216
rect 10822 5151 10942 5198
rect 11000 5198 11034 5216
rect 11086 5216 11102 5232
rect 11196 5232 11280 5248
rect 11196 5216 11212 5232
rect 11086 5198 11120 5216
rect 11000 5151 11120 5198
rect 11178 5198 11212 5216
rect 11264 5216 11280 5232
rect 11374 5232 11458 5248
rect 11374 5216 11390 5232
rect 11264 5198 11298 5216
rect 11178 5151 11298 5198
rect 11356 5198 11390 5216
rect 11442 5216 11458 5232
rect 11552 5232 11636 5248
rect 11552 5216 11568 5232
rect 11442 5198 11476 5216
rect 11356 5151 11476 5198
rect 11534 5198 11568 5216
rect 11620 5216 11636 5232
rect 11730 5232 11814 5248
rect 11730 5216 11746 5232
rect 11620 5198 11654 5216
rect 11534 5151 11654 5198
rect 11712 5198 11746 5216
rect 11798 5216 11814 5232
rect 11908 5232 11992 5248
rect 11908 5216 11924 5232
rect 11798 5198 11832 5216
rect 11712 5151 11832 5198
rect 11890 5198 11924 5216
rect 11976 5216 11992 5232
rect 12086 5232 12170 5248
rect 12086 5216 12102 5232
rect 11976 5198 12010 5216
rect 11890 5151 12010 5198
rect 12068 5198 12102 5216
rect 12154 5216 12170 5232
rect 12264 5232 12348 5248
rect 12264 5216 12280 5232
rect 12154 5198 12188 5216
rect 12068 5151 12188 5198
rect 12246 5198 12280 5216
rect 12332 5216 12348 5232
rect 12332 5198 12366 5216
rect 12246 5151 12366 5198
rect 7958 4824 8078 4871
rect 7958 4806 7992 4824
rect 7976 4790 7992 4806
rect 8044 4806 8078 4824
rect 8136 4824 8256 4871
rect 8136 4806 8170 4824
rect 8044 4790 8060 4806
rect 7976 4774 8060 4790
rect 8154 4790 8170 4806
rect 8222 4806 8256 4824
rect 8314 4824 8434 4871
rect 8314 4806 8348 4824
rect 8222 4790 8238 4806
rect 8154 4774 8238 4790
rect 8332 4790 8348 4806
rect 8400 4806 8434 4824
rect 8492 4824 8612 4871
rect 8492 4806 8526 4824
rect 8400 4790 8416 4806
rect 8332 4774 8416 4790
rect 8510 4790 8526 4806
rect 8578 4806 8612 4824
rect 8670 4824 8790 4871
rect 8670 4806 8704 4824
rect 8578 4790 8594 4806
rect 8510 4774 8594 4790
rect 8688 4790 8704 4806
rect 8756 4806 8790 4824
rect 8848 4824 8968 4871
rect 8848 4806 8882 4824
rect 8756 4790 8772 4806
rect 8688 4774 8772 4790
rect 8866 4790 8882 4806
rect 8934 4806 8968 4824
rect 9026 4824 9146 4871
rect 9026 4806 9060 4824
rect 8934 4790 8950 4806
rect 8866 4774 8950 4790
rect 9044 4790 9060 4806
rect 9112 4806 9146 4824
rect 9204 4824 9324 4871
rect 9204 4806 9238 4824
rect 9112 4790 9128 4806
rect 9044 4774 9128 4790
rect 9222 4790 9238 4806
rect 9290 4806 9324 4824
rect 9382 4824 9502 4871
rect 9382 4806 9416 4824
rect 9290 4790 9306 4806
rect 9222 4774 9306 4790
rect 9400 4790 9416 4806
rect 9468 4806 9502 4824
rect 9560 4824 9680 4871
rect 9560 4806 9594 4824
rect 9468 4790 9484 4806
rect 9400 4774 9484 4790
rect 9578 4790 9594 4806
rect 9646 4806 9680 4824
rect 9738 4824 9858 4871
rect 9738 4806 9772 4824
rect 9646 4790 9662 4806
rect 9578 4774 9662 4790
rect 9756 4790 9772 4806
rect 9824 4806 9858 4824
rect 9916 4824 10036 4871
rect 9916 4806 9950 4824
rect 9824 4790 9840 4806
rect 9756 4774 9840 4790
rect 9934 4790 9950 4806
rect 10002 4806 10036 4824
rect 10288 4824 10408 4871
rect 10288 4806 10322 4824
rect 10002 4790 10018 4806
rect 9934 4774 10018 4790
rect 10306 4790 10322 4806
rect 10374 4806 10408 4824
rect 10466 4824 10586 4871
rect 10466 4806 10500 4824
rect 10374 4790 10390 4806
rect 10306 4774 10390 4790
rect 10484 4790 10500 4806
rect 10552 4806 10586 4824
rect 10644 4824 10764 4871
rect 10644 4806 10678 4824
rect 10552 4790 10568 4806
rect 10484 4774 10568 4790
rect 10662 4790 10678 4806
rect 10730 4806 10764 4824
rect 10822 4824 10942 4871
rect 10822 4806 10856 4824
rect 10730 4790 10746 4806
rect 10662 4774 10746 4790
rect 10840 4790 10856 4806
rect 10908 4806 10942 4824
rect 11000 4824 11120 4871
rect 11000 4806 11034 4824
rect 10908 4790 10924 4806
rect 10840 4774 10924 4790
rect 11018 4790 11034 4806
rect 11086 4806 11120 4824
rect 11178 4824 11298 4871
rect 11178 4806 11212 4824
rect 11086 4790 11102 4806
rect 11018 4774 11102 4790
rect 11196 4790 11212 4806
rect 11264 4806 11298 4824
rect 11356 4824 11476 4871
rect 11356 4806 11390 4824
rect 11264 4790 11280 4806
rect 11196 4774 11280 4790
rect 11374 4790 11390 4806
rect 11442 4806 11476 4824
rect 11534 4824 11654 4871
rect 11534 4806 11568 4824
rect 11442 4790 11458 4806
rect 11374 4774 11458 4790
rect 11552 4790 11568 4806
rect 11620 4806 11654 4824
rect 11712 4824 11832 4871
rect 11712 4806 11746 4824
rect 11620 4790 11636 4806
rect 11552 4774 11636 4790
rect 11730 4790 11746 4806
rect 11798 4806 11832 4824
rect 11890 4824 12010 4871
rect 11890 4806 11924 4824
rect 11798 4790 11814 4806
rect 11730 4774 11814 4790
rect 11908 4790 11924 4806
rect 11976 4806 12010 4824
rect 12068 4824 12188 4871
rect 12068 4806 12102 4824
rect 11976 4790 11992 4806
rect 11908 4774 11992 4790
rect 12086 4790 12102 4806
rect 12154 4806 12188 4824
rect 12246 4824 12366 4871
rect 12246 4806 12280 4824
rect 12154 4790 12170 4806
rect 12086 4774 12170 4790
rect 12264 4790 12280 4806
rect 12332 4806 12366 4824
rect 12332 4790 12348 4806
rect 12264 4774 12348 4790
rect 7976 4662 8060 4678
rect 7976 4646 7992 4662
rect 7958 4628 7992 4646
rect 8044 4646 8060 4662
rect 8154 4662 8238 4678
rect 8154 4646 8170 4662
rect 8044 4628 8078 4646
rect 7958 4581 8078 4628
rect 8136 4628 8170 4646
rect 8222 4646 8238 4662
rect 8332 4662 8416 4678
rect 8332 4646 8348 4662
rect 8222 4628 8256 4646
rect 8136 4581 8256 4628
rect 8314 4628 8348 4646
rect 8400 4646 8416 4662
rect 8510 4662 8594 4678
rect 8510 4646 8526 4662
rect 8400 4628 8434 4646
rect 8314 4581 8434 4628
rect 8492 4628 8526 4646
rect 8578 4646 8594 4662
rect 8688 4662 8772 4678
rect 8688 4646 8704 4662
rect 8578 4628 8612 4646
rect 8492 4581 8612 4628
rect 8670 4628 8704 4646
rect 8756 4646 8772 4662
rect 8866 4662 8950 4678
rect 8866 4646 8882 4662
rect 8756 4628 8790 4646
rect 8670 4581 8790 4628
rect 8848 4628 8882 4646
rect 8934 4646 8950 4662
rect 9044 4662 9128 4678
rect 9044 4646 9060 4662
rect 8934 4628 8968 4646
rect 8848 4581 8968 4628
rect 9026 4628 9060 4646
rect 9112 4646 9128 4662
rect 9222 4662 9306 4678
rect 9222 4646 9238 4662
rect 9112 4628 9146 4646
rect 9026 4581 9146 4628
rect 9204 4628 9238 4646
rect 9290 4646 9306 4662
rect 9400 4662 9484 4678
rect 9400 4646 9416 4662
rect 9290 4628 9324 4646
rect 9204 4581 9324 4628
rect 9382 4628 9416 4646
rect 9468 4646 9484 4662
rect 9578 4662 9662 4678
rect 9578 4646 9594 4662
rect 9468 4628 9502 4646
rect 9382 4581 9502 4628
rect 9560 4628 9594 4646
rect 9646 4646 9662 4662
rect 9756 4662 9840 4678
rect 9756 4646 9772 4662
rect 9646 4628 9680 4646
rect 9560 4581 9680 4628
rect 9738 4628 9772 4646
rect 9824 4646 9840 4662
rect 9934 4662 10018 4678
rect 9934 4646 9950 4662
rect 9824 4628 9858 4646
rect 9738 4581 9858 4628
rect 9916 4628 9950 4646
rect 10002 4646 10018 4662
rect 10306 4662 10390 4678
rect 10306 4646 10322 4662
rect 10002 4628 10036 4646
rect 9916 4581 10036 4628
rect 10288 4628 10322 4646
rect 10374 4646 10390 4662
rect 10484 4662 10568 4678
rect 10484 4646 10500 4662
rect 10374 4628 10408 4646
rect 10288 4581 10408 4628
rect 10466 4628 10500 4646
rect 10552 4646 10568 4662
rect 10662 4662 10746 4678
rect 10662 4646 10678 4662
rect 10552 4628 10586 4646
rect 10466 4581 10586 4628
rect 10644 4628 10678 4646
rect 10730 4646 10746 4662
rect 10840 4662 10924 4678
rect 10840 4646 10856 4662
rect 10730 4628 10764 4646
rect 10644 4581 10764 4628
rect 10822 4628 10856 4646
rect 10908 4646 10924 4662
rect 11018 4662 11102 4678
rect 11018 4646 11034 4662
rect 10908 4628 10942 4646
rect 10822 4581 10942 4628
rect 11000 4628 11034 4646
rect 11086 4646 11102 4662
rect 11196 4662 11280 4678
rect 11196 4646 11212 4662
rect 11086 4628 11120 4646
rect 11000 4581 11120 4628
rect 11178 4628 11212 4646
rect 11264 4646 11280 4662
rect 11374 4662 11458 4678
rect 11374 4646 11390 4662
rect 11264 4628 11298 4646
rect 11178 4581 11298 4628
rect 11356 4628 11390 4646
rect 11442 4646 11458 4662
rect 11552 4662 11636 4678
rect 11552 4646 11568 4662
rect 11442 4628 11476 4646
rect 11356 4581 11476 4628
rect 11534 4628 11568 4646
rect 11620 4646 11636 4662
rect 11730 4662 11814 4678
rect 11730 4646 11746 4662
rect 11620 4628 11654 4646
rect 11534 4581 11654 4628
rect 11712 4628 11746 4646
rect 11798 4646 11814 4662
rect 11908 4662 11992 4678
rect 11908 4646 11924 4662
rect 11798 4628 11832 4646
rect 11712 4581 11832 4628
rect 11890 4628 11924 4646
rect 11976 4646 11992 4662
rect 12086 4662 12170 4678
rect 12086 4646 12102 4662
rect 11976 4628 12010 4646
rect 11890 4581 12010 4628
rect 12068 4628 12102 4646
rect 12154 4646 12170 4662
rect 12264 4662 12348 4678
rect 12264 4646 12280 4662
rect 12154 4628 12188 4646
rect 12068 4581 12188 4628
rect 12246 4628 12280 4646
rect 12332 4646 12348 4662
rect 12332 4628 12366 4646
rect 12246 4581 12366 4628
rect 7958 4254 8078 4301
rect 7958 4236 7992 4254
rect 7976 4220 7992 4236
rect 8044 4236 8078 4254
rect 8136 4254 8256 4301
rect 8136 4236 8170 4254
rect 8044 4220 8060 4236
rect 7976 4204 8060 4220
rect 8154 4220 8170 4236
rect 8222 4236 8256 4254
rect 8314 4254 8434 4301
rect 8314 4236 8348 4254
rect 8222 4220 8238 4236
rect 8154 4204 8238 4220
rect 8332 4220 8348 4236
rect 8400 4236 8434 4254
rect 8492 4254 8612 4301
rect 8492 4236 8526 4254
rect 8400 4220 8416 4236
rect 8332 4204 8416 4220
rect 8510 4220 8526 4236
rect 8578 4236 8612 4254
rect 8670 4254 8790 4301
rect 8670 4236 8704 4254
rect 8578 4220 8594 4236
rect 8510 4204 8594 4220
rect 8688 4220 8704 4236
rect 8756 4236 8790 4254
rect 8848 4254 8968 4301
rect 8848 4236 8882 4254
rect 8756 4220 8772 4236
rect 8688 4204 8772 4220
rect 8866 4220 8882 4236
rect 8934 4236 8968 4254
rect 9026 4254 9146 4301
rect 9026 4236 9060 4254
rect 8934 4220 8950 4236
rect 8866 4204 8950 4220
rect 9044 4220 9060 4236
rect 9112 4236 9146 4254
rect 9204 4254 9324 4301
rect 9204 4236 9238 4254
rect 9112 4220 9128 4236
rect 9044 4204 9128 4220
rect 9222 4220 9238 4236
rect 9290 4236 9324 4254
rect 9382 4254 9502 4301
rect 9382 4236 9416 4254
rect 9290 4220 9306 4236
rect 9222 4204 9306 4220
rect 9400 4220 9416 4236
rect 9468 4236 9502 4254
rect 9560 4254 9680 4301
rect 9560 4236 9594 4254
rect 9468 4220 9484 4236
rect 9400 4204 9484 4220
rect 9578 4220 9594 4236
rect 9646 4236 9680 4254
rect 9738 4254 9858 4301
rect 9738 4236 9772 4254
rect 9646 4220 9662 4236
rect 9578 4204 9662 4220
rect 9756 4220 9772 4236
rect 9824 4236 9858 4254
rect 9916 4254 10036 4301
rect 9916 4236 9950 4254
rect 9824 4220 9840 4236
rect 9756 4204 9840 4220
rect 9934 4220 9950 4236
rect 10002 4236 10036 4254
rect 10288 4254 10408 4301
rect 10288 4236 10322 4254
rect 10002 4220 10018 4236
rect 9934 4204 10018 4220
rect 10306 4220 10322 4236
rect 10374 4236 10408 4254
rect 10466 4254 10586 4301
rect 10466 4236 10500 4254
rect 10374 4220 10390 4236
rect 10306 4204 10390 4220
rect 10484 4220 10500 4236
rect 10552 4236 10586 4254
rect 10644 4254 10764 4301
rect 10644 4236 10678 4254
rect 10552 4220 10568 4236
rect 10484 4204 10568 4220
rect 10662 4220 10678 4236
rect 10730 4236 10764 4254
rect 10822 4254 10942 4301
rect 10822 4236 10856 4254
rect 10730 4220 10746 4236
rect 10662 4204 10746 4220
rect 10840 4220 10856 4236
rect 10908 4236 10942 4254
rect 11000 4254 11120 4301
rect 11000 4236 11034 4254
rect 10908 4220 10924 4236
rect 10840 4204 10924 4220
rect 11018 4220 11034 4236
rect 11086 4236 11120 4254
rect 11178 4254 11298 4301
rect 11178 4236 11212 4254
rect 11086 4220 11102 4236
rect 11018 4204 11102 4220
rect 11196 4220 11212 4236
rect 11264 4236 11298 4254
rect 11356 4254 11476 4301
rect 11356 4236 11390 4254
rect 11264 4220 11280 4236
rect 11196 4204 11280 4220
rect 11374 4220 11390 4236
rect 11442 4236 11476 4254
rect 11534 4254 11654 4301
rect 11534 4236 11568 4254
rect 11442 4220 11458 4236
rect 11374 4204 11458 4220
rect 11552 4220 11568 4236
rect 11620 4236 11654 4254
rect 11712 4254 11832 4301
rect 11712 4236 11746 4254
rect 11620 4220 11636 4236
rect 11552 4204 11636 4220
rect 11730 4220 11746 4236
rect 11798 4236 11832 4254
rect 11890 4254 12010 4301
rect 11890 4236 11924 4254
rect 11798 4220 11814 4236
rect 11730 4204 11814 4220
rect 11908 4220 11924 4236
rect 11976 4236 12010 4254
rect 12068 4254 12188 4301
rect 12068 4236 12102 4254
rect 11976 4220 11992 4236
rect 11908 4204 11992 4220
rect 12086 4220 12102 4236
rect 12154 4236 12188 4254
rect 12246 4254 12366 4301
rect 12246 4236 12280 4254
rect 12154 4220 12170 4236
rect 12086 4204 12170 4220
rect 12264 4220 12280 4236
rect 12332 4236 12366 4254
rect 12332 4220 12348 4236
rect 12264 4204 12348 4220
rect 7621 3723 7705 3739
rect 7621 3706 7637 3723
rect 7603 3689 7637 3706
rect 7689 3706 7705 3723
rect 7799 3723 7883 3739
rect 7799 3706 7815 3723
rect 7689 3689 7723 3706
rect 7603 3651 7723 3689
rect 7781 3689 7815 3706
rect 7867 3706 7883 3723
rect 7977 3723 8061 3739
rect 7977 3706 7993 3723
rect 7867 3689 7901 3706
rect 7781 3651 7901 3689
rect 7959 3689 7993 3706
rect 8045 3706 8061 3723
rect 8155 3723 8239 3739
rect 8155 3706 8171 3723
rect 8045 3689 8079 3706
rect 7959 3651 8079 3689
rect 8137 3689 8171 3706
rect 8223 3706 8239 3723
rect 8333 3723 8417 3739
rect 8333 3706 8349 3723
rect 8223 3689 8257 3706
rect 8137 3651 8257 3689
rect 8315 3689 8349 3706
rect 8401 3706 8417 3723
rect 8511 3723 8595 3739
rect 8511 3706 8527 3723
rect 8401 3689 8435 3706
rect 8315 3651 8435 3689
rect 8493 3689 8527 3706
rect 8579 3706 8595 3723
rect 8689 3723 8773 3739
rect 8689 3706 8705 3723
rect 8579 3689 8613 3706
rect 8493 3651 8613 3689
rect 8671 3689 8705 3706
rect 8757 3706 8773 3723
rect 8867 3723 8951 3739
rect 8867 3706 8883 3723
rect 8757 3689 8791 3706
rect 8671 3651 8791 3689
rect 8849 3689 8883 3706
rect 8935 3706 8951 3723
rect 9045 3723 9129 3739
rect 9045 3706 9061 3723
rect 8935 3689 8969 3706
rect 8849 3651 8969 3689
rect 9027 3689 9061 3706
rect 9113 3706 9129 3723
rect 9223 3723 9307 3739
rect 9223 3706 9239 3723
rect 9113 3689 9147 3706
rect 9027 3651 9147 3689
rect 9205 3689 9239 3706
rect 9291 3706 9307 3723
rect 9401 3723 9485 3739
rect 9401 3706 9417 3723
rect 9291 3689 9325 3706
rect 9205 3651 9325 3689
rect 9383 3689 9417 3706
rect 9469 3706 9485 3723
rect 9579 3723 9663 3739
rect 9579 3706 9595 3723
rect 9469 3689 9503 3706
rect 9383 3651 9503 3689
rect 9561 3689 9595 3706
rect 9647 3706 9663 3723
rect 9757 3723 9841 3739
rect 9757 3706 9773 3723
rect 9647 3689 9681 3706
rect 9561 3651 9681 3689
rect 9739 3689 9773 3706
rect 9825 3706 9841 3723
rect 9935 3723 10019 3739
rect 9935 3706 9951 3723
rect 9825 3689 9859 3706
rect 9739 3651 9859 3689
rect 9917 3689 9951 3706
rect 10003 3706 10019 3723
rect 10308 3723 10392 3739
rect 10308 3706 10324 3723
rect 10003 3689 10037 3706
rect 9917 3651 10037 3689
rect 10290 3689 10324 3706
rect 10376 3706 10392 3723
rect 10486 3723 10570 3739
rect 10486 3706 10502 3723
rect 10376 3689 10410 3706
rect 10290 3651 10410 3689
rect 10468 3689 10502 3706
rect 10554 3706 10570 3723
rect 10664 3723 10748 3739
rect 10664 3706 10680 3723
rect 10554 3689 10588 3706
rect 10468 3651 10588 3689
rect 10646 3689 10680 3706
rect 10732 3706 10748 3723
rect 10842 3723 10926 3739
rect 10842 3706 10858 3723
rect 10732 3689 10766 3706
rect 10646 3651 10766 3689
rect 10824 3689 10858 3706
rect 10910 3706 10926 3723
rect 11020 3723 11104 3739
rect 11020 3706 11036 3723
rect 10910 3689 10944 3706
rect 10824 3651 10944 3689
rect 11002 3689 11036 3706
rect 11088 3706 11104 3723
rect 11198 3723 11282 3739
rect 11198 3706 11214 3723
rect 11088 3689 11122 3706
rect 11002 3651 11122 3689
rect 11180 3689 11214 3706
rect 11266 3706 11282 3723
rect 11376 3723 11460 3739
rect 11376 3706 11392 3723
rect 11266 3689 11300 3706
rect 11180 3651 11300 3689
rect 11358 3689 11392 3706
rect 11444 3706 11460 3723
rect 11554 3723 11638 3739
rect 11554 3706 11570 3723
rect 11444 3689 11478 3706
rect 11358 3651 11478 3689
rect 11536 3689 11570 3706
rect 11622 3706 11638 3723
rect 11732 3723 11816 3739
rect 11732 3706 11748 3723
rect 11622 3689 11656 3706
rect 11536 3651 11656 3689
rect 11714 3689 11748 3706
rect 11800 3706 11816 3723
rect 11910 3723 11994 3739
rect 11910 3706 11926 3723
rect 11800 3689 11834 3706
rect 11714 3651 11834 3689
rect 11892 3689 11926 3706
rect 11978 3706 11994 3723
rect 12088 3723 12172 3739
rect 12088 3706 12104 3723
rect 11978 3689 12012 3706
rect 11892 3651 12012 3689
rect 12070 3689 12104 3706
rect 12156 3706 12172 3723
rect 12266 3723 12350 3739
rect 12266 3706 12282 3723
rect 12156 3689 12190 3706
rect 12070 3651 12190 3689
rect 12248 3689 12282 3706
rect 12334 3706 12350 3723
rect 12444 3723 12528 3739
rect 12444 3706 12460 3723
rect 12334 3689 12368 3706
rect 12248 3651 12368 3689
rect 12426 3689 12460 3706
rect 12512 3706 12528 3723
rect 12622 3723 12706 3739
rect 12622 3706 12638 3723
rect 12512 3689 12546 3706
rect 12426 3651 12546 3689
rect 12604 3689 12638 3706
rect 12690 3706 12706 3723
rect 12690 3689 12724 3706
rect 12604 3651 12724 3689
rect 492 3523 576 3539
rect 492 3505 508 3523
rect 474 3489 508 3505
rect 560 3505 576 3523
rect 670 3523 754 3539
rect 670 3505 686 3523
rect 560 3489 594 3505
rect 474 3451 594 3489
rect 652 3489 686 3505
rect 738 3505 754 3523
rect 848 3523 932 3539
rect 848 3505 864 3523
rect 738 3489 772 3505
rect 652 3451 772 3489
rect 830 3489 864 3505
rect 916 3505 932 3523
rect 1026 3523 1110 3539
rect 1026 3505 1042 3523
rect 916 3489 950 3505
rect 830 3451 950 3489
rect 1008 3489 1042 3505
rect 1094 3505 1110 3523
rect 1204 3523 1288 3539
rect 1204 3505 1220 3523
rect 1094 3489 1128 3505
rect 1008 3451 1128 3489
rect 1186 3489 1220 3505
rect 1272 3505 1288 3523
rect 1382 3523 1466 3539
rect 1382 3505 1398 3523
rect 1272 3489 1306 3505
rect 1186 3451 1306 3489
rect 1364 3489 1398 3505
rect 1450 3505 1466 3523
rect 1560 3523 1644 3539
rect 1560 3505 1576 3523
rect 1450 3489 1484 3505
rect 1364 3451 1484 3489
rect 1542 3489 1576 3505
rect 1628 3505 1644 3523
rect 1738 3523 1822 3539
rect 1738 3505 1754 3523
rect 1628 3489 1662 3505
rect 1542 3451 1662 3489
rect 1720 3489 1754 3505
rect 1806 3505 1822 3523
rect 1916 3523 2000 3539
rect 1916 3505 1932 3523
rect 1806 3489 1840 3505
rect 1720 3451 1840 3489
rect 1898 3489 1932 3505
rect 1984 3505 2000 3523
rect 2094 3523 2178 3539
rect 2094 3505 2110 3523
rect 1984 3489 2018 3505
rect 1898 3451 2018 3489
rect 2076 3489 2110 3505
rect 2162 3505 2178 3523
rect 2272 3523 2356 3539
rect 2272 3505 2288 3523
rect 2162 3489 2196 3505
rect 2076 3451 2196 3489
rect 2254 3489 2288 3505
rect 2340 3505 2356 3523
rect 2450 3523 2534 3539
rect 2450 3505 2466 3523
rect 2340 3489 2374 3505
rect 2254 3451 2374 3489
rect 2432 3489 2466 3505
rect 2518 3505 2534 3523
rect 2628 3523 2712 3539
rect 2628 3505 2644 3523
rect 2518 3489 2552 3505
rect 2432 3451 2552 3489
rect 2610 3489 2644 3505
rect 2696 3505 2712 3523
rect 2806 3523 2890 3539
rect 2806 3505 2822 3523
rect 2696 3489 2730 3505
rect 2610 3451 2730 3489
rect 2788 3489 2822 3505
rect 2874 3505 2890 3523
rect 2984 3523 3068 3539
rect 2984 3505 3000 3523
rect 2874 3489 2908 3505
rect 2788 3451 2908 3489
rect 2966 3489 3000 3505
rect 3052 3505 3068 3523
rect 3162 3523 3246 3539
rect 3162 3505 3178 3523
rect 3052 3489 3086 3505
rect 2966 3451 3086 3489
rect 3144 3489 3178 3505
rect 3230 3505 3246 3523
rect 3340 3523 3424 3539
rect 3340 3505 3356 3523
rect 3230 3489 3264 3505
rect 3144 3451 3264 3489
rect 3322 3489 3356 3505
rect 3408 3505 3424 3523
rect 3518 3523 3602 3539
rect 3518 3505 3534 3523
rect 3408 3489 3442 3505
rect 3322 3451 3442 3489
rect 3500 3489 3534 3505
rect 3586 3505 3602 3523
rect 3892 3523 3976 3539
rect 3892 3505 3908 3523
rect 3586 3489 3620 3505
rect 3500 3451 3620 3489
rect 3874 3489 3908 3505
rect 3960 3505 3976 3523
rect 4070 3523 4154 3539
rect 4070 3505 4086 3523
rect 3960 3489 3994 3505
rect 3874 3451 3994 3489
rect 4052 3489 4086 3505
rect 4138 3505 4154 3523
rect 4248 3523 4332 3539
rect 4248 3505 4264 3523
rect 4138 3489 4172 3505
rect 4052 3451 4172 3489
rect 4230 3489 4264 3505
rect 4316 3505 4332 3523
rect 4426 3523 4510 3539
rect 4426 3505 4442 3523
rect 4316 3489 4350 3505
rect 4230 3451 4350 3489
rect 4408 3489 4442 3505
rect 4494 3505 4510 3523
rect 4604 3523 4688 3539
rect 4604 3505 4620 3523
rect 4494 3489 4528 3505
rect 4408 3451 4528 3489
rect 4586 3489 4620 3505
rect 4672 3505 4688 3523
rect 4782 3523 4866 3539
rect 4782 3505 4798 3523
rect 4672 3489 4706 3505
rect 4586 3451 4706 3489
rect 4764 3489 4798 3505
rect 4850 3505 4866 3523
rect 4960 3523 5044 3539
rect 4960 3505 4976 3523
rect 4850 3489 4884 3505
rect 4764 3451 4884 3489
rect 4942 3489 4976 3505
rect 5028 3505 5044 3523
rect 5138 3523 5222 3539
rect 5138 3505 5154 3523
rect 5028 3489 5062 3505
rect 4942 3451 5062 3489
rect 5120 3489 5154 3505
rect 5206 3505 5222 3523
rect 5316 3523 5400 3539
rect 5316 3505 5332 3523
rect 5206 3489 5240 3505
rect 5120 3451 5240 3489
rect 5298 3489 5332 3505
rect 5384 3505 5400 3523
rect 5494 3523 5578 3539
rect 5494 3505 5510 3523
rect 5384 3489 5418 3505
rect 5298 3451 5418 3489
rect 5476 3489 5510 3505
rect 5562 3505 5578 3523
rect 5672 3523 5756 3539
rect 5672 3505 5688 3523
rect 5562 3489 5596 3505
rect 5476 3451 5596 3489
rect 5654 3489 5688 3505
rect 5740 3505 5756 3523
rect 5850 3523 5934 3539
rect 5850 3505 5866 3523
rect 5740 3489 5774 3505
rect 5654 3451 5774 3489
rect 5832 3489 5866 3505
rect 5918 3505 5934 3523
rect 6028 3523 6112 3539
rect 6028 3505 6044 3523
rect 5918 3489 5952 3505
rect 5832 3451 5952 3489
rect 6010 3489 6044 3505
rect 6096 3505 6112 3523
rect 6206 3523 6290 3539
rect 6206 3505 6222 3523
rect 6096 3489 6130 3505
rect 6010 3451 6130 3489
rect 6188 3489 6222 3505
rect 6274 3505 6290 3523
rect 6384 3523 6468 3539
rect 6384 3505 6400 3523
rect 6274 3489 6308 3505
rect 6188 3451 6308 3489
rect 6366 3489 6400 3505
rect 6452 3505 6468 3523
rect 6562 3523 6646 3539
rect 6562 3505 6578 3523
rect 6452 3489 6486 3505
rect 6366 3451 6486 3489
rect 6544 3489 6578 3505
rect 6630 3505 6646 3523
rect 6740 3523 6824 3539
rect 6740 3505 6756 3523
rect 6630 3489 6664 3505
rect 6544 3451 6664 3489
rect 6722 3489 6756 3505
rect 6808 3505 6824 3523
rect 6918 3523 7002 3539
rect 6918 3505 6934 3523
rect 6808 3489 6842 3505
rect 6722 3451 6842 3489
rect 6900 3489 6934 3505
rect 6986 3505 7002 3523
rect 6986 3489 7020 3505
rect 6900 3451 7020 3489
rect 7603 3333 7723 3371
rect 7603 3316 7637 3333
rect 7621 3299 7637 3316
rect 7689 3316 7723 3333
rect 7781 3333 7901 3371
rect 7781 3316 7815 3333
rect 7689 3299 7705 3316
rect 7621 3283 7705 3299
rect 7799 3299 7815 3316
rect 7867 3316 7901 3333
rect 7959 3333 8079 3371
rect 7959 3316 7993 3333
rect 7867 3299 7883 3316
rect 7799 3283 7883 3299
rect 7977 3299 7993 3316
rect 8045 3316 8079 3333
rect 8137 3333 8257 3371
rect 8137 3316 8171 3333
rect 8045 3299 8061 3316
rect 7977 3283 8061 3299
rect 8155 3299 8171 3316
rect 8223 3316 8257 3333
rect 8315 3333 8435 3371
rect 8315 3316 8349 3333
rect 8223 3299 8239 3316
rect 8155 3283 8239 3299
rect 8333 3299 8349 3316
rect 8401 3316 8435 3333
rect 8493 3333 8613 3371
rect 8493 3316 8527 3333
rect 8401 3299 8417 3316
rect 8333 3283 8417 3299
rect 8511 3299 8527 3316
rect 8579 3316 8613 3333
rect 8671 3333 8791 3371
rect 8671 3316 8705 3333
rect 8579 3299 8595 3316
rect 8511 3283 8595 3299
rect 8689 3299 8705 3316
rect 8757 3316 8791 3333
rect 8849 3333 8969 3371
rect 8849 3316 8883 3333
rect 8757 3299 8773 3316
rect 8689 3283 8773 3299
rect 8867 3299 8883 3316
rect 8935 3316 8969 3333
rect 9027 3333 9147 3371
rect 9027 3316 9061 3333
rect 8935 3299 8951 3316
rect 8867 3283 8951 3299
rect 9045 3299 9061 3316
rect 9113 3316 9147 3333
rect 9205 3333 9325 3371
rect 9205 3316 9239 3333
rect 9113 3299 9129 3316
rect 9045 3283 9129 3299
rect 9223 3299 9239 3316
rect 9291 3316 9325 3333
rect 9383 3333 9503 3371
rect 9383 3316 9417 3333
rect 9291 3299 9307 3316
rect 9223 3283 9307 3299
rect 9401 3299 9417 3316
rect 9469 3316 9503 3333
rect 9561 3333 9681 3371
rect 9561 3316 9595 3333
rect 9469 3299 9485 3316
rect 9401 3283 9485 3299
rect 9579 3299 9595 3316
rect 9647 3316 9681 3333
rect 9739 3333 9859 3371
rect 9739 3316 9773 3333
rect 9647 3299 9663 3316
rect 9579 3283 9663 3299
rect 9757 3299 9773 3316
rect 9825 3316 9859 3333
rect 9917 3333 10037 3371
rect 9917 3316 9951 3333
rect 9825 3299 9841 3316
rect 9757 3283 9841 3299
rect 9935 3299 9951 3316
rect 10003 3316 10037 3333
rect 10290 3333 10410 3371
rect 10290 3316 10324 3333
rect 10003 3299 10019 3316
rect 9935 3283 10019 3299
rect 10308 3299 10324 3316
rect 10376 3316 10410 3333
rect 10468 3333 10588 3371
rect 10468 3316 10502 3333
rect 10376 3299 10392 3316
rect 10308 3283 10392 3299
rect 10486 3299 10502 3316
rect 10554 3316 10588 3333
rect 10646 3333 10766 3371
rect 10646 3316 10680 3333
rect 10554 3299 10570 3316
rect 10486 3283 10570 3299
rect 10664 3299 10680 3316
rect 10732 3316 10766 3333
rect 10824 3333 10944 3371
rect 10824 3316 10858 3333
rect 10732 3299 10748 3316
rect 10664 3283 10748 3299
rect 10842 3299 10858 3316
rect 10910 3316 10944 3333
rect 11002 3333 11122 3371
rect 11002 3316 11036 3333
rect 10910 3299 10926 3316
rect 10842 3283 10926 3299
rect 11020 3299 11036 3316
rect 11088 3316 11122 3333
rect 11180 3333 11300 3371
rect 11180 3316 11214 3333
rect 11088 3299 11104 3316
rect 11020 3283 11104 3299
rect 11198 3299 11214 3316
rect 11266 3316 11300 3333
rect 11358 3333 11478 3371
rect 11358 3316 11392 3333
rect 11266 3299 11282 3316
rect 11198 3283 11282 3299
rect 11376 3299 11392 3316
rect 11444 3316 11478 3333
rect 11536 3333 11656 3371
rect 11536 3316 11570 3333
rect 11444 3299 11460 3316
rect 11376 3283 11460 3299
rect 11554 3299 11570 3316
rect 11622 3316 11656 3333
rect 11714 3333 11834 3371
rect 11714 3316 11748 3333
rect 11622 3299 11638 3316
rect 11554 3283 11638 3299
rect 11732 3299 11748 3316
rect 11800 3316 11834 3333
rect 11892 3333 12012 3371
rect 11892 3316 11926 3333
rect 11800 3299 11816 3316
rect 11732 3283 11816 3299
rect 11910 3299 11926 3316
rect 11978 3316 12012 3333
rect 12070 3333 12190 3371
rect 12070 3316 12104 3333
rect 11978 3299 11994 3316
rect 11910 3283 11994 3299
rect 12088 3299 12104 3316
rect 12156 3316 12190 3333
rect 12248 3333 12368 3371
rect 12248 3316 12282 3333
rect 12156 3299 12172 3316
rect 12088 3283 12172 3299
rect 12266 3299 12282 3316
rect 12334 3316 12368 3333
rect 12426 3333 12546 3371
rect 12426 3316 12460 3333
rect 12334 3299 12350 3316
rect 12266 3283 12350 3299
rect 12444 3299 12460 3316
rect 12512 3316 12546 3333
rect 12604 3333 12724 3371
rect 12604 3316 12638 3333
rect 12512 3299 12528 3316
rect 12444 3283 12528 3299
rect 12622 3299 12638 3316
rect 12690 3316 12724 3333
rect 12690 3299 12706 3316
rect 12622 3283 12706 3299
rect 7621 3223 7705 3239
rect 7621 3206 7637 3223
rect 7603 3189 7637 3206
rect 7689 3206 7705 3223
rect 7799 3223 7883 3239
rect 7799 3206 7815 3223
rect 7689 3189 7723 3206
rect 474 3133 594 3171
rect 474 3117 508 3133
rect 492 3099 508 3117
rect 560 3117 594 3133
rect 652 3133 772 3171
rect 652 3117 686 3133
rect 560 3099 576 3117
rect 492 3083 576 3099
rect 670 3099 686 3117
rect 738 3117 772 3133
rect 830 3133 950 3171
rect 830 3117 864 3133
rect 738 3099 754 3117
rect 670 3083 754 3099
rect 848 3099 864 3117
rect 916 3117 950 3133
rect 1008 3133 1128 3171
rect 1008 3117 1042 3133
rect 916 3099 932 3117
rect 848 3083 932 3099
rect 1026 3099 1042 3117
rect 1094 3117 1128 3133
rect 1186 3133 1306 3171
rect 1186 3117 1220 3133
rect 1094 3099 1110 3117
rect 1026 3083 1110 3099
rect 1204 3099 1220 3117
rect 1272 3117 1306 3133
rect 1364 3133 1484 3171
rect 1364 3117 1398 3133
rect 1272 3099 1288 3117
rect 1204 3083 1288 3099
rect 1382 3099 1398 3117
rect 1450 3117 1484 3133
rect 1542 3133 1662 3171
rect 1542 3117 1576 3133
rect 1450 3099 1466 3117
rect 1382 3083 1466 3099
rect 1560 3099 1576 3117
rect 1628 3117 1662 3133
rect 1720 3133 1840 3171
rect 1720 3117 1754 3133
rect 1628 3099 1644 3117
rect 1560 3083 1644 3099
rect 1738 3099 1754 3117
rect 1806 3117 1840 3133
rect 1898 3133 2018 3171
rect 1898 3117 1932 3133
rect 1806 3099 1822 3117
rect 1738 3083 1822 3099
rect 1916 3099 1932 3117
rect 1984 3117 2018 3133
rect 2076 3133 2196 3171
rect 2076 3117 2110 3133
rect 1984 3099 2000 3117
rect 1916 3083 2000 3099
rect 2094 3099 2110 3117
rect 2162 3117 2196 3133
rect 2254 3133 2374 3171
rect 2254 3117 2288 3133
rect 2162 3099 2178 3117
rect 2094 3083 2178 3099
rect 2272 3099 2288 3117
rect 2340 3117 2374 3133
rect 2432 3133 2552 3171
rect 2432 3117 2466 3133
rect 2340 3099 2356 3117
rect 2272 3083 2356 3099
rect 2450 3099 2466 3117
rect 2518 3117 2552 3133
rect 2610 3133 2730 3171
rect 2610 3117 2644 3133
rect 2518 3099 2534 3117
rect 2450 3083 2534 3099
rect 2628 3099 2644 3117
rect 2696 3117 2730 3133
rect 2788 3133 2908 3171
rect 2788 3117 2822 3133
rect 2696 3099 2712 3117
rect 2628 3083 2712 3099
rect 2806 3099 2822 3117
rect 2874 3117 2908 3133
rect 2966 3133 3086 3171
rect 2966 3117 3000 3133
rect 2874 3099 2890 3117
rect 2806 3083 2890 3099
rect 2984 3099 3000 3117
rect 3052 3117 3086 3133
rect 3144 3133 3264 3171
rect 3144 3117 3178 3133
rect 3052 3099 3068 3117
rect 2984 3083 3068 3099
rect 3162 3099 3178 3117
rect 3230 3117 3264 3133
rect 3322 3133 3442 3171
rect 3322 3117 3356 3133
rect 3230 3099 3246 3117
rect 3162 3083 3246 3099
rect 3340 3099 3356 3117
rect 3408 3117 3442 3133
rect 3500 3133 3620 3171
rect 3500 3117 3534 3133
rect 3408 3099 3424 3117
rect 3340 3083 3424 3099
rect 3518 3099 3534 3117
rect 3586 3117 3620 3133
rect 3874 3133 3994 3171
rect 3874 3117 3908 3133
rect 3586 3099 3602 3117
rect 3518 3083 3602 3099
rect 3892 3099 3908 3117
rect 3960 3117 3994 3133
rect 4052 3133 4172 3171
rect 4052 3117 4086 3133
rect 3960 3099 3976 3117
rect 3892 3083 3976 3099
rect 4070 3099 4086 3117
rect 4138 3117 4172 3133
rect 4230 3133 4350 3171
rect 4230 3117 4264 3133
rect 4138 3099 4154 3117
rect 4070 3083 4154 3099
rect 4248 3099 4264 3117
rect 4316 3117 4350 3133
rect 4408 3133 4528 3171
rect 4408 3117 4442 3133
rect 4316 3099 4332 3117
rect 4248 3083 4332 3099
rect 4426 3099 4442 3117
rect 4494 3117 4528 3133
rect 4586 3133 4706 3171
rect 4586 3117 4620 3133
rect 4494 3099 4510 3117
rect 4426 3083 4510 3099
rect 4604 3099 4620 3117
rect 4672 3117 4706 3133
rect 4764 3133 4884 3171
rect 4764 3117 4798 3133
rect 4672 3099 4688 3117
rect 4604 3083 4688 3099
rect 4782 3099 4798 3117
rect 4850 3117 4884 3133
rect 4942 3133 5062 3171
rect 4942 3117 4976 3133
rect 4850 3099 4866 3117
rect 4782 3083 4866 3099
rect 4960 3099 4976 3117
rect 5028 3117 5062 3133
rect 5120 3133 5240 3171
rect 5120 3117 5154 3133
rect 5028 3099 5044 3117
rect 4960 3083 5044 3099
rect 5138 3099 5154 3117
rect 5206 3117 5240 3133
rect 5298 3133 5418 3171
rect 5298 3117 5332 3133
rect 5206 3099 5222 3117
rect 5138 3083 5222 3099
rect 5316 3099 5332 3117
rect 5384 3117 5418 3133
rect 5476 3133 5596 3171
rect 5476 3117 5510 3133
rect 5384 3099 5400 3117
rect 5316 3083 5400 3099
rect 5494 3099 5510 3117
rect 5562 3117 5596 3133
rect 5654 3133 5774 3171
rect 5654 3117 5688 3133
rect 5562 3099 5578 3117
rect 5494 3083 5578 3099
rect 5672 3099 5688 3117
rect 5740 3117 5774 3133
rect 5832 3133 5952 3171
rect 5832 3117 5866 3133
rect 5740 3099 5756 3117
rect 5672 3083 5756 3099
rect 5850 3099 5866 3117
rect 5918 3117 5952 3133
rect 6010 3133 6130 3171
rect 6010 3117 6044 3133
rect 5918 3099 5934 3117
rect 5850 3083 5934 3099
rect 6028 3099 6044 3117
rect 6096 3117 6130 3133
rect 6188 3133 6308 3171
rect 6188 3117 6222 3133
rect 6096 3099 6112 3117
rect 6028 3083 6112 3099
rect 6206 3099 6222 3117
rect 6274 3117 6308 3133
rect 6366 3133 6486 3171
rect 6366 3117 6400 3133
rect 6274 3099 6290 3117
rect 6206 3083 6290 3099
rect 6384 3099 6400 3117
rect 6452 3117 6486 3133
rect 6544 3133 6664 3171
rect 6544 3117 6578 3133
rect 6452 3099 6468 3117
rect 6384 3083 6468 3099
rect 6562 3099 6578 3117
rect 6630 3117 6664 3133
rect 6722 3133 6842 3171
rect 6722 3117 6756 3133
rect 6630 3099 6646 3117
rect 6562 3083 6646 3099
rect 6740 3099 6756 3117
rect 6808 3117 6842 3133
rect 6900 3133 7020 3171
rect 7603 3151 7723 3189
rect 7781 3189 7815 3206
rect 7867 3206 7883 3223
rect 7977 3223 8061 3239
rect 7977 3206 7993 3223
rect 7867 3189 7901 3206
rect 7781 3151 7901 3189
rect 7959 3189 7993 3206
rect 8045 3206 8061 3223
rect 8155 3223 8239 3239
rect 8155 3206 8171 3223
rect 8045 3189 8079 3206
rect 7959 3151 8079 3189
rect 8137 3189 8171 3206
rect 8223 3206 8239 3223
rect 8333 3223 8417 3239
rect 8333 3206 8349 3223
rect 8223 3189 8257 3206
rect 8137 3151 8257 3189
rect 8315 3189 8349 3206
rect 8401 3206 8417 3223
rect 8511 3223 8595 3239
rect 8511 3206 8527 3223
rect 8401 3189 8435 3206
rect 8315 3151 8435 3189
rect 8493 3189 8527 3206
rect 8579 3206 8595 3223
rect 8689 3223 8773 3239
rect 8689 3206 8705 3223
rect 8579 3189 8613 3206
rect 8493 3151 8613 3189
rect 8671 3189 8705 3206
rect 8757 3206 8773 3223
rect 8867 3223 8951 3239
rect 8867 3206 8883 3223
rect 8757 3189 8791 3206
rect 8671 3151 8791 3189
rect 8849 3189 8883 3206
rect 8935 3206 8951 3223
rect 9045 3223 9129 3239
rect 9045 3206 9061 3223
rect 8935 3189 8969 3206
rect 8849 3151 8969 3189
rect 9027 3189 9061 3206
rect 9113 3206 9129 3223
rect 9223 3223 9307 3239
rect 9223 3206 9239 3223
rect 9113 3189 9147 3206
rect 9027 3151 9147 3189
rect 9205 3189 9239 3206
rect 9291 3206 9307 3223
rect 9401 3223 9485 3239
rect 9401 3206 9417 3223
rect 9291 3189 9325 3206
rect 9205 3151 9325 3189
rect 9383 3189 9417 3206
rect 9469 3206 9485 3223
rect 9579 3223 9663 3239
rect 9579 3206 9595 3223
rect 9469 3189 9503 3206
rect 9383 3151 9503 3189
rect 9561 3189 9595 3206
rect 9647 3206 9663 3223
rect 9757 3223 9841 3239
rect 9757 3206 9773 3223
rect 9647 3189 9681 3206
rect 9561 3151 9681 3189
rect 9739 3189 9773 3206
rect 9825 3206 9841 3223
rect 9935 3223 10019 3239
rect 9935 3206 9951 3223
rect 9825 3189 9859 3206
rect 9739 3151 9859 3189
rect 9917 3189 9951 3206
rect 10003 3206 10019 3223
rect 10308 3223 10392 3239
rect 10308 3206 10324 3223
rect 10003 3189 10037 3206
rect 9917 3151 10037 3189
rect 10290 3189 10324 3206
rect 10376 3206 10392 3223
rect 10486 3223 10570 3239
rect 10486 3206 10502 3223
rect 10376 3189 10410 3206
rect 10290 3151 10410 3189
rect 10468 3189 10502 3206
rect 10554 3206 10570 3223
rect 10664 3223 10748 3239
rect 10664 3206 10680 3223
rect 10554 3189 10588 3206
rect 10468 3151 10588 3189
rect 10646 3189 10680 3206
rect 10732 3206 10748 3223
rect 10842 3223 10926 3239
rect 10842 3206 10858 3223
rect 10732 3189 10766 3206
rect 10646 3151 10766 3189
rect 10824 3189 10858 3206
rect 10910 3206 10926 3223
rect 11020 3223 11104 3239
rect 11020 3206 11036 3223
rect 10910 3189 10944 3206
rect 10824 3151 10944 3189
rect 11002 3189 11036 3206
rect 11088 3206 11104 3223
rect 11198 3223 11282 3239
rect 11198 3206 11214 3223
rect 11088 3189 11122 3206
rect 11002 3151 11122 3189
rect 11180 3189 11214 3206
rect 11266 3206 11282 3223
rect 11376 3223 11460 3239
rect 11376 3206 11392 3223
rect 11266 3189 11300 3206
rect 11180 3151 11300 3189
rect 11358 3189 11392 3206
rect 11444 3206 11460 3223
rect 11554 3223 11638 3239
rect 11554 3206 11570 3223
rect 11444 3189 11478 3206
rect 11358 3151 11478 3189
rect 11536 3189 11570 3206
rect 11622 3206 11638 3223
rect 11732 3223 11816 3239
rect 11732 3206 11748 3223
rect 11622 3189 11656 3206
rect 11536 3151 11656 3189
rect 11714 3189 11748 3206
rect 11800 3206 11816 3223
rect 11910 3223 11994 3239
rect 11910 3206 11926 3223
rect 11800 3189 11834 3206
rect 11714 3151 11834 3189
rect 11892 3189 11926 3206
rect 11978 3206 11994 3223
rect 12088 3223 12172 3239
rect 12088 3206 12104 3223
rect 11978 3189 12012 3206
rect 11892 3151 12012 3189
rect 12070 3189 12104 3206
rect 12156 3206 12172 3223
rect 12266 3223 12350 3239
rect 12266 3206 12282 3223
rect 12156 3189 12190 3206
rect 12070 3151 12190 3189
rect 12248 3189 12282 3206
rect 12334 3206 12350 3223
rect 12444 3223 12528 3239
rect 12444 3206 12460 3223
rect 12334 3189 12368 3206
rect 12248 3151 12368 3189
rect 12426 3189 12460 3206
rect 12512 3206 12528 3223
rect 12622 3223 12706 3239
rect 12622 3206 12638 3223
rect 12512 3189 12546 3206
rect 12426 3151 12546 3189
rect 12604 3189 12638 3206
rect 12690 3206 12706 3223
rect 12690 3189 12724 3206
rect 12604 3151 12724 3189
rect 6900 3117 6934 3133
rect 6808 3099 6824 3117
rect 6740 3083 6824 3099
rect 6918 3099 6934 3117
rect 6986 3117 7020 3133
rect 6986 3099 7002 3117
rect 6918 3083 7002 3099
rect 492 3023 576 3039
rect 492 3005 508 3023
rect 474 2989 508 3005
rect 560 3005 576 3023
rect 670 3023 754 3039
rect 670 3005 686 3023
rect 560 2989 594 3005
rect 474 2951 594 2989
rect 652 2989 686 3005
rect 738 3005 754 3023
rect 848 3023 932 3039
rect 848 3005 864 3023
rect 738 2989 772 3005
rect 652 2951 772 2989
rect 830 2989 864 3005
rect 916 3005 932 3023
rect 1026 3023 1110 3039
rect 1026 3005 1042 3023
rect 916 2989 950 3005
rect 830 2951 950 2989
rect 1008 2989 1042 3005
rect 1094 3005 1110 3023
rect 1204 3023 1288 3039
rect 1204 3005 1220 3023
rect 1094 2989 1128 3005
rect 1008 2951 1128 2989
rect 1186 2989 1220 3005
rect 1272 3005 1288 3023
rect 1382 3023 1466 3039
rect 1382 3005 1398 3023
rect 1272 2989 1306 3005
rect 1186 2951 1306 2989
rect 1364 2989 1398 3005
rect 1450 3005 1466 3023
rect 1560 3023 1644 3039
rect 1560 3005 1576 3023
rect 1450 2989 1484 3005
rect 1364 2951 1484 2989
rect 1542 2989 1576 3005
rect 1628 3005 1644 3023
rect 1738 3023 1822 3039
rect 1738 3005 1754 3023
rect 1628 2989 1662 3005
rect 1542 2951 1662 2989
rect 1720 2989 1754 3005
rect 1806 3005 1822 3023
rect 1916 3023 2000 3039
rect 1916 3005 1932 3023
rect 1806 2989 1840 3005
rect 1720 2951 1840 2989
rect 1898 2989 1932 3005
rect 1984 3005 2000 3023
rect 2094 3023 2178 3039
rect 2094 3005 2110 3023
rect 1984 2989 2018 3005
rect 1898 2951 2018 2989
rect 2076 2989 2110 3005
rect 2162 3005 2178 3023
rect 2272 3023 2356 3039
rect 2272 3005 2288 3023
rect 2162 2989 2196 3005
rect 2076 2951 2196 2989
rect 2254 2989 2288 3005
rect 2340 3005 2356 3023
rect 2450 3023 2534 3039
rect 2450 3005 2466 3023
rect 2340 2989 2374 3005
rect 2254 2951 2374 2989
rect 2432 2989 2466 3005
rect 2518 3005 2534 3023
rect 2628 3023 2712 3039
rect 2628 3005 2644 3023
rect 2518 2989 2552 3005
rect 2432 2951 2552 2989
rect 2610 2989 2644 3005
rect 2696 3005 2712 3023
rect 2806 3023 2890 3039
rect 2806 3005 2822 3023
rect 2696 2989 2730 3005
rect 2610 2951 2730 2989
rect 2788 2989 2822 3005
rect 2874 3005 2890 3023
rect 2984 3023 3068 3039
rect 2984 3005 3000 3023
rect 2874 2989 2908 3005
rect 2788 2951 2908 2989
rect 2966 2989 3000 3005
rect 3052 3005 3068 3023
rect 3162 3023 3246 3039
rect 3162 3005 3178 3023
rect 3052 2989 3086 3005
rect 2966 2951 3086 2989
rect 3144 2989 3178 3005
rect 3230 3005 3246 3023
rect 3340 3023 3424 3039
rect 3340 3005 3356 3023
rect 3230 2989 3264 3005
rect 3144 2951 3264 2989
rect 3322 2989 3356 3005
rect 3408 3005 3424 3023
rect 3518 3023 3602 3039
rect 3518 3005 3534 3023
rect 3408 2989 3442 3005
rect 3322 2951 3442 2989
rect 3500 2989 3534 3005
rect 3586 3005 3602 3023
rect 3892 3023 3976 3039
rect 3892 3005 3908 3023
rect 3586 2989 3620 3005
rect 3500 2951 3620 2989
rect 3874 2989 3908 3005
rect 3960 3005 3976 3023
rect 4070 3023 4154 3039
rect 4070 3005 4086 3023
rect 3960 2989 3994 3005
rect 3874 2951 3994 2989
rect 4052 2989 4086 3005
rect 4138 3005 4154 3023
rect 4248 3023 4332 3039
rect 4248 3005 4264 3023
rect 4138 2989 4172 3005
rect 4052 2951 4172 2989
rect 4230 2989 4264 3005
rect 4316 3005 4332 3023
rect 4426 3023 4510 3039
rect 4426 3005 4442 3023
rect 4316 2989 4350 3005
rect 4230 2951 4350 2989
rect 4408 2989 4442 3005
rect 4494 3005 4510 3023
rect 4604 3023 4688 3039
rect 4604 3005 4620 3023
rect 4494 2989 4528 3005
rect 4408 2951 4528 2989
rect 4586 2989 4620 3005
rect 4672 3005 4688 3023
rect 4782 3023 4866 3039
rect 4782 3005 4798 3023
rect 4672 2989 4706 3005
rect 4586 2951 4706 2989
rect 4764 2989 4798 3005
rect 4850 3005 4866 3023
rect 4960 3023 5044 3039
rect 4960 3005 4976 3023
rect 4850 2989 4884 3005
rect 4764 2951 4884 2989
rect 4942 2989 4976 3005
rect 5028 3005 5044 3023
rect 5138 3023 5222 3039
rect 5138 3005 5154 3023
rect 5028 2989 5062 3005
rect 4942 2951 5062 2989
rect 5120 2989 5154 3005
rect 5206 3005 5222 3023
rect 5316 3023 5400 3039
rect 5316 3005 5332 3023
rect 5206 2989 5240 3005
rect 5120 2951 5240 2989
rect 5298 2989 5332 3005
rect 5384 3005 5400 3023
rect 5494 3023 5578 3039
rect 5494 3005 5510 3023
rect 5384 2989 5418 3005
rect 5298 2951 5418 2989
rect 5476 2989 5510 3005
rect 5562 3005 5578 3023
rect 5672 3023 5756 3039
rect 5672 3005 5688 3023
rect 5562 2989 5596 3005
rect 5476 2951 5596 2989
rect 5654 2989 5688 3005
rect 5740 3005 5756 3023
rect 5850 3023 5934 3039
rect 5850 3005 5866 3023
rect 5740 2989 5774 3005
rect 5654 2951 5774 2989
rect 5832 2989 5866 3005
rect 5918 3005 5934 3023
rect 6028 3023 6112 3039
rect 6028 3005 6044 3023
rect 5918 2989 5952 3005
rect 5832 2951 5952 2989
rect 6010 2989 6044 3005
rect 6096 3005 6112 3023
rect 6206 3023 6290 3039
rect 6206 3005 6222 3023
rect 6096 2989 6130 3005
rect 6010 2951 6130 2989
rect 6188 2989 6222 3005
rect 6274 3005 6290 3023
rect 6384 3023 6468 3039
rect 6384 3005 6400 3023
rect 6274 2989 6308 3005
rect 6188 2951 6308 2989
rect 6366 2989 6400 3005
rect 6452 3005 6468 3023
rect 6562 3023 6646 3039
rect 6562 3005 6578 3023
rect 6452 2989 6486 3005
rect 6366 2951 6486 2989
rect 6544 2989 6578 3005
rect 6630 3005 6646 3023
rect 6740 3023 6824 3039
rect 6740 3005 6756 3023
rect 6630 2989 6664 3005
rect 6544 2951 6664 2989
rect 6722 2989 6756 3005
rect 6808 3005 6824 3023
rect 6918 3023 7002 3039
rect 6918 3005 6934 3023
rect 6808 2989 6842 3005
rect 6722 2951 6842 2989
rect 6900 2989 6934 3005
rect 6986 3005 7002 3023
rect 6986 2989 7020 3005
rect 6900 2951 7020 2989
rect 7603 2833 7723 2871
rect 7603 2816 7637 2833
rect 7621 2799 7637 2816
rect 7689 2816 7723 2833
rect 7781 2833 7901 2871
rect 7781 2816 7815 2833
rect 7689 2799 7705 2816
rect 7621 2783 7705 2799
rect 7799 2799 7815 2816
rect 7867 2816 7901 2833
rect 7959 2833 8079 2871
rect 7959 2816 7993 2833
rect 7867 2799 7883 2816
rect 7799 2783 7883 2799
rect 7977 2799 7993 2816
rect 8045 2816 8079 2833
rect 8137 2833 8257 2871
rect 8137 2816 8171 2833
rect 8045 2799 8061 2816
rect 7977 2783 8061 2799
rect 8155 2799 8171 2816
rect 8223 2816 8257 2833
rect 8315 2833 8435 2871
rect 8315 2816 8349 2833
rect 8223 2799 8239 2816
rect 8155 2783 8239 2799
rect 8333 2799 8349 2816
rect 8401 2816 8435 2833
rect 8493 2833 8613 2871
rect 8493 2816 8527 2833
rect 8401 2799 8417 2816
rect 8333 2783 8417 2799
rect 8511 2799 8527 2816
rect 8579 2816 8613 2833
rect 8671 2833 8791 2871
rect 8671 2816 8705 2833
rect 8579 2799 8595 2816
rect 8511 2783 8595 2799
rect 8689 2799 8705 2816
rect 8757 2816 8791 2833
rect 8849 2833 8969 2871
rect 8849 2816 8883 2833
rect 8757 2799 8773 2816
rect 8689 2783 8773 2799
rect 8867 2799 8883 2816
rect 8935 2816 8969 2833
rect 9027 2833 9147 2871
rect 9027 2816 9061 2833
rect 8935 2799 8951 2816
rect 8867 2783 8951 2799
rect 9045 2799 9061 2816
rect 9113 2816 9147 2833
rect 9205 2833 9325 2871
rect 9205 2816 9239 2833
rect 9113 2799 9129 2816
rect 9045 2783 9129 2799
rect 9223 2799 9239 2816
rect 9291 2816 9325 2833
rect 9383 2833 9503 2871
rect 9383 2816 9417 2833
rect 9291 2799 9307 2816
rect 9223 2783 9307 2799
rect 9401 2799 9417 2816
rect 9469 2816 9503 2833
rect 9561 2833 9681 2871
rect 9561 2816 9595 2833
rect 9469 2799 9485 2816
rect 9401 2783 9485 2799
rect 9579 2799 9595 2816
rect 9647 2816 9681 2833
rect 9739 2833 9859 2871
rect 9739 2816 9773 2833
rect 9647 2799 9663 2816
rect 9579 2783 9663 2799
rect 9757 2799 9773 2816
rect 9825 2816 9859 2833
rect 9917 2833 10037 2871
rect 9917 2816 9951 2833
rect 9825 2799 9841 2816
rect 9757 2783 9841 2799
rect 9935 2799 9951 2816
rect 10003 2816 10037 2833
rect 10290 2833 10410 2871
rect 10290 2816 10324 2833
rect 10003 2799 10019 2816
rect 9935 2783 10019 2799
rect 10308 2799 10324 2816
rect 10376 2816 10410 2833
rect 10468 2833 10588 2871
rect 10468 2816 10502 2833
rect 10376 2799 10392 2816
rect 10308 2783 10392 2799
rect 10486 2799 10502 2816
rect 10554 2816 10588 2833
rect 10646 2833 10766 2871
rect 10646 2816 10680 2833
rect 10554 2799 10570 2816
rect 10486 2783 10570 2799
rect 10664 2799 10680 2816
rect 10732 2816 10766 2833
rect 10824 2833 10944 2871
rect 10824 2816 10858 2833
rect 10732 2799 10748 2816
rect 10664 2783 10748 2799
rect 10842 2799 10858 2816
rect 10910 2816 10944 2833
rect 11002 2833 11122 2871
rect 11002 2816 11036 2833
rect 10910 2799 10926 2816
rect 10842 2783 10926 2799
rect 11020 2799 11036 2816
rect 11088 2816 11122 2833
rect 11180 2833 11300 2871
rect 11180 2816 11214 2833
rect 11088 2799 11104 2816
rect 11020 2783 11104 2799
rect 11198 2799 11214 2816
rect 11266 2816 11300 2833
rect 11358 2833 11478 2871
rect 11358 2816 11392 2833
rect 11266 2799 11282 2816
rect 11198 2783 11282 2799
rect 11376 2799 11392 2816
rect 11444 2816 11478 2833
rect 11536 2833 11656 2871
rect 11536 2816 11570 2833
rect 11444 2799 11460 2816
rect 11376 2783 11460 2799
rect 11554 2799 11570 2816
rect 11622 2816 11656 2833
rect 11714 2833 11834 2871
rect 11714 2816 11748 2833
rect 11622 2799 11638 2816
rect 11554 2783 11638 2799
rect 11732 2799 11748 2816
rect 11800 2816 11834 2833
rect 11892 2833 12012 2871
rect 11892 2816 11926 2833
rect 11800 2799 11816 2816
rect 11732 2783 11816 2799
rect 11910 2799 11926 2816
rect 11978 2816 12012 2833
rect 12070 2833 12190 2871
rect 12070 2816 12104 2833
rect 11978 2799 11994 2816
rect 11910 2783 11994 2799
rect 12088 2799 12104 2816
rect 12156 2816 12190 2833
rect 12248 2833 12368 2871
rect 12248 2816 12282 2833
rect 12156 2799 12172 2816
rect 12088 2783 12172 2799
rect 12266 2799 12282 2816
rect 12334 2816 12368 2833
rect 12426 2833 12546 2871
rect 12426 2816 12460 2833
rect 12334 2799 12350 2816
rect 12266 2783 12350 2799
rect 12444 2799 12460 2816
rect 12512 2816 12546 2833
rect 12604 2833 12724 2871
rect 12604 2816 12638 2833
rect 12512 2799 12528 2816
rect 12444 2783 12528 2799
rect 12622 2799 12638 2816
rect 12690 2816 12724 2833
rect 12690 2799 12706 2816
rect 12622 2783 12706 2799
rect 7621 2723 7705 2739
rect 7621 2706 7637 2723
rect 7603 2689 7637 2706
rect 7689 2706 7705 2723
rect 7799 2723 7883 2739
rect 7799 2706 7815 2723
rect 7689 2689 7723 2706
rect 474 2633 594 2671
rect 474 2617 508 2633
rect 492 2599 508 2617
rect 560 2617 594 2633
rect 652 2633 772 2671
rect 652 2617 686 2633
rect 560 2599 576 2617
rect 492 2583 576 2599
rect 670 2599 686 2617
rect 738 2617 772 2633
rect 830 2633 950 2671
rect 830 2617 864 2633
rect 738 2599 754 2617
rect 670 2583 754 2599
rect 848 2599 864 2617
rect 916 2617 950 2633
rect 1008 2633 1128 2671
rect 1008 2617 1042 2633
rect 916 2599 932 2617
rect 848 2583 932 2599
rect 1026 2599 1042 2617
rect 1094 2617 1128 2633
rect 1186 2633 1306 2671
rect 1186 2617 1220 2633
rect 1094 2599 1110 2617
rect 1026 2583 1110 2599
rect 1204 2599 1220 2617
rect 1272 2617 1306 2633
rect 1364 2633 1484 2671
rect 1364 2617 1398 2633
rect 1272 2599 1288 2617
rect 1204 2583 1288 2599
rect 1382 2599 1398 2617
rect 1450 2617 1484 2633
rect 1542 2633 1662 2671
rect 1542 2617 1576 2633
rect 1450 2599 1466 2617
rect 1382 2583 1466 2599
rect 1560 2599 1576 2617
rect 1628 2617 1662 2633
rect 1720 2633 1840 2671
rect 1720 2617 1754 2633
rect 1628 2599 1644 2617
rect 1560 2583 1644 2599
rect 1738 2599 1754 2617
rect 1806 2617 1840 2633
rect 1898 2633 2018 2671
rect 1898 2617 1932 2633
rect 1806 2599 1822 2617
rect 1738 2583 1822 2599
rect 1916 2599 1932 2617
rect 1984 2617 2018 2633
rect 2076 2633 2196 2671
rect 2076 2617 2110 2633
rect 1984 2599 2000 2617
rect 1916 2583 2000 2599
rect 2094 2599 2110 2617
rect 2162 2617 2196 2633
rect 2254 2633 2374 2671
rect 2254 2617 2288 2633
rect 2162 2599 2178 2617
rect 2094 2583 2178 2599
rect 2272 2599 2288 2617
rect 2340 2617 2374 2633
rect 2432 2633 2552 2671
rect 2432 2617 2466 2633
rect 2340 2599 2356 2617
rect 2272 2583 2356 2599
rect 2450 2599 2466 2617
rect 2518 2617 2552 2633
rect 2610 2633 2730 2671
rect 2610 2617 2644 2633
rect 2518 2599 2534 2617
rect 2450 2583 2534 2599
rect 2628 2599 2644 2617
rect 2696 2617 2730 2633
rect 2788 2633 2908 2671
rect 2788 2617 2822 2633
rect 2696 2599 2712 2617
rect 2628 2583 2712 2599
rect 2806 2599 2822 2617
rect 2874 2617 2908 2633
rect 2966 2633 3086 2671
rect 2966 2617 3000 2633
rect 2874 2599 2890 2617
rect 2806 2583 2890 2599
rect 2984 2599 3000 2617
rect 3052 2617 3086 2633
rect 3144 2633 3264 2671
rect 3144 2617 3178 2633
rect 3052 2599 3068 2617
rect 2984 2583 3068 2599
rect 3162 2599 3178 2617
rect 3230 2617 3264 2633
rect 3322 2633 3442 2671
rect 3322 2617 3356 2633
rect 3230 2599 3246 2617
rect 3162 2583 3246 2599
rect 3340 2599 3356 2617
rect 3408 2617 3442 2633
rect 3500 2633 3620 2671
rect 3500 2617 3534 2633
rect 3408 2599 3424 2617
rect 3340 2583 3424 2599
rect 3518 2599 3534 2617
rect 3586 2617 3620 2633
rect 3874 2633 3994 2671
rect 3874 2617 3908 2633
rect 3586 2599 3602 2617
rect 3518 2583 3602 2599
rect 3892 2599 3908 2617
rect 3960 2617 3994 2633
rect 4052 2633 4172 2671
rect 4052 2617 4086 2633
rect 3960 2599 3976 2617
rect 3892 2583 3976 2599
rect 4070 2599 4086 2617
rect 4138 2617 4172 2633
rect 4230 2633 4350 2671
rect 4230 2617 4264 2633
rect 4138 2599 4154 2617
rect 4070 2583 4154 2599
rect 4248 2599 4264 2617
rect 4316 2617 4350 2633
rect 4408 2633 4528 2671
rect 4408 2617 4442 2633
rect 4316 2599 4332 2617
rect 4248 2583 4332 2599
rect 4426 2599 4442 2617
rect 4494 2617 4528 2633
rect 4586 2633 4706 2671
rect 4586 2617 4620 2633
rect 4494 2599 4510 2617
rect 4426 2583 4510 2599
rect 4604 2599 4620 2617
rect 4672 2617 4706 2633
rect 4764 2633 4884 2671
rect 4764 2617 4798 2633
rect 4672 2599 4688 2617
rect 4604 2583 4688 2599
rect 4782 2599 4798 2617
rect 4850 2617 4884 2633
rect 4942 2633 5062 2671
rect 4942 2617 4976 2633
rect 4850 2599 4866 2617
rect 4782 2583 4866 2599
rect 4960 2599 4976 2617
rect 5028 2617 5062 2633
rect 5120 2633 5240 2671
rect 5120 2617 5154 2633
rect 5028 2599 5044 2617
rect 4960 2583 5044 2599
rect 5138 2599 5154 2617
rect 5206 2617 5240 2633
rect 5298 2633 5418 2671
rect 5298 2617 5332 2633
rect 5206 2599 5222 2617
rect 5138 2583 5222 2599
rect 5316 2599 5332 2617
rect 5384 2617 5418 2633
rect 5476 2633 5596 2671
rect 5476 2617 5510 2633
rect 5384 2599 5400 2617
rect 5316 2583 5400 2599
rect 5494 2599 5510 2617
rect 5562 2617 5596 2633
rect 5654 2633 5774 2671
rect 5654 2617 5688 2633
rect 5562 2599 5578 2617
rect 5494 2583 5578 2599
rect 5672 2599 5688 2617
rect 5740 2617 5774 2633
rect 5832 2633 5952 2671
rect 5832 2617 5866 2633
rect 5740 2599 5756 2617
rect 5672 2583 5756 2599
rect 5850 2599 5866 2617
rect 5918 2617 5952 2633
rect 6010 2633 6130 2671
rect 6010 2617 6044 2633
rect 5918 2599 5934 2617
rect 5850 2583 5934 2599
rect 6028 2599 6044 2617
rect 6096 2617 6130 2633
rect 6188 2633 6308 2671
rect 6188 2617 6222 2633
rect 6096 2599 6112 2617
rect 6028 2583 6112 2599
rect 6206 2599 6222 2617
rect 6274 2617 6308 2633
rect 6366 2633 6486 2671
rect 6366 2617 6400 2633
rect 6274 2599 6290 2617
rect 6206 2583 6290 2599
rect 6384 2599 6400 2617
rect 6452 2617 6486 2633
rect 6544 2633 6664 2671
rect 6544 2617 6578 2633
rect 6452 2599 6468 2617
rect 6384 2583 6468 2599
rect 6562 2599 6578 2617
rect 6630 2617 6664 2633
rect 6722 2633 6842 2671
rect 6722 2617 6756 2633
rect 6630 2599 6646 2617
rect 6562 2583 6646 2599
rect 6740 2599 6756 2617
rect 6808 2617 6842 2633
rect 6900 2633 7020 2671
rect 7603 2651 7723 2689
rect 7781 2689 7815 2706
rect 7867 2706 7883 2723
rect 7977 2723 8061 2739
rect 7977 2706 7993 2723
rect 7867 2689 7901 2706
rect 7781 2651 7901 2689
rect 7959 2689 7993 2706
rect 8045 2706 8061 2723
rect 8155 2723 8239 2739
rect 8155 2706 8171 2723
rect 8045 2689 8079 2706
rect 7959 2651 8079 2689
rect 8137 2689 8171 2706
rect 8223 2706 8239 2723
rect 8333 2723 8417 2739
rect 8333 2706 8349 2723
rect 8223 2689 8257 2706
rect 8137 2651 8257 2689
rect 8315 2689 8349 2706
rect 8401 2706 8417 2723
rect 8511 2723 8595 2739
rect 8511 2706 8527 2723
rect 8401 2689 8435 2706
rect 8315 2651 8435 2689
rect 8493 2689 8527 2706
rect 8579 2706 8595 2723
rect 8689 2723 8773 2739
rect 8689 2706 8705 2723
rect 8579 2689 8613 2706
rect 8493 2651 8613 2689
rect 8671 2689 8705 2706
rect 8757 2706 8773 2723
rect 8867 2723 8951 2739
rect 8867 2706 8883 2723
rect 8757 2689 8791 2706
rect 8671 2651 8791 2689
rect 8849 2689 8883 2706
rect 8935 2706 8951 2723
rect 9045 2723 9129 2739
rect 9045 2706 9061 2723
rect 8935 2689 8969 2706
rect 8849 2651 8969 2689
rect 9027 2689 9061 2706
rect 9113 2706 9129 2723
rect 9223 2723 9307 2739
rect 9223 2706 9239 2723
rect 9113 2689 9147 2706
rect 9027 2651 9147 2689
rect 9205 2689 9239 2706
rect 9291 2706 9307 2723
rect 9401 2723 9485 2739
rect 9401 2706 9417 2723
rect 9291 2689 9325 2706
rect 9205 2651 9325 2689
rect 9383 2689 9417 2706
rect 9469 2706 9485 2723
rect 9579 2723 9663 2739
rect 9579 2706 9595 2723
rect 9469 2689 9503 2706
rect 9383 2651 9503 2689
rect 9561 2689 9595 2706
rect 9647 2706 9663 2723
rect 9757 2723 9841 2739
rect 9757 2706 9773 2723
rect 9647 2689 9681 2706
rect 9561 2651 9681 2689
rect 9739 2689 9773 2706
rect 9825 2706 9841 2723
rect 9935 2723 10019 2739
rect 9935 2706 9951 2723
rect 9825 2689 9859 2706
rect 9739 2651 9859 2689
rect 9917 2689 9951 2706
rect 10003 2706 10019 2723
rect 10308 2723 10392 2739
rect 10308 2706 10324 2723
rect 10003 2689 10037 2706
rect 9917 2651 10037 2689
rect 10290 2689 10324 2706
rect 10376 2706 10392 2723
rect 10486 2723 10570 2739
rect 10486 2706 10502 2723
rect 10376 2689 10410 2706
rect 10290 2651 10410 2689
rect 10468 2689 10502 2706
rect 10554 2706 10570 2723
rect 10664 2723 10748 2739
rect 10664 2706 10680 2723
rect 10554 2689 10588 2706
rect 10468 2651 10588 2689
rect 10646 2689 10680 2706
rect 10732 2706 10748 2723
rect 10842 2723 10926 2739
rect 10842 2706 10858 2723
rect 10732 2689 10766 2706
rect 10646 2651 10766 2689
rect 10824 2689 10858 2706
rect 10910 2706 10926 2723
rect 11020 2723 11104 2739
rect 11020 2706 11036 2723
rect 10910 2689 10944 2706
rect 10824 2651 10944 2689
rect 11002 2689 11036 2706
rect 11088 2706 11104 2723
rect 11198 2723 11282 2739
rect 11198 2706 11214 2723
rect 11088 2689 11122 2706
rect 11002 2651 11122 2689
rect 11180 2689 11214 2706
rect 11266 2706 11282 2723
rect 11376 2723 11460 2739
rect 11376 2706 11392 2723
rect 11266 2689 11300 2706
rect 11180 2651 11300 2689
rect 11358 2689 11392 2706
rect 11444 2706 11460 2723
rect 11554 2723 11638 2739
rect 11554 2706 11570 2723
rect 11444 2689 11478 2706
rect 11358 2651 11478 2689
rect 11536 2689 11570 2706
rect 11622 2706 11638 2723
rect 11732 2723 11816 2739
rect 11732 2706 11748 2723
rect 11622 2689 11656 2706
rect 11536 2651 11656 2689
rect 11714 2689 11748 2706
rect 11800 2706 11816 2723
rect 11910 2723 11994 2739
rect 11910 2706 11926 2723
rect 11800 2689 11834 2706
rect 11714 2651 11834 2689
rect 11892 2689 11926 2706
rect 11978 2706 11994 2723
rect 12088 2723 12172 2739
rect 12088 2706 12104 2723
rect 11978 2689 12012 2706
rect 11892 2651 12012 2689
rect 12070 2689 12104 2706
rect 12156 2706 12172 2723
rect 12266 2723 12350 2739
rect 12266 2706 12282 2723
rect 12156 2689 12190 2706
rect 12070 2651 12190 2689
rect 12248 2689 12282 2706
rect 12334 2706 12350 2723
rect 12444 2723 12528 2739
rect 12444 2706 12460 2723
rect 12334 2689 12368 2706
rect 12248 2651 12368 2689
rect 12426 2689 12460 2706
rect 12512 2706 12528 2723
rect 12622 2723 12706 2739
rect 12622 2706 12638 2723
rect 12512 2689 12546 2706
rect 12426 2651 12546 2689
rect 12604 2689 12638 2706
rect 12690 2706 12706 2723
rect 12690 2689 12724 2706
rect 12604 2651 12724 2689
rect 6900 2617 6934 2633
rect 6808 2599 6824 2617
rect 6740 2583 6824 2599
rect 6918 2599 6934 2617
rect 6986 2617 7020 2633
rect 6986 2599 7002 2617
rect 6918 2583 7002 2599
rect 492 2523 576 2539
rect 492 2505 508 2523
rect 474 2489 508 2505
rect 560 2505 576 2523
rect 670 2523 754 2539
rect 670 2505 686 2523
rect 560 2489 594 2505
rect 474 2451 594 2489
rect 652 2489 686 2505
rect 738 2505 754 2523
rect 848 2523 932 2539
rect 848 2505 864 2523
rect 738 2489 772 2505
rect 652 2451 772 2489
rect 830 2489 864 2505
rect 916 2505 932 2523
rect 1026 2523 1110 2539
rect 1026 2505 1042 2523
rect 916 2489 950 2505
rect 830 2451 950 2489
rect 1008 2489 1042 2505
rect 1094 2505 1110 2523
rect 1204 2523 1288 2539
rect 1204 2505 1220 2523
rect 1094 2489 1128 2505
rect 1008 2451 1128 2489
rect 1186 2489 1220 2505
rect 1272 2505 1288 2523
rect 1382 2523 1466 2539
rect 1382 2505 1398 2523
rect 1272 2489 1306 2505
rect 1186 2451 1306 2489
rect 1364 2489 1398 2505
rect 1450 2505 1466 2523
rect 1560 2523 1644 2539
rect 1560 2505 1576 2523
rect 1450 2489 1484 2505
rect 1364 2451 1484 2489
rect 1542 2489 1576 2505
rect 1628 2505 1644 2523
rect 1738 2523 1822 2539
rect 1738 2505 1754 2523
rect 1628 2489 1662 2505
rect 1542 2451 1662 2489
rect 1720 2489 1754 2505
rect 1806 2505 1822 2523
rect 1916 2523 2000 2539
rect 1916 2505 1932 2523
rect 1806 2489 1840 2505
rect 1720 2451 1840 2489
rect 1898 2489 1932 2505
rect 1984 2505 2000 2523
rect 2094 2523 2178 2539
rect 2094 2505 2110 2523
rect 1984 2489 2018 2505
rect 1898 2451 2018 2489
rect 2076 2489 2110 2505
rect 2162 2505 2178 2523
rect 2272 2523 2356 2539
rect 2272 2505 2288 2523
rect 2162 2489 2196 2505
rect 2076 2451 2196 2489
rect 2254 2489 2288 2505
rect 2340 2505 2356 2523
rect 2450 2523 2534 2539
rect 2450 2505 2466 2523
rect 2340 2489 2374 2505
rect 2254 2451 2374 2489
rect 2432 2489 2466 2505
rect 2518 2505 2534 2523
rect 2628 2523 2712 2539
rect 2628 2505 2644 2523
rect 2518 2489 2552 2505
rect 2432 2451 2552 2489
rect 2610 2489 2644 2505
rect 2696 2505 2712 2523
rect 2806 2523 2890 2539
rect 2806 2505 2822 2523
rect 2696 2489 2730 2505
rect 2610 2451 2730 2489
rect 2788 2489 2822 2505
rect 2874 2505 2890 2523
rect 2984 2523 3068 2539
rect 2984 2505 3000 2523
rect 2874 2489 2908 2505
rect 2788 2451 2908 2489
rect 2966 2489 3000 2505
rect 3052 2505 3068 2523
rect 3162 2523 3246 2539
rect 3162 2505 3178 2523
rect 3052 2489 3086 2505
rect 2966 2451 3086 2489
rect 3144 2489 3178 2505
rect 3230 2505 3246 2523
rect 3340 2523 3424 2539
rect 3340 2505 3356 2523
rect 3230 2489 3264 2505
rect 3144 2451 3264 2489
rect 3322 2489 3356 2505
rect 3408 2505 3424 2523
rect 3518 2523 3602 2539
rect 3518 2505 3534 2523
rect 3408 2489 3442 2505
rect 3322 2451 3442 2489
rect 3500 2489 3534 2505
rect 3586 2505 3602 2523
rect 3892 2523 3976 2539
rect 3892 2505 3908 2523
rect 3586 2489 3620 2505
rect 3500 2451 3620 2489
rect 3874 2489 3908 2505
rect 3960 2505 3976 2523
rect 4070 2523 4154 2539
rect 4070 2505 4086 2523
rect 3960 2489 3994 2505
rect 3874 2451 3994 2489
rect 4052 2489 4086 2505
rect 4138 2505 4154 2523
rect 4248 2523 4332 2539
rect 4248 2505 4264 2523
rect 4138 2489 4172 2505
rect 4052 2451 4172 2489
rect 4230 2489 4264 2505
rect 4316 2505 4332 2523
rect 4426 2523 4510 2539
rect 4426 2505 4442 2523
rect 4316 2489 4350 2505
rect 4230 2451 4350 2489
rect 4408 2489 4442 2505
rect 4494 2505 4510 2523
rect 4604 2523 4688 2539
rect 4604 2505 4620 2523
rect 4494 2489 4528 2505
rect 4408 2451 4528 2489
rect 4586 2489 4620 2505
rect 4672 2505 4688 2523
rect 4782 2523 4866 2539
rect 4782 2505 4798 2523
rect 4672 2489 4706 2505
rect 4586 2451 4706 2489
rect 4764 2489 4798 2505
rect 4850 2505 4866 2523
rect 4960 2523 5044 2539
rect 4960 2505 4976 2523
rect 4850 2489 4884 2505
rect 4764 2451 4884 2489
rect 4942 2489 4976 2505
rect 5028 2505 5044 2523
rect 5138 2523 5222 2539
rect 5138 2505 5154 2523
rect 5028 2489 5062 2505
rect 4942 2451 5062 2489
rect 5120 2489 5154 2505
rect 5206 2505 5222 2523
rect 5316 2523 5400 2539
rect 5316 2505 5332 2523
rect 5206 2489 5240 2505
rect 5120 2451 5240 2489
rect 5298 2489 5332 2505
rect 5384 2505 5400 2523
rect 5494 2523 5578 2539
rect 5494 2505 5510 2523
rect 5384 2489 5418 2505
rect 5298 2451 5418 2489
rect 5476 2489 5510 2505
rect 5562 2505 5578 2523
rect 5672 2523 5756 2539
rect 5672 2505 5688 2523
rect 5562 2489 5596 2505
rect 5476 2451 5596 2489
rect 5654 2489 5688 2505
rect 5740 2505 5756 2523
rect 5850 2523 5934 2539
rect 5850 2505 5866 2523
rect 5740 2489 5774 2505
rect 5654 2451 5774 2489
rect 5832 2489 5866 2505
rect 5918 2505 5934 2523
rect 6028 2523 6112 2539
rect 6028 2505 6044 2523
rect 5918 2489 5952 2505
rect 5832 2451 5952 2489
rect 6010 2489 6044 2505
rect 6096 2505 6112 2523
rect 6206 2523 6290 2539
rect 6206 2505 6222 2523
rect 6096 2489 6130 2505
rect 6010 2451 6130 2489
rect 6188 2489 6222 2505
rect 6274 2505 6290 2523
rect 6384 2523 6468 2539
rect 6384 2505 6400 2523
rect 6274 2489 6308 2505
rect 6188 2451 6308 2489
rect 6366 2489 6400 2505
rect 6452 2505 6468 2523
rect 6562 2523 6646 2539
rect 6562 2505 6578 2523
rect 6452 2489 6486 2505
rect 6366 2451 6486 2489
rect 6544 2489 6578 2505
rect 6630 2505 6646 2523
rect 6740 2523 6824 2539
rect 6740 2505 6756 2523
rect 6630 2489 6664 2505
rect 6544 2451 6664 2489
rect 6722 2489 6756 2505
rect 6808 2505 6824 2523
rect 6918 2523 7002 2539
rect 6918 2505 6934 2523
rect 6808 2489 6842 2505
rect 6722 2451 6842 2489
rect 6900 2489 6934 2505
rect 6986 2505 7002 2523
rect 6986 2489 7020 2505
rect 6900 2451 7020 2489
rect 7603 2333 7723 2371
rect 7603 2316 7637 2333
rect 7621 2299 7637 2316
rect 7689 2316 7723 2333
rect 7781 2333 7901 2371
rect 7781 2316 7815 2333
rect 7689 2299 7705 2316
rect 7621 2283 7705 2299
rect 7799 2299 7815 2316
rect 7867 2316 7901 2333
rect 7959 2333 8079 2371
rect 7959 2316 7993 2333
rect 7867 2299 7883 2316
rect 7799 2283 7883 2299
rect 7977 2299 7993 2316
rect 8045 2316 8079 2333
rect 8137 2333 8257 2371
rect 8137 2316 8171 2333
rect 8045 2299 8061 2316
rect 7977 2283 8061 2299
rect 8155 2299 8171 2316
rect 8223 2316 8257 2333
rect 8315 2333 8435 2371
rect 8315 2316 8349 2333
rect 8223 2299 8239 2316
rect 8155 2283 8239 2299
rect 8333 2299 8349 2316
rect 8401 2316 8435 2333
rect 8493 2333 8613 2371
rect 8493 2316 8527 2333
rect 8401 2299 8417 2316
rect 8333 2283 8417 2299
rect 8511 2299 8527 2316
rect 8579 2316 8613 2333
rect 8671 2333 8791 2371
rect 8671 2316 8705 2333
rect 8579 2299 8595 2316
rect 8511 2283 8595 2299
rect 8689 2299 8705 2316
rect 8757 2316 8791 2333
rect 8849 2333 8969 2371
rect 8849 2316 8883 2333
rect 8757 2299 8773 2316
rect 8689 2283 8773 2299
rect 8867 2299 8883 2316
rect 8935 2316 8969 2333
rect 9027 2333 9147 2371
rect 9027 2316 9061 2333
rect 8935 2299 8951 2316
rect 8867 2283 8951 2299
rect 9045 2299 9061 2316
rect 9113 2316 9147 2333
rect 9205 2333 9325 2371
rect 9205 2316 9239 2333
rect 9113 2299 9129 2316
rect 9045 2283 9129 2299
rect 9223 2299 9239 2316
rect 9291 2316 9325 2333
rect 9383 2333 9503 2371
rect 9383 2316 9417 2333
rect 9291 2299 9307 2316
rect 9223 2283 9307 2299
rect 9401 2299 9417 2316
rect 9469 2316 9503 2333
rect 9561 2333 9681 2371
rect 9561 2316 9595 2333
rect 9469 2299 9485 2316
rect 9401 2283 9485 2299
rect 9579 2299 9595 2316
rect 9647 2316 9681 2333
rect 9739 2333 9859 2371
rect 9739 2316 9773 2333
rect 9647 2299 9663 2316
rect 9579 2283 9663 2299
rect 9757 2299 9773 2316
rect 9825 2316 9859 2333
rect 9917 2333 10037 2371
rect 9917 2316 9951 2333
rect 9825 2299 9841 2316
rect 9757 2283 9841 2299
rect 9935 2299 9951 2316
rect 10003 2316 10037 2333
rect 10290 2333 10410 2371
rect 10290 2316 10324 2333
rect 10003 2299 10019 2316
rect 9935 2283 10019 2299
rect 10308 2299 10324 2316
rect 10376 2316 10410 2333
rect 10468 2333 10588 2371
rect 10468 2316 10502 2333
rect 10376 2299 10392 2316
rect 10308 2283 10392 2299
rect 10486 2299 10502 2316
rect 10554 2316 10588 2333
rect 10646 2333 10766 2371
rect 10646 2316 10680 2333
rect 10554 2299 10570 2316
rect 10486 2283 10570 2299
rect 10664 2299 10680 2316
rect 10732 2316 10766 2333
rect 10824 2333 10944 2371
rect 10824 2316 10858 2333
rect 10732 2299 10748 2316
rect 10664 2283 10748 2299
rect 10842 2299 10858 2316
rect 10910 2316 10944 2333
rect 11002 2333 11122 2371
rect 11002 2316 11036 2333
rect 10910 2299 10926 2316
rect 10842 2283 10926 2299
rect 11020 2299 11036 2316
rect 11088 2316 11122 2333
rect 11180 2333 11300 2371
rect 11180 2316 11214 2333
rect 11088 2299 11104 2316
rect 11020 2283 11104 2299
rect 11198 2299 11214 2316
rect 11266 2316 11300 2333
rect 11358 2333 11478 2371
rect 11358 2316 11392 2333
rect 11266 2299 11282 2316
rect 11198 2283 11282 2299
rect 11376 2299 11392 2316
rect 11444 2316 11478 2333
rect 11536 2333 11656 2371
rect 11536 2316 11570 2333
rect 11444 2299 11460 2316
rect 11376 2283 11460 2299
rect 11554 2299 11570 2316
rect 11622 2316 11656 2333
rect 11714 2333 11834 2371
rect 11714 2316 11748 2333
rect 11622 2299 11638 2316
rect 11554 2283 11638 2299
rect 11732 2299 11748 2316
rect 11800 2316 11834 2333
rect 11892 2333 12012 2371
rect 11892 2316 11926 2333
rect 11800 2299 11816 2316
rect 11732 2283 11816 2299
rect 11910 2299 11926 2316
rect 11978 2316 12012 2333
rect 12070 2333 12190 2371
rect 12070 2316 12104 2333
rect 11978 2299 11994 2316
rect 11910 2283 11994 2299
rect 12088 2299 12104 2316
rect 12156 2316 12190 2333
rect 12248 2333 12368 2371
rect 12248 2316 12282 2333
rect 12156 2299 12172 2316
rect 12088 2283 12172 2299
rect 12266 2299 12282 2316
rect 12334 2316 12368 2333
rect 12426 2333 12546 2371
rect 12426 2316 12460 2333
rect 12334 2299 12350 2316
rect 12266 2283 12350 2299
rect 12444 2299 12460 2316
rect 12512 2316 12546 2333
rect 12604 2333 12724 2371
rect 12604 2316 12638 2333
rect 12512 2299 12528 2316
rect 12444 2283 12528 2299
rect 12622 2299 12638 2316
rect 12690 2316 12724 2333
rect 12690 2299 12706 2316
rect 12622 2283 12706 2299
rect 474 2133 594 2171
rect 474 2117 508 2133
rect 492 2099 508 2117
rect 560 2117 594 2133
rect 652 2133 772 2171
rect 652 2117 686 2133
rect 560 2099 576 2117
rect 492 2083 576 2099
rect 670 2099 686 2117
rect 738 2117 772 2133
rect 830 2133 950 2171
rect 830 2117 864 2133
rect 738 2099 754 2117
rect 670 2083 754 2099
rect 848 2099 864 2117
rect 916 2117 950 2133
rect 1008 2133 1128 2171
rect 1008 2117 1042 2133
rect 916 2099 932 2117
rect 848 2083 932 2099
rect 1026 2099 1042 2117
rect 1094 2117 1128 2133
rect 1186 2133 1306 2171
rect 1186 2117 1220 2133
rect 1094 2099 1110 2117
rect 1026 2083 1110 2099
rect 1204 2099 1220 2117
rect 1272 2117 1306 2133
rect 1364 2133 1484 2171
rect 1364 2117 1398 2133
rect 1272 2099 1288 2117
rect 1204 2083 1288 2099
rect 1382 2099 1398 2117
rect 1450 2117 1484 2133
rect 1542 2133 1662 2171
rect 1542 2117 1576 2133
rect 1450 2099 1466 2117
rect 1382 2083 1466 2099
rect 1560 2099 1576 2117
rect 1628 2117 1662 2133
rect 1720 2133 1840 2171
rect 1720 2117 1754 2133
rect 1628 2099 1644 2117
rect 1560 2083 1644 2099
rect 1738 2099 1754 2117
rect 1806 2117 1840 2133
rect 1898 2133 2018 2171
rect 1898 2117 1932 2133
rect 1806 2099 1822 2117
rect 1738 2083 1822 2099
rect 1916 2099 1932 2117
rect 1984 2117 2018 2133
rect 2076 2133 2196 2171
rect 2076 2117 2110 2133
rect 1984 2099 2000 2117
rect 1916 2083 2000 2099
rect 2094 2099 2110 2117
rect 2162 2117 2196 2133
rect 2254 2133 2374 2171
rect 2254 2117 2288 2133
rect 2162 2099 2178 2117
rect 2094 2083 2178 2099
rect 2272 2099 2288 2117
rect 2340 2117 2374 2133
rect 2432 2133 2552 2171
rect 2432 2117 2466 2133
rect 2340 2099 2356 2117
rect 2272 2083 2356 2099
rect 2450 2099 2466 2117
rect 2518 2117 2552 2133
rect 2610 2133 2730 2171
rect 2610 2117 2644 2133
rect 2518 2099 2534 2117
rect 2450 2083 2534 2099
rect 2628 2099 2644 2117
rect 2696 2117 2730 2133
rect 2788 2133 2908 2171
rect 2788 2117 2822 2133
rect 2696 2099 2712 2117
rect 2628 2083 2712 2099
rect 2806 2099 2822 2117
rect 2874 2117 2908 2133
rect 2966 2133 3086 2171
rect 2966 2117 3000 2133
rect 2874 2099 2890 2117
rect 2806 2083 2890 2099
rect 2984 2099 3000 2117
rect 3052 2117 3086 2133
rect 3144 2133 3264 2171
rect 3144 2117 3178 2133
rect 3052 2099 3068 2117
rect 2984 2083 3068 2099
rect 3162 2099 3178 2117
rect 3230 2117 3264 2133
rect 3322 2133 3442 2171
rect 3322 2117 3356 2133
rect 3230 2099 3246 2117
rect 3162 2083 3246 2099
rect 3340 2099 3356 2117
rect 3408 2117 3442 2133
rect 3500 2133 3620 2171
rect 3500 2117 3534 2133
rect 3408 2099 3424 2117
rect 3340 2083 3424 2099
rect 3518 2099 3534 2117
rect 3586 2117 3620 2133
rect 3874 2133 3994 2171
rect 3874 2117 3908 2133
rect 3586 2099 3602 2117
rect 3518 2083 3602 2099
rect 3892 2099 3908 2117
rect 3960 2117 3994 2133
rect 4052 2133 4172 2171
rect 4052 2117 4086 2133
rect 3960 2099 3976 2117
rect 3892 2083 3976 2099
rect 4070 2099 4086 2117
rect 4138 2117 4172 2133
rect 4230 2133 4350 2171
rect 4230 2117 4264 2133
rect 4138 2099 4154 2117
rect 4070 2083 4154 2099
rect 4248 2099 4264 2117
rect 4316 2117 4350 2133
rect 4408 2133 4528 2171
rect 4408 2117 4442 2133
rect 4316 2099 4332 2117
rect 4248 2083 4332 2099
rect 4426 2099 4442 2117
rect 4494 2117 4528 2133
rect 4586 2133 4706 2171
rect 4586 2117 4620 2133
rect 4494 2099 4510 2117
rect 4426 2083 4510 2099
rect 4604 2099 4620 2117
rect 4672 2117 4706 2133
rect 4764 2133 4884 2171
rect 4764 2117 4798 2133
rect 4672 2099 4688 2117
rect 4604 2083 4688 2099
rect 4782 2099 4798 2117
rect 4850 2117 4884 2133
rect 4942 2133 5062 2171
rect 4942 2117 4976 2133
rect 4850 2099 4866 2117
rect 4782 2083 4866 2099
rect 4960 2099 4976 2117
rect 5028 2117 5062 2133
rect 5120 2133 5240 2171
rect 5120 2117 5154 2133
rect 5028 2099 5044 2117
rect 4960 2083 5044 2099
rect 5138 2099 5154 2117
rect 5206 2117 5240 2133
rect 5298 2133 5418 2171
rect 5298 2117 5332 2133
rect 5206 2099 5222 2117
rect 5138 2083 5222 2099
rect 5316 2099 5332 2117
rect 5384 2117 5418 2133
rect 5476 2133 5596 2171
rect 5476 2117 5510 2133
rect 5384 2099 5400 2117
rect 5316 2083 5400 2099
rect 5494 2099 5510 2117
rect 5562 2117 5596 2133
rect 5654 2133 5774 2171
rect 5654 2117 5688 2133
rect 5562 2099 5578 2117
rect 5494 2083 5578 2099
rect 5672 2099 5688 2117
rect 5740 2117 5774 2133
rect 5832 2133 5952 2171
rect 5832 2117 5866 2133
rect 5740 2099 5756 2117
rect 5672 2083 5756 2099
rect 5850 2099 5866 2117
rect 5918 2117 5952 2133
rect 6010 2133 6130 2171
rect 6010 2117 6044 2133
rect 5918 2099 5934 2117
rect 5850 2083 5934 2099
rect 6028 2099 6044 2117
rect 6096 2117 6130 2133
rect 6188 2133 6308 2171
rect 6188 2117 6222 2133
rect 6096 2099 6112 2117
rect 6028 2083 6112 2099
rect 6206 2099 6222 2117
rect 6274 2117 6308 2133
rect 6366 2133 6486 2171
rect 6366 2117 6400 2133
rect 6274 2099 6290 2117
rect 6206 2083 6290 2099
rect 6384 2099 6400 2117
rect 6452 2117 6486 2133
rect 6544 2133 6664 2171
rect 6544 2117 6578 2133
rect 6452 2099 6468 2117
rect 6384 2083 6468 2099
rect 6562 2099 6578 2117
rect 6630 2117 6664 2133
rect 6722 2133 6842 2171
rect 6722 2117 6756 2133
rect 6630 2099 6646 2117
rect 6562 2083 6646 2099
rect 6740 2099 6756 2117
rect 6808 2117 6842 2133
rect 6900 2133 7020 2171
rect 6900 2117 6934 2133
rect 6808 2099 6824 2117
rect 6740 2083 6824 2099
rect 6918 2099 6934 2117
rect 6986 2117 7020 2133
rect 6986 2099 7002 2117
rect 6918 2083 7002 2099
rect 492 2023 576 2039
rect 492 2005 508 2023
rect 474 1989 508 2005
rect 560 2005 576 2023
rect 670 2023 754 2039
rect 670 2005 686 2023
rect 560 1989 594 2005
rect 474 1951 594 1989
rect 652 1989 686 2005
rect 738 2005 754 2023
rect 848 2023 932 2039
rect 848 2005 864 2023
rect 738 1989 772 2005
rect 652 1951 772 1989
rect 830 1989 864 2005
rect 916 2005 932 2023
rect 1026 2023 1110 2039
rect 1026 2005 1042 2023
rect 916 1989 950 2005
rect 830 1951 950 1989
rect 1008 1989 1042 2005
rect 1094 2005 1110 2023
rect 1204 2023 1288 2039
rect 1204 2005 1220 2023
rect 1094 1989 1128 2005
rect 1008 1951 1128 1989
rect 1186 1989 1220 2005
rect 1272 2005 1288 2023
rect 1382 2023 1466 2039
rect 1382 2005 1398 2023
rect 1272 1989 1306 2005
rect 1186 1951 1306 1989
rect 1364 1989 1398 2005
rect 1450 2005 1466 2023
rect 1560 2023 1644 2039
rect 1560 2005 1576 2023
rect 1450 1989 1484 2005
rect 1364 1951 1484 1989
rect 1542 1989 1576 2005
rect 1628 2005 1644 2023
rect 1738 2023 1822 2039
rect 1738 2005 1754 2023
rect 1628 1989 1662 2005
rect 1542 1951 1662 1989
rect 1720 1989 1754 2005
rect 1806 2005 1822 2023
rect 1916 2023 2000 2039
rect 1916 2005 1932 2023
rect 1806 1989 1840 2005
rect 1720 1951 1840 1989
rect 1898 1989 1932 2005
rect 1984 2005 2000 2023
rect 2094 2023 2178 2039
rect 2094 2005 2110 2023
rect 1984 1989 2018 2005
rect 1898 1951 2018 1989
rect 2076 1989 2110 2005
rect 2162 2005 2178 2023
rect 2272 2023 2356 2039
rect 2272 2005 2288 2023
rect 2162 1989 2196 2005
rect 2076 1951 2196 1989
rect 2254 1989 2288 2005
rect 2340 2005 2356 2023
rect 2450 2023 2534 2039
rect 2450 2005 2466 2023
rect 2340 1989 2374 2005
rect 2254 1951 2374 1989
rect 2432 1989 2466 2005
rect 2518 2005 2534 2023
rect 2628 2023 2712 2039
rect 2628 2005 2644 2023
rect 2518 1989 2552 2005
rect 2432 1951 2552 1989
rect 2610 1989 2644 2005
rect 2696 2005 2712 2023
rect 2806 2023 2890 2039
rect 2806 2005 2822 2023
rect 2696 1989 2730 2005
rect 2610 1951 2730 1989
rect 2788 1989 2822 2005
rect 2874 2005 2890 2023
rect 2984 2023 3068 2039
rect 2984 2005 3000 2023
rect 2874 1989 2908 2005
rect 2788 1951 2908 1989
rect 2966 1989 3000 2005
rect 3052 2005 3068 2023
rect 3162 2023 3246 2039
rect 3162 2005 3178 2023
rect 3052 1989 3086 2005
rect 2966 1951 3086 1989
rect 3144 1989 3178 2005
rect 3230 2005 3246 2023
rect 3340 2023 3424 2039
rect 3340 2005 3356 2023
rect 3230 1989 3264 2005
rect 3144 1951 3264 1989
rect 3322 1989 3356 2005
rect 3408 2005 3424 2023
rect 3518 2023 3602 2039
rect 3518 2005 3534 2023
rect 3408 1989 3442 2005
rect 3322 1951 3442 1989
rect 3500 1989 3534 2005
rect 3586 2005 3602 2023
rect 3892 2023 3976 2039
rect 3892 2005 3908 2023
rect 3586 1989 3620 2005
rect 3500 1951 3620 1989
rect 3874 1989 3908 2005
rect 3960 2005 3976 2023
rect 4070 2023 4154 2039
rect 4070 2005 4086 2023
rect 3960 1989 3994 2005
rect 3874 1951 3994 1989
rect 4052 1989 4086 2005
rect 4138 2005 4154 2023
rect 4248 2023 4332 2039
rect 4248 2005 4264 2023
rect 4138 1989 4172 2005
rect 4052 1951 4172 1989
rect 4230 1989 4264 2005
rect 4316 2005 4332 2023
rect 4426 2023 4510 2039
rect 4426 2005 4442 2023
rect 4316 1989 4350 2005
rect 4230 1951 4350 1989
rect 4408 1989 4442 2005
rect 4494 2005 4510 2023
rect 4604 2023 4688 2039
rect 4604 2005 4620 2023
rect 4494 1989 4528 2005
rect 4408 1951 4528 1989
rect 4586 1989 4620 2005
rect 4672 2005 4688 2023
rect 4782 2023 4866 2039
rect 4782 2005 4798 2023
rect 4672 1989 4706 2005
rect 4586 1951 4706 1989
rect 4764 1989 4798 2005
rect 4850 2005 4866 2023
rect 4960 2023 5044 2039
rect 4960 2005 4976 2023
rect 4850 1989 4884 2005
rect 4764 1951 4884 1989
rect 4942 1989 4976 2005
rect 5028 2005 5044 2023
rect 5138 2023 5222 2039
rect 5138 2005 5154 2023
rect 5028 1989 5062 2005
rect 4942 1951 5062 1989
rect 5120 1989 5154 2005
rect 5206 2005 5222 2023
rect 5316 2023 5400 2039
rect 5316 2005 5332 2023
rect 5206 1989 5240 2005
rect 5120 1951 5240 1989
rect 5298 1989 5332 2005
rect 5384 2005 5400 2023
rect 5494 2023 5578 2039
rect 5494 2005 5510 2023
rect 5384 1989 5418 2005
rect 5298 1951 5418 1989
rect 5476 1989 5510 2005
rect 5562 2005 5578 2023
rect 5672 2023 5756 2039
rect 5672 2005 5688 2023
rect 5562 1989 5596 2005
rect 5476 1951 5596 1989
rect 5654 1989 5688 2005
rect 5740 2005 5756 2023
rect 5850 2023 5934 2039
rect 5850 2005 5866 2023
rect 5740 1989 5774 2005
rect 5654 1951 5774 1989
rect 5832 1989 5866 2005
rect 5918 2005 5934 2023
rect 6028 2023 6112 2039
rect 6028 2005 6044 2023
rect 5918 1989 5952 2005
rect 5832 1951 5952 1989
rect 6010 1989 6044 2005
rect 6096 2005 6112 2023
rect 6206 2023 6290 2039
rect 6206 2005 6222 2023
rect 6096 1989 6130 2005
rect 6010 1951 6130 1989
rect 6188 1989 6222 2005
rect 6274 2005 6290 2023
rect 6384 2023 6468 2039
rect 6384 2005 6400 2023
rect 6274 1989 6308 2005
rect 6188 1951 6308 1989
rect 6366 1989 6400 2005
rect 6452 2005 6468 2023
rect 6562 2023 6646 2039
rect 6562 2005 6578 2023
rect 6452 1989 6486 2005
rect 6366 1951 6486 1989
rect 6544 1989 6578 2005
rect 6630 2005 6646 2023
rect 6740 2023 6824 2039
rect 6740 2005 6756 2023
rect 6630 1989 6664 2005
rect 6544 1951 6664 1989
rect 6722 1989 6756 2005
rect 6808 2005 6824 2023
rect 6918 2023 7002 2039
rect 6918 2005 6934 2023
rect 6808 1989 6842 2005
rect 6722 1951 6842 1989
rect 6900 1989 6934 2005
rect 6986 2005 7002 2023
rect 7621 2023 7705 2039
rect 7621 2006 7637 2023
rect 6986 1989 7020 2005
rect 6900 1951 7020 1989
rect 7603 1989 7637 2006
rect 7689 2006 7705 2023
rect 7799 2023 7883 2039
rect 7799 2006 7815 2023
rect 7689 1989 7723 2006
rect 7603 1951 7723 1989
rect 7781 1989 7815 2006
rect 7867 2006 7883 2023
rect 7977 2023 8061 2039
rect 7977 2006 7993 2023
rect 7867 1989 7901 2006
rect 7781 1951 7901 1989
rect 7959 1989 7993 2006
rect 8045 2006 8061 2023
rect 8155 2023 8239 2039
rect 8155 2006 8171 2023
rect 8045 1989 8079 2006
rect 7959 1951 8079 1989
rect 8137 1989 8171 2006
rect 8223 2006 8239 2023
rect 8333 2023 8417 2039
rect 8333 2006 8349 2023
rect 8223 1989 8257 2006
rect 8137 1951 8257 1989
rect 8315 1989 8349 2006
rect 8401 2006 8417 2023
rect 8511 2023 8595 2039
rect 8511 2006 8527 2023
rect 8401 1989 8435 2006
rect 8315 1951 8435 1989
rect 8493 1989 8527 2006
rect 8579 2006 8595 2023
rect 8689 2023 8773 2039
rect 8689 2006 8705 2023
rect 8579 1989 8613 2006
rect 8493 1951 8613 1989
rect 8671 1989 8705 2006
rect 8757 2006 8773 2023
rect 8867 2023 8951 2039
rect 8867 2006 8883 2023
rect 8757 1989 8791 2006
rect 8671 1951 8791 1989
rect 8849 1989 8883 2006
rect 8935 2006 8951 2023
rect 9045 2023 9129 2039
rect 9045 2006 9061 2023
rect 8935 1989 8969 2006
rect 8849 1951 8969 1989
rect 9027 1989 9061 2006
rect 9113 2006 9129 2023
rect 9223 2023 9307 2039
rect 9223 2006 9239 2023
rect 9113 1989 9147 2006
rect 9027 1951 9147 1989
rect 9205 1989 9239 2006
rect 9291 2006 9307 2023
rect 9401 2023 9485 2039
rect 9401 2006 9417 2023
rect 9291 1989 9325 2006
rect 9205 1951 9325 1989
rect 9383 1989 9417 2006
rect 9469 2006 9485 2023
rect 9579 2023 9663 2039
rect 9579 2006 9595 2023
rect 9469 1989 9503 2006
rect 9383 1951 9503 1989
rect 9561 1989 9595 2006
rect 9647 2006 9663 2023
rect 9757 2023 9841 2039
rect 9757 2006 9773 2023
rect 9647 1989 9681 2006
rect 9561 1951 9681 1989
rect 9739 1989 9773 2006
rect 9825 2006 9841 2023
rect 9935 2023 10019 2039
rect 9935 2006 9951 2023
rect 9825 1989 9859 2006
rect 9739 1951 9859 1989
rect 9917 1989 9951 2006
rect 10003 2006 10019 2023
rect 10308 2023 10392 2039
rect 10308 2006 10324 2023
rect 10003 1989 10037 2006
rect 9917 1951 10037 1989
rect 10290 1989 10324 2006
rect 10376 2006 10392 2023
rect 10486 2023 10570 2039
rect 10486 2006 10502 2023
rect 10376 1989 10410 2006
rect 10290 1951 10410 1989
rect 10468 1989 10502 2006
rect 10554 2006 10570 2023
rect 10664 2023 10748 2039
rect 10664 2006 10680 2023
rect 10554 1989 10588 2006
rect 10468 1951 10588 1989
rect 10646 1989 10680 2006
rect 10732 2006 10748 2023
rect 10842 2023 10926 2039
rect 10842 2006 10858 2023
rect 10732 1989 10766 2006
rect 10646 1951 10766 1989
rect 10824 1989 10858 2006
rect 10910 2006 10926 2023
rect 11020 2023 11104 2039
rect 11020 2006 11036 2023
rect 10910 1989 10944 2006
rect 10824 1951 10944 1989
rect 11002 1989 11036 2006
rect 11088 2006 11104 2023
rect 11198 2023 11282 2039
rect 11198 2006 11214 2023
rect 11088 1989 11122 2006
rect 11002 1951 11122 1989
rect 11180 1989 11214 2006
rect 11266 2006 11282 2023
rect 11376 2023 11460 2039
rect 11376 2006 11392 2023
rect 11266 1989 11300 2006
rect 11180 1951 11300 1989
rect 11358 1989 11392 2006
rect 11444 2006 11460 2023
rect 11554 2023 11638 2039
rect 11554 2006 11570 2023
rect 11444 1989 11478 2006
rect 11358 1951 11478 1989
rect 11536 1989 11570 2006
rect 11622 2006 11638 2023
rect 11732 2023 11816 2039
rect 11732 2006 11748 2023
rect 11622 1989 11656 2006
rect 11536 1951 11656 1989
rect 11714 1989 11748 2006
rect 11800 2006 11816 2023
rect 11910 2023 11994 2039
rect 11910 2006 11926 2023
rect 11800 1989 11834 2006
rect 11714 1951 11834 1989
rect 11892 1989 11926 2006
rect 11978 2006 11994 2023
rect 12088 2023 12172 2039
rect 12088 2006 12104 2023
rect 11978 1989 12012 2006
rect 11892 1951 12012 1989
rect 12070 1989 12104 2006
rect 12156 2006 12172 2023
rect 12266 2023 12350 2039
rect 12266 2006 12282 2023
rect 12156 1989 12190 2006
rect 12070 1951 12190 1989
rect 12248 1989 12282 2006
rect 12334 2006 12350 2023
rect 12444 2023 12528 2039
rect 12444 2006 12460 2023
rect 12334 1989 12368 2006
rect 12248 1951 12368 1989
rect 12426 1989 12460 2006
rect 12512 2006 12528 2023
rect 12622 2023 12706 2039
rect 12622 2006 12638 2023
rect 12512 1989 12546 2006
rect 12426 1951 12546 1989
rect 12604 1989 12638 2006
rect 12690 2006 12706 2023
rect 12690 1989 12724 2006
rect 12604 1951 12724 1989
rect 474 1633 594 1671
rect 474 1617 508 1633
rect 492 1599 508 1617
rect 560 1617 594 1633
rect 652 1633 772 1671
rect 652 1617 686 1633
rect 560 1599 576 1617
rect 492 1583 576 1599
rect 670 1599 686 1617
rect 738 1617 772 1633
rect 830 1633 950 1671
rect 830 1617 864 1633
rect 738 1599 754 1617
rect 670 1583 754 1599
rect 848 1599 864 1617
rect 916 1617 950 1633
rect 1008 1633 1128 1671
rect 1008 1617 1042 1633
rect 916 1599 932 1617
rect 848 1583 932 1599
rect 1026 1599 1042 1617
rect 1094 1617 1128 1633
rect 1186 1633 1306 1671
rect 1186 1617 1220 1633
rect 1094 1599 1110 1617
rect 1026 1583 1110 1599
rect 1204 1599 1220 1617
rect 1272 1617 1306 1633
rect 1364 1633 1484 1671
rect 1364 1617 1398 1633
rect 1272 1599 1288 1617
rect 1204 1583 1288 1599
rect 1382 1599 1398 1617
rect 1450 1617 1484 1633
rect 1542 1633 1662 1671
rect 1542 1617 1576 1633
rect 1450 1599 1466 1617
rect 1382 1583 1466 1599
rect 1560 1599 1576 1617
rect 1628 1617 1662 1633
rect 1720 1633 1840 1671
rect 1720 1617 1754 1633
rect 1628 1599 1644 1617
rect 1560 1583 1644 1599
rect 1738 1599 1754 1617
rect 1806 1617 1840 1633
rect 1898 1633 2018 1671
rect 1898 1617 1932 1633
rect 1806 1599 1822 1617
rect 1738 1583 1822 1599
rect 1916 1599 1932 1617
rect 1984 1617 2018 1633
rect 2076 1633 2196 1671
rect 2076 1617 2110 1633
rect 1984 1599 2000 1617
rect 1916 1583 2000 1599
rect 2094 1599 2110 1617
rect 2162 1617 2196 1633
rect 2254 1633 2374 1671
rect 2254 1617 2288 1633
rect 2162 1599 2178 1617
rect 2094 1583 2178 1599
rect 2272 1599 2288 1617
rect 2340 1617 2374 1633
rect 2432 1633 2552 1671
rect 2432 1617 2466 1633
rect 2340 1599 2356 1617
rect 2272 1583 2356 1599
rect 2450 1599 2466 1617
rect 2518 1617 2552 1633
rect 2610 1633 2730 1671
rect 2610 1617 2644 1633
rect 2518 1599 2534 1617
rect 2450 1583 2534 1599
rect 2628 1599 2644 1617
rect 2696 1617 2730 1633
rect 2788 1633 2908 1671
rect 2788 1617 2822 1633
rect 2696 1599 2712 1617
rect 2628 1583 2712 1599
rect 2806 1599 2822 1617
rect 2874 1617 2908 1633
rect 2966 1633 3086 1671
rect 2966 1617 3000 1633
rect 2874 1599 2890 1617
rect 2806 1583 2890 1599
rect 2984 1599 3000 1617
rect 3052 1617 3086 1633
rect 3144 1633 3264 1671
rect 3144 1617 3178 1633
rect 3052 1599 3068 1617
rect 2984 1583 3068 1599
rect 3162 1599 3178 1617
rect 3230 1617 3264 1633
rect 3322 1633 3442 1671
rect 3322 1617 3356 1633
rect 3230 1599 3246 1617
rect 3162 1583 3246 1599
rect 3340 1599 3356 1617
rect 3408 1617 3442 1633
rect 3500 1633 3620 1671
rect 3500 1617 3534 1633
rect 3408 1599 3424 1617
rect 3340 1583 3424 1599
rect 3518 1599 3534 1617
rect 3586 1617 3620 1633
rect 3874 1633 3994 1671
rect 3874 1617 3908 1633
rect 3586 1599 3602 1617
rect 3518 1583 3602 1599
rect 3892 1599 3908 1617
rect 3960 1617 3994 1633
rect 4052 1633 4172 1671
rect 4052 1617 4086 1633
rect 3960 1599 3976 1617
rect 3892 1583 3976 1599
rect 4070 1599 4086 1617
rect 4138 1617 4172 1633
rect 4230 1633 4350 1671
rect 4230 1617 4264 1633
rect 4138 1599 4154 1617
rect 4070 1583 4154 1599
rect 4248 1599 4264 1617
rect 4316 1617 4350 1633
rect 4408 1633 4528 1671
rect 4408 1617 4442 1633
rect 4316 1599 4332 1617
rect 4248 1583 4332 1599
rect 4426 1599 4442 1617
rect 4494 1617 4528 1633
rect 4586 1633 4706 1671
rect 4586 1617 4620 1633
rect 4494 1599 4510 1617
rect 4426 1583 4510 1599
rect 4604 1599 4620 1617
rect 4672 1617 4706 1633
rect 4764 1633 4884 1671
rect 4764 1617 4798 1633
rect 4672 1599 4688 1617
rect 4604 1583 4688 1599
rect 4782 1599 4798 1617
rect 4850 1617 4884 1633
rect 4942 1633 5062 1671
rect 4942 1617 4976 1633
rect 4850 1599 4866 1617
rect 4782 1583 4866 1599
rect 4960 1599 4976 1617
rect 5028 1617 5062 1633
rect 5120 1633 5240 1671
rect 5120 1617 5154 1633
rect 5028 1599 5044 1617
rect 4960 1583 5044 1599
rect 5138 1599 5154 1617
rect 5206 1617 5240 1633
rect 5298 1633 5418 1671
rect 5298 1617 5332 1633
rect 5206 1599 5222 1617
rect 5138 1583 5222 1599
rect 5316 1599 5332 1617
rect 5384 1617 5418 1633
rect 5476 1633 5596 1671
rect 5476 1617 5510 1633
rect 5384 1599 5400 1617
rect 5316 1583 5400 1599
rect 5494 1599 5510 1617
rect 5562 1617 5596 1633
rect 5654 1633 5774 1671
rect 5654 1617 5688 1633
rect 5562 1599 5578 1617
rect 5494 1583 5578 1599
rect 5672 1599 5688 1617
rect 5740 1617 5774 1633
rect 5832 1633 5952 1671
rect 5832 1617 5866 1633
rect 5740 1599 5756 1617
rect 5672 1583 5756 1599
rect 5850 1599 5866 1617
rect 5918 1617 5952 1633
rect 6010 1633 6130 1671
rect 6010 1617 6044 1633
rect 5918 1599 5934 1617
rect 5850 1583 5934 1599
rect 6028 1599 6044 1617
rect 6096 1617 6130 1633
rect 6188 1633 6308 1671
rect 6188 1617 6222 1633
rect 6096 1599 6112 1617
rect 6028 1583 6112 1599
rect 6206 1599 6222 1617
rect 6274 1617 6308 1633
rect 6366 1633 6486 1671
rect 6366 1617 6400 1633
rect 6274 1599 6290 1617
rect 6206 1583 6290 1599
rect 6384 1599 6400 1617
rect 6452 1617 6486 1633
rect 6544 1633 6664 1671
rect 6544 1617 6578 1633
rect 6452 1599 6468 1617
rect 6384 1583 6468 1599
rect 6562 1599 6578 1617
rect 6630 1617 6664 1633
rect 6722 1633 6842 1671
rect 6722 1617 6756 1633
rect 6630 1599 6646 1617
rect 6562 1583 6646 1599
rect 6740 1599 6756 1617
rect 6808 1617 6842 1633
rect 6900 1633 7020 1671
rect 6900 1617 6934 1633
rect 6808 1599 6824 1617
rect 6740 1583 6824 1599
rect 6918 1599 6934 1617
rect 6986 1617 7020 1633
rect 7603 1633 7723 1671
rect 6986 1599 7002 1617
rect 7603 1616 7637 1633
rect 6918 1583 7002 1599
rect 7621 1599 7637 1616
rect 7689 1616 7723 1633
rect 7781 1633 7901 1671
rect 7781 1616 7815 1633
rect 7689 1599 7705 1616
rect 7621 1583 7705 1599
rect 7799 1599 7815 1616
rect 7867 1616 7901 1633
rect 7959 1633 8079 1671
rect 7959 1616 7993 1633
rect 7867 1599 7883 1616
rect 7799 1583 7883 1599
rect 7977 1599 7993 1616
rect 8045 1616 8079 1633
rect 8137 1633 8257 1671
rect 8137 1616 8171 1633
rect 8045 1599 8061 1616
rect 7977 1583 8061 1599
rect 8155 1599 8171 1616
rect 8223 1616 8257 1633
rect 8315 1633 8435 1671
rect 8315 1616 8349 1633
rect 8223 1599 8239 1616
rect 8155 1583 8239 1599
rect 8333 1599 8349 1616
rect 8401 1616 8435 1633
rect 8493 1633 8613 1671
rect 8493 1616 8527 1633
rect 8401 1599 8417 1616
rect 8333 1583 8417 1599
rect 8511 1599 8527 1616
rect 8579 1616 8613 1633
rect 8671 1633 8791 1671
rect 8671 1616 8705 1633
rect 8579 1599 8595 1616
rect 8511 1583 8595 1599
rect 8689 1599 8705 1616
rect 8757 1616 8791 1633
rect 8849 1633 8969 1671
rect 8849 1616 8883 1633
rect 8757 1599 8773 1616
rect 8689 1583 8773 1599
rect 8867 1599 8883 1616
rect 8935 1616 8969 1633
rect 9027 1633 9147 1671
rect 9027 1616 9061 1633
rect 8935 1599 8951 1616
rect 8867 1583 8951 1599
rect 9045 1599 9061 1616
rect 9113 1616 9147 1633
rect 9205 1633 9325 1671
rect 9205 1616 9239 1633
rect 9113 1599 9129 1616
rect 9045 1583 9129 1599
rect 9223 1599 9239 1616
rect 9291 1616 9325 1633
rect 9383 1633 9503 1671
rect 9383 1616 9417 1633
rect 9291 1599 9307 1616
rect 9223 1583 9307 1599
rect 9401 1599 9417 1616
rect 9469 1616 9503 1633
rect 9561 1633 9681 1671
rect 9561 1616 9595 1633
rect 9469 1599 9485 1616
rect 9401 1583 9485 1599
rect 9579 1599 9595 1616
rect 9647 1616 9681 1633
rect 9739 1633 9859 1671
rect 9739 1616 9773 1633
rect 9647 1599 9663 1616
rect 9579 1583 9663 1599
rect 9757 1599 9773 1616
rect 9825 1616 9859 1633
rect 9917 1633 10037 1671
rect 9917 1616 9951 1633
rect 9825 1599 9841 1616
rect 9757 1583 9841 1599
rect 9935 1599 9951 1616
rect 10003 1616 10037 1633
rect 10290 1633 10410 1671
rect 10290 1616 10324 1633
rect 10003 1599 10019 1616
rect 9935 1583 10019 1599
rect 10308 1599 10324 1616
rect 10376 1616 10410 1633
rect 10468 1633 10588 1671
rect 10468 1616 10502 1633
rect 10376 1599 10392 1616
rect 10308 1583 10392 1599
rect 10486 1599 10502 1616
rect 10554 1616 10588 1633
rect 10646 1633 10766 1671
rect 10646 1616 10680 1633
rect 10554 1599 10570 1616
rect 10486 1583 10570 1599
rect 10664 1599 10680 1616
rect 10732 1616 10766 1633
rect 10824 1633 10944 1671
rect 10824 1616 10858 1633
rect 10732 1599 10748 1616
rect 10664 1583 10748 1599
rect 10842 1599 10858 1616
rect 10910 1616 10944 1633
rect 11002 1633 11122 1671
rect 11002 1616 11036 1633
rect 10910 1599 10926 1616
rect 10842 1583 10926 1599
rect 11020 1599 11036 1616
rect 11088 1616 11122 1633
rect 11180 1633 11300 1671
rect 11180 1616 11214 1633
rect 11088 1599 11104 1616
rect 11020 1583 11104 1599
rect 11198 1599 11214 1616
rect 11266 1616 11300 1633
rect 11358 1633 11478 1671
rect 11358 1616 11392 1633
rect 11266 1599 11282 1616
rect 11198 1583 11282 1599
rect 11376 1599 11392 1616
rect 11444 1616 11478 1633
rect 11536 1633 11656 1671
rect 11536 1616 11570 1633
rect 11444 1599 11460 1616
rect 11376 1583 11460 1599
rect 11554 1599 11570 1616
rect 11622 1616 11656 1633
rect 11714 1633 11834 1671
rect 11714 1616 11748 1633
rect 11622 1599 11638 1616
rect 11554 1583 11638 1599
rect 11732 1599 11748 1616
rect 11800 1616 11834 1633
rect 11892 1633 12012 1671
rect 11892 1616 11926 1633
rect 11800 1599 11816 1616
rect 11732 1583 11816 1599
rect 11910 1599 11926 1616
rect 11978 1616 12012 1633
rect 12070 1633 12190 1671
rect 12070 1616 12104 1633
rect 11978 1599 11994 1616
rect 11910 1583 11994 1599
rect 12088 1599 12104 1616
rect 12156 1616 12190 1633
rect 12248 1633 12368 1671
rect 12248 1616 12282 1633
rect 12156 1599 12172 1616
rect 12088 1583 12172 1599
rect 12266 1599 12282 1616
rect 12334 1616 12368 1633
rect 12426 1633 12546 1671
rect 12426 1616 12460 1633
rect 12334 1599 12350 1616
rect 12266 1583 12350 1599
rect 12444 1599 12460 1616
rect 12512 1616 12546 1633
rect 12604 1633 12724 1671
rect 12604 1616 12638 1633
rect 12512 1599 12528 1616
rect 12444 1583 12528 1599
rect 12622 1599 12638 1616
rect 12690 1616 12724 1633
rect 12690 1599 12706 1616
rect 12622 1583 12706 1599
rect 492 1523 576 1539
rect 492 1505 508 1523
rect 474 1489 508 1505
rect 560 1505 576 1523
rect 670 1523 754 1539
rect 670 1505 686 1523
rect 560 1489 594 1505
rect 474 1451 594 1489
rect 652 1489 686 1505
rect 738 1505 754 1523
rect 848 1523 932 1539
rect 848 1505 864 1523
rect 738 1489 772 1505
rect 652 1451 772 1489
rect 830 1489 864 1505
rect 916 1505 932 1523
rect 1026 1523 1110 1539
rect 1026 1505 1042 1523
rect 916 1489 950 1505
rect 830 1451 950 1489
rect 1008 1489 1042 1505
rect 1094 1505 1110 1523
rect 1204 1523 1288 1539
rect 1204 1505 1220 1523
rect 1094 1489 1128 1505
rect 1008 1451 1128 1489
rect 1186 1489 1220 1505
rect 1272 1505 1288 1523
rect 1382 1523 1466 1539
rect 1382 1505 1398 1523
rect 1272 1489 1306 1505
rect 1186 1451 1306 1489
rect 1364 1489 1398 1505
rect 1450 1505 1466 1523
rect 1560 1523 1644 1539
rect 1560 1505 1576 1523
rect 1450 1489 1484 1505
rect 1364 1451 1484 1489
rect 1542 1489 1576 1505
rect 1628 1505 1644 1523
rect 1738 1523 1822 1539
rect 1738 1505 1754 1523
rect 1628 1489 1662 1505
rect 1542 1451 1662 1489
rect 1720 1489 1754 1505
rect 1806 1505 1822 1523
rect 1916 1523 2000 1539
rect 1916 1505 1932 1523
rect 1806 1489 1840 1505
rect 1720 1451 1840 1489
rect 1898 1489 1932 1505
rect 1984 1505 2000 1523
rect 2094 1523 2178 1539
rect 2094 1505 2110 1523
rect 1984 1489 2018 1505
rect 1898 1451 2018 1489
rect 2076 1489 2110 1505
rect 2162 1505 2178 1523
rect 2272 1523 2356 1539
rect 2272 1505 2288 1523
rect 2162 1489 2196 1505
rect 2076 1451 2196 1489
rect 2254 1489 2288 1505
rect 2340 1505 2356 1523
rect 2450 1523 2534 1539
rect 2450 1505 2466 1523
rect 2340 1489 2374 1505
rect 2254 1451 2374 1489
rect 2432 1489 2466 1505
rect 2518 1505 2534 1523
rect 2628 1523 2712 1539
rect 2628 1505 2644 1523
rect 2518 1489 2552 1505
rect 2432 1451 2552 1489
rect 2610 1489 2644 1505
rect 2696 1505 2712 1523
rect 2806 1523 2890 1539
rect 2806 1505 2822 1523
rect 2696 1489 2730 1505
rect 2610 1451 2730 1489
rect 2788 1489 2822 1505
rect 2874 1505 2890 1523
rect 2984 1523 3068 1539
rect 2984 1505 3000 1523
rect 2874 1489 2908 1505
rect 2788 1451 2908 1489
rect 2966 1489 3000 1505
rect 3052 1505 3068 1523
rect 3162 1523 3246 1539
rect 3162 1505 3178 1523
rect 3052 1489 3086 1505
rect 2966 1451 3086 1489
rect 3144 1489 3178 1505
rect 3230 1505 3246 1523
rect 3340 1523 3424 1539
rect 3340 1505 3356 1523
rect 3230 1489 3264 1505
rect 3144 1451 3264 1489
rect 3322 1489 3356 1505
rect 3408 1505 3424 1523
rect 3518 1523 3602 1539
rect 3518 1505 3534 1523
rect 3408 1489 3442 1505
rect 3322 1451 3442 1489
rect 3500 1489 3534 1505
rect 3586 1505 3602 1523
rect 3892 1523 3976 1539
rect 3892 1505 3908 1523
rect 3586 1489 3620 1505
rect 3500 1451 3620 1489
rect 3874 1489 3908 1505
rect 3960 1505 3976 1523
rect 4070 1523 4154 1539
rect 4070 1505 4086 1523
rect 3960 1489 3994 1505
rect 3874 1451 3994 1489
rect 4052 1489 4086 1505
rect 4138 1505 4154 1523
rect 4248 1523 4332 1539
rect 4248 1505 4264 1523
rect 4138 1489 4172 1505
rect 4052 1451 4172 1489
rect 4230 1489 4264 1505
rect 4316 1505 4332 1523
rect 4426 1523 4510 1539
rect 4426 1505 4442 1523
rect 4316 1489 4350 1505
rect 4230 1451 4350 1489
rect 4408 1489 4442 1505
rect 4494 1505 4510 1523
rect 4604 1523 4688 1539
rect 4604 1505 4620 1523
rect 4494 1489 4528 1505
rect 4408 1451 4528 1489
rect 4586 1489 4620 1505
rect 4672 1505 4688 1523
rect 4782 1523 4866 1539
rect 4782 1505 4798 1523
rect 4672 1489 4706 1505
rect 4586 1451 4706 1489
rect 4764 1489 4798 1505
rect 4850 1505 4866 1523
rect 4960 1523 5044 1539
rect 4960 1505 4976 1523
rect 4850 1489 4884 1505
rect 4764 1451 4884 1489
rect 4942 1489 4976 1505
rect 5028 1505 5044 1523
rect 5138 1523 5222 1539
rect 5138 1505 5154 1523
rect 5028 1489 5062 1505
rect 4942 1451 5062 1489
rect 5120 1489 5154 1505
rect 5206 1505 5222 1523
rect 5316 1523 5400 1539
rect 5316 1505 5332 1523
rect 5206 1489 5240 1505
rect 5120 1451 5240 1489
rect 5298 1489 5332 1505
rect 5384 1505 5400 1523
rect 5494 1523 5578 1539
rect 5494 1505 5510 1523
rect 5384 1489 5418 1505
rect 5298 1451 5418 1489
rect 5476 1489 5510 1505
rect 5562 1505 5578 1523
rect 5672 1523 5756 1539
rect 5672 1505 5688 1523
rect 5562 1489 5596 1505
rect 5476 1451 5596 1489
rect 5654 1489 5688 1505
rect 5740 1505 5756 1523
rect 5850 1523 5934 1539
rect 5850 1505 5866 1523
rect 5740 1489 5774 1505
rect 5654 1451 5774 1489
rect 5832 1489 5866 1505
rect 5918 1505 5934 1523
rect 6028 1523 6112 1539
rect 6028 1505 6044 1523
rect 5918 1489 5952 1505
rect 5832 1451 5952 1489
rect 6010 1489 6044 1505
rect 6096 1505 6112 1523
rect 6206 1523 6290 1539
rect 6206 1505 6222 1523
rect 6096 1489 6130 1505
rect 6010 1451 6130 1489
rect 6188 1489 6222 1505
rect 6274 1505 6290 1523
rect 6384 1523 6468 1539
rect 6384 1505 6400 1523
rect 6274 1489 6308 1505
rect 6188 1451 6308 1489
rect 6366 1489 6400 1505
rect 6452 1505 6468 1523
rect 6562 1523 6646 1539
rect 6562 1505 6578 1523
rect 6452 1489 6486 1505
rect 6366 1451 6486 1489
rect 6544 1489 6578 1505
rect 6630 1505 6646 1523
rect 6740 1523 6824 1539
rect 6740 1505 6756 1523
rect 6630 1489 6664 1505
rect 6544 1451 6664 1489
rect 6722 1489 6756 1505
rect 6808 1505 6824 1523
rect 6918 1523 7002 1539
rect 6918 1505 6934 1523
rect 6808 1489 6842 1505
rect 6722 1451 6842 1489
rect 6900 1489 6934 1505
rect 6986 1505 7002 1523
rect 7621 1523 7705 1539
rect 7621 1506 7637 1523
rect 6986 1489 7020 1505
rect 6900 1451 7020 1489
rect 7603 1489 7637 1506
rect 7689 1506 7705 1523
rect 7799 1523 7883 1539
rect 7799 1506 7815 1523
rect 7689 1489 7723 1506
rect 7603 1451 7723 1489
rect 7781 1489 7815 1506
rect 7867 1506 7883 1523
rect 7977 1523 8061 1539
rect 7977 1506 7993 1523
rect 7867 1489 7901 1506
rect 7781 1451 7901 1489
rect 7959 1489 7993 1506
rect 8045 1506 8061 1523
rect 8155 1523 8239 1539
rect 8155 1506 8171 1523
rect 8045 1489 8079 1506
rect 7959 1451 8079 1489
rect 8137 1489 8171 1506
rect 8223 1506 8239 1523
rect 8333 1523 8417 1539
rect 8333 1506 8349 1523
rect 8223 1489 8257 1506
rect 8137 1451 8257 1489
rect 8315 1489 8349 1506
rect 8401 1506 8417 1523
rect 8511 1523 8595 1539
rect 8511 1506 8527 1523
rect 8401 1489 8435 1506
rect 8315 1451 8435 1489
rect 8493 1489 8527 1506
rect 8579 1506 8595 1523
rect 8689 1523 8773 1539
rect 8689 1506 8705 1523
rect 8579 1489 8613 1506
rect 8493 1451 8613 1489
rect 8671 1489 8705 1506
rect 8757 1506 8773 1523
rect 8867 1523 8951 1539
rect 8867 1506 8883 1523
rect 8757 1489 8791 1506
rect 8671 1451 8791 1489
rect 8849 1489 8883 1506
rect 8935 1506 8951 1523
rect 9045 1523 9129 1539
rect 9045 1506 9061 1523
rect 8935 1489 8969 1506
rect 8849 1451 8969 1489
rect 9027 1489 9061 1506
rect 9113 1506 9129 1523
rect 9223 1523 9307 1539
rect 9223 1506 9239 1523
rect 9113 1489 9147 1506
rect 9027 1451 9147 1489
rect 9205 1489 9239 1506
rect 9291 1506 9307 1523
rect 9401 1523 9485 1539
rect 9401 1506 9417 1523
rect 9291 1489 9325 1506
rect 9205 1451 9325 1489
rect 9383 1489 9417 1506
rect 9469 1506 9485 1523
rect 9579 1523 9663 1539
rect 9579 1506 9595 1523
rect 9469 1489 9503 1506
rect 9383 1451 9503 1489
rect 9561 1489 9595 1506
rect 9647 1506 9663 1523
rect 9757 1523 9841 1539
rect 9757 1506 9773 1523
rect 9647 1489 9681 1506
rect 9561 1451 9681 1489
rect 9739 1489 9773 1506
rect 9825 1506 9841 1523
rect 9935 1523 10019 1539
rect 9935 1506 9951 1523
rect 9825 1489 9859 1506
rect 9739 1451 9859 1489
rect 9917 1489 9951 1506
rect 10003 1506 10019 1523
rect 10308 1523 10392 1539
rect 10308 1506 10324 1523
rect 10003 1489 10037 1506
rect 9917 1451 10037 1489
rect 10290 1489 10324 1506
rect 10376 1506 10392 1523
rect 10486 1523 10570 1539
rect 10486 1506 10502 1523
rect 10376 1489 10410 1506
rect 10290 1451 10410 1489
rect 10468 1489 10502 1506
rect 10554 1506 10570 1523
rect 10664 1523 10748 1539
rect 10664 1506 10680 1523
rect 10554 1489 10588 1506
rect 10468 1451 10588 1489
rect 10646 1489 10680 1506
rect 10732 1506 10748 1523
rect 10842 1523 10926 1539
rect 10842 1506 10858 1523
rect 10732 1489 10766 1506
rect 10646 1451 10766 1489
rect 10824 1489 10858 1506
rect 10910 1506 10926 1523
rect 11020 1523 11104 1539
rect 11020 1506 11036 1523
rect 10910 1489 10944 1506
rect 10824 1451 10944 1489
rect 11002 1489 11036 1506
rect 11088 1506 11104 1523
rect 11198 1523 11282 1539
rect 11198 1506 11214 1523
rect 11088 1489 11122 1506
rect 11002 1451 11122 1489
rect 11180 1489 11214 1506
rect 11266 1506 11282 1523
rect 11376 1523 11460 1539
rect 11376 1506 11392 1523
rect 11266 1489 11300 1506
rect 11180 1451 11300 1489
rect 11358 1489 11392 1506
rect 11444 1506 11460 1523
rect 11554 1523 11638 1539
rect 11554 1506 11570 1523
rect 11444 1489 11478 1506
rect 11358 1451 11478 1489
rect 11536 1489 11570 1506
rect 11622 1506 11638 1523
rect 11732 1523 11816 1539
rect 11732 1506 11748 1523
rect 11622 1489 11656 1506
rect 11536 1451 11656 1489
rect 11714 1489 11748 1506
rect 11800 1506 11816 1523
rect 11910 1523 11994 1539
rect 11910 1506 11926 1523
rect 11800 1489 11834 1506
rect 11714 1451 11834 1489
rect 11892 1489 11926 1506
rect 11978 1506 11994 1523
rect 12088 1523 12172 1539
rect 12088 1506 12104 1523
rect 11978 1489 12012 1506
rect 11892 1451 12012 1489
rect 12070 1489 12104 1506
rect 12156 1506 12172 1523
rect 12266 1523 12350 1539
rect 12266 1506 12282 1523
rect 12156 1489 12190 1506
rect 12070 1451 12190 1489
rect 12248 1489 12282 1506
rect 12334 1506 12350 1523
rect 12444 1523 12528 1539
rect 12444 1506 12460 1523
rect 12334 1489 12368 1506
rect 12248 1451 12368 1489
rect 12426 1489 12460 1506
rect 12512 1506 12528 1523
rect 12622 1523 12706 1539
rect 12622 1506 12638 1523
rect 12512 1489 12546 1506
rect 12426 1451 12546 1489
rect 12604 1489 12638 1506
rect 12690 1506 12706 1523
rect 12690 1489 12724 1506
rect 12604 1451 12724 1489
rect 474 1133 594 1171
rect 474 1117 508 1133
rect 492 1099 508 1117
rect 560 1117 594 1133
rect 652 1133 772 1171
rect 652 1117 686 1133
rect 560 1099 576 1117
rect 492 1083 576 1099
rect 670 1099 686 1117
rect 738 1117 772 1133
rect 830 1133 950 1171
rect 830 1117 864 1133
rect 738 1099 754 1117
rect 670 1083 754 1099
rect 848 1099 864 1117
rect 916 1117 950 1133
rect 1008 1133 1128 1171
rect 1008 1117 1042 1133
rect 916 1099 932 1117
rect 848 1083 932 1099
rect 1026 1099 1042 1117
rect 1094 1117 1128 1133
rect 1186 1133 1306 1171
rect 1186 1117 1220 1133
rect 1094 1099 1110 1117
rect 1026 1083 1110 1099
rect 1204 1099 1220 1117
rect 1272 1117 1306 1133
rect 1364 1133 1484 1171
rect 1364 1117 1398 1133
rect 1272 1099 1288 1117
rect 1204 1083 1288 1099
rect 1382 1099 1398 1117
rect 1450 1117 1484 1133
rect 1542 1133 1662 1171
rect 1542 1117 1576 1133
rect 1450 1099 1466 1117
rect 1382 1083 1466 1099
rect 1560 1099 1576 1117
rect 1628 1117 1662 1133
rect 1720 1133 1840 1171
rect 1720 1117 1754 1133
rect 1628 1099 1644 1117
rect 1560 1083 1644 1099
rect 1738 1099 1754 1117
rect 1806 1117 1840 1133
rect 1898 1133 2018 1171
rect 1898 1117 1932 1133
rect 1806 1099 1822 1117
rect 1738 1083 1822 1099
rect 1916 1099 1932 1117
rect 1984 1117 2018 1133
rect 2076 1133 2196 1171
rect 2076 1117 2110 1133
rect 1984 1099 2000 1117
rect 1916 1083 2000 1099
rect 2094 1099 2110 1117
rect 2162 1117 2196 1133
rect 2254 1133 2374 1171
rect 2254 1117 2288 1133
rect 2162 1099 2178 1117
rect 2094 1083 2178 1099
rect 2272 1099 2288 1117
rect 2340 1117 2374 1133
rect 2432 1133 2552 1171
rect 2432 1117 2466 1133
rect 2340 1099 2356 1117
rect 2272 1083 2356 1099
rect 2450 1099 2466 1117
rect 2518 1117 2552 1133
rect 2610 1133 2730 1171
rect 2610 1117 2644 1133
rect 2518 1099 2534 1117
rect 2450 1083 2534 1099
rect 2628 1099 2644 1117
rect 2696 1117 2730 1133
rect 2788 1133 2908 1171
rect 2788 1117 2822 1133
rect 2696 1099 2712 1117
rect 2628 1083 2712 1099
rect 2806 1099 2822 1117
rect 2874 1117 2908 1133
rect 2966 1133 3086 1171
rect 2966 1117 3000 1133
rect 2874 1099 2890 1117
rect 2806 1083 2890 1099
rect 2984 1099 3000 1117
rect 3052 1117 3086 1133
rect 3144 1133 3264 1171
rect 3144 1117 3178 1133
rect 3052 1099 3068 1117
rect 2984 1083 3068 1099
rect 3162 1099 3178 1117
rect 3230 1117 3264 1133
rect 3322 1133 3442 1171
rect 3322 1117 3356 1133
rect 3230 1099 3246 1117
rect 3162 1083 3246 1099
rect 3340 1099 3356 1117
rect 3408 1117 3442 1133
rect 3500 1133 3620 1171
rect 3500 1117 3534 1133
rect 3408 1099 3424 1117
rect 3340 1083 3424 1099
rect 3518 1099 3534 1117
rect 3586 1117 3620 1133
rect 3874 1133 3994 1171
rect 3874 1117 3908 1133
rect 3586 1099 3602 1117
rect 3518 1083 3602 1099
rect 3892 1099 3908 1117
rect 3960 1117 3994 1133
rect 4052 1133 4172 1171
rect 4052 1117 4086 1133
rect 3960 1099 3976 1117
rect 3892 1083 3976 1099
rect 4070 1099 4086 1117
rect 4138 1117 4172 1133
rect 4230 1133 4350 1171
rect 4230 1117 4264 1133
rect 4138 1099 4154 1117
rect 4070 1083 4154 1099
rect 4248 1099 4264 1117
rect 4316 1117 4350 1133
rect 4408 1133 4528 1171
rect 4408 1117 4442 1133
rect 4316 1099 4332 1117
rect 4248 1083 4332 1099
rect 4426 1099 4442 1117
rect 4494 1117 4528 1133
rect 4586 1133 4706 1171
rect 4586 1117 4620 1133
rect 4494 1099 4510 1117
rect 4426 1083 4510 1099
rect 4604 1099 4620 1117
rect 4672 1117 4706 1133
rect 4764 1133 4884 1171
rect 4764 1117 4798 1133
rect 4672 1099 4688 1117
rect 4604 1083 4688 1099
rect 4782 1099 4798 1117
rect 4850 1117 4884 1133
rect 4942 1133 5062 1171
rect 4942 1117 4976 1133
rect 4850 1099 4866 1117
rect 4782 1083 4866 1099
rect 4960 1099 4976 1117
rect 5028 1117 5062 1133
rect 5120 1133 5240 1171
rect 5120 1117 5154 1133
rect 5028 1099 5044 1117
rect 4960 1083 5044 1099
rect 5138 1099 5154 1117
rect 5206 1117 5240 1133
rect 5298 1133 5418 1171
rect 5298 1117 5332 1133
rect 5206 1099 5222 1117
rect 5138 1083 5222 1099
rect 5316 1099 5332 1117
rect 5384 1117 5418 1133
rect 5476 1133 5596 1171
rect 5476 1117 5510 1133
rect 5384 1099 5400 1117
rect 5316 1083 5400 1099
rect 5494 1099 5510 1117
rect 5562 1117 5596 1133
rect 5654 1133 5774 1171
rect 5654 1117 5688 1133
rect 5562 1099 5578 1117
rect 5494 1083 5578 1099
rect 5672 1099 5688 1117
rect 5740 1117 5774 1133
rect 5832 1133 5952 1171
rect 5832 1117 5866 1133
rect 5740 1099 5756 1117
rect 5672 1083 5756 1099
rect 5850 1099 5866 1117
rect 5918 1117 5952 1133
rect 6010 1133 6130 1171
rect 6010 1117 6044 1133
rect 5918 1099 5934 1117
rect 5850 1083 5934 1099
rect 6028 1099 6044 1117
rect 6096 1117 6130 1133
rect 6188 1133 6308 1171
rect 6188 1117 6222 1133
rect 6096 1099 6112 1117
rect 6028 1083 6112 1099
rect 6206 1099 6222 1117
rect 6274 1117 6308 1133
rect 6366 1133 6486 1171
rect 6366 1117 6400 1133
rect 6274 1099 6290 1117
rect 6206 1083 6290 1099
rect 6384 1099 6400 1117
rect 6452 1117 6486 1133
rect 6544 1133 6664 1171
rect 6544 1117 6578 1133
rect 6452 1099 6468 1117
rect 6384 1083 6468 1099
rect 6562 1099 6578 1117
rect 6630 1117 6664 1133
rect 6722 1133 6842 1171
rect 6722 1117 6756 1133
rect 6630 1099 6646 1117
rect 6562 1083 6646 1099
rect 6740 1099 6756 1117
rect 6808 1117 6842 1133
rect 6900 1133 7020 1171
rect 6900 1117 6934 1133
rect 6808 1099 6824 1117
rect 6740 1083 6824 1099
rect 6918 1099 6934 1117
rect 6986 1117 7020 1133
rect 7603 1133 7723 1171
rect 6986 1099 7002 1117
rect 7603 1116 7637 1133
rect 6918 1083 7002 1099
rect 7621 1099 7637 1116
rect 7689 1116 7723 1133
rect 7781 1133 7901 1171
rect 7781 1116 7815 1133
rect 7689 1099 7705 1116
rect 7621 1083 7705 1099
rect 7799 1099 7815 1116
rect 7867 1116 7901 1133
rect 7959 1133 8079 1171
rect 7959 1116 7993 1133
rect 7867 1099 7883 1116
rect 7799 1083 7883 1099
rect 7977 1099 7993 1116
rect 8045 1116 8079 1133
rect 8137 1133 8257 1171
rect 8137 1116 8171 1133
rect 8045 1099 8061 1116
rect 7977 1083 8061 1099
rect 8155 1099 8171 1116
rect 8223 1116 8257 1133
rect 8315 1133 8435 1171
rect 8315 1116 8349 1133
rect 8223 1099 8239 1116
rect 8155 1083 8239 1099
rect 8333 1099 8349 1116
rect 8401 1116 8435 1133
rect 8493 1133 8613 1171
rect 8493 1116 8527 1133
rect 8401 1099 8417 1116
rect 8333 1083 8417 1099
rect 8511 1099 8527 1116
rect 8579 1116 8613 1133
rect 8671 1133 8791 1171
rect 8671 1116 8705 1133
rect 8579 1099 8595 1116
rect 8511 1083 8595 1099
rect 8689 1099 8705 1116
rect 8757 1116 8791 1133
rect 8849 1133 8969 1171
rect 8849 1116 8883 1133
rect 8757 1099 8773 1116
rect 8689 1083 8773 1099
rect 8867 1099 8883 1116
rect 8935 1116 8969 1133
rect 9027 1133 9147 1171
rect 9027 1116 9061 1133
rect 8935 1099 8951 1116
rect 8867 1083 8951 1099
rect 9045 1099 9061 1116
rect 9113 1116 9147 1133
rect 9205 1133 9325 1171
rect 9205 1116 9239 1133
rect 9113 1099 9129 1116
rect 9045 1083 9129 1099
rect 9223 1099 9239 1116
rect 9291 1116 9325 1133
rect 9383 1133 9503 1171
rect 9383 1116 9417 1133
rect 9291 1099 9307 1116
rect 9223 1083 9307 1099
rect 9401 1099 9417 1116
rect 9469 1116 9503 1133
rect 9561 1133 9681 1171
rect 9561 1116 9595 1133
rect 9469 1099 9485 1116
rect 9401 1083 9485 1099
rect 9579 1099 9595 1116
rect 9647 1116 9681 1133
rect 9739 1133 9859 1171
rect 9739 1116 9773 1133
rect 9647 1099 9663 1116
rect 9579 1083 9663 1099
rect 9757 1099 9773 1116
rect 9825 1116 9859 1133
rect 9917 1133 10037 1171
rect 9917 1116 9951 1133
rect 9825 1099 9841 1116
rect 9757 1083 9841 1099
rect 9935 1099 9951 1116
rect 10003 1116 10037 1133
rect 10290 1133 10410 1171
rect 10290 1116 10324 1133
rect 10003 1099 10019 1116
rect 9935 1083 10019 1099
rect 10308 1099 10324 1116
rect 10376 1116 10410 1133
rect 10468 1133 10588 1171
rect 10468 1116 10502 1133
rect 10376 1099 10392 1116
rect 10308 1083 10392 1099
rect 10486 1099 10502 1116
rect 10554 1116 10588 1133
rect 10646 1133 10766 1171
rect 10646 1116 10680 1133
rect 10554 1099 10570 1116
rect 10486 1083 10570 1099
rect 10664 1099 10680 1116
rect 10732 1116 10766 1133
rect 10824 1133 10944 1171
rect 10824 1116 10858 1133
rect 10732 1099 10748 1116
rect 10664 1083 10748 1099
rect 10842 1099 10858 1116
rect 10910 1116 10944 1133
rect 11002 1133 11122 1171
rect 11002 1116 11036 1133
rect 10910 1099 10926 1116
rect 10842 1083 10926 1099
rect 11020 1099 11036 1116
rect 11088 1116 11122 1133
rect 11180 1133 11300 1171
rect 11180 1116 11214 1133
rect 11088 1099 11104 1116
rect 11020 1083 11104 1099
rect 11198 1099 11214 1116
rect 11266 1116 11300 1133
rect 11358 1133 11478 1171
rect 11358 1116 11392 1133
rect 11266 1099 11282 1116
rect 11198 1083 11282 1099
rect 11376 1099 11392 1116
rect 11444 1116 11478 1133
rect 11536 1133 11656 1171
rect 11536 1116 11570 1133
rect 11444 1099 11460 1116
rect 11376 1083 11460 1099
rect 11554 1099 11570 1116
rect 11622 1116 11656 1133
rect 11714 1133 11834 1171
rect 11714 1116 11748 1133
rect 11622 1099 11638 1116
rect 11554 1083 11638 1099
rect 11732 1099 11748 1116
rect 11800 1116 11834 1133
rect 11892 1133 12012 1171
rect 11892 1116 11926 1133
rect 11800 1099 11816 1116
rect 11732 1083 11816 1099
rect 11910 1099 11926 1116
rect 11978 1116 12012 1133
rect 12070 1133 12190 1171
rect 12070 1116 12104 1133
rect 11978 1099 11994 1116
rect 11910 1083 11994 1099
rect 12088 1099 12104 1116
rect 12156 1116 12190 1133
rect 12248 1133 12368 1171
rect 12248 1116 12282 1133
rect 12156 1099 12172 1116
rect 12088 1083 12172 1099
rect 12266 1099 12282 1116
rect 12334 1116 12368 1133
rect 12426 1133 12546 1171
rect 12426 1116 12460 1133
rect 12334 1099 12350 1116
rect 12266 1083 12350 1099
rect 12444 1099 12460 1116
rect 12512 1116 12546 1133
rect 12604 1133 12724 1171
rect 12604 1116 12638 1133
rect 12512 1099 12528 1116
rect 12444 1083 12528 1099
rect 12622 1099 12638 1116
rect 12690 1116 12724 1133
rect 12690 1099 12706 1116
rect 12622 1083 12706 1099
rect 492 1023 576 1039
rect 492 1005 508 1023
rect 474 989 508 1005
rect 560 1005 576 1023
rect 670 1023 754 1039
rect 670 1005 686 1023
rect 560 989 594 1005
rect 474 951 594 989
rect 652 989 686 1005
rect 738 1005 754 1023
rect 848 1023 932 1039
rect 848 1005 864 1023
rect 738 989 772 1005
rect 652 951 772 989
rect 830 989 864 1005
rect 916 1005 932 1023
rect 1026 1023 1110 1039
rect 1026 1005 1042 1023
rect 916 989 950 1005
rect 830 951 950 989
rect 1008 989 1042 1005
rect 1094 1005 1110 1023
rect 1204 1023 1288 1039
rect 1204 1005 1220 1023
rect 1094 989 1128 1005
rect 1008 951 1128 989
rect 1186 989 1220 1005
rect 1272 1005 1288 1023
rect 1382 1023 1466 1039
rect 1382 1005 1398 1023
rect 1272 989 1306 1005
rect 1186 951 1306 989
rect 1364 989 1398 1005
rect 1450 1005 1466 1023
rect 1560 1023 1644 1039
rect 1560 1005 1576 1023
rect 1450 989 1484 1005
rect 1364 951 1484 989
rect 1542 989 1576 1005
rect 1628 1005 1644 1023
rect 1738 1023 1822 1039
rect 1738 1005 1754 1023
rect 1628 989 1662 1005
rect 1542 951 1662 989
rect 1720 989 1754 1005
rect 1806 1005 1822 1023
rect 1916 1023 2000 1039
rect 1916 1005 1932 1023
rect 1806 989 1840 1005
rect 1720 951 1840 989
rect 1898 989 1932 1005
rect 1984 1005 2000 1023
rect 2094 1023 2178 1039
rect 2094 1005 2110 1023
rect 1984 989 2018 1005
rect 1898 951 2018 989
rect 2076 989 2110 1005
rect 2162 1005 2178 1023
rect 2272 1023 2356 1039
rect 2272 1005 2288 1023
rect 2162 989 2196 1005
rect 2076 951 2196 989
rect 2254 989 2288 1005
rect 2340 1005 2356 1023
rect 2450 1023 2534 1039
rect 2450 1005 2466 1023
rect 2340 989 2374 1005
rect 2254 951 2374 989
rect 2432 989 2466 1005
rect 2518 1005 2534 1023
rect 2628 1023 2712 1039
rect 2628 1005 2644 1023
rect 2518 989 2552 1005
rect 2432 951 2552 989
rect 2610 989 2644 1005
rect 2696 1005 2712 1023
rect 2806 1023 2890 1039
rect 2806 1005 2822 1023
rect 2696 989 2730 1005
rect 2610 951 2730 989
rect 2788 989 2822 1005
rect 2874 1005 2890 1023
rect 2984 1023 3068 1039
rect 2984 1005 3000 1023
rect 2874 989 2908 1005
rect 2788 951 2908 989
rect 2966 989 3000 1005
rect 3052 1005 3068 1023
rect 3162 1023 3246 1039
rect 3162 1005 3178 1023
rect 3052 989 3086 1005
rect 2966 951 3086 989
rect 3144 989 3178 1005
rect 3230 1005 3246 1023
rect 3340 1023 3424 1039
rect 3340 1005 3356 1023
rect 3230 989 3264 1005
rect 3144 951 3264 989
rect 3322 989 3356 1005
rect 3408 1005 3424 1023
rect 3518 1023 3602 1039
rect 3518 1005 3534 1023
rect 3408 989 3442 1005
rect 3322 951 3442 989
rect 3500 989 3534 1005
rect 3586 1005 3602 1023
rect 3892 1023 3976 1039
rect 3892 1005 3908 1023
rect 3586 989 3620 1005
rect 3500 951 3620 989
rect 3874 989 3908 1005
rect 3960 1005 3976 1023
rect 4070 1023 4154 1039
rect 4070 1005 4086 1023
rect 3960 989 3994 1005
rect 3874 951 3994 989
rect 4052 989 4086 1005
rect 4138 1005 4154 1023
rect 4248 1023 4332 1039
rect 4248 1005 4264 1023
rect 4138 989 4172 1005
rect 4052 951 4172 989
rect 4230 989 4264 1005
rect 4316 1005 4332 1023
rect 4426 1023 4510 1039
rect 4426 1005 4442 1023
rect 4316 989 4350 1005
rect 4230 951 4350 989
rect 4408 989 4442 1005
rect 4494 1005 4510 1023
rect 4604 1023 4688 1039
rect 4604 1005 4620 1023
rect 4494 989 4528 1005
rect 4408 951 4528 989
rect 4586 989 4620 1005
rect 4672 1005 4688 1023
rect 4782 1023 4866 1039
rect 4782 1005 4798 1023
rect 4672 989 4706 1005
rect 4586 951 4706 989
rect 4764 989 4798 1005
rect 4850 1005 4866 1023
rect 4960 1023 5044 1039
rect 4960 1005 4976 1023
rect 4850 989 4884 1005
rect 4764 951 4884 989
rect 4942 989 4976 1005
rect 5028 1005 5044 1023
rect 5138 1023 5222 1039
rect 5138 1005 5154 1023
rect 5028 989 5062 1005
rect 4942 951 5062 989
rect 5120 989 5154 1005
rect 5206 1005 5222 1023
rect 5316 1023 5400 1039
rect 5316 1005 5332 1023
rect 5206 989 5240 1005
rect 5120 951 5240 989
rect 5298 989 5332 1005
rect 5384 1005 5400 1023
rect 5494 1023 5578 1039
rect 5494 1005 5510 1023
rect 5384 989 5418 1005
rect 5298 951 5418 989
rect 5476 989 5510 1005
rect 5562 1005 5578 1023
rect 5672 1023 5756 1039
rect 5672 1005 5688 1023
rect 5562 989 5596 1005
rect 5476 951 5596 989
rect 5654 989 5688 1005
rect 5740 1005 5756 1023
rect 5850 1023 5934 1039
rect 5850 1005 5866 1023
rect 5740 989 5774 1005
rect 5654 951 5774 989
rect 5832 989 5866 1005
rect 5918 1005 5934 1023
rect 6028 1023 6112 1039
rect 6028 1005 6044 1023
rect 5918 989 5952 1005
rect 5832 951 5952 989
rect 6010 989 6044 1005
rect 6096 1005 6112 1023
rect 6206 1023 6290 1039
rect 6206 1005 6222 1023
rect 6096 989 6130 1005
rect 6010 951 6130 989
rect 6188 989 6222 1005
rect 6274 1005 6290 1023
rect 6384 1023 6468 1039
rect 6384 1005 6400 1023
rect 6274 989 6308 1005
rect 6188 951 6308 989
rect 6366 989 6400 1005
rect 6452 1005 6468 1023
rect 6562 1023 6646 1039
rect 6562 1005 6578 1023
rect 6452 989 6486 1005
rect 6366 951 6486 989
rect 6544 989 6578 1005
rect 6630 1005 6646 1023
rect 6740 1023 6824 1039
rect 6740 1005 6756 1023
rect 6630 989 6664 1005
rect 6544 951 6664 989
rect 6722 989 6756 1005
rect 6808 1005 6824 1023
rect 6918 1023 7002 1039
rect 6918 1005 6934 1023
rect 6808 989 6842 1005
rect 6722 951 6842 989
rect 6900 989 6934 1005
rect 6986 1005 7002 1023
rect 7621 1023 7705 1039
rect 7621 1006 7637 1023
rect 6986 989 7020 1005
rect 6900 951 7020 989
rect 7603 989 7637 1006
rect 7689 1006 7705 1023
rect 7799 1023 7883 1039
rect 7799 1006 7815 1023
rect 7689 989 7723 1006
rect 7603 951 7723 989
rect 7781 989 7815 1006
rect 7867 1006 7883 1023
rect 7977 1023 8061 1039
rect 7977 1006 7993 1023
rect 7867 989 7901 1006
rect 7781 951 7901 989
rect 7959 989 7993 1006
rect 8045 1006 8061 1023
rect 8155 1023 8239 1039
rect 8155 1006 8171 1023
rect 8045 989 8079 1006
rect 7959 951 8079 989
rect 8137 989 8171 1006
rect 8223 1006 8239 1023
rect 8333 1023 8417 1039
rect 8333 1006 8349 1023
rect 8223 989 8257 1006
rect 8137 951 8257 989
rect 8315 989 8349 1006
rect 8401 1006 8417 1023
rect 8511 1023 8595 1039
rect 8511 1006 8527 1023
rect 8401 989 8435 1006
rect 8315 951 8435 989
rect 8493 989 8527 1006
rect 8579 1006 8595 1023
rect 8689 1023 8773 1039
rect 8689 1006 8705 1023
rect 8579 989 8613 1006
rect 8493 951 8613 989
rect 8671 989 8705 1006
rect 8757 1006 8773 1023
rect 8867 1023 8951 1039
rect 8867 1006 8883 1023
rect 8757 989 8791 1006
rect 8671 951 8791 989
rect 8849 989 8883 1006
rect 8935 1006 8951 1023
rect 9045 1023 9129 1039
rect 9045 1006 9061 1023
rect 8935 989 8969 1006
rect 8849 951 8969 989
rect 9027 989 9061 1006
rect 9113 1006 9129 1023
rect 9223 1023 9307 1039
rect 9223 1006 9239 1023
rect 9113 989 9147 1006
rect 9027 951 9147 989
rect 9205 989 9239 1006
rect 9291 1006 9307 1023
rect 9401 1023 9485 1039
rect 9401 1006 9417 1023
rect 9291 989 9325 1006
rect 9205 951 9325 989
rect 9383 989 9417 1006
rect 9469 1006 9485 1023
rect 9579 1023 9663 1039
rect 9579 1006 9595 1023
rect 9469 989 9503 1006
rect 9383 951 9503 989
rect 9561 989 9595 1006
rect 9647 1006 9663 1023
rect 9757 1023 9841 1039
rect 9757 1006 9773 1023
rect 9647 989 9681 1006
rect 9561 951 9681 989
rect 9739 989 9773 1006
rect 9825 1006 9841 1023
rect 9935 1023 10019 1039
rect 9935 1006 9951 1023
rect 9825 989 9859 1006
rect 9739 951 9859 989
rect 9917 989 9951 1006
rect 10003 1006 10019 1023
rect 10308 1023 10392 1039
rect 10308 1006 10324 1023
rect 10003 989 10037 1006
rect 9917 951 10037 989
rect 10290 989 10324 1006
rect 10376 1006 10392 1023
rect 10486 1023 10570 1039
rect 10486 1006 10502 1023
rect 10376 989 10410 1006
rect 10290 951 10410 989
rect 10468 989 10502 1006
rect 10554 1006 10570 1023
rect 10664 1023 10748 1039
rect 10664 1006 10680 1023
rect 10554 989 10588 1006
rect 10468 951 10588 989
rect 10646 989 10680 1006
rect 10732 1006 10748 1023
rect 10842 1023 10926 1039
rect 10842 1006 10858 1023
rect 10732 989 10766 1006
rect 10646 951 10766 989
rect 10824 989 10858 1006
rect 10910 1006 10926 1023
rect 11020 1023 11104 1039
rect 11020 1006 11036 1023
rect 10910 989 10944 1006
rect 10824 951 10944 989
rect 11002 989 11036 1006
rect 11088 1006 11104 1023
rect 11198 1023 11282 1039
rect 11198 1006 11214 1023
rect 11088 989 11122 1006
rect 11002 951 11122 989
rect 11180 989 11214 1006
rect 11266 1006 11282 1023
rect 11376 1023 11460 1039
rect 11376 1006 11392 1023
rect 11266 989 11300 1006
rect 11180 951 11300 989
rect 11358 989 11392 1006
rect 11444 1006 11460 1023
rect 11554 1023 11638 1039
rect 11554 1006 11570 1023
rect 11444 989 11478 1006
rect 11358 951 11478 989
rect 11536 989 11570 1006
rect 11622 1006 11638 1023
rect 11732 1023 11816 1039
rect 11732 1006 11748 1023
rect 11622 989 11656 1006
rect 11536 951 11656 989
rect 11714 989 11748 1006
rect 11800 1006 11816 1023
rect 11910 1023 11994 1039
rect 11910 1006 11926 1023
rect 11800 989 11834 1006
rect 11714 951 11834 989
rect 11892 989 11926 1006
rect 11978 1006 11994 1023
rect 12088 1023 12172 1039
rect 12088 1006 12104 1023
rect 11978 989 12012 1006
rect 11892 951 12012 989
rect 12070 989 12104 1006
rect 12156 1006 12172 1023
rect 12266 1023 12350 1039
rect 12266 1006 12282 1023
rect 12156 989 12190 1006
rect 12070 951 12190 989
rect 12248 989 12282 1006
rect 12334 1006 12350 1023
rect 12444 1023 12528 1039
rect 12444 1006 12460 1023
rect 12334 989 12368 1006
rect 12248 951 12368 989
rect 12426 989 12460 1006
rect 12512 1006 12528 1023
rect 12622 1023 12706 1039
rect 12622 1006 12638 1023
rect 12512 989 12546 1006
rect 12426 951 12546 989
rect 12604 989 12638 1006
rect 12690 1006 12706 1023
rect 12690 989 12724 1006
rect 12604 951 12724 989
rect 474 633 594 671
rect 474 617 508 633
rect 492 599 508 617
rect 560 617 594 633
rect 652 633 772 671
rect 652 617 686 633
rect 560 599 576 617
rect 492 583 576 599
rect 670 599 686 617
rect 738 617 772 633
rect 830 633 950 671
rect 830 617 864 633
rect 738 599 754 617
rect 670 583 754 599
rect 848 599 864 617
rect 916 617 950 633
rect 1008 633 1128 671
rect 1008 617 1042 633
rect 916 599 932 617
rect 848 583 932 599
rect 1026 599 1042 617
rect 1094 617 1128 633
rect 1186 633 1306 671
rect 1186 617 1220 633
rect 1094 599 1110 617
rect 1026 583 1110 599
rect 1204 599 1220 617
rect 1272 617 1306 633
rect 1364 633 1484 671
rect 1364 617 1398 633
rect 1272 599 1288 617
rect 1204 583 1288 599
rect 1382 599 1398 617
rect 1450 617 1484 633
rect 1542 633 1662 671
rect 1542 617 1576 633
rect 1450 599 1466 617
rect 1382 583 1466 599
rect 1560 599 1576 617
rect 1628 617 1662 633
rect 1720 633 1840 671
rect 1720 617 1754 633
rect 1628 599 1644 617
rect 1560 583 1644 599
rect 1738 599 1754 617
rect 1806 617 1840 633
rect 1898 633 2018 671
rect 1898 617 1932 633
rect 1806 599 1822 617
rect 1738 583 1822 599
rect 1916 599 1932 617
rect 1984 617 2018 633
rect 2076 633 2196 671
rect 2076 617 2110 633
rect 1984 599 2000 617
rect 1916 583 2000 599
rect 2094 599 2110 617
rect 2162 617 2196 633
rect 2254 633 2374 671
rect 2254 617 2288 633
rect 2162 599 2178 617
rect 2094 583 2178 599
rect 2272 599 2288 617
rect 2340 617 2374 633
rect 2432 633 2552 671
rect 2432 617 2466 633
rect 2340 599 2356 617
rect 2272 583 2356 599
rect 2450 599 2466 617
rect 2518 617 2552 633
rect 2610 633 2730 671
rect 2610 617 2644 633
rect 2518 599 2534 617
rect 2450 583 2534 599
rect 2628 599 2644 617
rect 2696 617 2730 633
rect 2788 633 2908 671
rect 2788 617 2822 633
rect 2696 599 2712 617
rect 2628 583 2712 599
rect 2806 599 2822 617
rect 2874 617 2908 633
rect 2966 633 3086 671
rect 2966 617 3000 633
rect 2874 599 2890 617
rect 2806 583 2890 599
rect 2984 599 3000 617
rect 3052 617 3086 633
rect 3144 633 3264 671
rect 3144 617 3178 633
rect 3052 599 3068 617
rect 2984 583 3068 599
rect 3162 599 3178 617
rect 3230 617 3264 633
rect 3322 633 3442 671
rect 3322 617 3356 633
rect 3230 599 3246 617
rect 3162 583 3246 599
rect 3340 599 3356 617
rect 3408 617 3442 633
rect 3500 633 3620 671
rect 3500 617 3534 633
rect 3408 599 3424 617
rect 3340 583 3424 599
rect 3518 599 3534 617
rect 3586 617 3620 633
rect 3874 633 3994 671
rect 3874 617 3908 633
rect 3586 599 3602 617
rect 3518 583 3602 599
rect 3892 599 3908 617
rect 3960 617 3994 633
rect 4052 633 4172 671
rect 4052 617 4086 633
rect 3960 599 3976 617
rect 3892 583 3976 599
rect 4070 599 4086 617
rect 4138 617 4172 633
rect 4230 633 4350 671
rect 4230 617 4264 633
rect 4138 599 4154 617
rect 4070 583 4154 599
rect 4248 599 4264 617
rect 4316 617 4350 633
rect 4408 633 4528 671
rect 4408 617 4442 633
rect 4316 599 4332 617
rect 4248 583 4332 599
rect 4426 599 4442 617
rect 4494 617 4528 633
rect 4586 633 4706 671
rect 4586 617 4620 633
rect 4494 599 4510 617
rect 4426 583 4510 599
rect 4604 599 4620 617
rect 4672 617 4706 633
rect 4764 633 4884 671
rect 4764 617 4798 633
rect 4672 599 4688 617
rect 4604 583 4688 599
rect 4782 599 4798 617
rect 4850 617 4884 633
rect 4942 633 5062 671
rect 4942 617 4976 633
rect 4850 599 4866 617
rect 4782 583 4866 599
rect 4960 599 4976 617
rect 5028 617 5062 633
rect 5120 633 5240 671
rect 5120 617 5154 633
rect 5028 599 5044 617
rect 4960 583 5044 599
rect 5138 599 5154 617
rect 5206 617 5240 633
rect 5298 633 5418 671
rect 5298 617 5332 633
rect 5206 599 5222 617
rect 5138 583 5222 599
rect 5316 599 5332 617
rect 5384 617 5418 633
rect 5476 633 5596 671
rect 5476 617 5510 633
rect 5384 599 5400 617
rect 5316 583 5400 599
rect 5494 599 5510 617
rect 5562 617 5596 633
rect 5654 633 5774 671
rect 5654 617 5688 633
rect 5562 599 5578 617
rect 5494 583 5578 599
rect 5672 599 5688 617
rect 5740 617 5774 633
rect 5832 633 5952 671
rect 5832 617 5866 633
rect 5740 599 5756 617
rect 5672 583 5756 599
rect 5850 599 5866 617
rect 5918 617 5952 633
rect 6010 633 6130 671
rect 6010 617 6044 633
rect 5918 599 5934 617
rect 5850 583 5934 599
rect 6028 599 6044 617
rect 6096 617 6130 633
rect 6188 633 6308 671
rect 6188 617 6222 633
rect 6096 599 6112 617
rect 6028 583 6112 599
rect 6206 599 6222 617
rect 6274 617 6308 633
rect 6366 633 6486 671
rect 6366 617 6400 633
rect 6274 599 6290 617
rect 6206 583 6290 599
rect 6384 599 6400 617
rect 6452 617 6486 633
rect 6544 633 6664 671
rect 6544 617 6578 633
rect 6452 599 6468 617
rect 6384 583 6468 599
rect 6562 599 6578 617
rect 6630 617 6664 633
rect 6722 633 6842 671
rect 6722 617 6756 633
rect 6630 599 6646 617
rect 6562 583 6646 599
rect 6740 599 6756 617
rect 6808 617 6842 633
rect 6900 633 7020 671
rect 6900 617 6934 633
rect 6808 599 6824 617
rect 6740 583 6824 599
rect 6918 599 6934 617
rect 6986 617 7020 633
rect 7603 633 7723 671
rect 6986 599 7002 617
rect 7603 616 7637 633
rect 6918 583 7002 599
rect 7621 599 7637 616
rect 7689 616 7723 633
rect 7781 633 7901 671
rect 7781 616 7815 633
rect 7689 599 7705 616
rect 7621 583 7705 599
rect 7799 599 7815 616
rect 7867 616 7901 633
rect 7959 633 8079 671
rect 7959 616 7993 633
rect 7867 599 7883 616
rect 7799 583 7883 599
rect 7977 599 7993 616
rect 8045 616 8079 633
rect 8137 633 8257 671
rect 8137 616 8171 633
rect 8045 599 8061 616
rect 7977 583 8061 599
rect 8155 599 8171 616
rect 8223 616 8257 633
rect 8315 633 8435 671
rect 8315 616 8349 633
rect 8223 599 8239 616
rect 8155 583 8239 599
rect 8333 599 8349 616
rect 8401 616 8435 633
rect 8493 633 8613 671
rect 8493 616 8527 633
rect 8401 599 8417 616
rect 8333 583 8417 599
rect 8511 599 8527 616
rect 8579 616 8613 633
rect 8671 633 8791 671
rect 8671 616 8705 633
rect 8579 599 8595 616
rect 8511 583 8595 599
rect 8689 599 8705 616
rect 8757 616 8791 633
rect 8849 633 8969 671
rect 8849 616 8883 633
rect 8757 599 8773 616
rect 8689 583 8773 599
rect 8867 599 8883 616
rect 8935 616 8969 633
rect 9027 633 9147 671
rect 9027 616 9061 633
rect 8935 599 8951 616
rect 8867 583 8951 599
rect 9045 599 9061 616
rect 9113 616 9147 633
rect 9205 633 9325 671
rect 9205 616 9239 633
rect 9113 599 9129 616
rect 9045 583 9129 599
rect 9223 599 9239 616
rect 9291 616 9325 633
rect 9383 633 9503 671
rect 9383 616 9417 633
rect 9291 599 9307 616
rect 9223 583 9307 599
rect 9401 599 9417 616
rect 9469 616 9503 633
rect 9561 633 9681 671
rect 9561 616 9595 633
rect 9469 599 9485 616
rect 9401 583 9485 599
rect 9579 599 9595 616
rect 9647 616 9681 633
rect 9739 633 9859 671
rect 9739 616 9773 633
rect 9647 599 9663 616
rect 9579 583 9663 599
rect 9757 599 9773 616
rect 9825 616 9859 633
rect 9917 633 10037 671
rect 9917 616 9951 633
rect 9825 599 9841 616
rect 9757 583 9841 599
rect 9935 599 9951 616
rect 10003 616 10037 633
rect 10290 633 10410 671
rect 10290 616 10324 633
rect 10003 599 10019 616
rect 9935 583 10019 599
rect 10308 599 10324 616
rect 10376 616 10410 633
rect 10468 633 10588 671
rect 10468 616 10502 633
rect 10376 599 10392 616
rect 10308 583 10392 599
rect 10486 599 10502 616
rect 10554 616 10588 633
rect 10646 633 10766 671
rect 10646 616 10680 633
rect 10554 599 10570 616
rect 10486 583 10570 599
rect 10664 599 10680 616
rect 10732 616 10766 633
rect 10824 633 10944 671
rect 10824 616 10858 633
rect 10732 599 10748 616
rect 10664 583 10748 599
rect 10842 599 10858 616
rect 10910 616 10944 633
rect 11002 633 11122 671
rect 11002 616 11036 633
rect 10910 599 10926 616
rect 10842 583 10926 599
rect 11020 599 11036 616
rect 11088 616 11122 633
rect 11180 633 11300 671
rect 11180 616 11214 633
rect 11088 599 11104 616
rect 11020 583 11104 599
rect 11198 599 11214 616
rect 11266 616 11300 633
rect 11358 633 11478 671
rect 11358 616 11392 633
rect 11266 599 11282 616
rect 11198 583 11282 599
rect 11376 599 11392 616
rect 11444 616 11478 633
rect 11536 633 11656 671
rect 11536 616 11570 633
rect 11444 599 11460 616
rect 11376 583 11460 599
rect 11554 599 11570 616
rect 11622 616 11656 633
rect 11714 633 11834 671
rect 11714 616 11748 633
rect 11622 599 11638 616
rect 11554 583 11638 599
rect 11732 599 11748 616
rect 11800 616 11834 633
rect 11892 633 12012 671
rect 11892 616 11926 633
rect 11800 599 11816 616
rect 11732 583 11816 599
rect 11910 599 11926 616
rect 11978 616 12012 633
rect 12070 633 12190 671
rect 12070 616 12104 633
rect 11978 599 11994 616
rect 11910 583 11994 599
rect 12088 599 12104 616
rect 12156 616 12190 633
rect 12248 633 12368 671
rect 12248 616 12282 633
rect 12156 599 12172 616
rect 12088 583 12172 599
rect 12266 599 12282 616
rect 12334 616 12368 633
rect 12426 633 12546 671
rect 12426 616 12460 633
rect 12334 599 12350 616
rect 12266 583 12350 599
rect 12444 599 12460 616
rect 12512 616 12546 633
rect 12604 633 12724 671
rect 12604 616 12638 633
rect 12512 599 12528 616
rect 12444 583 12528 599
rect 12622 599 12638 616
rect 12690 616 12724 633
rect 12690 599 12706 616
rect 12622 583 12706 599
rect 13614 5131 13698 5147
rect 13614 5113 13630 5131
rect 13596 5097 13630 5113
rect 13682 5113 13698 5131
rect 13792 5131 13876 5147
rect 13792 5113 13808 5131
rect 13682 5097 13716 5113
rect 13596 5059 13716 5097
rect 13774 5097 13808 5113
rect 13860 5113 13876 5131
rect 13970 5131 14054 5147
rect 13970 5113 13986 5131
rect 13860 5097 13894 5113
rect 13774 5059 13894 5097
rect 13952 5097 13986 5113
rect 14038 5113 14054 5131
rect 14148 5131 14232 5147
rect 14148 5113 14164 5131
rect 14038 5097 14072 5113
rect 13952 5059 14072 5097
rect 14130 5097 14164 5113
rect 14216 5113 14232 5131
rect 14326 5131 14410 5147
rect 14326 5113 14342 5131
rect 14216 5097 14250 5113
rect 14130 5059 14250 5097
rect 14308 5097 14342 5113
rect 14394 5113 14410 5131
rect 14504 5131 14588 5147
rect 14504 5113 14520 5131
rect 14394 5097 14428 5113
rect 14308 5059 14428 5097
rect 14486 5097 14520 5113
rect 14572 5113 14588 5131
rect 14682 5131 14766 5147
rect 14682 5113 14698 5131
rect 14572 5097 14606 5113
rect 14486 5059 14606 5097
rect 14664 5097 14698 5113
rect 14750 5113 14766 5131
rect 14860 5131 14944 5147
rect 14860 5113 14876 5131
rect 14750 5097 14784 5113
rect 14664 5059 14784 5097
rect 14842 5097 14876 5113
rect 14928 5113 14944 5131
rect 15038 5131 15122 5147
rect 15038 5113 15054 5131
rect 14928 5097 14962 5113
rect 14842 5059 14962 5097
rect 15020 5097 15054 5113
rect 15106 5113 15122 5131
rect 15216 5131 15300 5147
rect 15216 5113 15232 5131
rect 15106 5097 15140 5113
rect 15020 5059 15140 5097
rect 15198 5097 15232 5113
rect 15284 5113 15300 5131
rect 15394 5131 15478 5147
rect 15394 5113 15410 5131
rect 15284 5097 15318 5113
rect 15198 5059 15318 5097
rect 15376 5097 15410 5113
rect 15462 5113 15478 5131
rect 15572 5131 15656 5147
rect 15572 5113 15588 5131
rect 15462 5097 15496 5113
rect 15376 5059 15496 5097
rect 15554 5097 15588 5113
rect 15640 5113 15656 5131
rect 15750 5131 15834 5147
rect 15750 5113 15766 5131
rect 15640 5097 15674 5113
rect 15554 5059 15674 5097
rect 15732 5097 15766 5113
rect 15818 5113 15834 5131
rect 15928 5131 16012 5147
rect 15928 5113 15944 5131
rect 15818 5097 15852 5113
rect 15732 5059 15852 5097
rect 15910 5097 15944 5113
rect 15996 5113 16012 5131
rect 16106 5131 16190 5147
rect 16106 5113 16122 5131
rect 15996 5097 16030 5113
rect 15910 5059 16030 5097
rect 16088 5097 16122 5113
rect 16174 5113 16190 5131
rect 16284 5131 16368 5147
rect 16284 5113 16300 5131
rect 16174 5097 16208 5113
rect 16088 5059 16208 5097
rect 16266 5097 16300 5113
rect 16352 5113 16368 5131
rect 16462 5131 16546 5147
rect 16462 5113 16478 5131
rect 16352 5097 16386 5113
rect 16266 5059 16386 5097
rect 16444 5097 16478 5113
rect 16530 5113 16546 5131
rect 16640 5131 16724 5147
rect 16640 5113 16656 5131
rect 16530 5097 16564 5113
rect 16444 5059 16564 5097
rect 16622 5097 16656 5113
rect 16708 5113 16724 5131
rect 16818 5131 16902 5147
rect 16818 5113 16834 5131
rect 16708 5097 16742 5113
rect 16622 5059 16742 5097
rect 16800 5097 16834 5113
rect 16886 5113 16902 5131
rect 16996 5131 17080 5147
rect 16996 5113 17012 5131
rect 16886 5097 16920 5113
rect 16800 5059 16920 5097
rect 16978 5097 17012 5113
rect 17064 5113 17080 5131
rect 17174 5131 17258 5147
rect 17174 5113 17190 5131
rect 17064 5097 17098 5113
rect 16978 5059 17098 5097
rect 17156 5097 17190 5113
rect 17242 5113 17258 5131
rect 17352 5131 17436 5147
rect 17352 5113 17368 5131
rect 17242 5097 17276 5113
rect 17156 5059 17276 5097
rect 17334 5097 17368 5113
rect 17420 5113 17436 5131
rect 17530 5131 17614 5147
rect 17530 5113 17546 5131
rect 17420 5097 17454 5113
rect 17334 5059 17454 5097
rect 17512 5097 17546 5113
rect 17598 5113 17614 5131
rect 17708 5131 17792 5147
rect 17708 5113 17724 5131
rect 17598 5097 17632 5113
rect 17512 5059 17632 5097
rect 17690 5097 17724 5113
rect 17776 5113 17792 5131
rect 17886 5131 17970 5147
rect 17886 5113 17902 5131
rect 17776 5097 17810 5113
rect 17690 5059 17810 5097
rect 17868 5097 17902 5113
rect 17954 5113 17970 5131
rect 18064 5131 18148 5147
rect 18064 5113 18080 5131
rect 17954 5097 17988 5113
rect 17868 5059 17988 5097
rect 18046 5097 18080 5113
rect 18132 5113 18148 5131
rect 18242 5131 18326 5147
rect 18242 5113 18258 5131
rect 18132 5097 18166 5113
rect 18046 5059 18166 5097
rect 18224 5097 18258 5113
rect 18310 5113 18326 5131
rect 18310 5097 18344 5113
rect 18224 5059 18344 5097
rect 13596 4741 13716 4779
rect 13596 4725 13630 4741
rect 13614 4707 13630 4725
rect 13682 4725 13716 4741
rect 13774 4741 13894 4779
rect 13774 4725 13808 4741
rect 13682 4707 13698 4725
rect 13614 4691 13698 4707
rect 13792 4707 13808 4725
rect 13860 4725 13894 4741
rect 13952 4741 14072 4779
rect 13952 4725 13986 4741
rect 13860 4707 13876 4725
rect 13792 4691 13876 4707
rect 13970 4707 13986 4725
rect 14038 4725 14072 4741
rect 14130 4741 14250 4779
rect 14130 4725 14164 4741
rect 14038 4707 14054 4725
rect 13970 4691 14054 4707
rect 14148 4707 14164 4725
rect 14216 4725 14250 4741
rect 14308 4741 14428 4779
rect 14308 4725 14342 4741
rect 14216 4707 14232 4725
rect 14148 4691 14232 4707
rect 14326 4707 14342 4725
rect 14394 4725 14428 4741
rect 14486 4741 14606 4779
rect 14486 4725 14520 4741
rect 14394 4707 14410 4725
rect 14326 4691 14410 4707
rect 14504 4707 14520 4725
rect 14572 4725 14606 4741
rect 14664 4741 14784 4779
rect 14664 4725 14698 4741
rect 14572 4707 14588 4725
rect 14504 4691 14588 4707
rect 14682 4707 14698 4725
rect 14750 4725 14784 4741
rect 14842 4741 14962 4779
rect 14842 4725 14876 4741
rect 14750 4707 14766 4725
rect 14682 4691 14766 4707
rect 14860 4707 14876 4725
rect 14928 4725 14962 4741
rect 15020 4741 15140 4779
rect 15020 4725 15054 4741
rect 14928 4707 14944 4725
rect 14860 4691 14944 4707
rect 15038 4707 15054 4725
rect 15106 4725 15140 4741
rect 15198 4741 15318 4779
rect 15198 4725 15232 4741
rect 15106 4707 15122 4725
rect 15038 4691 15122 4707
rect 15216 4707 15232 4725
rect 15284 4725 15318 4741
rect 15376 4741 15496 4779
rect 15376 4725 15410 4741
rect 15284 4707 15300 4725
rect 15216 4691 15300 4707
rect 15394 4707 15410 4725
rect 15462 4725 15496 4741
rect 15554 4741 15674 4779
rect 15554 4725 15588 4741
rect 15462 4707 15478 4725
rect 15394 4691 15478 4707
rect 15572 4707 15588 4725
rect 15640 4725 15674 4741
rect 15732 4741 15852 4779
rect 15732 4725 15766 4741
rect 15640 4707 15656 4725
rect 15572 4691 15656 4707
rect 15750 4707 15766 4725
rect 15818 4725 15852 4741
rect 15910 4741 16030 4779
rect 15910 4725 15944 4741
rect 15818 4707 15834 4725
rect 15750 4691 15834 4707
rect 15928 4707 15944 4725
rect 15996 4725 16030 4741
rect 16088 4741 16208 4779
rect 16088 4725 16122 4741
rect 15996 4707 16012 4725
rect 15928 4691 16012 4707
rect 16106 4707 16122 4725
rect 16174 4725 16208 4741
rect 16266 4741 16386 4779
rect 16266 4725 16300 4741
rect 16174 4707 16190 4725
rect 16106 4691 16190 4707
rect 16284 4707 16300 4725
rect 16352 4725 16386 4741
rect 16444 4741 16564 4779
rect 16444 4725 16478 4741
rect 16352 4707 16368 4725
rect 16284 4691 16368 4707
rect 16462 4707 16478 4725
rect 16530 4725 16564 4741
rect 16622 4741 16742 4779
rect 16622 4725 16656 4741
rect 16530 4707 16546 4725
rect 16462 4691 16546 4707
rect 16640 4707 16656 4725
rect 16708 4725 16742 4741
rect 16800 4741 16920 4779
rect 16800 4725 16834 4741
rect 16708 4707 16724 4725
rect 16640 4691 16724 4707
rect 16818 4707 16834 4725
rect 16886 4725 16920 4741
rect 16978 4741 17098 4779
rect 16978 4725 17012 4741
rect 16886 4707 16902 4725
rect 16818 4691 16902 4707
rect 16996 4707 17012 4725
rect 17064 4725 17098 4741
rect 17156 4741 17276 4779
rect 17156 4725 17190 4741
rect 17064 4707 17080 4725
rect 16996 4691 17080 4707
rect 17174 4707 17190 4725
rect 17242 4725 17276 4741
rect 17334 4741 17454 4779
rect 17334 4725 17368 4741
rect 17242 4707 17258 4725
rect 17174 4691 17258 4707
rect 17352 4707 17368 4725
rect 17420 4725 17454 4741
rect 17512 4741 17632 4779
rect 17512 4725 17546 4741
rect 17420 4707 17436 4725
rect 17352 4691 17436 4707
rect 17530 4707 17546 4725
rect 17598 4725 17632 4741
rect 17690 4741 17810 4779
rect 17690 4725 17724 4741
rect 17598 4707 17614 4725
rect 17530 4691 17614 4707
rect 17708 4707 17724 4725
rect 17776 4725 17810 4741
rect 17868 4741 17988 4779
rect 17868 4725 17902 4741
rect 17776 4707 17792 4725
rect 17708 4691 17792 4707
rect 17886 4707 17902 4725
rect 17954 4725 17988 4741
rect 18046 4741 18166 4779
rect 18046 4725 18080 4741
rect 17954 4707 17970 4725
rect 17886 4691 17970 4707
rect 18064 4707 18080 4725
rect 18132 4725 18166 4741
rect 18224 4741 18344 4779
rect 18224 4725 18258 4741
rect 18132 4707 18148 4725
rect 18064 4691 18148 4707
rect 18242 4707 18258 4725
rect 18310 4725 18344 4741
rect 18310 4707 18326 4725
rect 18242 4691 18326 4707
rect 13614 4631 13698 4647
rect 13614 4613 13630 4631
rect 13596 4597 13630 4613
rect 13682 4613 13698 4631
rect 13792 4631 13876 4647
rect 13792 4613 13808 4631
rect 13682 4597 13716 4613
rect 13596 4559 13716 4597
rect 13774 4597 13808 4613
rect 13860 4613 13876 4631
rect 13970 4631 14054 4647
rect 13970 4613 13986 4631
rect 13860 4597 13894 4613
rect 13774 4559 13894 4597
rect 13952 4597 13986 4613
rect 14038 4613 14054 4631
rect 14148 4631 14232 4647
rect 14148 4613 14164 4631
rect 14038 4597 14072 4613
rect 13952 4559 14072 4597
rect 14130 4597 14164 4613
rect 14216 4613 14232 4631
rect 14326 4631 14410 4647
rect 14326 4613 14342 4631
rect 14216 4597 14250 4613
rect 14130 4559 14250 4597
rect 14308 4597 14342 4613
rect 14394 4613 14410 4631
rect 14504 4631 14588 4647
rect 14504 4613 14520 4631
rect 14394 4597 14428 4613
rect 14308 4559 14428 4597
rect 14486 4597 14520 4613
rect 14572 4613 14588 4631
rect 14682 4631 14766 4647
rect 14682 4613 14698 4631
rect 14572 4597 14606 4613
rect 14486 4559 14606 4597
rect 14664 4597 14698 4613
rect 14750 4613 14766 4631
rect 14860 4631 14944 4647
rect 14860 4613 14876 4631
rect 14750 4597 14784 4613
rect 14664 4559 14784 4597
rect 14842 4597 14876 4613
rect 14928 4613 14944 4631
rect 15038 4631 15122 4647
rect 15038 4613 15054 4631
rect 14928 4597 14962 4613
rect 14842 4559 14962 4597
rect 15020 4597 15054 4613
rect 15106 4613 15122 4631
rect 15216 4631 15300 4647
rect 15216 4613 15232 4631
rect 15106 4597 15140 4613
rect 15020 4559 15140 4597
rect 15198 4597 15232 4613
rect 15284 4613 15300 4631
rect 15394 4631 15478 4647
rect 15394 4613 15410 4631
rect 15284 4597 15318 4613
rect 15198 4559 15318 4597
rect 15376 4597 15410 4613
rect 15462 4613 15478 4631
rect 15572 4631 15656 4647
rect 15572 4613 15588 4631
rect 15462 4597 15496 4613
rect 15376 4559 15496 4597
rect 15554 4597 15588 4613
rect 15640 4613 15656 4631
rect 15750 4631 15834 4647
rect 15750 4613 15766 4631
rect 15640 4597 15674 4613
rect 15554 4559 15674 4597
rect 15732 4597 15766 4613
rect 15818 4613 15834 4631
rect 15928 4631 16012 4647
rect 15928 4613 15944 4631
rect 15818 4597 15852 4613
rect 15732 4559 15852 4597
rect 15910 4597 15944 4613
rect 15996 4613 16012 4631
rect 16106 4631 16190 4647
rect 16106 4613 16122 4631
rect 15996 4597 16030 4613
rect 15910 4559 16030 4597
rect 16088 4597 16122 4613
rect 16174 4613 16190 4631
rect 16284 4631 16368 4647
rect 16284 4613 16300 4631
rect 16174 4597 16208 4613
rect 16088 4559 16208 4597
rect 16266 4597 16300 4613
rect 16352 4613 16368 4631
rect 16462 4631 16546 4647
rect 16462 4613 16478 4631
rect 16352 4597 16386 4613
rect 16266 4559 16386 4597
rect 16444 4597 16478 4613
rect 16530 4613 16546 4631
rect 16640 4631 16724 4647
rect 16640 4613 16656 4631
rect 16530 4597 16564 4613
rect 16444 4559 16564 4597
rect 16622 4597 16656 4613
rect 16708 4613 16724 4631
rect 16818 4631 16902 4647
rect 16818 4613 16834 4631
rect 16708 4597 16742 4613
rect 16622 4559 16742 4597
rect 16800 4597 16834 4613
rect 16886 4613 16902 4631
rect 16996 4631 17080 4647
rect 16996 4613 17012 4631
rect 16886 4597 16920 4613
rect 16800 4559 16920 4597
rect 16978 4597 17012 4613
rect 17064 4613 17080 4631
rect 17174 4631 17258 4647
rect 17174 4613 17190 4631
rect 17064 4597 17098 4613
rect 16978 4559 17098 4597
rect 17156 4597 17190 4613
rect 17242 4613 17258 4631
rect 17352 4631 17436 4647
rect 17352 4613 17368 4631
rect 17242 4597 17276 4613
rect 17156 4559 17276 4597
rect 17334 4597 17368 4613
rect 17420 4613 17436 4631
rect 17530 4631 17614 4647
rect 17530 4613 17546 4631
rect 17420 4597 17454 4613
rect 17334 4559 17454 4597
rect 17512 4597 17546 4613
rect 17598 4613 17614 4631
rect 17708 4631 17792 4647
rect 17708 4613 17724 4631
rect 17598 4597 17632 4613
rect 17512 4559 17632 4597
rect 17690 4597 17724 4613
rect 17776 4613 17792 4631
rect 17886 4631 17970 4647
rect 17886 4613 17902 4631
rect 17776 4597 17810 4613
rect 17690 4559 17810 4597
rect 17868 4597 17902 4613
rect 17954 4613 17970 4631
rect 18064 4631 18148 4647
rect 18064 4613 18080 4631
rect 17954 4597 17988 4613
rect 17868 4559 17988 4597
rect 18046 4597 18080 4613
rect 18132 4613 18148 4631
rect 18242 4631 18326 4647
rect 18242 4613 18258 4631
rect 18132 4597 18166 4613
rect 18046 4559 18166 4597
rect 18224 4597 18258 4613
rect 18310 4613 18326 4631
rect 18310 4597 18344 4613
rect 18224 4559 18344 4597
rect 13596 4241 13716 4279
rect 13596 4225 13630 4241
rect 13614 4207 13630 4225
rect 13682 4225 13716 4241
rect 13774 4241 13894 4279
rect 13774 4225 13808 4241
rect 13682 4207 13698 4225
rect 13614 4191 13698 4207
rect 13792 4207 13808 4225
rect 13860 4225 13894 4241
rect 13952 4241 14072 4279
rect 13952 4225 13986 4241
rect 13860 4207 13876 4225
rect 13792 4191 13876 4207
rect 13970 4207 13986 4225
rect 14038 4225 14072 4241
rect 14130 4241 14250 4279
rect 14130 4225 14164 4241
rect 14038 4207 14054 4225
rect 13970 4191 14054 4207
rect 14148 4207 14164 4225
rect 14216 4225 14250 4241
rect 14308 4241 14428 4279
rect 14308 4225 14342 4241
rect 14216 4207 14232 4225
rect 14148 4191 14232 4207
rect 14326 4207 14342 4225
rect 14394 4225 14428 4241
rect 14486 4241 14606 4279
rect 14486 4225 14520 4241
rect 14394 4207 14410 4225
rect 14326 4191 14410 4207
rect 14504 4207 14520 4225
rect 14572 4225 14606 4241
rect 14664 4241 14784 4279
rect 14664 4225 14698 4241
rect 14572 4207 14588 4225
rect 14504 4191 14588 4207
rect 14682 4207 14698 4225
rect 14750 4225 14784 4241
rect 14842 4241 14962 4279
rect 14842 4225 14876 4241
rect 14750 4207 14766 4225
rect 14682 4191 14766 4207
rect 14860 4207 14876 4225
rect 14928 4225 14962 4241
rect 15020 4241 15140 4279
rect 15020 4225 15054 4241
rect 14928 4207 14944 4225
rect 14860 4191 14944 4207
rect 15038 4207 15054 4225
rect 15106 4225 15140 4241
rect 15198 4241 15318 4279
rect 15198 4225 15232 4241
rect 15106 4207 15122 4225
rect 15038 4191 15122 4207
rect 15216 4207 15232 4225
rect 15284 4225 15318 4241
rect 15376 4241 15496 4279
rect 15376 4225 15410 4241
rect 15284 4207 15300 4225
rect 15216 4191 15300 4207
rect 15394 4207 15410 4225
rect 15462 4225 15496 4241
rect 15554 4241 15674 4279
rect 15554 4225 15588 4241
rect 15462 4207 15478 4225
rect 15394 4191 15478 4207
rect 15572 4207 15588 4225
rect 15640 4225 15674 4241
rect 15732 4241 15852 4279
rect 15732 4225 15766 4241
rect 15640 4207 15656 4225
rect 15572 4191 15656 4207
rect 15750 4207 15766 4225
rect 15818 4225 15852 4241
rect 15910 4241 16030 4279
rect 15910 4225 15944 4241
rect 15818 4207 15834 4225
rect 15750 4191 15834 4207
rect 15928 4207 15944 4225
rect 15996 4225 16030 4241
rect 16088 4241 16208 4279
rect 16088 4225 16122 4241
rect 15996 4207 16012 4225
rect 15928 4191 16012 4207
rect 16106 4207 16122 4225
rect 16174 4225 16208 4241
rect 16266 4241 16386 4279
rect 16266 4225 16300 4241
rect 16174 4207 16190 4225
rect 16106 4191 16190 4207
rect 16284 4207 16300 4225
rect 16352 4225 16386 4241
rect 16444 4241 16564 4279
rect 16444 4225 16478 4241
rect 16352 4207 16368 4225
rect 16284 4191 16368 4207
rect 16462 4207 16478 4225
rect 16530 4225 16564 4241
rect 16622 4241 16742 4279
rect 16622 4225 16656 4241
rect 16530 4207 16546 4225
rect 16462 4191 16546 4207
rect 16640 4207 16656 4225
rect 16708 4225 16742 4241
rect 16800 4241 16920 4279
rect 16800 4225 16834 4241
rect 16708 4207 16724 4225
rect 16640 4191 16724 4207
rect 16818 4207 16834 4225
rect 16886 4225 16920 4241
rect 16978 4241 17098 4279
rect 16978 4225 17012 4241
rect 16886 4207 16902 4225
rect 16818 4191 16902 4207
rect 16996 4207 17012 4225
rect 17064 4225 17098 4241
rect 17156 4241 17276 4279
rect 17156 4225 17190 4241
rect 17064 4207 17080 4225
rect 16996 4191 17080 4207
rect 17174 4207 17190 4225
rect 17242 4225 17276 4241
rect 17334 4241 17454 4279
rect 17334 4225 17368 4241
rect 17242 4207 17258 4225
rect 17174 4191 17258 4207
rect 17352 4207 17368 4225
rect 17420 4225 17454 4241
rect 17512 4241 17632 4279
rect 17512 4225 17546 4241
rect 17420 4207 17436 4225
rect 17352 4191 17436 4207
rect 17530 4207 17546 4225
rect 17598 4225 17632 4241
rect 17690 4241 17810 4279
rect 17690 4225 17724 4241
rect 17598 4207 17614 4225
rect 17530 4191 17614 4207
rect 17708 4207 17724 4225
rect 17776 4225 17810 4241
rect 17868 4241 17988 4279
rect 17868 4225 17902 4241
rect 17776 4207 17792 4225
rect 17708 4191 17792 4207
rect 17886 4207 17902 4225
rect 17954 4225 17988 4241
rect 18046 4241 18166 4279
rect 18046 4225 18080 4241
rect 17954 4207 17970 4225
rect 17886 4191 17970 4207
rect 18064 4207 18080 4225
rect 18132 4225 18166 4241
rect 18224 4241 18344 4279
rect 18224 4225 18258 4241
rect 18132 4207 18148 4225
rect 18064 4191 18148 4207
rect 18242 4207 18258 4225
rect 18310 4225 18344 4241
rect 18310 4207 18326 4225
rect 18242 4191 18326 4207
rect 17172 3627 17256 3643
rect 17172 3610 17188 3627
rect 17154 3593 17188 3610
rect 17240 3610 17256 3627
rect 17350 3627 17434 3643
rect 17350 3610 17366 3627
rect 17240 3593 17274 3610
rect 17154 3555 17274 3593
rect 17332 3593 17366 3610
rect 17418 3610 17434 3627
rect 17528 3627 17612 3643
rect 17528 3610 17544 3627
rect 17418 3593 17452 3610
rect 17332 3555 17452 3593
rect 17510 3593 17544 3610
rect 17596 3610 17612 3627
rect 17706 3627 17790 3643
rect 17706 3610 17722 3627
rect 17596 3593 17630 3610
rect 17510 3555 17630 3593
rect 17688 3593 17722 3610
rect 17774 3610 17790 3627
rect 17774 3593 17808 3610
rect 17688 3555 17808 3593
rect 17154 3237 17274 3275
rect 17154 3220 17188 3237
rect 17172 3203 17188 3220
rect 17240 3220 17274 3237
rect 17332 3237 17452 3275
rect 17332 3220 17366 3237
rect 17240 3203 17256 3220
rect 17172 3187 17256 3203
rect 17350 3203 17366 3220
rect 17418 3220 17452 3237
rect 17510 3237 17630 3275
rect 17510 3220 17544 3237
rect 17418 3203 17434 3220
rect 17350 3187 17434 3203
rect 17528 3203 17544 3220
rect 17596 3220 17630 3237
rect 17688 3237 17808 3275
rect 17688 3220 17722 3237
rect 17596 3203 17612 3220
rect 17528 3187 17612 3203
rect 17706 3203 17722 3220
rect 17774 3220 17808 3237
rect 17774 3203 17790 3220
rect 17706 3187 17790 3203
rect 16458 2688 16542 2704
rect 16458 2671 16474 2688
rect 16440 2654 16474 2671
rect 16526 2671 16542 2688
rect 16636 2688 16720 2704
rect 16636 2671 16652 2688
rect 16526 2654 16560 2671
rect 13740 2622 13824 2638
rect 13740 2606 13756 2622
rect 13722 2588 13756 2606
rect 13808 2606 13824 2622
rect 14032 2622 14116 2638
rect 14032 2606 14048 2622
rect 13808 2588 13842 2606
rect 13722 2550 13842 2588
rect 14014 2588 14048 2606
rect 14100 2606 14116 2622
rect 14324 2622 14408 2638
rect 14324 2606 14340 2622
rect 14100 2588 14134 2606
rect 14014 2550 14134 2588
rect 14306 2588 14340 2606
rect 14392 2606 14408 2622
rect 14616 2622 14700 2638
rect 14616 2606 14632 2622
rect 14392 2588 14426 2606
rect 14306 2550 14426 2588
rect 14598 2588 14632 2606
rect 14684 2606 14700 2622
rect 14908 2622 14992 2638
rect 14908 2606 14924 2622
rect 14684 2588 14718 2606
rect 14598 2550 14718 2588
rect 14890 2588 14924 2606
rect 14976 2606 14992 2622
rect 15200 2622 15284 2638
rect 15200 2606 15216 2622
rect 14976 2588 15010 2606
rect 14890 2550 15010 2588
rect 15182 2588 15216 2606
rect 15268 2606 15284 2622
rect 15492 2622 15576 2638
rect 15492 2606 15508 2622
rect 15268 2588 15302 2606
rect 15182 2550 15302 2588
rect 15474 2588 15508 2606
rect 15560 2606 15576 2622
rect 16440 2616 16560 2654
rect 16618 2654 16652 2671
rect 16704 2671 16720 2688
rect 16814 2688 16898 2704
rect 16814 2671 16830 2688
rect 16704 2654 16738 2671
rect 16618 2616 16738 2654
rect 16796 2654 16830 2671
rect 16882 2671 16898 2688
rect 16992 2688 17076 2704
rect 16992 2671 17008 2688
rect 16882 2654 16916 2671
rect 16796 2616 16916 2654
rect 16974 2654 17008 2671
rect 17060 2671 17076 2688
rect 17170 2688 17254 2704
rect 17170 2671 17186 2688
rect 17060 2654 17094 2671
rect 16974 2616 17094 2654
rect 17152 2654 17186 2671
rect 17238 2671 17254 2688
rect 17348 2688 17432 2704
rect 17348 2671 17364 2688
rect 17238 2654 17272 2671
rect 17152 2616 17272 2654
rect 17330 2654 17364 2671
rect 17416 2671 17432 2688
rect 17526 2688 17610 2704
rect 17526 2671 17542 2688
rect 17416 2654 17450 2671
rect 17330 2616 17450 2654
rect 17508 2654 17542 2671
rect 17594 2671 17610 2688
rect 17704 2688 17788 2704
rect 17704 2671 17720 2688
rect 17594 2654 17628 2671
rect 17508 2616 17628 2654
rect 17686 2654 17720 2671
rect 17772 2671 17788 2688
rect 17882 2688 17966 2704
rect 17882 2671 17898 2688
rect 17772 2654 17806 2671
rect 17686 2616 17806 2654
rect 17864 2654 17898 2671
rect 17950 2671 17966 2688
rect 18060 2688 18144 2704
rect 18060 2671 18076 2688
rect 17950 2654 17984 2671
rect 17864 2616 17984 2654
rect 18042 2654 18076 2671
rect 18128 2671 18144 2688
rect 18238 2688 18322 2704
rect 18238 2671 18254 2688
rect 18128 2654 18162 2671
rect 18042 2616 18162 2654
rect 18220 2654 18254 2671
rect 18306 2671 18322 2688
rect 18306 2654 18340 2671
rect 18220 2616 18340 2654
rect 15560 2588 15594 2606
rect 15474 2550 15594 2588
rect 16440 2298 16560 2336
rect 16440 2281 16474 2298
rect 13722 2232 13842 2270
rect 13722 2216 13756 2232
rect 13740 2198 13756 2216
rect 13808 2216 13842 2232
rect 14014 2232 14134 2270
rect 14014 2216 14048 2232
rect 13808 2198 13824 2216
rect 13740 2182 13824 2198
rect 14032 2198 14048 2216
rect 14100 2216 14134 2232
rect 14306 2232 14426 2270
rect 14306 2216 14340 2232
rect 14100 2198 14116 2216
rect 14032 2182 14116 2198
rect 14324 2198 14340 2216
rect 14392 2216 14426 2232
rect 14598 2232 14718 2270
rect 14598 2216 14632 2232
rect 14392 2198 14408 2216
rect 14324 2182 14408 2198
rect 14616 2198 14632 2216
rect 14684 2216 14718 2232
rect 14890 2232 15010 2270
rect 14890 2216 14924 2232
rect 14684 2198 14700 2216
rect 14616 2182 14700 2198
rect 14908 2198 14924 2216
rect 14976 2216 15010 2232
rect 15182 2232 15302 2270
rect 15182 2216 15216 2232
rect 14976 2198 14992 2216
rect 14908 2182 14992 2198
rect 15200 2198 15216 2216
rect 15268 2216 15302 2232
rect 15474 2232 15594 2270
rect 16458 2264 16474 2281
rect 16526 2281 16560 2298
rect 16618 2298 16738 2336
rect 16618 2281 16652 2298
rect 16526 2264 16542 2281
rect 16458 2248 16542 2264
rect 16636 2264 16652 2281
rect 16704 2281 16738 2298
rect 16796 2298 16916 2336
rect 16796 2281 16830 2298
rect 16704 2264 16720 2281
rect 16636 2248 16720 2264
rect 16814 2264 16830 2281
rect 16882 2281 16916 2298
rect 16974 2298 17094 2336
rect 16974 2281 17008 2298
rect 16882 2264 16898 2281
rect 16814 2248 16898 2264
rect 16992 2264 17008 2281
rect 17060 2281 17094 2298
rect 17152 2298 17272 2336
rect 17152 2281 17186 2298
rect 17060 2264 17076 2281
rect 16992 2248 17076 2264
rect 17170 2264 17186 2281
rect 17238 2281 17272 2298
rect 17330 2298 17450 2336
rect 17330 2281 17364 2298
rect 17238 2264 17254 2281
rect 17170 2248 17254 2264
rect 17348 2264 17364 2281
rect 17416 2281 17450 2298
rect 17508 2298 17628 2336
rect 17508 2281 17542 2298
rect 17416 2264 17432 2281
rect 17348 2248 17432 2264
rect 17526 2264 17542 2281
rect 17594 2281 17628 2298
rect 17686 2298 17806 2336
rect 17686 2281 17720 2298
rect 17594 2264 17610 2281
rect 17526 2248 17610 2264
rect 17704 2264 17720 2281
rect 17772 2281 17806 2298
rect 17864 2298 17984 2336
rect 17864 2281 17898 2298
rect 17772 2264 17788 2281
rect 17704 2248 17788 2264
rect 17882 2264 17898 2281
rect 17950 2281 17984 2298
rect 18042 2298 18162 2336
rect 18042 2281 18076 2298
rect 17950 2264 17966 2281
rect 17882 2248 17966 2264
rect 18060 2264 18076 2281
rect 18128 2281 18162 2298
rect 18220 2298 18340 2336
rect 18220 2281 18254 2298
rect 18128 2264 18144 2281
rect 18060 2248 18144 2264
rect 18238 2264 18254 2281
rect 18306 2281 18340 2298
rect 18306 2264 18322 2281
rect 18238 2248 18322 2264
rect 15474 2216 15508 2232
rect 15268 2198 15284 2216
rect 15200 2182 15284 2198
rect 15492 2198 15508 2216
rect 15560 2216 15594 2232
rect 15560 2198 15576 2216
rect 15492 2182 15576 2198
rect 16458 2188 16542 2204
rect 16458 2171 16474 2188
rect 16440 2154 16474 2171
rect 16526 2171 16542 2188
rect 16636 2188 16720 2204
rect 16636 2171 16652 2188
rect 16526 2154 16560 2171
rect 13740 2124 13824 2140
rect 13740 2108 13756 2124
rect 13722 2090 13756 2108
rect 13808 2108 13824 2124
rect 14032 2124 14116 2140
rect 14032 2108 14048 2124
rect 13808 2090 13842 2108
rect 13722 2052 13842 2090
rect 14014 2090 14048 2108
rect 14100 2108 14116 2124
rect 14324 2124 14408 2140
rect 14324 2108 14340 2124
rect 14100 2090 14134 2108
rect 14014 2052 14134 2090
rect 14306 2090 14340 2108
rect 14392 2108 14408 2124
rect 14616 2124 14700 2140
rect 14616 2108 14632 2124
rect 14392 2090 14426 2108
rect 14306 2052 14426 2090
rect 14598 2090 14632 2108
rect 14684 2108 14700 2124
rect 14908 2124 14992 2140
rect 14908 2108 14924 2124
rect 14684 2090 14718 2108
rect 14598 2052 14718 2090
rect 14890 2090 14924 2108
rect 14976 2108 14992 2124
rect 15200 2124 15284 2140
rect 15200 2108 15216 2124
rect 14976 2090 15010 2108
rect 14890 2052 15010 2090
rect 15182 2090 15216 2108
rect 15268 2108 15284 2124
rect 15492 2124 15576 2140
rect 15492 2108 15508 2124
rect 15268 2090 15302 2108
rect 15182 2052 15302 2090
rect 15474 2090 15508 2108
rect 15560 2108 15576 2124
rect 16440 2116 16560 2154
rect 16618 2154 16652 2171
rect 16704 2171 16720 2188
rect 16814 2188 16898 2204
rect 16814 2171 16830 2188
rect 16704 2154 16738 2171
rect 16618 2116 16738 2154
rect 16796 2154 16830 2171
rect 16882 2171 16898 2188
rect 16992 2188 17076 2204
rect 16992 2171 17008 2188
rect 16882 2154 16916 2171
rect 16796 2116 16916 2154
rect 16974 2154 17008 2171
rect 17060 2171 17076 2188
rect 17170 2188 17254 2204
rect 17170 2171 17186 2188
rect 17060 2154 17094 2171
rect 16974 2116 17094 2154
rect 17152 2154 17186 2171
rect 17238 2171 17254 2188
rect 17348 2188 17432 2204
rect 17348 2171 17364 2188
rect 17238 2154 17272 2171
rect 17152 2116 17272 2154
rect 17330 2154 17364 2171
rect 17416 2171 17432 2188
rect 17526 2188 17610 2204
rect 17526 2171 17542 2188
rect 17416 2154 17450 2171
rect 17330 2116 17450 2154
rect 17508 2154 17542 2171
rect 17594 2171 17610 2188
rect 17704 2188 17788 2204
rect 17704 2171 17720 2188
rect 17594 2154 17628 2171
rect 17508 2116 17628 2154
rect 17686 2154 17720 2171
rect 17772 2171 17788 2188
rect 17882 2188 17966 2204
rect 17882 2171 17898 2188
rect 17772 2154 17806 2171
rect 17686 2116 17806 2154
rect 17864 2154 17898 2171
rect 17950 2171 17966 2188
rect 18060 2188 18144 2204
rect 18060 2171 18076 2188
rect 17950 2154 17984 2171
rect 17864 2116 17984 2154
rect 18042 2154 18076 2171
rect 18128 2171 18144 2188
rect 18238 2188 18322 2204
rect 18238 2171 18254 2188
rect 18128 2154 18162 2171
rect 18042 2116 18162 2154
rect 18220 2154 18254 2171
rect 18306 2171 18322 2188
rect 18306 2154 18340 2171
rect 18220 2116 18340 2154
rect 15560 2090 15594 2108
rect 15474 2052 15594 2090
rect 16440 1798 16560 1836
rect 16440 1781 16474 1798
rect 13722 1734 13842 1772
rect 13722 1718 13756 1734
rect 13740 1700 13756 1718
rect 13808 1718 13842 1734
rect 14014 1734 14134 1772
rect 14014 1718 14048 1734
rect 13808 1700 13824 1718
rect 13740 1684 13824 1700
rect 14032 1700 14048 1718
rect 14100 1718 14134 1734
rect 14306 1734 14426 1772
rect 14306 1718 14340 1734
rect 14100 1700 14116 1718
rect 14032 1684 14116 1700
rect 14324 1700 14340 1718
rect 14392 1718 14426 1734
rect 14598 1734 14718 1772
rect 14598 1718 14632 1734
rect 14392 1700 14408 1718
rect 14324 1684 14408 1700
rect 14616 1700 14632 1718
rect 14684 1718 14718 1734
rect 14890 1734 15010 1772
rect 14890 1718 14924 1734
rect 14684 1700 14700 1718
rect 14616 1684 14700 1700
rect 14908 1700 14924 1718
rect 14976 1718 15010 1734
rect 15182 1734 15302 1772
rect 15182 1718 15216 1734
rect 14976 1700 14992 1718
rect 14908 1684 14992 1700
rect 15200 1700 15216 1718
rect 15268 1718 15302 1734
rect 15474 1734 15594 1772
rect 16458 1764 16474 1781
rect 16526 1781 16560 1798
rect 16618 1798 16738 1836
rect 16618 1781 16652 1798
rect 16526 1764 16542 1781
rect 16458 1748 16542 1764
rect 16636 1764 16652 1781
rect 16704 1781 16738 1798
rect 16796 1798 16916 1836
rect 16796 1781 16830 1798
rect 16704 1764 16720 1781
rect 16636 1748 16720 1764
rect 16814 1764 16830 1781
rect 16882 1781 16916 1798
rect 16974 1798 17094 1836
rect 16974 1781 17008 1798
rect 16882 1764 16898 1781
rect 16814 1748 16898 1764
rect 16992 1764 17008 1781
rect 17060 1781 17094 1798
rect 17152 1798 17272 1836
rect 17152 1781 17186 1798
rect 17060 1764 17076 1781
rect 16992 1748 17076 1764
rect 17170 1764 17186 1781
rect 17238 1781 17272 1798
rect 17330 1798 17450 1836
rect 17330 1781 17364 1798
rect 17238 1764 17254 1781
rect 17170 1748 17254 1764
rect 17348 1764 17364 1781
rect 17416 1781 17450 1798
rect 17508 1798 17628 1836
rect 17508 1781 17542 1798
rect 17416 1764 17432 1781
rect 17348 1748 17432 1764
rect 17526 1764 17542 1781
rect 17594 1781 17628 1798
rect 17686 1798 17806 1836
rect 17686 1781 17720 1798
rect 17594 1764 17610 1781
rect 17526 1748 17610 1764
rect 17704 1764 17720 1781
rect 17772 1781 17806 1798
rect 17864 1798 17984 1836
rect 17864 1781 17898 1798
rect 17772 1764 17788 1781
rect 17704 1748 17788 1764
rect 17882 1764 17898 1781
rect 17950 1781 17984 1798
rect 18042 1798 18162 1836
rect 18042 1781 18076 1798
rect 17950 1764 17966 1781
rect 17882 1748 17966 1764
rect 18060 1764 18076 1781
rect 18128 1781 18162 1798
rect 18220 1798 18340 1836
rect 18220 1781 18254 1798
rect 18128 1764 18144 1781
rect 18060 1748 18144 1764
rect 18238 1764 18254 1781
rect 18306 1781 18340 1798
rect 18306 1764 18322 1781
rect 18238 1748 18322 1764
rect 15474 1718 15508 1734
rect 15268 1700 15284 1718
rect 15200 1684 15284 1700
rect 15492 1700 15508 1718
rect 15560 1718 15594 1734
rect 15560 1700 15576 1718
rect 15492 1684 15576 1700
rect 13740 1626 13824 1642
rect 13740 1608 13756 1626
rect 13722 1592 13756 1608
rect 13808 1608 13824 1626
rect 14032 1626 14116 1642
rect 14032 1608 14048 1626
rect 13808 1592 13842 1608
rect 13722 1554 13842 1592
rect 14014 1592 14048 1608
rect 14100 1608 14116 1626
rect 14324 1626 14408 1642
rect 14324 1608 14340 1626
rect 14100 1592 14134 1608
rect 14014 1554 14134 1592
rect 14306 1592 14340 1608
rect 14392 1608 14408 1626
rect 14616 1626 14700 1642
rect 14616 1608 14632 1626
rect 14392 1592 14426 1608
rect 14306 1554 14426 1592
rect 14598 1592 14632 1608
rect 14684 1608 14700 1626
rect 14908 1626 14992 1642
rect 14908 1608 14924 1626
rect 14684 1592 14718 1608
rect 14598 1554 14718 1592
rect 14890 1592 14924 1608
rect 14976 1608 14992 1626
rect 15200 1626 15284 1642
rect 15200 1608 15216 1626
rect 14976 1592 15010 1608
rect 14890 1554 15010 1592
rect 15182 1592 15216 1608
rect 15268 1608 15284 1626
rect 15492 1626 15576 1642
rect 15492 1608 15508 1626
rect 15268 1592 15302 1608
rect 15182 1554 15302 1592
rect 15474 1592 15508 1608
rect 15560 1608 15576 1626
rect 16458 1628 16542 1644
rect 16458 1611 16474 1628
rect 15560 1592 15594 1608
rect 15474 1554 15594 1592
rect 16440 1594 16474 1611
rect 16526 1611 16542 1628
rect 16636 1628 16720 1644
rect 16636 1611 16652 1628
rect 16526 1594 16560 1611
rect 16440 1556 16560 1594
rect 16618 1594 16652 1611
rect 16704 1611 16720 1628
rect 16814 1628 16898 1644
rect 16814 1611 16830 1628
rect 16704 1594 16738 1611
rect 16618 1556 16738 1594
rect 16796 1594 16830 1611
rect 16882 1611 16898 1628
rect 16992 1628 17076 1644
rect 16992 1611 17008 1628
rect 16882 1594 16916 1611
rect 16796 1556 16916 1594
rect 16974 1594 17008 1611
rect 17060 1611 17076 1628
rect 17170 1628 17254 1644
rect 17170 1611 17186 1628
rect 17060 1594 17094 1611
rect 16974 1556 17094 1594
rect 17152 1594 17186 1611
rect 17238 1611 17254 1628
rect 17348 1628 17432 1644
rect 17348 1611 17364 1628
rect 17238 1594 17272 1611
rect 17152 1556 17272 1594
rect 17330 1594 17364 1611
rect 17416 1611 17432 1628
rect 17526 1628 17610 1644
rect 17526 1611 17542 1628
rect 17416 1594 17450 1611
rect 17330 1556 17450 1594
rect 17508 1594 17542 1611
rect 17594 1611 17610 1628
rect 17704 1628 17788 1644
rect 17704 1611 17720 1628
rect 17594 1594 17628 1611
rect 17508 1556 17628 1594
rect 17686 1594 17720 1611
rect 17772 1611 17788 1628
rect 17882 1628 17966 1644
rect 17882 1611 17898 1628
rect 17772 1594 17806 1611
rect 17686 1556 17806 1594
rect 17864 1594 17898 1611
rect 17950 1611 17966 1628
rect 18060 1628 18144 1644
rect 18060 1611 18076 1628
rect 17950 1594 17984 1611
rect 17864 1556 17984 1594
rect 18042 1594 18076 1611
rect 18128 1611 18144 1628
rect 18238 1628 18322 1644
rect 18238 1611 18254 1628
rect 18128 1594 18162 1611
rect 18042 1556 18162 1594
rect 18220 1594 18254 1611
rect 18306 1611 18322 1628
rect 18306 1594 18340 1611
rect 18220 1556 18340 1594
rect 13722 1236 13842 1274
rect 13722 1218 13756 1236
rect 13740 1202 13756 1218
rect 13808 1218 13842 1236
rect 14014 1236 14134 1274
rect 14014 1218 14048 1236
rect 13808 1202 13824 1218
rect 13740 1186 13824 1202
rect 14032 1202 14048 1218
rect 14100 1218 14134 1236
rect 14306 1236 14426 1274
rect 14306 1218 14340 1236
rect 14100 1202 14116 1218
rect 14032 1186 14116 1202
rect 14324 1202 14340 1218
rect 14392 1218 14426 1236
rect 14598 1236 14718 1274
rect 14598 1218 14632 1236
rect 14392 1202 14408 1218
rect 14324 1186 14408 1202
rect 14616 1202 14632 1218
rect 14684 1218 14718 1236
rect 14890 1236 15010 1274
rect 14890 1218 14924 1236
rect 14684 1202 14700 1218
rect 14616 1186 14700 1202
rect 14908 1202 14924 1218
rect 14976 1218 15010 1236
rect 15182 1236 15302 1274
rect 15182 1218 15216 1236
rect 14976 1202 14992 1218
rect 14908 1186 14992 1202
rect 15200 1202 15216 1218
rect 15268 1218 15302 1236
rect 15474 1236 15594 1274
rect 15474 1218 15508 1236
rect 15268 1202 15284 1218
rect 15200 1186 15284 1202
rect 15492 1202 15508 1218
rect 15560 1218 15594 1236
rect 16440 1238 16560 1276
rect 16440 1221 16474 1238
rect 15560 1202 15576 1218
rect 15492 1186 15576 1202
rect 16458 1204 16474 1221
rect 16526 1221 16560 1238
rect 16618 1238 16738 1276
rect 16618 1221 16652 1238
rect 16526 1204 16542 1221
rect 16458 1188 16542 1204
rect 16636 1204 16652 1221
rect 16704 1221 16738 1238
rect 16796 1238 16916 1276
rect 16796 1221 16830 1238
rect 16704 1204 16720 1221
rect 16636 1188 16720 1204
rect 16814 1204 16830 1221
rect 16882 1221 16916 1238
rect 16974 1238 17094 1276
rect 16974 1221 17008 1238
rect 16882 1204 16898 1221
rect 16814 1188 16898 1204
rect 16992 1204 17008 1221
rect 17060 1221 17094 1238
rect 17152 1238 17272 1276
rect 17152 1221 17186 1238
rect 17060 1204 17076 1221
rect 16992 1188 17076 1204
rect 17170 1204 17186 1221
rect 17238 1221 17272 1238
rect 17330 1238 17450 1276
rect 17330 1221 17364 1238
rect 17238 1204 17254 1221
rect 17170 1188 17254 1204
rect 17348 1204 17364 1221
rect 17416 1221 17450 1238
rect 17508 1238 17628 1276
rect 17508 1221 17542 1238
rect 17416 1204 17432 1221
rect 17348 1188 17432 1204
rect 17526 1204 17542 1221
rect 17594 1221 17628 1238
rect 17686 1238 17806 1276
rect 17686 1221 17720 1238
rect 17594 1204 17610 1221
rect 17526 1188 17610 1204
rect 17704 1204 17720 1221
rect 17772 1221 17806 1238
rect 17864 1238 17984 1276
rect 17864 1221 17898 1238
rect 17772 1204 17788 1221
rect 17704 1188 17788 1204
rect 17882 1204 17898 1221
rect 17950 1221 17984 1238
rect 18042 1238 18162 1276
rect 18042 1221 18076 1238
rect 17950 1204 17966 1221
rect 17882 1188 17966 1204
rect 18060 1204 18076 1221
rect 18128 1221 18162 1238
rect 18220 1238 18340 1276
rect 18220 1221 18254 1238
rect 18128 1204 18144 1221
rect 18060 1188 18144 1204
rect 18238 1204 18254 1221
rect 18306 1221 18340 1238
rect 18306 1204 18322 1221
rect 18238 1188 18322 1204
rect 13740 1128 13824 1144
rect 13740 1110 13756 1128
rect 13722 1094 13756 1110
rect 13808 1110 13824 1128
rect 14032 1128 14116 1144
rect 14032 1110 14048 1128
rect 13808 1094 13842 1110
rect 13722 1056 13842 1094
rect 14014 1094 14048 1110
rect 14100 1110 14116 1128
rect 14324 1128 14408 1144
rect 14324 1110 14340 1128
rect 14100 1094 14134 1110
rect 14014 1056 14134 1094
rect 14306 1094 14340 1110
rect 14392 1110 14408 1128
rect 14616 1128 14700 1144
rect 14616 1110 14632 1128
rect 14392 1094 14426 1110
rect 14306 1056 14426 1094
rect 14598 1094 14632 1110
rect 14684 1110 14700 1128
rect 14908 1128 14992 1144
rect 14908 1110 14924 1128
rect 14684 1094 14718 1110
rect 14598 1056 14718 1094
rect 14890 1094 14924 1110
rect 14976 1110 14992 1128
rect 15200 1128 15284 1144
rect 15200 1110 15216 1128
rect 14976 1094 15010 1110
rect 14890 1056 15010 1094
rect 15182 1094 15216 1110
rect 15268 1110 15284 1128
rect 15492 1128 15576 1144
rect 15492 1110 15508 1128
rect 15268 1094 15302 1110
rect 15182 1056 15302 1094
rect 15474 1094 15508 1110
rect 15560 1110 15576 1128
rect 16458 1128 16542 1144
rect 16458 1111 16474 1128
rect 15560 1094 15594 1110
rect 15474 1056 15594 1094
rect 16440 1094 16474 1111
rect 16526 1111 16542 1128
rect 16636 1128 16720 1144
rect 16636 1111 16652 1128
rect 16526 1094 16560 1111
rect 16440 1056 16560 1094
rect 16618 1094 16652 1111
rect 16704 1111 16720 1128
rect 16814 1128 16898 1144
rect 16814 1111 16830 1128
rect 16704 1094 16738 1111
rect 16618 1056 16738 1094
rect 16796 1094 16830 1111
rect 16882 1111 16898 1128
rect 16992 1128 17076 1144
rect 16992 1111 17008 1128
rect 16882 1094 16916 1111
rect 16796 1056 16916 1094
rect 16974 1094 17008 1111
rect 17060 1111 17076 1128
rect 17170 1128 17254 1144
rect 17170 1111 17186 1128
rect 17060 1094 17094 1111
rect 16974 1056 17094 1094
rect 17152 1094 17186 1111
rect 17238 1111 17254 1128
rect 17348 1128 17432 1144
rect 17348 1111 17364 1128
rect 17238 1094 17272 1111
rect 17152 1056 17272 1094
rect 17330 1094 17364 1111
rect 17416 1111 17432 1128
rect 17526 1128 17610 1144
rect 17526 1111 17542 1128
rect 17416 1094 17450 1111
rect 17330 1056 17450 1094
rect 17508 1094 17542 1111
rect 17594 1111 17610 1128
rect 17704 1128 17788 1144
rect 17704 1111 17720 1128
rect 17594 1094 17628 1111
rect 17508 1056 17628 1094
rect 17686 1094 17720 1111
rect 17772 1111 17788 1128
rect 17882 1128 17966 1144
rect 17882 1111 17898 1128
rect 17772 1094 17806 1111
rect 17686 1056 17806 1094
rect 17864 1094 17898 1111
rect 17950 1111 17966 1128
rect 18060 1128 18144 1144
rect 18060 1111 18076 1128
rect 17950 1094 17984 1111
rect 17864 1056 17984 1094
rect 18042 1094 18076 1111
rect 18128 1111 18144 1128
rect 18238 1128 18322 1144
rect 18238 1111 18254 1128
rect 18128 1094 18162 1111
rect 18042 1056 18162 1094
rect 18220 1094 18254 1111
rect 18306 1111 18322 1128
rect 18306 1094 18340 1111
rect 18220 1056 18340 1094
rect 13722 738 13842 776
rect 13722 720 13756 738
rect 13740 704 13756 720
rect 13808 720 13842 738
rect 14014 738 14134 776
rect 14014 720 14048 738
rect 13808 704 13824 720
rect 13740 688 13824 704
rect 14032 704 14048 720
rect 14100 720 14134 738
rect 14306 738 14426 776
rect 14306 720 14340 738
rect 14100 704 14116 720
rect 14032 688 14116 704
rect 14324 704 14340 720
rect 14392 720 14426 738
rect 14598 738 14718 776
rect 14598 720 14632 738
rect 14392 704 14408 720
rect 14324 688 14408 704
rect 14616 704 14632 720
rect 14684 720 14718 738
rect 14890 738 15010 776
rect 14890 720 14924 738
rect 14684 704 14700 720
rect 14616 688 14700 704
rect 14908 704 14924 720
rect 14976 720 15010 738
rect 15182 738 15302 776
rect 15182 720 15216 738
rect 14976 704 14992 720
rect 14908 688 14992 704
rect 15200 704 15216 720
rect 15268 720 15302 738
rect 15474 738 15594 776
rect 15474 720 15508 738
rect 15268 704 15284 720
rect 15200 688 15284 704
rect 15492 704 15508 720
rect 15560 720 15594 738
rect 16440 738 16560 776
rect 16440 721 16474 738
rect 15560 704 15576 720
rect 15492 688 15576 704
rect 16458 704 16474 721
rect 16526 721 16560 738
rect 16618 738 16738 776
rect 16618 721 16652 738
rect 16526 704 16542 721
rect 16458 688 16542 704
rect 16636 704 16652 721
rect 16704 721 16738 738
rect 16796 738 16916 776
rect 16796 721 16830 738
rect 16704 704 16720 721
rect 16636 688 16720 704
rect 16814 704 16830 721
rect 16882 721 16916 738
rect 16974 738 17094 776
rect 16974 721 17008 738
rect 16882 704 16898 721
rect 16814 688 16898 704
rect 16992 704 17008 721
rect 17060 721 17094 738
rect 17152 738 17272 776
rect 17152 721 17186 738
rect 17060 704 17076 721
rect 16992 688 17076 704
rect 17170 704 17186 721
rect 17238 721 17272 738
rect 17330 738 17450 776
rect 17330 721 17364 738
rect 17238 704 17254 721
rect 17170 688 17254 704
rect 17348 704 17364 721
rect 17416 721 17450 738
rect 17508 738 17628 776
rect 17508 721 17542 738
rect 17416 704 17432 721
rect 17348 688 17432 704
rect 17526 704 17542 721
rect 17594 721 17628 738
rect 17686 738 17806 776
rect 17686 721 17720 738
rect 17594 704 17610 721
rect 17526 688 17610 704
rect 17704 704 17720 721
rect 17772 721 17806 738
rect 17864 738 17984 776
rect 17864 721 17898 738
rect 17772 704 17788 721
rect 17704 688 17788 704
rect 17882 704 17898 721
rect 17950 721 17984 738
rect 18042 738 18162 776
rect 18042 721 18076 738
rect 17950 704 17966 721
rect 17882 688 17966 704
rect 18060 704 18076 721
rect 18128 721 18162 738
rect 18220 738 18340 776
rect 18220 721 18254 738
rect 18128 704 18144 721
rect 18060 688 18144 704
rect 18238 704 18254 721
rect 18306 721 18340 738
rect 18306 704 18322 721
rect 18238 688 18322 704
rect 19073 5122 19157 5138
rect 19073 5106 19089 5122
rect 19055 5088 19089 5106
rect 19141 5106 19157 5122
rect 19251 5122 19335 5138
rect 19251 5106 19267 5122
rect 19141 5088 19175 5106
rect 19055 5050 19175 5088
rect 19233 5088 19267 5106
rect 19319 5106 19335 5122
rect 19429 5122 19513 5138
rect 19429 5106 19445 5122
rect 19319 5088 19353 5106
rect 19233 5050 19353 5088
rect 19411 5088 19445 5106
rect 19497 5106 19513 5122
rect 19607 5122 19691 5138
rect 19607 5106 19623 5122
rect 19497 5088 19531 5106
rect 19411 5050 19531 5088
rect 19589 5088 19623 5106
rect 19675 5106 19691 5122
rect 19785 5122 19869 5138
rect 19785 5106 19801 5122
rect 19675 5088 19709 5106
rect 19589 5050 19709 5088
rect 19767 5088 19801 5106
rect 19853 5106 19869 5122
rect 19963 5122 20047 5138
rect 19963 5106 19979 5122
rect 19853 5088 19887 5106
rect 19767 5050 19887 5088
rect 19945 5088 19979 5106
rect 20031 5106 20047 5122
rect 20141 5122 20225 5138
rect 20141 5106 20157 5122
rect 20031 5088 20065 5106
rect 19945 5050 20065 5088
rect 20123 5088 20157 5106
rect 20209 5106 20225 5122
rect 20319 5122 20403 5138
rect 20319 5106 20335 5122
rect 20209 5088 20243 5106
rect 20123 5050 20243 5088
rect 20301 5088 20335 5106
rect 20387 5106 20403 5122
rect 20497 5122 20581 5138
rect 20497 5106 20513 5122
rect 20387 5088 20421 5106
rect 20301 5050 20421 5088
rect 20479 5088 20513 5106
rect 20565 5106 20581 5122
rect 20675 5122 20759 5138
rect 20675 5106 20691 5122
rect 20565 5088 20599 5106
rect 20479 5050 20599 5088
rect 20657 5088 20691 5106
rect 20743 5106 20759 5122
rect 20853 5122 20937 5138
rect 20853 5106 20869 5122
rect 20743 5088 20777 5106
rect 20657 5050 20777 5088
rect 20835 5088 20869 5106
rect 20921 5106 20937 5122
rect 21031 5122 21115 5138
rect 21031 5106 21047 5122
rect 20921 5088 20955 5106
rect 20835 5050 20955 5088
rect 21013 5088 21047 5106
rect 21099 5106 21115 5122
rect 21209 5122 21293 5138
rect 21209 5106 21225 5122
rect 21099 5088 21133 5106
rect 21013 5050 21133 5088
rect 21191 5088 21225 5106
rect 21277 5106 21293 5122
rect 21387 5122 21471 5138
rect 21387 5106 21403 5122
rect 21277 5088 21311 5106
rect 21191 5050 21311 5088
rect 21369 5088 21403 5106
rect 21455 5106 21471 5122
rect 21565 5122 21649 5138
rect 21565 5106 21581 5122
rect 21455 5088 21489 5106
rect 21369 5050 21489 5088
rect 21547 5088 21581 5106
rect 21633 5106 21649 5122
rect 21743 5122 21827 5138
rect 21743 5106 21759 5122
rect 21633 5088 21667 5106
rect 21547 5050 21667 5088
rect 21725 5088 21759 5106
rect 21811 5106 21827 5122
rect 21811 5088 21845 5106
rect 21725 5050 21845 5088
rect 19055 4732 19175 4770
rect 19055 4716 19089 4732
rect 19073 4698 19089 4716
rect 19141 4716 19175 4732
rect 19233 4732 19353 4770
rect 19233 4716 19267 4732
rect 19141 4698 19157 4716
rect 19073 4682 19157 4698
rect 19251 4698 19267 4716
rect 19319 4716 19353 4732
rect 19411 4732 19531 4770
rect 19411 4716 19445 4732
rect 19319 4698 19335 4716
rect 19251 4682 19335 4698
rect 19429 4698 19445 4716
rect 19497 4716 19531 4732
rect 19589 4732 19709 4770
rect 19589 4716 19623 4732
rect 19497 4698 19513 4716
rect 19429 4682 19513 4698
rect 19607 4698 19623 4716
rect 19675 4716 19709 4732
rect 19767 4732 19887 4770
rect 19767 4716 19801 4732
rect 19675 4698 19691 4716
rect 19607 4682 19691 4698
rect 19785 4698 19801 4716
rect 19853 4716 19887 4732
rect 19945 4732 20065 4770
rect 19945 4716 19979 4732
rect 19853 4698 19869 4716
rect 19785 4682 19869 4698
rect 19963 4698 19979 4716
rect 20031 4716 20065 4732
rect 20123 4732 20243 4770
rect 20123 4716 20157 4732
rect 20031 4698 20047 4716
rect 19963 4682 20047 4698
rect 20141 4698 20157 4716
rect 20209 4716 20243 4732
rect 20301 4732 20421 4770
rect 20301 4716 20335 4732
rect 20209 4698 20225 4716
rect 20141 4682 20225 4698
rect 20319 4698 20335 4716
rect 20387 4716 20421 4732
rect 20479 4732 20599 4770
rect 20479 4716 20513 4732
rect 20387 4698 20403 4716
rect 20319 4682 20403 4698
rect 20497 4698 20513 4716
rect 20565 4716 20599 4732
rect 20657 4732 20777 4770
rect 20657 4716 20691 4732
rect 20565 4698 20581 4716
rect 20497 4682 20581 4698
rect 20675 4698 20691 4716
rect 20743 4716 20777 4732
rect 20835 4732 20955 4770
rect 20835 4716 20869 4732
rect 20743 4698 20759 4716
rect 20675 4682 20759 4698
rect 20853 4698 20869 4716
rect 20921 4716 20955 4732
rect 21013 4732 21133 4770
rect 21013 4716 21047 4732
rect 20921 4698 20937 4716
rect 20853 4682 20937 4698
rect 21031 4698 21047 4716
rect 21099 4716 21133 4732
rect 21191 4732 21311 4770
rect 21191 4716 21225 4732
rect 21099 4698 21115 4716
rect 21031 4682 21115 4698
rect 21209 4698 21225 4716
rect 21277 4716 21311 4732
rect 21369 4732 21489 4770
rect 21369 4716 21403 4732
rect 21277 4698 21293 4716
rect 21209 4682 21293 4698
rect 21387 4698 21403 4716
rect 21455 4716 21489 4732
rect 21547 4732 21667 4770
rect 21547 4716 21581 4732
rect 21455 4698 21471 4716
rect 21387 4682 21471 4698
rect 21565 4698 21581 4716
rect 21633 4716 21667 4732
rect 21725 4732 21845 4770
rect 21725 4716 21759 4732
rect 21633 4698 21649 4716
rect 21565 4682 21649 4698
rect 21743 4698 21759 4716
rect 21811 4716 21845 4732
rect 21811 4698 21827 4716
rect 21743 4682 21827 4698
rect 19073 4624 19157 4640
rect 19073 4608 19089 4624
rect 19055 4590 19089 4608
rect 19141 4608 19157 4624
rect 19251 4624 19335 4640
rect 19251 4608 19267 4624
rect 19141 4590 19175 4608
rect 19055 4552 19175 4590
rect 19233 4590 19267 4608
rect 19319 4608 19335 4624
rect 19429 4624 19513 4640
rect 19429 4608 19445 4624
rect 19319 4590 19353 4608
rect 19233 4552 19353 4590
rect 19411 4590 19445 4608
rect 19497 4608 19513 4624
rect 19607 4624 19691 4640
rect 19607 4608 19623 4624
rect 19497 4590 19531 4608
rect 19411 4552 19531 4590
rect 19589 4590 19623 4608
rect 19675 4608 19691 4624
rect 19785 4624 19869 4640
rect 19785 4608 19801 4624
rect 19675 4590 19709 4608
rect 19589 4552 19709 4590
rect 19767 4590 19801 4608
rect 19853 4608 19869 4624
rect 19963 4624 20047 4640
rect 19963 4608 19979 4624
rect 19853 4590 19887 4608
rect 19767 4552 19887 4590
rect 19945 4590 19979 4608
rect 20031 4608 20047 4624
rect 20141 4624 20225 4640
rect 20141 4608 20157 4624
rect 20031 4590 20065 4608
rect 19945 4552 20065 4590
rect 20123 4590 20157 4608
rect 20209 4608 20225 4624
rect 20319 4624 20403 4640
rect 20319 4608 20335 4624
rect 20209 4590 20243 4608
rect 20123 4552 20243 4590
rect 20301 4590 20335 4608
rect 20387 4608 20403 4624
rect 20497 4624 20581 4640
rect 20497 4608 20513 4624
rect 20387 4590 20421 4608
rect 20301 4552 20421 4590
rect 20479 4590 20513 4608
rect 20565 4608 20581 4624
rect 20675 4624 20759 4640
rect 20675 4608 20691 4624
rect 20565 4590 20599 4608
rect 20479 4552 20599 4590
rect 20657 4590 20691 4608
rect 20743 4608 20759 4624
rect 20853 4624 20937 4640
rect 20853 4608 20869 4624
rect 20743 4590 20777 4608
rect 20657 4552 20777 4590
rect 20835 4590 20869 4608
rect 20921 4608 20937 4624
rect 21031 4624 21115 4640
rect 21031 4608 21047 4624
rect 20921 4590 20955 4608
rect 20835 4552 20955 4590
rect 21013 4590 21047 4608
rect 21099 4608 21115 4624
rect 21209 4624 21293 4640
rect 21209 4608 21225 4624
rect 21099 4590 21133 4608
rect 21013 4552 21133 4590
rect 21191 4590 21225 4608
rect 21277 4608 21293 4624
rect 21387 4624 21471 4640
rect 21387 4608 21403 4624
rect 21277 4590 21311 4608
rect 21191 4552 21311 4590
rect 21369 4590 21403 4608
rect 21455 4608 21471 4624
rect 21565 4624 21649 4640
rect 21565 4608 21581 4624
rect 21455 4590 21489 4608
rect 21369 4552 21489 4590
rect 21547 4590 21581 4608
rect 21633 4608 21649 4624
rect 21743 4624 21827 4640
rect 21743 4608 21759 4624
rect 21633 4590 21667 4608
rect 21547 4552 21667 4590
rect 21725 4590 21759 4608
rect 21811 4608 21827 4624
rect 21811 4590 21845 4608
rect 21725 4552 21845 4590
rect 19055 4234 19175 4272
rect 19055 4218 19089 4234
rect 19073 4200 19089 4218
rect 19141 4218 19175 4234
rect 19233 4234 19353 4272
rect 19233 4218 19267 4234
rect 19141 4200 19157 4218
rect 19073 4184 19157 4200
rect 19251 4200 19267 4218
rect 19319 4218 19353 4234
rect 19411 4234 19531 4272
rect 19411 4218 19445 4234
rect 19319 4200 19335 4218
rect 19251 4184 19335 4200
rect 19429 4200 19445 4218
rect 19497 4218 19531 4234
rect 19589 4234 19709 4272
rect 19589 4218 19623 4234
rect 19497 4200 19513 4218
rect 19429 4184 19513 4200
rect 19607 4200 19623 4218
rect 19675 4218 19709 4234
rect 19767 4234 19887 4272
rect 19767 4218 19801 4234
rect 19675 4200 19691 4218
rect 19607 4184 19691 4200
rect 19785 4200 19801 4218
rect 19853 4218 19887 4234
rect 19945 4234 20065 4272
rect 19945 4218 19979 4234
rect 19853 4200 19869 4218
rect 19785 4184 19869 4200
rect 19963 4200 19979 4218
rect 20031 4218 20065 4234
rect 20123 4234 20243 4272
rect 20123 4218 20157 4234
rect 20031 4200 20047 4218
rect 19963 4184 20047 4200
rect 20141 4200 20157 4218
rect 20209 4218 20243 4234
rect 20301 4234 20421 4272
rect 20301 4218 20335 4234
rect 20209 4200 20225 4218
rect 20141 4184 20225 4200
rect 20319 4200 20335 4218
rect 20387 4218 20421 4234
rect 20479 4234 20599 4272
rect 20479 4218 20513 4234
rect 20387 4200 20403 4218
rect 20319 4184 20403 4200
rect 20497 4200 20513 4218
rect 20565 4218 20599 4234
rect 20657 4234 20777 4272
rect 20657 4218 20691 4234
rect 20565 4200 20581 4218
rect 20497 4184 20581 4200
rect 20675 4200 20691 4218
rect 20743 4218 20777 4234
rect 20835 4234 20955 4272
rect 20835 4218 20869 4234
rect 20743 4200 20759 4218
rect 20675 4184 20759 4200
rect 20853 4200 20869 4218
rect 20921 4218 20955 4234
rect 21013 4234 21133 4272
rect 21013 4218 21047 4234
rect 20921 4200 20937 4218
rect 20853 4184 20937 4200
rect 21031 4200 21047 4218
rect 21099 4218 21133 4234
rect 21191 4234 21311 4272
rect 21191 4218 21225 4234
rect 21099 4200 21115 4218
rect 21031 4184 21115 4200
rect 21209 4200 21225 4218
rect 21277 4218 21311 4234
rect 21369 4234 21489 4272
rect 21369 4218 21403 4234
rect 21277 4200 21293 4218
rect 21209 4184 21293 4200
rect 21387 4200 21403 4218
rect 21455 4218 21489 4234
rect 21547 4234 21667 4272
rect 21547 4218 21581 4234
rect 21455 4200 21471 4218
rect 21387 4184 21471 4200
rect 21565 4200 21581 4218
rect 21633 4218 21667 4234
rect 21725 4234 21845 4272
rect 21725 4218 21759 4234
rect 21633 4200 21649 4218
rect 21565 4184 21649 4200
rect 21743 4200 21759 4218
rect 21811 4218 21845 4234
rect 21811 4200 21827 4218
rect 21743 4184 21827 4200
rect 19073 4126 19157 4142
rect 19073 4108 19089 4126
rect 19055 4092 19089 4108
rect 19141 4108 19157 4126
rect 19251 4126 19335 4142
rect 19251 4108 19267 4126
rect 19141 4092 19175 4108
rect 19055 4054 19175 4092
rect 19233 4092 19267 4108
rect 19319 4108 19335 4126
rect 19429 4126 19513 4142
rect 19429 4108 19445 4126
rect 19319 4092 19353 4108
rect 19233 4054 19353 4092
rect 19411 4092 19445 4108
rect 19497 4108 19513 4126
rect 19607 4126 19691 4142
rect 19607 4108 19623 4126
rect 19497 4092 19531 4108
rect 19411 4054 19531 4092
rect 19589 4092 19623 4108
rect 19675 4108 19691 4126
rect 19785 4126 19869 4142
rect 19785 4108 19801 4126
rect 19675 4092 19709 4108
rect 19589 4054 19709 4092
rect 19767 4092 19801 4108
rect 19853 4108 19869 4126
rect 19963 4126 20047 4142
rect 19963 4108 19979 4126
rect 19853 4092 19887 4108
rect 19767 4054 19887 4092
rect 19945 4092 19979 4108
rect 20031 4108 20047 4126
rect 20141 4126 20225 4142
rect 20141 4108 20157 4126
rect 20031 4092 20065 4108
rect 19945 4054 20065 4092
rect 20123 4092 20157 4108
rect 20209 4108 20225 4126
rect 20319 4126 20403 4142
rect 20319 4108 20335 4126
rect 20209 4092 20243 4108
rect 20123 4054 20243 4092
rect 20301 4092 20335 4108
rect 20387 4108 20403 4126
rect 20497 4126 20581 4142
rect 20497 4108 20513 4126
rect 20387 4092 20421 4108
rect 20301 4054 20421 4092
rect 20479 4092 20513 4108
rect 20565 4108 20581 4126
rect 20675 4126 20759 4142
rect 20675 4108 20691 4126
rect 20565 4092 20599 4108
rect 20479 4054 20599 4092
rect 20657 4092 20691 4108
rect 20743 4108 20759 4126
rect 20853 4126 20937 4142
rect 20853 4108 20869 4126
rect 20743 4092 20777 4108
rect 20657 4054 20777 4092
rect 20835 4092 20869 4108
rect 20921 4108 20937 4126
rect 21031 4126 21115 4142
rect 21031 4108 21047 4126
rect 20921 4092 20955 4108
rect 20835 4054 20955 4092
rect 21013 4092 21047 4108
rect 21099 4108 21115 4126
rect 21209 4126 21293 4142
rect 21209 4108 21225 4126
rect 21099 4092 21133 4108
rect 21013 4054 21133 4092
rect 21191 4092 21225 4108
rect 21277 4108 21293 4126
rect 21387 4126 21471 4142
rect 21387 4108 21403 4126
rect 21277 4092 21311 4108
rect 21191 4054 21311 4092
rect 21369 4092 21403 4108
rect 21455 4108 21471 4126
rect 21565 4126 21649 4142
rect 21565 4108 21581 4126
rect 21455 4092 21489 4108
rect 21369 4054 21489 4092
rect 21547 4092 21581 4108
rect 21633 4108 21649 4126
rect 21743 4126 21827 4142
rect 21743 4108 21759 4126
rect 21633 4092 21667 4108
rect 21547 4054 21667 4092
rect 21725 4092 21759 4108
rect 21811 4108 21827 4126
rect 21811 4092 21845 4108
rect 21725 4054 21845 4092
rect 19055 3736 19175 3774
rect 19055 3718 19089 3736
rect 19073 3702 19089 3718
rect 19141 3718 19175 3736
rect 19233 3736 19353 3774
rect 19233 3718 19267 3736
rect 19141 3702 19157 3718
rect 19073 3686 19157 3702
rect 19251 3702 19267 3718
rect 19319 3718 19353 3736
rect 19411 3736 19531 3774
rect 19411 3718 19445 3736
rect 19319 3702 19335 3718
rect 19251 3686 19335 3702
rect 19429 3702 19445 3718
rect 19497 3718 19531 3736
rect 19589 3736 19709 3774
rect 19589 3718 19623 3736
rect 19497 3702 19513 3718
rect 19429 3686 19513 3702
rect 19607 3702 19623 3718
rect 19675 3718 19709 3736
rect 19767 3736 19887 3774
rect 19767 3718 19801 3736
rect 19675 3702 19691 3718
rect 19607 3686 19691 3702
rect 19785 3702 19801 3718
rect 19853 3718 19887 3736
rect 19945 3736 20065 3774
rect 19945 3718 19979 3736
rect 19853 3702 19869 3718
rect 19785 3686 19869 3702
rect 19963 3702 19979 3718
rect 20031 3718 20065 3736
rect 20123 3736 20243 3774
rect 20123 3718 20157 3736
rect 20031 3702 20047 3718
rect 19963 3686 20047 3702
rect 20141 3702 20157 3718
rect 20209 3718 20243 3736
rect 20301 3736 20421 3774
rect 20301 3718 20335 3736
rect 20209 3702 20225 3718
rect 20141 3686 20225 3702
rect 20319 3702 20335 3718
rect 20387 3718 20421 3736
rect 20479 3736 20599 3774
rect 20479 3718 20513 3736
rect 20387 3702 20403 3718
rect 20319 3686 20403 3702
rect 20497 3702 20513 3718
rect 20565 3718 20599 3736
rect 20657 3736 20777 3774
rect 20657 3718 20691 3736
rect 20565 3702 20581 3718
rect 20497 3686 20581 3702
rect 20675 3702 20691 3718
rect 20743 3718 20777 3736
rect 20835 3736 20955 3774
rect 20835 3718 20869 3736
rect 20743 3702 20759 3718
rect 20675 3686 20759 3702
rect 20853 3702 20869 3718
rect 20921 3718 20955 3736
rect 21013 3736 21133 3774
rect 21013 3718 21047 3736
rect 20921 3702 20937 3718
rect 20853 3686 20937 3702
rect 21031 3702 21047 3718
rect 21099 3718 21133 3736
rect 21191 3736 21311 3774
rect 21191 3718 21225 3736
rect 21099 3702 21115 3718
rect 21031 3686 21115 3702
rect 21209 3702 21225 3718
rect 21277 3718 21311 3736
rect 21369 3736 21489 3774
rect 21369 3718 21403 3736
rect 21277 3702 21293 3718
rect 21209 3686 21293 3702
rect 21387 3702 21403 3718
rect 21455 3718 21489 3736
rect 21547 3736 21667 3774
rect 21547 3718 21581 3736
rect 21455 3702 21471 3718
rect 21387 3686 21471 3702
rect 21565 3702 21581 3718
rect 21633 3718 21667 3736
rect 21725 3736 21845 3774
rect 21725 3718 21759 3736
rect 21633 3702 21649 3718
rect 21565 3686 21649 3702
rect 21743 3702 21759 3718
rect 21811 3718 21845 3736
rect 21811 3702 21827 3718
rect 21743 3686 21827 3702
rect 19073 3628 19157 3644
rect 19073 3610 19089 3628
rect 19055 3594 19089 3610
rect 19141 3610 19157 3628
rect 19251 3628 19335 3644
rect 19251 3610 19267 3628
rect 19141 3594 19175 3610
rect 19055 3556 19175 3594
rect 19233 3594 19267 3610
rect 19319 3610 19335 3628
rect 19429 3628 19513 3644
rect 19429 3610 19445 3628
rect 19319 3594 19353 3610
rect 19233 3556 19353 3594
rect 19411 3594 19445 3610
rect 19497 3610 19513 3628
rect 19607 3628 19691 3644
rect 19607 3610 19623 3628
rect 19497 3594 19531 3610
rect 19411 3556 19531 3594
rect 19589 3594 19623 3610
rect 19675 3610 19691 3628
rect 19785 3628 19869 3644
rect 19785 3610 19801 3628
rect 19675 3594 19709 3610
rect 19589 3556 19709 3594
rect 19767 3594 19801 3610
rect 19853 3610 19869 3628
rect 19963 3628 20047 3644
rect 19963 3610 19979 3628
rect 19853 3594 19887 3610
rect 19767 3556 19887 3594
rect 19945 3594 19979 3610
rect 20031 3610 20047 3628
rect 20141 3628 20225 3644
rect 20141 3610 20157 3628
rect 20031 3594 20065 3610
rect 19945 3556 20065 3594
rect 20123 3594 20157 3610
rect 20209 3610 20225 3628
rect 20319 3628 20403 3644
rect 20319 3610 20335 3628
rect 20209 3594 20243 3610
rect 20123 3556 20243 3594
rect 20301 3594 20335 3610
rect 20387 3610 20403 3628
rect 20497 3628 20581 3644
rect 20497 3610 20513 3628
rect 20387 3594 20421 3610
rect 20301 3556 20421 3594
rect 20479 3594 20513 3610
rect 20565 3610 20581 3628
rect 20675 3628 20759 3644
rect 20675 3610 20691 3628
rect 20565 3594 20599 3610
rect 20479 3556 20599 3594
rect 20657 3594 20691 3610
rect 20743 3610 20759 3628
rect 20853 3628 20937 3644
rect 20853 3610 20869 3628
rect 20743 3594 20777 3610
rect 20657 3556 20777 3594
rect 20835 3594 20869 3610
rect 20921 3610 20937 3628
rect 21031 3628 21115 3644
rect 21031 3610 21047 3628
rect 20921 3594 20955 3610
rect 20835 3556 20955 3594
rect 21013 3594 21047 3610
rect 21099 3610 21115 3628
rect 21209 3628 21293 3644
rect 21209 3610 21225 3628
rect 21099 3594 21133 3610
rect 21013 3556 21133 3594
rect 21191 3594 21225 3610
rect 21277 3610 21293 3628
rect 21387 3628 21471 3644
rect 21387 3610 21403 3628
rect 21277 3594 21311 3610
rect 21191 3556 21311 3594
rect 21369 3594 21403 3610
rect 21455 3610 21471 3628
rect 21565 3628 21649 3644
rect 21565 3610 21581 3628
rect 21455 3594 21489 3610
rect 21369 3556 21489 3594
rect 21547 3594 21581 3610
rect 21633 3610 21649 3628
rect 21743 3628 21827 3644
rect 21743 3610 21759 3628
rect 21633 3594 21667 3610
rect 21547 3556 21667 3594
rect 21725 3594 21759 3610
rect 21811 3610 21827 3628
rect 21811 3594 21845 3610
rect 21725 3556 21845 3594
rect 19055 3238 19175 3276
rect 19055 3220 19089 3238
rect 19073 3204 19089 3220
rect 19141 3220 19175 3238
rect 19233 3238 19353 3276
rect 19233 3220 19267 3238
rect 19141 3204 19157 3220
rect 19073 3188 19157 3204
rect 19251 3204 19267 3220
rect 19319 3220 19353 3238
rect 19411 3238 19531 3276
rect 19411 3220 19445 3238
rect 19319 3204 19335 3220
rect 19251 3188 19335 3204
rect 19429 3204 19445 3220
rect 19497 3220 19531 3238
rect 19589 3238 19709 3276
rect 19589 3220 19623 3238
rect 19497 3204 19513 3220
rect 19429 3188 19513 3204
rect 19607 3204 19623 3220
rect 19675 3220 19709 3238
rect 19767 3238 19887 3276
rect 19767 3220 19801 3238
rect 19675 3204 19691 3220
rect 19607 3188 19691 3204
rect 19785 3204 19801 3220
rect 19853 3220 19887 3238
rect 19945 3238 20065 3276
rect 19945 3220 19979 3238
rect 19853 3204 19869 3220
rect 19785 3188 19869 3204
rect 19963 3204 19979 3220
rect 20031 3220 20065 3238
rect 20123 3238 20243 3276
rect 20123 3220 20157 3238
rect 20031 3204 20047 3220
rect 19963 3188 20047 3204
rect 20141 3204 20157 3220
rect 20209 3220 20243 3238
rect 20301 3238 20421 3276
rect 20301 3220 20335 3238
rect 20209 3204 20225 3220
rect 20141 3188 20225 3204
rect 20319 3204 20335 3220
rect 20387 3220 20421 3238
rect 20479 3238 20599 3276
rect 20479 3220 20513 3238
rect 20387 3204 20403 3220
rect 20319 3188 20403 3204
rect 20497 3204 20513 3220
rect 20565 3220 20599 3238
rect 20657 3238 20777 3276
rect 20657 3220 20691 3238
rect 20565 3204 20581 3220
rect 20497 3188 20581 3204
rect 20675 3204 20691 3220
rect 20743 3220 20777 3238
rect 20835 3238 20955 3276
rect 20835 3220 20869 3238
rect 20743 3204 20759 3220
rect 20675 3188 20759 3204
rect 20853 3204 20869 3220
rect 20921 3220 20955 3238
rect 21013 3238 21133 3276
rect 21013 3220 21047 3238
rect 20921 3204 20937 3220
rect 20853 3188 20937 3204
rect 21031 3204 21047 3220
rect 21099 3220 21133 3238
rect 21191 3238 21311 3276
rect 21191 3220 21225 3238
rect 21099 3204 21115 3220
rect 21031 3188 21115 3204
rect 21209 3204 21225 3220
rect 21277 3220 21311 3238
rect 21369 3238 21489 3276
rect 21369 3220 21403 3238
rect 21277 3204 21293 3220
rect 21209 3188 21293 3204
rect 21387 3204 21403 3220
rect 21455 3220 21489 3238
rect 21547 3238 21667 3276
rect 21547 3220 21581 3238
rect 21455 3204 21471 3220
rect 21387 3188 21471 3204
rect 21565 3204 21581 3220
rect 21633 3220 21667 3238
rect 21725 3238 21845 3276
rect 21725 3220 21759 3238
rect 21633 3204 21649 3220
rect 21565 3188 21649 3204
rect 21743 3204 21759 3220
rect 21811 3220 21845 3238
rect 21811 3204 21827 3220
rect 21743 3188 21827 3204
rect 19431 2614 19515 2630
rect 19431 2598 19447 2614
rect 19413 2580 19447 2598
rect 19499 2598 19515 2614
rect 19609 2614 19693 2630
rect 19609 2598 19625 2614
rect 19499 2580 19533 2598
rect 19413 2542 19533 2580
rect 19591 2580 19625 2598
rect 19677 2598 19693 2614
rect 19787 2614 19871 2630
rect 19787 2598 19803 2614
rect 19677 2580 19711 2598
rect 19591 2542 19711 2580
rect 19769 2580 19803 2598
rect 19855 2598 19871 2614
rect 19965 2614 20049 2630
rect 19965 2598 19981 2614
rect 19855 2580 19889 2598
rect 19769 2542 19889 2580
rect 19947 2580 19981 2598
rect 20033 2598 20049 2614
rect 20143 2614 20227 2630
rect 20143 2598 20159 2614
rect 20033 2580 20067 2598
rect 19947 2542 20067 2580
rect 20125 2580 20159 2598
rect 20211 2598 20227 2614
rect 20321 2614 20405 2630
rect 20321 2598 20337 2614
rect 20211 2580 20245 2598
rect 20125 2542 20245 2580
rect 20303 2580 20337 2598
rect 20389 2598 20405 2614
rect 20499 2614 20583 2630
rect 20499 2598 20515 2614
rect 20389 2580 20423 2598
rect 20303 2542 20423 2580
rect 20481 2580 20515 2598
rect 20567 2598 20583 2614
rect 20677 2614 20761 2630
rect 20677 2598 20693 2614
rect 20567 2580 20601 2598
rect 20481 2542 20601 2580
rect 20659 2580 20693 2598
rect 20745 2598 20761 2614
rect 20855 2614 20939 2630
rect 20855 2598 20871 2614
rect 20745 2580 20779 2598
rect 20659 2542 20779 2580
rect 20837 2580 20871 2598
rect 20923 2598 20939 2614
rect 21033 2614 21117 2630
rect 21033 2598 21049 2614
rect 20923 2580 20957 2598
rect 20837 2542 20957 2580
rect 21015 2580 21049 2598
rect 21101 2598 21117 2614
rect 21211 2614 21295 2630
rect 21211 2598 21227 2614
rect 21101 2580 21135 2598
rect 21015 2542 21135 2580
rect 21193 2580 21227 2598
rect 21279 2598 21295 2614
rect 21279 2580 21313 2598
rect 21193 2542 21313 2580
rect 19413 2224 19533 2262
rect 19413 2208 19447 2224
rect 19431 2190 19447 2208
rect 19499 2208 19533 2224
rect 19591 2224 19711 2262
rect 19591 2208 19625 2224
rect 19499 2190 19515 2208
rect 19431 2174 19515 2190
rect 19609 2190 19625 2208
rect 19677 2208 19711 2224
rect 19769 2224 19889 2262
rect 19769 2208 19803 2224
rect 19677 2190 19693 2208
rect 19609 2174 19693 2190
rect 19787 2190 19803 2208
rect 19855 2208 19889 2224
rect 19947 2224 20067 2262
rect 19947 2208 19981 2224
rect 19855 2190 19871 2208
rect 19787 2174 19871 2190
rect 19965 2190 19981 2208
rect 20033 2208 20067 2224
rect 20125 2224 20245 2262
rect 20125 2208 20159 2224
rect 20033 2190 20049 2208
rect 19965 2174 20049 2190
rect 20143 2190 20159 2208
rect 20211 2208 20245 2224
rect 20303 2224 20423 2262
rect 20303 2208 20337 2224
rect 20211 2190 20227 2208
rect 20143 2174 20227 2190
rect 20321 2190 20337 2208
rect 20389 2208 20423 2224
rect 20481 2224 20601 2262
rect 20481 2208 20515 2224
rect 20389 2190 20405 2208
rect 20321 2174 20405 2190
rect 20499 2190 20515 2208
rect 20567 2208 20601 2224
rect 20659 2224 20779 2262
rect 20659 2208 20693 2224
rect 20567 2190 20583 2208
rect 20499 2174 20583 2190
rect 20677 2190 20693 2208
rect 20745 2208 20779 2224
rect 20837 2224 20957 2262
rect 20837 2208 20871 2224
rect 20745 2190 20761 2208
rect 20677 2174 20761 2190
rect 20855 2190 20871 2208
rect 20923 2208 20957 2224
rect 21015 2224 21135 2262
rect 21015 2208 21049 2224
rect 20923 2190 20939 2208
rect 20855 2174 20939 2190
rect 21033 2190 21049 2208
rect 21101 2208 21135 2224
rect 21193 2224 21313 2262
rect 21193 2208 21227 2224
rect 21101 2190 21117 2208
rect 21033 2174 21117 2190
rect 21211 2190 21227 2208
rect 21279 2208 21313 2224
rect 21279 2190 21295 2208
rect 21211 2174 21295 2190
rect 19431 2116 19515 2132
rect 19431 2100 19447 2116
rect 19413 2082 19447 2100
rect 19499 2100 19515 2116
rect 19609 2116 19693 2132
rect 19609 2100 19625 2116
rect 19499 2082 19533 2100
rect 19413 2044 19533 2082
rect 19591 2082 19625 2100
rect 19677 2100 19693 2116
rect 19787 2116 19871 2132
rect 19787 2100 19803 2116
rect 19677 2082 19711 2100
rect 19591 2044 19711 2082
rect 19769 2082 19803 2100
rect 19855 2100 19871 2116
rect 19965 2116 20049 2132
rect 19965 2100 19981 2116
rect 19855 2082 19889 2100
rect 19769 2044 19889 2082
rect 19947 2082 19981 2100
rect 20033 2100 20049 2116
rect 20143 2116 20227 2132
rect 20143 2100 20159 2116
rect 20033 2082 20067 2100
rect 19947 2044 20067 2082
rect 20125 2082 20159 2100
rect 20211 2100 20227 2116
rect 20321 2116 20405 2132
rect 20321 2100 20337 2116
rect 20211 2082 20245 2100
rect 20125 2044 20245 2082
rect 20303 2082 20337 2100
rect 20389 2100 20405 2116
rect 20499 2116 20583 2132
rect 20499 2100 20515 2116
rect 20389 2082 20423 2100
rect 20303 2044 20423 2082
rect 20481 2082 20515 2100
rect 20567 2100 20583 2116
rect 20677 2116 20761 2132
rect 20677 2100 20693 2116
rect 20567 2082 20601 2100
rect 20481 2044 20601 2082
rect 20659 2082 20693 2100
rect 20745 2100 20761 2116
rect 20855 2116 20939 2132
rect 20855 2100 20871 2116
rect 20745 2082 20779 2100
rect 20659 2044 20779 2082
rect 20837 2082 20871 2100
rect 20923 2100 20939 2116
rect 21033 2116 21117 2132
rect 21033 2100 21049 2116
rect 20923 2082 20957 2100
rect 20837 2044 20957 2082
rect 21015 2082 21049 2100
rect 21101 2100 21117 2116
rect 21211 2116 21295 2132
rect 21211 2100 21227 2116
rect 21101 2082 21135 2100
rect 21015 2044 21135 2082
rect 21193 2082 21227 2100
rect 21279 2100 21295 2116
rect 21279 2082 21313 2100
rect 21193 2044 21313 2082
rect 19413 1726 19533 1764
rect 19413 1710 19447 1726
rect 19431 1692 19447 1710
rect 19499 1710 19533 1726
rect 19591 1726 19711 1764
rect 19591 1710 19625 1726
rect 19499 1692 19515 1710
rect 19431 1676 19515 1692
rect 19609 1692 19625 1710
rect 19677 1710 19711 1726
rect 19769 1726 19889 1764
rect 19769 1710 19803 1726
rect 19677 1692 19693 1710
rect 19609 1676 19693 1692
rect 19787 1692 19803 1710
rect 19855 1710 19889 1726
rect 19947 1726 20067 1764
rect 19947 1710 19981 1726
rect 19855 1692 19871 1710
rect 19787 1676 19871 1692
rect 19965 1692 19981 1710
rect 20033 1710 20067 1726
rect 20125 1726 20245 1764
rect 20125 1710 20159 1726
rect 20033 1692 20049 1710
rect 19965 1676 20049 1692
rect 20143 1692 20159 1710
rect 20211 1710 20245 1726
rect 20303 1726 20423 1764
rect 20303 1710 20337 1726
rect 20211 1692 20227 1710
rect 20143 1676 20227 1692
rect 20321 1692 20337 1710
rect 20389 1710 20423 1726
rect 20481 1726 20601 1764
rect 20481 1710 20515 1726
rect 20389 1692 20405 1710
rect 20321 1676 20405 1692
rect 20499 1692 20515 1710
rect 20567 1710 20601 1726
rect 20659 1726 20779 1764
rect 20659 1710 20693 1726
rect 20567 1692 20583 1710
rect 20499 1676 20583 1692
rect 20677 1692 20693 1710
rect 20745 1710 20779 1726
rect 20837 1726 20957 1764
rect 20837 1710 20871 1726
rect 20745 1692 20761 1710
rect 20677 1676 20761 1692
rect 20855 1692 20871 1710
rect 20923 1710 20957 1726
rect 21015 1726 21135 1764
rect 21015 1710 21049 1726
rect 20923 1692 20939 1710
rect 20855 1676 20939 1692
rect 21033 1692 21049 1710
rect 21101 1710 21135 1726
rect 21193 1726 21313 1764
rect 21193 1710 21227 1726
rect 21101 1692 21117 1710
rect 21033 1676 21117 1692
rect 21211 1692 21227 1710
rect 21279 1710 21313 1726
rect 21279 1692 21295 1710
rect 21211 1676 21295 1692
rect 19431 1618 19515 1634
rect 19431 1600 19447 1618
rect 19413 1584 19447 1600
rect 19499 1600 19515 1618
rect 19609 1618 19693 1634
rect 19609 1600 19625 1618
rect 19499 1584 19533 1600
rect 19413 1546 19533 1584
rect 19591 1584 19625 1600
rect 19677 1600 19693 1618
rect 19787 1618 19871 1634
rect 19787 1600 19803 1618
rect 19677 1584 19711 1600
rect 19591 1546 19711 1584
rect 19769 1584 19803 1600
rect 19855 1600 19871 1618
rect 19965 1618 20049 1634
rect 19965 1600 19981 1618
rect 19855 1584 19889 1600
rect 19769 1546 19889 1584
rect 19947 1584 19981 1600
rect 20033 1600 20049 1618
rect 20143 1618 20227 1634
rect 20143 1600 20159 1618
rect 20033 1584 20067 1600
rect 19947 1546 20067 1584
rect 20125 1584 20159 1600
rect 20211 1600 20227 1618
rect 20321 1618 20405 1634
rect 20321 1600 20337 1618
rect 20211 1584 20245 1600
rect 20125 1546 20245 1584
rect 20303 1584 20337 1600
rect 20389 1600 20405 1618
rect 20499 1618 20583 1634
rect 20499 1600 20515 1618
rect 20389 1584 20423 1600
rect 20303 1546 20423 1584
rect 20481 1584 20515 1600
rect 20567 1600 20583 1618
rect 20677 1618 20761 1634
rect 20677 1600 20693 1618
rect 20567 1584 20601 1600
rect 20481 1546 20601 1584
rect 20659 1584 20693 1600
rect 20745 1600 20761 1618
rect 20855 1618 20939 1634
rect 20855 1600 20871 1618
rect 20745 1584 20779 1600
rect 20659 1546 20779 1584
rect 20837 1584 20871 1600
rect 20923 1600 20939 1618
rect 21033 1618 21117 1634
rect 21033 1600 21049 1618
rect 20923 1584 20957 1600
rect 20837 1546 20957 1584
rect 21015 1584 21049 1600
rect 21101 1600 21117 1618
rect 21211 1618 21295 1634
rect 21211 1600 21227 1618
rect 21101 1584 21135 1600
rect 21015 1546 21135 1584
rect 21193 1584 21227 1600
rect 21279 1600 21295 1618
rect 21279 1584 21313 1600
rect 21193 1546 21313 1584
rect 19413 1228 19533 1266
rect 19413 1210 19447 1228
rect 19431 1194 19447 1210
rect 19499 1210 19533 1228
rect 19591 1228 19711 1266
rect 19591 1210 19625 1228
rect 19499 1194 19515 1210
rect 19431 1178 19515 1194
rect 19609 1194 19625 1210
rect 19677 1210 19711 1228
rect 19769 1228 19889 1266
rect 19769 1210 19803 1228
rect 19677 1194 19693 1210
rect 19609 1178 19693 1194
rect 19787 1194 19803 1210
rect 19855 1210 19889 1228
rect 19947 1228 20067 1266
rect 19947 1210 19981 1228
rect 19855 1194 19871 1210
rect 19787 1178 19871 1194
rect 19965 1194 19981 1210
rect 20033 1210 20067 1228
rect 20125 1228 20245 1266
rect 20125 1210 20159 1228
rect 20033 1194 20049 1210
rect 19965 1178 20049 1194
rect 20143 1194 20159 1210
rect 20211 1210 20245 1228
rect 20303 1228 20423 1266
rect 20303 1210 20337 1228
rect 20211 1194 20227 1210
rect 20143 1178 20227 1194
rect 20321 1194 20337 1210
rect 20389 1210 20423 1228
rect 20481 1228 20601 1266
rect 20481 1210 20515 1228
rect 20389 1194 20405 1210
rect 20321 1178 20405 1194
rect 20499 1194 20515 1210
rect 20567 1210 20601 1228
rect 20659 1228 20779 1266
rect 20659 1210 20693 1228
rect 20567 1194 20583 1210
rect 20499 1178 20583 1194
rect 20677 1194 20693 1210
rect 20745 1210 20779 1228
rect 20837 1228 20957 1266
rect 20837 1210 20871 1228
rect 20745 1194 20761 1210
rect 20677 1178 20761 1194
rect 20855 1194 20871 1210
rect 20923 1210 20957 1228
rect 21015 1228 21135 1266
rect 21015 1210 21049 1228
rect 20923 1194 20939 1210
rect 20855 1178 20939 1194
rect 21033 1194 21049 1210
rect 21101 1210 21135 1228
rect 21193 1228 21313 1266
rect 21193 1210 21227 1228
rect 21101 1194 21117 1210
rect 21033 1178 21117 1194
rect 21211 1194 21227 1210
rect 21279 1210 21313 1228
rect 21279 1194 21295 1210
rect 21211 1178 21295 1194
rect 19431 1120 19515 1136
rect 19431 1102 19447 1120
rect 19413 1086 19447 1102
rect 19499 1102 19515 1120
rect 19609 1120 19693 1136
rect 19609 1102 19625 1120
rect 19499 1086 19533 1102
rect 19413 1048 19533 1086
rect 19591 1086 19625 1102
rect 19677 1102 19693 1120
rect 19787 1120 19871 1136
rect 19787 1102 19803 1120
rect 19677 1086 19711 1102
rect 19591 1048 19711 1086
rect 19769 1086 19803 1102
rect 19855 1102 19871 1120
rect 19965 1120 20049 1136
rect 19965 1102 19981 1120
rect 19855 1086 19889 1102
rect 19769 1048 19889 1086
rect 19947 1086 19981 1102
rect 20033 1102 20049 1120
rect 20143 1120 20227 1136
rect 20143 1102 20159 1120
rect 20033 1086 20067 1102
rect 19947 1048 20067 1086
rect 20125 1086 20159 1102
rect 20211 1102 20227 1120
rect 20321 1120 20405 1136
rect 20321 1102 20337 1120
rect 20211 1086 20245 1102
rect 20125 1048 20245 1086
rect 20303 1086 20337 1102
rect 20389 1102 20405 1120
rect 20499 1120 20583 1136
rect 20499 1102 20515 1120
rect 20389 1086 20423 1102
rect 20303 1048 20423 1086
rect 20481 1086 20515 1102
rect 20567 1102 20583 1120
rect 20677 1120 20761 1136
rect 20677 1102 20693 1120
rect 20567 1086 20601 1102
rect 20481 1048 20601 1086
rect 20659 1086 20693 1102
rect 20745 1102 20761 1120
rect 20855 1120 20939 1136
rect 20855 1102 20871 1120
rect 20745 1086 20779 1102
rect 20659 1048 20779 1086
rect 20837 1086 20871 1102
rect 20923 1102 20939 1120
rect 21033 1120 21117 1136
rect 21033 1102 21049 1120
rect 20923 1086 20957 1102
rect 20837 1048 20957 1086
rect 21015 1086 21049 1102
rect 21101 1102 21117 1120
rect 21211 1120 21295 1136
rect 21211 1102 21227 1120
rect 21101 1086 21135 1102
rect 21015 1048 21135 1086
rect 21193 1086 21227 1102
rect 21279 1102 21295 1120
rect 21279 1086 21313 1102
rect 21193 1048 21313 1086
rect 19413 730 19533 768
rect 19413 712 19447 730
rect 19431 696 19447 712
rect 19499 712 19533 730
rect 19591 730 19711 768
rect 19591 712 19625 730
rect 19499 696 19515 712
rect 19431 680 19515 696
rect 19609 696 19625 712
rect 19677 712 19711 730
rect 19769 730 19889 768
rect 19769 712 19803 730
rect 19677 696 19693 712
rect 19609 680 19693 696
rect 19787 696 19803 712
rect 19855 712 19889 730
rect 19947 730 20067 768
rect 19947 712 19981 730
rect 19855 696 19871 712
rect 19787 680 19871 696
rect 19965 696 19981 712
rect 20033 712 20067 730
rect 20125 730 20245 768
rect 20125 712 20159 730
rect 20033 696 20049 712
rect 19965 680 20049 696
rect 20143 696 20159 712
rect 20211 712 20245 730
rect 20303 730 20423 768
rect 20303 712 20337 730
rect 20211 696 20227 712
rect 20143 680 20227 696
rect 20321 696 20337 712
rect 20389 712 20423 730
rect 20481 730 20601 768
rect 20481 712 20515 730
rect 20389 696 20405 712
rect 20321 680 20405 696
rect 20499 696 20515 712
rect 20567 712 20601 730
rect 20659 730 20779 768
rect 20659 712 20693 730
rect 20567 696 20583 712
rect 20499 680 20583 696
rect 20677 696 20693 712
rect 20745 712 20779 730
rect 20837 730 20957 768
rect 20837 712 20871 730
rect 20745 696 20761 712
rect 20677 680 20761 696
rect 20855 696 20871 712
rect 20923 712 20957 730
rect 21015 730 21135 768
rect 21015 712 21049 730
rect 20923 696 20939 712
rect 20855 680 20939 696
rect 21033 696 21049 712
rect 21101 712 21135 730
rect 21193 730 21313 768
rect 21193 712 21227 730
rect 21101 696 21117 712
rect 21033 680 21117 696
rect 21211 696 21227 712
rect 21279 712 21313 730
rect 21279 696 21295 712
rect 21211 680 21295 696
<< polycont >>
rect 7303 18801 7337 18835
rect 7495 18801 7529 18835
rect 7687 18801 7721 18835
rect 7879 18801 7913 18835
rect 8071 18801 8105 18835
rect 8263 18801 8297 18835
rect 20233 18801 20267 18835
rect 20425 18801 20459 18835
rect 20617 18801 20651 18835
rect 20809 18801 20843 18835
rect 21001 18801 21035 18835
rect 21193 18801 21227 18835
rect 7303 17990 7337 18024
rect 7495 17990 7529 18024
rect 7687 17990 7721 18024
rect 7879 17990 7913 18024
rect 8071 17990 8105 18024
rect 8263 17990 8297 18024
rect 20233 17990 20267 18024
rect 20425 17990 20459 18024
rect 20617 17990 20651 18024
rect 20809 17990 20843 18024
rect 21001 17990 21035 18024
rect 21193 17990 21227 18024
rect 7303 17001 7337 17035
rect 7495 17001 7529 17035
rect 7687 17001 7721 17035
rect 7879 17001 7913 17035
rect 8071 17001 8105 17035
rect 8263 17001 8297 17035
rect 20233 17001 20267 17035
rect 20425 17001 20459 17035
rect 20617 17001 20651 17035
rect 20809 17001 20843 17035
rect 21001 17001 21035 17035
rect 21193 17001 21227 17035
rect 7303 16190 7337 16224
rect 7495 16190 7529 16224
rect 7687 16190 7721 16224
rect 7879 16190 7913 16224
rect 8071 16190 8105 16224
rect 8263 16190 8297 16224
rect 20233 16190 20267 16224
rect 20425 16190 20459 16224
rect 20617 16190 20651 16224
rect 20809 16190 20843 16224
rect 21001 16190 21035 16224
rect 21193 16190 21227 16224
rect 7303 15201 7337 15235
rect 7495 15201 7529 15235
rect 7687 15201 7721 15235
rect 7879 15201 7913 15235
rect 8071 15201 8105 15235
rect 8263 15201 8297 15235
rect 20233 15201 20267 15235
rect 20425 15201 20459 15235
rect 20617 15201 20651 15235
rect 20809 15201 20843 15235
rect 21001 15201 21035 15235
rect 21193 15201 21227 15235
rect 7303 14390 7337 14424
rect 7495 14390 7529 14424
rect 7687 14390 7721 14424
rect 7879 14390 7913 14424
rect 8071 14390 8105 14424
rect 8263 14390 8297 14424
rect 20233 14390 20267 14424
rect 20425 14390 20459 14424
rect 20617 14390 20651 14424
rect 20809 14390 20843 14424
rect 21001 14390 21035 14424
rect 21193 14390 21227 14424
rect 7303 13401 7337 13435
rect 7495 13401 7529 13435
rect 7687 13401 7721 13435
rect 7879 13401 7913 13435
rect 8071 13401 8105 13435
rect 8263 13401 8297 13435
rect 20233 13401 20267 13435
rect 20425 13401 20459 13435
rect 20617 13401 20651 13435
rect 20809 13401 20843 13435
rect 21001 13401 21035 13435
rect 21193 13401 21227 13435
rect 7303 12590 7337 12624
rect 7495 12590 7529 12624
rect 7687 12590 7721 12624
rect 7879 12590 7913 12624
rect 8071 12590 8105 12624
rect 8263 12590 8297 12624
rect 20233 12590 20267 12624
rect 20425 12590 20459 12624
rect 20617 12590 20651 12624
rect 20809 12590 20843 12624
rect 21001 12590 21035 12624
rect 21193 12590 21227 12624
rect 7303 11601 7337 11635
rect 7495 11601 7529 11635
rect 7687 11601 7721 11635
rect 7879 11601 7913 11635
rect 8071 11601 8105 11635
rect 8263 11601 8297 11635
rect 20233 11601 20267 11635
rect 20425 11601 20459 11635
rect 20617 11601 20651 11635
rect 20809 11601 20843 11635
rect 21001 11601 21035 11635
rect 21193 11601 21227 11635
rect 7303 10790 7337 10824
rect 7495 10790 7529 10824
rect 7687 10790 7721 10824
rect 7879 10790 7913 10824
rect 8071 10790 8105 10824
rect 8263 10790 8297 10824
rect 20233 10790 20267 10824
rect 20425 10790 20459 10824
rect 20617 10790 20651 10824
rect 20809 10790 20843 10824
rect 21001 10790 21035 10824
rect 21193 10790 21227 10824
rect 7303 9801 7337 9835
rect 7495 9801 7529 9835
rect 7687 9801 7721 9835
rect 7879 9801 7913 9835
rect 8071 9801 8105 9835
rect 8263 9801 8297 9835
rect 20233 9801 20267 9835
rect 20425 9801 20459 9835
rect 20617 9801 20651 9835
rect 20809 9801 20843 9835
rect 21001 9801 21035 9835
rect 21193 9801 21227 9835
rect 7303 8990 7337 9024
rect 7495 8990 7529 9024
rect 7687 8990 7721 9024
rect 7879 8990 7913 9024
rect 8071 8990 8105 9024
rect 8263 8990 8297 9024
rect 20233 8990 20267 9024
rect 20425 8990 20459 9024
rect 20617 8990 20651 9024
rect 20809 8990 20843 9024
rect 21001 8990 21035 9024
rect 21193 8990 21227 9024
rect 2100 4269 2134 4303
rect 2524 4269 2558 4303
rect 2946 4269 2980 4303
rect 3370 4269 3404 4303
rect 3880 4269 3914 4303
rect 4304 4269 4338 4303
rect 4726 4269 4760 4303
rect 5150 4269 5184 4303
rect 2312 3919 2346 3953
rect 2736 3919 2770 3953
rect 3158 3919 3192 3953
rect 3582 3919 3616 3953
rect 4092 3919 4126 3953
rect 4516 3919 4550 3953
rect 4938 3919 4972 3953
rect 5362 3919 5396 3953
rect 7636 6656 7688 6690
rect 7814 6656 7866 6690
rect 7992 6656 8044 6690
rect 8170 6656 8222 6690
rect 8348 6656 8400 6690
rect 8526 6656 8578 6690
rect 8704 6656 8756 6690
rect 8882 6656 8934 6690
rect 9060 6656 9112 6690
rect 9238 6656 9290 6690
rect 9416 6656 9468 6690
rect 9594 6656 9646 6690
rect 9772 6656 9824 6690
rect 9950 6656 10002 6690
rect 10322 6656 10374 6690
rect 10500 6656 10552 6690
rect 10678 6656 10730 6690
rect 10856 6656 10908 6690
rect 11034 6656 11086 6690
rect 11212 6656 11264 6690
rect 11390 6656 11442 6690
rect 11568 6656 11620 6690
rect 11746 6656 11798 6690
rect 11924 6656 11976 6690
rect 12102 6656 12154 6690
rect 12280 6656 12332 6690
rect 12458 6656 12510 6690
rect 12636 6656 12688 6690
rect 7636 6248 7688 6282
rect 7814 6248 7866 6282
rect 7992 6248 8044 6282
rect 8170 6248 8222 6282
rect 8348 6248 8400 6282
rect 8526 6248 8578 6282
rect 8704 6248 8756 6282
rect 8882 6248 8934 6282
rect 9060 6248 9112 6282
rect 9238 6248 9290 6282
rect 9416 6248 9468 6282
rect 9594 6248 9646 6282
rect 9772 6248 9824 6282
rect 9950 6248 10002 6282
rect 10322 6248 10374 6282
rect 10500 6248 10552 6282
rect 10678 6248 10730 6282
rect 10856 6248 10908 6282
rect 11034 6248 11086 6282
rect 11212 6248 11264 6282
rect 11390 6248 11442 6282
rect 11568 6248 11620 6282
rect 11746 6248 11798 6282
rect 11924 6248 11976 6282
rect 12102 6248 12154 6282
rect 12280 6248 12332 6282
rect 12458 6248 12510 6282
rect 12636 6248 12688 6282
rect 7636 6078 7688 6112
rect 7814 6078 7866 6112
rect 7992 6078 8044 6112
rect 8170 6078 8222 6112
rect 8348 6078 8400 6112
rect 8526 6078 8578 6112
rect 8704 6078 8756 6112
rect 8882 6078 8934 6112
rect 9060 6078 9112 6112
rect 9238 6078 9290 6112
rect 9416 6078 9468 6112
rect 9594 6078 9646 6112
rect 9772 6078 9824 6112
rect 9950 6078 10002 6112
rect 10322 6079 10374 6113
rect 10500 6079 10552 6113
rect 10678 6079 10730 6113
rect 10856 6079 10908 6113
rect 11034 6079 11086 6113
rect 11212 6079 11264 6113
rect 11390 6079 11442 6113
rect 11568 6079 11620 6113
rect 11746 6079 11798 6113
rect 11924 6079 11976 6113
rect 12102 6079 12154 6113
rect 12280 6079 12332 6113
rect 12458 6079 12510 6113
rect 12636 6079 12688 6113
rect 7636 5670 7688 5704
rect 7814 5670 7866 5704
rect 7992 5670 8044 5704
rect 8170 5670 8222 5704
rect 8348 5670 8400 5704
rect 8526 5670 8578 5704
rect 8704 5670 8756 5704
rect 8882 5670 8934 5704
rect 9060 5670 9112 5704
rect 9238 5670 9290 5704
rect 9416 5670 9468 5704
rect 9594 5670 9646 5704
rect 9772 5670 9824 5704
rect 9950 5670 10002 5704
rect 10322 5671 10374 5705
rect 10500 5671 10552 5705
rect 10678 5671 10730 5705
rect 10856 5671 10908 5705
rect 11034 5671 11086 5705
rect 11212 5671 11264 5705
rect 11390 5671 11442 5705
rect 11568 5671 11620 5705
rect 11746 5671 11798 5705
rect 11924 5671 11976 5705
rect 12102 5671 12154 5705
rect 12280 5671 12332 5705
rect 12458 5671 12510 5705
rect 12636 5671 12688 5705
rect 14776 6725 14828 6759
rect 14954 6725 15006 6759
rect 15132 6725 15184 6759
rect 15310 6725 15362 6759
rect 15488 6725 15540 6759
rect 15666 6725 15718 6759
rect 15844 6725 15896 6759
rect 16022 6725 16074 6759
rect 16976 6725 17028 6759
rect 17154 6725 17206 6759
rect 17332 6725 17384 6759
rect 17510 6725 17562 6759
rect 17688 6725 17740 6759
rect 17866 6725 17918 6759
rect 18044 6725 18096 6759
rect 18222 6725 18274 6759
rect 19176 6725 19228 6759
rect 19354 6725 19406 6759
rect 19532 6725 19584 6759
rect 19710 6725 19762 6759
rect 19888 6725 19940 6759
rect 20066 6725 20118 6759
rect 20244 6725 20296 6759
rect 20422 6725 20474 6759
rect 14776 6317 14828 6351
rect 14954 6317 15006 6351
rect 15132 6317 15184 6351
rect 15310 6317 15362 6351
rect 15488 6317 15540 6351
rect 15666 6317 15718 6351
rect 15844 6317 15896 6351
rect 16022 6317 16074 6351
rect 16976 6317 17028 6351
rect 17154 6317 17206 6351
rect 17332 6317 17384 6351
rect 17510 6317 17562 6351
rect 17688 6317 17740 6351
rect 17866 6317 17918 6351
rect 18044 6317 18096 6351
rect 18222 6317 18274 6351
rect 19176 6317 19228 6351
rect 19354 6317 19406 6351
rect 19532 6317 19584 6351
rect 19710 6317 19762 6351
rect 19888 6317 19940 6351
rect 20066 6317 20118 6351
rect 20244 6317 20296 6351
rect 20422 6317 20474 6351
rect 14777 5958 14829 5992
rect 14955 5958 15007 5992
rect 15133 5958 15185 5992
rect 15311 5958 15363 5992
rect 15489 5958 15541 5992
rect 15667 5958 15719 5992
rect 15845 5958 15897 5992
rect 16023 5958 16075 5992
rect 16977 5958 17029 5992
rect 17155 5958 17207 5992
rect 17333 5958 17385 5992
rect 17511 5958 17563 5992
rect 17689 5958 17741 5992
rect 17867 5958 17919 5992
rect 18045 5958 18097 5992
rect 18223 5958 18275 5992
rect 19177 5958 19229 5992
rect 19355 5958 19407 5992
rect 19533 5958 19585 5992
rect 19711 5958 19763 5992
rect 19889 5958 19941 5992
rect 20067 5958 20119 5992
rect 20245 5958 20297 5992
rect 20423 5958 20475 5992
rect 14777 5550 14829 5584
rect 14955 5550 15007 5584
rect 15133 5550 15185 5584
rect 15311 5550 15363 5584
rect 15489 5550 15541 5584
rect 15667 5550 15719 5584
rect 15845 5550 15897 5584
rect 16023 5550 16075 5584
rect 16977 5550 17029 5584
rect 17155 5550 17207 5584
rect 17333 5550 17385 5584
rect 17511 5550 17563 5584
rect 17689 5550 17741 5584
rect 17867 5550 17919 5584
rect 18045 5550 18097 5584
rect 18223 5550 18275 5584
rect 19177 5550 19229 5584
rect 19355 5550 19407 5584
rect 19533 5550 19585 5584
rect 19711 5550 19763 5584
rect 19889 5550 19941 5584
rect 20067 5550 20119 5584
rect 20245 5550 20297 5584
rect 20423 5550 20475 5584
rect 7992 5198 8044 5232
rect 8170 5198 8222 5232
rect 8348 5198 8400 5232
rect 8526 5198 8578 5232
rect 8704 5198 8756 5232
rect 8882 5198 8934 5232
rect 9060 5198 9112 5232
rect 9238 5198 9290 5232
rect 9416 5198 9468 5232
rect 9594 5198 9646 5232
rect 9772 5198 9824 5232
rect 9950 5198 10002 5232
rect 10322 5198 10374 5232
rect 10500 5198 10552 5232
rect 10678 5198 10730 5232
rect 10856 5198 10908 5232
rect 11034 5198 11086 5232
rect 11212 5198 11264 5232
rect 11390 5198 11442 5232
rect 11568 5198 11620 5232
rect 11746 5198 11798 5232
rect 11924 5198 11976 5232
rect 12102 5198 12154 5232
rect 12280 5198 12332 5232
rect 7992 4790 8044 4824
rect 8170 4790 8222 4824
rect 8348 4790 8400 4824
rect 8526 4790 8578 4824
rect 8704 4790 8756 4824
rect 8882 4790 8934 4824
rect 9060 4790 9112 4824
rect 9238 4790 9290 4824
rect 9416 4790 9468 4824
rect 9594 4790 9646 4824
rect 9772 4790 9824 4824
rect 9950 4790 10002 4824
rect 10322 4790 10374 4824
rect 10500 4790 10552 4824
rect 10678 4790 10730 4824
rect 10856 4790 10908 4824
rect 11034 4790 11086 4824
rect 11212 4790 11264 4824
rect 11390 4790 11442 4824
rect 11568 4790 11620 4824
rect 11746 4790 11798 4824
rect 11924 4790 11976 4824
rect 12102 4790 12154 4824
rect 12280 4790 12332 4824
rect 7992 4628 8044 4662
rect 8170 4628 8222 4662
rect 8348 4628 8400 4662
rect 8526 4628 8578 4662
rect 8704 4628 8756 4662
rect 8882 4628 8934 4662
rect 9060 4628 9112 4662
rect 9238 4628 9290 4662
rect 9416 4628 9468 4662
rect 9594 4628 9646 4662
rect 9772 4628 9824 4662
rect 9950 4628 10002 4662
rect 10322 4628 10374 4662
rect 10500 4628 10552 4662
rect 10678 4628 10730 4662
rect 10856 4628 10908 4662
rect 11034 4628 11086 4662
rect 11212 4628 11264 4662
rect 11390 4628 11442 4662
rect 11568 4628 11620 4662
rect 11746 4628 11798 4662
rect 11924 4628 11976 4662
rect 12102 4628 12154 4662
rect 12280 4628 12332 4662
rect 7992 4220 8044 4254
rect 8170 4220 8222 4254
rect 8348 4220 8400 4254
rect 8526 4220 8578 4254
rect 8704 4220 8756 4254
rect 8882 4220 8934 4254
rect 9060 4220 9112 4254
rect 9238 4220 9290 4254
rect 9416 4220 9468 4254
rect 9594 4220 9646 4254
rect 9772 4220 9824 4254
rect 9950 4220 10002 4254
rect 10322 4220 10374 4254
rect 10500 4220 10552 4254
rect 10678 4220 10730 4254
rect 10856 4220 10908 4254
rect 11034 4220 11086 4254
rect 11212 4220 11264 4254
rect 11390 4220 11442 4254
rect 11568 4220 11620 4254
rect 11746 4220 11798 4254
rect 11924 4220 11976 4254
rect 12102 4220 12154 4254
rect 12280 4220 12332 4254
rect 7637 3689 7689 3723
rect 7815 3689 7867 3723
rect 7993 3689 8045 3723
rect 8171 3689 8223 3723
rect 8349 3689 8401 3723
rect 8527 3689 8579 3723
rect 8705 3689 8757 3723
rect 8883 3689 8935 3723
rect 9061 3689 9113 3723
rect 9239 3689 9291 3723
rect 9417 3689 9469 3723
rect 9595 3689 9647 3723
rect 9773 3689 9825 3723
rect 9951 3689 10003 3723
rect 10324 3689 10376 3723
rect 10502 3689 10554 3723
rect 10680 3689 10732 3723
rect 10858 3689 10910 3723
rect 11036 3689 11088 3723
rect 11214 3689 11266 3723
rect 11392 3689 11444 3723
rect 11570 3689 11622 3723
rect 11748 3689 11800 3723
rect 11926 3689 11978 3723
rect 12104 3689 12156 3723
rect 12282 3689 12334 3723
rect 12460 3689 12512 3723
rect 12638 3689 12690 3723
rect 508 3489 560 3523
rect 686 3489 738 3523
rect 864 3489 916 3523
rect 1042 3489 1094 3523
rect 1220 3489 1272 3523
rect 1398 3489 1450 3523
rect 1576 3489 1628 3523
rect 1754 3489 1806 3523
rect 1932 3489 1984 3523
rect 2110 3489 2162 3523
rect 2288 3489 2340 3523
rect 2466 3489 2518 3523
rect 2644 3489 2696 3523
rect 2822 3489 2874 3523
rect 3000 3489 3052 3523
rect 3178 3489 3230 3523
rect 3356 3489 3408 3523
rect 3534 3489 3586 3523
rect 3908 3489 3960 3523
rect 4086 3489 4138 3523
rect 4264 3489 4316 3523
rect 4442 3489 4494 3523
rect 4620 3489 4672 3523
rect 4798 3489 4850 3523
rect 4976 3489 5028 3523
rect 5154 3489 5206 3523
rect 5332 3489 5384 3523
rect 5510 3489 5562 3523
rect 5688 3489 5740 3523
rect 5866 3489 5918 3523
rect 6044 3489 6096 3523
rect 6222 3489 6274 3523
rect 6400 3489 6452 3523
rect 6578 3489 6630 3523
rect 6756 3489 6808 3523
rect 6934 3489 6986 3523
rect 7637 3299 7689 3333
rect 7815 3299 7867 3333
rect 7993 3299 8045 3333
rect 8171 3299 8223 3333
rect 8349 3299 8401 3333
rect 8527 3299 8579 3333
rect 8705 3299 8757 3333
rect 8883 3299 8935 3333
rect 9061 3299 9113 3333
rect 9239 3299 9291 3333
rect 9417 3299 9469 3333
rect 9595 3299 9647 3333
rect 9773 3299 9825 3333
rect 9951 3299 10003 3333
rect 10324 3299 10376 3333
rect 10502 3299 10554 3333
rect 10680 3299 10732 3333
rect 10858 3299 10910 3333
rect 11036 3299 11088 3333
rect 11214 3299 11266 3333
rect 11392 3299 11444 3333
rect 11570 3299 11622 3333
rect 11748 3299 11800 3333
rect 11926 3299 11978 3333
rect 12104 3299 12156 3333
rect 12282 3299 12334 3333
rect 12460 3299 12512 3333
rect 12638 3299 12690 3333
rect 7637 3189 7689 3223
rect 508 3099 560 3133
rect 686 3099 738 3133
rect 864 3099 916 3133
rect 1042 3099 1094 3133
rect 1220 3099 1272 3133
rect 1398 3099 1450 3133
rect 1576 3099 1628 3133
rect 1754 3099 1806 3133
rect 1932 3099 1984 3133
rect 2110 3099 2162 3133
rect 2288 3099 2340 3133
rect 2466 3099 2518 3133
rect 2644 3099 2696 3133
rect 2822 3099 2874 3133
rect 3000 3099 3052 3133
rect 3178 3099 3230 3133
rect 3356 3099 3408 3133
rect 3534 3099 3586 3133
rect 3908 3099 3960 3133
rect 4086 3099 4138 3133
rect 4264 3099 4316 3133
rect 4442 3099 4494 3133
rect 4620 3099 4672 3133
rect 4798 3099 4850 3133
rect 4976 3099 5028 3133
rect 5154 3099 5206 3133
rect 5332 3099 5384 3133
rect 5510 3099 5562 3133
rect 5688 3099 5740 3133
rect 5866 3099 5918 3133
rect 6044 3099 6096 3133
rect 6222 3099 6274 3133
rect 6400 3099 6452 3133
rect 6578 3099 6630 3133
rect 6756 3099 6808 3133
rect 7815 3189 7867 3223
rect 7993 3189 8045 3223
rect 8171 3189 8223 3223
rect 8349 3189 8401 3223
rect 8527 3189 8579 3223
rect 8705 3189 8757 3223
rect 8883 3189 8935 3223
rect 9061 3189 9113 3223
rect 9239 3189 9291 3223
rect 9417 3189 9469 3223
rect 9595 3189 9647 3223
rect 9773 3189 9825 3223
rect 9951 3189 10003 3223
rect 10324 3189 10376 3223
rect 10502 3189 10554 3223
rect 10680 3189 10732 3223
rect 10858 3189 10910 3223
rect 11036 3189 11088 3223
rect 11214 3189 11266 3223
rect 11392 3189 11444 3223
rect 11570 3189 11622 3223
rect 11748 3189 11800 3223
rect 11926 3189 11978 3223
rect 12104 3189 12156 3223
rect 12282 3189 12334 3223
rect 12460 3189 12512 3223
rect 12638 3189 12690 3223
rect 6934 3099 6986 3133
rect 508 2989 560 3023
rect 686 2989 738 3023
rect 864 2989 916 3023
rect 1042 2989 1094 3023
rect 1220 2989 1272 3023
rect 1398 2989 1450 3023
rect 1576 2989 1628 3023
rect 1754 2989 1806 3023
rect 1932 2989 1984 3023
rect 2110 2989 2162 3023
rect 2288 2989 2340 3023
rect 2466 2989 2518 3023
rect 2644 2989 2696 3023
rect 2822 2989 2874 3023
rect 3000 2989 3052 3023
rect 3178 2989 3230 3023
rect 3356 2989 3408 3023
rect 3534 2989 3586 3023
rect 3908 2989 3960 3023
rect 4086 2989 4138 3023
rect 4264 2989 4316 3023
rect 4442 2989 4494 3023
rect 4620 2989 4672 3023
rect 4798 2989 4850 3023
rect 4976 2989 5028 3023
rect 5154 2989 5206 3023
rect 5332 2989 5384 3023
rect 5510 2989 5562 3023
rect 5688 2989 5740 3023
rect 5866 2989 5918 3023
rect 6044 2989 6096 3023
rect 6222 2989 6274 3023
rect 6400 2989 6452 3023
rect 6578 2989 6630 3023
rect 6756 2989 6808 3023
rect 6934 2989 6986 3023
rect 7637 2799 7689 2833
rect 7815 2799 7867 2833
rect 7993 2799 8045 2833
rect 8171 2799 8223 2833
rect 8349 2799 8401 2833
rect 8527 2799 8579 2833
rect 8705 2799 8757 2833
rect 8883 2799 8935 2833
rect 9061 2799 9113 2833
rect 9239 2799 9291 2833
rect 9417 2799 9469 2833
rect 9595 2799 9647 2833
rect 9773 2799 9825 2833
rect 9951 2799 10003 2833
rect 10324 2799 10376 2833
rect 10502 2799 10554 2833
rect 10680 2799 10732 2833
rect 10858 2799 10910 2833
rect 11036 2799 11088 2833
rect 11214 2799 11266 2833
rect 11392 2799 11444 2833
rect 11570 2799 11622 2833
rect 11748 2799 11800 2833
rect 11926 2799 11978 2833
rect 12104 2799 12156 2833
rect 12282 2799 12334 2833
rect 12460 2799 12512 2833
rect 12638 2799 12690 2833
rect 7637 2689 7689 2723
rect 508 2599 560 2633
rect 686 2599 738 2633
rect 864 2599 916 2633
rect 1042 2599 1094 2633
rect 1220 2599 1272 2633
rect 1398 2599 1450 2633
rect 1576 2599 1628 2633
rect 1754 2599 1806 2633
rect 1932 2599 1984 2633
rect 2110 2599 2162 2633
rect 2288 2599 2340 2633
rect 2466 2599 2518 2633
rect 2644 2599 2696 2633
rect 2822 2599 2874 2633
rect 3000 2599 3052 2633
rect 3178 2599 3230 2633
rect 3356 2599 3408 2633
rect 3534 2599 3586 2633
rect 3908 2599 3960 2633
rect 4086 2599 4138 2633
rect 4264 2599 4316 2633
rect 4442 2599 4494 2633
rect 4620 2599 4672 2633
rect 4798 2599 4850 2633
rect 4976 2599 5028 2633
rect 5154 2599 5206 2633
rect 5332 2599 5384 2633
rect 5510 2599 5562 2633
rect 5688 2599 5740 2633
rect 5866 2599 5918 2633
rect 6044 2599 6096 2633
rect 6222 2599 6274 2633
rect 6400 2599 6452 2633
rect 6578 2599 6630 2633
rect 6756 2599 6808 2633
rect 7815 2689 7867 2723
rect 7993 2689 8045 2723
rect 8171 2689 8223 2723
rect 8349 2689 8401 2723
rect 8527 2689 8579 2723
rect 8705 2689 8757 2723
rect 8883 2689 8935 2723
rect 9061 2689 9113 2723
rect 9239 2689 9291 2723
rect 9417 2689 9469 2723
rect 9595 2689 9647 2723
rect 9773 2689 9825 2723
rect 9951 2689 10003 2723
rect 10324 2689 10376 2723
rect 10502 2689 10554 2723
rect 10680 2689 10732 2723
rect 10858 2689 10910 2723
rect 11036 2689 11088 2723
rect 11214 2689 11266 2723
rect 11392 2689 11444 2723
rect 11570 2689 11622 2723
rect 11748 2689 11800 2723
rect 11926 2689 11978 2723
rect 12104 2689 12156 2723
rect 12282 2689 12334 2723
rect 12460 2689 12512 2723
rect 12638 2689 12690 2723
rect 6934 2599 6986 2633
rect 508 2489 560 2523
rect 686 2489 738 2523
rect 864 2489 916 2523
rect 1042 2489 1094 2523
rect 1220 2489 1272 2523
rect 1398 2489 1450 2523
rect 1576 2489 1628 2523
rect 1754 2489 1806 2523
rect 1932 2489 1984 2523
rect 2110 2489 2162 2523
rect 2288 2489 2340 2523
rect 2466 2489 2518 2523
rect 2644 2489 2696 2523
rect 2822 2489 2874 2523
rect 3000 2489 3052 2523
rect 3178 2489 3230 2523
rect 3356 2489 3408 2523
rect 3534 2489 3586 2523
rect 3908 2489 3960 2523
rect 4086 2489 4138 2523
rect 4264 2489 4316 2523
rect 4442 2489 4494 2523
rect 4620 2489 4672 2523
rect 4798 2489 4850 2523
rect 4976 2489 5028 2523
rect 5154 2489 5206 2523
rect 5332 2489 5384 2523
rect 5510 2489 5562 2523
rect 5688 2489 5740 2523
rect 5866 2489 5918 2523
rect 6044 2489 6096 2523
rect 6222 2489 6274 2523
rect 6400 2489 6452 2523
rect 6578 2489 6630 2523
rect 6756 2489 6808 2523
rect 6934 2489 6986 2523
rect 7637 2299 7689 2333
rect 7815 2299 7867 2333
rect 7993 2299 8045 2333
rect 8171 2299 8223 2333
rect 8349 2299 8401 2333
rect 8527 2299 8579 2333
rect 8705 2299 8757 2333
rect 8883 2299 8935 2333
rect 9061 2299 9113 2333
rect 9239 2299 9291 2333
rect 9417 2299 9469 2333
rect 9595 2299 9647 2333
rect 9773 2299 9825 2333
rect 9951 2299 10003 2333
rect 10324 2299 10376 2333
rect 10502 2299 10554 2333
rect 10680 2299 10732 2333
rect 10858 2299 10910 2333
rect 11036 2299 11088 2333
rect 11214 2299 11266 2333
rect 11392 2299 11444 2333
rect 11570 2299 11622 2333
rect 11748 2299 11800 2333
rect 11926 2299 11978 2333
rect 12104 2299 12156 2333
rect 12282 2299 12334 2333
rect 12460 2299 12512 2333
rect 12638 2299 12690 2333
rect 508 2099 560 2133
rect 686 2099 738 2133
rect 864 2099 916 2133
rect 1042 2099 1094 2133
rect 1220 2099 1272 2133
rect 1398 2099 1450 2133
rect 1576 2099 1628 2133
rect 1754 2099 1806 2133
rect 1932 2099 1984 2133
rect 2110 2099 2162 2133
rect 2288 2099 2340 2133
rect 2466 2099 2518 2133
rect 2644 2099 2696 2133
rect 2822 2099 2874 2133
rect 3000 2099 3052 2133
rect 3178 2099 3230 2133
rect 3356 2099 3408 2133
rect 3534 2099 3586 2133
rect 3908 2099 3960 2133
rect 4086 2099 4138 2133
rect 4264 2099 4316 2133
rect 4442 2099 4494 2133
rect 4620 2099 4672 2133
rect 4798 2099 4850 2133
rect 4976 2099 5028 2133
rect 5154 2099 5206 2133
rect 5332 2099 5384 2133
rect 5510 2099 5562 2133
rect 5688 2099 5740 2133
rect 5866 2099 5918 2133
rect 6044 2099 6096 2133
rect 6222 2099 6274 2133
rect 6400 2099 6452 2133
rect 6578 2099 6630 2133
rect 6756 2099 6808 2133
rect 6934 2099 6986 2133
rect 508 1989 560 2023
rect 686 1989 738 2023
rect 864 1989 916 2023
rect 1042 1989 1094 2023
rect 1220 1989 1272 2023
rect 1398 1989 1450 2023
rect 1576 1989 1628 2023
rect 1754 1989 1806 2023
rect 1932 1989 1984 2023
rect 2110 1989 2162 2023
rect 2288 1989 2340 2023
rect 2466 1989 2518 2023
rect 2644 1989 2696 2023
rect 2822 1989 2874 2023
rect 3000 1989 3052 2023
rect 3178 1989 3230 2023
rect 3356 1989 3408 2023
rect 3534 1989 3586 2023
rect 3908 1989 3960 2023
rect 4086 1989 4138 2023
rect 4264 1989 4316 2023
rect 4442 1989 4494 2023
rect 4620 1989 4672 2023
rect 4798 1989 4850 2023
rect 4976 1989 5028 2023
rect 5154 1989 5206 2023
rect 5332 1989 5384 2023
rect 5510 1989 5562 2023
rect 5688 1989 5740 2023
rect 5866 1989 5918 2023
rect 6044 1989 6096 2023
rect 6222 1989 6274 2023
rect 6400 1989 6452 2023
rect 6578 1989 6630 2023
rect 6756 1989 6808 2023
rect 6934 1989 6986 2023
rect 7637 1989 7689 2023
rect 7815 1989 7867 2023
rect 7993 1989 8045 2023
rect 8171 1989 8223 2023
rect 8349 1989 8401 2023
rect 8527 1989 8579 2023
rect 8705 1989 8757 2023
rect 8883 1989 8935 2023
rect 9061 1989 9113 2023
rect 9239 1989 9291 2023
rect 9417 1989 9469 2023
rect 9595 1989 9647 2023
rect 9773 1989 9825 2023
rect 9951 1989 10003 2023
rect 10324 1989 10376 2023
rect 10502 1989 10554 2023
rect 10680 1989 10732 2023
rect 10858 1989 10910 2023
rect 11036 1989 11088 2023
rect 11214 1989 11266 2023
rect 11392 1989 11444 2023
rect 11570 1989 11622 2023
rect 11748 1989 11800 2023
rect 11926 1989 11978 2023
rect 12104 1989 12156 2023
rect 12282 1989 12334 2023
rect 12460 1989 12512 2023
rect 12638 1989 12690 2023
rect 508 1599 560 1633
rect 686 1599 738 1633
rect 864 1599 916 1633
rect 1042 1599 1094 1633
rect 1220 1599 1272 1633
rect 1398 1599 1450 1633
rect 1576 1599 1628 1633
rect 1754 1599 1806 1633
rect 1932 1599 1984 1633
rect 2110 1599 2162 1633
rect 2288 1599 2340 1633
rect 2466 1599 2518 1633
rect 2644 1599 2696 1633
rect 2822 1599 2874 1633
rect 3000 1599 3052 1633
rect 3178 1599 3230 1633
rect 3356 1599 3408 1633
rect 3534 1599 3586 1633
rect 3908 1599 3960 1633
rect 4086 1599 4138 1633
rect 4264 1599 4316 1633
rect 4442 1599 4494 1633
rect 4620 1599 4672 1633
rect 4798 1599 4850 1633
rect 4976 1599 5028 1633
rect 5154 1599 5206 1633
rect 5332 1599 5384 1633
rect 5510 1599 5562 1633
rect 5688 1599 5740 1633
rect 5866 1599 5918 1633
rect 6044 1599 6096 1633
rect 6222 1599 6274 1633
rect 6400 1599 6452 1633
rect 6578 1599 6630 1633
rect 6756 1599 6808 1633
rect 6934 1599 6986 1633
rect 7637 1599 7689 1633
rect 7815 1599 7867 1633
rect 7993 1599 8045 1633
rect 8171 1599 8223 1633
rect 8349 1599 8401 1633
rect 8527 1599 8579 1633
rect 8705 1599 8757 1633
rect 8883 1599 8935 1633
rect 9061 1599 9113 1633
rect 9239 1599 9291 1633
rect 9417 1599 9469 1633
rect 9595 1599 9647 1633
rect 9773 1599 9825 1633
rect 9951 1599 10003 1633
rect 10324 1599 10376 1633
rect 10502 1599 10554 1633
rect 10680 1599 10732 1633
rect 10858 1599 10910 1633
rect 11036 1599 11088 1633
rect 11214 1599 11266 1633
rect 11392 1599 11444 1633
rect 11570 1599 11622 1633
rect 11748 1599 11800 1633
rect 11926 1599 11978 1633
rect 12104 1599 12156 1633
rect 12282 1599 12334 1633
rect 12460 1599 12512 1633
rect 12638 1599 12690 1633
rect 508 1489 560 1523
rect 686 1489 738 1523
rect 864 1489 916 1523
rect 1042 1489 1094 1523
rect 1220 1489 1272 1523
rect 1398 1489 1450 1523
rect 1576 1489 1628 1523
rect 1754 1489 1806 1523
rect 1932 1489 1984 1523
rect 2110 1489 2162 1523
rect 2288 1489 2340 1523
rect 2466 1489 2518 1523
rect 2644 1489 2696 1523
rect 2822 1489 2874 1523
rect 3000 1489 3052 1523
rect 3178 1489 3230 1523
rect 3356 1489 3408 1523
rect 3534 1489 3586 1523
rect 3908 1489 3960 1523
rect 4086 1489 4138 1523
rect 4264 1489 4316 1523
rect 4442 1489 4494 1523
rect 4620 1489 4672 1523
rect 4798 1489 4850 1523
rect 4976 1489 5028 1523
rect 5154 1489 5206 1523
rect 5332 1489 5384 1523
rect 5510 1489 5562 1523
rect 5688 1489 5740 1523
rect 5866 1489 5918 1523
rect 6044 1489 6096 1523
rect 6222 1489 6274 1523
rect 6400 1489 6452 1523
rect 6578 1489 6630 1523
rect 6756 1489 6808 1523
rect 6934 1489 6986 1523
rect 7637 1489 7689 1523
rect 7815 1489 7867 1523
rect 7993 1489 8045 1523
rect 8171 1489 8223 1523
rect 8349 1489 8401 1523
rect 8527 1489 8579 1523
rect 8705 1489 8757 1523
rect 8883 1489 8935 1523
rect 9061 1489 9113 1523
rect 9239 1489 9291 1523
rect 9417 1489 9469 1523
rect 9595 1489 9647 1523
rect 9773 1489 9825 1523
rect 9951 1489 10003 1523
rect 10324 1489 10376 1523
rect 10502 1489 10554 1523
rect 10680 1489 10732 1523
rect 10858 1489 10910 1523
rect 11036 1489 11088 1523
rect 11214 1489 11266 1523
rect 11392 1489 11444 1523
rect 11570 1489 11622 1523
rect 11748 1489 11800 1523
rect 11926 1489 11978 1523
rect 12104 1489 12156 1523
rect 12282 1489 12334 1523
rect 12460 1489 12512 1523
rect 12638 1489 12690 1523
rect 508 1099 560 1133
rect 686 1099 738 1133
rect 864 1099 916 1133
rect 1042 1099 1094 1133
rect 1220 1099 1272 1133
rect 1398 1099 1450 1133
rect 1576 1099 1628 1133
rect 1754 1099 1806 1133
rect 1932 1099 1984 1133
rect 2110 1099 2162 1133
rect 2288 1099 2340 1133
rect 2466 1099 2518 1133
rect 2644 1099 2696 1133
rect 2822 1099 2874 1133
rect 3000 1099 3052 1133
rect 3178 1099 3230 1133
rect 3356 1099 3408 1133
rect 3534 1099 3586 1133
rect 3908 1099 3960 1133
rect 4086 1099 4138 1133
rect 4264 1099 4316 1133
rect 4442 1099 4494 1133
rect 4620 1099 4672 1133
rect 4798 1099 4850 1133
rect 4976 1099 5028 1133
rect 5154 1099 5206 1133
rect 5332 1099 5384 1133
rect 5510 1099 5562 1133
rect 5688 1099 5740 1133
rect 5866 1099 5918 1133
rect 6044 1099 6096 1133
rect 6222 1099 6274 1133
rect 6400 1099 6452 1133
rect 6578 1099 6630 1133
rect 6756 1099 6808 1133
rect 6934 1099 6986 1133
rect 7637 1099 7689 1133
rect 7815 1099 7867 1133
rect 7993 1099 8045 1133
rect 8171 1099 8223 1133
rect 8349 1099 8401 1133
rect 8527 1099 8579 1133
rect 8705 1099 8757 1133
rect 8883 1099 8935 1133
rect 9061 1099 9113 1133
rect 9239 1099 9291 1133
rect 9417 1099 9469 1133
rect 9595 1099 9647 1133
rect 9773 1099 9825 1133
rect 9951 1099 10003 1133
rect 10324 1099 10376 1133
rect 10502 1099 10554 1133
rect 10680 1099 10732 1133
rect 10858 1099 10910 1133
rect 11036 1099 11088 1133
rect 11214 1099 11266 1133
rect 11392 1099 11444 1133
rect 11570 1099 11622 1133
rect 11748 1099 11800 1133
rect 11926 1099 11978 1133
rect 12104 1099 12156 1133
rect 12282 1099 12334 1133
rect 12460 1099 12512 1133
rect 12638 1099 12690 1133
rect 508 989 560 1023
rect 686 989 738 1023
rect 864 989 916 1023
rect 1042 989 1094 1023
rect 1220 989 1272 1023
rect 1398 989 1450 1023
rect 1576 989 1628 1023
rect 1754 989 1806 1023
rect 1932 989 1984 1023
rect 2110 989 2162 1023
rect 2288 989 2340 1023
rect 2466 989 2518 1023
rect 2644 989 2696 1023
rect 2822 989 2874 1023
rect 3000 989 3052 1023
rect 3178 989 3230 1023
rect 3356 989 3408 1023
rect 3534 989 3586 1023
rect 3908 989 3960 1023
rect 4086 989 4138 1023
rect 4264 989 4316 1023
rect 4442 989 4494 1023
rect 4620 989 4672 1023
rect 4798 989 4850 1023
rect 4976 989 5028 1023
rect 5154 989 5206 1023
rect 5332 989 5384 1023
rect 5510 989 5562 1023
rect 5688 989 5740 1023
rect 5866 989 5918 1023
rect 6044 989 6096 1023
rect 6222 989 6274 1023
rect 6400 989 6452 1023
rect 6578 989 6630 1023
rect 6756 989 6808 1023
rect 6934 989 6986 1023
rect 7637 989 7689 1023
rect 7815 989 7867 1023
rect 7993 989 8045 1023
rect 8171 989 8223 1023
rect 8349 989 8401 1023
rect 8527 989 8579 1023
rect 8705 989 8757 1023
rect 8883 989 8935 1023
rect 9061 989 9113 1023
rect 9239 989 9291 1023
rect 9417 989 9469 1023
rect 9595 989 9647 1023
rect 9773 989 9825 1023
rect 9951 989 10003 1023
rect 10324 989 10376 1023
rect 10502 989 10554 1023
rect 10680 989 10732 1023
rect 10858 989 10910 1023
rect 11036 989 11088 1023
rect 11214 989 11266 1023
rect 11392 989 11444 1023
rect 11570 989 11622 1023
rect 11748 989 11800 1023
rect 11926 989 11978 1023
rect 12104 989 12156 1023
rect 12282 989 12334 1023
rect 12460 989 12512 1023
rect 12638 989 12690 1023
rect 508 599 560 633
rect 686 599 738 633
rect 864 599 916 633
rect 1042 599 1094 633
rect 1220 599 1272 633
rect 1398 599 1450 633
rect 1576 599 1628 633
rect 1754 599 1806 633
rect 1932 599 1984 633
rect 2110 599 2162 633
rect 2288 599 2340 633
rect 2466 599 2518 633
rect 2644 599 2696 633
rect 2822 599 2874 633
rect 3000 599 3052 633
rect 3178 599 3230 633
rect 3356 599 3408 633
rect 3534 599 3586 633
rect 3908 599 3960 633
rect 4086 599 4138 633
rect 4264 599 4316 633
rect 4442 599 4494 633
rect 4620 599 4672 633
rect 4798 599 4850 633
rect 4976 599 5028 633
rect 5154 599 5206 633
rect 5332 599 5384 633
rect 5510 599 5562 633
rect 5688 599 5740 633
rect 5866 599 5918 633
rect 6044 599 6096 633
rect 6222 599 6274 633
rect 6400 599 6452 633
rect 6578 599 6630 633
rect 6756 599 6808 633
rect 6934 599 6986 633
rect 7637 599 7689 633
rect 7815 599 7867 633
rect 7993 599 8045 633
rect 8171 599 8223 633
rect 8349 599 8401 633
rect 8527 599 8579 633
rect 8705 599 8757 633
rect 8883 599 8935 633
rect 9061 599 9113 633
rect 9239 599 9291 633
rect 9417 599 9469 633
rect 9595 599 9647 633
rect 9773 599 9825 633
rect 9951 599 10003 633
rect 10324 599 10376 633
rect 10502 599 10554 633
rect 10680 599 10732 633
rect 10858 599 10910 633
rect 11036 599 11088 633
rect 11214 599 11266 633
rect 11392 599 11444 633
rect 11570 599 11622 633
rect 11748 599 11800 633
rect 11926 599 11978 633
rect 12104 599 12156 633
rect 12282 599 12334 633
rect 12460 599 12512 633
rect 12638 599 12690 633
rect 13630 5097 13682 5131
rect 13808 5097 13860 5131
rect 13986 5097 14038 5131
rect 14164 5097 14216 5131
rect 14342 5097 14394 5131
rect 14520 5097 14572 5131
rect 14698 5097 14750 5131
rect 14876 5097 14928 5131
rect 15054 5097 15106 5131
rect 15232 5097 15284 5131
rect 15410 5097 15462 5131
rect 15588 5097 15640 5131
rect 15766 5097 15818 5131
rect 15944 5097 15996 5131
rect 16122 5097 16174 5131
rect 16300 5097 16352 5131
rect 16478 5097 16530 5131
rect 16656 5097 16708 5131
rect 16834 5097 16886 5131
rect 17012 5097 17064 5131
rect 17190 5097 17242 5131
rect 17368 5097 17420 5131
rect 17546 5097 17598 5131
rect 17724 5097 17776 5131
rect 17902 5097 17954 5131
rect 18080 5097 18132 5131
rect 18258 5097 18310 5131
rect 13630 4707 13682 4741
rect 13808 4707 13860 4741
rect 13986 4707 14038 4741
rect 14164 4707 14216 4741
rect 14342 4707 14394 4741
rect 14520 4707 14572 4741
rect 14698 4707 14750 4741
rect 14876 4707 14928 4741
rect 15054 4707 15106 4741
rect 15232 4707 15284 4741
rect 15410 4707 15462 4741
rect 15588 4707 15640 4741
rect 15766 4707 15818 4741
rect 15944 4707 15996 4741
rect 16122 4707 16174 4741
rect 16300 4707 16352 4741
rect 16478 4707 16530 4741
rect 16656 4707 16708 4741
rect 16834 4707 16886 4741
rect 17012 4707 17064 4741
rect 17190 4707 17242 4741
rect 17368 4707 17420 4741
rect 17546 4707 17598 4741
rect 17724 4707 17776 4741
rect 17902 4707 17954 4741
rect 18080 4707 18132 4741
rect 18258 4707 18310 4741
rect 13630 4597 13682 4631
rect 13808 4597 13860 4631
rect 13986 4597 14038 4631
rect 14164 4597 14216 4631
rect 14342 4597 14394 4631
rect 14520 4597 14572 4631
rect 14698 4597 14750 4631
rect 14876 4597 14928 4631
rect 15054 4597 15106 4631
rect 15232 4597 15284 4631
rect 15410 4597 15462 4631
rect 15588 4597 15640 4631
rect 15766 4597 15818 4631
rect 15944 4597 15996 4631
rect 16122 4597 16174 4631
rect 16300 4597 16352 4631
rect 16478 4597 16530 4631
rect 16656 4597 16708 4631
rect 16834 4597 16886 4631
rect 17012 4597 17064 4631
rect 17190 4597 17242 4631
rect 17368 4597 17420 4631
rect 17546 4597 17598 4631
rect 17724 4597 17776 4631
rect 17902 4597 17954 4631
rect 18080 4597 18132 4631
rect 18258 4597 18310 4631
rect 13630 4207 13682 4241
rect 13808 4207 13860 4241
rect 13986 4207 14038 4241
rect 14164 4207 14216 4241
rect 14342 4207 14394 4241
rect 14520 4207 14572 4241
rect 14698 4207 14750 4241
rect 14876 4207 14928 4241
rect 15054 4207 15106 4241
rect 15232 4207 15284 4241
rect 15410 4207 15462 4241
rect 15588 4207 15640 4241
rect 15766 4207 15818 4241
rect 15944 4207 15996 4241
rect 16122 4207 16174 4241
rect 16300 4207 16352 4241
rect 16478 4207 16530 4241
rect 16656 4207 16708 4241
rect 16834 4207 16886 4241
rect 17012 4207 17064 4241
rect 17190 4207 17242 4241
rect 17368 4207 17420 4241
rect 17546 4207 17598 4241
rect 17724 4207 17776 4241
rect 17902 4207 17954 4241
rect 18080 4207 18132 4241
rect 18258 4207 18310 4241
rect 17188 3593 17240 3627
rect 17366 3593 17418 3627
rect 17544 3593 17596 3627
rect 17722 3593 17774 3627
rect 17188 3203 17240 3237
rect 17366 3203 17418 3237
rect 17544 3203 17596 3237
rect 17722 3203 17774 3237
rect 16474 2654 16526 2688
rect 13756 2588 13808 2622
rect 14048 2588 14100 2622
rect 14340 2588 14392 2622
rect 14632 2588 14684 2622
rect 14924 2588 14976 2622
rect 15216 2588 15268 2622
rect 15508 2588 15560 2622
rect 16652 2654 16704 2688
rect 16830 2654 16882 2688
rect 17008 2654 17060 2688
rect 17186 2654 17238 2688
rect 17364 2654 17416 2688
rect 17542 2654 17594 2688
rect 17720 2654 17772 2688
rect 17898 2654 17950 2688
rect 18076 2654 18128 2688
rect 18254 2654 18306 2688
rect 13756 2198 13808 2232
rect 14048 2198 14100 2232
rect 14340 2198 14392 2232
rect 14632 2198 14684 2232
rect 14924 2198 14976 2232
rect 15216 2198 15268 2232
rect 16474 2264 16526 2298
rect 16652 2264 16704 2298
rect 16830 2264 16882 2298
rect 17008 2264 17060 2298
rect 17186 2264 17238 2298
rect 17364 2264 17416 2298
rect 17542 2264 17594 2298
rect 17720 2264 17772 2298
rect 17898 2264 17950 2298
rect 18076 2264 18128 2298
rect 18254 2264 18306 2298
rect 15508 2198 15560 2232
rect 16474 2154 16526 2188
rect 13756 2090 13808 2124
rect 14048 2090 14100 2124
rect 14340 2090 14392 2124
rect 14632 2090 14684 2124
rect 14924 2090 14976 2124
rect 15216 2090 15268 2124
rect 15508 2090 15560 2124
rect 16652 2154 16704 2188
rect 16830 2154 16882 2188
rect 17008 2154 17060 2188
rect 17186 2154 17238 2188
rect 17364 2154 17416 2188
rect 17542 2154 17594 2188
rect 17720 2154 17772 2188
rect 17898 2154 17950 2188
rect 18076 2154 18128 2188
rect 18254 2154 18306 2188
rect 13756 1700 13808 1734
rect 14048 1700 14100 1734
rect 14340 1700 14392 1734
rect 14632 1700 14684 1734
rect 14924 1700 14976 1734
rect 15216 1700 15268 1734
rect 16474 1764 16526 1798
rect 16652 1764 16704 1798
rect 16830 1764 16882 1798
rect 17008 1764 17060 1798
rect 17186 1764 17238 1798
rect 17364 1764 17416 1798
rect 17542 1764 17594 1798
rect 17720 1764 17772 1798
rect 17898 1764 17950 1798
rect 18076 1764 18128 1798
rect 18254 1764 18306 1798
rect 15508 1700 15560 1734
rect 13756 1592 13808 1626
rect 14048 1592 14100 1626
rect 14340 1592 14392 1626
rect 14632 1592 14684 1626
rect 14924 1592 14976 1626
rect 15216 1592 15268 1626
rect 15508 1592 15560 1626
rect 16474 1594 16526 1628
rect 16652 1594 16704 1628
rect 16830 1594 16882 1628
rect 17008 1594 17060 1628
rect 17186 1594 17238 1628
rect 17364 1594 17416 1628
rect 17542 1594 17594 1628
rect 17720 1594 17772 1628
rect 17898 1594 17950 1628
rect 18076 1594 18128 1628
rect 18254 1594 18306 1628
rect 13756 1202 13808 1236
rect 14048 1202 14100 1236
rect 14340 1202 14392 1236
rect 14632 1202 14684 1236
rect 14924 1202 14976 1236
rect 15216 1202 15268 1236
rect 15508 1202 15560 1236
rect 16474 1204 16526 1238
rect 16652 1204 16704 1238
rect 16830 1204 16882 1238
rect 17008 1204 17060 1238
rect 17186 1204 17238 1238
rect 17364 1204 17416 1238
rect 17542 1204 17594 1238
rect 17720 1204 17772 1238
rect 17898 1204 17950 1238
rect 18076 1204 18128 1238
rect 18254 1204 18306 1238
rect 13756 1094 13808 1128
rect 14048 1094 14100 1128
rect 14340 1094 14392 1128
rect 14632 1094 14684 1128
rect 14924 1094 14976 1128
rect 15216 1094 15268 1128
rect 15508 1094 15560 1128
rect 16474 1094 16526 1128
rect 16652 1094 16704 1128
rect 16830 1094 16882 1128
rect 17008 1094 17060 1128
rect 17186 1094 17238 1128
rect 17364 1094 17416 1128
rect 17542 1094 17594 1128
rect 17720 1094 17772 1128
rect 17898 1094 17950 1128
rect 18076 1094 18128 1128
rect 18254 1094 18306 1128
rect 13756 704 13808 738
rect 14048 704 14100 738
rect 14340 704 14392 738
rect 14632 704 14684 738
rect 14924 704 14976 738
rect 15216 704 15268 738
rect 15508 704 15560 738
rect 16474 704 16526 738
rect 16652 704 16704 738
rect 16830 704 16882 738
rect 17008 704 17060 738
rect 17186 704 17238 738
rect 17364 704 17416 738
rect 17542 704 17594 738
rect 17720 704 17772 738
rect 17898 704 17950 738
rect 18076 704 18128 738
rect 18254 704 18306 738
rect 19089 5088 19141 5122
rect 19267 5088 19319 5122
rect 19445 5088 19497 5122
rect 19623 5088 19675 5122
rect 19801 5088 19853 5122
rect 19979 5088 20031 5122
rect 20157 5088 20209 5122
rect 20335 5088 20387 5122
rect 20513 5088 20565 5122
rect 20691 5088 20743 5122
rect 20869 5088 20921 5122
rect 21047 5088 21099 5122
rect 21225 5088 21277 5122
rect 21403 5088 21455 5122
rect 21581 5088 21633 5122
rect 21759 5088 21811 5122
rect 19089 4698 19141 4732
rect 19267 4698 19319 4732
rect 19445 4698 19497 4732
rect 19623 4698 19675 4732
rect 19801 4698 19853 4732
rect 19979 4698 20031 4732
rect 20157 4698 20209 4732
rect 20335 4698 20387 4732
rect 20513 4698 20565 4732
rect 20691 4698 20743 4732
rect 20869 4698 20921 4732
rect 21047 4698 21099 4732
rect 21225 4698 21277 4732
rect 21403 4698 21455 4732
rect 21581 4698 21633 4732
rect 21759 4698 21811 4732
rect 19089 4590 19141 4624
rect 19267 4590 19319 4624
rect 19445 4590 19497 4624
rect 19623 4590 19675 4624
rect 19801 4590 19853 4624
rect 19979 4590 20031 4624
rect 20157 4590 20209 4624
rect 20335 4590 20387 4624
rect 20513 4590 20565 4624
rect 20691 4590 20743 4624
rect 20869 4590 20921 4624
rect 21047 4590 21099 4624
rect 21225 4590 21277 4624
rect 21403 4590 21455 4624
rect 21581 4590 21633 4624
rect 21759 4590 21811 4624
rect 19089 4200 19141 4234
rect 19267 4200 19319 4234
rect 19445 4200 19497 4234
rect 19623 4200 19675 4234
rect 19801 4200 19853 4234
rect 19979 4200 20031 4234
rect 20157 4200 20209 4234
rect 20335 4200 20387 4234
rect 20513 4200 20565 4234
rect 20691 4200 20743 4234
rect 20869 4200 20921 4234
rect 21047 4200 21099 4234
rect 21225 4200 21277 4234
rect 21403 4200 21455 4234
rect 21581 4200 21633 4234
rect 21759 4200 21811 4234
rect 19089 4092 19141 4126
rect 19267 4092 19319 4126
rect 19445 4092 19497 4126
rect 19623 4092 19675 4126
rect 19801 4092 19853 4126
rect 19979 4092 20031 4126
rect 20157 4092 20209 4126
rect 20335 4092 20387 4126
rect 20513 4092 20565 4126
rect 20691 4092 20743 4126
rect 20869 4092 20921 4126
rect 21047 4092 21099 4126
rect 21225 4092 21277 4126
rect 21403 4092 21455 4126
rect 21581 4092 21633 4126
rect 21759 4092 21811 4126
rect 19089 3702 19141 3736
rect 19267 3702 19319 3736
rect 19445 3702 19497 3736
rect 19623 3702 19675 3736
rect 19801 3702 19853 3736
rect 19979 3702 20031 3736
rect 20157 3702 20209 3736
rect 20335 3702 20387 3736
rect 20513 3702 20565 3736
rect 20691 3702 20743 3736
rect 20869 3702 20921 3736
rect 21047 3702 21099 3736
rect 21225 3702 21277 3736
rect 21403 3702 21455 3736
rect 21581 3702 21633 3736
rect 21759 3702 21811 3736
rect 19089 3594 19141 3628
rect 19267 3594 19319 3628
rect 19445 3594 19497 3628
rect 19623 3594 19675 3628
rect 19801 3594 19853 3628
rect 19979 3594 20031 3628
rect 20157 3594 20209 3628
rect 20335 3594 20387 3628
rect 20513 3594 20565 3628
rect 20691 3594 20743 3628
rect 20869 3594 20921 3628
rect 21047 3594 21099 3628
rect 21225 3594 21277 3628
rect 21403 3594 21455 3628
rect 21581 3594 21633 3628
rect 21759 3594 21811 3628
rect 19089 3204 19141 3238
rect 19267 3204 19319 3238
rect 19445 3204 19497 3238
rect 19623 3204 19675 3238
rect 19801 3204 19853 3238
rect 19979 3204 20031 3238
rect 20157 3204 20209 3238
rect 20335 3204 20387 3238
rect 20513 3204 20565 3238
rect 20691 3204 20743 3238
rect 20869 3204 20921 3238
rect 21047 3204 21099 3238
rect 21225 3204 21277 3238
rect 21403 3204 21455 3238
rect 21581 3204 21633 3238
rect 21759 3204 21811 3238
rect 19447 2580 19499 2614
rect 19625 2580 19677 2614
rect 19803 2580 19855 2614
rect 19981 2580 20033 2614
rect 20159 2580 20211 2614
rect 20337 2580 20389 2614
rect 20515 2580 20567 2614
rect 20693 2580 20745 2614
rect 20871 2580 20923 2614
rect 21049 2580 21101 2614
rect 21227 2580 21279 2614
rect 19447 2190 19499 2224
rect 19625 2190 19677 2224
rect 19803 2190 19855 2224
rect 19981 2190 20033 2224
rect 20159 2190 20211 2224
rect 20337 2190 20389 2224
rect 20515 2190 20567 2224
rect 20693 2190 20745 2224
rect 20871 2190 20923 2224
rect 21049 2190 21101 2224
rect 21227 2190 21279 2224
rect 19447 2082 19499 2116
rect 19625 2082 19677 2116
rect 19803 2082 19855 2116
rect 19981 2082 20033 2116
rect 20159 2082 20211 2116
rect 20337 2082 20389 2116
rect 20515 2082 20567 2116
rect 20693 2082 20745 2116
rect 20871 2082 20923 2116
rect 21049 2082 21101 2116
rect 21227 2082 21279 2116
rect 19447 1692 19499 1726
rect 19625 1692 19677 1726
rect 19803 1692 19855 1726
rect 19981 1692 20033 1726
rect 20159 1692 20211 1726
rect 20337 1692 20389 1726
rect 20515 1692 20567 1726
rect 20693 1692 20745 1726
rect 20871 1692 20923 1726
rect 21049 1692 21101 1726
rect 21227 1692 21279 1726
rect 19447 1584 19499 1618
rect 19625 1584 19677 1618
rect 19803 1584 19855 1618
rect 19981 1584 20033 1618
rect 20159 1584 20211 1618
rect 20337 1584 20389 1618
rect 20515 1584 20567 1618
rect 20693 1584 20745 1618
rect 20871 1584 20923 1618
rect 21049 1584 21101 1618
rect 21227 1584 21279 1618
rect 19447 1194 19499 1228
rect 19625 1194 19677 1228
rect 19803 1194 19855 1228
rect 19981 1194 20033 1228
rect 20159 1194 20211 1228
rect 20337 1194 20389 1228
rect 20515 1194 20567 1228
rect 20693 1194 20745 1228
rect 20871 1194 20923 1228
rect 21049 1194 21101 1228
rect 21227 1194 21279 1228
rect 19447 1086 19499 1120
rect 19625 1086 19677 1120
rect 19803 1086 19855 1120
rect 19981 1086 20033 1120
rect 20159 1086 20211 1120
rect 20337 1086 20389 1120
rect 20515 1086 20567 1120
rect 20693 1086 20745 1120
rect 20871 1086 20923 1120
rect 21049 1086 21101 1120
rect 21227 1086 21279 1120
rect 19447 696 19499 730
rect 19625 696 19677 730
rect 19803 696 19855 730
rect 19981 696 20033 730
rect 20159 696 20211 730
rect 20337 696 20389 730
rect 20515 696 20567 730
rect 20693 696 20745 730
rect 20871 696 20923 730
rect 21049 696 21101 730
rect 21227 696 21279 730
<< locali >>
rect 6609 19960 21840 20216
rect 6609 18784 6865 19960
rect 21584 19254 21840 19960
rect 8715 18998 19906 19254
rect 7189 18903 7285 18937
rect 8315 18903 8411 18937
rect 7189 18841 7223 18903
rect 6609 18528 7189 18784
rect 6609 16983 6865 18528
rect 7287 18835 8313 18843
rect 7287 18801 7303 18835
rect 7337 18801 7495 18835
rect 7529 18801 7687 18835
rect 7721 18801 7879 18835
rect 7913 18801 8071 18835
rect 8105 18801 8262 18835
rect 8297 18801 8313 18835
rect 7287 18793 8313 18801
rect 8377 18841 8411 18903
rect 7303 18741 7337 18757
rect 7303 18477 7337 18493
rect 7399 18741 7433 18757
rect 7399 18477 7433 18493
rect 7495 18741 7529 18757
rect 7495 18477 7529 18493
rect 7591 18741 7625 18757
rect 7591 18477 7625 18493
rect 7687 18741 7721 18757
rect 7687 18477 7721 18493
rect 7783 18741 7817 18757
rect 7783 18477 7817 18493
rect 7879 18741 7913 18757
rect 7879 18477 7913 18493
rect 7975 18741 8009 18757
rect 7975 18477 8009 18493
rect 8071 18741 8105 18757
rect 8071 18477 8105 18493
rect 8167 18741 8201 18757
rect 8167 18477 8201 18493
rect 8263 18741 8297 18757
rect 8263 18477 8297 18493
rect 7189 18393 7223 18455
rect 8377 18393 8411 18455
rect 7189 18359 7285 18393
rect 8315 18359 8411 18393
rect 7189 18253 7285 18287
rect 8315 18253 8411 18287
rect 7189 18191 7223 18253
rect 8377 18205 8411 18253
rect 8715 18205 8971 18998
rect 8377 18191 8971 18205
rect 7303 18163 7337 18179
rect 7303 18067 7337 18083
rect 7399 18163 7433 18179
rect 7399 18067 7433 18083
rect 7495 18163 7529 18179
rect 7495 18067 7529 18083
rect 7591 18163 7625 18179
rect 7591 18067 7625 18083
rect 7687 18163 7721 18179
rect 7687 18067 7721 18083
rect 7783 18163 7817 18179
rect 7783 18067 7817 18083
rect 7879 18163 7913 18179
rect 7879 18067 7913 18083
rect 7975 18163 8009 18179
rect 7975 18067 8009 18083
rect 8071 18163 8105 18179
rect 8071 18067 8105 18083
rect 8167 18163 8201 18179
rect 8167 18067 8201 18083
rect 8263 18163 8297 18179
rect 8263 18067 8297 18083
rect 7189 17931 7223 17993
rect 7287 18024 8313 18032
rect 7287 17989 7303 18024
rect 7337 17990 7495 18024
rect 7529 17990 7687 18024
rect 7721 17990 7879 18024
rect 7913 17990 8071 18024
rect 8105 17990 8263 18024
rect 8298 17990 8313 18024
rect 7337 17989 8313 17990
rect 7287 17982 8313 17989
rect 8411 17993 8971 18191
rect 8377 17949 8971 17993
rect 8377 17931 8411 17949
rect 7189 17897 7285 17931
rect 8315 17897 8411 17931
rect 7189 17103 7285 17137
rect 8315 17103 8411 17137
rect 7189 17041 7223 17103
rect 6609 16727 7189 16983
rect 6609 15188 6865 16727
rect 7287 17036 8313 17043
rect 7287 17001 7303 17036
rect 7337 17035 8313 17036
rect 7337 17001 7495 17035
rect 7529 17001 7687 17035
rect 7721 17001 7879 17035
rect 7913 17001 8071 17035
rect 8105 17001 8263 17035
rect 8297 17001 8313 17035
rect 7287 16993 8313 17001
rect 8377 17041 8411 17103
rect 7303 16941 7337 16957
rect 7303 16677 7337 16693
rect 7399 16941 7433 16957
rect 7399 16677 7433 16693
rect 7495 16941 7529 16957
rect 7495 16677 7529 16693
rect 7591 16941 7625 16957
rect 7591 16677 7625 16693
rect 7687 16941 7721 16957
rect 7687 16677 7721 16693
rect 7783 16941 7817 16957
rect 7783 16677 7817 16693
rect 7879 16941 7913 16957
rect 7879 16677 7913 16693
rect 7975 16941 8009 16957
rect 7975 16677 8009 16693
rect 8071 16941 8105 16957
rect 8071 16677 8105 16693
rect 8167 16941 8201 16957
rect 8167 16677 8201 16693
rect 8263 16941 8297 16957
rect 8263 16677 8297 16693
rect 7189 16593 7223 16655
rect 8377 16593 8411 16655
rect 7189 16559 7285 16593
rect 8315 16559 8411 16593
rect 7189 16453 7285 16487
rect 8315 16453 8411 16487
rect 7189 16391 7223 16453
rect 8377 16427 8411 16453
rect 8715 16427 8971 17949
rect 8377 16391 8971 16427
rect 7303 16363 7337 16379
rect 7303 16267 7337 16283
rect 7399 16363 7433 16379
rect 7399 16267 7433 16283
rect 7495 16363 7529 16379
rect 7495 16267 7529 16283
rect 7591 16363 7625 16379
rect 7591 16267 7625 16283
rect 7687 16363 7721 16379
rect 7687 16267 7721 16283
rect 7783 16363 7817 16379
rect 7783 16267 7817 16283
rect 7879 16363 7913 16379
rect 7879 16267 7913 16283
rect 7975 16363 8009 16379
rect 7975 16267 8009 16283
rect 8071 16363 8105 16379
rect 8071 16267 8105 16283
rect 8167 16363 8201 16379
rect 8167 16267 8201 16283
rect 8263 16363 8297 16379
rect 8263 16267 8297 16283
rect 7189 16131 7223 16193
rect 7287 16224 8313 16232
rect 7287 16190 7303 16224
rect 7337 16223 7495 16224
rect 7338 16190 7495 16223
rect 7529 16190 7687 16224
rect 7721 16190 7879 16224
rect 7913 16190 8071 16224
rect 8105 16223 8263 16224
rect 8105 16190 8261 16223
rect 8297 16190 8313 16224
rect 7287 16189 7304 16190
rect 7338 16189 8261 16190
rect 8295 16189 8313 16190
rect 7287 16182 8313 16189
rect 8411 16193 8971 16391
rect 8377 16171 8971 16193
rect 8377 16131 8411 16171
rect 7189 16097 7285 16131
rect 8315 16097 8411 16131
rect 7189 15303 7285 15337
rect 8315 15303 8411 15337
rect 7189 15241 7223 15303
rect 6609 14932 7189 15188
rect 6609 13387 6865 14932
rect 7287 15235 8313 15243
rect 7287 15201 7301 15235
rect 7337 15201 7495 15235
rect 7529 15201 7687 15235
rect 7721 15201 7879 15235
rect 7913 15201 8071 15235
rect 8105 15201 8263 15235
rect 8299 15201 8313 15235
rect 7287 15193 8313 15201
rect 8377 15241 8411 15303
rect 7303 15141 7337 15157
rect 7303 14877 7337 14893
rect 7399 15141 7433 15157
rect 7399 14877 7433 14893
rect 7495 15141 7529 15157
rect 7495 14877 7529 14893
rect 7591 15141 7625 15157
rect 7591 14877 7625 14893
rect 7687 15141 7721 15157
rect 7687 14877 7721 14893
rect 7783 15141 7817 15157
rect 7783 14877 7817 14893
rect 7879 15141 7913 15157
rect 7879 14877 7913 14893
rect 7975 15141 8009 15157
rect 7975 14877 8009 14893
rect 8071 15141 8105 15157
rect 8071 14877 8105 14893
rect 8167 15141 8201 15157
rect 8167 14877 8201 14893
rect 8263 15141 8297 15157
rect 8263 14877 8297 14893
rect 7189 14793 7223 14855
rect 8377 14793 8411 14855
rect 7189 14759 7285 14793
rect 8315 14759 8411 14793
rect 7189 14653 7285 14687
rect 8315 14653 8411 14687
rect 7189 14591 7223 14653
rect 8377 14629 8411 14653
rect 8715 14629 8971 16171
rect 8377 14591 8971 14629
rect 7303 14563 7337 14579
rect 7303 14467 7337 14483
rect 7399 14563 7433 14579
rect 7399 14467 7433 14483
rect 7495 14563 7529 14579
rect 7495 14467 7529 14483
rect 7591 14563 7625 14579
rect 7591 14467 7625 14483
rect 7687 14563 7721 14579
rect 7687 14467 7721 14483
rect 7783 14563 7817 14579
rect 7783 14467 7817 14483
rect 7879 14563 7913 14579
rect 7879 14467 7913 14483
rect 7975 14563 8009 14579
rect 7975 14467 8009 14483
rect 8071 14563 8105 14579
rect 8071 14467 8105 14483
rect 8167 14563 8201 14579
rect 8167 14467 8201 14483
rect 8263 14563 8297 14579
rect 8263 14467 8297 14483
rect 7189 14331 7223 14393
rect 7287 14424 8313 14432
rect 7287 14390 7303 14424
rect 7337 14423 7495 14424
rect 7338 14390 7495 14423
rect 7529 14390 7687 14424
rect 7721 14390 7879 14424
rect 7913 14390 8071 14424
rect 8105 14390 8263 14424
rect 8297 14390 8313 14424
rect 7287 14389 7304 14390
rect 7338 14389 8313 14390
rect 7287 14382 8313 14389
rect 8411 14393 8971 14591
rect 8377 14373 8971 14393
rect 8377 14331 8411 14373
rect 7189 14297 7285 14331
rect 8315 14297 8411 14331
rect 7189 13503 7285 13537
rect 8315 13503 8411 13537
rect 7189 13441 7223 13503
rect 6609 13131 7189 13387
rect 6609 11552 6865 13131
rect 7287 13436 8313 13443
rect 7287 13435 7304 13436
rect 7338 13435 8262 13436
rect 8296 13435 8313 13436
rect 7287 13401 7303 13435
rect 7338 13402 7495 13435
rect 7337 13401 7495 13402
rect 7529 13401 7687 13435
rect 7721 13401 7879 13435
rect 7913 13401 8071 13435
rect 8105 13402 8262 13435
rect 8105 13401 8263 13402
rect 8297 13401 8313 13435
rect 7287 13393 8313 13401
rect 8377 13441 8411 13503
rect 7303 13341 7337 13357
rect 7303 13077 7337 13093
rect 7399 13341 7433 13357
rect 7399 13077 7433 13093
rect 7495 13341 7529 13357
rect 7495 13077 7529 13093
rect 7591 13341 7625 13357
rect 7591 13077 7625 13093
rect 7687 13341 7721 13357
rect 7687 13077 7721 13093
rect 7783 13341 7817 13357
rect 7783 13077 7817 13093
rect 7879 13341 7913 13357
rect 7879 13077 7913 13093
rect 7975 13341 8009 13357
rect 7975 13077 8009 13093
rect 8071 13341 8105 13357
rect 8071 13077 8105 13093
rect 8167 13341 8201 13357
rect 8167 13077 8201 13093
rect 8263 13341 8297 13357
rect 8263 13077 8297 13093
rect 7189 12993 7223 13055
rect 8377 12993 8411 13055
rect 7189 12959 7285 12993
rect 8315 12959 8411 12993
rect 7189 12853 7285 12887
rect 8315 12853 8411 12887
rect 7189 12791 7223 12853
rect 8377 12828 8411 12853
rect 8715 12828 8971 14373
rect 8377 12791 8971 12828
rect 7303 12763 7337 12779
rect 7303 12667 7337 12683
rect 7399 12763 7433 12779
rect 7399 12667 7433 12683
rect 7495 12763 7529 12779
rect 7495 12667 7529 12683
rect 7591 12763 7625 12779
rect 7591 12667 7625 12683
rect 7687 12763 7721 12779
rect 7687 12667 7721 12683
rect 7783 12763 7817 12779
rect 7783 12667 7817 12683
rect 7879 12763 7913 12779
rect 7879 12667 7913 12683
rect 7975 12763 8009 12779
rect 7975 12667 8009 12683
rect 8071 12763 8105 12779
rect 8071 12667 8105 12683
rect 8167 12763 8201 12779
rect 8167 12667 8201 12683
rect 8263 12763 8297 12779
rect 8263 12667 8297 12683
rect 7189 12531 7223 12593
rect 7287 12624 8313 12632
rect 7287 12623 7303 12624
rect 7287 12589 7301 12623
rect 7337 12590 7495 12624
rect 7529 12590 7687 12624
rect 7721 12590 7879 12624
rect 7913 12590 8071 12624
rect 8105 12590 8263 12624
rect 8297 12623 8313 12624
rect 7335 12589 8264 12590
rect 8298 12589 8313 12623
rect 7287 12582 8313 12589
rect 8411 12593 8971 12791
rect 8377 12572 8971 12593
rect 8377 12531 8411 12572
rect 7189 12497 7285 12531
rect 8315 12497 8411 12531
rect 7189 11703 7285 11737
rect 8315 11703 8411 11737
rect 7189 11641 7223 11703
rect 6609 11296 7189 11552
rect 6609 9779 6865 11296
rect 7287 11636 8313 11643
rect 7287 11635 8262 11636
rect 8296 11635 8313 11636
rect 7287 11601 7301 11635
rect 7337 11601 7495 11635
rect 7529 11601 7687 11635
rect 7721 11601 7879 11635
rect 7913 11601 8071 11635
rect 8105 11602 8262 11635
rect 8105 11601 8263 11602
rect 8297 11601 8313 11635
rect 7287 11593 8313 11601
rect 8377 11641 8411 11703
rect 7303 11541 7337 11557
rect 7303 11277 7337 11293
rect 7399 11541 7433 11557
rect 7399 11277 7433 11293
rect 7495 11541 7529 11557
rect 7495 11277 7529 11293
rect 7591 11541 7625 11557
rect 7591 11277 7625 11293
rect 7687 11541 7721 11557
rect 7687 11277 7721 11293
rect 7783 11541 7817 11557
rect 7783 11277 7817 11293
rect 7879 11541 7913 11557
rect 7879 11277 7913 11293
rect 7975 11541 8009 11557
rect 7975 11277 8009 11293
rect 8071 11541 8105 11557
rect 8071 11277 8105 11293
rect 8167 11541 8201 11557
rect 8167 11277 8201 11293
rect 8263 11541 8297 11557
rect 8263 11277 8297 11293
rect 7189 11193 7223 11255
rect 8377 11193 8411 11255
rect 7189 11159 7285 11193
rect 8315 11159 8411 11193
rect 7189 11053 7285 11087
rect 8315 11053 8411 11087
rect 7189 10991 7223 11053
rect 8377 11019 8411 11053
rect 8715 11019 8971 12572
rect 8377 10991 8971 11019
rect 7303 10963 7337 10979
rect 7303 10867 7337 10883
rect 7399 10963 7433 10979
rect 7399 10867 7433 10883
rect 7495 10963 7529 10979
rect 7495 10867 7529 10883
rect 7591 10963 7625 10979
rect 7591 10867 7625 10883
rect 7687 10963 7721 10979
rect 7687 10867 7721 10883
rect 7783 10963 7817 10979
rect 7783 10867 7817 10883
rect 7879 10963 7913 10979
rect 7879 10867 7913 10883
rect 7975 10963 8009 10979
rect 7975 10867 8009 10883
rect 8071 10963 8105 10979
rect 8071 10867 8105 10883
rect 8167 10963 8201 10979
rect 8167 10867 8201 10883
rect 8263 10963 8297 10979
rect 8263 10867 8297 10883
rect 7189 10731 7223 10793
rect 7287 10824 8313 10832
rect 7287 10823 7303 10824
rect 7287 10789 7300 10823
rect 7337 10790 7495 10824
rect 7529 10790 7687 10824
rect 7721 10790 7879 10824
rect 7913 10790 8071 10824
rect 8105 10823 8263 10824
rect 8105 10790 8262 10823
rect 8297 10790 8313 10824
rect 7334 10789 8262 10790
rect 8296 10789 8313 10790
rect 7287 10782 8313 10789
rect 8411 10793 8971 10991
rect 8377 10763 8971 10793
rect 8377 10731 8411 10763
rect 7189 10697 7285 10731
rect 8315 10697 8411 10731
rect 7189 9903 7285 9937
rect 8315 9903 8411 9937
rect 7189 9841 7223 9903
rect 6609 9523 7189 9779
rect 6609 8868 6865 9523
rect 7287 9837 8313 9843
rect 7287 9835 8262 9837
rect 8296 9835 8313 9837
rect 7287 9834 7303 9835
rect 7287 9800 7302 9834
rect 7337 9801 7495 9835
rect 7529 9801 7687 9835
rect 7721 9801 7879 9835
rect 7913 9801 8071 9835
rect 8105 9803 8262 9835
rect 8105 9801 8263 9803
rect 8297 9801 8313 9835
rect 7336 9800 8313 9801
rect 7287 9793 8313 9800
rect 8377 9841 8411 9903
rect 7303 9741 7337 9757
rect 7303 9477 7337 9493
rect 7399 9741 7433 9757
rect 7399 9477 7433 9493
rect 7495 9741 7529 9757
rect 7495 9477 7529 9493
rect 7591 9741 7625 9757
rect 7591 9477 7625 9493
rect 7687 9741 7721 9757
rect 7687 9477 7721 9493
rect 7783 9741 7817 9757
rect 7783 9477 7817 9493
rect 7879 9741 7913 9757
rect 7879 9477 7913 9493
rect 7975 9741 8009 9757
rect 7975 9477 8009 9493
rect 8071 9741 8105 9757
rect 8071 9477 8105 9493
rect 8167 9741 8201 9757
rect 8167 9477 8201 9493
rect 8263 9741 8297 9757
rect 8263 9477 8297 9493
rect 7189 9393 7223 9455
rect 8377 9393 8411 9455
rect 7189 9359 7285 9393
rect 8315 9359 8411 9393
rect 7189 9253 7285 9287
rect 8315 9253 8411 9287
rect 7189 9191 7223 9253
rect 8377 9239 8411 9253
rect 8715 9239 8971 10763
rect 8377 9191 8971 9239
rect 7303 9163 7337 9179
rect 7303 9067 7337 9083
rect 7399 9163 7433 9179
rect 7399 9067 7433 9083
rect 7495 9163 7529 9179
rect 7495 9067 7529 9083
rect 7591 9163 7625 9179
rect 7591 9067 7625 9083
rect 7687 9163 7721 9179
rect 7687 9067 7721 9083
rect 7783 9163 7817 9179
rect 7783 9067 7817 9083
rect 7879 9163 7913 9179
rect 7879 9067 7913 9083
rect 7975 9163 8009 9179
rect 7975 9067 8009 9083
rect 8071 9163 8105 9179
rect 8071 9067 8105 9083
rect 8167 9163 8201 9179
rect 8167 9067 8201 9083
rect 8263 9163 8297 9179
rect 8263 9067 8297 9083
rect 7189 8931 7223 8993
rect 7287 9026 8313 9032
rect 7287 8990 7303 9026
rect 7337 9024 8260 9026
rect 8294 9024 8313 9026
rect 7337 8990 7495 9024
rect 7529 8990 7687 9024
rect 7721 8990 7879 9024
rect 7913 8990 8071 9024
rect 8105 8992 8260 9024
rect 8105 8990 8263 8992
rect 8297 8990 8313 9024
rect 7287 8982 8313 8990
rect 8411 9017 8971 9191
rect 8411 8993 8715 9017
rect 8377 8983 8715 8993
rect 8377 8931 8411 8983
rect 7189 8897 7285 8931
rect 8315 8897 8411 8931
rect 6609 8734 6868 8868
rect 19650 18221 19906 18998
rect 21581 18966 21840 19254
rect 20119 18903 20215 18937
rect 21245 18903 21341 18937
rect 20119 18841 20153 18903
rect 20217 18837 21243 18843
rect 20217 18803 20224 18837
rect 20258 18835 21243 18837
rect 20217 18801 20233 18803
rect 20267 18801 20425 18835
rect 20459 18801 20617 18835
rect 20651 18801 20809 18835
rect 20843 18801 21001 18835
rect 21035 18801 21192 18835
rect 21227 18801 21243 18835
rect 20217 18793 21243 18801
rect 21307 18841 21341 18903
rect 20233 18741 20267 18757
rect 20233 18477 20267 18493
rect 20329 18741 20363 18757
rect 20329 18477 20363 18493
rect 20425 18741 20459 18757
rect 20425 18477 20459 18493
rect 20521 18741 20555 18757
rect 20521 18477 20555 18493
rect 20617 18741 20651 18757
rect 20617 18477 20651 18493
rect 20713 18741 20747 18757
rect 20713 18477 20747 18493
rect 20809 18741 20843 18757
rect 20809 18477 20843 18493
rect 20905 18741 20939 18757
rect 20905 18477 20939 18493
rect 21001 18741 21035 18757
rect 21001 18477 21035 18493
rect 21097 18741 21131 18757
rect 21097 18477 21131 18493
rect 21193 18741 21227 18757
rect 21193 18477 21227 18493
rect 20119 18393 20153 18455
rect 21581 18777 21837 18966
rect 21341 18521 21837 18777
rect 21307 18393 21341 18455
rect 20119 18359 20215 18393
rect 21245 18359 21341 18393
rect 20119 18253 20215 18287
rect 21245 18253 21341 18287
rect 20119 18221 20153 18253
rect 19650 18191 20153 18221
rect 19650 17993 20119 18191
rect 21307 18191 21341 18253
rect 20233 18163 20267 18179
rect 20233 18067 20267 18083
rect 20329 18163 20363 18179
rect 20329 18067 20363 18083
rect 20425 18163 20459 18179
rect 20425 18067 20459 18083
rect 20521 18163 20555 18179
rect 20521 18067 20555 18083
rect 20617 18163 20651 18179
rect 20617 18067 20651 18083
rect 20713 18163 20747 18179
rect 20713 18067 20747 18083
rect 20809 18163 20843 18179
rect 20809 18067 20843 18083
rect 20905 18163 20939 18179
rect 20905 18067 20939 18083
rect 21001 18163 21035 18179
rect 21001 18067 21035 18083
rect 21097 18163 21131 18179
rect 21097 18067 21131 18083
rect 21193 18163 21227 18179
rect 21193 18067 21227 18083
rect 19650 17965 20153 17993
rect 20217 18026 21243 18032
rect 20217 18024 21196 18026
rect 20217 17990 20233 18024
rect 20267 17990 20425 18024
rect 20459 17990 20617 18024
rect 20651 17990 20809 18024
rect 20843 17990 21001 18024
rect 21035 17990 21193 18024
rect 21230 17992 21243 18026
rect 21227 17990 21243 17992
rect 20217 17982 21243 17990
rect 19650 16417 19906 17965
rect 20119 17931 20153 17965
rect 21307 17931 21341 17993
rect 20119 17897 20215 17931
rect 21245 17897 21341 17931
rect 20119 17103 20215 17137
rect 21245 17103 21341 17137
rect 20119 17041 20153 17103
rect 20217 17039 21243 17043
rect 20217 17005 20229 17039
rect 20263 17035 21243 17039
rect 20217 17001 20233 17005
rect 20267 17001 20425 17035
rect 20459 17001 20617 17035
rect 20651 17001 20809 17035
rect 20843 17001 21001 17035
rect 21035 17001 21193 17035
rect 21228 17001 21243 17035
rect 20217 16993 21243 17001
rect 21307 17041 21341 17103
rect 20233 16941 20267 16957
rect 20233 16677 20267 16693
rect 20329 16941 20363 16957
rect 20329 16677 20363 16693
rect 20425 16941 20459 16957
rect 20425 16677 20459 16693
rect 20521 16941 20555 16957
rect 20521 16677 20555 16693
rect 20617 16941 20651 16957
rect 20617 16677 20651 16693
rect 20713 16941 20747 16957
rect 20713 16677 20747 16693
rect 20809 16941 20843 16957
rect 20809 16677 20843 16693
rect 20905 16941 20939 16957
rect 20905 16677 20939 16693
rect 21001 16941 21035 16957
rect 21001 16677 21035 16693
rect 21097 16941 21131 16957
rect 21097 16677 21131 16693
rect 21193 16941 21227 16957
rect 21193 16677 21227 16693
rect 20119 16593 20153 16655
rect 21581 16994 21837 18521
rect 21341 16738 21837 16994
rect 21307 16593 21341 16655
rect 20119 16559 20215 16593
rect 21245 16559 21341 16593
rect 20119 16453 20215 16487
rect 21245 16453 21341 16487
rect 20119 16417 20153 16453
rect 19650 16391 20153 16417
rect 19650 16193 20119 16391
rect 21307 16391 21341 16453
rect 20233 16363 20267 16379
rect 20233 16267 20267 16283
rect 20329 16363 20363 16379
rect 20329 16267 20363 16283
rect 20425 16363 20459 16379
rect 20425 16267 20459 16283
rect 20521 16363 20555 16379
rect 20521 16267 20555 16283
rect 20617 16363 20651 16379
rect 20617 16267 20651 16283
rect 20713 16363 20747 16379
rect 20713 16267 20747 16283
rect 20809 16363 20843 16379
rect 20809 16267 20843 16283
rect 20905 16363 20939 16379
rect 20905 16267 20939 16283
rect 21001 16363 21035 16379
rect 21001 16267 21035 16283
rect 21097 16363 21131 16379
rect 21097 16267 21131 16283
rect 21193 16363 21227 16379
rect 21193 16267 21227 16283
rect 19650 16161 20153 16193
rect 20217 16228 21243 16232
rect 20217 16226 21194 16228
rect 20217 16192 20229 16226
rect 20263 16224 21194 16226
rect 20217 16190 20233 16192
rect 20267 16190 20425 16224
rect 20459 16190 20617 16224
rect 20651 16190 20809 16224
rect 20843 16190 21001 16224
rect 21035 16190 21193 16224
rect 21228 16194 21243 16228
rect 21227 16190 21243 16194
rect 20217 16182 21243 16190
rect 19650 14629 19906 16161
rect 20119 16131 20153 16161
rect 21307 16131 21341 16193
rect 20119 16097 20215 16131
rect 21245 16097 21341 16131
rect 20119 15303 20215 15337
rect 21245 15303 21341 15337
rect 20119 15241 20153 15303
rect 20217 15235 21243 15243
rect 20217 15201 20233 15235
rect 20269 15201 20425 15235
rect 20459 15201 20617 15235
rect 20651 15201 20809 15235
rect 20843 15201 21001 15235
rect 21035 15201 21193 15235
rect 21230 15201 21243 15235
rect 20217 15193 21243 15201
rect 21307 15241 21341 15303
rect 20233 15141 20267 15157
rect 20233 14877 20267 14893
rect 20329 15141 20363 15157
rect 20329 14877 20363 14893
rect 20425 15141 20459 15157
rect 20425 14877 20459 14893
rect 20521 15141 20555 15157
rect 20521 14877 20555 14893
rect 20617 15141 20651 15157
rect 20617 14877 20651 14893
rect 20713 15141 20747 15157
rect 20713 14877 20747 14893
rect 20809 15141 20843 15157
rect 20809 14877 20843 14893
rect 20905 15141 20939 15157
rect 20905 14877 20939 14893
rect 21001 15141 21035 15157
rect 21001 14877 21035 14893
rect 21097 15141 21131 15157
rect 21097 14877 21131 14893
rect 21193 15141 21227 15157
rect 21193 14877 21227 14893
rect 20119 14793 20153 14855
rect 21581 15180 21837 16738
rect 21341 14924 21837 15180
rect 21307 14793 21341 14855
rect 20119 14759 20215 14793
rect 21245 14759 21341 14793
rect 20119 14653 20215 14687
rect 21245 14653 21341 14687
rect 20119 14629 20153 14653
rect 19650 14591 20153 14629
rect 19650 14393 20119 14591
rect 21307 14591 21341 14653
rect 20233 14563 20267 14579
rect 20233 14467 20267 14483
rect 20329 14563 20363 14579
rect 20329 14467 20363 14483
rect 20425 14563 20459 14579
rect 20425 14467 20459 14483
rect 20521 14563 20555 14579
rect 20521 14467 20555 14483
rect 20617 14563 20651 14579
rect 20617 14467 20651 14483
rect 20713 14563 20747 14579
rect 20713 14467 20747 14483
rect 20809 14563 20843 14579
rect 20809 14467 20843 14483
rect 20905 14563 20939 14579
rect 20905 14467 20939 14483
rect 21001 14563 21035 14579
rect 21001 14467 21035 14483
rect 21097 14563 21131 14579
rect 21097 14467 21131 14483
rect 21193 14563 21227 14579
rect 21193 14467 21227 14483
rect 19650 14373 20153 14393
rect 20217 14426 21243 14432
rect 20217 14424 21200 14426
rect 20217 14422 20233 14424
rect 20217 14388 20231 14422
rect 20267 14390 20425 14424
rect 20459 14390 20617 14424
rect 20651 14390 20809 14424
rect 20843 14390 21001 14424
rect 21035 14390 21193 14424
rect 21234 14392 21243 14426
rect 21227 14390 21243 14392
rect 20265 14388 21243 14390
rect 20217 14382 21243 14388
rect 19650 12825 19906 14373
rect 20119 14331 20153 14373
rect 21307 14331 21341 14393
rect 20119 14297 20215 14331
rect 21245 14297 21341 14331
rect 20119 13503 20215 13537
rect 21245 13503 21341 13537
rect 20119 13441 20153 13503
rect 20217 13439 21243 13443
rect 20217 13405 20231 13439
rect 20265 13435 21192 13439
rect 21226 13435 21243 13439
rect 20217 13401 20233 13405
rect 20267 13401 20425 13435
rect 20459 13401 20617 13435
rect 20651 13401 20809 13435
rect 20843 13401 21001 13435
rect 21035 13405 21192 13435
rect 21035 13401 21193 13405
rect 21227 13401 21243 13435
rect 20217 13393 21243 13401
rect 21307 13441 21341 13503
rect 20233 13341 20267 13357
rect 20233 13077 20267 13093
rect 20329 13341 20363 13357
rect 20329 13077 20363 13093
rect 20425 13341 20459 13357
rect 20425 13077 20459 13093
rect 20521 13341 20555 13357
rect 20521 13077 20555 13093
rect 20617 13341 20651 13357
rect 20617 13077 20651 13093
rect 20713 13341 20747 13357
rect 20713 13077 20747 13093
rect 20809 13341 20843 13357
rect 20809 13077 20843 13093
rect 20905 13341 20939 13357
rect 20905 13077 20939 13093
rect 21001 13341 21035 13357
rect 21001 13077 21035 13093
rect 21097 13341 21131 13357
rect 21097 13077 21131 13093
rect 21193 13341 21227 13357
rect 21193 13077 21227 13093
rect 20119 12993 20153 13055
rect 21581 13379 21837 14924
rect 21341 13123 21837 13379
rect 21307 12993 21341 13055
rect 20119 12959 20215 12993
rect 21245 12959 21341 12993
rect 20119 12853 20215 12887
rect 21245 12853 21341 12887
rect 20119 12825 20153 12853
rect 19650 12791 20153 12825
rect 19650 12593 20119 12791
rect 21307 12791 21341 12853
rect 20233 12763 20267 12779
rect 20233 12667 20267 12683
rect 20329 12763 20363 12779
rect 20329 12667 20363 12683
rect 20425 12763 20459 12779
rect 20425 12667 20459 12683
rect 20521 12763 20555 12779
rect 20521 12667 20555 12683
rect 20617 12763 20651 12779
rect 20617 12667 20651 12683
rect 20713 12763 20747 12779
rect 20713 12667 20747 12683
rect 20809 12763 20843 12779
rect 20809 12667 20843 12683
rect 20905 12763 20939 12779
rect 20905 12667 20939 12683
rect 21001 12763 21035 12779
rect 21001 12667 21035 12683
rect 21097 12763 21131 12779
rect 21097 12667 21131 12683
rect 21193 12763 21227 12779
rect 21193 12667 21227 12683
rect 19650 12569 20153 12593
rect 20217 12624 21243 12632
rect 20217 12590 20229 12624
rect 20267 12590 20425 12624
rect 20459 12590 20617 12624
rect 20651 12590 20809 12624
rect 20843 12590 21001 12624
rect 21035 12590 21193 12624
rect 21227 12620 21243 12624
rect 20217 12586 21196 12590
rect 21230 12586 21243 12620
rect 20217 12582 21243 12586
rect 19650 11014 19906 12569
rect 20119 12531 20153 12569
rect 21307 12531 21341 12593
rect 20119 12497 20215 12531
rect 21245 12497 21341 12531
rect 20119 11703 20215 11737
rect 21245 11703 21341 11737
rect 20119 11641 20153 11703
rect 20217 11639 21243 11643
rect 20217 11605 20231 11639
rect 20265 11635 21243 11639
rect 20217 11601 20233 11605
rect 20267 11601 20425 11635
rect 20459 11601 20617 11635
rect 20651 11601 20809 11635
rect 20843 11601 21001 11635
rect 21035 11601 21193 11635
rect 21227 11633 21243 11635
rect 20217 11599 21196 11601
rect 21230 11599 21243 11633
rect 20217 11593 21243 11599
rect 21307 11641 21341 11703
rect 20233 11541 20267 11557
rect 20233 11277 20267 11293
rect 20329 11541 20363 11557
rect 20329 11277 20363 11293
rect 20425 11541 20459 11557
rect 20425 11277 20459 11293
rect 20521 11541 20555 11557
rect 20521 11277 20555 11293
rect 20617 11541 20651 11557
rect 20617 11277 20651 11293
rect 20713 11541 20747 11557
rect 20713 11277 20747 11293
rect 20809 11541 20843 11557
rect 20809 11277 20843 11293
rect 20905 11541 20939 11557
rect 20905 11277 20939 11293
rect 21001 11541 21035 11557
rect 21001 11277 21035 11293
rect 21097 11541 21131 11557
rect 21097 11277 21131 11293
rect 21193 11541 21227 11557
rect 21193 11277 21227 11293
rect 20119 11193 20153 11255
rect 21581 11580 21837 13123
rect 21341 11324 21837 11580
rect 21307 11193 21341 11255
rect 20119 11159 20215 11193
rect 21245 11159 21341 11193
rect 20119 11053 20215 11087
rect 21245 11053 21341 11087
rect 20119 11014 20153 11053
rect 19650 10991 20153 11014
rect 19650 10793 20119 10991
rect 21307 10991 21341 11053
rect 20233 10963 20267 10979
rect 20233 10867 20267 10883
rect 20329 10963 20363 10979
rect 20329 10867 20363 10883
rect 20425 10963 20459 10979
rect 20425 10867 20459 10883
rect 20521 10963 20555 10979
rect 20521 10867 20555 10883
rect 20617 10963 20651 10979
rect 20617 10867 20651 10883
rect 20713 10963 20747 10979
rect 20713 10867 20747 10883
rect 20809 10963 20843 10979
rect 20809 10867 20843 10883
rect 20905 10963 20939 10979
rect 20905 10867 20939 10883
rect 21001 10963 21035 10979
rect 21001 10867 21035 10883
rect 21097 10963 21131 10979
rect 21097 10867 21131 10883
rect 21193 10963 21227 10979
rect 21193 10867 21227 10883
rect 19650 10758 20153 10793
rect 20217 10824 21243 10832
rect 20217 10819 20233 10824
rect 20217 10785 20231 10819
rect 20267 10790 20425 10824
rect 20459 10790 20617 10824
rect 20651 10790 20809 10824
rect 20843 10790 21001 10824
rect 21035 10790 21190 10824
rect 21227 10790 21243 10824
rect 20265 10785 21243 10790
rect 20217 10782 21243 10785
rect 19650 9229 19906 10758
rect 20119 10731 20153 10758
rect 21307 10731 21341 10793
rect 20119 10697 20215 10731
rect 21245 10697 21341 10731
rect 20119 9903 20215 9937
rect 21245 9903 21341 9937
rect 20119 9841 20153 9903
rect 20217 9839 21243 9843
rect 20217 9835 21194 9839
rect 20217 9801 20233 9835
rect 20267 9801 20425 9835
rect 20459 9801 20617 9835
rect 20651 9801 20809 9835
rect 20843 9801 21001 9835
rect 21035 9801 21193 9835
rect 21228 9805 21243 9839
rect 21227 9801 21243 9805
rect 20217 9793 21243 9801
rect 21307 9841 21341 9903
rect 20233 9741 20267 9757
rect 20233 9477 20267 9493
rect 20329 9741 20363 9757
rect 20329 9477 20363 9493
rect 20425 9741 20459 9757
rect 20425 9477 20459 9493
rect 20521 9741 20555 9757
rect 20521 9477 20555 9493
rect 20617 9741 20651 9757
rect 20617 9477 20651 9493
rect 20713 9741 20747 9757
rect 20713 9477 20747 9493
rect 20809 9741 20843 9757
rect 20809 9477 20843 9493
rect 20905 9741 20939 9757
rect 20905 9477 20939 9493
rect 21001 9741 21035 9757
rect 21001 9477 21035 9493
rect 21097 9741 21131 9757
rect 21097 9477 21131 9493
rect 21193 9741 21227 9757
rect 21193 9477 21227 9493
rect 20119 9393 20153 9455
rect 21581 9795 21837 11324
rect 21341 9539 21837 9795
rect 21307 9393 21341 9455
rect 20119 9359 20215 9393
rect 21245 9359 21341 9393
rect 20119 9253 20215 9287
rect 21245 9253 21341 9287
rect 20119 9229 20153 9253
rect 19650 9191 20153 9229
rect 19650 9005 20119 9191
rect 8971 8761 19650 8990
rect 8715 8749 19650 8761
rect 19906 8993 20119 9005
rect 21307 9191 21341 9253
rect 20233 9163 20267 9179
rect 20233 9067 20267 9083
rect 20329 9163 20363 9179
rect 20329 9067 20363 9083
rect 20425 9163 20459 9179
rect 20425 9067 20459 9083
rect 20521 9163 20555 9179
rect 20521 9067 20555 9083
rect 20617 9163 20651 9179
rect 20617 9067 20651 9083
rect 20713 9163 20747 9179
rect 20713 9067 20747 9083
rect 20809 9163 20843 9179
rect 20809 9067 20843 9083
rect 20905 9163 20939 9179
rect 20905 9067 20939 9083
rect 21001 9163 21035 9179
rect 21001 9067 21035 9083
rect 21097 9163 21131 9179
rect 21097 9067 21131 9083
rect 21193 9163 21227 9179
rect 21193 9067 21227 9083
rect 19906 8973 20153 8993
rect 20217 9024 21243 9032
rect 20217 8990 20233 9024
rect 20267 9023 20425 9024
rect 20271 8990 20425 9023
rect 20459 8990 20617 9024
rect 20651 8990 20809 9024
rect 20843 8990 21001 9024
rect 21035 8990 21193 9024
rect 21227 9021 21243 9024
rect 20217 8989 20237 8990
rect 20271 8989 21196 8990
rect 20217 8987 21196 8989
rect 21230 8987 21243 9021
rect 20217 8982 21243 8987
rect 20119 8931 20153 8973
rect 21307 8931 21341 8993
rect 20119 8897 20215 8931
rect 21245 8897 21341 8931
rect 8715 8734 19906 8749
rect -61 8576 5805 8582
rect -61 8332 5555 8576
rect 5799 8332 5805 8576
rect -61 8326 5805 8332
rect -61 4649 195 8326
rect 6612 7996 6868 8734
rect 21581 7996 21837 9539
rect 6612 7740 21837 7996
rect 7193 7047 7449 7740
rect 11584 7047 11840 7740
rect 16315 7047 16571 7740
rect 21581 7047 21837 7740
rect 23491 8569 23747 8575
rect 23491 8325 23497 8569
rect 23741 8325 23747 8569
rect 7193 6991 22071 7047
rect 7193 6957 7445 6991
rect 14299 6957 14467 6991
rect 20872 6957 22071 6991
rect 7193 6919 22071 6957
rect 7193 6918 7575 6919
rect 7310 6852 7344 6918
rect -61 4600 272 4649
rect 6855 4600 6973 4649
rect -61 4548 210 4600
rect -61 149 161 4548
rect 1928 4303 2065 4600
rect 3649 4303 3843 4600
rect 1928 4269 2100 4303
rect 2134 4269 2182 4303
rect 2508 4269 2524 4303
rect 2558 4269 2574 4303
rect 2930 4269 2946 4303
rect 2980 4269 2996 4303
rect 3354 4269 3370 4303
rect 3404 4269 3420 4303
rect 3649 4269 3880 4303
rect 3914 4269 3962 4303
rect 4288 4269 4304 4303
rect 4338 4269 4354 4303
rect 4710 4269 4726 4303
rect 4760 4269 4776 4303
rect 5134 4269 5150 4303
rect 5184 4269 5200 4303
rect 1928 4219 2084 4269
rect 1928 4003 2050 4219
rect 1928 3987 2084 4003
rect 2148 4219 2182 4269
rect 3649 4235 3864 4269
rect 2148 3987 2182 4003
rect 2262 4219 2296 4235
rect 2262 3987 2296 4003
rect 2360 4219 2394 4235
rect 2360 3987 2394 4003
rect 2474 4219 2508 4235
rect 2474 3987 2508 4003
rect 2572 4219 2606 4235
rect 2572 3987 2606 4003
rect 2686 4219 2720 4235
rect 2686 3987 2720 4003
rect 2784 4219 2818 4235
rect 2784 3987 2818 4003
rect 2898 4219 2932 4235
rect 2898 3987 2932 4003
rect 2996 4219 3030 4235
rect 2996 3987 3030 4003
rect 3110 4219 3144 4235
rect 3110 3987 3144 4003
rect 3208 4219 3242 4235
rect 3208 3987 3242 4003
rect 3322 4219 3356 4235
rect 3322 3987 3356 4003
rect 3420 4219 3454 4235
rect 3420 3987 3454 4003
rect 3534 4219 3568 4235
rect 1928 3928 2065 3987
rect 3534 3953 3568 4003
rect 3632 4219 3864 4235
rect 3666 4003 3830 4219
rect 3632 3987 3864 4003
rect 3928 4219 3962 4269
rect 5436 4235 5573 4600
rect 3928 3987 3962 4003
rect 4042 4219 4076 4235
rect 4042 3987 4076 4003
rect 4140 4219 4174 4235
rect 4140 3987 4174 4003
rect 4254 4219 4288 4235
rect 4254 3987 4288 4003
rect 4352 4219 4386 4235
rect 4352 3987 4386 4003
rect 4466 4219 4500 4235
rect 4466 3987 4500 4003
rect 4564 4219 4598 4235
rect 4564 3987 4598 4003
rect 4678 4219 4712 4235
rect 4678 3987 4712 4003
rect 4776 4219 4810 4235
rect 4776 3987 4810 4003
rect 4890 4219 4924 4235
rect 4890 3987 4924 4003
rect 4988 4219 5022 4235
rect 4988 3987 5022 4003
rect 5102 4219 5136 4235
rect 5102 3987 5136 4003
rect 5200 4219 5234 4235
rect 5200 3987 5234 4003
rect 5314 4219 5348 4235
rect 3632 3953 3843 3987
rect 5314 3953 5348 4003
rect 5412 4219 5573 4235
rect 5446 4003 5573 4219
rect 5412 3953 5573 4003
rect 2296 3919 2312 3953
rect 2346 3919 2362 3953
rect 2720 3919 2736 3953
rect 2770 3919 2786 3953
rect 3142 3919 3158 3953
rect 3192 3919 3208 3953
rect 3534 3919 3582 3953
rect 3616 3919 3843 3953
rect 4076 3919 4092 3953
rect 4126 3919 4142 3953
rect 4500 3919 4516 3953
rect 4550 3919 4566 3953
rect 4922 3919 4938 3953
rect 4972 3919 4988 3953
rect 5314 3919 5362 3953
rect 5396 3919 5573 3953
rect 3649 3523 3843 3919
rect 5436 3909 5573 3919
rect 6924 4564 6973 4600
rect 7447 6690 7575 6918
rect 10053 6779 10258 6919
rect 10052 6690 10258 6779
rect 12746 6690 12874 6919
rect 7447 6656 7636 6690
rect 7688 6656 7704 6690
rect 7798 6656 7814 6690
rect 7866 6656 7882 6690
rect 7976 6656 7992 6690
rect 8044 6656 8060 6690
rect 8154 6656 8170 6690
rect 8222 6656 8238 6690
rect 8332 6656 8348 6690
rect 8400 6656 8416 6690
rect 8510 6656 8526 6690
rect 8578 6656 8594 6690
rect 8688 6656 8704 6690
rect 8756 6656 8772 6690
rect 8866 6656 8882 6690
rect 8934 6656 8950 6690
rect 9044 6656 9060 6690
rect 9112 6656 9128 6690
rect 9222 6656 9238 6690
rect 9290 6656 9306 6690
rect 9400 6656 9416 6690
rect 9468 6656 9484 6690
rect 9578 6656 9594 6690
rect 9646 6656 9662 6690
rect 9756 6656 9772 6690
rect 9824 6656 9840 6690
rect 9934 6656 9950 6690
rect 10002 6656 10322 6690
rect 10374 6656 10390 6690
rect 10484 6656 10500 6690
rect 10552 6656 10568 6690
rect 10662 6656 10678 6690
rect 10730 6656 10746 6690
rect 10840 6656 10856 6690
rect 10908 6656 10924 6690
rect 11018 6656 11034 6690
rect 11086 6656 11102 6690
rect 11196 6656 11212 6690
rect 11264 6656 11280 6690
rect 11374 6656 11390 6690
rect 11442 6656 11458 6690
rect 11552 6656 11568 6690
rect 11620 6656 11636 6690
rect 11730 6656 11746 6690
rect 11798 6656 11814 6690
rect 11908 6656 11924 6690
rect 11976 6656 11992 6690
rect 12086 6656 12102 6690
rect 12154 6656 12170 6690
rect 12264 6656 12280 6690
rect 12332 6656 12348 6690
rect 12442 6656 12458 6690
rect 12510 6656 12526 6690
rect 12620 6656 12636 6690
rect 12688 6656 12874 6690
rect 7447 6597 7590 6656
rect 7447 6341 7556 6597
rect 7447 6282 7590 6341
rect 7734 6597 7768 6613
rect 7734 6325 7768 6341
rect 7912 6597 7946 6613
rect 7912 6325 7946 6341
rect 8090 6597 8124 6613
rect 8090 6325 8124 6341
rect 8268 6597 8302 6613
rect 8268 6325 8302 6341
rect 8446 6597 8480 6613
rect 8446 6325 8480 6341
rect 8624 6597 8658 6613
rect 8624 6325 8658 6341
rect 8802 6597 8836 6613
rect 8802 6325 8836 6341
rect 8980 6597 9014 6613
rect 8980 6325 9014 6341
rect 9158 6597 9192 6613
rect 9158 6325 9192 6341
rect 9336 6597 9370 6613
rect 9336 6325 9370 6341
rect 9514 6597 9548 6613
rect 9514 6325 9548 6341
rect 9692 6597 9726 6613
rect 9692 6325 9726 6341
rect 9870 6597 9904 6613
rect 9870 6325 9904 6341
rect 10048 6597 10276 6656
rect 10082 6341 10242 6597
rect 10048 6282 10276 6341
rect 10420 6597 10454 6613
rect 10420 6325 10454 6341
rect 10598 6597 10632 6613
rect 10598 6325 10632 6341
rect 10776 6597 10810 6613
rect 10776 6325 10810 6341
rect 10954 6597 10988 6613
rect 10954 6325 10988 6341
rect 11132 6597 11166 6613
rect 11132 6325 11166 6341
rect 11310 6597 11344 6613
rect 11310 6325 11344 6341
rect 11488 6597 11522 6613
rect 11488 6325 11522 6341
rect 11666 6597 11700 6613
rect 11666 6325 11700 6341
rect 11844 6597 11878 6613
rect 11844 6325 11878 6341
rect 12022 6597 12056 6613
rect 12022 6325 12056 6341
rect 12200 6597 12234 6613
rect 12200 6325 12234 6341
rect 12378 6597 12412 6613
rect 12378 6325 12412 6341
rect 12556 6597 12590 6613
rect 12556 6325 12590 6341
rect 12734 6597 12874 6656
rect 12768 6341 12874 6597
rect 12734 6282 12874 6341
rect 7447 6248 7636 6282
rect 7688 6248 7704 6282
rect 7798 6248 7814 6282
rect 7866 6248 7882 6282
rect 7976 6248 7992 6282
rect 8044 6248 8060 6282
rect 8154 6248 8170 6282
rect 8222 6248 8238 6282
rect 8332 6248 8348 6282
rect 8400 6248 8416 6282
rect 8510 6248 8526 6282
rect 8578 6248 8594 6282
rect 8688 6248 8704 6282
rect 8756 6248 8772 6282
rect 8866 6248 8882 6282
rect 8934 6248 8950 6282
rect 9044 6248 9060 6282
rect 9112 6248 9128 6282
rect 9222 6248 9238 6282
rect 9290 6248 9306 6282
rect 9400 6248 9416 6282
rect 9468 6248 9484 6282
rect 9578 6248 9594 6282
rect 9646 6248 9662 6282
rect 9756 6248 9772 6282
rect 9824 6248 9840 6282
rect 9934 6248 9950 6282
rect 10002 6248 10322 6282
rect 10374 6248 10390 6282
rect 10484 6248 10500 6282
rect 10552 6248 10568 6282
rect 10662 6248 10678 6282
rect 10730 6248 10746 6282
rect 10840 6248 10856 6282
rect 10908 6248 10924 6282
rect 11018 6248 11034 6282
rect 11086 6248 11102 6282
rect 11196 6248 11212 6282
rect 11264 6248 11280 6282
rect 11374 6248 11390 6282
rect 11442 6248 11458 6282
rect 11552 6248 11568 6282
rect 11620 6248 11636 6282
rect 11730 6248 11746 6282
rect 11798 6248 11814 6282
rect 11908 6248 11924 6282
rect 11976 6248 11992 6282
rect 12086 6248 12102 6282
rect 12154 6248 12170 6282
rect 12264 6248 12280 6282
rect 12332 6248 12348 6282
rect 12442 6248 12458 6282
rect 12510 6248 12526 6282
rect 12620 6248 12636 6282
rect 12688 6248 12874 6282
rect 7447 6112 7575 6248
rect 10053 6113 10258 6248
rect 12746 6113 12874 6248
rect 10053 6112 10322 6113
rect 7447 6078 7636 6112
rect 7688 6078 7704 6112
rect 7798 6078 7814 6112
rect 7866 6078 7882 6112
rect 7976 6078 7992 6112
rect 8044 6078 8060 6112
rect 8154 6078 8170 6112
rect 8222 6078 8238 6112
rect 8332 6078 8348 6112
rect 8400 6078 8416 6112
rect 8510 6078 8526 6112
rect 8578 6078 8594 6112
rect 8688 6078 8704 6112
rect 8756 6078 8772 6112
rect 8866 6078 8882 6112
rect 8934 6078 8950 6112
rect 9044 6078 9060 6112
rect 9112 6078 9128 6112
rect 9222 6078 9238 6112
rect 9290 6078 9306 6112
rect 9400 6078 9416 6112
rect 9468 6078 9484 6112
rect 9578 6078 9594 6112
rect 9646 6078 9662 6112
rect 9756 6078 9772 6112
rect 9824 6078 9840 6112
rect 9934 6078 9950 6112
rect 10002 6079 10322 6112
rect 10374 6079 10390 6113
rect 10484 6079 10500 6113
rect 10552 6079 10568 6113
rect 10662 6079 10678 6113
rect 10730 6079 10746 6113
rect 10840 6079 10856 6113
rect 10908 6079 10924 6113
rect 11018 6079 11034 6113
rect 11086 6079 11102 6113
rect 11196 6079 11212 6113
rect 11264 6079 11280 6113
rect 11374 6079 11390 6113
rect 11442 6079 11458 6113
rect 11552 6079 11568 6113
rect 11620 6079 11636 6113
rect 11730 6079 11746 6113
rect 11798 6079 11814 6113
rect 11908 6079 11924 6113
rect 11976 6079 11992 6113
rect 12086 6079 12102 6113
rect 12154 6079 12170 6113
rect 12264 6079 12280 6113
rect 12332 6079 12348 6113
rect 12442 6079 12458 6113
rect 12510 6079 12526 6113
rect 12620 6079 12636 6113
rect 12688 6079 12874 6113
rect 10002 6078 10276 6079
rect 7447 6019 7590 6078
rect 7447 5763 7556 6019
rect 7447 5704 7590 5763
rect 7734 6019 7768 6035
rect 7734 5747 7768 5763
rect 7912 6019 7946 6035
rect 7912 5747 7946 5763
rect 8090 6019 8124 6035
rect 8090 5747 8124 5763
rect 8268 6019 8302 6035
rect 8268 5747 8302 5763
rect 8446 6019 8480 6035
rect 8446 5747 8480 5763
rect 8624 6019 8658 6035
rect 8624 5747 8658 5763
rect 8802 6019 8836 6035
rect 8802 5747 8836 5763
rect 8980 6019 9014 6035
rect 8980 5747 9014 5763
rect 9158 6019 9192 6035
rect 9158 5747 9192 5763
rect 9336 6019 9370 6035
rect 9336 5747 9370 5763
rect 9514 6019 9548 6035
rect 9514 5747 9548 5763
rect 9692 6019 9726 6035
rect 9692 5747 9726 5763
rect 9870 6019 9904 6035
rect 9870 5747 9904 5763
rect 10048 6020 10276 6078
rect 10048 6019 10242 6020
rect 10082 5764 10242 6019
rect 10082 5763 10276 5764
rect 10048 5705 10276 5763
rect 10420 6020 10454 6036
rect 10420 5748 10454 5764
rect 10598 6020 10632 6036
rect 10598 5748 10632 5764
rect 10776 6020 10810 6036
rect 10776 5748 10810 5764
rect 10954 6020 10988 6036
rect 10954 5748 10988 5764
rect 11132 6020 11166 6036
rect 11132 5748 11166 5764
rect 11310 6020 11344 6036
rect 11310 5748 11344 5764
rect 11488 6020 11522 6036
rect 11488 5748 11522 5764
rect 11666 6020 11700 6036
rect 11666 5748 11700 5764
rect 11844 6020 11878 6036
rect 11844 5748 11878 5764
rect 12022 6020 12056 6036
rect 12022 5748 12056 5764
rect 12200 6020 12234 6036
rect 12200 5748 12234 5764
rect 12378 6020 12412 6036
rect 12378 5748 12412 5764
rect 12556 6020 12590 6036
rect 12556 5748 12590 5764
rect 12734 6020 12874 6079
rect 12768 5764 12874 6020
rect 12734 5705 12874 5764
rect 10048 5704 10322 5705
rect 7447 5670 7636 5704
rect 7688 5670 7704 5704
rect 7798 5670 7814 5704
rect 7866 5670 7882 5704
rect 7976 5670 7992 5704
rect 8044 5670 8060 5704
rect 8154 5670 8170 5704
rect 8222 5670 8238 5704
rect 8332 5670 8348 5704
rect 8400 5670 8416 5704
rect 8510 5670 8526 5704
rect 8578 5670 8594 5704
rect 8688 5670 8704 5704
rect 8756 5670 8772 5704
rect 8866 5670 8882 5704
rect 8934 5670 8950 5704
rect 9044 5670 9060 5704
rect 9112 5670 9128 5704
rect 9222 5670 9238 5704
rect 9290 5670 9306 5704
rect 9400 5670 9416 5704
rect 9468 5670 9484 5704
rect 9578 5670 9594 5704
rect 9646 5670 9662 5704
rect 9756 5670 9772 5704
rect 9824 5670 9840 5704
rect 9934 5670 9950 5704
rect 10002 5671 10322 5704
rect 10374 5671 10390 5705
rect 10484 5671 10500 5705
rect 10552 5671 10568 5705
rect 10662 5671 10678 5705
rect 10730 5671 10746 5705
rect 10840 5671 10856 5705
rect 10908 5671 10924 5705
rect 11018 5671 11034 5705
rect 11086 5671 11102 5705
rect 11196 5671 11212 5705
rect 11264 5671 11280 5705
rect 11374 5671 11390 5705
rect 11442 5671 11458 5705
rect 11552 5671 11568 5705
rect 11620 5671 11636 5705
rect 11730 5671 11746 5705
rect 11798 5671 11814 5705
rect 11908 5671 11924 5705
rect 11976 5671 11992 5705
rect 12086 5671 12102 5705
rect 12154 5671 12170 5705
rect 12264 5671 12280 5705
rect 12332 5671 12348 5705
rect 12442 5671 12458 5705
rect 12510 5671 12526 5705
rect 12620 5671 12636 5705
rect 12688 5671 12874 5705
rect 10002 5670 10258 5671
rect 12746 5670 12874 5671
rect 14358 6892 14392 6919
rect 7447 5653 7575 5670
rect 10053 5232 10258 5670
rect 14603 6759 14731 6919
rect 16144 6759 16272 6919
rect 14603 6725 14776 6759
rect 14828 6725 14844 6759
rect 14938 6725 14954 6759
rect 15006 6725 15022 6759
rect 15116 6725 15132 6759
rect 15184 6725 15200 6759
rect 15294 6725 15310 6759
rect 15362 6725 15378 6759
rect 15472 6725 15488 6759
rect 15540 6725 15556 6759
rect 15650 6725 15666 6759
rect 15718 6725 15734 6759
rect 15828 6725 15844 6759
rect 15896 6725 15912 6759
rect 16006 6725 16022 6759
rect 16074 6725 16272 6759
rect 14603 6666 14731 6725
rect 14603 6410 14696 6666
rect 14730 6410 14731 6666
rect 14603 6351 14731 6410
rect 14874 6666 14908 6682
rect 14874 6394 14908 6410
rect 15052 6666 15086 6682
rect 15052 6394 15086 6410
rect 15230 6666 15264 6682
rect 15230 6394 15264 6410
rect 15408 6666 15442 6682
rect 15408 6394 15442 6410
rect 15586 6666 15620 6682
rect 15586 6394 15620 6410
rect 15764 6666 15798 6682
rect 15764 6394 15798 6410
rect 15942 6666 15976 6682
rect 15942 6394 15976 6410
rect 16120 6666 16272 6725
rect 16154 6410 16272 6666
rect 16120 6351 16272 6410
rect 14603 6317 14776 6351
rect 14828 6317 14844 6351
rect 14938 6317 14954 6351
rect 15006 6317 15022 6351
rect 15116 6317 15132 6351
rect 15184 6317 15200 6351
rect 15294 6317 15310 6351
rect 15362 6317 15378 6351
rect 15472 6317 15488 6351
rect 15540 6317 15556 6351
rect 15650 6317 15666 6351
rect 15718 6317 15734 6351
rect 15828 6317 15844 6351
rect 15896 6317 15912 6351
rect 16006 6317 16022 6351
rect 16074 6317 16272 6351
rect 14603 5992 14731 6317
rect 16144 5992 16272 6317
rect 14603 5958 14777 5992
rect 14829 5958 14845 5992
rect 14939 5958 14955 5992
rect 15007 5958 15023 5992
rect 15117 5958 15133 5992
rect 15185 5958 15201 5992
rect 15295 5958 15311 5992
rect 15363 5958 15379 5992
rect 15473 5958 15489 5992
rect 15541 5958 15557 5992
rect 15651 5958 15667 5992
rect 15719 5958 15735 5992
rect 15829 5958 15845 5992
rect 15897 5958 15913 5992
rect 16007 5958 16023 5992
rect 16075 5958 16272 5992
rect 14603 5899 14731 5958
rect 14603 5643 14697 5899
rect 14603 5584 14731 5643
rect 14875 5899 14909 5915
rect 14875 5627 14909 5643
rect 15053 5899 15087 5915
rect 15053 5627 15087 5643
rect 15231 5899 15265 5915
rect 15231 5627 15265 5643
rect 15409 5899 15443 5915
rect 15409 5627 15443 5643
rect 15587 5899 15621 5915
rect 15587 5627 15621 5643
rect 15765 5899 15799 5915
rect 15765 5627 15799 5643
rect 15943 5899 15977 5915
rect 15943 5627 15977 5643
rect 16121 5899 16272 5958
rect 16155 5643 16272 5899
rect 16121 5584 16272 5643
rect 14603 5553 14777 5584
rect 14697 5550 14777 5553
rect 14829 5550 14845 5584
rect 14939 5550 14955 5584
rect 15007 5550 15023 5584
rect 15117 5550 15133 5584
rect 15185 5550 15201 5584
rect 15295 5550 15311 5584
rect 15363 5550 15379 5584
rect 15473 5550 15489 5584
rect 15541 5550 15557 5584
rect 15651 5550 15667 5584
rect 15719 5550 15735 5584
rect 15829 5550 15845 5584
rect 15897 5550 15913 5584
rect 16007 5550 16023 5584
rect 16075 5556 16272 5584
rect 16796 6759 16924 6919
rect 18336 6759 18464 6919
rect 16796 6725 16976 6759
rect 17028 6725 17044 6759
rect 17138 6725 17154 6759
rect 17206 6725 17222 6759
rect 17316 6725 17332 6759
rect 17384 6725 17400 6759
rect 17494 6725 17510 6759
rect 17562 6725 17578 6759
rect 17672 6725 17688 6759
rect 17740 6725 17756 6759
rect 17850 6725 17866 6759
rect 17918 6725 17934 6759
rect 18028 6725 18044 6759
rect 18096 6725 18112 6759
rect 18206 6725 18222 6759
rect 18274 6725 18464 6759
rect 16796 6666 16930 6725
rect 16796 6410 16896 6666
rect 16796 6351 16930 6410
rect 17074 6666 17108 6682
rect 17074 6394 17108 6410
rect 17252 6666 17286 6682
rect 17252 6394 17286 6410
rect 17430 6666 17464 6682
rect 17430 6394 17464 6410
rect 17608 6666 17642 6682
rect 17608 6394 17642 6410
rect 17786 6666 17820 6682
rect 17786 6394 17820 6410
rect 17964 6666 17998 6682
rect 17964 6394 17998 6410
rect 18142 6666 18176 6682
rect 18142 6394 18176 6410
rect 18320 6666 18464 6725
rect 18354 6410 18464 6666
rect 18320 6351 18464 6410
rect 16796 6317 16976 6351
rect 17028 6317 17044 6351
rect 17138 6317 17154 6351
rect 17206 6317 17222 6351
rect 17316 6317 17332 6351
rect 17384 6317 17400 6351
rect 17494 6317 17510 6351
rect 17562 6317 17578 6351
rect 17672 6317 17688 6351
rect 17740 6317 17756 6351
rect 17850 6317 17866 6351
rect 17918 6317 17934 6351
rect 18028 6317 18044 6351
rect 18096 6317 18112 6351
rect 18206 6317 18222 6351
rect 18274 6317 18464 6351
rect 16796 5992 16924 6317
rect 18336 5992 18464 6317
rect 16796 5958 16977 5992
rect 17029 5958 17045 5992
rect 17139 5958 17155 5992
rect 17207 5958 17223 5992
rect 17317 5958 17333 5992
rect 17385 5958 17401 5992
rect 17495 5958 17511 5992
rect 17563 5958 17579 5992
rect 17673 5958 17689 5992
rect 17741 5958 17757 5992
rect 17851 5958 17867 5992
rect 17919 5958 17935 5992
rect 18029 5958 18045 5992
rect 18097 5958 18113 5992
rect 18207 5958 18223 5992
rect 18275 5958 18464 5992
rect 16796 5899 16931 5958
rect 16796 5643 16897 5899
rect 16796 5584 16931 5643
rect 17075 5899 17109 5915
rect 17075 5627 17109 5643
rect 17253 5899 17287 5915
rect 17253 5627 17287 5643
rect 17431 5899 17465 5915
rect 17431 5627 17465 5643
rect 17609 5899 17643 5915
rect 17609 5627 17643 5643
rect 17787 5899 17821 5915
rect 17787 5627 17821 5643
rect 17965 5899 17999 5915
rect 17965 5627 17999 5643
rect 18143 5899 18177 5915
rect 18143 5627 18177 5643
rect 18321 5899 18464 5958
rect 18355 5643 18464 5899
rect 18321 5584 18464 5643
rect 16075 5550 16155 5556
rect 16796 5550 16977 5584
rect 17029 5550 17045 5584
rect 17139 5550 17155 5584
rect 17207 5550 17223 5584
rect 17317 5550 17333 5584
rect 17385 5550 17401 5584
rect 17495 5550 17511 5584
rect 17563 5550 17579 5584
rect 17673 5550 17689 5584
rect 17741 5550 17757 5584
rect 17851 5550 17867 5584
rect 17919 5550 17935 5584
rect 18029 5550 18045 5584
rect 18097 5550 18113 5584
rect 18207 5550 18223 5584
rect 18275 5554 18464 5584
rect 18992 6759 19120 6919
rect 20541 6759 20669 6919
rect 18992 6725 19176 6759
rect 19228 6725 19244 6759
rect 19338 6725 19354 6759
rect 19406 6725 19422 6759
rect 19516 6725 19532 6759
rect 19584 6725 19600 6759
rect 19694 6725 19710 6759
rect 19762 6725 19778 6759
rect 19872 6725 19888 6759
rect 19940 6725 19956 6759
rect 20050 6725 20066 6759
rect 20118 6725 20134 6759
rect 20228 6725 20244 6759
rect 20296 6725 20312 6759
rect 20406 6725 20422 6759
rect 20474 6725 20669 6759
rect 18992 6666 19130 6725
rect 18992 6410 19096 6666
rect 18992 6351 19130 6410
rect 19274 6666 19308 6682
rect 19274 6394 19308 6410
rect 19452 6666 19486 6682
rect 19452 6394 19486 6410
rect 19630 6666 19664 6682
rect 19630 6394 19664 6410
rect 19808 6666 19842 6682
rect 19808 6394 19842 6410
rect 19986 6666 20020 6682
rect 19986 6394 20020 6410
rect 20164 6666 20198 6682
rect 20164 6394 20198 6410
rect 20342 6666 20376 6682
rect 20342 6394 20376 6410
rect 20520 6666 20669 6725
rect 20554 6410 20669 6666
rect 20520 6351 20669 6410
rect 18992 6317 19176 6351
rect 19228 6317 19244 6351
rect 19338 6317 19354 6351
rect 19406 6317 19422 6351
rect 19516 6317 19532 6351
rect 19584 6317 19600 6351
rect 19694 6317 19710 6351
rect 19762 6317 19778 6351
rect 19872 6317 19888 6351
rect 19940 6317 19956 6351
rect 20050 6317 20066 6351
rect 20118 6317 20134 6351
rect 20228 6317 20244 6351
rect 20296 6317 20312 6351
rect 20406 6317 20422 6351
rect 20474 6317 20669 6351
rect 18992 5992 19120 6317
rect 20541 5992 20669 6317
rect 18992 5958 19177 5992
rect 19229 5958 19245 5992
rect 19339 5958 19355 5992
rect 19407 5958 19423 5992
rect 19517 5958 19533 5992
rect 19585 5958 19601 5992
rect 19695 5958 19711 5992
rect 19763 5958 19779 5992
rect 19873 5958 19889 5992
rect 19941 5958 19957 5992
rect 20051 5958 20067 5992
rect 20119 5958 20135 5992
rect 20229 5958 20245 5992
rect 20297 5958 20313 5992
rect 20407 5958 20423 5992
rect 20475 5958 20669 5992
rect 18992 5899 19131 5958
rect 18992 5643 19097 5899
rect 18992 5584 19131 5643
rect 19275 5899 19309 5915
rect 19275 5627 19309 5643
rect 19453 5899 19487 5915
rect 19453 5627 19487 5643
rect 19631 5899 19665 5915
rect 19631 5627 19665 5643
rect 19809 5899 19843 5915
rect 19809 5627 19843 5643
rect 19987 5899 20021 5915
rect 19987 5627 20021 5643
rect 20165 5899 20199 5915
rect 20165 5627 20199 5643
rect 20343 5899 20377 5915
rect 20343 5627 20377 5643
rect 20521 5899 20669 5958
rect 20555 5643 20669 5899
rect 20521 5584 20669 5643
rect 18275 5550 18355 5554
rect 18992 5553 19177 5584
rect 19097 5550 19177 5553
rect 19229 5550 19245 5584
rect 19339 5550 19355 5584
rect 19407 5550 19423 5584
rect 19517 5550 19533 5584
rect 19585 5550 19601 5584
rect 19695 5550 19711 5584
rect 19763 5550 19779 5584
rect 19873 5550 19889 5584
rect 19941 5550 19957 5584
rect 20051 5550 20067 5584
rect 20119 5550 20135 5584
rect 20229 5550 20245 5584
rect 20297 5550 20313 5584
rect 20407 5550 20423 5584
rect 20475 5553 20669 5584
rect 20475 5550 20555 5553
rect 16796 5547 16924 5550
rect 14358 5413 14392 5525
rect 20943 5413 20977 5483
rect 12999 5379 13108 5413
rect 14264 5379 14464 5413
rect 20857 5379 20977 5413
rect 12999 5315 13033 5379
rect 12397 5232 12505 5240
rect 7912 5209 7992 5232
rect 7310 4124 7344 4198
rect 7805 5198 7992 5209
rect 8044 5198 8060 5232
rect 8154 5198 8170 5232
rect 8222 5198 8238 5232
rect 8332 5198 8348 5232
rect 8400 5198 8416 5232
rect 8510 5198 8526 5232
rect 8578 5198 8594 5232
rect 8688 5198 8704 5232
rect 8756 5198 8772 5232
rect 8866 5198 8882 5232
rect 8934 5198 8950 5232
rect 9044 5198 9060 5232
rect 9112 5198 9128 5232
rect 9222 5198 9238 5232
rect 9290 5198 9306 5232
rect 9400 5198 9416 5232
rect 9468 5198 9484 5232
rect 9578 5198 9594 5232
rect 9646 5198 9662 5232
rect 9756 5198 9772 5232
rect 9824 5198 9840 5232
rect 9934 5198 9950 5232
rect 10002 5198 10322 5232
rect 10374 5198 10390 5232
rect 10484 5198 10500 5232
rect 10552 5198 10568 5232
rect 10662 5198 10678 5232
rect 10730 5198 10746 5232
rect 10840 5198 10856 5232
rect 10908 5198 10924 5232
rect 11018 5198 11034 5232
rect 11086 5198 11102 5232
rect 11196 5198 11212 5232
rect 11264 5198 11280 5232
rect 11374 5198 11390 5232
rect 11442 5198 11458 5232
rect 11552 5198 11568 5232
rect 11620 5198 11636 5232
rect 11730 5198 11746 5232
rect 11798 5198 11814 5232
rect 11908 5198 11924 5232
rect 11976 5198 11992 5232
rect 12086 5198 12102 5232
rect 12154 5198 12170 5232
rect 12264 5198 12280 5232
rect 12332 5198 12505 5232
rect 7805 5139 7946 5198
rect 7805 4883 7912 5139
rect 7805 4824 7946 4883
rect 8090 5139 8124 5155
rect 8090 4867 8124 4883
rect 8268 5139 8302 5155
rect 8268 4867 8302 4883
rect 8446 5139 8480 5155
rect 8446 4867 8480 4883
rect 8624 5139 8658 5155
rect 8624 4867 8658 4883
rect 8802 5139 8836 5155
rect 8802 4867 8836 4883
rect 8980 5139 9014 5155
rect 8980 4867 9014 4883
rect 9158 5139 9192 5155
rect 9158 4867 9192 4883
rect 9336 5139 9370 5155
rect 9336 4867 9370 4883
rect 9514 5139 9548 5155
rect 9514 4867 9548 4883
rect 9692 5139 9726 5155
rect 9692 4867 9726 4883
rect 9870 5139 9904 5155
rect 9870 4867 9904 4883
rect 10048 5139 10276 5198
rect 10082 4883 10242 5139
rect 10048 4824 10276 4883
rect 10420 5139 10454 5155
rect 10420 4867 10454 4883
rect 10598 5139 10632 5155
rect 10598 4867 10632 4883
rect 10776 5139 10810 5155
rect 10776 4867 10810 4883
rect 10954 5139 10988 5155
rect 10954 4867 10988 4883
rect 11132 5139 11166 5155
rect 11132 4867 11166 4883
rect 11310 5139 11344 5155
rect 11310 4867 11344 4883
rect 11488 5139 11522 5155
rect 11488 4867 11522 4883
rect 11666 5139 11700 5155
rect 11666 4867 11700 4883
rect 11844 5139 11878 5155
rect 11844 4867 11878 4883
rect 12022 5139 12056 5155
rect 12022 4867 12056 4883
rect 12200 5139 12234 5155
rect 12200 4867 12234 4883
rect 12378 5139 12505 5198
rect 12412 4883 12505 5139
rect 12378 4824 12505 4883
rect 7805 4790 7992 4824
rect 8044 4790 8060 4824
rect 8154 4790 8170 4824
rect 8222 4790 8238 4824
rect 8332 4790 8348 4824
rect 8400 4790 8416 4824
rect 8510 4790 8526 4824
rect 8578 4790 8594 4824
rect 8688 4790 8704 4824
rect 8756 4790 8772 4824
rect 8866 4790 8882 4824
rect 8934 4790 8950 4824
rect 9044 4790 9060 4824
rect 9112 4790 9128 4824
rect 9222 4790 9238 4824
rect 9290 4790 9306 4824
rect 9400 4790 9416 4824
rect 9468 4790 9484 4824
rect 9578 4790 9594 4824
rect 9646 4790 9662 4824
rect 9756 4790 9772 4824
rect 9824 4790 9840 4824
rect 9934 4790 9950 4824
rect 10002 4790 10322 4824
rect 10374 4790 10390 4824
rect 10484 4790 10500 4824
rect 10552 4790 10568 4824
rect 10662 4790 10678 4824
rect 10730 4790 10746 4824
rect 10840 4790 10856 4824
rect 10908 4790 10924 4824
rect 11018 4790 11034 4824
rect 11086 4790 11102 4824
rect 11196 4790 11212 4824
rect 11264 4790 11280 4824
rect 11374 4790 11390 4824
rect 11442 4790 11458 4824
rect 11552 4790 11568 4824
rect 11620 4790 11636 4824
rect 11730 4790 11746 4824
rect 11798 4790 11814 4824
rect 11908 4790 11924 4824
rect 11976 4790 11992 4824
rect 12086 4790 12102 4824
rect 12154 4790 12170 4824
rect 12264 4790 12280 4824
rect 12332 4790 12505 4824
rect 7805 4662 7933 4790
rect 10053 4662 10258 4790
rect 12397 4662 12505 4790
rect 7805 4628 7992 4662
rect 8044 4628 8060 4662
rect 8154 4628 8170 4662
rect 8222 4628 8238 4662
rect 8332 4628 8348 4662
rect 8400 4628 8416 4662
rect 8510 4628 8526 4662
rect 8578 4628 8594 4662
rect 8688 4628 8704 4662
rect 8756 4628 8772 4662
rect 8866 4628 8882 4662
rect 8934 4628 8950 4662
rect 9044 4628 9060 4662
rect 9112 4628 9128 4662
rect 9222 4628 9238 4662
rect 9290 4628 9306 4662
rect 9400 4628 9416 4662
rect 9468 4628 9484 4662
rect 9578 4628 9594 4662
rect 9646 4628 9662 4662
rect 9756 4628 9772 4662
rect 9824 4628 9840 4662
rect 9934 4628 9950 4662
rect 10002 4628 10322 4662
rect 10374 4628 10390 4662
rect 10484 4628 10500 4662
rect 10552 4628 10568 4662
rect 10662 4628 10678 4662
rect 10730 4628 10746 4662
rect 10840 4628 10856 4662
rect 10908 4628 10924 4662
rect 11018 4628 11034 4662
rect 11086 4628 11102 4662
rect 11196 4628 11212 4662
rect 11264 4628 11280 4662
rect 11374 4628 11390 4662
rect 11442 4628 11458 4662
rect 11552 4628 11568 4662
rect 11620 4628 11636 4662
rect 11730 4628 11746 4662
rect 11798 4628 11814 4662
rect 11908 4628 11924 4662
rect 11976 4628 11992 4662
rect 12086 4628 12102 4662
rect 12154 4628 12170 4662
rect 12264 4628 12280 4662
rect 12332 4628 12505 4662
rect 7805 4569 7946 4628
rect 7805 4313 7912 4569
rect 7805 4254 7946 4313
rect 8090 4569 8124 4585
rect 8090 4297 8124 4313
rect 8268 4569 8302 4585
rect 8268 4297 8302 4313
rect 8446 4569 8480 4585
rect 8446 4297 8480 4313
rect 8624 4569 8658 4585
rect 8624 4297 8658 4313
rect 8802 4569 8836 4585
rect 8802 4297 8836 4313
rect 8980 4569 9014 4585
rect 8980 4297 9014 4313
rect 9158 4569 9192 4585
rect 9158 4297 9192 4313
rect 9336 4569 9370 4585
rect 9336 4297 9370 4313
rect 9514 4569 9548 4585
rect 9514 4297 9548 4313
rect 9692 4569 9726 4585
rect 9692 4297 9726 4313
rect 9870 4569 9904 4585
rect 9870 4297 9904 4313
rect 10048 4569 10276 4628
rect 10082 4313 10242 4569
rect 10048 4254 10276 4313
rect 10420 4569 10454 4585
rect 10420 4297 10454 4313
rect 10598 4569 10632 4585
rect 10598 4297 10632 4313
rect 10776 4569 10810 4585
rect 10776 4297 10810 4313
rect 10954 4569 10988 4585
rect 10954 4297 10988 4313
rect 11132 4569 11166 4585
rect 11132 4297 11166 4313
rect 11310 4569 11344 4585
rect 11310 4297 11344 4313
rect 11488 4569 11522 4585
rect 11488 4297 11522 4313
rect 11666 4569 11700 4585
rect 11666 4297 11700 4313
rect 11844 4569 11878 4585
rect 11844 4297 11878 4313
rect 12022 4569 12056 4585
rect 12022 4297 12056 4313
rect 12200 4569 12234 4585
rect 12200 4297 12234 4313
rect 12378 4569 12505 4628
rect 12412 4313 12505 4569
rect 12378 4254 12505 4313
rect 7805 4220 7992 4254
rect 8044 4220 8060 4254
rect 8154 4220 8170 4254
rect 8222 4220 8238 4254
rect 8332 4220 8348 4254
rect 8400 4220 8416 4254
rect 8510 4220 8526 4254
rect 8578 4220 8594 4254
rect 8688 4220 8704 4254
rect 8756 4220 8772 4254
rect 8866 4220 8882 4254
rect 8934 4220 8950 4254
rect 9044 4220 9060 4254
rect 9112 4220 9128 4254
rect 9222 4220 9238 4254
rect 9290 4220 9306 4254
rect 9400 4220 9416 4254
rect 9468 4220 9484 4254
rect 9578 4220 9594 4254
rect 9646 4220 9662 4254
rect 9756 4220 9772 4254
rect 9824 4220 9840 4254
rect 9934 4220 9950 4254
rect 10002 4220 10322 4254
rect 10374 4220 10390 4254
rect 10484 4220 10500 4254
rect 10552 4220 10568 4254
rect 10662 4220 10678 4254
rect 10730 4220 10746 4254
rect 10840 4220 10856 4254
rect 10908 4220 10924 4254
rect 11018 4220 11034 4254
rect 11086 4220 11102 4254
rect 11196 4220 11212 4254
rect 11264 4220 11280 4254
rect 11374 4220 11390 4254
rect 11442 4220 11458 4254
rect 11552 4220 11568 4254
rect 11620 4220 11636 4254
rect 11730 4220 11746 4254
rect 11798 4220 11814 4254
rect 11908 4220 11924 4254
rect 11976 4220 11992 4254
rect 12086 4220 12102 4254
rect 12154 4220 12170 4254
rect 12264 4220 12280 4254
rect 12332 4220 12505 4254
rect 7805 4124 7933 4220
rect 10053 4124 10258 4220
rect 12397 4124 12505 4220
rect 12999 4124 13033 4221
rect 7310 4090 7453 4124
rect 12924 4090 13033 4124
rect 13318 5260 13367 5261
rect 13318 5211 13584 5260
rect 13318 5128 13367 5211
rect 7805 4083 7933 4090
rect 6924 3934 6973 3960
rect 6924 3885 7001 3934
rect 13229 3885 13318 3934
rect 7047 3523 7184 3885
rect 428 3511 508 3523
rect 313 3489 508 3511
rect 560 3489 576 3523
rect 670 3489 686 3523
rect 738 3489 754 3523
rect 848 3489 864 3523
rect 916 3489 932 3523
rect 1026 3489 1042 3523
rect 1094 3489 1110 3523
rect 1204 3489 1220 3523
rect 1272 3489 1288 3523
rect 1382 3489 1398 3523
rect 1450 3489 1466 3523
rect 1560 3489 1576 3523
rect 1628 3489 1644 3523
rect 1738 3489 1754 3523
rect 1806 3489 1822 3523
rect 1916 3489 1932 3523
rect 1984 3489 2000 3523
rect 2094 3489 2110 3523
rect 2162 3489 2178 3523
rect 2272 3489 2288 3523
rect 2340 3489 2356 3523
rect 2450 3489 2466 3523
rect 2518 3489 2534 3523
rect 2628 3489 2644 3523
rect 2696 3489 2712 3523
rect 2806 3489 2822 3523
rect 2874 3489 2890 3523
rect 2984 3489 3000 3523
rect 3052 3489 3068 3523
rect 3162 3489 3178 3523
rect 3230 3489 3246 3523
rect 3340 3489 3356 3523
rect 3408 3489 3424 3523
rect 3518 3489 3534 3523
rect 3586 3489 3908 3523
rect 3960 3489 3976 3523
rect 4070 3489 4086 3523
rect 4138 3489 4154 3523
rect 4248 3489 4264 3523
rect 4316 3489 4332 3523
rect 4426 3489 4442 3523
rect 4494 3489 4510 3523
rect 4604 3489 4620 3523
rect 4672 3489 4688 3523
rect 4782 3489 4798 3523
rect 4850 3489 4866 3523
rect 4960 3489 4976 3523
rect 5028 3489 5044 3523
rect 5138 3489 5154 3523
rect 5206 3489 5222 3523
rect 5316 3489 5332 3523
rect 5384 3489 5400 3523
rect 5494 3489 5510 3523
rect 5562 3489 5578 3523
rect 5672 3489 5688 3523
rect 5740 3489 5756 3523
rect 5850 3489 5866 3523
rect 5918 3489 5934 3523
rect 6028 3489 6044 3523
rect 6096 3489 6112 3523
rect 6206 3489 6222 3523
rect 6274 3489 6290 3523
rect 6384 3489 6400 3523
rect 6452 3489 6468 3523
rect 6562 3489 6578 3523
rect 6630 3489 6646 3523
rect 6740 3489 6756 3523
rect 6808 3489 6824 3523
rect 6918 3489 6934 3523
rect 6986 3489 7184 3523
rect 313 3439 462 3489
rect 313 3183 428 3439
rect 313 3133 462 3183
rect 606 3439 640 3455
rect 606 3167 640 3183
rect 784 3439 818 3455
rect 784 3167 818 3183
rect 962 3439 996 3455
rect 962 3167 996 3183
rect 1140 3439 1174 3455
rect 1140 3167 1174 3183
rect 1318 3439 1352 3455
rect 1318 3167 1352 3183
rect 1496 3439 1530 3455
rect 1496 3167 1530 3183
rect 1674 3439 1708 3455
rect 1674 3167 1708 3183
rect 1852 3439 1886 3455
rect 1852 3167 1886 3183
rect 2030 3439 2064 3455
rect 2030 3167 2064 3183
rect 2208 3439 2242 3455
rect 2208 3167 2242 3183
rect 2386 3439 2420 3455
rect 2386 3167 2420 3183
rect 2564 3439 2598 3455
rect 2564 3167 2598 3183
rect 2742 3439 2776 3455
rect 2742 3167 2776 3183
rect 2920 3439 2954 3455
rect 2920 3167 2954 3183
rect 3098 3439 3132 3455
rect 3098 3167 3132 3183
rect 3276 3439 3310 3455
rect 3276 3167 3310 3183
rect 3454 3439 3488 3455
rect 3454 3167 3488 3183
rect 3632 3439 3862 3489
rect 3666 3183 3828 3439
rect 3632 3133 3862 3183
rect 4006 3439 4040 3455
rect 4006 3167 4040 3183
rect 4184 3439 4218 3455
rect 4184 3167 4218 3183
rect 4362 3439 4396 3455
rect 4362 3167 4396 3183
rect 4540 3439 4574 3455
rect 4540 3167 4574 3183
rect 4718 3439 4752 3455
rect 4718 3167 4752 3183
rect 4896 3439 4930 3455
rect 4896 3167 4930 3183
rect 5074 3439 5108 3455
rect 5074 3167 5108 3183
rect 5252 3439 5286 3455
rect 5252 3167 5286 3183
rect 5430 3439 5464 3455
rect 5430 3167 5464 3183
rect 5608 3439 5642 3455
rect 5608 3167 5642 3183
rect 5786 3439 5820 3455
rect 5786 3167 5820 3183
rect 5964 3439 5998 3455
rect 5964 3167 5998 3183
rect 6142 3439 6176 3455
rect 6142 3167 6176 3183
rect 6320 3439 6354 3455
rect 6320 3167 6354 3183
rect 6498 3439 6532 3455
rect 6498 3167 6532 3183
rect 6676 3439 6710 3455
rect 6676 3167 6710 3183
rect 6854 3439 6888 3455
rect 6854 3167 6888 3183
rect 7032 3439 7184 3489
rect 7066 3183 7184 3439
rect 7032 3133 7184 3183
rect 313 3099 508 3133
rect 560 3099 576 3133
rect 670 3099 686 3133
rect 738 3099 754 3133
rect 848 3099 864 3133
rect 916 3099 932 3133
rect 1026 3099 1042 3133
rect 1094 3099 1110 3133
rect 1204 3099 1220 3133
rect 1272 3099 1288 3133
rect 1382 3099 1398 3133
rect 1450 3099 1466 3133
rect 1560 3099 1576 3133
rect 1628 3099 1644 3133
rect 1738 3099 1754 3133
rect 1806 3099 1822 3133
rect 1916 3099 1932 3133
rect 1984 3099 2000 3133
rect 2094 3099 2110 3133
rect 2162 3099 2178 3133
rect 2272 3099 2288 3133
rect 2340 3099 2356 3133
rect 2450 3099 2466 3133
rect 2518 3099 2534 3133
rect 2628 3099 2644 3133
rect 2696 3099 2712 3133
rect 2806 3099 2822 3133
rect 2874 3099 2890 3133
rect 2984 3099 3000 3133
rect 3052 3099 3068 3133
rect 3162 3099 3178 3133
rect 3230 3099 3246 3133
rect 3340 3099 3356 3133
rect 3408 3099 3424 3133
rect 3518 3099 3534 3133
rect 3586 3099 3908 3133
rect 3960 3099 3976 3133
rect 4070 3099 4086 3133
rect 4138 3099 4154 3133
rect 4248 3099 4264 3133
rect 4316 3099 4332 3133
rect 4426 3099 4442 3133
rect 4494 3099 4510 3133
rect 4604 3099 4620 3133
rect 4672 3099 4688 3133
rect 4782 3099 4798 3133
rect 4850 3099 4866 3133
rect 4960 3099 4976 3133
rect 5028 3099 5044 3133
rect 5138 3099 5154 3133
rect 5206 3099 5222 3133
rect 5316 3099 5332 3133
rect 5384 3099 5400 3133
rect 5494 3099 5510 3133
rect 5562 3099 5578 3133
rect 5672 3099 5688 3133
rect 5740 3099 5756 3133
rect 5850 3099 5866 3133
rect 5918 3099 5934 3133
rect 6028 3099 6044 3133
rect 6096 3099 6112 3133
rect 6206 3099 6222 3133
rect 6274 3099 6290 3133
rect 6384 3099 6400 3133
rect 6452 3099 6468 3133
rect 6562 3099 6578 3133
rect 6630 3099 6646 3133
rect 6740 3099 6756 3133
rect 6808 3099 6824 3133
rect 6918 3099 6934 3133
rect 6986 3099 7184 3133
rect 313 3023 450 3099
rect 3649 3023 3843 3099
rect 7047 3023 7184 3099
rect 313 2989 508 3023
rect 560 2989 576 3023
rect 670 2989 686 3023
rect 738 2989 754 3023
rect 848 2989 864 3023
rect 916 2989 932 3023
rect 1026 2989 1042 3023
rect 1094 2989 1110 3023
rect 1204 2989 1220 3023
rect 1272 2989 1288 3023
rect 1382 2989 1398 3023
rect 1450 2989 1466 3023
rect 1560 2989 1576 3023
rect 1628 2989 1644 3023
rect 1738 2989 1754 3023
rect 1806 2989 1822 3023
rect 1916 2989 1932 3023
rect 1984 2989 2000 3023
rect 2094 2989 2110 3023
rect 2162 2989 2178 3023
rect 2272 2989 2288 3023
rect 2340 2989 2356 3023
rect 2450 2989 2466 3023
rect 2518 2989 2534 3023
rect 2628 2989 2644 3023
rect 2696 2989 2712 3023
rect 2806 2989 2822 3023
rect 2874 2989 2890 3023
rect 2984 2989 3000 3023
rect 3052 2989 3068 3023
rect 3162 2989 3178 3023
rect 3230 2989 3246 3023
rect 3340 2989 3356 3023
rect 3408 2989 3424 3023
rect 3518 2989 3534 3023
rect 3586 2989 3908 3023
rect 3960 2989 3976 3023
rect 4070 2989 4086 3023
rect 4138 2989 4154 3023
rect 4248 2989 4264 3023
rect 4316 2989 4332 3023
rect 4426 2989 4442 3023
rect 4494 2989 4510 3023
rect 4604 2989 4620 3023
rect 4672 2989 4688 3023
rect 4782 2989 4798 3023
rect 4850 2989 4866 3023
rect 4960 2989 4976 3023
rect 5028 2989 5044 3023
rect 5138 2989 5154 3023
rect 5206 2989 5222 3023
rect 5316 2989 5332 3023
rect 5384 2989 5400 3023
rect 5494 2989 5510 3023
rect 5562 2989 5578 3023
rect 5672 2989 5688 3023
rect 5740 2989 5756 3023
rect 5850 2989 5866 3023
rect 5918 2989 5934 3023
rect 6028 2989 6044 3023
rect 6096 2989 6112 3023
rect 6206 2989 6222 3023
rect 6274 2989 6290 3023
rect 6384 2989 6400 3023
rect 6452 2989 6468 3023
rect 6562 2989 6578 3023
rect 6630 2989 6646 3023
rect 6740 2989 6756 3023
rect 6808 2989 6824 3023
rect 6918 2989 6934 3023
rect 6986 2989 7184 3023
rect 313 2939 462 2989
rect 313 2683 428 2939
rect 313 2633 462 2683
rect 606 2939 640 2955
rect 606 2667 640 2683
rect 784 2939 818 2955
rect 784 2667 818 2683
rect 962 2939 996 2955
rect 962 2667 996 2683
rect 1140 2939 1174 2955
rect 1140 2667 1174 2683
rect 1318 2939 1352 2955
rect 1318 2667 1352 2683
rect 1496 2939 1530 2955
rect 1496 2667 1530 2683
rect 1674 2939 1708 2955
rect 1674 2667 1708 2683
rect 1852 2939 1886 2955
rect 1852 2667 1886 2683
rect 2030 2939 2064 2955
rect 2030 2667 2064 2683
rect 2208 2939 2242 2955
rect 2208 2667 2242 2683
rect 2386 2939 2420 2955
rect 2386 2667 2420 2683
rect 2564 2939 2598 2955
rect 2564 2667 2598 2683
rect 2742 2939 2776 2955
rect 2742 2667 2776 2683
rect 2920 2939 2954 2955
rect 2920 2667 2954 2683
rect 3098 2939 3132 2955
rect 3098 2667 3132 2683
rect 3276 2939 3310 2955
rect 3276 2667 3310 2683
rect 3454 2939 3488 2955
rect 3454 2667 3488 2683
rect 3632 2939 3862 2989
rect 3666 2683 3828 2939
rect 3632 2633 3862 2683
rect 4006 2939 4040 2955
rect 4006 2667 4040 2683
rect 4184 2939 4218 2955
rect 4184 2667 4218 2683
rect 4362 2939 4396 2955
rect 4362 2667 4396 2683
rect 4540 2939 4574 2955
rect 4540 2667 4574 2683
rect 4718 2939 4752 2955
rect 4718 2667 4752 2683
rect 4896 2939 4930 2955
rect 4896 2667 4930 2683
rect 5074 2939 5108 2955
rect 5074 2667 5108 2683
rect 5252 2939 5286 2955
rect 5252 2667 5286 2683
rect 5430 2939 5464 2955
rect 5430 2667 5464 2683
rect 5608 2939 5642 2955
rect 5608 2667 5642 2683
rect 5786 2939 5820 2955
rect 5786 2667 5820 2683
rect 5964 2939 5998 2955
rect 5964 2667 5998 2683
rect 6142 2939 6176 2955
rect 6142 2667 6176 2683
rect 6320 2939 6354 2955
rect 6320 2667 6354 2683
rect 6498 2939 6532 2955
rect 6498 2667 6532 2683
rect 6676 2939 6710 2955
rect 6676 2667 6710 2683
rect 6854 2939 6888 2955
rect 6854 2667 6888 2683
rect 7032 2939 7184 2989
rect 7066 2683 7184 2939
rect 7032 2633 7184 2683
rect 313 2599 508 2633
rect 560 2599 576 2633
rect 670 2599 686 2633
rect 738 2599 754 2633
rect 848 2599 864 2633
rect 916 2599 932 2633
rect 1026 2599 1042 2633
rect 1094 2599 1110 2633
rect 1204 2599 1220 2633
rect 1272 2599 1288 2633
rect 1382 2599 1398 2633
rect 1450 2599 1466 2633
rect 1560 2599 1576 2633
rect 1628 2599 1644 2633
rect 1738 2599 1754 2633
rect 1806 2599 1822 2633
rect 1916 2599 1932 2633
rect 1984 2599 2000 2633
rect 2094 2599 2110 2633
rect 2162 2599 2178 2633
rect 2272 2599 2288 2633
rect 2340 2599 2356 2633
rect 2450 2599 2466 2633
rect 2518 2599 2534 2633
rect 2628 2599 2644 2633
rect 2696 2599 2712 2633
rect 2806 2599 2822 2633
rect 2874 2599 2890 2633
rect 2984 2599 3000 2633
rect 3052 2599 3068 2633
rect 3162 2599 3178 2633
rect 3230 2599 3246 2633
rect 3340 2599 3356 2633
rect 3408 2599 3424 2633
rect 3518 2599 3534 2633
rect 3586 2599 3908 2633
rect 3960 2599 3976 2633
rect 4070 2599 4086 2633
rect 4138 2599 4154 2633
rect 4248 2599 4264 2633
rect 4316 2599 4332 2633
rect 4426 2599 4442 2633
rect 4494 2599 4510 2633
rect 4604 2599 4620 2633
rect 4672 2599 4688 2633
rect 4782 2599 4798 2633
rect 4850 2599 4866 2633
rect 4960 2599 4976 2633
rect 5028 2599 5044 2633
rect 5138 2599 5154 2633
rect 5206 2599 5222 2633
rect 5316 2599 5332 2633
rect 5384 2599 5400 2633
rect 5494 2599 5510 2633
rect 5562 2599 5578 2633
rect 5672 2599 5688 2633
rect 5740 2599 5756 2633
rect 5850 2599 5866 2633
rect 5918 2599 5934 2633
rect 6028 2599 6044 2633
rect 6096 2599 6112 2633
rect 6206 2599 6222 2633
rect 6274 2599 6290 2633
rect 6384 2599 6400 2633
rect 6452 2599 6468 2633
rect 6562 2599 6578 2633
rect 6630 2599 6646 2633
rect 6740 2599 6756 2633
rect 6808 2599 6824 2633
rect 6918 2599 6934 2633
rect 6986 2599 7184 2633
rect 313 2523 450 2599
rect 3649 2523 3843 2599
rect 7047 2523 7184 2599
rect 313 2489 508 2523
rect 560 2489 576 2523
rect 670 2489 686 2523
rect 738 2489 754 2523
rect 848 2489 864 2523
rect 916 2489 932 2523
rect 1026 2489 1042 2523
rect 1094 2489 1110 2523
rect 1204 2489 1220 2523
rect 1272 2489 1288 2523
rect 1382 2489 1398 2523
rect 1450 2489 1466 2523
rect 1560 2489 1576 2523
rect 1628 2489 1644 2523
rect 1738 2489 1754 2523
rect 1806 2489 1822 2523
rect 1916 2489 1932 2523
rect 1984 2489 2000 2523
rect 2094 2489 2110 2523
rect 2162 2489 2178 2523
rect 2272 2489 2288 2523
rect 2340 2489 2356 2523
rect 2450 2489 2466 2523
rect 2518 2489 2534 2523
rect 2628 2489 2644 2523
rect 2696 2489 2712 2523
rect 2806 2489 2822 2523
rect 2874 2489 2890 2523
rect 2984 2489 3000 2523
rect 3052 2489 3068 2523
rect 3162 2489 3178 2523
rect 3230 2489 3246 2523
rect 3340 2489 3356 2523
rect 3408 2489 3424 2523
rect 3518 2489 3534 2523
rect 3586 2489 3908 2523
rect 3960 2489 3976 2523
rect 4070 2489 4086 2523
rect 4138 2489 4154 2523
rect 4248 2489 4264 2523
rect 4316 2489 4332 2523
rect 4426 2489 4442 2523
rect 4494 2489 4510 2523
rect 4604 2489 4620 2523
rect 4672 2489 4688 2523
rect 4782 2489 4798 2523
rect 4850 2489 4866 2523
rect 4960 2489 4976 2523
rect 5028 2489 5044 2523
rect 5138 2489 5154 2523
rect 5206 2489 5222 2523
rect 5316 2489 5332 2523
rect 5384 2489 5400 2523
rect 5494 2489 5510 2523
rect 5562 2489 5578 2523
rect 5672 2489 5688 2523
rect 5740 2489 5756 2523
rect 5850 2489 5866 2523
rect 5918 2489 5934 2523
rect 6028 2489 6044 2523
rect 6096 2489 6112 2523
rect 6206 2489 6222 2523
rect 6274 2489 6290 2523
rect 6384 2489 6400 2523
rect 6452 2489 6468 2523
rect 6562 2489 6578 2523
rect 6630 2489 6646 2523
rect 6740 2489 6756 2523
rect 6808 2489 6824 2523
rect 6918 2489 6934 2523
rect 6986 2489 7184 2523
rect 313 2439 462 2489
rect 313 2183 428 2439
rect 313 2133 462 2183
rect 606 2439 640 2455
rect 606 2167 640 2183
rect 784 2439 818 2455
rect 784 2167 818 2183
rect 962 2439 996 2455
rect 962 2167 996 2183
rect 1140 2439 1174 2455
rect 1140 2167 1174 2183
rect 1318 2439 1352 2455
rect 1318 2167 1352 2183
rect 1496 2439 1530 2455
rect 1496 2167 1530 2183
rect 1674 2439 1708 2455
rect 1674 2167 1708 2183
rect 1852 2439 1886 2455
rect 1852 2167 1886 2183
rect 2030 2439 2064 2455
rect 2030 2167 2064 2183
rect 2208 2439 2242 2455
rect 2208 2167 2242 2183
rect 2386 2439 2420 2455
rect 2386 2167 2420 2183
rect 2564 2439 2598 2455
rect 2564 2167 2598 2183
rect 2742 2439 2776 2455
rect 2742 2167 2776 2183
rect 2920 2439 2954 2455
rect 2920 2167 2954 2183
rect 3098 2439 3132 2455
rect 3098 2167 3132 2183
rect 3276 2439 3310 2455
rect 3276 2167 3310 2183
rect 3454 2439 3488 2455
rect 3454 2167 3488 2183
rect 3632 2439 3862 2489
rect 3666 2183 3828 2439
rect 3632 2133 3862 2183
rect 4006 2439 4040 2455
rect 4006 2167 4040 2183
rect 4184 2439 4218 2455
rect 4184 2167 4218 2183
rect 4362 2439 4396 2455
rect 4362 2167 4396 2183
rect 4540 2439 4574 2455
rect 4540 2167 4574 2183
rect 4718 2439 4752 2455
rect 4718 2167 4752 2183
rect 4896 2439 4930 2455
rect 4896 2167 4930 2183
rect 5074 2439 5108 2455
rect 5074 2167 5108 2183
rect 5252 2439 5286 2455
rect 5252 2167 5286 2183
rect 5430 2439 5464 2455
rect 5430 2167 5464 2183
rect 5608 2439 5642 2455
rect 5608 2167 5642 2183
rect 5786 2439 5820 2455
rect 5786 2167 5820 2183
rect 5964 2439 5998 2455
rect 5964 2167 5998 2183
rect 6142 2439 6176 2455
rect 6142 2167 6176 2183
rect 6320 2439 6354 2455
rect 6320 2167 6354 2183
rect 6498 2439 6532 2455
rect 6498 2167 6532 2183
rect 6676 2439 6710 2455
rect 6676 2167 6710 2183
rect 6854 2439 6888 2455
rect 6854 2167 6888 2183
rect 7032 2439 7184 2489
rect 7066 2183 7184 2439
rect 7032 2133 7184 2183
rect 313 2099 508 2133
rect 560 2099 576 2133
rect 670 2099 686 2133
rect 738 2099 754 2133
rect 848 2099 864 2133
rect 916 2099 932 2133
rect 1026 2099 1042 2133
rect 1094 2099 1110 2133
rect 1204 2099 1220 2133
rect 1272 2099 1288 2133
rect 1382 2099 1398 2133
rect 1450 2099 1466 2133
rect 1560 2099 1576 2133
rect 1628 2099 1644 2133
rect 1738 2099 1754 2133
rect 1806 2099 1822 2133
rect 1916 2099 1932 2133
rect 1984 2099 2000 2133
rect 2094 2099 2110 2133
rect 2162 2099 2178 2133
rect 2272 2099 2288 2133
rect 2340 2099 2356 2133
rect 2450 2099 2466 2133
rect 2518 2099 2534 2133
rect 2628 2099 2644 2133
rect 2696 2099 2712 2133
rect 2806 2099 2822 2133
rect 2874 2099 2890 2133
rect 2984 2099 3000 2133
rect 3052 2099 3068 2133
rect 3162 2099 3178 2133
rect 3230 2099 3246 2133
rect 3340 2099 3356 2133
rect 3408 2099 3424 2133
rect 3518 2099 3534 2133
rect 3586 2099 3908 2133
rect 3960 2099 3976 2133
rect 4070 2099 4086 2133
rect 4138 2099 4154 2133
rect 4248 2099 4264 2133
rect 4316 2099 4332 2133
rect 4426 2099 4442 2133
rect 4494 2099 4510 2133
rect 4604 2099 4620 2133
rect 4672 2099 4688 2133
rect 4782 2099 4798 2133
rect 4850 2099 4866 2133
rect 4960 2099 4976 2133
rect 5028 2099 5044 2133
rect 5138 2099 5154 2133
rect 5206 2099 5222 2133
rect 5316 2099 5332 2133
rect 5384 2099 5400 2133
rect 5494 2099 5510 2133
rect 5562 2099 5578 2133
rect 5672 2099 5688 2133
rect 5740 2099 5756 2133
rect 5850 2099 5866 2133
rect 5918 2099 5934 2133
rect 6028 2099 6044 2133
rect 6096 2099 6112 2133
rect 6206 2099 6222 2133
rect 6274 2099 6290 2133
rect 6384 2099 6400 2133
rect 6452 2099 6468 2133
rect 6562 2099 6578 2133
rect 6630 2099 6646 2133
rect 6740 2099 6756 2133
rect 6808 2099 6824 2133
rect 6918 2099 6934 2133
rect 6986 2099 7184 2133
rect 313 2023 450 2099
rect 3649 2023 3843 2099
rect 7047 2023 7184 2099
rect 313 1989 508 2023
rect 560 1989 576 2023
rect 670 1989 686 2023
rect 738 1989 754 2023
rect 848 1989 864 2023
rect 916 1989 932 2023
rect 1026 1989 1042 2023
rect 1094 1989 1110 2023
rect 1204 1989 1220 2023
rect 1272 1989 1288 2023
rect 1382 1989 1398 2023
rect 1450 1989 1466 2023
rect 1560 1989 1576 2023
rect 1628 1989 1644 2023
rect 1738 1989 1754 2023
rect 1806 1989 1822 2023
rect 1916 1989 1932 2023
rect 1984 1989 2000 2023
rect 2094 1989 2110 2023
rect 2162 1989 2178 2023
rect 2272 1989 2288 2023
rect 2340 1989 2356 2023
rect 2450 1989 2466 2023
rect 2518 1989 2534 2023
rect 2628 1989 2644 2023
rect 2696 1989 2712 2023
rect 2806 1989 2822 2023
rect 2874 1989 2890 2023
rect 2984 1989 3000 2023
rect 3052 1989 3068 2023
rect 3162 1989 3178 2023
rect 3230 1989 3246 2023
rect 3340 1989 3356 2023
rect 3408 1989 3424 2023
rect 3518 1989 3534 2023
rect 3586 1989 3908 2023
rect 3960 1989 3976 2023
rect 4070 1989 4086 2023
rect 4138 1989 4154 2023
rect 4248 1989 4264 2023
rect 4316 1989 4332 2023
rect 4426 1989 4442 2023
rect 4494 1989 4510 2023
rect 4604 1989 4620 2023
rect 4672 1989 4688 2023
rect 4782 1989 4798 2023
rect 4850 1989 4866 2023
rect 4960 1989 4976 2023
rect 5028 1989 5044 2023
rect 5138 1989 5154 2023
rect 5206 1989 5222 2023
rect 5316 1989 5332 2023
rect 5384 1989 5400 2023
rect 5494 1989 5510 2023
rect 5562 1989 5578 2023
rect 5672 1989 5688 2023
rect 5740 1989 5756 2023
rect 5850 1989 5866 2023
rect 5918 1989 5934 2023
rect 6028 1989 6044 2023
rect 6096 1989 6112 2023
rect 6206 1989 6222 2023
rect 6274 1989 6290 2023
rect 6384 1989 6400 2023
rect 6452 1989 6468 2023
rect 6562 1989 6578 2023
rect 6630 1989 6646 2023
rect 6740 1989 6756 2023
rect 6808 1989 6824 2023
rect 6918 1989 6934 2023
rect 6986 1989 7184 2023
rect 313 1939 462 1989
rect 313 1683 428 1939
rect 313 1633 462 1683
rect 606 1939 640 1955
rect 606 1667 640 1683
rect 784 1939 818 1955
rect 784 1667 818 1683
rect 962 1939 996 1955
rect 962 1667 996 1683
rect 1140 1939 1174 1955
rect 1140 1667 1174 1683
rect 1318 1939 1352 1955
rect 1318 1667 1352 1683
rect 1496 1939 1530 1955
rect 1496 1667 1530 1683
rect 1674 1939 1708 1955
rect 1674 1667 1708 1683
rect 1852 1939 1886 1955
rect 1852 1667 1886 1683
rect 2030 1939 2064 1955
rect 2030 1667 2064 1683
rect 2208 1939 2242 1955
rect 2208 1667 2242 1683
rect 2386 1939 2420 1955
rect 2386 1667 2420 1683
rect 2564 1939 2598 1955
rect 2564 1667 2598 1683
rect 2742 1939 2776 1955
rect 2742 1667 2776 1683
rect 2920 1939 2954 1955
rect 2920 1667 2954 1683
rect 3098 1939 3132 1955
rect 3098 1667 3132 1683
rect 3276 1939 3310 1955
rect 3276 1667 3310 1683
rect 3454 1939 3488 1955
rect 3454 1667 3488 1683
rect 3632 1939 3862 1989
rect 3666 1683 3828 1939
rect 3632 1633 3862 1683
rect 4006 1939 4040 1955
rect 4006 1667 4040 1683
rect 4184 1939 4218 1955
rect 4184 1667 4218 1683
rect 4362 1939 4396 1955
rect 4362 1667 4396 1683
rect 4540 1939 4574 1955
rect 4540 1667 4574 1683
rect 4718 1939 4752 1955
rect 4718 1667 4752 1683
rect 4896 1939 4930 1955
rect 4896 1667 4930 1683
rect 5074 1939 5108 1955
rect 5074 1667 5108 1683
rect 5252 1939 5286 1955
rect 5252 1667 5286 1683
rect 5430 1939 5464 1955
rect 5430 1667 5464 1683
rect 5608 1939 5642 1955
rect 5608 1667 5642 1683
rect 5786 1939 5820 1955
rect 5786 1667 5820 1683
rect 5964 1939 5998 1955
rect 5964 1667 5998 1683
rect 6142 1939 6176 1955
rect 6142 1667 6176 1683
rect 6320 1939 6354 1955
rect 6320 1667 6354 1683
rect 6498 1939 6532 1955
rect 6498 1667 6532 1683
rect 6676 1939 6710 1955
rect 6676 1667 6710 1683
rect 6854 1939 6888 1955
rect 6854 1667 6888 1683
rect 7032 1939 7184 1989
rect 7066 1683 7184 1939
rect 7032 1633 7184 1683
rect 313 1599 508 1633
rect 560 1599 576 1633
rect 670 1599 686 1633
rect 738 1599 754 1633
rect 848 1599 864 1633
rect 916 1599 932 1633
rect 1026 1599 1042 1633
rect 1094 1599 1110 1633
rect 1204 1599 1220 1633
rect 1272 1599 1288 1633
rect 1382 1599 1398 1633
rect 1450 1599 1466 1633
rect 1560 1599 1576 1633
rect 1628 1599 1644 1633
rect 1738 1599 1754 1633
rect 1806 1599 1822 1633
rect 1916 1599 1932 1633
rect 1984 1599 2000 1633
rect 2094 1599 2110 1633
rect 2162 1599 2178 1633
rect 2272 1599 2288 1633
rect 2340 1599 2356 1633
rect 2450 1599 2466 1633
rect 2518 1599 2534 1633
rect 2628 1599 2644 1633
rect 2696 1599 2712 1633
rect 2806 1599 2822 1633
rect 2874 1599 2890 1633
rect 2984 1599 3000 1633
rect 3052 1599 3068 1633
rect 3162 1599 3178 1633
rect 3230 1599 3246 1633
rect 3340 1599 3356 1633
rect 3408 1599 3424 1633
rect 3518 1599 3534 1633
rect 3586 1599 3908 1633
rect 3960 1599 3976 1633
rect 4070 1599 4086 1633
rect 4138 1599 4154 1633
rect 4248 1599 4264 1633
rect 4316 1599 4332 1633
rect 4426 1599 4442 1633
rect 4494 1599 4510 1633
rect 4604 1599 4620 1633
rect 4672 1599 4688 1633
rect 4782 1599 4798 1633
rect 4850 1599 4866 1633
rect 4960 1599 4976 1633
rect 5028 1599 5044 1633
rect 5138 1599 5154 1633
rect 5206 1599 5222 1633
rect 5316 1599 5332 1633
rect 5384 1599 5400 1633
rect 5494 1599 5510 1633
rect 5562 1599 5578 1633
rect 5672 1599 5688 1633
rect 5740 1599 5756 1633
rect 5850 1599 5866 1633
rect 5918 1599 5934 1633
rect 6028 1599 6044 1633
rect 6096 1599 6112 1633
rect 6206 1599 6222 1633
rect 6274 1599 6290 1633
rect 6384 1599 6400 1633
rect 6452 1599 6468 1633
rect 6562 1599 6578 1633
rect 6630 1599 6646 1633
rect 6740 1599 6756 1633
rect 6808 1599 6824 1633
rect 6918 1599 6934 1633
rect 6986 1599 7184 1633
rect 313 1523 450 1599
rect 3649 1523 3843 1599
rect 7047 1523 7184 1599
rect 313 1489 508 1523
rect 560 1489 576 1523
rect 670 1489 686 1523
rect 738 1489 754 1523
rect 848 1489 864 1523
rect 916 1489 932 1523
rect 1026 1489 1042 1523
rect 1094 1489 1110 1523
rect 1204 1489 1220 1523
rect 1272 1489 1288 1523
rect 1382 1489 1398 1523
rect 1450 1489 1466 1523
rect 1560 1489 1576 1523
rect 1628 1489 1644 1523
rect 1738 1489 1754 1523
rect 1806 1489 1822 1523
rect 1916 1489 1932 1523
rect 1984 1489 2000 1523
rect 2094 1489 2110 1523
rect 2162 1489 2178 1523
rect 2272 1489 2288 1523
rect 2340 1489 2356 1523
rect 2450 1489 2466 1523
rect 2518 1489 2534 1523
rect 2628 1489 2644 1523
rect 2696 1489 2712 1523
rect 2806 1489 2822 1523
rect 2874 1489 2890 1523
rect 2984 1489 3000 1523
rect 3052 1489 3068 1523
rect 3162 1489 3178 1523
rect 3230 1489 3246 1523
rect 3340 1489 3356 1523
rect 3408 1489 3424 1523
rect 3518 1489 3534 1523
rect 3586 1489 3908 1523
rect 3960 1489 3976 1523
rect 4070 1489 4086 1523
rect 4138 1489 4154 1523
rect 4248 1489 4264 1523
rect 4316 1489 4332 1523
rect 4426 1489 4442 1523
rect 4494 1489 4510 1523
rect 4604 1489 4620 1523
rect 4672 1489 4688 1523
rect 4782 1489 4798 1523
rect 4850 1489 4866 1523
rect 4960 1489 4976 1523
rect 5028 1489 5044 1523
rect 5138 1489 5154 1523
rect 5206 1489 5222 1523
rect 5316 1489 5332 1523
rect 5384 1489 5400 1523
rect 5494 1489 5510 1523
rect 5562 1489 5578 1523
rect 5672 1489 5688 1523
rect 5740 1489 5756 1523
rect 5850 1489 5866 1523
rect 5918 1489 5934 1523
rect 6028 1489 6044 1523
rect 6096 1489 6112 1523
rect 6206 1489 6222 1523
rect 6274 1489 6290 1523
rect 6384 1489 6400 1523
rect 6452 1489 6468 1523
rect 6562 1489 6578 1523
rect 6630 1489 6646 1523
rect 6740 1489 6756 1523
rect 6808 1489 6824 1523
rect 6918 1489 6934 1523
rect 6986 1489 7184 1523
rect 313 1439 462 1489
rect 313 1183 428 1439
rect 313 1133 462 1183
rect 606 1439 640 1455
rect 606 1167 640 1183
rect 784 1439 818 1455
rect 784 1167 818 1183
rect 962 1439 996 1455
rect 962 1167 996 1183
rect 1140 1439 1174 1455
rect 1140 1167 1174 1183
rect 1318 1439 1352 1455
rect 1318 1167 1352 1183
rect 1496 1439 1530 1455
rect 1496 1167 1530 1183
rect 1674 1439 1708 1455
rect 1674 1167 1708 1183
rect 1852 1439 1886 1455
rect 1852 1167 1886 1183
rect 2030 1439 2064 1455
rect 2030 1167 2064 1183
rect 2208 1439 2242 1455
rect 2208 1167 2242 1183
rect 2386 1439 2420 1455
rect 2386 1167 2420 1183
rect 2564 1439 2598 1455
rect 2564 1167 2598 1183
rect 2742 1439 2776 1455
rect 2742 1167 2776 1183
rect 2920 1439 2954 1455
rect 2920 1167 2954 1183
rect 3098 1439 3132 1455
rect 3098 1167 3132 1183
rect 3276 1439 3310 1455
rect 3276 1167 3310 1183
rect 3454 1439 3488 1455
rect 3454 1167 3488 1183
rect 3632 1439 3862 1489
rect 3666 1183 3828 1439
rect 3632 1133 3862 1183
rect 4006 1439 4040 1455
rect 4006 1167 4040 1183
rect 4184 1439 4218 1455
rect 4184 1167 4218 1183
rect 4362 1439 4396 1455
rect 4362 1167 4396 1183
rect 4540 1439 4574 1455
rect 4540 1167 4574 1183
rect 4718 1439 4752 1455
rect 4718 1167 4752 1183
rect 4896 1439 4930 1455
rect 4896 1167 4930 1183
rect 5074 1439 5108 1455
rect 5074 1167 5108 1183
rect 5252 1439 5286 1455
rect 5252 1167 5286 1183
rect 5430 1439 5464 1455
rect 5430 1167 5464 1183
rect 5608 1439 5642 1455
rect 5608 1167 5642 1183
rect 5786 1439 5820 1455
rect 5786 1167 5820 1183
rect 5964 1439 5998 1455
rect 5964 1167 5998 1183
rect 6142 1439 6176 1455
rect 6142 1167 6176 1183
rect 6320 1439 6354 1455
rect 6320 1167 6354 1183
rect 6498 1439 6532 1455
rect 6498 1167 6532 1183
rect 6676 1439 6710 1455
rect 6676 1167 6710 1183
rect 6854 1439 6888 1455
rect 6854 1167 6888 1183
rect 7032 1439 7184 1489
rect 7066 1183 7184 1439
rect 7032 1133 7184 1183
rect 313 1099 508 1133
rect 560 1099 576 1133
rect 670 1099 686 1133
rect 738 1099 754 1133
rect 848 1099 864 1133
rect 916 1099 932 1133
rect 1026 1099 1042 1133
rect 1094 1099 1110 1133
rect 1204 1099 1220 1133
rect 1272 1099 1288 1133
rect 1382 1099 1398 1133
rect 1450 1099 1466 1133
rect 1560 1099 1576 1133
rect 1628 1099 1644 1133
rect 1738 1099 1754 1133
rect 1806 1099 1822 1133
rect 1916 1099 1932 1133
rect 1984 1099 2000 1133
rect 2094 1099 2110 1133
rect 2162 1099 2178 1133
rect 2272 1099 2288 1133
rect 2340 1099 2356 1133
rect 2450 1099 2466 1133
rect 2518 1099 2534 1133
rect 2628 1099 2644 1133
rect 2696 1099 2712 1133
rect 2806 1099 2822 1133
rect 2874 1099 2890 1133
rect 2984 1099 3000 1133
rect 3052 1099 3068 1133
rect 3162 1099 3178 1133
rect 3230 1099 3246 1133
rect 3340 1099 3356 1133
rect 3408 1099 3424 1133
rect 3518 1099 3534 1133
rect 3586 1099 3908 1133
rect 3960 1099 3976 1133
rect 4070 1099 4086 1133
rect 4138 1099 4154 1133
rect 4248 1099 4264 1133
rect 4316 1099 4332 1133
rect 4426 1099 4442 1133
rect 4494 1099 4510 1133
rect 4604 1099 4620 1133
rect 4672 1099 4688 1133
rect 4782 1099 4798 1133
rect 4850 1099 4866 1133
rect 4960 1099 4976 1133
rect 5028 1099 5044 1133
rect 5138 1099 5154 1133
rect 5206 1099 5222 1133
rect 5316 1099 5332 1133
rect 5384 1099 5400 1133
rect 5494 1099 5510 1133
rect 5562 1099 5578 1133
rect 5672 1099 5688 1133
rect 5740 1099 5756 1133
rect 5850 1099 5866 1133
rect 5918 1099 5934 1133
rect 6028 1099 6044 1133
rect 6096 1099 6112 1133
rect 6206 1099 6222 1133
rect 6274 1099 6290 1133
rect 6384 1099 6400 1133
rect 6452 1099 6468 1133
rect 6562 1099 6578 1133
rect 6630 1099 6646 1133
rect 6740 1099 6756 1133
rect 6808 1099 6824 1133
rect 6918 1099 6934 1133
rect 6986 1099 7184 1133
rect 313 1023 450 1099
rect 3649 1023 3843 1099
rect 7047 1023 7184 1099
rect 313 989 508 1023
rect 560 989 576 1023
rect 670 989 686 1023
rect 738 989 754 1023
rect 848 989 864 1023
rect 916 989 932 1023
rect 1026 989 1042 1023
rect 1094 989 1110 1023
rect 1204 989 1220 1023
rect 1272 989 1288 1023
rect 1382 989 1398 1023
rect 1450 989 1466 1023
rect 1560 989 1576 1023
rect 1628 989 1644 1023
rect 1738 989 1754 1023
rect 1806 989 1822 1023
rect 1916 989 1932 1023
rect 1984 989 2000 1023
rect 2094 989 2110 1023
rect 2162 989 2178 1023
rect 2272 989 2288 1023
rect 2340 989 2356 1023
rect 2450 989 2466 1023
rect 2518 989 2534 1023
rect 2628 989 2644 1023
rect 2696 989 2712 1023
rect 2806 989 2822 1023
rect 2874 989 2890 1023
rect 2984 989 3000 1023
rect 3052 989 3068 1023
rect 3162 989 3178 1023
rect 3230 989 3246 1023
rect 3340 989 3356 1023
rect 3408 989 3424 1023
rect 3518 989 3534 1023
rect 3586 989 3908 1023
rect 3960 989 3976 1023
rect 4070 989 4086 1023
rect 4138 989 4154 1023
rect 4248 989 4264 1023
rect 4316 989 4332 1023
rect 4426 989 4442 1023
rect 4494 989 4510 1023
rect 4604 989 4620 1023
rect 4672 989 4688 1023
rect 4782 989 4798 1023
rect 4850 989 4866 1023
rect 4960 989 4976 1023
rect 5028 989 5044 1023
rect 5138 989 5154 1023
rect 5206 989 5222 1023
rect 5316 989 5332 1023
rect 5384 989 5400 1023
rect 5494 989 5510 1023
rect 5562 989 5578 1023
rect 5672 989 5688 1023
rect 5740 989 5756 1023
rect 5850 989 5866 1023
rect 5918 989 5934 1023
rect 6028 989 6044 1023
rect 6096 989 6112 1023
rect 6206 989 6222 1023
rect 6274 989 6290 1023
rect 6384 989 6400 1023
rect 6452 989 6468 1023
rect 6562 989 6578 1023
rect 6630 989 6646 1023
rect 6740 989 6756 1023
rect 6808 989 6824 1023
rect 6918 989 6934 1023
rect 6986 989 7184 1023
rect 313 939 462 989
rect 313 683 428 939
rect 313 633 462 683
rect 606 939 640 955
rect 606 667 640 683
rect 784 939 818 955
rect 784 667 818 683
rect 962 939 996 955
rect 962 667 996 683
rect 1140 939 1174 955
rect 1140 667 1174 683
rect 1318 939 1352 955
rect 1318 667 1352 683
rect 1496 939 1530 955
rect 1496 667 1530 683
rect 1674 939 1708 955
rect 1674 667 1708 683
rect 1852 939 1886 955
rect 1852 667 1886 683
rect 2030 939 2064 955
rect 2030 667 2064 683
rect 2208 939 2242 955
rect 2208 667 2242 683
rect 2386 939 2420 955
rect 2386 667 2420 683
rect 2564 939 2598 955
rect 2564 667 2598 683
rect 2742 939 2776 955
rect 2742 667 2776 683
rect 2920 939 2954 955
rect 2920 667 2954 683
rect 3098 939 3132 955
rect 3098 667 3132 683
rect 3276 939 3310 955
rect 3276 667 3310 683
rect 3454 939 3488 955
rect 3454 667 3488 683
rect 3632 939 3862 989
rect 3666 683 3828 939
rect 3632 633 3862 683
rect 4006 939 4040 955
rect 4006 667 4040 683
rect 4184 939 4218 955
rect 4184 667 4218 683
rect 4362 939 4396 955
rect 4362 667 4396 683
rect 4540 939 4574 955
rect 4540 667 4574 683
rect 4718 939 4752 955
rect 4718 667 4752 683
rect 4896 939 4930 955
rect 4896 667 4930 683
rect 5074 939 5108 955
rect 5074 667 5108 683
rect 5252 939 5286 955
rect 5252 667 5286 683
rect 5430 939 5464 955
rect 5430 667 5464 683
rect 5608 939 5642 955
rect 5608 667 5642 683
rect 5786 939 5820 955
rect 5786 667 5820 683
rect 5964 939 5998 955
rect 5964 667 5998 683
rect 6142 939 6176 955
rect 6142 667 6176 683
rect 6320 939 6354 955
rect 6320 667 6354 683
rect 6498 939 6532 955
rect 6498 667 6532 683
rect 6676 939 6710 955
rect 6676 667 6710 683
rect 6854 939 6888 955
rect 6854 667 6888 683
rect 7032 939 7184 989
rect 7066 683 7184 939
rect 7032 633 7184 683
rect 313 599 508 633
rect 560 599 576 633
rect 670 599 686 633
rect 738 599 754 633
rect 848 599 864 633
rect 916 599 932 633
rect 1026 599 1042 633
rect 1094 599 1110 633
rect 1204 599 1220 633
rect 1272 599 1288 633
rect 1382 599 1398 633
rect 1450 599 1466 633
rect 1560 599 1576 633
rect 1628 599 1644 633
rect 1738 599 1754 633
rect 1806 599 1822 633
rect 1916 599 1932 633
rect 1984 599 2000 633
rect 2094 599 2110 633
rect 2162 599 2178 633
rect 2272 599 2288 633
rect 2340 599 2356 633
rect 2450 599 2466 633
rect 2518 599 2534 633
rect 2628 599 2644 633
rect 2696 599 2712 633
rect 2806 599 2822 633
rect 2874 599 2890 633
rect 2984 599 3000 633
rect 3052 599 3068 633
rect 3162 599 3178 633
rect 3230 599 3246 633
rect 3340 599 3356 633
rect 3408 599 3424 633
rect 3518 599 3534 633
rect 3586 599 3908 633
rect 3960 599 3976 633
rect 4070 599 4086 633
rect 4138 599 4154 633
rect 4248 599 4264 633
rect 4316 599 4332 633
rect 4426 599 4442 633
rect 4494 599 4510 633
rect 4604 599 4620 633
rect 4672 599 4688 633
rect 4782 599 4798 633
rect 4850 599 4866 633
rect 4960 599 4976 633
rect 5028 599 5044 633
rect 5138 599 5154 633
rect 5206 599 5222 633
rect 5316 599 5332 633
rect 5384 599 5400 633
rect 5494 599 5510 633
rect 5562 599 5578 633
rect 5672 599 5688 633
rect 5740 599 5756 633
rect 5850 599 5866 633
rect 5918 599 5934 633
rect 6028 599 6044 633
rect 6096 599 6112 633
rect 6206 599 6222 633
rect 6274 599 6290 633
rect 6384 599 6400 633
rect 6452 599 6468 633
rect 6562 599 6578 633
rect 6630 599 6646 633
rect 6740 599 6756 633
rect 6808 599 6824 633
rect 6918 599 6934 633
rect 6986 599 7184 633
rect 313 149 450 599
rect 3649 149 3843 599
rect 7047 149 7184 599
rect 7442 3723 7579 3885
rect 10067 3723 10261 3885
rect 12757 3723 12894 3885
rect 7442 3689 7637 3723
rect 7689 3689 7705 3723
rect 7799 3689 7815 3723
rect 7867 3689 7883 3723
rect 7977 3689 7993 3723
rect 8045 3689 8061 3723
rect 8155 3689 8171 3723
rect 8223 3689 8239 3723
rect 8333 3689 8349 3723
rect 8401 3689 8417 3723
rect 8511 3689 8527 3723
rect 8579 3689 8595 3723
rect 8689 3689 8705 3723
rect 8757 3689 8773 3723
rect 8867 3689 8883 3723
rect 8935 3689 8951 3723
rect 9045 3689 9061 3723
rect 9113 3689 9129 3723
rect 9223 3689 9239 3723
rect 9291 3689 9307 3723
rect 9401 3689 9417 3723
rect 9469 3689 9485 3723
rect 9579 3689 9595 3723
rect 9647 3689 9663 3723
rect 9757 3689 9773 3723
rect 9825 3689 9841 3723
rect 9935 3689 9951 3723
rect 10003 3689 10324 3723
rect 10376 3689 10392 3723
rect 10486 3689 10502 3723
rect 10554 3689 10570 3723
rect 10664 3689 10680 3723
rect 10732 3689 10748 3723
rect 10842 3689 10858 3723
rect 10910 3689 10926 3723
rect 11020 3689 11036 3723
rect 11088 3689 11104 3723
rect 11198 3689 11214 3723
rect 11266 3689 11282 3723
rect 11376 3689 11392 3723
rect 11444 3689 11460 3723
rect 11554 3689 11570 3723
rect 11622 3689 11638 3723
rect 11732 3689 11748 3723
rect 11800 3689 11816 3723
rect 11910 3689 11926 3723
rect 11978 3689 11994 3723
rect 12088 3689 12104 3723
rect 12156 3689 12172 3723
rect 12266 3689 12282 3723
rect 12334 3689 12350 3723
rect 12444 3689 12460 3723
rect 12512 3689 12528 3723
rect 12622 3689 12638 3723
rect 12690 3689 12894 3723
rect 7442 3639 7591 3689
rect 7442 3383 7557 3639
rect 7442 3333 7591 3383
rect 7735 3639 7769 3655
rect 7735 3367 7769 3383
rect 7913 3639 7947 3655
rect 7913 3367 7947 3383
rect 8091 3639 8125 3655
rect 8091 3367 8125 3383
rect 8269 3639 8303 3655
rect 8269 3367 8303 3383
rect 8447 3639 8481 3655
rect 8447 3367 8481 3383
rect 8625 3639 8659 3655
rect 8625 3367 8659 3383
rect 8803 3639 8837 3655
rect 8803 3367 8837 3383
rect 8981 3639 9015 3655
rect 8981 3367 9015 3383
rect 9159 3639 9193 3655
rect 9159 3367 9193 3383
rect 9337 3639 9371 3655
rect 9337 3367 9371 3383
rect 9515 3639 9549 3655
rect 9515 3367 9549 3383
rect 9693 3639 9727 3655
rect 9693 3367 9727 3383
rect 9871 3639 9905 3655
rect 9871 3367 9905 3383
rect 10049 3639 10278 3689
rect 10083 3383 10244 3639
rect 10049 3333 10278 3383
rect 10422 3639 10456 3655
rect 10422 3367 10456 3383
rect 10600 3639 10634 3655
rect 10600 3367 10634 3383
rect 10778 3639 10812 3655
rect 10778 3367 10812 3383
rect 10956 3639 10990 3655
rect 10956 3367 10990 3383
rect 11134 3639 11168 3655
rect 11134 3367 11168 3383
rect 11312 3639 11346 3655
rect 11312 3367 11346 3383
rect 11490 3639 11524 3655
rect 11490 3367 11524 3383
rect 11668 3639 11702 3655
rect 11668 3367 11702 3383
rect 11846 3639 11880 3655
rect 11846 3367 11880 3383
rect 12024 3639 12058 3655
rect 12024 3367 12058 3383
rect 12202 3639 12236 3655
rect 12202 3367 12236 3383
rect 12380 3639 12414 3655
rect 12380 3367 12414 3383
rect 12558 3639 12592 3655
rect 12558 3367 12592 3383
rect 12736 3639 12894 3689
rect 12770 3383 12894 3639
rect 12736 3333 12894 3383
rect 7442 3299 7637 3333
rect 7689 3299 7705 3333
rect 7799 3299 7815 3333
rect 7867 3299 7883 3333
rect 7977 3299 7993 3333
rect 8045 3299 8061 3333
rect 8155 3299 8171 3333
rect 8223 3299 8239 3333
rect 8333 3299 8349 3333
rect 8401 3299 8417 3333
rect 8511 3299 8527 3333
rect 8579 3299 8595 3333
rect 8689 3299 8705 3333
rect 8757 3299 8773 3333
rect 8867 3299 8883 3333
rect 8935 3299 8951 3333
rect 9045 3299 9061 3333
rect 9113 3299 9129 3333
rect 9223 3299 9239 3333
rect 9291 3299 9307 3333
rect 9401 3299 9417 3333
rect 9469 3299 9485 3333
rect 9579 3299 9595 3333
rect 9647 3299 9663 3333
rect 9757 3299 9773 3333
rect 9825 3299 9841 3333
rect 9935 3299 9951 3333
rect 10003 3299 10324 3333
rect 10376 3299 10392 3333
rect 10486 3299 10502 3333
rect 10554 3299 10570 3333
rect 10664 3299 10680 3333
rect 10732 3299 10748 3333
rect 10842 3299 10858 3333
rect 10910 3299 10926 3333
rect 11020 3299 11036 3333
rect 11088 3299 11104 3333
rect 11198 3299 11214 3333
rect 11266 3299 11282 3333
rect 11376 3299 11392 3333
rect 11444 3299 11460 3333
rect 11554 3299 11570 3333
rect 11622 3299 11638 3333
rect 11732 3299 11748 3333
rect 11800 3299 11816 3333
rect 11910 3299 11926 3333
rect 11978 3299 11994 3333
rect 12088 3299 12104 3333
rect 12156 3299 12172 3333
rect 12266 3299 12282 3333
rect 12334 3299 12350 3333
rect 12444 3299 12460 3333
rect 12512 3299 12528 3333
rect 12622 3299 12638 3333
rect 12690 3299 12894 3333
rect 7442 3223 7579 3299
rect 10067 3223 10261 3299
rect 12757 3223 12894 3299
rect 7442 3189 7637 3223
rect 7689 3189 7705 3223
rect 7799 3189 7815 3223
rect 7867 3189 7883 3223
rect 7977 3189 7993 3223
rect 8045 3189 8061 3223
rect 8155 3189 8171 3223
rect 8223 3189 8239 3223
rect 8333 3189 8349 3223
rect 8401 3189 8417 3223
rect 8511 3189 8527 3223
rect 8579 3189 8595 3223
rect 8689 3189 8705 3223
rect 8757 3189 8773 3223
rect 8867 3189 8883 3223
rect 8935 3189 8951 3223
rect 9045 3189 9061 3223
rect 9113 3189 9129 3223
rect 9223 3189 9239 3223
rect 9291 3189 9307 3223
rect 9401 3189 9417 3223
rect 9469 3189 9485 3223
rect 9579 3189 9595 3223
rect 9647 3189 9663 3223
rect 9757 3189 9773 3223
rect 9825 3189 9841 3223
rect 9935 3189 9951 3223
rect 10003 3189 10324 3223
rect 10376 3189 10392 3223
rect 10486 3189 10502 3223
rect 10554 3189 10570 3223
rect 10664 3189 10680 3223
rect 10732 3189 10748 3223
rect 10842 3189 10858 3223
rect 10910 3189 10926 3223
rect 11020 3189 11036 3223
rect 11088 3189 11104 3223
rect 11198 3189 11214 3223
rect 11266 3189 11282 3223
rect 11376 3189 11392 3223
rect 11444 3189 11460 3223
rect 11554 3189 11570 3223
rect 11622 3189 11638 3223
rect 11732 3189 11748 3223
rect 11800 3189 11816 3223
rect 11910 3189 11926 3223
rect 11978 3189 11994 3223
rect 12088 3189 12104 3223
rect 12156 3189 12172 3223
rect 12266 3189 12282 3223
rect 12334 3189 12350 3223
rect 12444 3189 12460 3223
rect 12512 3189 12528 3223
rect 12622 3189 12638 3223
rect 12690 3189 12894 3223
rect 7442 3139 7591 3189
rect 7442 2883 7557 3139
rect 7442 2833 7591 2883
rect 7735 3139 7769 3155
rect 7735 2867 7769 2883
rect 7913 3139 7947 3155
rect 7913 2867 7947 2883
rect 8091 3139 8125 3155
rect 8091 2867 8125 2883
rect 8269 3139 8303 3155
rect 8269 2867 8303 2883
rect 8447 3139 8481 3155
rect 8447 2867 8481 2883
rect 8625 3139 8659 3155
rect 8625 2867 8659 2883
rect 8803 3139 8837 3155
rect 8803 2867 8837 2883
rect 8981 3139 9015 3155
rect 8981 2867 9015 2883
rect 9159 3139 9193 3155
rect 9159 2867 9193 2883
rect 9337 3139 9371 3155
rect 9337 2867 9371 2883
rect 9515 3139 9549 3155
rect 9515 2867 9549 2883
rect 9693 3139 9727 3155
rect 9693 2867 9727 2883
rect 9871 3139 9905 3155
rect 9871 2867 9905 2883
rect 10049 3139 10278 3189
rect 10083 2883 10244 3139
rect 10049 2833 10278 2883
rect 10422 3139 10456 3155
rect 10422 2867 10456 2883
rect 10600 3139 10634 3155
rect 10600 2867 10634 2883
rect 10778 3139 10812 3155
rect 10778 2867 10812 2883
rect 10956 3139 10990 3155
rect 10956 2867 10990 2883
rect 11134 3139 11168 3155
rect 11134 2867 11168 2883
rect 11312 3139 11346 3155
rect 11312 2867 11346 2883
rect 11490 3139 11524 3155
rect 11490 2867 11524 2883
rect 11668 3139 11702 3155
rect 11668 2867 11702 2883
rect 11846 3139 11880 3155
rect 11846 2867 11880 2883
rect 12024 3139 12058 3155
rect 12024 2867 12058 2883
rect 12202 3139 12236 3155
rect 12202 2867 12236 2883
rect 12380 3139 12414 3155
rect 12380 2867 12414 2883
rect 12558 3139 12592 3155
rect 12558 2867 12592 2883
rect 12736 3139 12894 3189
rect 12770 2883 12894 3139
rect 12736 2833 12894 2883
rect 7442 2799 7637 2833
rect 7689 2799 7705 2833
rect 7799 2799 7815 2833
rect 7867 2799 7883 2833
rect 7977 2799 7993 2833
rect 8045 2799 8061 2833
rect 8155 2799 8171 2833
rect 8223 2799 8239 2833
rect 8333 2799 8349 2833
rect 8401 2799 8417 2833
rect 8511 2799 8527 2833
rect 8579 2799 8595 2833
rect 8689 2799 8705 2833
rect 8757 2799 8773 2833
rect 8867 2799 8883 2833
rect 8935 2799 8951 2833
rect 9045 2799 9061 2833
rect 9113 2799 9129 2833
rect 9223 2799 9239 2833
rect 9291 2799 9307 2833
rect 9401 2799 9417 2833
rect 9469 2799 9485 2833
rect 9579 2799 9595 2833
rect 9647 2799 9663 2833
rect 9757 2799 9773 2833
rect 9825 2799 9841 2833
rect 9935 2799 9951 2833
rect 10003 2799 10324 2833
rect 10376 2799 10392 2833
rect 10486 2799 10502 2833
rect 10554 2799 10570 2833
rect 10664 2799 10680 2833
rect 10732 2799 10748 2833
rect 10842 2799 10858 2833
rect 10910 2799 10926 2833
rect 11020 2799 11036 2833
rect 11088 2799 11104 2833
rect 11198 2799 11214 2833
rect 11266 2799 11282 2833
rect 11376 2799 11392 2833
rect 11444 2799 11460 2833
rect 11554 2799 11570 2833
rect 11622 2799 11638 2833
rect 11732 2799 11748 2833
rect 11800 2799 11816 2833
rect 11910 2799 11926 2833
rect 11978 2799 11994 2833
rect 12088 2799 12104 2833
rect 12156 2799 12172 2833
rect 12266 2799 12282 2833
rect 12334 2799 12350 2833
rect 12444 2799 12460 2833
rect 12512 2799 12528 2833
rect 12622 2799 12638 2833
rect 12690 2799 12894 2833
rect 7442 2723 7579 2799
rect 10067 2723 10261 2799
rect 12757 2723 12894 2799
rect 7442 2689 7637 2723
rect 7689 2689 7705 2723
rect 7799 2689 7815 2723
rect 7867 2689 7883 2723
rect 7977 2689 7993 2723
rect 8045 2689 8061 2723
rect 8155 2689 8171 2723
rect 8223 2689 8239 2723
rect 8333 2689 8349 2723
rect 8401 2689 8417 2723
rect 8511 2689 8527 2723
rect 8579 2689 8595 2723
rect 8689 2689 8705 2723
rect 8757 2689 8773 2723
rect 8867 2689 8883 2723
rect 8935 2689 8951 2723
rect 9045 2689 9061 2723
rect 9113 2689 9129 2723
rect 9223 2689 9239 2723
rect 9291 2689 9307 2723
rect 9401 2689 9417 2723
rect 9469 2689 9485 2723
rect 9579 2689 9595 2723
rect 9647 2689 9663 2723
rect 9757 2689 9773 2723
rect 9825 2689 9841 2723
rect 9935 2689 9951 2723
rect 10003 2689 10324 2723
rect 10376 2689 10392 2723
rect 10486 2689 10502 2723
rect 10554 2689 10570 2723
rect 10664 2689 10680 2723
rect 10732 2689 10748 2723
rect 10842 2689 10858 2723
rect 10910 2689 10926 2723
rect 11020 2689 11036 2723
rect 11088 2689 11104 2723
rect 11198 2689 11214 2723
rect 11266 2689 11282 2723
rect 11376 2689 11392 2723
rect 11444 2689 11460 2723
rect 11554 2689 11570 2723
rect 11622 2689 11638 2723
rect 11732 2689 11748 2723
rect 11800 2689 11816 2723
rect 11910 2689 11926 2723
rect 11978 2689 11994 2723
rect 12088 2689 12104 2723
rect 12156 2689 12172 2723
rect 12266 2689 12282 2723
rect 12334 2689 12350 2723
rect 12444 2689 12460 2723
rect 12512 2689 12528 2723
rect 12622 2689 12638 2723
rect 12690 2689 12894 2723
rect 7442 2639 7591 2689
rect 7442 2383 7557 2639
rect 7442 2333 7591 2383
rect 7735 2639 7769 2655
rect 7735 2367 7769 2383
rect 7913 2639 7947 2655
rect 7913 2367 7947 2383
rect 8091 2639 8125 2655
rect 8091 2367 8125 2383
rect 8269 2639 8303 2655
rect 8269 2367 8303 2383
rect 8447 2639 8481 2655
rect 8447 2367 8481 2383
rect 8625 2639 8659 2655
rect 8625 2367 8659 2383
rect 8803 2639 8837 2655
rect 8803 2367 8837 2383
rect 8981 2639 9015 2655
rect 8981 2367 9015 2383
rect 9159 2639 9193 2655
rect 9159 2367 9193 2383
rect 9337 2639 9371 2655
rect 9337 2367 9371 2383
rect 9515 2639 9549 2655
rect 9515 2367 9549 2383
rect 9693 2639 9727 2655
rect 9693 2367 9727 2383
rect 9871 2639 9905 2655
rect 9871 2367 9905 2383
rect 10049 2639 10278 2689
rect 10083 2383 10244 2639
rect 10049 2333 10278 2383
rect 10422 2639 10456 2655
rect 10422 2367 10456 2383
rect 10600 2639 10634 2655
rect 10600 2367 10634 2383
rect 10778 2639 10812 2655
rect 10778 2367 10812 2383
rect 10956 2639 10990 2655
rect 10956 2367 10990 2383
rect 11134 2639 11168 2655
rect 11134 2367 11168 2383
rect 11312 2639 11346 2655
rect 11312 2367 11346 2383
rect 11490 2639 11524 2655
rect 11490 2367 11524 2383
rect 11668 2639 11702 2655
rect 11668 2367 11702 2383
rect 11846 2639 11880 2655
rect 11846 2367 11880 2383
rect 12024 2639 12058 2655
rect 12024 2367 12058 2383
rect 12202 2639 12236 2655
rect 12202 2367 12236 2383
rect 12380 2639 12414 2655
rect 12380 2367 12414 2383
rect 12558 2639 12592 2655
rect 12558 2367 12592 2383
rect 12736 2639 12894 2689
rect 12770 2383 12894 2639
rect 12736 2333 12894 2383
rect 7442 2299 7637 2333
rect 7689 2299 7705 2333
rect 7799 2299 7815 2333
rect 7867 2299 7883 2333
rect 7977 2299 7993 2333
rect 8045 2299 8061 2333
rect 8155 2299 8171 2333
rect 8223 2299 8239 2333
rect 8333 2299 8349 2333
rect 8401 2299 8417 2333
rect 8511 2299 8527 2333
rect 8579 2299 8595 2333
rect 8689 2299 8705 2333
rect 8757 2299 8773 2333
rect 8867 2299 8883 2333
rect 8935 2299 8951 2333
rect 9045 2299 9061 2333
rect 9113 2299 9129 2333
rect 9223 2299 9239 2333
rect 9291 2299 9307 2333
rect 9401 2299 9417 2333
rect 9469 2299 9485 2333
rect 9579 2299 9595 2333
rect 9647 2299 9663 2333
rect 9757 2299 9773 2333
rect 9825 2299 9841 2333
rect 9935 2299 9951 2333
rect 10003 2299 10324 2333
rect 10376 2299 10392 2333
rect 10486 2299 10502 2333
rect 10554 2299 10570 2333
rect 10664 2299 10680 2333
rect 10732 2299 10748 2333
rect 10842 2299 10858 2333
rect 10910 2299 10926 2333
rect 11020 2299 11036 2333
rect 11088 2299 11104 2333
rect 11198 2299 11214 2333
rect 11266 2299 11282 2333
rect 11376 2299 11392 2333
rect 11444 2299 11460 2333
rect 11554 2299 11570 2333
rect 11622 2299 11638 2333
rect 11732 2299 11748 2333
rect 11800 2299 11816 2333
rect 11910 2299 11926 2333
rect 11978 2299 11994 2333
rect 12088 2299 12104 2333
rect 12156 2299 12172 2333
rect 12266 2299 12282 2333
rect 12334 2299 12350 2333
rect 12444 2299 12460 2333
rect 12512 2299 12528 2333
rect 12622 2299 12638 2333
rect 12690 2299 12894 2333
rect 7442 2023 7579 2299
rect 10067 2023 10261 2299
rect 12757 2023 12894 2299
rect 7442 1989 7637 2023
rect 7689 1989 7705 2023
rect 7799 1989 7815 2023
rect 7867 1989 7883 2023
rect 7977 1989 7993 2023
rect 8045 1989 8061 2023
rect 8155 1989 8171 2023
rect 8223 1989 8239 2023
rect 8333 1989 8349 2023
rect 8401 1989 8417 2023
rect 8511 1989 8527 2023
rect 8579 1989 8595 2023
rect 8689 1989 8705 2023
rect 8757 1989 8773 2023
rect 8867 1989 8883 2023
rect 8935 1989 8951 2023
rect 9045 1989 9061 2023
rect 9113 1989 9129 2023
rect 9223 1989 9239 2023
rect 9291 1989 9307 2023
rect 9401 1989 9417 2023
rect 9469 1989 9485 2023
rect 9579 1989 9595 2023
rect 9647 1989 9663 2023
rect 9757 1989 9773 2023
rect 9825 1989 9841 2023
rect 9935 1989 9951 2023
rect 10003 1989 10324 2023
rect 10376 1989 10392 2023
rect 10486 1989 10502 2023
rect 10554 1989 10570 2023
rect 10664 1989 10680 2023
rect 10732 1989 10748 2023
rect 10842 1989 10858 2023
rect 10910 1989 10926 2023
rect 11020 1989 11036 2023
rect 11088 1989 11104 2023
rect 11198 1989 11214 2023
rect 11266 1989 11282 2023
rect 11376 1989 11392 2023
rect 11444 1989 11460 2023
rect 11554 1989 11570 2023
rect 11622 1989 11638 2023
rect 11732 1989 11748 2023
rect 11800 1989 11816 2023
rect 11910 1989 11926 2023
rect 11978 1989 11994 2023
rect 12088 1989 12104 2023
rect 12156 1989 12172 2023
rect 12266 1989 12282 2023
rect 12334 1989 12350 2023
rect 12444 1989 12460 2023
rect 12512 1989 12528 2023
rect 12622 1989 12638 2023
rect 12690 1989 12894 2023
rect 7442 1939 7591 1989
rect 7442 1683 7557 1939
rect 7442 1633 7591 1683
rect 7735 1939 7769 1955
rect 7735 1667 7769 1683
rect 7913 1939 7947 1955
rect 7913 1667 7947 1683
rect 8091 1939 8125 1955
rect 8091 1667 8125 1683
rect 8269 1939 8303 1955
rect 8269 1667 8303 1683
rect 8447 1939 8481 1955
rect 8447 1667 8481 1683
rect 8625 1939 8659 1955
rect 8625 1667 8659 1683
rect 8803 1939 8837 1955
rect 8803 1667 8837 1683
rect 8981 1939 9015 1955
rect 8981 1667 9015 1683
rect 9159 1939 9193 1955
rect 9159 1667 9193 1683
rect 9337 1939 9371 1955
rect 9337 1667 9371 1683
rect 9515 1939 9549 1955
rect 9515 1667 9549 1683
rect 9693 1939 9727 1955
rect 9693 1667 9727 1683
rect 9871 1939 9905 1955
rect 9871 1667 9905 1683
rect 10049 1939 10278 1989
rect 10083 1683 10244 1939
rect 10049 1633 10278 1683
rect 10422 1939 10456 1955
rect 10422 1667 10456 1683
rect 10600 1939 10634 1955
rect 10600 1667 10634 1683
rect 10778 1939 10812 1955
rect 10778 1667 10812 1683
rect 10956 1939 10990 1955
rect 10956 1667 10990 1683
rect 11134 1939 11168 1955
rect 11134 1667 11168 1683
rect 11312 1939 11346 1955
rect 11312 1667 11346 1683
rect 11490 1939 11524 1955
rect 11490 1667 11524 1683
rect 11668 1939 11702 1955
rect 11668 1667 11702 1683
rect 11846 1939 11880 1955
rect 11846 1667 11880 1683
rect 12024 1939 12058 1955
rect 12024 1667 12058 1683
rect 12202 1939 12236 1955
rect 12202 1667 12236 1683
rect 12380 1939 12414 1955
rect 12380 1667 12414 1683
rect 12558 1939 12592 1955
rect 12558 1667 12592 1683
rect 12736 1939 12894 1989
rect 12770 1683 12894 1939
rect 12736 1633 12894 1683
rect 7442 1599 7637 1633
rect 7689 1599 7705 1633
rect 7799 1599 7815 1633
rect 7867 1599 7883 1633
rect 7977 1599 7993 1633
rect 8045 1599 8061 1633
rect 8155 1599 8171 1633
rect 8223 1599 8239 1633
rect 8333 1599 8349 1633
rect 8401 1599 8417 1633
rect 8511 1599 8527 1633
rect 8579 1599 8595 1633
rect 8689 1599 8705 1633
rect 8757 1599 8773 1633
rect 8867 1599 8883 1633
rect 8935 1599 8951 1633
rect 9045 1599 9061 1633
rect 9113 1599 9129 1633
rect 9223 1599 9239 1633
rect 9291 1599 9307 1633
rect 9401 1599 9417 1633
rect 9469 1599 9485 1633
rect 9579 1599 9595 1633
rect 9647 1599 9663 1633
rect 9757 1599 9773 1633
rect 9825 1599 9841 1633
rect 9935 1599 9951 1633
rect 10003 1599 10324 1633
rect 10376 1599 10392 1633
rect 10486 1599 10502 1633
rect 10554 1599 10570 1633
rect 10664 1599 10680 1633
rect 10732 1599 10748 1633
rect 10842 1599 10858 1633
rect 10910 1599 10926 1633
rect 11020 1599 11036 1633
rect 11088 1599 11104 1633
rect 11198 1599 11214 1633
rect 11266 1599 11282 1633
rect 11376 1599 11392 1633
rect 11444 1599 11460 1633
rect 11554 1599 11570 1633
rect 11622 1599 11638 1633
rect 11732 1599 11748 1633
rect 11800 1599 11816 1633
rect 11910 1599 11926 1633
rect 11978 1599 11994 1633
rect 12088 1599 12104 1633
rect 12156 1599 12172 1633
rect 12266 1599 12282 1633
rect 12334 1599 12350 1633
rect 12444 1599 12460 1633
rect 12512 1599 12528 1633
rect 12622 1599 12638 1633
rect 12690 1599 12894 1633
rect 7442 1523 7579 1599
rect 10067 1523 10261 1599
rect 12757 1523 12894 1599
rect 7442 1489 7637 1523
rect 7689 1489 7705 1523
rect 7799 1489 7815 1523
rect 7867 1489 7883 1523
rect 7977 1489 7993 1523
rect 8045 1489 8061 1523
rect 8155 1489 8171 1523
rect 8223 1489 8239 1523
rect 8333 1489 8349 1523
rect 8401 1489 8417 1523
rect 8511 1489 8527 1523
rect 8579 1489 8595 1523
rect 8689 1489 8705 1523
rect 8757 1489 8773 1523
rect 8867 1489 8883 1523
rect 8935 1489 8951 1523
rect 9045 1489 9061 1523
rect 9113 1489 9129 1523
rect 9223 1489 9239 1523
rect 9291 1489 9307 1523
rect 9401 1489 9417 1523
rect 9469 1489 9485 1523
rect 9579 1489 9595 1523
rect 9647 1489 9663 1523
rect 9757 1489 9773 1523
rect 9825 1489 9841 1523
rect 9935 1489 9951 1523
rect 10003 1489 10324 1523
rect 10376 1489 10392 1523
rect 10486 1489 10502 1523
rect 10554 1489 10570 1523
rect 10664 1489 10680 1523
rect 10732 1489 10748 1523
rect 10842 1489 10858 1523
rect 10910 1489 10926 1523
rect 11020 1489 11036 1523
rect 11088 1489 11104 1523
rect 11198 1489 11214 1523
rect 11266 1489 11282 1523
rect 11376 1489 11392 1523
rect 11444 1489 11460 1523
rect 11554 1489 11570 1523
rect 11622 1489 11638 1523
rect 11732 1489 11748 1523
rect 11800 1489 11816 1523
rect 11910 1489 11926 1523
rect 11978 1489 11994 1523
rect 12088 1489 12104 1523
rect 12156 1489 12172 1523
rect 12266 1489 12282 1523
rect 12334 1489 12350 1523
rect 12444 1489 12460 1523
rect 12512 1489 12528 1523
rect 12622 1489 12638 1523
rect 12690 1489 12894 1523
rect 7442 1439 7591 1489
rect 7442 1183 7557 1439
rect 7442 1133 7591 1183
rect 7735 1439 7769 1455
rect 7735 1167 7769 1183
rect 7913 1439 7947 1455
rect 7913 1167 7947 1183
rect 8091 1439 8125 1455
rect 8091 1167 8125 1183
rect 8269 1439 8303 1455
rect 8269 1167 8303 1183
rect 8447 1439 8481 1455
rect 8447 1167 8481 1183
rect 8625 1439 8659 1455
rect 8625 1167 8659 1183
rect 8803 1439 8837 1455
rect 8803 1167 8837 1183
rect 8981 1439 9015 1455
rect 8981 1167 9015 1183
rect 9159 1439 9193 1455
rect 9159 1167 9193 1183
rect 9337 1439 9371 1455
rect 9337 1167 9371 1183
rect 9515 1439 9549 1455
rect 9515 1167 9549 1183
rect 9693 1439 9727 1455
rect 9693 1167 9727 1183
rect 9871 1439 9905 1455
rect 9871 1167 9905 1183
rect 10049 1439 10278 1489
rect 10083 1183 10244 1439
rect 10049 1133 10278 1183
rect 10422 1439 10456 1455
rect 10422 1167 10456 1183
rect 10600 1439 10634 1455
rect 10600 1167 10634 1183
rect 10778 1439 10812 1455
rect 10778 1167 10812 1183
rect 10956 1439 10990 1455
rect 10956 1167 10990 1183
rect 11134 1439 11168 1455
rect 11134 1167 11168 1183
rect 11312 1439 11346 1455
rect 11312 1167 11346 1183
rect 11490 1439 11524 1455
rect 11490 1167 11524 1183
rect 11668 1439 11702 1455
rect 11668 1167 11702 1183
rect 11846 1439 11880 1455
rect 11846 1167 11880 1183
rect 12024 1439 12058 1455
rect 12024 1167 12058 1183
rect 12202 1439 12236 1455
rect 12202 1167 12236 1183
rect 12380 1439 12414 1455
rect 12380 1167 12414 1183
rect 12558 1439 12592 1455
rect 12558 1167 12592 1183
rect 12736 1439 12894 1489
rect 12770 1183 12894 1439
rect 12736 1133 12894 1183
rect 7442 1099 7637 1133
rect 7689 1099 7705 1133
rect 7799 1099 7815 1133
rect 7867 1099 7883 1133
rect 7977 1099 7993 1133
rect 8045 1099 8061 1133
rect 8155 1099 8171 1133
rect 8223 1099 8239 1133
rect 8333 1099 8349 1133
rect 8401 1099 8417 1133
rect 8511 1099 8527 1133
rect 8579 1099 8595 1133
rect 8689 1099 8705 1133
rect 8757 1099 8773 1133
rect 8867 1099 8883 1133
rect 8935 1099 8951 1133
rect 9045 1099 9061 1133
rect 9113 1099 9129 1133
rect 9223 1099 9239 1133
rect 9291 1099 9307 1133
rect 9401 1099 9417 1133
rect 9469 1099 9485 1133
rect 9579 1099 9595 1133
rect 9647 1099 9663 1133
rect 9757 1099 9773 1133
rect 9825 1099 9841 1133
rect 9935 1099 9951 1133
rect 10003 1099 10324 1133
rect 10376 1099 10392 1133
rect 10486 1099 10502 1133
rect 10554 1099 10570 1133
rect 10664 1099 10680 1133
rect 10732 1099 10748 1133
rect 10842 1099 10858 1133
rect 10910 1099 10926 1133
rect 11020 1099 11036 1133
rect 11088 1099 11104 1133
rect 11198 1099 11214 1133
rect 11266 1099 11282 1133
rect 11376 1099 11392 1133
rect 11444 1099 11460 1133
rect 11554 1099 11570 1133
rect 11622 1099 11638 1133
rect 11732 1099 11748 1133
rect 11800 1099 11816 1133
rect 11910 1099 11926 1133
rect 11978 1099 11994 1133
rect 12088 1099 12104 1133
rect 12156 1099 12172 1133
rect 12266 1099 12282 1133
rect 12334 1099 12350 1133
rect 12444 1099 12460 1133
rect 12512 1099 12528 1133
rect 12622 1099 12638 1133
rect 12690 1099 12894 1133
rect 7442 1023 7579 1099
rect 10067 1023 10261 1099
rect 12757 1023 12894 1099
rect 7442 989 7637 1023
rect 7689 989 7705 1023
rect 7799 989 7815 1023
rect 7867 989 7883 1023
rect 7977 989 7993 1023
rect 8045 989 8061 1023
rect 8155 989 8171 1023
rect 8223 989 8239 1023
rect 8333 989 8349 1023
rect 8401 989 8417 1023
rect 8511 989 8527 1023
rect 8579 989 8595 1023
rect 8689 989 8705 1023
rect 8757 989 8773 1023
rect 8867 989 8883 1023
rect 8935 989 8951 1023
rect 9045 989 9061 1023
rect 9113 989 9129 1023
rect 9223 989 9239 1023
rect 9291 989 9307 1023
rect 9401 989 9417 1023
rect 9469 989 9485 1023
rect 9579 989 9595 1023
rect 9647 989 9663 1023
rect 9757 989 9773 1023
rect 9825 989 9841 1023
rect 9935 989 9951 1023
rect 10003 989 10324 1023
rect 10376 989 10392 1023
rect 10486 989 10502 1023
rect 10554 989 10570 1023
rect 10664 989 10680 1023
rect 10732 989 10748 1023
rect 10842 989 10858 1023
rect 10910 989 10926 1023
rect 11020 989 11036 1023
rect 11088 989 11104 1023
rect 11198 989 11214 1023
rect 11266 989 11282 1023
rect 11376 989 11392 1023
rect 11444 989 11460 1023
rect 11554 989 11570 1023
rect 11622 989 11638 1023
rect 11732 989 11748 1023
rect 11800 989 11816 1023
rect 11910 989 11926 1023
rect 11978 989 11994 1023
rect 12088 989 12104 1023
rect 12156 989 12172 1023
rect 12266 989 12282 1023
rect 12334 989 12350 1023
rect 12444 989 12460 1023
rect 12512 989 12528 1023
rect 12622 989 12638 1023
rect 12690 989 12894 1023
rect 7442 939 7591 989
rect 7442 683 7557 939
rect 7442 633 7591 683
rect 7735 939 7769 955
rect 7735 667 7769 683
rect 7913 939 7947 955
rect 7913 667 7947 683
rect 8091 939 8125 955
rect 8091 667 8125 683
rect 8269 939 8303 955
rect 8269 667 8303 683
rect 8447 939 8481 955
rect 8447 667 8481 683
rect 8625 939 8659 955
rect 8625 667 8659 683
rect 8803 939 8837 955
rect 8803 667 8837 683
rect 8981 939 9015 955
rect 8981 667 9015 683
rect 9159 939 9193 955
rect 9159 667 9193 683
rect 9337 939 9371 955
rect 9337 667 9371 683
rect 9515 939 9549 955
rect 9515 667 9549 683
rect 9693 939 9727 955
rect 9693 667 9727 683
rect 9871 939 9905 955
rect 9871 667 9905 683
rect 10049 939 10278 989
rect 10083 683 10244 939
rect 10049 633 10278 683
rect 10422 939 10456 955
rect 10422 667 10456 683
rect 10600 939 10634 955
rect 10600 667 10634 683
rect 10778 939 10812 955
rect 10778 667 10812 683
rect 10956 939 10990 955
rect 10956 667 10990 683
rect 11134 939 11168 955
rect 11134 667 11168 683
rect 11312 939 11346 955
rect 11312 667 11346 683
rect 11490 939 11524 955
rect 11490 667 11524 683
rect 11668 939 11702 955
rect 11668 667 11702 683
rect 11846 939 11880 955
rect 11846 667 11880 683
rect 12024 939 12058 955
rect 12024 667 12058 683
rect 12202 939 12236 955
rect 12202 667 12236 683
rect 12380 939 12414 955
rect 12380 667 12414 683
rect 12558 939 12592 955
rect 12558 667 12592 683
rect 12736 939 12894 989
rect 12770 683 12894 939
rect 12736 633 12894 683
rect 7442 599 7637 633
rect 7689 599 7705 633
rect 7799 599 7815 633
rect 7867 599 7883 633
rect 7977 599 7993 633
rect 8045 599 8061 633
rect 8155 599 8171 633
rect 8223 599 8239 633
rect 8333 599 8349 633
rect 8401 599 8417 633
rect 8511 599 8527 633
rect 8579 599 8595 633
rect 8689 599 8705 633
rect 8757 599 8773 633
rect 8867 599 8883 633
rect 8935 599 8951 633
rect 9045 599 9061 633
rect 9113 599 9129 633
rect 9223 599 9239 633
rect 9291 599 9307 633
rect 9401 599 9417 633
rect 9469 599 9485 633
rect 9579 599 9595 633
rect 9647 599 9663 633
rect 9757 599 9773 633
rect 9825 599 9841 633
rect 9935 599 9951 633
rect 10003 599 10324 633
rect 10376 599 10392 633
rect 10486 599 10502 633
rect 10554 599 10570 633
rect 10664 599 10680 633
rect 10732 599 10748 633
rect 10842 599 10858 633
rect 10910 599 10926 633
rect 11020 599 11036 633
rect 11088 599 11104 633
rect 11198 599 11214 633
rect 11266 599 11282 633
rect 11376 599 11392 633
rect 11444 599 11460 633
rect 11554 599 11570 633
rect 11622 599 11638 633
rect 11732 599 11748 633
rect 11800 599 11816 633
rect 11910 599 11926 633
rect 11978 599 11994 633
rect 12088 599 12104 633
rect 12156 599 12172 633
rect 12266 599 12282 633
rect 12334 599 12350 633
rect 12444 599 12460 633
rect 12512 599 12528 633
rect 12622 599 12638 633
rect 12690 599 12894 633
rect 7442 149 7579 599
rect 10067 149 10261 599
rect 12757 149 12894 599
rect -61 113 13318 149
rect 13438 5131 13575 5211
rect 18360 5145 18506 5260
rect 18360 5131 18457 5145
rect 13438 5097 13630 5131
rect 13682 5097 13698 5131
rect 13792 5097 13808 5131
rect 13860 5097 13876 5131
rect 13970 5097 13986 5131
rect 14038 5097 14054 5131
rect 14148 5097 14164 5131
rect 14216 5097 14232 5131
rect 14326 5097 14342 5131
rect 14394 5097 14410 5131
rect 14504 5097 14520 5131
rect 14572 5097 14588 5131
rect 14682 5097 14698 5131
rect 14750 5097 14766 5131
rect 14860 5097 14876 5131
rect 14928 5097 14944 5131
rect 15038 5097 15054 5131
rect 15106 5097 15122 5131
rect 15216 5097 15232 5131
rect 15284 5097 15300 5131
rect 15394 5097 15410 5131
rect 15462 5097 15478 5131
rect 15572 5097 15588 5131
rect 15640 5097 15656 5131
rect 15750 5097 15766 5131
rect 15818 5097 15834 5131
rect 15928 5097 15944 5131
rect 15996 5097 16012 5131
rect 16106 5097 16122 5131
rect 16174 5097 16190 5131
rect 16284 5097 16300 5131
rect 16352 5097 16368 5131
rect 16462 5097 16478 5131
rect 16530 5097 16546 5131
rect 16640 5097 16656 5131
rect 16708 5097 16724 5131
rect 16818 5097 16834 5131
rect 16886 5097 16902 5131
rect 16996 5097 17012 5131
rect 17064 5097 17080 5131
rect 17174 5097 17190 5131
rect 17242 5097 17258 5131
rect 17352 5097 17368 5131
rect 17420 5097 17436 5131
rect 17530 5097 17546 5131
rect 17598 5097 17614 5131
rect 17708 5097 17724 5131
rect 17776 5097 17792 5131
rect 17886 5097 17902 5131
rect 17954 5097 17970 5131
rect 18064 5097 18080 5131
rect 18132 5097 18148 5131
rect 18242 5097 18258 5131
rect 18310 5097 18457 5131
rect 13438 5047 13584 5097
rect 13438 4791 13550 5047
rect 13438 4741 13584 4791
rect 13728 5047 13762 5063
rect 13728 4775 13762 4791
rect 13906 5047 13940 5063
rect 13906 4775 13940 4791
rect 14084 5047 14118 5063
rect 14084 4775 14118 4791
rect 14262 5047 14296 5063
rect 14262 4775 14296 4791
rect 14440 5047 14474 5063
rect 14440 4775 14474 4791
rect 14618 5047 14652 5063
rect 14618 4775 14652 4791
rect 14796 5047 14830 5063
rect 14796 4775 14830 4791
rect 14974 5047 15008 5063
rect 14974 4775 15008 4791
rect 15152 5047 15186 5063
rect 15152 4775 15186 4791
rect 15330 5047 15364 5063
rect 15330 4775 15364 4791
rect 15508 5047 15542 5063
rect 15508 4775 15542 4791
rect 15686 5047 15720 5063
rect 15686 4775 15720 4791
rect 15864 5047 15898 5063
rect 15864 4775 15898 4791
rect 16042 5047 16076 5063
rect 16042 4775 16076 4791
rect 16220 5047 16254 5063
rect 16220 4775 16254 4791
rect 16398 5047 16432 5063
rect 16398 4775 16432 4791
rect 16576 5047 16610 5063
rect 16576 4775 16610 4791
rect 16754 5047 16788 5063
rect 16754 4775 16788 4791
rect 16932 5047 16966 5063
rect 16932 4775 16966 4791
rect 17110 5047 17144 5063
rect 17110 4775 17144 4791
rect 17288 5047 17322 5063
rect 17288 4775 17322 4791
rect 17466 5047 17500 5063
rect 17466 4775 17500 4791
rect 17644 5047 17678 5063
rect 17644 4775 17678 4791
rect 17822 5047 17856 5063
rect 17822 4775 17856 4791
rect 18000 5047 18034 5063
rect 18000 4775 18034 4791
rect 18178 5047 18212 5063
rect 18178 4775 18212 4791
rect 18356 5047 18457 5097
rect 18390 4791 18457 5047
rect 18356 4741 18457 4791
rect 13438 4707 13630 4741
rect 13682 4707 13698 4741
rect 13792 4707 13808 4741
rect 13860 4707 13876 4741
rect 13970 4707 13986 4741
rect 14038 4707 14054 4741
rect 14148 4707 14164 4741
rect 14216 4707 14232 4741
rect 14326 4707 14342 4741
rect 14394 4707 14410 4741
rect 14504 4707 14520 4741
rect 14572 4707 14588 4741
rect 14682 4707 14698 4741
rect 14750 4707 14766 4741
rect 14860 4707 14876 4741
rect 14928 4707 14944 4741
rect 15038 4707 15054 4741
rect 15106 4707 15122 4741
rect 15216 4707 15232 4741
rect 15284 4707 15300 4741
rect 15394 4707 15410 4741
rect 15462 4707 15478 4741
rect 15572 4707 15588 4741
rect 15640 4707 15656 4741
rect 15750 4707 15766 4741
rect 15818 4707 15834 4741
rect 15928 4707 15944 4741
rect 15996 4707 16012 4741
rect 16106 4707 16122 4741
rect 16174 4707 16190 4741
rect 16284 4707 16300 4741
rect 16352 4707 16368 4741
rect 16462 4707 16478 4741
rect 16530 4707 16546 4741
rect 16640 4707 16656 4741
rect 16708 4707 16724 4741
rect 16818 4707 16834 4741
rect 16886 4707 16902 4741
rect 16996 4707 17012 4741
rect 17064 4707 17080 4741
rect 17174 4707 17190 4741
rect 17242 4707 17258 4741
rect 17352 4707 17368 4741
rect 17420 4707 17436 4741
rect 17530 4707 17546 4741
rect 17598 4707 17614 4741
rect 17708 4707 17724 4741
rect 17776 4707 17792 4741
rect 17886 4707 17902 4741
rect 17954 4707 17970 4741
rect 18064 4707 18080 4741
rect 18132 4707 18148 4741
rect 18242 4707 18258 4741
rect 18310 4707 18457 4741
rect 13438 4631 13575 4707
rect 18360 4631 18457 4707
rect 13438 4597 13630 4631
rect 13682 4597 13698 4631
rect 13792 4597 13808 4631
rect 13860 4597 13876 4631
rect 13970 4597 13986 4631
rect 14038 4597 14054 4631
rect 14148 4597 14164 4631
rect 14216 4597 14232 4631
rect 14326 4597 14342 4631
rect 14394 4597 14410 4631
rect 14504 4597 14520 4631
rect 14572 4597 14588 4631
rect 14682 4597 14698 4631
rect 14750 4597 14766 4631
rect 14860 4597 14876 4631
rect 14928 4597 14944 4631
rect 15038 4597 15054 4631
rect 15106 4597 15122 4631
rect 15216 4597 15232 4631
rect 15284 4597 15300 4631
rect 15394 4597 15410 4631
rect 15462 4597 15478 4631
rect 15572 4597 15588 4631
rect 15640 4597 15656 4631
rect 15750 4597 15766 4631
rect 15818 4597 15834 4631
rect 15928 4597 15944 4631
rect 15996 4597 16012 4631
rect 16106 4597 16122 4631
rect 16174 4597 16190 4631
rect 16284 4597 16300 4631
rect 16352 4597 16368 4631
rect 16462 4597 16478 4631
rect 16530 4597 16546 4631
rect 16640 4597 16656 4631
rect 16708 4597 16724 4631
rect 16818 4597 16834 4631
rect 16886 4597 16902 4631
rect 16996 4597 17012 4631
rect 17064 4597 17080 4631
rect 17174 4597 17190 4631
rect 17242 4597 17258 4631
rect 17352 4597 17368 4631
rect 17420 4597 17436 4631
rect 17530 4597 17546 4631
rect 17598 4597 17614 4631
rect 17708 4597 17724 4631
rect 17776 4597 17792 4631
rect 17886 4597 17902 4631
rect 17954 4597 17970 4631
rect 18064 4597 18080 4631
rect 18132 4597 18148 4631
rect 18242 4597 18258 4631
rect 18310 4597 18457 4631
rect 13438 4547 13584 4597
rect 13438 4291 13550 4547
rect 13438 4241 13584 4291
rect 13728 4547 13762 4563
rect 13728 4275 13762 4291
rect 13906 4547 13940 4563
rect 13906 4275 13940 4291
rect 14084 4547 14118 4563
rect 14084 4275 14118 4291
rect 14262 4547 14296 4563
rect 14262 4275 14296 4291
rect 14440 4547 14474 4563
rect 14440 4275 14474 4291
rect 14618 4547 14652 4563
rect 14618 4275 14652 4291
rect 14796 4547 14830 4563
rect 14796 4275 14830 4291
rect 14974 4547 15008 4563
rect 14974 4275 15008 4291
rect 15152 4547 15186 4563
rect 15152 4275 15186 4291
rect 15330 4547 15364 4563
rect 15330 4275 15364 4291
rect 15508 4547 15542 4563
rect 15508 4275 15542 4291
rect 15686 4547 15720 4563
rect 15686 4275 15720 4291
rect 15864 4547 15898 4563
rect 15864 4275 15898 4291
rect 16042 4547 16076 4563
rect 16042 4275 16076 4291
rect 16220 4547 16254 4563
rect 16220 4275 16254 4291
rect 16398 4547 16432 4563
rect 16398 4275 16432 4291
rect 16576 4547 16610 4563
rect 16576 4275 16610 4291
rect 16754 4547 16788 4563
rect 16754 4275 16788 4291
rect 16932 4547 16966 4563
rect 16932 4275 16966 4291
rect 17110 4547 17144 4563
rect 17110 4275 17144 4291
rect 17288 4547 17322 4563
rect 17288 4275 17322 4291
rect 17466 4547 17500 4563
rect 17466 4275 17500 4291
rect 17644 4547 17678 4563
rect 17644 4275 17678 4291
rect 17822 4547 17856 4563
rect 17822 4275 17856 4291
rect 18000 4547 18034 4563
rect 18000 4275 18034 4291
rect 18178 4547 18212 4563
rect 18178 4275 18212 4291
rect 18356 4547 18457 4597
rect 18390 4291 18457 4547
rect 18356 4241 18457 4291
rect 13438 4207 13630 4241
rect 13682 4207 13698 4241
rect 13792 4207 13808 4241
rect 13860 4207 13876 4241
rect 13970 4207 13986 4241
rect 14038 4207 14054 4241
rect 14148 4207 14164 4241
rect 14216 4207 14232 4241
rect 14326 4207 14342 4241
rect 14394 4207 14410 4241
rect 14504 4207 14520 4241
rect 14572 4207 14588 4241
rect 14682 4207 14698 4241
rect 14750 4207 14766 4241
rect 14860 4207 14876 4241
rect 14928 4207 14944 4241
rect 15038 4207 15054 4241
rect 15106 4207 15122 4241
rect 15216 4207 15232 4241
rect 15284 4207 15300 4241
rect 15394 4207 15410 4241
rect 15462 4207 15478 4241
rect 15572 4207 15588 4241
rect 15640 4207 15656 4241
rect 15750 4207 15766 4241
rect 15818 4207 15834 4241
rect 15928 4207 15944 4241
rect 15996 4207 16012 4241
rect 16106 4207 16122 4241
rect 16174 4207 16190 4241
rect 16284 4207 16300 4241
rect 16352 4207 16368 4241
rect 16462 4207 16478 4241
rect 16530 4207 16546 4241
rect 16640 4207 16656 4241
rect 16708 4207 16724 4241
rect 16818 4207 16834 4241
rect 16886 4207 16902 4241
rect 16996 4207 17012 4241
rect 17064 4207 17080 4241
rect 17174 4207 17190 4241
rect 17242 4207 17258 4241
rect 17352 4207 17368 4241
rect 17420 4207 17436 4241
rect 17530 4207 17546 4241
rect 17598 4207 17614 4241
rect 17708 4207 17724 4241
rect 17776 4207 17792 4241
rect 17886 4207 17902 4241
rect 17954 4207 17970 4241
rect 18064 4207 18080 4241
rect 18132 4207 18148 4241
rect 18242 4207 18258 4241
rect 18310 4207 18457 4241
rect 13438 3474 13575 4207
rect 17108 3593 17188 3627
rect 17240 3593 17256 3627
rect 17350 3593 17366 3627
rect 17418 3593 17434 3627
rect 17528 3593 17544 3627
rect 17596 3593 17612 3627
rect 17706 3593 17722 3627
rect 17774 3593 17854 3627
rect 17108 3543 17142 3593
rect 13438 3346 17108 3474
rect 13438 2499 13575 3346
rect 13740 2588 13756 2622
rect 13808 2588 13824 2622
rect 14032 2588 14048 2622
rect 14100 2588 14116 2622
rect 14324 2588 14340 2622
rect 14392 2588 14408 2622
rect 14616 2588 14632 2622
rect 14684 2588 14700 2622
rect 14908 2588 14924 2622
rect 14976 2588 14992 2622
rect 15200 2588 15216 2622
rect 15268 2588 15284 2622
rect 15492 2588 15508 2622
rect 15560 2588 15576 2622
rect 15639 2554 15767 3346
rect 13676 2538 13710 2554
rect 13438 2362 13676 2499
rect 13438 1982 13575 2362
rect 13676 2266 13710 2282
rect 13854 2538 13888 2554
rect 13854 2266 13888 2282
rect 13968 2538 14002 2554
rect 13968 2266 14002 2282
rect 14146 2538 14180 2554
rect 14146 2266 14180 2282
rect 14260 2538 14294 2554
rect 14260 2266 14294 2282
rect 14438 2538 14472 2554
rect 14438 2266 14472 2282
rect 14552 2538 14586 2554
rect 14552 2266 14586 2282
rect 14730 2538 14764 2554
rect 14730 2266 14764 2282
rect 14844 2538 14878 2554
rect 14844 2266 14878 2282
rect 15022 2538 15056 2554
rect 15022 2266 15056 2282
rect 15136 2538 15170 2554
rect 15136 2266 15170 2282
rect 15314 2538 15348 2554
rect 15314 2266 15348 2282
rect 15428 2538 15462 2554
rect 15428 2266 15462 2282
rect 15606 2538 15767 2554
rect 15640 2282 15767 2538
rect 15606 2266 15767 2282
rect 13740 2198 13756 2232
rect 13808 2198 13824 2232
rect 14032 2198 14048 2232
rect 14100 2198 14116 2232
rect 14324 2198 14340 2232
rect 14392 2198 14408 2232
rect 14616 2198 14632 2232
rect 14684 2198 14700 2232
rect 14908 2198 14924 2232
rect 14976 2198 14992 2232
rect 15200 2198 15216 2232
rect 15268 2198 15284 2232
rect 15492 2198 15508 2232
rect 15560 2198 15576 2232
rect 13740 2090 13756 2124
rect 13808 2090 13824 2124
rect 14032 2090 14048 2124
rect 14100 2090 14116 2124
rect 14324 2090 14340 2124
rect 14392 2090 14408 2124
rect 14616 2090 14632 2124
rect 14684 2090 14700 2124
rect 14908 2090 14924 2124
rect 14976 2090 14992 2124
rect 15200 2090 15216 2124
rect 15268 2090 15284 2124
rect 15492 2090 15508 2124
rect 15560 2090 15576 2124
rect 15639 2056 15767 2266
rect 13676 2040 13710 2056
rect 13438 1845 13676 1982
rect 13438 1496 13575 1845
rect 13676 1768 13710 1784
rect 13854 2040 13888 2056
rect 13854 1768 13888 1784
rect 13968 2040 14002 2056
rect 13968 1768 14002 1784
rect 14146 2040 14180 2056
rect 14146 1768 14180 1784
rect 14260 2040 14294 2056
rect 14260 1768 14294 1784
rect 14438 2040 14472 2056
rect 14438 1768 14472 1784
rect 14552 2040 14586 2056
rect 14552 1768 14586 1784
rect 14730 2040 14764 2056
rect 14730 1768 14764 1784
rect 14844 2040 14878 2056
rect 14844 1768 14878 1784
rect 15022 2040 15056 2056
rect 15022 1768 15056 1784
rect 15136 2040 15170 2056
rect 15136 1768 15170 1784
rect 15314 2040 15348 2056
rect 15314 1768 15348 1784
rect 15428 2040 15462 2056
rect 15428 1768 15462 1784
rect 15606 2040 15767 2056
rect 15640 1784 15767 2040
rect 15606 1768 15767 1784
rect 13740 1700 13756 1734
rect 13808 1700 13824 1734
rect 14032 1700 14048 1734
rect 14100 1700 14116 1734
rect 14324 1700 14340 1734
rect 14392 1700 14408 1734
rect 14616 1700 14632 1734
rect 14684 1700 14700 1734
rect 14908 1700 14924 1734
rect 14976 1700 14992 1734
rect 15200 1700 15216 1734
rect 15268 1700 15284 1734
rect 15492 1700 15508 1734
rect 15560 1700 15576 1734
rect 13740 1592 13756 1626
rect 13808 1592 13824 1626
rect 14032 1592 14048 1626
rect 14100 1592 14116 1626
rect 14324 1592 14340 1626
rect 14392 1592 14408 1626
rect 14616 1592 14632 1626
rect 14684 1592 14700 1626
rect 14908 1592 14924 1626
rect 14976 1592 14992 1626
rect 15200 1592 15216 1626
rect 15268 1592 15284 1626
rect 15492 1592 15508 1626
rect 15560 1592 15576 1626
rect 15639 1558 15767 1768
rect 13676 1542 13710 1558
rect 13438 1359 13676 1496
rect 13438 994 13575 1359
rect 13676 1270 13710 1286
rect 13854 1542 13888 1558
rect 13854 1270 13888 1286
rect 13968 1542 14002 1558
rect 13968 1270 14002 1286
rect 14146 1542 14180 1558
rect 14146 1270 14180 1286
rect 14260 1542 14294 1558
rect 14260 1270 14294 1286
rect 14438 1542 14472 1558
rect 14438 1270 14472 1286
rect 14552 1542 14586 1558
rect 14552 1270 14586 1286
rect 14730 1542 14764 1558
rect 14730 1270 14764 1286
rect 14844 1542 14878 1558
rect 14844 1270 14878 1286
rect 15022 1542 15056 1558
rect 15022 1270 15056 1286
rect 15136 1542 15170 1558
rect 15136 1270 15170 1286
rect 15314 1542 15348 1558
rect 15314 1270 15348 1286
rect 15428 1542 15462 1558
rect 15428 1270 15462 1286
rect 15606 1542 15767 1558
rect 15640 1286 15767 1542
rect 15606 1270 15767 1286
rect 13740 1202 13756 1236
rect 13808 1202 13824 1236
rect 14032 1202 14048 1236
rect 14100 1202 14116 1236
rect 14324 1202 14340 1236
rect 14392 1202 14408 1236
rect 14616 1202 14632 1236
rect 14684 1202 14700 1236
rect 14908 1202 14924 1236
rect 14976 1202 14992 1236
rect 15200 1202 15216 1236
rect 15268 1202 15284 1236
rect 15492 1202 15508 1236
rect 15560 1202 15576 1236
rect 13740 1094 13756 1128
rect 13808 1094 13824 1128
rect 14032 1094 14048 1128
rect 14100 1094 14116 1128
rect 14324 1094 14340 1128
rect 14392 1094 14408 1128
rect 14616 1094 14632 1128
rect 14684 1094 14700 1128
rect 14908 1094 14924 1128
rect 14976 1094 14992 1128
rect 15200 1094 15216 1128
rect 15268 1094 15284 1128
rect 15492 1094 15508 1128
rect 15560 1094 15576 1128
rect 15639 1060 15767 1270
rect 13676 1044 13710 1060
rect 13438 857 13676 994
rect 13438 632 13575 857
rect 13676 772 13710 788
rect 13854 1044 13888 1060
rect 13854 772 13888 788
rect 13968 1044 14002 1060
rect 13968 772 14002 788
rect 14146 1044 14180 1060
rect 14146 772 14180 788
rect 14260 1044 14294 1060
rect 14260 772 14294 788
rect 14438 1044 14472 1060
rect 14438 772 14472 788
rect 14552 1044 14586 1060
rect 14552 772 14586 788
rect 14730 1044 14764 1060
rect 14730 772 14764 788
rect 14844 1044 14878 1060
rect 14844 772 14878 788
rect 15022 1044 15056 1060
rect 15022 772 15056 788
rect 15136 1044 15170 1060
rect 15136 772 15170 788
rect 15314 1044 15348 1060
rect 15314 772 15348 788
rect 15428 1044 15462 1060
rect 15428 772 15462 788
rect 15606 1044 15767 1060
rect 15640 788 15767 1044
rect 15606 772 15767 788
rect 13740 704 13756 738
rect 13808 704 13824 738
rect 14032 704 14048 738
rect 14100 704 14116 738
rect 14324 704 14340 738
rect 14392 704 14408 738
rect 14616 704 14632 738
rect 14684 704 14700 738
rect 14908 704 14924 738
rect 14976 704 14992 738
rect 15200 704 15216 738
rect 15268 704 15284 738
rect 15492 704 15508 738
rect 15560 704 15576 738
rect 15639 632 15767 772
rect 13438 614 15767 632
rect 13438 613 15279 614
rect 13438 516 14109 613
rect 14212 517 15279 613
rect 15382 517 15767 614
rect 14212 516 15767 517
rect 13438 504 15767 516
rect 13438 149 13575 504
rect 15639 149 15767 504
rect 16279 2688 16407 3346
rect 17108 3237 17142 3287
rect 17286 3543 17320 3559
rect 17286 3271 17320 3287
rect 17464 3543 17498 3559
rect 17464 3271 17498 3287
rect 17642 3543 17676 3559
rect 17642 3271 17676 3287
rect 17820 3543 17854 3593
rect 18360 3474 18457 4207
rect 17854 3346 18457 3474
rect 17820 3237 17854 3287
rect 17108 3203 17188 3237
rect 17240 3203 17256 3237
rect 17350 3203 17366 3237
rect 17418 3203 17434 3237
rect 17528 3203 17544 3237
rect 17596 3203 17612 3237
rect 17706 3203 17722 3237
rect 17774 3203 17854 3237
rect 18360 2688 18457 3346
rect 16279 2654 16474 2688
rect 16526 2654 16542 2688
rect 16636 2654 16652 2688
rect 16704 2654 16720 2688
rect 16814 2654 16830 2688
rect 16882 2654 16898 2688
rect 16992 2654 17008 2688
rect 17060 2654 17076 2688
rect 17170 2654 17186 2688
rect 17238 2654 17254 2688
rect 17348 2654 17364 2688
rect 17416 2654 17432 2688
rect 17526 2654 17542 2688
rect 17594 2654 17610 2688
rect 17704 2654 17720 2688
rect 17772 2654 17788 2688
rect 17882 2654 17898 2688
rect 17950 2654 17966 2688
rect 18060 2654 18076 2688
rect 18128 2654 18144 2688
rect 18238 2654 18254 2688
rect 18306 2654 18457 2688
rect 16279 2604 16428 2654
rect 16279 2348 16394 2604
rect 16279 2298 16428 2348
rect 16572 2604 16606 2620
rect 16572 2332 16606 2348
rect 16750 2604 16784 2620
rect 16750 2332 16784 2348
rect 16928 2604 16962 2620
rect 16928 2332 16962 2348
rect 17106 2604 17140 2620
rect 17106 2332 17140 2348
rect 17284 2604 17318 2620
rect 17284 2332 17318 2348
rect 17462 2604 17496 2620
rect 17462 2332 17496 2348
rect 17640 2604 17674 2620
rect 17640 2332 17674 2348
rect 17818 2604 17852 2620
rect 17818 2332 17852 2348
rect 17996 2604 18030 2620
rect 17996 2332 18030 2348
rect 18174 2604 18208 2620
rect 18174 2332 18208 2348
rect 18352 2604 18457 2654
rect 18386 2348 18457 2604
rect 18352 2298 18457 2348
rect 16279 2264 16474 2298
rect 16526 2264 16542 2298
rect 16636 2264 16652 2298
rect 16704 2264 16720 2298
rect 16814 2264 16830 2298
rect 16882 2264 16898 2298
rect 16992 2264 17008 2298
rect 17060 2264 17076 2298
rect 17170 2264 17186 2298
rect 17238 2264 17254 2298
rect 17348 2264 17364 2298
rect 17416 2264 17432 2298
rect 17526 2264 17542 2298
rect 17594 2264 17610 2298
rect 17704 2264 17720 2298
rect 17772 2264 17788 2298
rect 17882 2264 17898 2298
rect 17950 2264 17966 2298
rect 18060 2264 18076 2298
rect 18128 2264 18144 2298
rect 18238 2264 18254 2298
rect 18306 2264 18457 2298
rect 16279 2188 16407 2264
rect 18360 2188 18457 2264
rect 16279 2154 16474 2188
rect 16526 2154 16542 2188
rect 16636 2154 16652 2188
rect 16704 2154 16720 2188
rect 16814 2154 16830 2188
rect 16882 2154 16898 2188
rect 16992 2154 17008 2188
rect 17060 2154 17076 2188
rect 17170 2154 17186 2188
rect 17238 2154 17254 2188
rect 17348 2154 17364 2188
rect 17416 2154 17432 2188
rect 17526 2154 17542 2188
rect 17594 2154 17610 2188
rect 17704 2154 17720 2188
rect 17772 2154 17788 2188
rect 17882 2154 17898 2188
rect 17950 2154 17966 2188
rect 18060 2154 18076 2188
rect 18128 2154 18144 2188
rect 18238 2154 18254 2188
rect 18306 2154 18457 2188
rect 16279 2104 16428 2154
rect 16279 1848 16394 2104
rect 16279 1798 16428 1848
rect 16572 2104 16606 2120
rect 16572 1832 16606 1848
rect 16750 2104 16784 2120
rect 16750 1832 16784 1848
rect 16928 2104 16962 2120
rect 16928 1832 16962 1848
rect 17106 2104 17140 2120
rect 17106 1832 17140 1848
rect 17284 2104 17318 2120
rect 17284 1832 17318 1848
rect 17462 2104 17496 2120
rect 17462 1832 17496 1848
rect 17640 2104 17674 2120
rect 17640 1832 17674 1848
rect 17818 2104 17852 2120
rect 17818 1832 17852 1848
rect 17996 2104 18030 2120
rect 17996 1832 18030 1848
rect 18174 2104 18208 2120
rect 18174 1832 18208 1848
rect 18352 2104 18457 2154
rect 18386 1848 18457 2104
rect 18352 1798 18457 1848
rect 16279 1764 16474 1798
rect 16526 1764 16542 1798
rect 16636 1764 16652 1798
rect 16704 1764 16720 1798
rect 16814 1764 16830 1798
rect 16882 1764 16898 1798
rect 16992 1764 17008 1798
rect 17060 1764 17076 1798
rect 17170 1764 17186 1798
rect 17238 1764 17254 1798
rect 17348 1764 17364 1798
rect 17416 1764 17432 1798
rect 17526 1764 17542 1798
rect 17594 1764 17610 1798
rect 17704 1764 17720 1798
rect 17772 1764 17788 1798
rect 17882 1764 17898 1798
rect 17950 1764 17966 1798
rect 18060 1764 18076 1798
rect 18128 1764 18144 1798
rect 18238 1764 18254 1798
rect 18306 1764 18457 1798
rect 16279 1628 16407 1764
rect 18360 1628 18457 1764
rect 16279 1594 16474 1628
rect 16526 1594 16542 1628
rect 16636 1594 16652 1628
rect 16704 1594 16720 1628
rect 16814 1594 16830 1628
rect 16882 1594 16898 1628
rect 16992 1594 17008 1628
rect 17060 1594 17076 1628
rect 17170 1594 17186 1628
rect 17238 1594 17254 1628
rect 17348 1594 17364 1628
rect 17416 1594 17432 1628
rect 17526 1594 17542 1628
rect 17594 1594 17610 1628
rect 17704 1594 17720 1628
rect 17772 1594 17788 1628
rect 17882 1594 17898 1628
rect 17950 1594 17966 1628
rect 18060 1594 18076 1628
rect 18128 1594 18144 1628
rect 18238 1594 18254 1628
rect 18306 1594 18457 1628
rect 16279 1544 16428 1594
rect 16279 1288 16394 1544
rect 16279 1238 16428 1288
rect 16572 1544 16606 1560
rect 16572 1272 16606 1288
rect 16750 1544 16784 1560
rect 16750 1272 16784 1288
rect 16928 1544 16962 1560
rect 16928 1272 16962 1288
rect 17106 1544 17140 1560
rect 17106 1272 17140 1288
rect 17284 1544 17318 1560
rect 17284 1272 17318 1288
rect 17462 1544 17496 1560
rect 17462 1272 17496 1288
rect 17640 1544 17674 1560
rect 17640 1272 17674 1288
rect 17818 1544 17852 1560
rect 17818 1272 17852 1288
rect 17996 1544 18030 1560
rect 17996 1272 18030 1288
rect 18174 1544 18208 1560
rect 18174 1272 18208 1288
rect 18352 1544 18457 1594
rect 18386 1288 18457 1544
rect 18352 1238 18457 1288
rect 16279 1204 16474 1238
rect 16526 1204 16542 1238
rect 16636 1204 16652 1238
rect 16704 1204 16720 1238
rect 16814 1204 16830 1238
rect 16882 1204 16898 1238
rect 16992 1204 17008 1238
rect 17060 1204 17076 1238
rect 17170 1204 17186 1238
rect 17238 1204 17254 1238
rect 17348 1204 17364 1238
rect 17416 1204 17432 1238
rect 17526 1204 17542 1238
rect 17594 1204 17610 1238
rect 17704 1204 17720 1238
rect 17772 1204 17788 1238
rect 17882 1204 17898 1238
rect 17950 1204 17966 1238
rect 18060 1204 18076 1238
rect 18128 1204 18144 1238
rect 18238 1204 18254 1238
rect 18306 1204 18457 1238
rect 16279 1128 16407 1204
rect 18360 1128 18457 1204
rect 16279 1094 16474 1128
rect 16526 1094 16542 1128
rect 16636 1094 16652 1128
rect 16704 1094 16720 1128
rect 16814 1094 16830 1128
rect 16882 1094 16898 1128
rect 16992 1094 17008 1128
rect 17060 1094 17076 1128
rect 17170 1094 17186 1128
rect 17238 1094 17254 1128
rect 17348 1094 17364 1128
rect 17416 1094 17432 1128
rect 17526 1094 17542 1128
rect 17594 1094 17610 1128
rect 17704 1094 17720 1128
rect 17772 1094 17788 1128
rect 17882 1094 17898 1128
rect 17950 1094 17966 1128
rect 18060 1094 18076 1128
rect 18128 1094 18144 1128
rect 18238 1094 18254 1128
rect 18306 1094 18457 1128
rect 16279 1044 16428 1094
rect 16279 788 16394 1044
rect 16279 738 16428 788
rect 16572 1044 16606 1060
rect 16572 772 16606 788
rect 16750 1044 16784 1060
rect 16750 772 16784 788
rect 16928 1044 16962 1060
rect 16928 772 16962 788
rect 17106 1044 17140 1060
rect 17106 772 17140 788
rect 17284 1044 17318 1060
rect 17284 772 17318 788
rect 17462 1044 17496 1060
rect 17462 772 17496 788
rect 17640 1044 17674 1060
rect 17640 772 17674 788
rect 17818 1044 17852 1060
rect 17818 772 17852 788
rect 17996 1044 18030 1060
rect 17996 772 18030 788
rect 18174 1044 18208 1060
rect 18174 772 18208 788
rect 18352 1044 18457 1094
rect 18386 788 18457 1044
rect 18352 738 18457 788
rect 16279 704 16474 738
rect 16526 704 16542 738
rect 16636 704 16652 738
rect 16704 704 16720 738
rect 16814 704 16830 738
rect 16882 704 16898 738
rect 16992 704 17008 738
rect 17060 704 17076 738
rect 17170 704 17186 738
rect 17238 704 17254 738
rect 17348 704 17364 738
rect 17416 704 17432 738
rect 17526 704 17542 738
rect 17594 704 17610 738
rect 17704 704 17720 738
rect 17772 704 17788 738
rect 17882 704 17898 738
rect 17950 704 17966 738
rect 18060 704 18076 738
rect 18128 704 18144 738
rect 18238 704 18254 738
rect 18306 704 18457 738
rect 16279 149 16407 704
rect 16529 611 16657 630
rect 16529 524 16547 611
rect 16640 524 16657 611
rect 16529 149 16657 524
rect 17948 600 18076 621
rect 17948 513 17969 600
rect 18062 513 18076 600
rect 17948 149 18076 513
rect 18360 149 18457 704
rect 18888 5224 19016 5228
rect 21891 5224 22019 5236
rect 18888 5190 18991 5224
rect 21909 5190 22019 5224
rect 18888 5128 19016 5190
rect 18888 3198 18895 5128
rect 18929 5122 19016 5128
rect 21891 5128 22019 5190
rect 21891 5122 21971 5128
rect 18929 5088 19089 5122
rect 19141 5088 19157 5122
rect 19251 5088 19267 5122
rect 19319 5088 19335 5122
rect 19429 5088 19445 5122
rect 19497 5088 19513 5122
rect 19607 5088 19623 5122
rect 19675 5088 19691 5122
rect 19785 5088 19801 5122
rect 19853 5088 19869 5122
rect 19963 5088 19979 5122
rect 20031 5088 20047 5122
rect 20141 5088 20157 5122
rect 20209 5088 20225 5122
rect 20319 5088 20335 5122
rect 20387 5088 20403 5122
rect 20497 5088 20513 5122
rect 20565 5088 20581 5122
rect 20675 5088 20691 5122
rect 20743 5088 20759 5122
rect 20853 5088 20869 5122
rect 20921 5088 20937 5122
rect 21031 5088 21047 5122
rect 21099 5088 21115 5122
rect 21209 5088 21225 5122
rect 21277 5088 21293 5122
rect 21387 5088 21403 5122
rect 21455 5088 21471 5122
rect 21565 5088 21581 5122
rect 21633 5088 21649 5122
rect 21743 5088 21759 5122
rect 21811 5088 21971 5122
rect 18929 5038 19043 5088
rect 18929 4782 19009 5038
rect 18929 4732 19043 4782
rect 19187 5038 19221 5054
rect 19187 4766 19221 4782
rect 19365 5038 19399 5054
rect 19365 4766 19399 4782
rect 19543 5038 19577 5054
rect 19543 4766 19577 4782
rect 19721 5038 19755 5054
rect 19721 4766 19755 4782
rect 19899 5038 19933 5054
rect 19899 4766 19933 4782
rect 20077 5038 20111 5054
rect 20077 4766 20111 4782
rect 20255 5038 20289 5054
rect 20255 4766 20289 4782
rect 20433 5038 20467 5054
rect 20433 4766 20467 4782
rect 20611 5038 20645 5054
rect 20611 4766 20645 4782
rect 20789 5038 20823 5054
rect 20789 4766 20823 4782
rect 20967 5038 21001 5054
rect 20967 4766 21001 4782
rect 21145 5038 21179 5054
rect 21145 4766 21179 4782
rect 21323 5038 21357 5054
rect 21323 4766 21357 4782
rect 21501 5038 21535 5054
rect 21501 4766 21535 4782
rect 21679 5038 21713 5054
rect 21679 4766 21713 4782
rect 21857 5038 21971 5088
rect 21891 4782 21971 5038
rect 21857 4732 21971 4782
rect 18929 4698 19089 4732
rect 19141 4698 19157 4732
rect 19251 4698 19267 4732
rect 19319 4698 19335 4732
rect 19429 4698 19445 4732
rect 19497 4698 19513 4732
rect 19607 4698 19623 4732
rect 19675 4698 19691 4732
rect 19785 4698 19801 4732
rect 19853 4698 19869 4732
rect 19963 4698 19979 4732
rect 20031 4698 20047 4732
rect 20141 4698 20157 4732
rect 20209 4698 20225 4732
rect 20319 4698 20335 4732
rect 20387 4698 20403 4732
rect 20497 4698 20513 4732
rect 20565 4698 20581 4732
rect 20675 4698 20691 4732
rect 20743 4698 20759 4732
rect 20853 4698 20869 4732
rect 20921 4698 20937 4732
rect 21031 4698 21047 4732
rect 21099 4698 21115 4732
rect 21209 4698 21225 4732
rect 21277 4698 21293 4732
rect 21387 4698 21403 4732
rect 21455 4698 21471 4732
rect 21565 4698 21581 4732
rect 21633 4698 21649 4732
rect 21743 4698 21759 4732
rect 21811 4698 21971 4732
rect 18929 4624 19016 4698
rect 21891 4624 21971 4698
rect 18929 4590 19089 4624
rect 19141 4590 19157 4624
rect 19251 4590 19267 4624
rect 19319 4590 19335 4624
rect 19429 4590 19445 4624
rect 19497 4590 19513 4624
rect 19607 4590 19623 4624
rect 19675 4590 19691 4624
rect 19785 4590 19801 4624
rect 19853 4590 19869 4624
rect 19963 4590 19979 4624
rect 20031 4590 20047 4624
rect 20141 4590 20157 4624
rect 20209 4590 20225 4624
rect 20319 4590 20335 4624
rect 20387 4590 20403 4624
rect 20497 4590 20513 4624
rect 20565 4590 20581 4624
rect 20675 4590 20691 4624
rect 20743 4590 20759 4624
rect 20853 4590 20869 4624
rect 20921 4590 20937 4624
rect 21031 4590 21047 4624
rect 21099 4590 21115 4624
rect 21209 4590 21225 4624
rect 21277 4590 21293 4624
rect 21387 4590 21403 4624
rect 21455 4590 21471 4624
rect 21565 4590 21581 4624
rect 21633 4590 21649 4624
rect 21743 4590 21759 4624
rect 21811 4590 21971 4624
rect 18929 4540 19043 4590
rect 18929 4284 19009 4540
rect 18929 4234 19043 4284
rect 19187 4540 19221 4556
rect 19187 4268 19221 4284
rect 19365 4540 19399 4556
rect 19365 4268 19399 4284
rect 19543 4540 19577 4556
rect 19543 4268 19577 4284
rect 19721 4540 19755 4556
rect 19721 4268 19755 4284
rect 19899 4540 19933 4556
rect 19899 4268 19933 4284
rect 20077 4540 20111 4556
rect 20077 4268 20111 4284
rect 20255 4540 20289 4556
rect 20255 4268 20289 4284
rect 20433 4540 20467 4556
rect 20433 4268 20467 4284
rect 20611 4540 20645 4556
rect 20611 4268 20645 4284
rect 20789 4540 20823 4556
rect 20789 4268 20823 4284
rect 20967 4540 21001 4556
rect 20967 4268 21001 4284
rect 21145 4540 21179 4556
rect 21145 4268 21179 4284
rect 21323 4540 21357 4556
rect 21323 4268 21357 4284
rect 21501 4540 21535 4556
rect 21501 4268 21535 4284
rect 21679 4540 21713 4556
rect 21679 4268 21713 4284
rect 21857 4540 21971 4590
rect 21891 4284 21971 4540
rect 21857 4234 21971 4284
rect 18929 4200 19089 4234
rect 19141 4200 19157 4234
rect 19251 4200 19267 4234
rect 19319 4200 19335 4234
rect 19429 4200 19445 4234
rect 19497 4200 19513 4234
rect 19607 4200 19623 4234
rect 19675 4200 19691 4234
rect 19785 4200 19801 4234
rect 19853 4200 19869 4234
rect 19963 4200 19979 4234
rect 20031 4200 20047 4234
rect 20141 4200 20157 4234
rect 20209 4200 20225 4234
rect 20319 4200 20335 4234
rect 20387 4200 20403 4234
rect 20497 4200 20513 4234
rect 20565 4200 20581 4234
rect 20675 4200 20691 4234
rect 20743 4200 20759 4234
rect 20853 4200 20869 4234
rect 20921 4200 20937 4234
rect 21031 4200 21047 4234
rect 21099 4200 21115 4234
rect 21209 4200 21225 4234
rect 21277 4200 21293 4234
rect 21387 4200 21403 4234
rect 21455 4200 21471 4234
rect 21565 4200 21581 4234
rect 21633 4200 21649 4234
rect 21743 4200 21759 4234
rect 21811 4200 21971 4234
rect 18929 4126 19016 4200
rect 21891 4126 21971 4200
rect 18929 4092 19089 4126
rect 19141 4092 19157 4126
rect 19251 4092 19267 4126
rect 19319 4092 19335 4126
rect 19429 4092 19445 4126
rect 19497 4092 19513 4126
rect 19607 4092 19623 4126
rect 19675 4092 19691 4126
rect 19785 4092 19801 4126
rect 19853 4092 19869 4126
rect 19963 4092 19979 4126
rect 20031 4092 20047 4126
rect 20141 4092 20157 4126
rect 20209 4092 20225 4126
rect 20319 4092 20335 4126
rect 20387 4092 20403 4126
rect 20497 4092 20513 4126
rect 20565 4092 20581 4126
rect 20675 4092 20691 4126
rect 20743 4092 20759 4126
rect 20853 4092 20869 4126
rect 20921 4092 20937 4126
rect 21031 4092 21047 4126
rect 21099 4092 21115 4126
rect 21209 4092 21225 4126
rect 21277 4092 21293 4126
rect 21387 4092 21403 4126
rect 21455 4092 21471 4126
rect 21565 4092 21581 4126
rect 21633 4092 21649 4126
rect 21743 4092 21759 4126
rect 21811 4092 21971 4126
rect 18929 4042 19043 4092
rect 18929 3786 19009 4042
rect 18929 3736 19043 3786
rect 19187 4042 19221 4058
rect 19187 3770 19221 3786
rect 19365 4042 19399 4058
rect 19365 3770 19399 3786
rect 19543 4042 19577 4058
rect 19543 3770 19577 3786
rect 19721 4042 19755 4058
rect 19721 3770 19755 3786
rect 19899 4042 19933 4058
rect 19899 3770 19933 3786
rect 20077 4042 20111 4058
rect 20077 3770 20111 3786
rect 20255 4042 20289 4058
rect 20255 3770 20289 3786
rect 20433 4042 20467 4058
rect 20433 3770 20467 3786
rect 20611 4042 20645 4058
rect 20611 3770 20645 3786
rect 20789 4042 20823 4058
rect 20789 3770 20823 3786
rect 20967 4042 21001 4058
rect 20967 3770 21001 3786
rect 21145 4042 21179 4058
rect 21145 3770 21179 3786
rect 21323 4042 21357 4058
rect 21323 3770 21357 3786
rect 21501 4042 21535 4058
rect 21501 3770 21535 3786
rect 21679 4042 21713 4058
rect 21679 3770 21713 3786
rect 21857 4042 21971 4092
rect 21891 3786 21971 4042
rect 21857 3736 21971 3786
rect 18929 3702 19089 3736
rect 19141 3702 19157 3736
rect 19251 3702 19267 3736
rect 19319 3702 19335 3736
rect 19429 3702 19445 3736
rect 19497 3702 19513 3736
rect 19607 3702 19623 3736
rect 19675 3702 19691 3736
rect 19785 3702 19801 3736
rect 19853 3702 19869 3736
rect 19963 3702 19979 3736
rect 20031 3702 20047 3736
rect 20141 3702 20157 3736
rect 20209 3702 20225 3736
rect 20319 3702 20335 3736
rect 20387 3702 20403 3736
rect 20497 3702 20513 3736
rect 20565 3702 20581 3736
rect 20675 3702 20691 3736
rect 20743 3702 20759 3736
rect 20853 3702 20869 3736
rect 20921 3702 20937 3736
rect 21031 3702 21047 3736
rect 21099 3702 21115 3736
rect 21209 3702 21225 3736
rect 21277 3702 21293 3736
rect 21387 3702 21403 3736
rect 21455 3702 21471 3736
rect 21565 3702 21581 3736
rect 21633 3702 21649 3736
rect 21743 3702 21759 3736
rect 21811 3702 21971 3736
rect 18929 3628 19016 3702
rect 21891 3628 21971 3702
rect 18929 3594 19089 3628
rect 19141 3594 19157 3628
rect 19251 3594 19267 3628
rect 19319 3594 19335 3628
rect 19429 3594 19445 3628
rect 19497 3594 19513 3628
rect 19607 3594 19623 3628
rect 19675 3594 19691 3628
rect 19785 3594 19801 3628
rect 19853 3594 19869 3628
rect 19963 3594 19979 3628
rect 20031 3594 20047 3628
rect 20141 3594 20157 3628
rect 20209 3594 20225 3628
rect 20319 3594 20335 3628
rect 20387 3594 20403 3628
rect 20497 3594 20513 3628
rect 20565 3594 20581 3628
rect 20675 3594 20691 3628
rect 20743 3594 20759 3628
rect 20853 3594 20869 3628
rect 20921 3594 20937 3628
rect 21031 3594 21047 3628
rect 21099 3594 21115 3628
rect 21209 3594 21225 3628
rect 21277 3594 21293 3628
rect 21387 3594 21403 3628
rect 21455 3594 21471 3628
rect 21565 3594 21581 3628
rect 21633 3594 21649 3628
rect 21743 3594 21759 3628
rect 21811 3594 21971 3628
rect 18929 3544 19043 3594
rect 18929 3288 19009 3544
rect 18929 3238 19043 3288
rect 19187 3544 19221 3560
rect 19187 3272 19221 3288
rect 19365 3544 19399 3560
rect 19365 3272 19399 3288
rect 19543 3544 19577 3560
rect 19543 3272 19577 3288
rect 19721 3544 19755 3560
rect 19721 3272 19755 3288
rect 19899 3544 19933 3560
rect 19899 3272 19933 3288
rect 20077 3544 20111 3560
rect 20077 3272 20111 3288
rect 20255 3544 20289 3560
rect 20255 3272 20289 3288
rect 20433 3544 20467 3560
rect 20433 3272 20467 3288
rect 20611 3544 20645 3560
rect 20611 3272 20645 3288
rect 20789 3544 20823 3560
rect 20789 3272 20823 3288
rect 20967 3544 21001 3560
rect 20967 3272 21001 3288
rect 21145 3544 21179 3560
rect 21145 3272 21179 3288
rect 21323 3544 21357 3560
rect 21323 3272 21357 3288
rect 21501 3544 21535 3560
rect 21501 3272 21535 3288
rect 21679 3544 21713 3560
rect 21679 3272 21713 3288
rect 21857 3544 21971 3594
rect 21891 3288 21971 3544
rect 21857 3238 21971 3288
rect 18929 3204 19089 3238
rect 19141 3204 19157 3238
rect 19251 3204 19267 3238
rect 19319 3204 19335 3238
rect 19429 3204 19445 3238
rect 19497 3204 19513 3238
rect 19607 3204 19623 3238
rect 19675 3204 19691 3238
rect 19785 3204 19801 3238
rect 19853 3204 19869 3238
rect 19963 3204 19979 3238
rect 20031 3204 20047 3238
rect 20141 3204 20157 3238
rect 20209 3204 20225 3238
rect 20319 3204 20335 3238
rect 20387 3204 20403 3238
rect 20497 3204 20513 3238
rect 20565 3204 20581 3238
rect 20675 3204 20691 3238
rect 20743 3204 20759 3238
rect 20853 3204 20869 3238
rect 20921 3204 20937 3238
rect 21031 3204 21047 3238
rect 21099 3204 21115 3238
rect 21209 3204 21225 3238
rect 21277 3204 21293 3238
rect 21387 3204 21403 3238
rect 21455 3204 21471 3238
rect 21565 3204 21581 3238
rect 21633 3204 21649 3238
rect 21743 3204 21759 3238
rect 21811 3204 21971 3238
rect 18929 3198 19016 3204
rect 18888 3136 19016 3198
rect 21891 3198 21971 3204
rect 22005 3198 22019 5128
rect 21891 3136 22019 3198
rect 18888 3102 18991 3136
rect 21909 3102 22019 3136
rect 18888 149 19016 3102
rect 19254 2716 19382 2723
rect 21398 2716 21526 2720
rect 19253 2702 19349 2716
rect 19196 2682 19349 2702
rect 21377 2682 21526 2716
rect 19196 2620 19382 2682
rect 19196 690 19253 2620
rect 19287 2614 19382 2620
rect 21332 2620 21526 2682
rect 21332 2614 21439 2620
rect 19287 2580 19447 2614
rect 19499 2580 19515 2614
rect 19609 2580 19625 2614
rect 19677 2580 19693 2614
rect 19787 2580 19803 2614
rect 19855 2580 19871 2614
rect 19965 2580 19981 2614
rect 20033 2580 20049 2614
rect 20143 2580 20159 2614
rect 20211 2580 20227 2614
rect 20321 2580 20337 2614
rect 20389 2580 20405 2614
rect 20499 2580 20515 2614
rect 20567 2580 20583 2614
rect 20677 2580 20693 2614
rect 20745 2580 20761 2614
rect 20855 2580 20871 2614
rect 20923 2580 20939 2614
rect 21033 2580 21049 2614
rect 21101 2580 21117 2614
rect 21211 2580 21227 2614
rect 21279 2580 21439 2614
rect 19287 2530 19401 2580
rect 19287 2274 19367 2530
rect 19287 2224 19401 2274
rect 19545 2530 19579 2546
rect 19545 2258 19579 2274
rect 19723 2530 19757 2546
rect 19723 2258 19757 2274
rect 19901 2530 19935 2546
rect 19901 2258 19935 2274
rect 20079 2530 20113 2546
rect 20079 2258 20113 2274
rect 20257 2530 20291 2546
rect 20257 2258 20291 2274
rect 20435 2530 20469 2546
rect 20435 2258 20469 2274
rect 20613 2530 20647 2546
rect 20613 2258 20647 2274
rect 20791 2530 20825 2546
rect 20791 2258 20825 2274
rect 20969 2530 21003 2546
rect 20969 2258 21003 2274
rect 21147 2530 21181 2546
rect 21147 2258 21181 2274
rect 21325 2530 21439 2580
rect 21359 2274 21439 2530
rect 21325 2224 21439 2274
rect 19287 2190 19447 2224
rect 19499 2190 19515 2224
rect 19609 2190 19625 2224
rect 19677 2190 19693 2224
rect 19787 2190 19803 2224
rect 19855 2190 19871 2224
rect 19965 2190 19981 2224
rect 20033 2190 20049 2224
rect 20143 2190 20159 2224
rect 20211 2190 20227 2224
rect 20321 2190 20337 2224
rect 20389 2190 20405 2224
rect 20499 2190 20515 2224
rect 20567 2190 20583 2224
rect 20677 2190 20693 2224
rect 20745 2190 20761 2224
rect 20855 2190 20871 2224
rect 20923 2190 20939 2224
rect 21033 2190 21049 2224
rect 21101 2190 21117 2224
rect 21211 2190 21227 2224
rect 21279 2190 21439 2224
rect 19287 2116 19382 2190
rect 21332 2116 21439 2190
rect 19287 2082 19447 2116
rect 19499 2082 19515 2116
rect 19609 2082 19625 2116
rect 19677 2082 19693 2116
rect 19787 2082 19803 2116
rect 19855 2082 19871 2116
rect 19965 2082 19981 2116
rect 20033 2082 20049 2116
rect 20143 2082 20159 2116
rect 20211 2082 20227 2116
rect 20321 2082 20337 2116
rect 20389 2082 20405 2116
rect 20499 2082 20515 2116
rect 20567 2082 20583 2116
rect 20677 2082 20693 2116
rect 20745 2082 20761 2116
rect 20855 2082 20871 2116
rect 20923 2082 20939 2116
rect 21033 2082 21049 2116
rect 21101 2082 21117 2116
rect 21211 2082 21227 2116
rect 21279 2082 21439 2116
rect 19287 2032 19401 2082
rect 19287 1776 19367 2032
rect 19287 1726 19401 1776
rect 19545 2032 19579 2048
rect 19545 1760 19579 1776
rect 19723 2032 19757 2048
rect 19723 1760 19757 1776
rect 19901 2032 19935 2048
rect 19901 1760 19935 1776
rect 20079 2032 20113 2048
rect 20079 1760 20113 1776
rect 20257 2032 20291 2048
rect 20257 1760 20291 1776
rect 20435 2032 20469 2048
rect 20435 1760 20469 1776
rect 20613 2032 20647 2048
rect 20613 1760 20647 1776
rect 20791 2032 20825 2048
rect 20791 1760 20825 1776
rect 20969 2032 21003 2048
rect 20969 1760 21003 1776
rect 21147 2032 21181 2048
rect 21147 1760 21181 1776
rect 21325 2032 21439 2082
rect 21359 1776 21439 2032
rect 21325 1726 21439 1776
rect 19287 1692 19447 1726
rect 19499 1692 19515 1726
rect 19609 1692 19625 1726
rect 19677 1692 19693 1726
rect 19787 1692 19803 1726
rect 19855 1692 19871 1726
rect 19965 1692 19981 1726
rect 20033 1692 20049 1726
rect 20143 1692 20159 1726
rect 20211 1692 20227 1726
rect 20321 1692 20337 1726
rect 20389 1692 20405 1726
rect 20499 1692 20515 1726
rect 20567 1692 20583 1726
rect 20677 1692 20693 1726
rect 20745 1692 20761 1726
rect 20855 1692 20871 1726
rect 20923 1692 20939 1726
rect 21033 1692 21049 1726
rect 21101 1692 21117 1726
rect 21211 1692 21227 1726
rect 21279 1692 21439 1726
rect 19287 1618 19382 1692
rect 21332 1618 21439 1692
rect 19287 1584 19447 1618
rect 19499 1584 19515 1618
rect 19609 1584 19625 1618
rect 19677 1584 19693 1618
rect 19787 1584 19803 1618
rect 19855 1584 19871 1618
rect 19965 1584 19981 1618
rect 20033 1584 20049 1618
rect 20143 1584 20159 1618
rect 20211 1584 20227 1618
rect 20321 1584 20337 1618
rect 20389 1584 20405 1618
rect 20499 1584 20515 1618
rect 20567 1584 20583 1618
rect 20677 1584 20693 1618
rect 20745 1584 20761 1618
rect 20855 1584 20871 1618
rect 20923 1584 20939 1618
rect 21033 1584 21049 1618
rect 21101 1584 21117 1618
rect 21211 1584 21227 1618
rect 21279 1584 21439 1618
rect 19287 1534 19401 1584
rect 19287 1278 19367 1534
rect 19287 1228 19401 1278
rect 19545 1534 19579 1550
rect 19545 1262 19579 1278
rect 19723 1534 19757 1550
rect 19723 1262 19757 1278
rect 19901 1534 19935 1550
rect 19901 1262 19935 1278
rect 20079 1534 20113 1550
rect 20079 1262 20113 1278
rect 20257 1534 20291 1550
rect 20257 1262 20291 1278
rect 20435 1534 20469 1550
rect 20435 1262 20469 1278
rect 20613 1534 20647 1550
rect 20613 1262 20647 1278
rect 20791 1534 20825 1550
rect 20791 1262 20825 1278
rect 20969 1534 21003 1550
rect 20969 1262 21003 1278
rect 21147 1534 21181 1550
rect 21147 1262 21181 1278
rect 21325 1534 21439 1584
rect 21359 1278 21439 1534
rect 21325 1228 21439 1278
rect 19287 1194 19447 1228
rect 19499 1194 19515 1228
rect 19609 1194 19625 1228
rect 19677 1194 19693 1228
rect 19787 1194 19803 1228
rect 19855 1194 19871 1228
rect 19965 1194 19981 1228
rect 20033 1194 20049 1228
rect 20143 1194 20159 1228
rect 20211 1194 20227 1228
rect 20321 1194 20337 1228
rect 20389 1194 20405 1228
rect 20499 1194 20515 1228
rect 20567 1194 20583 1228
rect 20677 1194 20693 1228
rect 20745 1194 20761 1228
rect 20855 1194 20871 1228
rect 20923 1194 20939 1228
rect 21033 1194 21049 1228
rect 21101 1194 21117 1228
rect 21211 1194 21227 1228
rect 21279 1194 21439 1228
rect 19287 1120 19382 1194
rect 21332 1120 21439 1194
rect 19287 1086 19447 1120
rect 19499 1086 19515 1120
rect 19609 1086 19625 1120
rect 19677 1086 19693 1120
rect 19787 1086 19803 1120
rect 19855 1086 19871 1120
rect 19965 1086 19981 1120
rect 20033 1086 20049 1120
rect 20143 1086 20159 1120
rect 20211 1086 20227 1120
rect 20321 1086 20337 1120
rect 20389 1086 20405 1120
rect 20499 1086 20515 1120
rect 20567 1086 20583 1120
rect 20677 1086 20693 1120
rect 20745 1086 20761 1120
rect 20855 1086 20871 1120
rect 20923 1086 20939 1120
rect 21033 1086 21049 1120
rect 21101 1086 21117 1120
rect 21211 1086 21227 1120
rect 21279 1086 21439 1120
rect 19287 1036 19401 1086
rect 19287 780 19367 1036
rect 19287 730 19401 780
rect 19545 1036 19579 1052
rect 19545 764 19579 780
rect 19723 1036 19757 1052
rect 19723 764 19757 780
rect 19901 1036 19935 1052
rect 19901 764 19935 780
rect 20079 1036 20113 1052
rect 20079 764 20113 780
rect 20257 1036 20291 1052
rect 20257 764 20291 780
rect 20435 1036 20469 1052
rect 20435 764 20469 780
rect 20613 1036 20647 1052
rect 20613 764 20647 780
rect 20791 1036 20825 1052
rect 20791 764 20825 780
rect 20969 1036 21003 1052
rect 20969 764 21003 780
rect 21147 1036 21181 1052
rect 21147 764 21181 780
rect 21325 1036 21439 1086
rect 21359 780 21439 1036
rect 21325 730 21439 780
rect 19287 696 19447 730
rect 19499 696 19515 730
rect 19609 696 19625 730
rect 19677 696 19693 730
rect 19787 696 19803 730
rect 19855 696 19871 730
rect 19965 696 19981 730
rect 20033 696 20049 730
rect 20143 696 20159 730
rect 20211 696 20227 730
rect 20321 696 20337 730
rect 20389 696 20405 730
rect 20499 696 20515 730
rect 20567 696 20583 730
rect 20677 696 20693 730
rect 20745 696 20761 730
rect 20855 696 20871 730
rect 20923 696 20939 730
rect 21033 696 21049 730
rect 21101 696 21117 730
rect 21211 696 21227 730
rect 21279 696 21439 730
rect 19287 690 19382 696
rect 19196 628 19382 690
rect 21332 690 21439 696
rect 21473 690 21526 2620
rect 21332 628 21526 690
rect 19196 594 19349 628
rect 21377 594 21526 628
rect 19196 149 19382 594
rect 19855 149 19983 594
rect 20566 149 20694 594
rect 21332 149 21526 594
rect 21891 280 22019 3102
rect 23491 280 23747 8325
rect 21891 149 23747 280
rect 13367 129 23747 149
rect 13367 113 14118 129
rect -61 71 14118 113
rect -61 22 304 71
rect 13205 70 14118 71
rect 14211 127 23747 129
rect 14211 123 16542 127
rect 14211 70 15279 123
rect 15372 70 16542 123
rect 16635 122 23747 127
rect 16635 70 17969 122
rect 18062 70 23747 122
rect 13205 22 13476 70
rect -61 21 13476 22
rect 18366 24 23747 70
rect 18366 21 22071 24
rect -61 18 195 21
<< viali >>
rect 7303 18801 7337 18835
rect 8262 18801 8263 18835
rect 8263 18801 8296 18835
rect 7303 18493 7337 18741
rect 7399 18493 7433 18741
rect 7495 18493 7529 18741
rect 7591 18493 7625 18741
rect 7687 18493 7721 18741
rect 7783 18493 7817 18741
rect 7879 18493 7913 18741
rect 7975 18493 8009 18741
rect 8071 18493 8105 18741
rect 8167 18493 8201 18741
rect 8263 18493 8297 18741
rect 7303 18083 7337 18163
rect 7399 18083 7433 18163
rect 7495 18083 7529 18163
rect 7591 18083 7625 18163
rect 7687 18083 7721 18163
rect 7783 18083 7817 18163
rect 7879 18083 7913 18163
rect 7975 18083 8009 18163
rect 8071 18083 8105 18163
rect 8167 18083 8201 18163
rect 8263 18083 8297 18163
rect 7303 17990 7337 18023
rect 8264 17990 8297 18024
rect 8297 17990 8298 18024
rect 7303 17989 7337 17990
rect 7303 17035 7337 17036
rect 7303 17002 7337 17035
rect 8263 17001 8297 17035
rect 7303 16693 7337 16941
rect 7399 16693 7433 16941
rect 7495 16693 7529 16941
rect 7591 16693 7625 16941
rect 7687 16693 7721 16941
rect 7783 16693 7817 16941
rect 7879 16693 7913 16941
rect 7975 16693 8009 16941
rect 8071 16693 8105 16941
rect 8167 16693 8201 16941
rect 8263 16693 8297 16941
rect 7303 16283 7337 16363
rect 7399 16283 7433 16363
rect 7495 16283 7529 16363
rect 7591 16283 7625 16363
rect 7687 16283 7721 16363
rect 7783 16283 7817 16363
rect 7879 16283 7913 16363
rect 7975 16283 8009 16363
rect 8071 16283 8105 16363
rect 8167 16283 8201 16363
rect 8263 16283 8297 16363
rect 7304 16190 7337 16223
rect 7337 16190 7338 16223
rect 8261 16190 8263 16223
rect 8263 16190 8295 16223
rect 7304 16189 7338 16190
rect 8261 16189 8295 16190
rect 7301 15201 7303 15235
rect 7303 15201 7335 15235
rect 8265 15201 8297 15235
rect 8297 15201 8299 15235
rect 7303 14893 7337 15141
rect 7399 14893 7433 15141
rect 7495 14893 7529 15141
rect 7591 14893 7625 15141
rect 7687 14893 7721 15141
rect 7783 14893 7817 15141
rect 7879 14893 7913 15141
rect 7975 14893 8009 15141
rect 8071 14893 8105 15141
rect 8167 14893 8201 15141
rect 8263 14893 8297 15141
rect 7303 14483 7337 14563
rect 7399 14483 7433 14563
rect 7495 14483 7529 14563
rect 7591 14483 7625 14563
rect 7687 14483 7721 14563
rect 7783 14483 7817 14563
rect 7879 14483 7913 14563
rect 7975 14483 8009 14563
rect 8071 14483 8105 14563
rect 8167 14483 8201 14563
rect 8263 14483 8297 14563
rect 7304 14390 7337 14423
rect 7337 14390 7338 14423
rect 8263 14390 8297 14424
rect 7304 14389 7338 14390
rect 7304 13435 7338 13436
rect 8262 13435 8296 13436
rect 7304 13402 7337 13435
rect 7337 13402 7338 13435
rect 8262 13402 8263 13435
rect 8263 13402 8296 13435
rect 7303 13093 7337 13341
rect 7399 13093 7433 13341
rect 7495 13093 7529 13341
rect 7591 13093 7625 13341
rect 7687 13093 7721 13341
rect 7783 13093 7817 13341
rect 7879 13093 7913 13341
rect 7975 13093 8009 13341
rect 8071 13093 8105 13341
rect 8167 13093 8201 13341
rect 8263 13093 8297 13341
rect 7303 12683 7337 12763
rect 7399 12683 7433 12763
rect 7495 12683 7529 12763
rect 7591 12683 7625 12763
rect 7687 12683 7721 12763
rect 7783 12683 7817 12763
rect 7879 12683 7913 12763
rect 7975 12683 8009 12763
rect 8071 12683 8105 12763
rect 8167 12683 8201 12763
rect 8263 12683 8297 12763
rect 7301 12590 7303 12623
rect 7303 12590 7335 12623
rect 8264 12590 8297 12623
rect 8297 12590 8298 12623
rect 7301 12589 7335 12590
rect 8264 12589 8298 12590
rect 8262 11635 8296 11636
rect 7301 11601 7303 11635
rect 7303 11601 7335 11635
rect 8262 11602 8263 11635
rect 8263 11602 8296 11635
rect 7303 11293 7337 11541
rect 7399 11293 7433 11541
rect 7495 11293 7529 11541
rect 7591 11293 7625 11541
rect 7687 11293 7721 11541
rect 7783 11293 7817 11541
rect 7879 11293 7913 11541
rect 7975 11293 8009 11541
rect 8071 11293 8105 11541
rect 8167 11293 8201 11541
rect 8263 11293 8297 11541
rect 7303 10883 7337 10963
rect 7399 10883 7433 10963
rect 7495 10883 7529 10963
rect 7591 10883 7625 10963
rect 7687 10883 7721 10963
rect 7783 10883 7817 10963
rect 7879 10883 7913 10963
rect 7975 10883 8009 10963
rect 8071 10883 8105 10963
rect 8167 10883 8201 10963
rect 8263 10883 8297 10963
rect 7300 10790 7303 10823
rect 7303 10790 7334 10823
rect 8262 10790 8263 10823
rect 8263 10790 8296 10823
rect 7300 10789 7334 10790
rect 8262 10789 8296 10790
rect 8262 9835 8296 9837
rect 7302 9801 7303 9834
rect 7303 9801 7336 9834
rect 8262 9803 8263 9835
rect 8263 9803 8296 9835
rect 7302 9800 7336 9801
rect 7303 9493 7337 9741
rect 7399 9493 7433 9741
rect 7495 9493 7529 9741
rect 7591 9493 7625 9741
rect 7687 9493 7721 9741
rect 7783 9493 7817 9741
rect 7879 9493 7913 9741
rect 7975 9493 8009 9741
rect 8071 9493 8105 9741
rect 8167 9493 8201 9741
rect 8263 9493 8297 9741
rect 7303 9083 7337 9163
rect 7399 9083 7433 9163
rect 7495 9083 7529 9163
rect 7591 9083 7625 9163
rect 7687 9083 7721 9163
rect 7783 9083 7817 9163
rect 7879 9083 7913 9163
rect 7975 9083 8009 9163
rect 8071 9083 8105 9163
rect 8167 9083 8201 9163
rect 8263 9083 8297 9163
rect 7303 9024 7337 9026
rect 8260 9024 8294 9026
rect 7303 8992 7337 9024
rect 8260 8992 8263 9024
rect 8263 8992 8294 9024
rect 8715 8761 8971 9017
rect 20224 18835 20258 18837
rect 20224 18803 20233 18835
rect 20233 18803 20258 18835
rect 21192 18801 21193 18835
rect 21193 18801 21226 18835
rect 20233 18493 20267 18741
rect 20329 18493 20363 18741
rect 20425 18493 20459 18741
rect 20521 18493 20555 18741
rect 20617 18493 20651 18741
rect 20713 18493 20747 18741
rect 20809 18493 20843 18741
rect 20905 18493 20939 18741
rect 21001 18493 21035 18741
rect 21097 18493 21131 18741
rect 21193 18493 21227 18741
rect 20233 18083 20267 18163
rect 20329 18083 20363 18163
rect 20425 18083 20459 18163
rect 20521 18083 20555 18163
rect 20617 18083 20651 18163
rect 20713 18083 20747 18163
rect 20809 18083 20843 18163
rect 20905 18083 20939 18163
rect 21001 18083 21035 18163
rect 21097 18083 21131 18163
rect 21193 18083 21227 18163
rect 21196 18024 21230 18026
rect 20233 17990 20267 18024
rect 21196 17992 21227 18024
rect 21227 17992 21230 18024
rect 20229 17035 20263 17039
rect 20229 17005 20233 17035
rect 20233 17005 20263 17035
rect 21194 17001 21227 17035
rect 21227 17001 21228 17035
rect 20233 16693 20267 16941
rect 20329 16693 20363 16941
rect 20425 16693 20459 16941
rect 20521 16693 20555 16941
rect 20617 16693 20651 16941
rect 20713 16693 20747 16941
rect 20809 16693 20843 16941
rect 20905 16693 20939 16941
rect 21001 16693 21035 16941
rect 21097 16693 21131 16941
rect 21193 16693 21227 16941
rect 20233 16283 20267 16363
rect 20329 16283 20363 16363
rect 20425 16283 20459 16363
rect 20521 16283 20555 16363
rect 20617 16283 20651 16363
rect 20713 16283 20747 16363
rect 20809 16283 20843 16363
rect 20905 16283 20939 16363
rect 21001 16283 21035 16363
rect 21097 16283 21131 16363
rect 21193 16283 21227 16363
rect 20229 16224 20263 16226
rect 21194 16224 21228 16228
rect 20229 16192 20233 16224
rect 20233 16192 20263 16224
rect 21194 16194 21227 16224
rect 21227 16194 21228 16224
rect 20235 15201 20267 15235
rect 20267 15201 20269 15235
rect 21196 15201 21227 15235
rect 21227 15201 21230 15235
rect 20233 14893 20267 15141
rect 20329 14893 20363 15141
rect 20425 14893 20459 15141
rect 20521 14893 20555 15141
rect 20617 14893 20651 15141
rect 20713 14893 20747 15141
rect 20809 14893 20843 15141
rect 20905 14893 20939 15141
rect 21001 14893 21035 15141
rect 21097 14893 21131 15141
rect 21193 14893 21227 15141
rect 20233 14483 20267 14563
rect 20329 14483 20363 14563
rect 20425 14483 20459 14563
rect 20521 14483 20555 14563
rect 20617 14483 20651 14563
rect 20713 14483 20747 14563
rect 20809 14483 20843 14563
rect 20905 14483 20939 14563
rect 21001 14483 21035 14563
rect 21097 14483 21131 14563
rect 21193 14483 21227 14563
rect 21200 14424 21234 14426
rect 20231 14390 20233 14422
rect 20233 14390 20265 14422
rect 21200 14392 21227 14424
rect 21227 14392 21234 14424
rect 20231 14388 20265 14390
rect 20231 13435 20265 13439
rect 21192 13435 21226 13439
rect 20231 13405 20233 13435
rect 20233 13405 20265 13435
rect 21192 13405 21193 13435
rect 21193 13405 21226 13435
rect 20233 13093 20267 13341
rect 20329 13093 20363 13341
rect 20425 13093 20459 13341
rect 20521 13093 20555 13341
rect 20617 13093 20651 13341
rect 20713 13093 20747 13341
rect 20809 13093 20843 13341
rect 20905 13093 20939 13341
rect 21001 13093 21035 13341
rect 21097 13093 21131 13341
rect 21193 13093 21227 13341
rect 20233 12683 20267 12763
rect 20329 12683 20363 12763
rect 20425 12683 20459 12763
rect 20521 12683 20555 12763
rect 20617 12683 20651 12763
rect 20713 12683 20747 12763
rect 20809 12683 20843 12763
rect 20905 12683 20939 12763
rect 21001 12683 21035 12763
rect 21097 12683 21131 12763
rect 21193 12683 21227 12763
rect 20229 12590 20233 12624
rect 20233 12590 20263 12624
rect 21196 12590 21227 12620
rect 21227 12590 21230 12620
rect 21196 12586 21230 12590
rect 20231 11635 20265 11639
rect 20231 11605 20233 11635
rect 20233 11605 20265 11635
rect 21196 11601 21227 11633
rect 21227 11601 21230 11633
rect 21196 11599 21230 11601
rect 20233 11293 20267 11541
rect 20329 11293 20363 11541
rect 20425 11293 20459 11541
rect 20521 11293 20555 11541
rect 20617 11293 20651 11541
rect 20713 11293 20747 11541
rect 20809 11293 20843 11541
rect 20905 11293 20939 11541
rect 21001 11293 21035 11541
rect 21097 11293 21131 11541
rect 21193 11293 21227 11541
rect 20233 10883 20267 10963
rect 20329 10883 20363 10963
rect 20425 10883 20459 10963
rect 20521 10883 20555 10963
rect 20617 10883 20651 10963
rect 20713 10883 20747 10963
rect 20809 10883 20843 10963
rect 20905 10883 20939 10963
rect 21001 10883 21035 10963
rect 21097 10883 21131 10963
rect 21193 10883 21227 10963
rect 20231 10790 20233 10819
rect 20233 10790 20265 10819
rect 21190 10790 21193 10824
rect 21193 10790 21224 10824
rect 20231 10785 20265 10790
rect 21194 9835 21228 9839
rect 20233 9801 20267 9835
rect 21194 9805 21227 9835
rect 21227 9805 21228 9835
rect 20233 9493 20267 9741
rect 20329 9493 20363 9741
rect 20425 9493 20459 9741
rect 20521 9493 20555 9741
rect 20617 9493 20651 9741
rect 20713 9493 20747 9741
rect 20809 9493 20843 9741
rect 20905 9493 20939 9741
rect 21001 9493 21035 9741
rect 21097 9493 21131 9741
rect 21193 9493 21227 9741
rect 19650 8749 19906 9005
rect 20233 9083 20267 9163
rect 20329 9083 20363 9163
rect 20425 9083 20459 9163
rect 20521 9083 20555 9163
rect 20617 9083 20651 9163
rect 20713 9083 20747 9163
rect 20809 9083 20843 9163
rect 20905 9083 20939 9163
rect 21001 9083 21035 9163
rect 21097 9083 21131 9163
rect 21193 9083 21227 9163
rect 20237 8990 20267 9023
rect 20267 8990 20271 9023
rect 21196 8990 21227 9021
rect 21227 8990 21230 9021
rect 20237 8989 20271 8990
rect 21196 8987 21230 8990
rect 5555 8332 5799 8576
rect 23497 8325 23741 8569
rect 7445 6957 14299 6991
rect 14467 6957 20872 6991
rect 2524 4269 2558 4303
rect 2946 4269 2980 4303
rect 3370 4269 3404 4303
rect 4304 4269 4338 4303
rect 4726 4269 4760 4303
rect 5150 4269 5184 4303
rect 2262 4003 2296 4037
rect 2360 4185 2394 4219
rect 2474 4003 2508 4037
rect 2572 4185 2606 4219
rect 2686 4003 2720 4037
rect 2784 4185 2818 4219
rect 2898 4003 2932 4037
rect 2996 4185 3030 4219
rect 3110 4003 3144 4037
rect 3208 4185 3242 4219
rect 3322 4003 3356 4037
rect 3420 4185 3454 4219
rect 4042 4003 4076 4037
rect 4140 4185 4174 4219
rect 4254 4003 4288 4037
rect 4352 4185 4386 4219
rect 4466 4003 4500 4037
rect 4564 4185 4598 4219
rect 4678 4003 4712 4037
rect 4776 4185 4810 4219
rect 4890 4003 4924 4037
rect 4988 4185 5022 4219
rect 5102 4003 5136 4037
rect 5200 4185 5234 4219
rect 2312 3919 2346 3953
rect 2736 3919 2770 3953
rect 3158 3919 3192 3953
rect 4092 3919 4126 3953
rect 4516 3919 4550 3953
rect 4938 3919 4972 3953
rect 7814 6656 7866 6690
rect 7992 6656 8044 6690
rect 8170 6656 8222 6690
rect 8348 6656 8400 6690
rect 8526 6656 8578 6690
rect 8704 6656 8756 6690
rect 8882 6656 8934 6690
rect 9060 6656 9112 6690
rect 9238 6656 9290 6690
rect 9416 6656 9468 6690
rect 9594 6656 9646 6690
rect 9772 6656 9824 6690
rect 10500 6656 10552 6690
rect 10678 6656 10730 6690
rect 10856 6656 10908 6690
rect 11034 6656 11086 6690
rect 11212 6656 11264 6690
rect 11390 6656 11442 6690
rect 11568 6656 11620 6690
rect 11746 6656 11798 6690
rect 11924 6656 11976 6690
rect 12102 6656 12154 6690
rect 12280 6656 12332 6690
rect 12458 6656 12510 6690
rect 7734 6563 7768 6597
rect 7912 6341 7946 6375
rect 8090 6563 8124 6597
rect 8268 6341 8302 6375
rect 8446 6563 8480 6597
rect 8624 6341 8658 6375
rect 8802 6563 8836 6597
rect 8980 6341 9014 6375
rect 9158 6563 9192 6597
rect 9336 6341 9370 6375
rect 9514 6563 9548 6597
rect 9692 6341 9726 6375
rect 9870 6563 9904 6597
rect 10420 6563 10454 6597
rect 10598 6341 10632 6375
rect 10776 6563 10810 6597
rect 10954 6341 10988 6375
rect 11132 6563 11166 6597
rect 11310 6341 11344 6375
rect 11488 6563 11522 6597
rect 11666 6341 11700 6375
rect 11844 6563 11878 6597
rect 12022 6341 12056 6375
rect 12200 6563 12234 6597
rect 12378 6341 12412 6375
rect 12556 6563 12590 6597
rect 7814 6248 7866 6282
rect 7992 6248 8044 6282
rect 8170 6248 8222 6282
rect 8348 6248 8400 6282
rect 8526 6248 8578 6282
rect 8704 6248 8756 6282
rect 8882 6248 8934 6282
rect 9060 6248 9112 6282
rect 9238 6248 9290 6282
rect 9416 6248 9468 6282
rect 9594 6248 9646 6282
rect 9772 6248 9824 6282
rect 10500 6248 10552 6282
rect 10678 6248 10730 6282
rect 10856 6248 10908 6282
rect 11034 6248 11086 6282
rect 11212 6248 11264 6282
rect 11390 6248 11442 6282
rect 11568 6248 11620 6282
rect 11746 6248 11798 6282
rect 11924 6248 11976 6282
rect 12102 6248 12154 6282
rect 12280 6248 12332 6282
rect 12458 6248 12510 6282
rect 7814 6078 7866 6112
rect 7992 6078 8044 6112
rect 8170 6078 8222 6112
rect 8348 6078 8400 6112
rect 8526 6078 8578 6112
rect 8704 6078 8756 6112
rect 8882 6078 8934 6112
rect 9060 6078 9112 6112
rect 9238 6078 9290 6112
rect 9416 6078 9468 6112
rect 9594 6078 9646 6112
rect 9772 6078 9824 6112
rect 10500 6079 10552 6113
rect 10678 6079 10730 6113
rect 10856 6079 10908 6113
rect 11034 6079 11086 6113
rect 11212 6079 11264 6113
rect 11390 6079 11442 6113
rect 11568 6079 11620 6113
rect 11746 6079 11798 6113
rect 11924 6079 11976 6113
rect 12102 6079 12154 6113
rect 12280 6079 12332 6113
rect 12458 6079 12510 6113
rect 7734 5985 7768 6019
rect 7912 5763 7946 5797
rect 8090 5985 8124 6019
rect 8268 5763 8302 5797
rect 8446 5985 8480 6019
rect 8624 5763 8658 5797
rect 8802 5985 8836 6019
rect 8980 5763 9014 5797
rect 9158 5985 9192 6019
rect 9336 5763 9370 5797
rect 9514 5985 9548 6019
rect 9692 5763 9726 5797
rect 9870 5985 9904 6019
rect 10420 5986 10454 6020
rect 10598 5764 10632 5798
rect 10776 5986 10810 6020
rect 10954 5764 10988 5798
rect 11132 5986 11166 6020
rect 11310 5764 11344 5798
rect 11488 5986 11522 6020
rect 11666 5764 11700 5798
rect 11844 5986 11878 6020
rect 12022 5764 12056 5798
rect 12200 5986 12234 6020
rect 12378 5764 12412 5798
rect 12556 5986 12590 6020
rect 7814 5670 7866 5704
rect 7992 5670 8044 5704
rect 8170 5670 8222 5704
rect 8348 5670 8400 5704
rect 8526 5670 8578 5704
rect 8704 5670 8756 5704
rect 8882 5670 8934 5704
rect 9060 5670 9112 5704
rect 9238 5670 9290 5704
rect 9416 5670 9468 5704
rect 9594 5670 9646 5704
rect 9772 5670 9824 5704
rect 10500 5671 10552 5705
rect 10678 5671 10730 5705
rect 10856 5671 10908 5705
rect 11034 5671 11086 5705
rect 11212 5671 11264 5705
rect 11390 5671 11442 5705
rect 11568 5671 11620 5705
rect 11746 5671 11798 5705
rect 11924 5671 11976 5705
rect 12102 5671 12154 5705
rect 12280 5671 12332 5705
rect 12458 5671 12510 5705
rect 14954 6725 15006 6759
rect 15132 6725 15184 6759
rect 15310 6725 15362 6759
rect 15488 6725 15540 6759
rect 15666 6725 15718 6759
rect 15844 6725 15896 6759
rect 14874 6410 14908 6666
rect 15052 6410 15086 6666
rect 15230 6410 15264 6666
rect 15408 6410 15442 6666
rect 15586 6410 15620 6666
rect 15764 6410 15798 6666
rect 15942 6410 15976 6666
rect 14954 6317 15006 6351
rect 15132 6317 15184 6351
rect 15310 6317 15362 6351
rect 15488 6317 15540 6351
rect 15666 6317 15718 6351
rect 15844 6317 15896 6351
rect 14955 5958 15007 5992
rect 15133 5958 15185 5992
rect 15311 5958 15363 5992
rect 15489 5958 15541 5992
rect 15667 5958 15719 5992
rect 15845 5958 15897 5992
rect 14875 5643 14909 5899
rect 15053 5643 15087 5899
rect 15231 5643 15265 5899
rect 15409 5643 15443 5899
rect 15587 5643 15621 5899
rect 15765 5643 15799 5899
rect 15943 5643 15977 5899
rect 14955 5550 15007 5584
rect 15133 5550 15185 5584
rect 15311 5550 15363 5584
rect 15489 5550 15541 5584
rect 15667 5550 15719 5584
rect 15845 5550 15897 5584
rect 17154 6725 17206 6759
rect 17332 6725 17384 6759
rect 17510 6725 17562 6759
rect 17688 6725 17740 6759
rect 17866 6725 17918 6759
rect 18044 6725 18096 6759
rect 17074 6410 17108 6666
rect 17252 6410 17286 6666
rect 17430 6410 17464 6666
rect 17608 6410 17642 6666
rect 17786 6410 17820 6666
rect 17964 6410 17998 6666
rect 18142 6410 18176 6666
rect 17154 6317 17206 6351
rect 17332 6317 17384 6351
rect 17510 6317 17562 6351
rect 17688 6317 17740 6351
rect 17866 6317 17918 6351
rect 18044 6317 18096 6351
rect 17155 5958 17207 5992
rect 17333 5958 17385 5992
rect 17511 5958 17563 5992
rect 17689 5958 17741 5992
rect 17867 5958 17919 5992
rect 18045 5958 18097 5992
rect 17075 5643 17109 5899
rect 17253 5643 17287 5899
rect 17431 5643 17465 5899
rect 17609 5643 17643 5899
rect 17787 5643 17821 5899
rect 17965 5643 17999 5899
rect 18143 5643 18177 5899
rect 17155 5550 17207 5584
rect 17333 5550 17385 5584
rect 17511 5550 17563 5584
rect 17689 5550 17741 5584
rect 17867 5550 17919 5584
rect 18045 5550 18097 5584
rect 19354 6725 19406 6759
rect 19532 6725 19584 6759
rect 19710 6725 19762 6759
rect 19888 6725 19940 6759
rect 20066 6725 20118 6759
rect 20244 6725 20296 6759
rect 19274 6410 19308 6666
rect 19452 6410 19486 6666
rect 19630 6410 19664 6666
rect 19808 6410 19842 6666
rect 19986 6410 20020 6666
rect 20164 6410 20198 6666
rect 20342 6410 20376 6666
rect 19354 6317 19406 6351
rect 19532 6317 19584 6351
rect 19710 6317 19762 6351
rect 19888 6317 19940 6351
rect 20066 6317 20118 6351
rect 20244 6317 20296 6351
rect 19355 5958 19407 5992
rect 19533 5958 19585 5992
rect 19711 5958 19763 5992
rect 19889 5958 19941 5992
rect 20067 5958 20119 5992
rect 20245 5958 20297 5992
rect 19275 5643 19309 5899
rect 19453 5643 19487 5899
rect 19631 5643 19665 5899
rect 19809 5643 19843 5899
rect 19987 5643 20021 5899
rect 20165 5643 20199 5899
rect 20343 5643 20377 5899
rect 19355 5550 19407 5584
rect 19533 5550 19585 5584
rect 19711 5550 19763 5584
rect 19889 5550 19941 5584
rect 20067 5550 20119 5584
rect 20245 5550 20297 5584
rect 8170 5198 8222 5232
rect 8348 5198 8400 5232
rect 8526 5198 8578 5232
rect 8704 5198 8756 5232
rect 8882 5198 8934 5232
rect 9060 5198 9112 5232
rect 9238 5198 9290 5232
rect 9416 5198 9468 5232
rect 9594 5198 9646 5232
rect 9772 5198 9824 5232
rect 10500 5198 10552 5232
rect 10678 5198 10730 5232
rect 10856 5198 10908 5232
rect 11034 5198 11086 5232
rect 11212 5198 11264 5232
rect 11390 5198 11442 5232
rect 11568 5198 11620 5232
rect 11746 5198 11798 5232
rect 11924 5198 11976 5232
rect 12102 5198 12154 5232
rect 8090 5105 8124 5139
rect 8268 4883 8302 4917
rect 8446 5105 8480 5139
rect 8624 4883 8658 4917
rect 8802 5105 8836 5139
rect 8980 4883 9014 4917
rect 9158 5105 9192 5139
rect 9336 4883 9370 4917
rect 9514 5105 9548 5139
rect 9692 4883 9726 4917
rect 9870 5105 9904 5139
rect 10420 5105 10454 5139
rect 10598 4883 10632 4917
rect 10776 5105 10810 5139
rect 10954 4883 10988 4917
rect 11132 5105 11166 5139
rect 11310 4883 11344 4917
rect 11488 5105 11522 5139
rect 11666 4883 11700 4917
rect 11844 5105 11878 5139
rect 12022 4883 12056 4917
rect 12200 5105 12234 5139
rect 8170 4790 8222 4824
rect 8348 4790 8400 4824
rect 8526 4790 8578 4824
rect 8704 4790 8756 4824
rect 8882 4790 8934 4824
rect 9060 4790 9112 4824
rect 9238 4790 9290 4824
rect 9416 4790 9468 4824
rect 9594 4790 9646 4824
rect 9772 4790 9824 4824
rect 10500 4790 10552 4824
rect 10678 4790 10730 4824
rect 10856 4790 10908 4824
rect 11034 4790 11086 4824
rect 11212 4790 11264 4824
rect 11390 4790 11442 4824
rect 11568 4790 11620 4824
rect 11746 4790 11798 4824
rect 11924 4790 11976 4824
rect 12102 4790 12154 4824
rect 8170 4628 8222 4662
rect 8348 4628 8400 4662
rect 8526 4628 8578 4662
rect 8704 4628 8756 4662
rect 8882 4628 8934 4662
rect 9060 4628 9112 4662
rect 9238 4628 9290 4662
rect 9416 4628 9468 4662
rect 9594 4628 9646 4662
rect 9772 4628 9824 4662
rect 10500 4628 10552 4662
rect 10678 4628 10730 4662
rect 10856 4628 10908 4662
rect 11034 4628 11086 4662
rect 11212 4628 11264 4662
rect 11390 4628 11442 4662
rect 11568 4628 11620 4662
rect 11746 4628 11798 4662
rect 11924 4628 11976 4662
rect 12102 4628 12154 4662
rect 8090 4535 8124 4569
rect 8268 4313 8302 4347
rect 8446 4535 8480 4569
rect 8624 4313 8658 4347
rect 8802 4535 8836 4569
rect 8980 4313 9014 4347
rect 9158 4535 9192 4569
rect 9336 4313 9370 4347
rect 9514 4535 9548 4569
rect 9692 4313 9726 4347
rect 9870 4535 9904 4569
rect 10420 4535 10454 4569
rect 10598 4313 10632 4347
rect 10776 4535 10810 4569
rect 10954 4313 10988 4347
rect 11132 4535 11166 4569
rect 11310 4313 11344 4347
rect 11488 4535 11522 4569
rect 11666 4313 11700 4347
rect 11844 4535 11878 4569
rect 12022 4313 12056 4347
rect 12200 4535 12234 4569
rect 8170 4220 8222 4254
rect 8348 4220 8400 4254
rect 8526 4220 8578 4254
rect 8704 4220 8756 4254
rect 8882 4220 8934 4254
rect 9060 4220 9112 4254
rect 9238 4220 9290 4254
rect 9416 4220 9468 4254
rect 9594 4220 9646 4254
rect 9772 4220 9824 4254
rect 10500 4220 10552 4254
rect 10678 4220 10730 4254
rect 10856 4220 10908 4254
rect 11034 4220 11086 4254
rect 11212 4220 11264 4254
rect 11390 4220 11442 4254
rect 11568 4220 11620 4254
rect 11746 4220 11798 4254
rect 11924 4220 11976 4254
rect 12102 4220 12154 4254
rect 686 3489 738 3523
rect 864 3489 916 3523
rect 1042 3489 1094 3523
rect 1220 3489 1272 3523
rect 1398 3489 1450 3523
rect 1576 3489 1628 3523
rect 1754 3489 1806 3523
rect 1932 3489 1984 3523
rect 2110 3489 2162 3523
rect 2288 3489 2340 3523
rect 2466 3489 2518 3523
rect 2644 3489 2696 3523
rect 2822 3489 2874 3523
rect 3000 3489 3052 3523
rect 3178 3489 3230 3523
rect 3356 3489 3408 3523
rect 4086 3489 4138 3523
rect 4264 3489 4316 3523
rect 4442 3489 4494 3523
rect 4620 3489 4672 3523
rect 4798 3489 4850 3523
rect 4976 3489 5028 3523
rect 5154 3489 5206 3523
rect 5332 3489 5384 3523
rect 5510 3489 5562 3523
rect 5688 3489 5740 3523
rect 5866 3489 5918 3523
rect 6044 3489 6096 3523
rect 6222 3489 6274 3523
rect 6400 3489 6452 3523
rect 6578 3489 6630 3523
rect 6756 3489 6808 3523
rect 606 3405 640 3439
rect 784 3183 818 3217
rect 962 3405 996 3439
rect 1140 3183 1174 3217
rect 1318 3405 1352 3439
rect 1496 3183 1530 3217
rect 1674 3405 1708 3439
rect 1852 3183 1886 3217
rect 2030 3405 2064 3439
rect 2208 3183 2242 3217
rect 2386 3405 2420 3439
rect 2564 3183 2598 3217
rect 2742 3405 2776 3439
rect 2920 3183 2954 3217
rect 3098 3405 3132 3439
rect 3276 3183 3310 3217
rect 3454 3405 3488 3439
rect 4006 3405 4040 3439
rect 4184 3183 4218 3217
rect 4362 3405 4396 3439
rect 4540 3183 4574 3217
rect 4718 3405 4752 3439
rect 4896 3183 4930 3217
rect 5074 3405 5108 3439
rect 5252 3183 5286 3217
rect 5430 3405 5464 3439
rect 5608 3183 5642 3217
rect 5786 3405 5820 3439
rect 5964 3183 5998 3217
rect 6142 3405 6176 3439
rect 6320 3183 6354 3217
rect 6498 3405 6532 3439
rect 6676 3183 6710 3217
rect 6854 3405 6888 3439
rect 686 3099 738 3133
rect 864 3099 916 3133
rect 1042 3099 1094 3133
rect 1220 3099 1272 3133
rect 1398 3099 1450 3133
rect 1576 3099 1628 3133
rect 1754 3099 1806 3133
rect 1932 3099 1984 3133
rect 2110 3099 2162 3133
rect 2288 3099 2340 3133
rect 2466 3099 2518 3133
rect 2644 3099 2696 3133
rect 2822 3099 2874 3133
rect 3000 3099 3052 3133
rect 3178 3099 3230 3133
rect 3356 3099 3408 3133
rect 4086 3099 4138 3133
rect 4264 3099 4316 3133
rect 4442 3099 4494 3133
rect 4620 3099 4672 3133
rect 4798 3099 4850 3133
rect 4976 3099 5028 3133
rect 5154 3099 5206 3133
rect 5332 3099 5384 3133
rect 5510 3099 5562 3133
rect 5688 3099 5740 3133
rect 5866 3099 5918 3133
rect 6044 3099 6096 3133
rect 6222 3099 6274 3133
rect 6400 3099 6452 3133
rect 6578 3099 6630 3133
rect 6756 3099 6808 3133
rect 686 2989 738 3023
rect 864 2989 916 3023
rect 1042 2989 1094 3023
rect 1220 2989 1272 3023
rect 1398 2989 1450 3023
rect 1576 2989 1628 3023
rect 1754 2989 1806 3023
rect 1932 2989 1984 3023
rect 2110 2989 2162 3023
rect 2288 2989 2340 3023
rect 2466 2989 2518 3023
rect 2644 2989 2696 3023
rect 2822 2989 2874 3023
rect 3000 2989 3052 3023
rect 3178 2989 3230 3023
rect 3356 2989 3408 3023
rect 4086 2989 4138 3023
rect 4264 2989 4316 3023
rect 4442 2989 4494 3023
rect 4620 2989 4672 3023
rect 4798 2989 4850 3023
rect 4976 2989 5028 3023
rect 5154 2989 5206 3023
rect 5332 2989 5384 3023
rect 5510 2989 5562 3023
rect 5688 2989 5740 3023
rect 5866 2989 5918 3023
rect 6044 2989 6096 3023
rect 6222 2989 6274 3023
rect 6400 2989 6452 3023
rect 6578 2989 6630 3023
rect 6756 2989 6808 3023
rect 606 2905 640 2939
rect 784 2683 818 2717
rect 962 2905 996 2939
rect 1140 2683 1174 2717
rect 1318 2905 1352 2939
rect 1496 2683 1530 2717
rect 1674 2905 1708 2939
rect 1852 2683 1886 2717
rect 2030 2905 2064 2939
rect 2208 2683 2242 2717
rect 2386 2905 2420 2939
rect 2564 2683 2598 2717
rect 2742 2905 2776 2939
rect 2920 2683 2954 2717
rect 3098 2905 3132 2939
rect 3276 2683 3310 2717
rect 3454 2905 3488 2939
rect 4006 2905 4040 2939
rect 4184 2683 4218 2717
rect 4362 2905 4396 2939
rect 4540 2683 4574 2717
rect 4718 2905 4752 2939
rect 4896 2683 4930 2717
rect 5074 2905 5108 2939
rect 5252 2683 5286 2717
rect 5430 2905 5464 2939
rect 5608 2683 5642 2717
rect 5786 2905 5820 2939
rect 5964 2683 5998 2717
rect 6142 2905 6176 2939
rect 6320 2683 6354 2717
rect 6498 2905 6532 2939
rect 6676 2683 6710 2717
rect 6854 2905 6888 2939
rect 686 2599 738 2633
rect 864 2599 916 2633
rect 1042 2599 1094 2633
rect 1220 2599 1272 2633
rect 1398 2599 1450 2633
rect 1576 2599 1628 2633
rect 1754 2599 1806 2633
rect 1932 2599 1984 2633
rect 2110 2599 2162 2633
rect 2288 2599 2340 2633
rect 2466 2599 2518 2633
rect 2644 2599 2696 2633
rect 2822 2599 2874 2633
rect 3000 2599 3052 2633
rect 3178 2599 3230 2633
rect 3356 2599 3408 2633
rect 4086 2599 4138 2633
rect 4264 2599 4316 2633
rect 4442 2599 4494 2633
rect 4620 2599 4672 2633
rect 4798 2599 4850 2633
rect 4976 2599 5028 2633
rect 5154 2599 5206 2633
rect 5332 2599 5384 2633
rect 5510 2599 5562 2633
rect 5688 2599 5740 2633
rect 5866 2599 5918 2633
rect 6044 2599 6096 2633
rect 6222 2599 6274 2633
rect 6400 2599 6452 2633
rect 6578 2599 6630 2633
rect 6756 2599 6808 2633
rect 686 2489 738 2523
rect 864 2489 916 2523
rect 1042 2489 1094 2523
rect 1220 2489 1272 2523
rect 1398 2489 1450 2523
rect 1576 2489 1628 2523
rect 1754 2489 1806 2523
rect 1932 2489 1984 2523
rect 2110 2489 2162 2523
rect 2288 2489 2340 2523
rect 2466 2489 2518 2523
rect 2644 2489 2696 2523
rect 2822 2489 2874 2523
rect 3000 2489 3052 2523
rect 3178 2489 3230 2523
rect 3356 2489 3408 2523
rect 4086 2489 4138 2523
rect 4264 2489 4316 2523
rect 4442 2489 4494 2523
rect 4620 2489 4672 2523
rect 4798 2489 4850 2523
rect 4976 2489 5028 2523
rect 5154 2489 5206 2523
rect 5332 2489 5384 2523
rect 5510 2489 5562 2523
rect 5688 2489 5740 2523
rect 5866 2489 5918 2523
rect 6044 2489 6096 2523
rect 6222 2489 6274 2523
rect 6400 2489 6452 2523
rect 6578 2489 6630 2523
rect 6756 2489 6808 2523
rect 606 2405 640 2439
rect 784 2183 818 2217
rect 962 2405 996 2439
rect 1140 2183 1174 2217
rect 1318 2405 1352 2439
rect 1496 2183 1530 2217
rect 1674 2405 1708 2439
rect 1852 2183 1886 2217
rect 2030 2405 2064 2439
rect 2208 2183 2242 2217
rect 2386 2405 2420 2439
rect 2564 2183 2598 2217
rect 2742 2405 2776 2439
rect 2920 2183 2954 2217
rect 3098 2405 3132 2439
rect 3276 2183 3310 2217
rect 3454 2405 3488 2439
rect 4006 2405 4040 2439
rect 4184 2183 4218 2217
rect 4362 2405 4396 2439
rect 4540 2183 4574 2217
rect 4718 2405 4752 2439
rect 4896 2183 4930 2217
rect 5074 2405 5108 2439
rect 5252 2183 5286 2217
rect 5430 2405 5464 2439
rect 5608 2183 5642 2217
rect 5786 2405 5820 2439
rect 5964 2183 5998 2217
rect 6142 2405 6176 2439
rect 6320 2183 6354 2217
rect 6498 2405 6532 2439
rect 6676 2183 6710 2217
rect 6854 2405 6888 2439
rect 686 2099 738 2133
rect 864 2099 916 2133
rect 1042 2099 1094 2133
rect 1220 2099 1272 2133
rect 1398 2099 1450 2133
rect 1576 2099 1628 2133
rect 1754 2099 1806 2133
rect 1932 2099 1984 2133
rect 2110 2099 2162 2133
rect 2288 2099 2340 2133
rect 2466 2099 2518 2133
rect 2644 2099 2696 2133
rect 2822 2099 2874 2133
rect 3000 2099 3052 2133
rect 3178 2099 3230 2133
rect 3356 2099 3408 2133
rect 4086 2099 4138 2133
rect 4264 2099 4316 2133
rect 4442 2099 4494 2133
rect 4620 2099 4672 2133
rect 4798 2099 4850 2133
rect 4976 2099 5028 2133
rect 5154 2099 5206 2133
rect 5332 2099 5384 2133
rect 5510 2099 5562 2133
rect 5688 2099 5740 2133
rect 5866 2099 5918 2133
rect 6044 2099 6096 2133
rect 6222 2099 6274 2133
rect 6400 2099 6452 2133
rect 6578 2099 6630 2133
rect 6756 2099 6808 2133
rect 686 1989 738 2023
rect 864 1989 916 2023
rect 1042 1989 1094 2023
rect 1220 1989 1272 2023
rect 1398 1989 1450 2023
rect 1576 1989 1628 2023
rect 1754 1989 1806 2023
rect 1932 1989 1984 2023
rect 2110 1989 2162 2023
rect 2288 1989 2340 2023
rect 2466 1989 2518 2023
rect 2644 1989 2696 2023
rect 2822 1989 2874 2023
rect 3000 1989 3052 2023
rect 3178 1989 3230 2023
rect 3356 1989 3408 2023
rect 4086 1989 4138 2023
rect 4264 1989 4316 2023
rect 4442 1989 4494 2023
rect 4620 1989 4672 2023
rect 4798 1989 4850 2023
rect 4976 1989 5028 2023
rect 5154 1989 5206 2023
rect 5332 1989 5384 2023
rect 5510 1989 5562 2023
rect 5688 1989 5740 2023
rect 5866 1989 5918 2023
rect 6044 1989 6096 2023
rect 6222 1989 6274 2023
rect 6400 1989 6452 2023
rect 6578 1989 6630 2023
rect 6756 1989 6808 2023
rect 606 1905 640 1939
rect 784 1683 818 1717
rect 962 1905 996 1939
rect 1140 1683 1174 1717
rect 1318 1905 1352 1939
rect 1496 1683 1530 1717
rect 1674 1905 1708 1939
rect 1852 1683 1886 1717
rect 2030 1905 2064 1939
rect 2208 1683 2242 1717
rect 2386 1905 2420 1939
rect 2564 1683 2598 1717
rect 2742 1905 2776 1939
rect 2920 1683 2954 1717
rect 3098 1905 3132 1939
rect 3276 1683 3310 1717
rect 3454 1905 3488 1939
rect 4006 1905 4040 1939
rect 4184 1683 4218 1717
rect 4362 1905 4396 1939
rect 4540 1683 4574 1717
rect 4718 1905 4752 1939
rect 4896 1683 4930 1717
rect 5074 1905 5108 1939
rect 5252 1683 5286 1717
rect 5430 1905 5464 1939
rect 5608 1683 5642 1717
rect 5786 1905 5820 1939
rect 5964 1683 5998 1717
rect 6142 1905 6176 1939
rect 6320 1683 6354 1717
rect 6498 1905 6532 1939
rect 6676 1683 6710 1717
rect 6854 1905 6888 1939
rect 686 1599 738 1633
rect 864 1599 916 1633
rect 1042 1599 1094 1633
rect 1220 1599 1272 1633
rect 1398 1599 1450 1633
rect 1576 1599 1628 1633
rect 1754 1599 1806 1633
rect 1932 1599 1984 1633
rect 2110 1599 2162 1633
rect 2288 1599 2340 1633
rect 2466 1599 2518 1633
rect 2644 1599 2696 1633
rect 2822 1599 2874 1633
rect 3000 1599 3052 1633
rect 3178 1599 3230 1633
rect 3356 1599 3408 1633
rect 4086 1599 4138 1633
rect 4264 1599 4316 1633
rect 4442 1599 4494 1633
rect 4620 1599 4672 1633
rect 4798 1599 4850 1633
rect 4976 1599 5028 1633
rect 5154 1599 5206 1633
rect 5332 1599 5384 1633
rect 5510 1599 5562 1633
rect 5688 1599 5740 1633
rect 5866 1599 5918 1633
rect 6044 1599 6096 1633
rect 6222 1599 6274 1633
rect 6400 1599 6452 1633
rect 6578 1599 6630 1633
rect 6756 1599 6808 1633
rect 686 1489 738 1523
rect 864 1489 916 1523
rect 1042 1489 1094 1523
rect 1220 1489 1272 1523
rect 1398 1489 1450 1523
rect 1576 1489 1628 1523
rect 1754 1489 1806 1523
rect 1932 1489 1984 1523
rect 2110 1489 2162 1523
rect 2288 1489 2340 1523
rect 2466 1489 2518 1523
rect 2644 1489 2696 1523
rect 2822 1489 2874 1523
rect 3000 1489 3052 1523
rect 3178 1489 3230 1523
rect 3356 1489 3408 1523
rect 4086 1489 4138 1523
rect 4264 1489 4316 1523
rect 4442 1489 4494 1523
rect 4620 1489 4672 1523
rect 4798 1489 4850 1523
rect 4976 1489 5028 1523
rect 5154 1489 5206 1523
rect 5332 1489 5384 1523
rect 5510 1489 5562 1523
rect 5688 1489 5740 1523
rect 5866 1489 5918 1523
rect 6044 1489 6096 1523
rect 6222 1489 6274 1523
rect 6400 1489 6452 1523
rect 6578 1489 6630 1523
rect 6756 1489 6808 1523
rect 606 1405 640 1439
rect 784 1183 818 1217
rect 962 1405 996 1439
rect 1140 1183 1174 1217
rect 1318 1405 1352 1439
rect 1496 1183 1530 1217
rect 1674 1405 1708 1439
rect 1852 1183 1886 1217
rect 2030 1405 2064 1439
rect 2208 1183 2242 1217
rect 2386 1405 2420 1439
rect 2564 1183 2598 1217
rect 2742 1405 2776 1439
rect 2920 1183 2954 1217
rect 3098 1405 3132 1439
rect 3276 1183 3310 1217
rect 3454 1405 3488 1439
rect 4006 1405 4040 1439
rect 4184 1183 4218 1217
rect 4362 1405 4396 1439
rect 4540 1183 4574 1217
rect 4718 1405 4752 1439
rect 4896 1183 4930 1217
rect 5074 1405 5108 1439
rect 5252 1183 5286 1217
rect 5430 1405 5464 1439
rect 5608 1183 5642 1217
rect 5786 1405 5820 1439
rect 5964 1183 5998 1217
rect 6142 1405 6176 1439
rect 6320 1183 6354 1217
rect 6498 1405 6532 1439
rect 6676 1183 6710 1217
rect 6854 1405 6888 1439
rect 686 1099 738 1133
rect 864 1099 916 1133
rect 1042 1099 1094 1133
rect 1220 1099 1272 1133
rect 1398 1099 1450 1133
rect 1576 1099 1628 1133
rect 1754 1099 1806 1133
rect 1932 1099 1984 1133
rect 2110 1099 2162 1133
rect 2288 1099 2340 1133
rect 2466 1099 2518 1133
rect 2644 1099 2696 1133
rect 2822 1099 2874 1133
rect 3000 1099 3052 1133
rect 3178 1099 3230 1133
rect 3356 1099 3408 1133
rect 4086 1099 4138 1133
rect 4264 1099 4316 1133
rect 4442 1099 4494 1133
rect 4620 1099 4672 1133
rect 4798 1099 4850 1133
rect 4976 1099 5028 1133
rect 5154 1099 5206 1133
rect 5332 1099 5384 1133
rect 5510 1099 5562 1133
rect 5688 1099 5740 1133
rect 5866 1099 5918 1133
rect 6044 1099 6096 1133
rect 6222 1099 6274 1133
rect 6400 1099 6452 1133
rect 6578 1099 6630 1133
rect 6756 1099 6808 1133
rect 686 989 738 1023
rect 864 989 916 1023
rect 1042 989 1094 1023
rect 1220 989 1272 1023
rect 1398 989 1450 1023
rect 1576 989 1628 1023
rect 1754 989 1806 1023
rect 1932 989 1984 1023
rect 2110 989 2162 1023
rect 2288 989 2340 1023
rect 2466 989 2518 1023
rect 2644 989 2696 1023
rect 2822 989 2874 1023
rect 3000 989 3052 1023
rect 3178 989 3230 1023
rect 3356 989 3408 1023
rect 4086 989 4138 1023
rect 4264 989 4316 1023
rect 4442 989 4494 1023
rect 4620 989 4672 1023
rect 4798 989 4850 1023
rect 4976 989 5028 1023
rect 5154 989 5206 1023
rect 5332 989 5384 1023
rect 5510 989 5562 1023
rect 5688 989 5740 1023
rect 5866 989 5918 1023
rect 6044 989 6096 1023
rect 6222 989 6274 1023
rect 6400 989 6452 1023
rect 6578 989 6630 1023
rect 6756 989 6808 1023
rect 606 905 640 939
rect 784 683 818 717
rect 962 905 996 939
rect 1140 683 1174 717
rect 1318 905 1352 939
rect 1496 683 1530 717
rect 1674 905 1708 939
rect 1852 683 1886 717
rect 2030 905 2064 939
rect 2208 683 2242 717
rect 2386 905 2420 939
rect 2564 683 2598 717
rect 2742 905 2776 939
rect 2920 683 2954 717
rect 3098 905 3132 939
rect 3276 683 3310 717
rect 3454 905 3488 939
rect 4006 905 4040 939
rect 4184 683 4218 717
rect 4362 905 4396 939
rect 4540 683 4574 717
rect 4718 905 4752 939
rect 4896 683 4930 717
rect 5074 905 5108 939
rect 5252 683 5286 717
rect 5430 905 5464 939
rect 5608 683 5642 717
rect 5786 905 5820 939
rect 5964 683 5998 717
rect 6142 905 6176 939
rect 6320 683 6354 717
rect 6498 905 6532 939
rect 6676 683 6710 717
rect 6854 905 6888 939
rect 686 599 738 633
rect 864 599 916 633
rect 1042 599 1094 633
rect 1220 599 1272 633
rect 1398 599 1450 633
rect 1576 599 1628 633
rect 1754 599 1806 633
rect 1932 599 1984 633
rect 2110 599 2162 633
rect 2288 599 2340 633
rect 2466 599 2518 633
rect 2644 599 2696 633
rect 2822 599 2874 633
rect 3000 599 3052 633
rect 3178 599 3230 633
rect 3356 599 3408 633
rect 4086 599 4138 633
rect 4264 599 4316 633
rect 4442 599 4494 633
rect 4620 599 4672 633
rect 4798 599 4850 633
rect 4976 599 5028 633
rect 5154 599 5206 633
rect 5332 599 5384 633
rect 5510 599 5562 633
rect 5688 599 5740 633
rect 5866 599 5918 633
rect 6044 599 6096 633
rect 6222 599 6274 633
rect 6400 599 6452 633
rect 6578 599 6630 633
rect 6756 599 6808 633
rect 7815 3689 7867 3723
rect 7993 3689 8045 3723
rect 8171 3689 8223 3723
rect 8349 3689 8401 3723
rect 8527 3689 8579 3723
rect 8705 3689 8757 3723
rect 8883 3689 8935 3723
rect 9061 3689 9113 3723
rect 9239 3689 9291 3723
rect 9417 3689 9469 3723
rect 9595 3689 9647 3723
rect 9773 3689 9825 3723
rect 10502 3689 10554 3723
rect 10680 3689 10732 3723
rect 10858 3689 10910 3723
rect 11036 3689 11088 3723
rect 11214 3689 11266 3723
rect 11392 3689 11444 3723
rect 11570 3689 11622 3723
rect 11748 3689 11800 3723
rect 11926 3689 11978 3723
rect 12104 3689 12156 3723
rect 12282 3689 12334 3723
rect 12460 3689 12512 3723
rect 7735 3605 7769 3639
rect 7913 3383 7947 3417
rect 8091 3605 8125 3639
rect 8269 3383 8303 3417
rect 8447 3605 8481 3639
rect 8625 3383 8659 3417
rect 8803 3605 8837 3639
rect 8981 3383 9015 3417
rect 9159 3605 9193 3639
rect 9337 3383 9371 3417
rect 9515 3605 9549 3639
rect 9693 3383 9727 3417
rect 9871 3605 9905 3639
rect 10422 3605 10456 3639
rect 10600 3383 10634 3417
rect 10778 3605 10812 3639
rect 10956 3383 10990 3417
rect 11134 3605 11168 3639
rect 11312 3383 11346 3417
rect 11490 3605 11524 3639
rect 11668 3383 11702 3417
rect 11846 3605 11880 3639
rect 12024 3383 12058 3417
rect 12202 3605 12236 3639
rect 12380 3383 12414 3417
rect 12558 3605 12592 3639
rect 7815 3299 7867 3333
rect 7993 3299 8045 3333
rect 8171 3299 8223 3333
rect 8349 3299 8401 3333
rect 8527 3299 8579 3333
rect 8705 3299 8757 3333
rect 8883 3299 8935 3333
rect 9061 3299 9113 3333
rect 9239 3299 9291 3333
rect 9417 3299 9469 3333
rect 9595 3299 9647 3333
rect 9773 3299 9825 3333
rect 10502 3299 10554 3333
rect 10680 3299 10732 3333
rect 10858 3299 10910 3333
rect 11036 3299 11088 3333
rect 11214 3299 11266 3333
rect 11392 3299 11444 3333
rect 11570 3299 11622 3333
rect 11748 3299 11800 3333
rect 11926 3299 11978 3333
rect 12104 3299 12156 3333
rect 12282 3299 12334 3333
rect 12460 3299 12512 3333
rect 7815 3189 7867 3223
rect 7993 3189 8045 3223
rect 8171 3189 8223 3223
rect 8349 3189 8401 3223
rect 8527 3189 8579 3223
rect 8705 3189 8757 3223
rect 8883 3189 8935 3223
rect 9061 3189 9113 3223
rect 9239 3189 9291 3223
rect 9417 3189 9469 3223
rect 9595 3189 9647 3223
rect 9773 3189 9825 3223
rect 10502 3189 10554 3223
rect 10680 3189 10732 3223
rect 10858 3189 10910 3223
rect 11036 3189 11088 3223
rect 11214 3189 11266 3223
rect 11392 3189 11444 3223
rect 11570 3189 11622 3223
rect 11748 3189 11800 3223
rect 11926 3189 11978 3223
rect 12104 3189 12156 3223
rect 12282 3189 12334 3223
rect 12460 3189 12512 3223
rect 7735 3105 7769 3139
rect 7913 2883 7947 2917
rect 8091 3105 8125 3139
rect 8269 2883 8303 2917
rect 8447 3105 8481 3139
rect 8625 2883 8659 2917
rect 8803 3105 8837 3139
rect 8981 2883 9015 2917
rect 9159 3105 9193 3139
rect 9337 2883 9371 2917
rect 9515 3105 9549 3139
rect 9693 2883 9727 2917
rect 9871 3105 9905 3139
rect 10422 3105 10456 3139
rect 10600 2883 10634 2917
rect 10778 3105 10812 3139
rect 10956 2883 10990 2917
rect 11134 3105 11168 3139
rect 11312 2883 11346 2917
rect 11490 3105 11524 3139
rect 11668 2883 11702 2917
rect 11846 3105 11880 3139
rect 12024 2883 12058 2917
rect 12202 3105 12236 3139
rect 12380 2883 12414 2917
rect 12558 3105 12592 3139
rect 7815 2799 7867 2833
rect 7993 2799 8045 2833
rect 8171 2799 8223 2833
rect 8349 2799 8401 2833
rect 8527 2799 8579 2833
rect 8705 2799 8757 2833
rect 8883 2799 8935 2833
rect 9061 2799 9113 2833
rect 9239 2799 9291 2833
rect 9417 2799 9469 2833
rect 9595 2799 9647 2833
rect 9773 2799 9825 2833
rect 10502 2799 10554 2833
rect 10680 2799 10732 2833
rect 10858 2799 10910 2833
rect 11036 2799 11088 2833
rect 11214 2799 11266 2833
rect 11392 2799 11444 2833
rect 11570 2799 11622 2833
rect 11748 2799 11800 2833
rect 11926 2799 11978 2833
rect 12104 2799 12156 2833
rect 12282 2799 12334 2833
rect 12460 2799 12512 2833
rect 7815 2689 7867 2723
rect 7993 2689 8045 2723
rect 8171 2689 8223 2723
rect 8349 2689 8401 2723
rect 8527 2689 8579 2723
rect 8705 2689 8757 2723
rect 8883 2689 8935 2723
rect 9061 2689 9113 2723
rect 9239 2689 9291 2723
rect 9417 2689 9469 2723
rect 9595 2689 9647 2723
rect 9773 2689 9825 2723
rect 10502 2689 10554 2723
rect 10680 2689 10732 2723
rect 10858 2689 10910 2723
rect 11036 2689 11088 2723
rect 11214 2689 11266 2723
rect 11392 2689 11444 2723
rect 11570 2689 11622 2723
rect 11748 2689 11800 2723
rect 11926 2689 11978 2723
rect 12104 2689 12156 2723
rect 12282 2689 12334 2723
rect 12460 2689 12512 2723
rect 7735 2605 7769 2639
rect 7913 2383 7947 2417
rect 8091 2605 8125 2639
rect 8269 2383 8303 2417
rect 8447 2605 8481 2639
rect 8625 2383 8659 2417
rect 8803 2605 8837 2639
rect 8981 2383 9015 2417
rect 9159 2605 9193 2639
rect 9337 2383 9371 2417
rect 9515 2605 9549 2639
rect 9693 2383 9727 2417
rect 9871 2605 9905 2639
rect 10422 2605 10456 2639
rect 10600 2383 10634 2417
rect 10778 2605 10812 2639
rect 10956 2383 10990 2417
rect 11134 2605 11168 2639
rect 11312 2383 11346 2417
rect 11490 2605 11524 2639
rect 11668 2383 11702 2417
rect 11846 2605 11880 2639
rect 12024 2383 12058 2417
rect 12202 2605 12236 2639
rect 12380 2383 12414 2417
rect 12558 2605 12592 2639
rect 7815 2299 7867 2333
rect 7993 2299 8045 2333
rect 8171 2299 8223 2333
rect 8349 2299 8401 2333
rect 8527 2299 8579 2333
rect 8705 2299 8757 2333
rect 8883 2299 8935 2333
rect 9061 2299 9113 2333
rect 9239 2299 9291 2333
rect 9417 2299 9469 2333
rect 9595 2299 9647 2333
rect 9773 2299 9825 2333
rect 10502 2299 10554 2333
rect 10680 2299 10732 2333
rect 10858 2299 10910 2333
rect 11036 2299 11088 2333
rect 11214 2299 11266 2333
rect 11392 2299 11444 2333
rect 11570 2299 11622 2333
rect 11748 2299 11800 2333
rect 11926 2299 11978 2333
rect 12104 2299 12156 2333
rect 12282 2299 12334 2333
rect 12460 2299 12512 2333
rect 7815 1989 7867 2023
rect 7993 1989 8045 2023
rect 8171 1989 8223 2023
rect 8349 1989 8401 2023
rect 8527 1989 8579 2023
rect 8705 1989 8757 2023
rect 8883 1989 8935 2023
rect 9061 1989 9113 2023
rect 9239 1989 9291 2023
rect 9417 1989 9469 2023
rect 9595 1989 9647 2023
rect 9773 1989 9825 2023
rect 10502 1989 10554 2023
rect 10680 1989 10732 2023
rect 10858 1989 10910 2023
rect 11036 1989 11088 2023
rect 11214 1989 11266 2023
rect 11392 1989 11444 2023
rect 11570 1989 11622 2023
rect 11748 1989 11800 2023
rect 11926 1989 11978 2023
rect 12104 1989 12156 2023
rect 12282 1989 12334 2023
rect 12460 1989 12512 2023
rect 7735 1905 7769 1939
rect 7913 1683 7947 1717
rect 8091 1905 8125 1939
rect 8269 1683 8303 1717
rect 8447 1905 8481 1939
rect 8625 1683 8659 1717
rect 8803 1905 8837 1939
rect 8981 1683 9015 1717
rect 9159 1905 9193 1939
rect 9337 1683 9371 1717
rect 9515 1905 9549 1939
rect 9693 1683 9727 1717
rect 9871 1905 9905 1939
rect 10422 1905 10456 1939
rect 10600 1683 10634 1717
rect 10778 1905 10812 1939
rect 10956 1683 10990 1717
rect 11134 1905 11168 1939
rect 11312 1683 11346 1717
rect 11490 1905 11524 1939
rect 11668 1683 11702 1717
rect 11846 1905 11880 1939
rect 12024 1683 12058 1717
rect 12202 1905 12236 1939
rect 12380 1683 12414 1717
rect 12558 1905 12592 1939
rect 7815 1599 7867 1633
rect 7993 1599 8045 1633
rect 8171 1599 8223 1633
rect 8349 1599 8401 1633
rect 8527 1599 8579 1633
rect 8705 1599 8757 1633
rect 8883 1599 8935 1633
rect 9061 1599 9113 1633
rect 9239 1599 9291 1633
rect 9417 1599 9469 1633
rect 9595 1599 9647 1633
rect 9773 1599 9825 1633
rect 10502 1599 10554 1633
rect 10680 1599 10732 1633
rect 10858 1599 10910 1633
rect 11036 1599 11088 1633
rect 11214 1599 11266 1633
rect 11392 1599 11444 1633
rect 11570 1599 11622 1633
rect 11748 1599 11800 1633
rect 11926 1599 11978 1633
rect 12104 1599 12156 1633
rect 12282 1599 12334 1633
rect 12460 1599 12512 1633
rect 7815 1489 7867 1523
rect 7993 1489 8045 1523
rect 8171 1489 8223 1523
rect 8349 1489 8401 1523
rect 8527 1489 8579 1523
rect 8705 1489 8757 1523
rect 8883 1489 8935 1523
rect 9061 1489 9113 1523
rect 9239 1489 9291 1523
rect 9417 1489 9469 1523
rect 9595 1489 9647 1523
rect 9773 1489 9825 1523
rect 10502 1489 10554 1523
rect 10680 1489 10732 1523
rect 10858 1489 10910 1523
rect 11036 1489 11088 1523
rect 11214 1489 11266 1523
rect 11392 1489 11444 1523
rect 11570 1489 11622 1523
rect 11748 1489 11800 1523
rect 11926 1489 11978 1523
rect 12104 1489 12156 1523
rect 12282 1489 12334 1523
rect 12460 1489 12512 1523
rect 7735 1405 7769 1439
rect 7913 1183 7947 1217
rect 8091 1405 8125 1439
rect 8269 1183 8303 1217
rect 8447 1405 8481 1439
rect 8625 1183 8659 1217
rect 8803 1405 8837 1439
rect 8981 1183 9015 1217
rect 9159 1405 9193 1439
rect 9337 1183 9371 1217
rect 9515 1405 9549 1439
rect 9693 1183 9727 1217
rect 9871 1405 9905 1439
rect 10422 1405 10456 1439
rect 10600 1183 10634 1217
rect 10778 1405 10812 1439
rect 10956 1183 10990 1217
rect 11134 1405 11168 1439
rect 11312 1183 11346 1217
rect 11490 1405 11524 1439
rect 11668 1183 11702 1217
rect 11846 1405 11880 1439
rect 12024 1183 12058 1217
rect 12202 1405 12236 1439
rect 12380 1183 12414 1217
rect 12558 1405 12592 1439
rect 7815 1099 7867 1133
rect 7993 1099 8045 1133
rect 8171 1099 8223 1133
rect 8349 1099 8401 1133
rect 8527 1099 8579 1133
rect 8705 1099 8757 1133
rect 8883 1099 8935 1133
rect 9061 1099 9113 1133
rect 9239 1099 9291 1133
rect 9417 1099 9469 1133
rect 9595 1099 9647 1133
rect 9773 1099 9825 1133
rect 10502 1099 10554 1133
rect 10680 1099 10732 1133
rect 10858 1099 10910 1133
rect 11036 1099 11088 1133
rect 11214 1099 11266 1133
rect 11392 1099 11444 1133
rect 11570 1099 11622 1133
rect 11748 1099 11800 1133
rect 11926 1099 11978 1133
rect 12104 1099 12156 1133
rect 12282 1099 12334 1133
rect 12460 1099 12512 1133
rect 7815 989 7867 1023
rect 7993 989 8045 1023
rect 8171 989 8223 1023
rect 8349 989 8401 1023
rect 8527 989 8579 1023
rect 8705 989 8757 1023
rect 8883 989 8935 1023
rect 9061 989 9113 1023
rect 9239 989 9291 1023
rect 9417 989 9469 1023
rect 9595 989 9647 1023
rect 9773 989 9825 1023
rect 10502 989 10554 1023
rect 10680 989 10732 1023
rect 10858 989 10910 1023
rect 11036 989 11088 1023
rect 11214 989 11266 1023
rect 11392 989 11444 1023
rect 11570 989 11622 1023
rect 11748 989 11800 1023
rect 11926 989 11978 1023
rect 12104 989 12156 1023
rect 12282 989 12334 1023
rect 12460 989 12512 1023
rect 7735 905 7769 939
rect 7913 683 7947 717
rect 8091 905 8125 939
rect 8269 683 8303 717
rect 8447 905 8481 939
rect 8625 683 8659 717
rect 8803 905 8837 939
rect 8981 683 9015 717
rect 9159 905 9193 939
rect 9337 683 9371 717
rect 9515 905 9549 939
rect 9693 683 9727 717
rect 9871 905 9905 939
rect 10422 905 10456 939
rect 10600 683 10634 717
rect 10778 905 10812 939
rect 10956 683 10990 717
rect 11134 905 11168 939
rect 11312 683 11346 717
rect 11490 905 11524 939
rect 11668 683 11702 717
rect 11846 905 11880 939
rect 12024 683 12058 717
rect 12202 905 12236 939
rect 12380 683 12414 717
rect 12558 905 12592 939
rect 7815 599 7867 633
rect 7993 599 8045 633
rect 8171 599 8223 633
rect 8349 599 8401 633
rect 8527 599 8579 633
rect 8705 599 8757 633
rect 8883 599 8935 633
rect 9061 599 9113 633
rect 9239 599 9291 633
rect 9417 599 9469 633
rect 9595 599 9647 633
rect 9773 599 9825 633
rect 10502 599 10554 633
rect 10680 599 10732 633
rect 10858 599 10910 633
rect 11036 599 11088 633
rect 11214 599 11266 633
rect 11392 599 11444 633
rect 11570 599 11622 633
rect 11748 599 11800 633
rect 11926 599 11978 633
rect 12104 599 12156 633
rect 12282 599 12334 633
rect 12460 599 12512 633
rect 13808 5097 13860 5131
rect 13986 5097 14038 5131
rect 14164 5097 14216 5131
rect 14342 5097 14394 5131
rect 14520 5097 14572 5131
rect 14698 5097 14750 5131
rect 14876 5097 14928 5131
rect 15054 5097 15106 5131
rect 15232 5097 15284 5131
rect 15410 5097 15462 5131
rect 15588 5097 15640 5131
rect 15766 5097 15818 5131
rect 15944 5097 15996 5131
rect 16122 5097 16174 5131
rect 16300 5097 16352 5131
rect 16478 5097 16530 5131
rect 16656 5097 16708 5131
rect 16834 5097 16886 5131
rect 17012 5097 17064 5131
rect 17190 5097 17242 5131
rect 17368 5097 17420 5131
rect 17546 5097 17598 5131
rect 17724 5097 17776 5131
rect 17902 5097 17954 5131
rect 18080 5097 18132 5131
rect 13728 4791 13762 4825
rect 13906 5013 13940 5047
rect 14084 4791 14118 4825
rect 14262 5013 14296 5047
rect 14440 4791 14474 4825
rect 14618 5013 14652 5047
rect 14796 4791 14830 4825
rect 14974 5013 15008 5047
rect 15152 4791 15186 4825
rect 15330 5013 15364 5047
rect 15508 4791 15542 4825
rect 15686 5013 15720 5047
rect 15864 4791 15898 4825
rect 16042 5013 16076 5047
rect 16220 4791 16254 4825
rect 16398 5013 16432 5047
rect 16576 4791 16610 4825
rect 16754 5013 16788 5047
rect 16932 4791 16966 4825
rect 17110 5013 17144 5047
rect 17288 4791 17322 4825
rect 17466 5013 17500 5047
rect 17644 4791 17678 4825
rect 17822 5013 17856 5047
rect 18000 4791 18034 4825
rect 18178 5013 18212 5047
rect 13808 4707 13860 4741
rect 13986 4707 14038 4741
rect 14164 4707 14216 4741
rect 14342 4707 14394 4741
rect 14520 4707 14572 4741
rect 14698 4707 14750 4741
rect 14876 4707 14928 4741
rect 15054 4707 15106 4741
rect 15232 4707 15284 4741
rect 15410 4707 15462 4741
rect 15588 4707 15640 4741
rect 15766 4707 15818 4741
rect 15944 4707 15996 4741
rect 16122 4707 16174 4741
rect 16300 4707 16352 4741
rect 16478 4707 16530 4741
rect 16656 4707 16708 4741
rect 16834 4707 16886 4741
rect 17012 4707 17064 4741
rect 17190 4707 17242 4741
rect 17368 4707 17420 4741
rect 17546 4707 17598 4741
rect 17724 4707 17776 4741
rect 17902 4707 17954 4741
rect 18080 4707 18132 4741
rect 13808 4597 13860 4631
rect 13986 4597 14038 4631
rect 14164 4597 14216 4631
rect 14342 4597 14394 4631
rect 14520 4597 14572 4631
rect 14698 4597 14750 4631
rect 14876 4597 14928 4631
rect 15054 4597 15106 4631
rect 15232 4597 15284 4631
rect 15410 4597 15462 4631
rect 15588 4597 15640 4631
rect 15766 4597 15818 4631
rect 15944 4597 15996 4631
rect 16122 4597 16174 4631
rect 16300 4597 16352 4631
rect 16478 4597 16530 4631
rect 16656 4597 16708 4631
rect 16834 4597 16886 4631
rect 17012 4597 17064 4631
rect 17190 4597 17242 4631
rect 17368 4597 17420 4631
rect 17546 4597 17598 4631
rect 17724 4597 17776 4631
rect 17902 4597 17954 4631
rect 18080 4597 18132 4631
rect 13728 4291 13762 4325
rect 13906 4513 13940 4547
rect 14084 4291 14118 4325
rect 14262 4513 14296 4547
rect 14440 4291 14474 4325
rect 14618 4513 14652 4547
rect 14796 4291 14830 4325
rect 14974 4513 15008 4547
rect 15152 4291 15186 4325
rect 15330 4513 15364 4547
rect 15508 4291 15542 4325
rect 15686 4513 15720 4547
rect 15864 4291 15898 4325
rect 16042 4513 16076 4547
rect 16220 4291 16254 4325
rect 16398 4513 16432 4547
rect 16576 4291 16610 4325
rect 16754 4513 16788 4547
rect 16932 4291 16966 4325
rect 17110 4513 17144 4547
rect 17288 4291 17322 4325
rect 17466 4513 17500 4547
rect 17644 4291 17678 4325
rect 17822 4513 17856 4547
rect 18000 4291 18034 4325
rect 18178 4513 18212 4547
rect 13808 4207 13860 4241
rect 13986 4207 14038 4241
rect 14164 4207 14216 4241
rect 14342 4207 14394 4241
rect 14520 4207 14572 4241
rect 14698 4207 14750 4241
rect 14876 4207 14928 4241
rect 15054 4207 15106 4241
rect 15232 4207 15284 4241
rect 15410 4207 15462 4241
rect 15588 4207 15640 4241
rect 15766 4207 15818 4241
rect 15944 4207 15996 4241
rect 16122 4207 16174 4241
rect 16300 4207 16352 4241
rect 16478 4207 16530 4241
rect 16656 4207 16708 4241
rect 16834 4207 16886 4241
rect 17012 4207 17064 4241
rect 17190 4207 17242 4241
rect 17368 4207 17420 4241
rect 17546 4207 17598 4241
rect 17724 4207 17776 4241
rect 17902 4207 17954 4241
rect 18080 4207 18132 4241
rect 17366 3593 17418 3627
rect 17544 3593 17596 3627
rect 13756 2588 13808 2622
rect 14048 2588 14100 2622
rect 14340 2588 14392 2622
rect 14632 2588 14684 2622
rect 14924 2588 14976 2622
rect 15216 2588 15268 2622
rect 15508 2588 15560 2622
rect 13676 2282 13710 2538
rect 13854 2282 13888 2538
rect 13968 2282 14002 2538
rect 14146 2282 14180 2538
rect 14260 2282 14294 2538
rect 14438 2282 14472 2538
rect 14552 2282 14586 2538
rect 14730 2282 14764 2538
rect 14844 2282 14878 2538
rect 15022 2282 15056 2538
rect 15136 2282 15170 2538
rect 15314 2282 15348 2538
rect 15428 2282 15462 2538
rect 15606 2282 15640 2538
rect 13756 2198 13808 2232
rect 14048 2198 14100 2232
rect 14340 2198 14392 2232
rect 14632 2198 14684 2232
rect 14924 2198 14976 2232
rect 15216 2198 15268 2232
rect 15508 2198 15560 2232
rect 13756 2090 13808 2124
rect 14048 2090 14100 2124
rect 14340 2090 14392 2124
rect 14632 2090 14684 2124
rect 14924 2090 14976 2124
rect 15216 2090 15268 2124
rect 15508 2090 15560 2124
rect 13676 1784 13710 2040
rect 13854 1784 13888 2040
rect 13968 1784 14002 2040
rect 14146 1784 14180 2040
rect 14260 1784 14294 2040
rect 14438 1784 14472 2040
rect 14552 1784 14586 2040
rect 14730 1784 14764 2040
rect 14844 1784 14878 2040
rect 15022 1784 15056 2040
rect 15136 1784 15170 2040
rect 15314 1784 15348 2040
rect 15428 1784 15462 2040
rect 15606 1784 15640 2040
rect 13756 1700 13808 1734
rect 14048 1700 14100 1734
rect 14340 1700 14392 1734
rect 14632 1700 14684 1734
rect 14924 1700 14976 1734
rect 15216 1700 15268 1734
rect 15508 1700 15560 1734
rect 13756 1592 13808 1626
rect 14048 1592 14100 1626
rect 14340 1592 14392 1626
rect 14632 1592 14684 1626
rect 14924 1592 14976 1626
rect 15216 1592 15268 1626
rect 15508 1592 15560 1626
rect 13676 1286 13710 1542
rect 13854 1286 13888 1542
rect 13968 1286 14002 1542
rect 14146 1286 14180 1542
rect 14260 1286 14294 1542
rect 14438 1286 14472 1542
rect 14552 1286 14586 1542
rect 14730 1286 14764 1542
rect 14844 1286 14878 1542
rect 15022 1286 15056 1542
rect 15136 1286 15170 1542
rect 15314 1286 15348 1542
rect 15428 1286 15462 1542
rect 15606 1286 15640 1542
rect 13756 1202 13808 1236
rect 14048 1202 14100 1236
rect 14340 1202 14392 1236
rect 14632 1202 14684 1236
rect 14924 1202 14976 1236
rect 15216 1202 15268 1236
rect 15508 1202 15560 1236
rect 13756 1094 13808 1128
rect 14048 1094 14100 1128
rect 14340 1094 14392 1128
rect 14632 1094 14684 1128
rect 14924 1094 14976 1128
rect 15216 1094 15268 1128
rect 15508 1094 15560 1128
rect 13676 788 13710 1044
rect 13854 788 13888 1044
rect 13968 788 14002 1044
rect 14146 788 14180 1044
rect 14260 788 14294 1044
rect 14438 788 14472 1044
rect 14552 788 14586 1044
rect 14730 788 14764 1044
rect 14844 788 14878 1044
rect 15022 788 15056 1044
rect 15136 788 15170 1044
rect 15314 788 15348 1044
rect 15428 788 15462 1044
rect 15606 788 15640 1044
rect 13756 704 13808 738
rect 14048 704 14100 738
rect 14340 704 14392 738
rect 14632 704 14684 738
rect 14924 704 14976 738
rect 15216 704 15268 738
rect 15508 704 15560 738
rect 14109 516 14212 613
rect 15279 517 15382 614
rect 17286 3287 17320 3543
rect 17464 3287 17498 3404
rect 17642 3447 17676 3543
rect 17366 3203 17418 3237
rect 17544 3203 17596 3237
rect 16652 2654 16704 2688
rect 16830 2654 16882 2688
rect 17008 2654 17060 2688
rect 17186 2654 17238 2688
rect 17364 2654 17416 2688
rect 17542 2654 17594 2688
rect 17720 2654 17772 2688
rect 17898 2654 17950 2688
rect 18076 2654 18128 2688
rect 16572 2348 16606 2382
rect 16750 2570 16784 2604
rect 16928 2348 16962 2382
rect 17106 2570 17140 2604
rect 17284 2348 17318 2382
rect 17462 2570 17496 2604
rect 17640 2348 17674 2382
rect 17818 2570 17852 2604
rect 17996 2348 18030 2382
rect 18174 2570 18208 2604
rect 16652 2264 16704 2298
rect 16830 2264 16882 2298
rect 17008 2264 17060 2298
rect 17186 2264 17238 2298
rect 17364 2264 17416 2298
rect 17542 2264 17594 2298
rect 17720 2264 17772 2298
rect 17898 2264 17950 2298
rect 18076 2264 18128 2298
rect 16652 2154 16704 2188
rect 16830 2154 16882 2188
rect 17008 2154 17060 2188
rect 17186 2154 17238 2188
rect 17364 2154 17416 2188
rect 17542 2154 17594 2188
rect 17720 2154 17772 2188
rect 17898 2154 17950 2188
rect 18076 2154 18128 2188
rect 16572 1848 16606 1882
rect 16750 2070 16784 2104
rect 16928 1848 16962 1882
rect 17106 2070 17140 2104
rect 17284 1848 17318 1882
rect 17462 2070 17496 2104
rect 17640 1848 17674 1882
rect 17818 2070 17852 2104
rect 17996 1848 18030 1882
rect 18174 2070 18208 2104
rect 16652 1764 16704 1798
rect 16830 1764 16882 1798
rect 17008 1764 17060 1798
rect 17186 1764 17238 1798
rect 17364 1764 17416 1798
rect 17542 1764 17594 1798
rect 17720 1764 17772 1798
rect 17898 1764 17950 1798
rect 18076 1764 18128 1798
rect 16652 1594 16704 1628
rect 16830 1594 16882 1628
rect 17008 1594 17060 1628
rect 17186 1594 17238 1628
rect 17364 1594 17416 1628
rect 17542 1594 17594 1628
rect 17720 1594 17772 1628
rect 17898 1594 17950 1628
rect 18076 1594 18128 1628
rect 16572 1288 16606 1322
rect 16750 1510 16784 1544
rect 16928 1288 16962 1322
rect 17106 1510 17140 1544
rect 17284 1288 17318 1322
rect 17462 1510 17496 1544
rect 17640 1288 17674 1322
rect 17818 1510 17852 1544
rect 17996 1288 18030 1322
rect 18174 1510 18208 1544
rect 16652 1204 16704 1238
rect 16830 1204 16882 1238
rect 17008 1204 17060 1238
rect 17186 1204 17238 1238
rect 17364 1204 17416 1238
rect 17542 1204 17594 1238
rect 17720 1204 17772 1238
rect 17898 1204 17950 1238
rect 18076 1204 18128 1238
rect 16652 1094 16704 1128
rect 16830 1094 16882 1128
rect 17008 1094 17060 1128
rect 17186 1094 17238 1128
rect 17364 1094 17416 1128
rect 17542 1094 17594 1128
rect 17720 1094 17772 1128
rect 17898 1094 17950 1128
rect 18076 1094 18128 1128
rect 16572 788 16606 822
rect 16750 1010 16784 1044
rect 16928 788 16962 822
rect 17106 1010 17140 1044
rect 17284 788 17318 822
rect 17462 1010 17496 1044
rect 17640 788 17674 822
rect 17818 1010 17852 1044
rect 17996 788 18030 822
rect 18174 1010 18208 1044
rect 16652 704 16704 738
rect 16830 704 16882 738
rect 17008 704 17060 738
rect 17186 704 17238 738
rect 17364 704 17416 738
rect 17542 704 17594 738
rect 17720 704 17772 738
rect 17898 704 17950 738
rect 18076 704 18128 738
rect 16547 524 16640 611
rect 17969 513 18062 600
rect 19267 5088 19319 5122
rect 19445 5088 19497 5122
rect 19623 5088 19675 5122
rect 19801 5088 19853 5122
rect 19979 5088 20031 5122
rect 20157 5088 20209 5122
rect 20335 5088 20387 5122
rect 20513 5088 20565 5122
rect 20691 5088 20743 5122
rect 20869 5088 20921 5122
rect 21047 5088 21099 5122
rect 21225 5088 21277 5122
rect 21403 5088 21455 5122
rect 21581 5088 21633 5122
rect 19187 5004 19221 5038
rect 19365 4782 19399 4816
rect 19543 5004 19577 5038
rect 19721 4782 19755 4816
rect 19899 5004 19933 5038
rect 20077 4782 20111 4816
rect 20255 5004 20289 5038
rect 20433 4782 20467 4816
rect 20611 5004 20645 5038
rect 20789 4782 20823 4816
rect 20967 5004 21001 5038
rect 21145 4782 21179 4816
rect 21323 5004 21357 5038
rect 21501 4782 21535 4816
rect 21679 5004 21713 5038
rect 19267 4698 19319 4732
rect 19445 4698 19497 4732
rect 19623 4698 19675 4732
rect 19801 4698 19853 4732
rect 19979 4698 20031 4732
rect 20157 4698 20209 4732
rect 20335 4698 20387 4732
rect 20513 4698 20565 4732
rect 20691 4698 20743 4732
rect 20869 4698 20921 4732
rect 21047 4698 21099 4732
rect 21225 4698 21277 4732
rect 21403 4698 21455 4732
rect 21581 4698 21633 4732
rect 19267 4590 19319 4624
rect 19445 4590 19497 4624
rect 19623 4590 19675 4624
rect 19801 4590 19853 4624
rect 19979 4590 20031 4624
rect 20157 4590 20209 4624
rect 20335 4590 20387 4624
rect 20513 4590 20565 4624
rect 20691 4590 20743 4624
rect 20869 4590 20921 4624
rect 21047 4590 21099 4624
rect 21225 4590 21277 4624
rect 21403 4590 21455 4624
rect 21581 4590 21633 4624
rect 19187 4506 19221 4540
rect 19365 4284 19399 4318
rect 19543 4506 19577 4540
rect 19721 4284 19755 4318
rect 19899 4506 19933 4540
rect 20077 4284 20111 4318
rect 20255 4506 20289 4540
rect 20433 4284 20467 4318
rect 20611 4506 20645 4540
rect 20789 4284 20823 4318
rect 20967 4506 21001 4540
rect 21145 4284 21179 4318
rect 21323 4506 21357 4540
rect 21501 4284 21535 4318
rect 21679 4506 21713 4540
rect 19267 4200 19319 4234
rect 19445 4200 19497 4234
rect 19623 4200 19675 4234
rect 19801 4200 19853 4234
rect 19979 4200 20031 4234
rect 20157 4200 20209 4234
rect 20335 4200 20387 4234
rect 20513 4200 20565 4234
rect 20691 4200 20743 4234
rect 20869 4200 20921 4234
rect 21047 4200 21099 4234
rect 21225 4200 21277 4234
rect 21403 4200 21455 4234
rect 21581 4200 21633 4234
rect 19267 4092 19319 4126
rect 19445 4092 19497 4126
rect 19623 4092 19675 4126
rect 19801 4092 19853 4126
rect 19979 4092 20031 4126
rect 20157 4092 20209 4126
rect 20335 4092 20387 4126
rect 20513 4092 20565 4126
rect 20691 4092 20743 4126
rect 20869 4092 20921 4126
rect 21047 4092 21099 4126
rect 21225 4092 21277 4126
rect 21403 4092 21455 4126
rect 21581 4092 21633 4126
rect 19187 4008 19221 4042
rect 19365 3786 19399 3820
rect 19543 4008 19577 4042
rect 19721 3786 19755 3820
rect 19899 4008 19933 4042
rect 20077 3786 20111 3820
rect 20255 4008 20289 4042
rect 20433 3786 20467 3820
rect 20611 4008 20645 4042
rect 20789 3786 20823 3820
rect 20967 4008 21001 4042
rect 21145 3786 21179 3820
rect 21323 4008 21357 4042
rect 21501 3786 21535 3820
rect 21679 4008 21713 4042
rect 19267 3702 19319 3736
rect 19445 3702 19497 3736
rect 19623 3702 19675 3736
rect 19801 3702 19853 3736
rect 19979 3702 20031 3736
rect 20157 3702 20209 3736
rect 20335 3702 20387 3736
rect 20513 3702 20565 3736
rect 20691 3702 20743 3736
rect 20869 3702 20921 3736
rect 21047 3702 21099 3736
rect 21225 3702 21277 3736
rect 21403 3702 21455 3736
rect 21581 3702 21633 3736
rect 19267 3594 19319 3628
rect 19445 3594 19497 3628
rect 19623 3594 19675 3628
rect 19801 3594 19853 3628
rect 19979 3594 20031 3628
rect 20157 3594 20209 3628
rect 20335 3594 20387 3628
rect 20513 3594 20565 3628
rect 20691 3594 20743 3628
rect 20869 3594 20921 3628
rect 21047 3594 21099 3628
rect 21225 3594 21277 3628
rect 21403 3594 21455 3628
rect 21581 3594 21633 3628
rect 19187 3510 19221 3544
rect 19365 3288 19399 3322
rect 19543 3510 19577 3544
rect 19721 3288 19755 3322
rect 19899 3510 19933 3544
rect 20077 3288 20111 3322
rect 20255 3510 20289 3544
rect 20433 3288 20467 3322
rect 20611 3510 20645 3544
rect 20789 3288 20823 3322
rect 20967 3510 21001 3544
rect 21145 3288 21179 3322
rect 21323 3510 21357 3544
rect 21501 3288 21535 3322
rect 21679 3510 21713 3544
rect 19267 3204 19319 3238
rect 19445 3204 19497 3238
rect 19623 3204 19675 3238
rect 19801 3204 19853 3238
rect 19979 3204 20031 3238
rect 20157 3204 20209 3238
rect 20335 3204 20387 3238
rect 20513 3204 20565 3238
rect 20691 3204 20743 3238
rect 20869 3204 20921 3238
rect 21047 3204 21099 3238
rect 21225 3204 21277 3238
rect 21403 3204 21455 3238
rect 21581 3204 21633 3238
rect 19053 3102 21864 3136
rect 19625 2580 19677 2614
rect 19803 2580 19855 2614
rect 19981 2580 20033 2614
rect 20159 2580 20211 2614
rect 20337 2580 20389 2614
rect 20515 2580 20567 2614
rect 20693 2580 20745 2614
rect 20871 2580 20923 2614
rect 21049 2580 21101 2614
rect 19545 2274 19579 2308
rect 19723 2496 19757 2530
rect 19901 2274 19935 2308
rect 20079 2496 20113 2530
rect 20257 2274 20291 2308
rect 20435 2496 20469 2530
rect 20613 2274 20647 2308
rect 20791 2496 20825 2530
rect 20969 2274 21003 2308
rect 21147 2496 21181 2530
rect 19625 2190 19677 2224
rect 19803 2190 19855 2224
rect 19981 2190 20033 2224
rect 20159 2190 20211 2224
rect 20337 2190 20389 2224
rect 20515 2190 20567 2224
rect 20693 2190 20745 2224
rect 20871 2190 20923 2224
rect 21049 2190 21101 2224
rect 19625 2082 19677 2116
rect 19803 2082 19855 2116
rect 19981 2082 20033 2116
rect 20159 2082 20211 2116
rect 20337 2082 20389 2116
rect 20515 2082 20567 2116
rect 20693 2082 20745 2116
rect 20871 2082 20923 2116
rect 21049 2082 21101 2116
rect 19545 1776 19579 1810
rect 19723 1998 19757 2032
rect 19901 1776 19935 1810
rect 20079 1998 20113 2032
rect 20257 1776 20291 1810
rect 20435 1998 20469 2032
rect 20613 1776 20647 1810
rect 20791 1998 20825 2032
rect 20969 1776 21003 1810
rect 21147 1998 21181 2032
rect 19625 1692 19677 1726
rect 19803 1692 19855 1726
rect 19981 1692 20033 1726
rect 20159 1692 20211 1726
rect 20337 1692 20389 1726
rect 20515 1692 20567 1726
rect 20693 1692 20745 1726
rect 20871 1692 20923 1726
rect 21049 1692 21101 1726
rect 19625 1584 19677 1618
rect 19803 1584 19855 1618
rect 19981 1584 20033 1618
rect 20159 1584 20211 1618
rect 20337 1584 20389 1618
rect 20515 1584 20567 1618
rect 20693 1584 20745 1618
rect 20871 1584 20923 1618
rect 21049 1584 21101 1618
rect 19545 1308 19579 1342
rect 19723 1470 19757 1504
rect 19901 1308 19935 1342
rect 20079 1470 20113 1504
rect 20257 1308 20291 1342
rect 20435 1470 20469 1504
rect 20613 1308 20647 1342
rect 20791 1470 20825 1504
rect 20969 1308 21003 1342
rect 21147 1470 21181 1504
rect 19625 1194 19677 1228
rect 19803 1194 19855 1228
rect 19981 1194 20033 1228
rect 20159 1194 20211 1228
rect 20337 1194 20389 1228
rect 20515 1194 20567 1228
rect 20693 1194 20745 1228
rect 20871 1194 20923 1228
rect 21049 1194 21101 1228
rect 19625 1086 19677 1120
rect 19803 1086 19855 1120
rect 19981 1086 20033 1120
rect 20159 1086 20211 1120
rect 20337 1086 20389 1120
rect 20515 1086 20567 1120
rect 20693 1086 20745 1120
rect 20871 1086 20923 1120
rect 21049 1086 21101 1120
rect 19545 810 19579 844
rect 19723 972 19757 1006
rect 19901 810 19935 844
rect 20079 972 20113 1006
rect 20257 810 20291 844
rect 20435 972 20469 1006
rect 20613 810 20647 844
rect 20791 972 20825 1006
rect 20969 810 21003 844
rect 21147 972 21181 1006
rect 19625 696 19677 730
rect 19803 696 19855 730
rect 19981 696 20033 730
rect 20159 696 20211 730
rect 20337 696 20389 730
rect 20515 696 20567 730
rect 20693 696 20745 730
rect 20871 696 20923 730
rect 21049 696 21101 730
rect 19349 594 21377 628
rect 304 22 13205 71
rect 14118 70 14211 129
rect 15279 70 15372 123
rect 16542 70 16635 127
rect 17969 70 18062 122
rect 13476 21 18366 70
<< metal1 >>
rect 7399 18903 8447 18937
rect 7276 18783 7286 18847
rect 7350 18783 7360 18847
rect 7399 18753 7433 18903
rect 7591 18753 7625 18903
rect 7783 18753 7817 18903
rect 7975 18753 8009 18903
rect 8167 18753 8201 18903
rect 8236 18783 8246 18847
rect 8310 18783 8320 18847
rect 7297 18741 7343 18753
rect 7297 18493 7303 18741
rect 7337 18493 7343 18741
rect 7297 18481 7343 18493
rect 7393 18741 7439 18753
rect 7393 18493 7399 18741
rect 7433 18493 7439 18741
rect 7393 18481 7439 18493
rect 7489 18741 7535 18753
rect 7489 18493 7495 18741
rect 7529 18493 7535 18741
rect 7489 18481 7535 18493
rect 7585 18741 7631 18753
rect 7585 18493 7591 18741
rect 7625 18493 7631 18741
rect 7585 18481 7631 18493
rect 7681 18741 7727 18753
rect 7681 18493 7687 18741
rect 7721 18493 7727 18741
rect 7681 18481 7727 18493
rect 7777 18741 7823 18753
rect 7777 18493 7783 18741
rect 7817 18493 7823 18741
rect 7777 18481 7823 18493
rect 7873 18741 7919 18753
rect 7873 18493 7879 18741
rect 7913 18493 7919 18741
rect 7873 18481 7919 18493
rect 7969 18741 8015 18753
rect 7969 18493 7975 18741
rect 8009 18493 8015 18741
rect 7969 18481 8015 18493
rect 8065 18741 8111 18753
rect 8065 18493 8071 18741
rect 8105 18493 8111 18741
rect 8065 18481 8111 18493
rect 8161 18741 8207 18753
rect 8161 18493 8167 18741
rect 8201 18493 8207 18741
rect 8161 18481 8207 18493
rect 8257 18741 8303 18753
rect 8257 18493 8263 18741
rect 8297 18493 8303 18741
rect 8257 18481 8303 18493
rect 5695 18360 7067 18432
rect 7303 18360 7337 18481
rect 5695 18340 7337 18360
rect 7495 18340 7529 18481
rect 7687 18340 7721 18481
rect 7879 18340 7913 18481
rect 8071 18340 8105 18481
rect 8263 18354 8297 18481
rect 8413 18360 8447 18903
rect 20329 18903 21377 18937
rect 20206 18787 20216 18851
rect 20280 18787 20290 18851
rect 20329 18753 20363 18903
rect 20521 18753 20555 18903
rect 20713 18753 20747 18903
rect 20905 18753 20939 18903
rect 21097 18753 21131 18903
rect 21170 18790 21180 18854
rect 21244 18790 21254 18854
rect 20227 18741 20273 18753
rect 20227 18493 20233 18741
rect 20267 18493 20273 18741
rect 20227 18481 20273 18493
rect 20323 18741 20369 18753
rect 20323 18493 20329 18741
rect 20363 18493 20369 18741
rect 20323 18481 20369 18493
rect 20419 18741 20465 18753
rect 20419 18493 20425 18741
rect 20459 18493 20465 18741
rect 20419 18481 20465 18493
rect 20515 18741 20561 18753
rect 20515 18493 20521 18741
rect 20555 18493 20561 18741
rect 20515 18481 20561 18493
rect 20611 18741 20657 18753
rect 20611 18493 20617 18741
rect 20651 18493 20657 18741
rect 20611 18481 20657 18493
rect 20707 18741 20753 18753
rect 20707 18493 20713 18741
rect 20747 18493 20753 18741
rect 20707 18481 20753 18493
rect 20803 18741 20849 18753
rect 20803 18493 20809 18741
rect 20843 18493 20849 18741
rect 20803 18481 20849 18493
rect 20899 18741 20945 18753
rect 20899 18493 20905 18741
rect 20939 18493 20945 18741
rect 20899 18481 20945 18493
rect 20995 18741 21041 18753
rect 20995 18493 21001 18741
rect 21035 18493 21041 18741
rect 20995 18481 21041 18493
rect 21091 18741 21137 18753
rect 21091 18493 21097 18741
rect 21131 18493 21137 18741
rect 21091 18481 21137 18493
rect 21187 18741 21233 18753
rect 21187 18493 21193 18741
rect 21227 18493 21233 18741
rect 21187 18481 21233 18493
rect 8413 18356 10736 18360
rect 20233 18356 20267 18481
rect 8219 18340 8229 18354
rect 5695 18306 8229 18340
rect 5695 18296 7337 18306
rect 5695 18225 7067 18296
rect 5695 13485 5902 18225
rect 7303 18175 7337 18296
rect 7495 18175 7529 18306
rect 7687 18175 7721 18306
rect 7879 18175 7913 18306
rect 8071 18175 8105 18306
rect 8219 18290 8229 18306
rect 8293 18290 8303 18354
rect 8413 18296 13482 18356
rect 8263 18175 8297 18290
rect 7297 18163 7343 18175
rect 7297 18083 7303 18163
rect 7337 18083 7343 18163
rect 7297 18071 7343 18083
rect 7393 18163 7439 18175
rect 7393 18083 7399 18163
rect 7433 18083 7439 18163
rect 7393 18071 7439 18083
rect 7489 18163 7535 18175
rect 7489 18083 7495 18163
rect 7529 18083 7535 18163
rect 7489 18071 7535 18083
rect 7585 18163 7631 18175
rect 7585 18083 7591 18163
rect 7625 18083 7631 18163
rect 7585 18071 7631 18083
rect 7681 18163 7727 18175
rect 7681 18083 7687 18163
rect 7721 18083 7727 18163
rect 7681 18071 7727 18083
rect 7777 18163 7823 18175
rect 7777 18083 7783 18163
rect 7817 18083 7823 18163
rect 7777 18071 7823 18083
rect 7873 18163 7919 18175
rect 7873 18083 7879 18163
rect 7913 18083 7919 18163
rect 7873 18071 7919 18083
rect 7969 18163 8015 18175
rect 7969 18083 7975 18163
rect 8009 18083 8015 18163
rect 7969 18071 8015 18083
rect 8065 18163 8111 18175
rect 8065 18083 8071 18163
rect 8105 18083 8111 18163
rect 8065 18071 8111 18083
rect 8161 18163 8207 18175
rect 8161 18083 8167 18163
rect 8201 18083 8207 18163
rect 8161 18071 8207 18083
rect 8257 18163 8303 18175
rect 8257 18083 8263 18163
rect 8297 18083 8303 18163
rect 8257 18071 8303 18083
rect 7282 17977 7292 18041
rect 7356 17977 7366 18041
rect 7399 17929 7433 18071
rect 7591 17929 7625 18071
rect 7783 17929 7817 18071
rect 7975 17929 8009 18071
rect 8167 17929 8201 18071
rect 8237 17973 8247 18037
rect 8311 17973 8321 18037
rect 8413 17929 8447 18296
rect 10586 18292 13482 18296
rect 17752 18292 17762 18356
rect 17826 18340 20267 18356
rect 20425 18340 20459 18481
rect 20617 18340 20651 18481
rect 20809 18340 20843 18481
rect 21001 18340 21035 18481
rect 21193 18340 21227 18481
rect 17826 18306 21227 18340
rect 17826 18292 20267 18306
rect 7399 17895 8447 17929
rect 7399 17103 8447 17137
rect 7277 16987 7287 17051
rect 7351 16987 7361 17051
rect 7399 16953 7433 17103
rect 7591 16953 7625 17103
rect 7783 16953 7817 17103
rect 7975 16953 8009 17103
rect 8167 16953 8201 17103
rect 8239 16990 8249 17054
rect 8313 16990 8323 17054
rect 7297 16941 7343 16953
rect 7297 16693 7303 16941
rect 7337 16693 7343 16941
rect 7297 16681 7343 16693
rect 7393 16941 7439 16953
rect 7393 16693 7399 16941
rect 7433 16693 7439 16941
rect 7393 16681 7439 16693
rect 7489 16941 7535 16953
rect 7489 16693 7495 16941
rect 7529 16693 7535 16941
rect 7489 16681 7535 16693
rect 7585 16941 7631 16953
rect 7585 16693 7591 16941
rect 7625 16693 7631 16941
rect 7585 16681 7631 16693
rect 7681 16941 7727 16953
rect 7681 16693 7687 16941
rect 7721 16693 7727 16941
rect 7681 16681 7727 16693
rect 7777 16941 7823 16953
rect 7777 16693 7783 16941
rect 7817 16693 7823 16941
rect 7777 16681 7823 16693
rect 7873 16941 7919 16953
rect 7873 16693 7879 16941
rect 7913 16693 7919 16941
rect 7873 16681 7919 16693
rect 7969 16941 8015 16953
rect 7969 16693 7975 16941
rect 8009 16693 8015 16941
rect 7969 16681 8015 16693
rect 8065 16941 8111 16953
rect 8065 16693 8071 16941
rect 8105 16693 8111 16941
rect 8065 16681 8111 16693
rect 8161 16941 8207 16953
rect 8161 16693 8167 16941
rect 8201 16693 8207 16941
rect 8161 16681 8207 16693
rect 8257 16941 8303 16953
rect 8257 16693 8263 16941
rect 8297 16693 8303 16941
rect 8257 16681 8303 16693
rect 5451 13073 5457 13485
rect 5869 13073 5902 13485
rect 5695 9392 5902 13073
rect 6307 16558 7075 16612
rect 7303 16558 7337 16681
rect 6307 16540 7337 16558
rect 7495 16540 7529 16681
rect 7687 16540 7721 16681
rect 7879 16540 7913 16681
rect 8071 16540 8105 16681
rect 8263 16554 8297 16681
rect 8213 16540 8223 16554
rect 6307 16506 8223 16540
rect 6307 16494 7337 16506
rect 6307 16405 7075 16494
rect 6307 11637 6514 16405
rect 7303 16375 7337 16494
rect 7495 16375 7529 16506
rect 7687 16375 7721 16506
rect 7879 16375 7913 16506
rect 8071 16375 8105 16506
rect 8213 16490 8223 16506
rect 8287 16490 8297 16554
rect 8263 16375 8297 16490
rect 8413 16553 8447 17103
rect 12689 17071 12699 17135
rect 12763 17071 12773 17135
rect 8413 16552 10640 16553
rect 8413 16489 10594 16552
rect 7297 16363 7343 16375
rect 7297 16283 7303 16363
rect 7337 16283 7343 16363
rect 7297 16271 7343 16283
rect 7393 16363 7439 16375
rect 7393 16283 7399 16363
rect 7433 16283 7439 16363
rect 7393 16271 7439 16283
rect 7489 16363 7535 16375
rect 7489 16283 7495 16363
rect 7529 16283 7535 16363
rect 7489 16271 7535 16283
rect 7585 16363 7631 16375
rect 7585 16283 7591 16363
rect 7625 16283 7631 16363
rect 7585 16271 7631 16283
rect 7681 16363 7727 16375
rect 7681 16283 7687 16363
rect 7721 16283 7727 16363
rect 7681 16271 7727 16283
rect 7777 16363 7823 16375
rect 7777 16283 7783 16363
rect 7817 16283 7823 16363
rect 7777 16271 7823 16283
rect 7873 16363 7919 16375
rect 7873 16283 7879 16363
rect 7913 16283 7919 16363
rect 7873 16271 7919 16283
rect 7969 16363 8015 16375
rect 7969 16283 7975 16363
rect 8009 16283 8015 16363
rect 7969 16271 8015 16283
rect 8065 16363 8111 16375
rect 8065 16283 8071 16363
rect 8105 16283 8111 16363
rect 8065 16271 8111 16283
rect 8161 16363 8207 16375
rect 8161 16283 8167 16363
rect 8201 16283 8207 16363
rect 8161 16271 8207 16283
rect 8257 16363 8303 16375
rect 8257 16283 8263 16363
rect 8297 16283 8303 16363
rect 8257 16271 8303 16283
rect 7280 16176 7290 16240
rect 7354 16176 7364 16240
rect 7399 16129 7433 16271
rect 7591 16129 7625 16271
rect 7783 16129 7817 16271
rect 7975 16129 8009 16271
rect 8167 16129 8201 16271
rect 8238 16176 8248 16240
rect 8312 16176 8322 16240
rect 8413 16129 8447 16489
rect 10584 16488 10594 16489
rect 10658 16488 10668 16552
rect 7399 16095 8447 16129
rect 7399 15303 8447 15337
rect 7276 15186 7286 15250
rect 7350 15186 7360 15250
rect 7399 15153 7433 15303
rect 7591 15153 7625 15303
rect 7783 15153 7817 15303
rect 7975 15153 8009 15303
rect 8167 15153 8201 15303
rect 8237 15186 8247 15250
rect 8311 15186 8321 15250
rect 7297 15141 7343 15153
rect 7297 14893 7303 15141
rect 7337 14893 7343 15141
rect 7297 14881 7343 14893
rect 7393 15141 7439 15153
rect 7393 14893 7399 15141
rect 7433 14893 7439 15141
rect 7393 14881 7439 14893
rect 7489 15141 7535 15153
rect 7489 14893 7495 15141
rect 7529 14893 7535 15141
rect 7489 14881 7535 14893
rect 7585 15141 7631 15153
rect 7585 14893 7591 15141
rect 7625 14893 7631 15141
rect 7585 14881 7631 14893
rect 7681 15141 7727 15153
rect 7681 14893 7687 15141
rect 7721 14893 7727 15141
rect 7681 14881 7727 14893
rect 7777 15141 7823 15153
rect 7777 14893 7783 15141
rect 7817 14893 7823 15141
rect 7777 14881 7823 14893
rect 7873 15141 7919 15153
rect 7873 14893 7879 15141
rect 7913 14893 7919 15141
rect 7873 14881 7919 14893
rect 7969 15141 8015 15153
rect 7969 14893 7975 15141
rect 8009 14893 8015 15141
rect 7969 14881 8015 14893
rect 8065 15141 8111 15153
rect 8065 14893 8071 15141
rect 8105 14893 8111 15141
rect 8065 14881 8111 14893
rect 8161 15141 8207 15153
rect 8161 14893 8167 15141
rect 8201 14893 8207 15141
rect 8161 14881 8207 14893
rect 8257 15141 8303 15153
rect 8257 14893 8263 15141
rect 8297 14893 8303 15141
rect 8257 14881 8303 14893
rect 6792 14759 6999 14827
rect 7303 14759 7337 14881
rect 6792 14740 7337 14759
rect 7495 14740 7529 14881
rect 7687 14740 7721 14881
rect 7879 14740 7913 14881
rect 8071 14740 8105 14881
rect 8263 14754 8297 14881
rect 8413 14757 8447 15303
rect 8217 14740 8227 14754
rect 6792 14706 8227 14740
rect 6792 14695 7337 14706
rect 6792 14689 6999 14695
rect 6792 14170 6815 14689
rect 6910 14170 6999 14689
rect 7303 14575 7337 14695
rect 7495 14575 7529 14706
rect 7687 14575 7721 14706
rect 7879 14575 7913 14706
rect 8071 14575 8105 14706
rect 8217 14690 8227 14706
rect 8291 14690 8301 14754
rect 8413 14753 10697 14757
rect 8413 14693 10637 14753
rect 8263 14575 8297 14690
rect 7297 14563 7343 14575
rect 7297 14483 7303 14563
rect 7337 14483 7343 14563
rect 7297 14471 7343 14483
rect 7393 14563 7439 14575
rect 7393 14483 7399 14563
rect 7433 14483 7439 14563
rect 7393 14471 7439 14483
rect 7489 14563 7535 14575
rect 7489 14483 7495 14563
rect 7529 14483 7535 14563
rect 7489 14471 7535 14483
rect 7585 14563 7631 14575
rect 7585 14483 7591 14563
rect 7625 14483 7631 14563
rect 7585 14471 7631 14483
rect 7681 14563 7727 14575
rect 7681 14483 7687 14563
rect 7721 14483 7727 14563
rect 7681 14471 7727 14483
rect 7777 14563 7823 14575
rect 7777 14483 7783 14563
rect 7817 14483 7823 14563
rect 7777 14471 7823 14483
rect 7873 14563 7919 14575
rect 7873 14483 7879 14563
rect 7913 14483 7919 14563
rect 7873 14471 7919 14483
rect 7969 14563 8015 14575
rect 7969 14483 7975 14563
rect 8009 14483 8015 14563
rect 7969 14471 8015 14483
rect 8065 14563 8111 14575
rect 8065 14483 8071 14563
rect 8105 14483 8111 14563
rect 8065 14471 8111 14483
rect 8161 14563 8207 14575
rect 8161 14483 8167 14563
rect 8201 14483 8207 14563
rect 8161 14471 8207 14483
rect 8257 14563 8303 14575
rect 8257 14483 8263 14563
rect 8297 14483 8303 14563
rect 8257 14471 8303 14483
rect 7278 14373 7288 14437
rect 7352 14373 7362 14437
rect 7399 14329 7433 14471
rect 7591 14329 7625 14471
rect 7783 14329 7817 14471
rect 7975 14329 8009 14471
rect 8167 14329 8201 14471
rect 8240 14376 8250 14440
rect 8314 14376 8324 14440
rect 8413 14329 8447 14693
rect 10627 14689 10637 14693
rect 10701 14689 10711 14753
rect 12699 14505 12763 17071
rect 13418 15222 13482 18292
rect 20233 18175 20267 18292
rect 20425 18175 20459 18306
rect 20617 18175 20651 18306
rect 20809 18175 20843 18306
rect 21001 18175 21035 18306
rect 21193 18175 21227 18306
rect 21343 18427 21377 18903
rect 21343 18220 22617 18427
rect 20227 18163 20273 18175
rect 20227 18083 20233 18163
rect 20267 18083 20273 18163
rect 20227 18071 20273 18083
rect 20323 18163 20369 18175
rect 20323 18083 20329 18163
rect 20363 18083 20369 18163
rect 20323 18071 20369 18083
rect 20419 18163 20465 18175
rect 20419 18083 20425 18163
rect 20459 18083 20465 18163
rect 20419 18071 20465 18083
rect 20515 18163 20561 18175
rect 20515 18083 20521 18163
rect 20555 18083 20561 18163
rect 20515 18071 20561 18083
rect 20611 18163 20657 18175
rect 20611 18083 20617 18163
rect 20651 18083 20657 18163
rect 20611 18071 20657 18083
rect 20707 18163 20753 18175
rect 20707 18083 20713 18163
rect 20747 18083 20753 18163
rect 20707 18071 20753 18083
rect 20803 18163 20849 18175
rect 20803 18083 20809 18163
rect 20843 18083 20849 18163
rect 20803 18071 20849 18083
rect 20899 18163 20945 18175
rect 20899 18083 20905 18163
rect 20939 18083 20945 18163
rect 20899 18071 20945 18083
rect 20995 18163 21041 18175
rect 20995 18083 21001 18163
rect 21035 18083 21041 18163
rect 20995 18071 21041 18083
rect 21091 18163 21137 18175
rect 21091 18083 21097 18163
rect 21131 18083 21137 18163
rect 21091 18071 21137 18083
rect 21187 18163 21233 18175
rect 21187 18083 21193 18163
rect 21227 18083 21233 18163
rect 21187 18071 21233 18083
rect 20205 17971 20215 18035
rect 20279 17971 20289 18035
rect 20329 17929 20363 18071
rect 20521 17929 20555 18071
rect 20713 17929 20747 18071
rect 20905 17929 20939 18071
rect 21097 17929 21131 18071
rect 21172 17974 21182 18038
rect 21246 17974 21256 18038
rect 21343 17929 21377 18220
rect 20329 17895 21377 17929
rect 20329 17103 21377 17137
rect 20209 16991 20219 17055
rect 20283 16991 20293 17055
rect 20329 16953 20363 17103
rect 20521 16953 20555 17103
rect 20713 16953 20747 17103
rect 20905 16953 20939 17103
rect 21097 16953 21131 17103
rect 21169 16989 21179 17053
rect 21243 16989 21253 17053
rect 20227 16941 20273 16953
rect 20227 16693 20233 16941
rect 20267 16693 20273 16941
rect 20227 16681 20273 16693
rect 20323 16941 20369 16953
rect 20323 16693 20329 16941
rect 20363 16693 20369 16941
rect 20323 16681 20369 16693
rect 20419 16941 20465 16953
rect 20419 16693 20425 16941
rect 20459 16693 20465 16941
rect 20419 16681 20465 16693
rect 20515 16941 20561 16953
rect 20515 16693 20521 16941
rect 20555 16693 20561 16941
rect 20515 16681 20561 16693
rect 20611 16941 20657 16953
rect 20611 16693 20617 16941
rect 20651 16693 20657 16941
rect 20611 16681 20657 16693
rect 20707 16941 20753 16953
rect 20707 16693 20713 16941
rect 20747 16693 20753 16941
rect 20707 16681 20753 16693
rect 20803 16941 20849 16953
rect 20803 16693 20809 16941
rect 20843 16693 20849 16941
rect 20803 16681 20849 16693
rect 20899 16941 20945 16953
rect 20899 16693 20905 16941
rect 20939 16693 20945 16941
rect 20899 16681 20945 16693
rect 20995 16941 21041 16953
rect 20995 16693 21001 16941
rect 21035 16693 21041 16941
rect 20995 16681 21041 16693
rect 21091 16941 21137 16953
rect 21091 16693 21097 16941
rect 21131 16693 21137 16941
rect 21091 16681 21137 16693
rect 21187 16941 21233 16953
rect 21187 16693 21193 16941
rect 21227 16693 21233 16941
rect 21187 16681 21233 16693
rect 17799 16554 17893 16555
rect 17765 16490 17775 16554
rect 17839 16552 17893 16554
rect 20233 16552 20267 16681
rect 17839 16540 20267 16552
rect 20425 16540 20459 16681
rect 20617 16540 20651 16681
rect 20809 16540 20843 16681
rect 21001 16540 21035 16681
rect 21193 16540 21227 16681
rect 17839 16506 21227 16540
rect 17839 16490 20267 16506
rect 17799 16488 20267 16490
rect 20233 16375 20267 16488
rect 20425 16375 20459 16506
rect 20617 16375 20651 16506
rect 20809 16375 20843 16506
rect 21001 16375 21035 16506
rect 21193 16375 21227 16506
rect 21343 16624 21377 17103
rect 21343 16417 22051 16624
rect 20227 16363 20273 16375
rect 20227 16283 20233 16363
rect 20267 16283 20273 16363
rect 20227 16271 20273 16283
rect 20323 16363 20369 16375
rect 20323 16283 20329 16363
rect 20363 16283 20369 16363
rect 20323 16271 20369 16283
rect 20419 16363 20465 16375
rect 20419 16283 20425 16363
rect 20459 16283 20465 16363
rect 20419 16271 20465 16283
rect 20515 16363 20561 16375
rect 20515 16283 20521 16363
rect 20555 16283 20561 16363
rect 20515 16271 20561 16283
rect 20611 16363 20657 16375
rect 20611 16283 20617 16363
rect 20651 16283 20657 16363
rect 20611 16271 20657 16283
rect 20707 16363 20753 16375
rect 20707 16283 20713 16363
rect 20747 16283 20753 16363
rect 20707 16271 20753 16283
rect 20803 16363 20849 16375
rect 20803 16283 20809 16363
rect 20843 16283 20849 16363
rect 20803 16271 20849 16283
rect 20899 16363 20945 16375
rect 20899 16283 20905 16363
rect 20939 16283 20945 16363
rect 20899 16271 20945 16283
rect 20995 16363 21041 16375
rect 20995 16283 21001 16363
rect 21035 16283 21041 16363
rect 20995 16271 21041 16283
rect 21091 16363 21137 16375
rect 21091 16283 21097 16363
rect 21131 16283 21137 16363
rect 21091 16271 21137 16283
rect 21187 16363 21233 16375
rect 21187 16283 21193 16363
rect 21227 16283 21233 16363
rect 21187 16271 21233 16283
rect 14218 16153 14228 16217
rect 14292 16153 14302 16217
rect 20208 16175 20218 16239
rect 20282 16175 20292 16239
rect 14228 15743 14292 16153
rect 20329 16129 20363 16271
rect 20521 16129 20555 16271
rect 20713 16129 20747 16271
rect 20905 16129 20939 16271
rect 21097 16129 21131 16271
rect 21167 16174 21177 16238
rect 21241 16174 21251 16238
rect 21343 16129 21377 16417
rect 20329 16095 21377 16129
rect 14218 15679 14228 15743
rect 14292 15679 14302 15743
rect 14902 15587 17237 15591
rect 14829 15523 14839 15587
rect 14903 15527 17237 15587
rect 17301 15527 17311 15591
rect 14903 15523 14913 15527
rect 20329 15303 21377 15337
rect 13418 15158 14177 15222
rect 14241 15158 14251 15222
rect 20208 15189 20218 15253
rect 20282 15189 20292 15253
rect 20329 15153 20363 15303
rect 20521 15153 20555 15303
rect 20713 15153 20747 15303
rect 20905 15153 20939 15303
rect 21097 15153 21131 15303
rect 21169 15188 21179 15252
rect 21243 15188 21253 15252
rect 20227 15141 20273 15153
rect 15945 14985 16278 15049
rect 16342 14985 16352 15049
rect 14369 14807 14379 14871
rect 14443 14807 14453 14871
rect 14379 14744 14443 14807
rect 12699 14441 12937 14505
rect 7399 14295 8447 14329
rect 6792 12960 6999 14170
rect 11394 14078 11404 14142
rect 11468 14078 12702 14142
rect 12766 14078 12776 14142
rect 12873 13813 12937 14441
rect 11394 13749 11404 13813
rect 11468 13749 12937 13813
rect 7399 13503 8447 13537
rect 7275 13384 7285 13448
rect 7349 13384 7359 13448
rect 7399 13353 7433 13503
rect 7591 13353 7625 13503
rect 7783 13353 7817 13503
rect 7975 13353 8009 13503
rect 8167 13353 8201 13503
rect 8242 13386 8252 13450
rect 8316 13386 8326 13450
rect 7297 13341 7343 13353
rect 7297 13093 7303 13341
rect 7337 13093 7343 13341
rect 7297 13081 7343 13093
rect 7393 13341 7439 13353
rect 7393 13093 7399 13341
rect 7433 13093 7439 13341
rect 7393 13081 7439 13093
rect 7489 13341 7535 13353
rect 7489 13093 7495 13341
rect 7529 13093 7535 13341
rect 7489 13081 7535 13093
rect 7585 13341 7631 13353
rect 7585 13093 7591 13341
rect 7625 13093 7631 13341
rect 7585 13081 7631 13093
rect 7681 13341 7727 13353
rect 7681 13093 7687 13341
rect 7721 13093 7727 13341
rect 7681 13081 7727 13093
rect 7777 13341 7823 13353
rect 7777 13093 7783 13341
rect 7817 13093 7823 13341
rect 7777 13081 7823 13093
rect 7873 13341 7919 13353
rect 7873 13093 7879 13341
rect 7913 13093 7919 13341
rect 7873 13081 7919 13093
rect 7969 13341 8015 13353
rect 7969 13093 7975 13341
rect 8009 13093 8015 13341
rect 7969 13081 8015 13093
rect 8065 13341 8111 13353
rect 8065 13093 8071 13341
rect 8105 13093 8111 13341
rect 8065 13081 8111 13093
rect 8161 13341 8207 13353
rect 8161 13093 8167 13341
rect 8201 13093 8207 13341
rect 8161 13081 8207 13093
rect 8257 13341 8303 13353
rect 8257 13093 8263 13341
rect 8297 13093 8303 13341
rect 8257 13081 8303 13093
rect 7303 12960 7337 13081
rect 6792 12940 7337 12960
rect 7495 12940 7529 13081
rect 7687 12940 7721 13081
rect 7879 12940 7913 13081
rect 8071 12940 8105 13081
rect 8263 12954 8297 13081
rect 8413 12957 8447 13503
rect 8214 12940 8224 12954
rect 6792 12906 8224 12940
rect 6792 12896 7337 12906
rect 6792 12852 6999 12896
rect 7303 12775 7337 12896
rect 7495 12775 7529 12906
rect 7687 12775 7721 12906
rect 7879 12775 7913 12906
rect 8071 12775 8105 12906
rect 8214 12890 8224 12906
rect 8288 12890 8298 12954
rect 8413 12950 10684 12957
rect 8413 12893 10637 12950
rect 8263 12775 8297 12890
rect 7297 12763 7343 12775
rect 7297 12683 7303 12763
rect 7337 12683 7343 12763
rect 7297 12671 7343 12683
rect 7393 12763 7439 12775
rect 7393 12683 7399 12763
rect 7433 12683 7439 12763
rect 7393 12671 7439 12683
rect 7489 12763 7535 12775
rect 7489 12683 7495 12763
rect 7529 12683 7535 12763
rect 7489 12671 7535 12683
rect 7585 12763 7631 12775
rect 7585 12683 7591 12763
rect 7625 12683 7631 12763
rect 7585 12671 7631 12683
rect 7681 12763 7727 12775
rect 7681 12683 7687 12763
rect 7721 12683 7727 12763
rect 7681 12671 7727 12683
rect 7777 12763 7823 12775
rect 7777 12683 7783 12763
rect 7817 12683 7823 12763
rect 7777 12671 7823 12683
rect 7873 12763 7919 12775
rect 7873 12683 7879 12763
rect 7913 12683 7919 12763
rect 7873 12671 7919 12683
rect 7969 12763 8015 12775
rect 7969 12683 7975 12763
rect 8009 12683 8015 12763
rect 7969 12671 8015 12683
rect 8065 12763 8111 12775
rect 8065 12683 8071 12763
rect 8105 12683 8111 12763
rect 8065 12671 8111 12683
rect 8161 12763 8207 12775
rect 8161 12683 8167 12763
rect 8201 12683 8207 12763
rect 8161 12671 8207 12683
rect 8257 12763 8303 12775
rect 8257 12683 8263 12763
rect 8297 12683 8303 12763
rect 8257 12671 8303 12683
rect 7277 12576 7287 12640
rect 7351 12576 7361 12640
rect 7399 12529 7433 12671
rect 7591 12529 7625 12671
rect 7783 12529 7817 12671
rect 7975 12529 8009 12671
rect 8167 12529 8201 12671
rect 8243 12578 8253 12642
rect 8317 12578 8327 12642
rect 8413 12529 8447 12893
rect 10627 12886 10637 12893
rect 10701 12886 10711 12950
rect 14379 12882 14442 14744
rect 15945 14301 16009 14985
rect 20227 14893 20233 15141
rect 20267 14893 20273 15141
rect 20227 14881 20273 14893
rect 20323 15141 20369 15153
rect 20323 14893 20329 15141
rect 20363 14893 20369 15141
rect 20323 14881 20369 14893
rect 20419 15141 20465 15153
rect 20419 14893 20425 15141
rect 20459 14893 20465 15141
rect 20419 14881 20465 14893
rect 20515 15141 20561 15153
rect 20515 14893 20521 15141
rect 20555 14893 20561 15141
rect 20515 14881 20561 14893
rect 20611 15141 20657 15153
rect 20611 14893 20617 15141
rect 20651 14893 20657 15141
rect 20611 14881 20657 14893
rect 20707 15141 20753 15153
rect 20707 14893 20713 15141
rect 20747 14893 20753 15141
rect 20707 14881 20753 14893
rect 20803 15141 20849 15153
rect 20803 14893 20809 15141
rect 20843 14893 20849 15141
rect 20803 14881 20849 14893
rect 20899 15141 20945 15153
rect 20899 14893 20905 15141
rect 20939 14893 20945 15141
rect 20899 14881 20945 14893
rect 20995 15141 21041 15153
rect 20995 14893 21001 15141
rect 21035 14893 21041 15141
rect 20995 14881 21041 14893
rect 21091 15141 21137 15153
rect 21091 14893 21097 15141
rect 21131 14893 21137 15141
rect 21091 14881 21137 14893
rect 21187 15141 21233 15153
rect 21187 14893 21193 15141
rect 21227 14893 21233 15141
rect 21187 14881 21233 14893
rect 20233 14754 20267 14881
rect 17820 14690 17830 14754
rect 17894 14740 20267 14754
rect 20425 14740 20459 14881
rect 20617 14740 20651 14881
rect 20809 14740 20843 14881
rect 21001 14740 21035 14881
rect 21193 14740 21227 14881
rect 17894 14706 21227 14740
rect 17894 14690 20267 14706
rect 20233 14575 20267 14690
rect 20425 14575 20459 14706
rect 20617 14575 20651 14706
rect 20809 14575 20843 14706
rect 21001 14575 21035 14706
rect 21193 14575 21227 14706
rect 21343 14818 21377 15303
rect 21844 14818 22051 16417
rect 21343 14611 22051 14818
rect 20227 14563 20273 14575
rect 20227 14483 20233 14563
rect 20267 14483 20273 14563
rect 20227 14471 20273 14483
rect 20323 14563 20369 14575
rect 20323 14483 20329 14563
rect 20363 14483 20369 14563
rect 20323 14471 20369 14483
rect 20419 14563 20465 14575
rect 20419 14483 20425 14563
rect 20459 14483 20465 14563
rect 20419 14471 20465 14483
rect 20515 14563 20561 14575
rect 20515 14483 20521 14563
rect 20555 14483 20561 14563
rect 20515 14471 20561 14483
rect 20611 14563 20657 14575
rect 20611 14483 20617 14563
rect 20651 14483 20657 14563
rect 20611 14471 20657 14483
rect 20707 14563 20753 14575
rect 20707 14483 20713 14563
rect 20747 14483 20753 14563
rect 20707 14471 20753 14483
rect 20803 14563 20849 14575
rect 20803 14483 20809 14563
rect 20843 14483 20849 14563
rect 20803 14471 20849 14483
rect 20899 14563 20945 14575
rect 20899 14483 20905 14563
rect 20939 14483 20945 14563
rect 20899 14471 20945 14483
rect 20995 14563 21041 14575
rect 20995 14483 21001 14563
rect 21035 14483 21041 14563
rect 20995 14471 21041 14483
rect 21091 14563 21137 14575
rect 21091 14483 21097 14563
rect 21131 14483 21137 14563
rect 21091 14471 21137 14483
rect 21187 14563 21233 14575
rect 21187 14483 21193 14563
rect 21227 14483 21233 14563
rect 21187 14471 21233 14483
rect 20207 14373 20217 14437
rect 20281 14373 20291 14437
rect 20329 14329 20363 14471
rect 20521 14329 20555 14471
rect 20713 14329 20747 14471
rect 20905 14329 20939 14471
rect 21097 14329 21131 14471
rect 21170 14378 21180 14442
rect 21244 14378 21254 14442
rect 21343 14329 21377 14611
rect 15935 14237 15945 14301
rect 16009 14237 16019 14301
rect 20329 14295 21377 14329
rect 20329 13503 21377 13537
rect 20208 13386 20218 13450
rect 20282 13386 20292 13450
rect 20329 13353 20363 13503
rect 20521 13353 20555 13503
rect 20713 13353 20747 13503
rect 20905 13353 20939 13503
rect 21097 13353 21131 13503
rect 21168 13386 21178 13450
rect 21242 13386 21252 13450
rect 20227 13341 20273 13353
rect 20227 13093 20233 13341
rect 20267 13093 20273 13341
rect 20227 13081 20273 13093
rect 20323 13341 20369 13353
rect 20323 13093 20329 13341
rect 20363 13093 20369 13341
rect 20323 13081 20369 13093
rect 20419 13341 20465 13353
rect 20419 13093 20425 13341
rect 20459 13093 20465 13341
rect 20419 13081 20465 13093
rect 20515 13341 20561 13353
rect 20515 13093 20521 13341
rect 20555 13093 20561 13341
rect 20515 13081 20561 13093
rect 20611 13341 20657 13353
rect 20611 13093 20617 13341
rect 20651 13093 20657 13341
rect 20611 13081 20657 13093
rect 20707 13341 20753 13353
rect 20707 13093 20713 13341
rect 20747 13093 20753 13341
rect 20707 13081 20753 13093
rect 20803 13341 20849 13353
rect 20803 13093 20809 13341
rect 20843 13093 20849 13341
rect 20803 13081 20849 13093
rect 20899 13341 20945 13353
rect 20899 13093 20905 13341
rect 20939 13093 20945 13341
rect 20899 13081 20945 13093
rect 20995 13341 21041 13353
rect 20995 13093 21001 13341
rect 21035 13093 21041 13341
rect 20995 13081 21041 13093
rect 21091 13341 21137 13353
rect 21091 13093 21097 13341
rect 21131 13093 21137 13341
rect 21091 13081 21137 13093
rect 21187 13341 21233 13353
rect 21187 13093 21193 13341
rect 21227 13093 21233 13341
rect 21187 13081 21233 13093
rect 20233 12956 20267 13081
rect 17825 12892 17835 12956
rect 17899 12940 20267 12956
rect 20425 12940 20459 13081
rect 20617 12940 20651 13081
rect 20809 12940 20843 13081
rect 21001 12940 21035 13081
rect 21193 12940 21227 13081
rect 17899 12906 21227 12940
rect 17899 12892 20267 12906
rect 14369 12818 14379 12882
rect 14443 12818 14453 12882
rect 20233 12775 20267 12892
rect 20425 12775 20459 12906
rect 20617 12775 20651 12906
rect 20809 12775 20843 12906
rect 21001 12775 21035 12906
rect 21193 12775 21227 12906
rect 21343 13014 21377 13503
rect 21844 13014 22051 14611
rect 21343 12807 22051 13014
rect 20227 12763 20273 12775
rect 20227 12683 20233 12763
rect 20267 12683 20273 12763
rect 20227 12671 20273 12683
rect 20323 12763 20369 12775
rect 20323 12683 20329 12763
rect 20363 12683 20369 12763
rect 20323 12671 20369 12683
rect 20419 12763 20465 12775
rect 20419 12683 20425 12763
rect 20459 12683 20465 12763
rect 20419 12671 20465 12683
rect 20515 12763 20561 12775
rect 20515 12683 20521 12763
rect 20555 12683 20561 12763
rect 20515 12671 20561 12683
rect 20611 12763 20657 12775
rect 20611 12683 20617 12763
rect 20651 12683 20657 12763
rect 20611 12671 20657 12683
rect 20707 12763 20753 12775
rect 20707 12683 20713 12763
rect 20747 12683 20753 12763
rect 20707 12671 20753 12683
rect 20803 12763 20849 12775
rect 20803 12683 20809 12763
rect 20843 12683 20849 12763
rect 20803 12671 20849 12683
rect 20899 12763 20945 12775
rect 20899 12683 20905 12763
rect 20939 12683 20945 12763
rect 20899 12671 20945 12683
rect 20995 12763 21041 12775
rect 20995 12683 21001 12763
rect 21035 12683 21041 12763
rect 20995 12671 21041 12683
rect 21091 12763 21137 12775
rect 21091 12683 21097 12763
rect 21131 12683 21137 12763
rect 21091 12671 21137 12683
rect 21187 12763 21233 12775
rect 21187 12683 21193 12763
rect 21227 12683 21233 12763
rect 21187 12671 21233 12683
rect 20205 12572 20215 12636
rect 20279 12572 20289 12636
rect 7399 12495 8447 12529
rect 20329 12529 20363 12671
rect 20521 12529 20555 12671
rect 20713 12529 20747 12671
rect 20905 12529 20939 12671
rect 21097 12529 21131 12671
rect 21170 12574 21180 12638
rect 21244 12574 21254 12638
rect 21343 12529 21377 12807
rect 20329 12495 21377 12529
rect 10707 12235 13401 12299
rect 13465 12235 13475 12299
rect 7399 11703 8447 11737
rect 6307 11514 6348 11637
rect 6458 11514 6514 11637
rect 7277 11587 7287 11651
rect 7351 11587 7361 11651
rect 7399 11553 7433 11703
rect 7591 11553 7625 11703
rect 7783 11553 7817 11703
rect 7975 11553 8009 11703
rect 8167 11553 8201 11703
rect 8240 11587 8250 11651
rect 8314 11587 8324 11651
rect 7297 11541 7343 11553
rect 6307 11102 6335 11514
rect 6747 11236 6753 11514
rect 7297 11293 7303 11541
rect 7337 11293 7343 11541
rect 7297 11281 7343 11293
rect 7393 11541 7439 11553
rect 7393 11293 7399 11541
rect 7433 11293 7439 11541
rect 7393 11281 7439 11293
rect 7489 11541 7535 11553
rect 7489 11293 7495 11541
rect 7529 11293 7535 11541
rect 7489 11281 7535 11293
rect 7585 11541 7631 11553
rect 7585 11293 7591 11541
rect 7625 11293 7631 11541
rect 7585 11281 7631 11293
rect 7681 11541 7727 11553
rect 7681 11293 7687 11541
rect 7721 11293 7727 11541
rect 7681 11281 7727 11293
rect 7777 11541 7823 11553
rect 7777 11293 7783 11541
rect 7817 11293 7823 11541
rect 7777 11281 7823 11293
rect 7873 11541 7919 11553
rect 7873 11293 7879 11541
rect 7913 11293 7919 11541
rect 7873 11281 7919 11293
rect 7969 11541 8015 11553
rect 7969 11293 7975 11541
rect 8009 11293 8015 11541
rect 7969 11281 8015 11293
rect 8065 11541 8111 11553
rect 8065 11293 8071 11541
rect 8105 11293 8111 11541
rect 8065 11281 8111 11293
rect 8161 11541 8207 11553
rect 8161 11293 8167 11541
rect 8201 11293 8207 11541
rect 8161 11281 8207 11293
rect 8257 11541 8303 11553
rect 8257 11293 8263 11541
rect 8297 11293 8303 11541
rect 8257 11281 8303 11293
rect 6747 11156 6956 11236
rect 7303 11156 7337 11281
rect 6747 11140 7337 11156
rect 7495 11140 7529 11281
rect 7687 11140 7721 11281
rect 7879 11140 7913 11281
rect 8071 11140 8105 11281
rect 8263 11156 8297 11281
rect 8221 11140 8231 11156
rect 6747 11106 8231 11140
rect 6747 11102 7337 11106
rect 6307 11097 6348 11102
rect 6458 11097 7337 11102
rect 6307 11092 7337 11097
rect 6307 11029 6956 11092
rect 7303 10975 7337 11092
rect 7495 10975 7529 11106
rect 7687 10975 7721 11106
rect 7879 10975 7913 11106
rect 8071 10975 8105 11106
rect 8221 11092 8231 11106
rect 8295 11092 8305 11156
rect 8413 11153 8447 11703
rect 10707 11153 10771 12235
rect 14663 12121 14673 12185
rect 14737 12121 17223 12185
rect 17287 12121 17297 12185
rect 11231 11936 11241 12000
rect 11305 11936 15397 12000
rect 15461 11936 15471 12000
rect 20329 11703 21377 11737
rect 20207 11585 20217 11649
rect 20281 11585 20291 11649
rect 20329 11553 20363 11703
rect 20521 11553 20555 11703
rect 20713 11553 20747 11703
rect 20905 11553 20939 11703
rect 21097 11553 21131 11703
rect 21172 11586 21182 11650
rect 21246 11586 21256 11650
rect 20227 11541 20273 11553
rect 20227 11293 20233 11541
rect 20267 11293 20273 11541
rect 20227 11281 20273 11293
rect 20323 11541 20369 11553
rect 20323 11293 20329 11541
rect 20363 11293 20369 11541
rect 20323 11281 20369 11293
rect 20419 11541 20465 11553
rect 20419 11293 20425 11541
rect 20459 11293 20465 11541
rect 20419 11281 20465 11293
rect 20515 11541 20561 11553
rect 20515 11293 20521 11541
rect 20555 11293 20561 11541
rect 20515 11281 20561 11293
rect 20611 11541 20657 11553
rect 20611 11293 20617 11541
rect 20651 11293 20657 11541
rect 20611 11281 20657 11293
rect 20707 11541 20753 11553
rect 20707 11293 20713 11541
rect 20747 11293 20753 11541
rect 20707 11281 20753 11293
rect 20803 11541 20849 11553
rect 20803 11293 20809 11541
rect 20843 11293 20849 11541
rect 20803 11281 20849 11293
rect 20899 11541 20945 11553
rect 20899 11293 20905 11541
rect 20939 11293 20945 11541
rect 20899 11281 20945 11293
rect 20995 11541 21041 11553
rect 20995 11293 21001 11541
rect 21035 11293 21041 11541
rect 20995 11281 21041 11293
rect 21091 11541 21137 11553
rect 21091 11293 21097 11541
rect 21131 11293 21137 11541
rect 21091 11281 21137 11293
rect 21187 11541 21233 11553
rect 21187 11293 21193 11541
rect 21227 11293 21233 11541
rect 21187 11281 21233 11293
rect 20233 11156 20267 11281
rect 8263 10975 8297 11092
rect 8413 11089 10772 11153
rect 17793 11152 20267 11156
rect 7297 10963 7343 10975
rect 7297 10883 7303 10963
rect 7337 10883 7343 10963
rect 7297 10871 7343 10883
rect 7393 10963 7439 10975
rect 7393 10883 7399 10963
rect 7433 10883 7439 10963
rect 7393 10871 7439 10883
rect 7489 10963 7535 10975
rect 7489 10883 7495 10963
rect 7529 10883 7535 10963
rect 7489 10871 7535 10883
rect 7585 10963 7631 10975
rect 7585 10883 7591 10963
rect 7625 10883 7631 10963
rect 7585 10871 7631 10883
rect 7681 10963 7727 10975
rect 7681 10883 7687 10963
rect 7721 10883 7727 10963
rect 7681 10871 7727 10883
rect 7777 10963 7823 10975
rect 7777 10883 7783 10963
rect 7817 10883 7823 10963
rect 7777 10871 7823 10883
rect 7873 10963 7919 10975
rect 7873 10883 7879 10963
rect 7913 10883 7919 10963
rect 7873 10871 7919 10883
rect 7969 10963 8015 10975
rect 7969 10883 7975 10963
rect 8009 10883 8015 10963
rect 7969 10871 8015 10883
rect 8065 10963 8111 10975
rect 8065 10883 8071 10963
rect 8105 10883 8111 10963
rect 8065 10871 8111 10883
rect 8161 10963 8207 10975
rect 8161 10883 8167 10963
rect 8201 10883 8207 10963
rect 8161 10871 8207 10883
rect 8257 10963 8303 10975
rect 8257 10883 8263 10963
rect 8297 10883 8303 10963
rect 8257 10871 8303 10883
rect 7277 10773 7287 10837
rect 7351 10773 7361 10837
rect 7399 10729 7433 10871
rect 7591 10729 7625 10871
rect 7783 10729 7817 10871
rect 7975 10729 8009 10871
rect 8167 10729 8201 10871
rect 8240 10777 8250 10841
rect 8314 10777 8324 10841
rect 8413 10729 8447 11089
rect 17761 11088 17771 11152
rect 17835 11140 20267 11152
rect 20425 11140 20459 11281
rect 20617 11140 20651 11281
rect 20809 11140 20843 11281
rect 21001 11140 21035 11281
rect 21193 11140 21227 11281
rect 17835 11106 21227 11140
rect 17835 11092 20267 11106
rect 17835 11088 17845 11092
rect 20233 10975 20267 11092
rect 20425 10975 20459 11106
rect 20617 10975 20651 11106
rect 20809 10975 20843 11106
rect 21001 10975 21035 11106
rect 21193 10975 21227 11106
rect 21343 11261 21377 11703
rect 21844 11732 22051 12807
rect 21844 11261 21885 11732
rect 21996 11539 22051 11732
rect 21997 11429 22051 11539
rect 21343 11225 21885 11261
rect 21996 11225 22051 11429
rect 21343 11054 22051 11225
rect 20227 10963 20273 10975
rect 20227 10883 20233 10963
rect 20267 10883 20273 10963
rect 20227 10871 20273 10883
rect 20323 10963 20369 10975
rect 20323 10883 20329 10963
rect 20363 10883 20369 10963
rect 20323 10871 20369 10883
rect 20419 10963 20465 10975
rect 20419 10883 20425 10963
rect 20459 10883 20465 10963
rect 20419 10871 20465 10883
rect 20515 10963 20561 10975
rect 20515 10883 20521 10963
rect 20555 10883 20561 10963
rect 20515 10871 20561 10883
rect 20611 10963 20657 10975
rect 20611 10883 20617 10963
rect 20651 10883 20657 10963
rect 20611 10871 20657 10883
rect 20707 10963 20753 10975
rect 20707 10883 20713 10963
rect 20747 10883 20753 10963
rect 20707 10871 20753 10883
rect 20803 10963 20849 10975
rect 20803 10883 20809 10963
rect 20843 10883 20849 10963
rect 20803 10871 20849 10883
rect 20899 10963 20945 10975
rect 20899 10883 20905 10963
rect 20939 10883 20945 10963
rect 20899 10871 20945 10883
rect 20995 10963 21041 10975
rect 20995 10883 21001 10963
rect 21035 10883 21041 10963
rect 20995 10871 21041 10883
rect 21091 10963 21137 10975
rect 21091 10883 21097 10963
rect 21131 10883 21137 10963
rect 21091 10871 21137 10883
rect 21187 10963 21233 10975
rect 21187 10883 21193 10963
rect 21227 10883 21233 10963
rect 21187 10871 21233 10883
rect 20207 10774 20217 10838
rect 20281 10774 20291 10838
rect 7399 10695 8447 10729
rect 20329 10729 20363 10871
rect 20521 10729 20555 10871
rect 20713 10729 20747 10871
rect 20905 10729 20939 10871
rect 21097 10729 21131 10871
rect 21169 10775 21179 10839
rect 21243 10775 21253 10839
rect 21343 10729 21377 11054
rect 20329 10695 21377 10729
rect 7399 9903 8447 9937
rect 7277 9787 7287 9851
rect 7351 9787 7361 9851
rect 7399 9753 7433 9903
rect 7591 9753 7625 9903
rect 7783 9753 7817 9903
rect 7975 9753 8009 9903
rect 8167 9753 8201 9903
rect 8238 9788 8248 9852
rect 8312 9788 8322 9852
rect 7297 9741 7343 9753
rect 7297 9493 7303 9741
rect 7337 9493 7343 9741
rect 7297 9481 7343 9493
rect 7393 9741 7439 9753
rect 7393 9493 7399 9741
rect 7433 9493 7439 9741
rect 7393 9481 7439 9493
rect 7489 9741 7535 9753
rect 7489 9493 7495 9741
rect 7529 9493 7535 9741
rect 7489 9481 7535 9493
rect 7585 9741 7631 9753
rect 7585 9493 7591 9741
rect 7625 9493 7631 9741
rect 7585 9481 7631 9493
rect 7681 9741 7727 9753
rect 7681 9493 7687 9741
rect 7721 9493 7727 9741
rect 7681 9481 7727 9493
rect 7777 9741 7823 9753
rect 7777 9493 7783 9741
rect 7817 9493 7823 9741
rect 7777 9481 7823 9493
rect 7873 9741 7919 9753
rect 7873 9493 7879 9741
rect 7913 9493 7919 9741
rect 7873 9481 7919 9493
rect 7969 9741 8015 9753
rect 7969 9493 7975 9741
rect 8009 9493 8015 9741
rect 7969 9481 8015 9493
rect 8065 9741 8111 9753
rect 8065 9493 8071 9741
rect 8105 9493 8111 9741
rect 8065 9481 8111 9493
rect 8161 9741 8207 9753
rect 8161 9493 8167 9741
rect 8201 9493 8207 9741
rect 8161 9481 8207 9493
rect 8257 9741 8303 9753
rect 8257 9493 8263 9741
rect 8297 9493 8303 9741
rect 8257 9481 8303 9493
rect 5695 9358 6958 9392
rect 7303 9358 7337 9481
rect 5695 9340 7337 9358
rect 7495 9340 7529 9481
rect 7687 9340 7721 9481
rect 7879 9340 7913 9481
rect 8071 9340 8105 9481
rect 8263 9355 8297 9481
rect 8413 9357 8447 9903
rect 20329 9903 21377 9937
rect 20209 9786 20219 9850
rect 20283 9786 20293 9850
rect 20329 9753 20363 9903
rect 20521 9753 20555 9903
rect 20713 9753 20747 9903
rect 20905 9753 20939 9903
rect 21097 9753 21131 9903
rect 21169 9786 21179 9850
rect 21243 9786 21253 9850
rect 20227 9741 20273 9753
rect 20227 9493 20233 9741
rect 20267 9493 20273 9741
rect 20227 9481 20273 9493
rect 20323 9741 20369 9753
rect 20323 9493 20329 9741
rect 20363 9493 20369 9741
rect 20323 9481 20369 9493
rect 20419 9741 20465 9753
rect 20419 9493 20425 9741
rect 20459 9493 20465 9741
rect 20419 9481 20465 9493
rect 20515 9741 20561 9753
rect 20515 9493 20521 9741
rect 20555 9493 20561 9741
rect 20515 9481 20561 9493
rect 20611 9741 20657 9753
rect 20611 9493 20617 9741
rect 20651 9493 20657 9741
rect 20611 9481 20657 9493
rect 20707 9741 20753 9753
rect 20707 9493 20713 9741
rect 20747 9493 20753 9741
rect 20707 9481 20753 9493
rect 20803 9741 20849 9753
rect 20803 9493 20809 9741
rect 20843 9493 20849 9741
rect 20803 9481 20849 9493
rect 20899 9741 20945 9753
rect 20899 9493 20905 9741
rect 20939 9493 20945 9741
rect 20899 9481 20945 9493
rect 20995 9741 21041 9753
rect 20995 9493 21001 9741
rect 21035 9493 21041 9741
rect 20995 9481 21041 9493
rect 21091 9741 21137 9753
rect 21091 9493 21097 9741
rect 21131 9493 21137 9741
rect 21091 9481 21137 9493
rect 21187 9741 21233 9753
rect 21187 9493 21193 9741
rect 21227 9493 21233 9741
rect 21187 9481 21233 9493
rect 10559 9357 10569 9358
rect 8222 9340 8232 9355
rect 5695 9306 8232 9340
rect 5695 9294 7337 9306
rect 5695 9185 6958 9294
rect 7303 9175 7337 9294
rect 7495 9175 7529 9306
rect 7687 9175 7721 9306
rect 7879 9175 7913 9306
rect 8071 9175 8105 9306
rect 8222 9291 8232 9306
rect 8296 9291 8306 9355
rect 8413 9294 10569 9357
rect 10633 9294 10643 9358
rect 17779 9296 17789 9360
rect 17853 9359 17863 9360
rect 20233 9359 20267 9481
rect 17853 9340 20267 9359
rect 20425 9340 20459 9481
rect 20617 9340 20651 9481
rect 20809 9340 20843 9481
rect 21001 9340 21035 9481
rect 21193 9340 21227 9481
rect 17853 9306 21227 9340
rect 17853 9296 20267 9306
rect 17838 9295 20267 9296
rect 8413 9293 10631 9294
rect 8263 9175 8297 9291
rect 7297 9163 7343 9175
rect 7297 9083 7303 9163
rect 7337 9083 7343 9163
rect 7297 9071 7343 9083
rect 7393 9163 7439 9175
rect 7393 9083 7399 9163
rect 7433 9083 7439 9163
rect 7393 9071 7439 9083
rect 7489 9163 7535 9175
rect 7489 9083 7495 9163
rect 7529 9083 7535 9163
rect 7489 9071 7535 9083
rect 7585 9163 7631 9175
rect 7585 9083 7591 9163
rect 7625 9083 7631 9163
rect 7585 9071 7631 9083
rect 7681 9163 7727 9175
rect 7681 9083 7687 9163
rect 7721 9083 7727 9163
rect 7681 9071 7727 9083
rect 7777 9163 7823 9175
rect 7777 9083 7783 9163
rect 7817 9083 7823 9163
rect 7777 9071 7823 9083
rect 7873 9163 7919 9175
rect 7873 9083 7879 9163
rect 7913 9083 7919 9163
rect 7873 9071 7919 9083
rect 7969 9163 8015 9175
rect 7969 9083 7975 9163
rect 8009 9083 8015 9163
rect 7969 9071 8015 9083
rect 8065 9163 8111 9175
rect 8065 9083 8071 9163
rect 8105 9083 8111 9163
rect 8065 9071 8111 9083
rect 8161 9163 8207 9175
rect 8161 9083 8167 9163
rect 8201 9083 8207 9163
rect 8161 9071 8207 9083
rect 8257 9163 8303 9175
rect 8257 9083 8263 9163
rect 8297 9083 8303 9163
rect 8257 9071 8303 9083
rect 7280 8973 7290 9037
rect 7354 8973 7364 9037
rect 7399 8929 7433 9071
rect 7591 8929 7625 9071
rect 7783 8929 7817 9071
rect 7975 8929 8009 9071
rect 8167 8929 8201 9071
rect 8237 8975 8247 9039
rect 8311 8975 8321 9039
rect 8413 8929 8447 9293
rect 20233 9175 20267 9295
rect 20425 9175 20459 9306
rect 20617 9175 20651 9306
rect 20809 9175 20843 9306
rect 21001 9175 21035 9306
rect 21193 9175 21227 9306
rect 21343 9462 21377 9903
rect 22410 9835 22617 18220
rect 22389 9462 22399 9835
rect 21343 9295 22399 9462
rect 22509 9295 22617 9835
rect 21343 9255 22617 9295
rect 20227 9163 20273 9175
rect 20227 9083 20233 9163
rect 20267 9083 20273 9163
rect 20227 9071 20273 9083
rect 20323 9163 20369 9175
rect 20323 9083 20329 9163
rect 20363 9083 20369 9163
rect 20323 9071 20369 9083
rect 20419 9163 20465 9175
rect 20419 9083 20425 9163
rect 20459 9083 20465 9163
rect 20419 9071 20465 9083
rect 20515 9163 20561 9175
rect 20515 9083 20521 9163
rect 20555 9083 20561 9163
rect 20515 9071 20561 9083
rect 20611 9163 20657 9175
rect 20611 9083 20617 9163
rect 20651 9083 20657 9163
rect 20611 9071 20657 9083
rect 20707 9163 20753 9175
rect 20707 9083 20713 9163
rect 20747 9083 20753 9163
rect 20707 9071 20753 9083
rect 20803 9163 20849 9175
rect 20803 9083 20809 9163
rect 20843 9083 20849 9163
rect 20803 9071 20849 9083
rect 20899 9163 20945 9175
rect 20899 9083 20905 9163
rect 20939 9083 20945 9163
rect 20899 9071 20945 9083
rect 20995 9163 21041 9175
rect 20995 9083 21001 9163
rect 21035 9083 21041 9163
rect 20995 9071 21041 9083
rect 21091 9163 21137 9175
rect 21091 9083 21097 9163
rect 21131 9083 21137 9163
rect 21091 9071 21137 9083
rect 21187 9163 21233 9175
rect 21187 9083 21193 9163
rect 21227 9083 21233 9163
rect 21187 9071 21233 9083
rect 7399 8895 8447 8929
rect 8703 9017 8983 9023
rect 8703 8761 8715 9017
rect 8971 8761 8983 9017
rect 8703 8755 8983 8761
rect 19638 9005 19918 9011
rect 8715 8582 8971 8755
rect 19638 8749 19650 9005
rect 19906 8749 19918 9005
rect 20206 8976 20216 9040
rect 20280 8976 20290 9040
rect 20329 8929 20363 9071
rect 20521 8929 20555 9071
rect 20713 8929 20747 9071
rect 20905 8929 20939 9071
rect 21097 8929 21131 9071
rect 21171 8975 21181 9039
rect 21245 8975 21255 9039
rect 21343 8929 21377 9255
rect 20329 8895 21377 8929
rect 19638 8743 19918 8749
rect 5543 8576 8971 8582
rect 5543 8332 5555 8576
rect 5799 8332 8971 8576
rect 5543 8326 8971 8332
rect 19650 8575 19906 8743
rect 19650 8569 23753 8575
rect 19650 8325 23497 8569
rect 23741 8325 23753 8569
rect 19650 8319 23753 8325
rect 7238 7007 22063 7047
rect 7238 7005 12010 7007
rect 7238 7002 9324 7005
rect 7238 6991 8256 7002
rect 8314 6991 9324 7002
rect 9382 7002 12010 7005
rect 9382 6991 10942 7002
rect 11000 6991 12010 7002
rect 12068 6991 22063 7007
rect 7238 6957 7445 6991
rect 14299 6957 14467 6991
rect 20872 6957 22063 6991
rect 7238 6944 8256 6957
rect 8314 6947 9324 6957
rect 9382 6947 10942 6957
rect 8314 6944 10942 6947
rect 11000 6949 12010 6957
rect 12068 6949 22063 6957
rect 11000 6944 22063 6949
rect 7238 6919 22063 6944
rect 15050 6813 15798 6919
rect 14942 6759 15018 6765
rect 14942 6725 14954 6759
rect 15006 6725 15018 6759
rect 14942 6719 15018 6725
rect 7802 6690 7878 6696
rect 7802 6656 7814 6690
rect 7866 6656 7878 6690
rect 7802 6650 7878 6656
rect 7980 6690 8056 6696
rect 7980 6656 7992 6690
rect 8044 6656 8056 6690
rect 7980 6650 8056 6656
rect 8158 6690 8234 6696
rect 8158 6656 8170 6690
rect 8222 6656 8234 6690
rect 8158 6650 8234 6656
rect 8336 6690 8412 6696
rect 8336 6656 8348 6690
rect 8400 6656 8412 6690
rect 8336 6650 8412 6656
rect 8514 6690 8590 6696
rect 8514 6656 8526 6690
rect 8578 6656 8590 6690
rect 8514 6650 8590 6656
rect 8692 6690 8768 6696
rect 8692 6656 8704 6690
rect 8756 6656 8768 6690
rect 8692 6650 8768 6656
rect 8870 6690 8946 6696
rect 8870 6656 8882 6690
rect 8934 6656 8946 6690
rect 8870 6650 8946 6656
rect 9048 6690 9124 6696
rect 9048 6656 9060 6690
rect 9112 6656 9124 6690
rect 9048 6650 9124 6656
rect 9226 6690 9302 6696
rect 9226 6656 9238 6690
rect 9290 6656 9302 6690
rect 9226 6650 9302 6656
rect 9404 6690 9480 6696
rect 9404 6656 9416 6690
rect 9468 6656 9480 6690
rect 9404 6650 9480 6656
rect 9582 6690 9658 6696
rect 9582 6656 9594 6690
rect 9646 6656 9658 6690
rect 9582 6650 9658 6656
rect 9760 6690 9836 6696
rect 9760 6656 9772 6690
rect 9824 6656 9836 6690
rect 9760 6650 9836 6656
rect 10488 6690 10564 6696
rect 10488 6656 10500 6690
rect 10552 6656 10564 6690
rect 10488 6650 10564 6656
rect 10666 6690 10742 6696
rect 10666 6656 10678 6690
rect 10730 6656 10742 6690
rect 10666 6650 10742 6656
rect 10844 6690 10920 6696
rect 10844 6656 10856 6690
rect 10908 6656 10920 6690
rect 10844 6650 10920 6656
rect 11022 6690 11098 6696
rect 11022 6656 11034 6690
rect 11086 6656 11098 6690
rect 11022 6650 11098 6656
rect 11200 6690 11276 6696
rect 11200 6656 11212 6690
rect 11264 6656 11276 6690
rect 11200 6650 11276 6656
rect 11378 6690 11454 6696
rect 11378 6656 11390 6690
rect 11442 6656 11454 6690
rect 11378 6650 11454 6656
rect 11556 6690 11632 6696
rect 11556 6656 11568 6690
rect 11620 6656 11632 6690
rect 11556 6650 11632 6656
rect 11734 6690 11810 6696
rect 11734 6656 11746 6690
rect 11798 6656 11810 6690
rect 11734 6650 11810 6656
rect 11912 6690 11988 6696
rect 11912 6656 11924 6690
rect 11976 6656 11988 6690
rect 11912 6650 11988 6656
rect 12090 6690 12166 6696
rect 12090 6656 12102 6690
rect 12154 6656 12166 6690
rect 12090 6650 12166 6656
rect 12268 6690 12344 6696
rect 12268 6656 12280 6690
rect 12332 6656 12344 6690
rect 12268 6650 12344 6656
rect 12446 6690 12522 6696
rect 12446 6656 12458 6690
rect 12510 6656 12522 6690
rect 15051 6678 15086 6813
rect 15120 6759 15196 6765
rect 15120 6725 15132 6759
rect 15184 6725 15196 6759
rect 15120 6719 15196 6725
rect 15298 6759 15374 6765
rect 15298 6725 15310 6759
rect 15362 6725 15374 6759
rect 15298 6719 15374 6725
rect 15407 6678 15442 6813
rect 15476 6759 15552 6765
rect 15476 6725 15488 6759
rect 15540 6725 15552 6759
rect 15476 6719 15552 6725
rect 15654 6759 15730 6765
rect 15654 6725 15666 6759
rect 15718 6725 15730 6759
rect 15654 6719 15730 6725
rect 15763 6678 15798 6813
rect 17251 6803 17999 6919
rect 15832 6759 15908 6765
rect 15832 6725 15844 6759
rect 15896 6725 15908 6759
rect 15832 6719 15908 6725
rect 17142 6759 17218 6765
rect 17142 6725 17154 6759
rect 17206 6725 17218 6759
rect 17142 6719 17218 6725
rect 17251 6678 17286 6803
rect 17320 6759 17396 6765
rect 17320 6725 17332 6759
rect 17384 6725 17396 6759
rect 17320 6719 17396 6725
rect 17498 6759 17574 6765
rect 17498 6725 17510 6759
rect 17562 6725 17574 6759
rect 17498 6719 17574 6725
rect 17608 6678 17643 6803
rect 17676 6759 17752 6765
rect 17676 6725 17688 6759
rect 17740 6725 17752 6759
rect 17676 6719 17752 6725
rect 17854 6759 17930 6765
rect 17854 6725 17866 6759
rect 17918 6725 17930 6759
rect 17854 6719 17930 6725
rect 17964 6678 17999 6803
rect 19451 6839 20199 6919
rect 19451 6804 20198 6839
rect 18032 6759 18108 6765
rect 18032 6725 18044 6759
rect 18096 6725 18108 6759
rect 18032 6719 18108 6725
rect 19342 6759 19418 6765
rect 19342 6725 19354 6759
rect 19406 6725 19418 6759
rect 19342 6719 19418 6725
rect 19451 6678 19486 6804
rect 19520 6759 19596 6765
rect 19520 6725 19532 6759
rect 19584 6725 19596 6759
rect 19520 6719 19596 6725
rect 19698 6759 19774 6765
rect 19698 6725 19710 6759
rect 19762 6725 19774 6759
rect 19698 6719 19774 6725
rect 19808 6678 19843 6804
rect 19876 6759 19952 6765
rect 19876 6725 19888 6759
rect 19940 6725 19952 6759
rect 19876 6719 19952 6725
rect 20054 6759 20130 6765
rect 20054 6725 20066 6759
rect 20118 6725 20130 6759
rect 20054 6719 20130 6725
rect 20163 6678 20198 6804
rect 20232 6759 20308 6765
rect 20232 6725 20244 6759
rect 20296 6725 20308 6759
rect 20232 6719 20308 6725
rect 14868 6666 14914 6678
rect 15046 6666 15092 6678
rect 15224 6666 15270 6678
rect 15402 6666 15448 6678
rect 15580 6666 15626 6678
rect 15758 6666 15804 6678
rect 15936 6666 15982 6678
rect 17068 6666 17114 6678
rect 17246 6666 17292 6678
rect 17424 6666 17470 6678
rect 17602 6666 17648 6678
rect 17780 6666 17826 6678
rect 17958 6666 18004 6678
rect 18136 6666 18182 6678
rect 19268 6666 19314 6678
rect 19446 6666 19492 6678
rect 19624 6666 19670 6678
rect 19802 6666 19848 6678
rect 19980 6666 20026 6678
rect 20158 6666 20204 6678
rect 20336 6666 20382 6678
rect 12446 6650 12522 6656
rect 14852 6608 14862 6666
rect 14920 6608 14930 6666
rect 12178 6603 12188 6604
rect 7722 6598 9502 6603
rect 7722 6597 8078 6598
rect 8136 6597 9502 6598
rect 9560 6597 9916 6603
rect 7722 6563 7734 6597
rect 7768 6563 8078 6597
rect 8136 6563 8446 6597
rect 8480 6563 8802 6597
rect 8836 6563 9158 6597
rect 9192 6563 9502 6597
rect 9560 6563 9870 6597
rect 9904 6563 9916 6597
rect 7722 6557 8078 6563
rect 8068 6540 8078 6557
rect 8136 6557 9502 6563
rect 8136 6540 8146 6557
rect 9492 6545 9502 6557
rect 9560 6557 9916 6563
rect 10408 6597 12188 6603
rect 12246 6603 12256 6604
rect 12246 6597 12602 6603
rect 10408 6563 10420 6597
rect 10454 6563 10764 6597
rect 10822 6563 11132 6597
rect 11166 6563 11488 6597
rect 11522 6563 11844 6597
rect 11878 6563 12188 6597
rect 12246 6563 12556 6597
rect 12590 6563 12602 6597
rect 10408 6557 10764 6563
rect 9560 6545 9570 6557
rect 10754 6539 10764 6557
rect 10822 6557 12188 6563
rect 10822 6539 10832 6557
rect 12178 6546 12188 6557
rect 12246 6557 12602 6563
rect 12246 6546 12256 6557
rect 14868 6410 14874 6608
rect 14908 6410 14914 6608
rect 15046 6468 15052 6666
rect 15086 6468 15092 6666
rect 15208 6608 15218 6666
rect 15276 6608 15286 6666
rect 15030 6410 15040 6468
rect 15098 6410 15108 6468
rect 15224 6410 15230 6608
rect 15264 6410 15270 6608
rect 15402 6468 15408 6666
rect 15442 6468 15448 6666
rect 15564 6608 15574 6666
rect 15632 6608 15642 6666
rect 15386 6410 15396 6468
rect 15454 6410 15464 6468
rect 15580 6410 15586 6608
rect 15620 6410 15626 6608
rect 15758 6468 15764 6666
rect 15798 6468 15804 6666
rect 15920 6608 15930 6666
rect 15988 6608 15998 6666
rect 17053 6608 17063 6666
rect 17121 6608 17131 6666
rect 15742 6410 15752 6468
rect 15810 6410 15820 6468
rect 15936 6410 15942 6608
rect 15976 6410 15982 6608
rect 14868 6398 14914 6410
rect 15046 6398 15092 6410
rect 15224 6398 15270 6410
rect 15402 6398 15448 6410
rect 15580 6398 15626 6410
rect 15758 6398 15804 6410
rect 15936 6398 15982 6410
rect 17068 6410 17074 6608
rect 17108 6410 17114 6608
rect 17246 6468 17252 6666
rect 17286 6468 17292 6666
rect 17408 6608 17418 6666
rect 17476 6608 17486 6666
rect 17230 6410 17240 6468
rect 17298 6410 17308 6468
rect 17424 6410 17430 6608
rect 17464 6410 17470 6608
rect 17602 6467 17608 6666
rect 17642 6467 17648 6666
rect 17764 6608 17774 6666
rect 17832 6608 17842 6666
rect 17068 6398 17114 6410
rect 17246 6398 17292 6410
rect 17424 6398 17470 6410
rect 17586 6409 17596 6467
rect 17654 6409 17664 6467
rect 17780 6410 17786 6608
rect 17820 6410 17826 6608
rect 17958 6468 17964 6666
rect 17998 6468 18004 6666
rect 18120 6608 18130 6666
rect 18188 6608 18198 6666
rect 19252 6608 19262 6666
rect 19320 6608 19330 6666
rect 17942 6410 17952 6468
rect 18010 6410 18020 6468
rect 18136 6410 18142 6608
rect 18176 6410 18182 6608
rect 17602 6398 17648 6409
rect 17780 6398 17826 6410
rect 17958 6398 18004 6410
rect 18136 6398 18182 6410
rect 19268 6410 19274 6608
rect 19308 6410 19314 6608
rect 19446 6468 19452 6666
rect 19486 6468 19492 6666
rect 19608 6608 19618 6666
rect 19676 6608 19686 6666
rect 19430 6410 19440 6468
rect 19498 6410 19508 6468
rect 19624 6410 19630 6608
rect 19664 6410 19670 6608
rect 19802 6468 19808 6666
rect 19842 6468 19848 6666
rect 19964 6608 19974 6666
rect 20032 6608 20042 6666
rect 19786 6410 19796 6468
rect 19854 6410 19864 6468
rect 19980 6410 19986 6608
rect 20020 6410 20026 6608
rect 20158 6468 20164 6666
rect 20198 6468 20204 6666
rect 20320 6608 20330 6666
rect 20388 6608 20398 6666
rect 20142 6410 20152 6468
rect 20210 6410 20220 6468
rect 20336 6410 20342 6608
rect 20376 6410 20382 6608
rect 19268 6398 19314 6410
rect 19446 6398 19492 6410
rect 19624 6398 19670 6410
rect 19802 6398 19848 6410
rect 19980 6398 20026 6410
rect 20158 6398 20204 6410
rect 20336 6398 20382 6410
rect 8246 6381 8256 6393
rect 7900 6375 8256 6381
rect 8314 6381 8324 6393
rect 9314 6381 9324 6393
rect 8314 6375 9324 6381
rect 9382 6381 9392 6393
rect 10932 6381 10942 6393
rect 9382 6375 9738 6381
rect 7900 6341 7912 6375
rect 7946 6341 8256 6375
rect 8314 6341 8624 6375
rect 8658 6341 8980 6375
rect 9014 6341 9324 6375
rect 9382 6341 9692 6375
rect 9726 6341 9738 6375
rect 7900 6335 8256 6341
rect 8314 6335 9324 6341
rect 9382 6335 9738 6341
rect 10586 6375 10942 6381
rect 11000 6381 11010 6393
rect 12000 6381 12010 6393
rect 11000 6375 12010 6381
rect 12068 6381 12078 6393
rect 12068 6375 12424 6381
rect 10586 6341 10598 6375
rect 10632 6341 10942 6375
rect 11000 6341 11310 6375
rect 11344 6341 11666 6375
rect 11700 6341 12010 6375
rect 12068 6341 12378 6375
rect 12412 6341 12424 6375
rect 10586 6335 10942 6341
rect 11000 6335 12010 6341
rect 12068 6335 12424 6341
rect 14942 6351 15018 6357
rect 15120 6351 15196 6357
rect 15298 6351 15374 6357
rect 15407 6351 15442 6352
rect 15476 6351 15552 6357
rect 15654 6351 15730 6357
rect 15832 6351 15908 6357
rect 14942 6317 14954 6351
rect 15006 6317 15132 6351
rect 15184 6317 15310 6351
rect 15362 6317 15488 6351
rect 15540 6317 15666 6351
rect 15718 6317 15844 6351
rect 15896 6317 15908 6351
rect 14942 6311 15018 6317
rect 15120 6311 15196 6317
rect 15298 6311 15552 6317
rect 15654 6311 15730 6317
rect 15832 6311 15908 6317
rect 17142 6351 17218 6357
rect 17320 6351 17396 6357
rect 17498 6351 17574 6357
rect 17676 6351 17752 6357
rect 17854 6351 17930 6357
rect 18032 6351 18108 6357
rect 17142 6317 17154 6351
rect 17206 6317 17332 6351
rect 17384 6317 17510 6351
rect 17562 6317 17688 6351
rect 17740 6317 17866 6351
rect 17918 6317 18044 6351
rect 18096 6317 18108 6351
rect 17142 6311 17218 6317
rect 17320 6311 17396 6317
rect 17498 6311 17752 6317
rect 17854 6311 17930 6317
rect 18032 6311 18108 6317
rect 19342 6351 19418 6357
rect 19520 6351 19596 6357
rect 19698 6351 19774 6357
rect 19876 6351 19952 6357
rect 20054 6351 20130 6357
rect 20231 6351 20241 6357
rect 19342 6317 19354 6351
rect 19406 6317 19532 6351
rect 19584 6317 19710 6351
rect 19762 6317 19888 6351
rect 19940 6317 20066 6351
rect 20118 6317 20241 6351
rect 19342 6311 19418 6317
rect 19520 6311 19596 6317
rect 19698 6311 19843 6317
rect 19876 6311 19952 6317
rect 20054 6311 20130 6317
rect 7802 6282 7878 6288
rect 7980 6282 8056 6288
rect 8158 6282 8234 6288
rect 8336 6282 8412 6288
rect 8514 6282 8590 6288
rect 8692 6282 8768 6288
rect 8870 6282 8946 6288
rect 9048 6282 9124 6288
rect 9226 6282 9302 6288
rect 9404 6282 9480 6288
rect 9582 6282 9658 6288
rect 9760 6282 9836 6288
rect 7802 6248 7814 6282
rect 7866 6248 7992 6282
rect 8044 6248 8170 6282
rect 8222 6248 8348 6282
rect 8400 6248 8526 6282
rect 8578 6248 8704 6282
rect 8756 6248 8882 6282
rect 8934 6248 9060 6282
rect 9112 6248 9238 6282
rect 9290 6248 9416 6282
rect 9468 6248 9594 6282
rect 9646 6248 9772 6282
rect 9824 6248 9836 6282
rect 7802 6112 7878 6248
rect 7980 6242 8056 6248
rect 8158 6242 8234 6248
rect 8336 6242 8412 6248
rect 8514 6242 8590 6248
rect 8692 6242 8768 6248
rect 8870 6242 8946 6248
rect 9048 6242 9124 6248
rect 9226 6242 9302 6248
rect 9404 6242 9480 6248
rect 9582 6242 9658 6248
rect 9760 6209 9836 6248
rect 10488 6282 10564 6288
rect 10666 6282 10742 6288
rect 10844 6282 10920 6288
rect 11022 6282 11098 6288
rect 11200 6282 11276 6288
rect 11378 6282 11454 6288
rect 11556 6282 11632 6288
rect 11734 6282 11810 6288
rect 11912 6282 11988 6288
rect 12090 6282 12166 6288
rect 12268 6282 12344 6288
rect 12446 6282 12522 6288
rect 10488 6248 10500 6282
rect 10552 6248 10678 6282
rect 10730 6248 10856 6282
rect 10908 6248 11034 6282
rect 11086 6248 11212 6282
rect 11264 6248 11390 6282
rect 11442 6248 11568 6282
rect 11620 6248 11746 6282
rect 11798 6248 11924 6282
rect 11976 6248 12102 6282
rect 12154 6248 12280 6282
rect 12332 6280 12458 6282
rect 12510 6280 12522 6282
rect 12332 6248 12446 6280
rect 10488 6209 10564 6248
rect 10666 6242 10742 6248
rect 10844 6242 10920 6248
rect 11022 6242 11098 6248
rect 11200 6242 11276 6248
rect 11378 6242 11454 6248
rect 11556 6242 11632 6248
rect 11734 6242 11810 6248
rect 11912 6242 11988 6248
rect 12090 6242 12166 6248
rect 12268 6242 12344 6248
rect 9758 6151 9768 6209
rect 9826 6151 9836 6209
rect 10487 6151 10497 6209
rect 10555 6151 10565 6209
rect 7980 6112 8056 6118
rect 8158 6112 8234 6118
rect 8336 6112 8412 6118
rect 8514 6112 8590 6118
rect 8692 6112 8768 6118
rect 8870 6112 8946 6118
rect 9048 6112 9124 6118
rect 9226 6112 9302 6118
rect 9404 6112 9480 6118
rect 9582 6112 9658 6118
rect 9760 6112 9836 6151
rect 7802 6078 7814 6112
rect 7866 6078 7992 6112
rect 8044 6078 8170 6112
rect 8222 6078 8348 6112
rect 8400 6078 8526 6112
rect 8578 6078 8704 6112
rect 8756 6078 8882 6112
rect 8934 6078 9060 6112
rect 9112 6078 9238 6112
rect 9290 6078 9416 6112
rect 9468 6078 9594 6112
rect 9646 6078 9772 6112
rect 9824 6078 9836 6112
rect 7802 6072 7878 6078
rect 7980 6072 8056 6078
rect 8158 6072 8234 6078
rect 8336 6072 8412 6078
rect 8514 6072 8590 6078
rect 8692 6072 8768 6078
rect 8870 6072 8946 6078
rect 9048 6072 9124 6078
rect 9226 6072 9302 6078
rect 9404 6072 9480 6078
rect 9582 6072 9658 6078
rect 9760 6072 9836 6078
rect 10488 6113 10564 6151
rect 10666 6113 10742 6119
rect 10844 6113 10920 6119
rect 11022 6113 11098 6119
rect 11200 6113 11276 6119
rect 11378 6113 11454 6119
rect 11556 6113 11632 6119
rect 11734 6113 11810 6119
rect 11912 6113 11988 6119
rect 12090 6113 12166 6119
rect 12268 6113 12344 6119
rect 12436 6113 12446 6248
rect 10488 6079 10500 6113
rect 10552 6079 10678 6113
rect 10730 6079 10856 6113
rect 10908 6079 11034 6113
rect 11086 6079 11212 6113
rect 11264 6079 11390 6113
rect 11442 6079 11568 6113
rect 11620 6079 11746 6113
rect 11798 6079 11924 6113
rect 11976 6079 12102 6113
rect 12154 6079 12280 6113
rect 12332 6080 12446 6113
rect 12525 6080 12535 6280
rect 15366 6228 15483 6311
rect 17568 6228 17685 6311
rect 19726 6228 19843 6311
rect 20231 6299 20241 6317
rect 20299 6299 20309 6357
rect 12834 6111 12844 6228
rect 12957 6111 19843 6228
rect 12332 6079 12458 6080
rect 12510 6079 12522 6080
rect 10488 6073 10564 6079
rect 10666 6073 10742 6079
rect 10844 6073 10920 6079
rect 11022 6073 11098 6079
rect 11200 6073 11276 6079
rect 11378 6073 11454 6079
rect 11556 6073 11632 6079
rect 11734 6073 11810 6079
rect 11912 6073 11988 6079
rect 12090 6073 12166 6079
rect 12268 6073 12344 6079
rect 12446 6073 12522 6079
rect 8712 6025 8722 6032
rect 7722 6019 8078 6025
rect 8136 6019 8722 6025
rect 8914 6025 8924 6032
rect 11398 6026 11408 6030
rect 8914 6019 9502 6025
rect 9560 6019 9916 6025
rect 7722 5985 7734 6019
rect 7768 5985 8078 6019
rect 8136 5985 8446 6019
rect 8480 5985 8722 6019
rect 8914 5985 9158 6019
rect 9192 5985 9502 6019
rect 9560 5985 9870 6019
rect 9904 5985 9916 6019
rect 7722 5979 8078 5985
rect 8068 5967 8078 5979
rect 8136 5979 8722 5985
rect 8136 5967 8146 5979
rect 8712 5974 8722 5979
rect 8914 5979 9502 5985
rect 8914 5974 8924 5979
rect 8780 5967 8790 5974
rect 8848 5967 8858 5974
rect 9492 5967 9502 5979
rect 9560 5979 9916 5985
rect 10408 6020 10764 6026
rect 10822 6020 11408 6026
rect 11600 6026 11610 6030
rect 11600 6020 12188 6026
rect 12246 6020 12602 6026
rect 10408 5986 10420 6020
rect 10454 5986 10764 6020
rect 10822 5986 11132 6020
rect 11166 5986 11408 6020
rect 11600 5986 11844 6020
rect 11878 5986 12188 6020
rect 12246 5986 12556 6020
rect 12590 5986 12602 6020
rect 10408 5980 10764 5986
rect 9560 5967 9570 5979
rect 10754 5968 10764 5980
rect 10822 5980 11408 5986
rect 10822 5968 10832 5980
rect 11398 5972 11408 5980
rect 11600 5980 12188 5986
rect 11600 5972 11610 5980
rect 11466 5968 11476 5972
rect 11534 5968 11544 5972
rect 12178 5968 12188 5980
rect 12246 5980 12602 5986
rect 14943 5992 15019 5998
rect 12246 5968 12256 5980
rect 14943 5958 14955 5992
rect 15007 5958 15019 5992
rect 14943 5952 15019 5958
rect 15121 5992 15197 5998
rect 15121 5958 15133 5992
rect 15185 5958 15197 5992
rect 15121 5952 15197 5958
rect 15299 5992 15375 5998
rect 15299 5958 15311 5992
rect 15363 5958 15375 5992
rect 15299 5952 15375 5958
rect 15477 5992 15553 5998
rect 15477 5958 15489 5992
rect 15541 5958 15553 5992
rect 15477 5952 15553 5958
rect 15655 5992 15731 5998
rect 15655 5958 15667 5992
rect 15719 5958 15731 5992
rect 15655 5952 15731 5958
rect 15833 5992 15909 5998
rect 15833 5958 15845 5992
rect 15897 5958 15909 5992
rect 15833 5952 15909 5958
rect 17143 5992 17219 5998
rect 17143 5958 17155 5992
rect 17207 5958 17219 5992
rect 17143 5952 17219 5958
rect 17321 5992 17397 5998
rect 17321 5958 17333 5992
rect 17385 5958 17397 5992
rect 17321 5952 17397 5958
rect 17499 5992 17575 5998
rect 17499 5958 17511 5992
rect 17563 5958 17575 5992
rect 17499 5952 17575 5958
rect 17677 5992 17753 5998
rect 17677 5958 17689 5992
rect 17741 5958 17753 5992
rect 17677 5952 17753 5958
rect 17855 5992 17931 5998
rect 17855 5958 17867 5992
rect 17919 5958 17931 5992
rect 17855 5952 17931 5958
rect 18033 5992 18109 5998
rect 18033 5958 18045 5992
rect 18097 5958 18109 5992
rect 18033 5952 18109 5958
rect 19343 5992 19419 5998
rect 19343 5958 19355 5992
rect 19407 5958 19419 5992
rect 19343 5952 19419 5958
rect 19521 5992 19597 5998
rect 19521 5958 19533 5992
rect 19585 5958 19597 5992
rect 19521 5952 19597 5958
rect 19699 5992 19775 5998
rect 19699 5958 19711 5992
rect 19763 5958 19775 5992
rect 19699 5952 19775 5958
rect 19877 5992 19953 5998
rect 19877 5958 19889 5992
rect 19941 5958 19953 5992
rect 19877 5952 19953 5958
rect 20055 5992 20131 5998
rect 20055 5958 20067 5992
rect 20119 5958 20131 5992
rect 20055 5952 20131 5958
rect 20233 5992 20309 5998
rect 20233 5958 20245 5992
rect 20297 5958 20309 5992
rect 20233 5952 20309 5958
rect 14869 5899 14915 5911
rect 15047 5899 15093 5911
rect 15225 5899 15271 5911
rect 15403 5899 15449 5911
rect 15581 5899 15627 5911
rect 15759 5899 15805 5911
rect 15937 5899 15983 5911
rect 17069 5899 17115 5911
rect 17247 5899 17293 5911
rect 17425 5899 17471 5911
rect 17603 5899 17649 5911
rect 17781 5899 17827 5911
rect 17959 5899 18005 5911
rect 18137 5899 18183 5911
rect 19269 5899 19315 5911
rect 19447 5899 19493 5911
rect 19625 5899 19671 5911
rect 19803 5899 19849 5911
rect 19981 5899 20027 5911
rect 20159 5899 20205 5911
rect 20337 5899 20383 5911
rect 14853 5841 14863 5899
rect 14921 5841 14931 5899
rect 8246 5803 8256 5815
rect 7900 5797 8256 5803
rect 8314 5803 8324 5815
rect 9314 5803 9324 5815
rect 8314 5797 9324 5803
rect 9382 5803 9392 5815
rect 10932 5804 10942 5816
rect 9382 5797 9738 5803
rect 7900 5763 7912 5797
rect 7946 5763 8256 5797
rect 8314 5763 8624 5797
rect 8658 5763 8980 5797
rect 9014 5763 9324 5797
rect 9382 5763 9692 5797
rect 9726 5763 9738 5797
rect 7900 5757 8256 5763
rect 8314 5757 9324 5763
rect 9382 5757 9738 5763
rect 10586 5798 10942 5804
rect 11000 5804 11010 5816
rect 12000 5804 12010 5816
rect 11000 5798 12010 5804
rect 12068 5804 12078 5816
rect 12068 5798 12424 5804
rect 10586 5764 10598 5798
rect 10632 5764 10942 5798
rect 11000 5764 11310 5798
rect 11344 5764 11666 5798
rect 11700 5764 12010 5798
rect 12068 5764 12378 5798
rect 12412 5764 12424 5798
rect 10586 5758 10942 5764
rect 11000 5758 12010 5764
rect 12068 5758 12424 5764
rect 7802 5704 7878 5710
rect 7802 5670 7814 5704
rect 7866 5670 7878 5704
rect 7802 5664 7878 5670
rect 7980 5704 8056 5710
rect 7980 5670 7992 5704
rect 8044 5670 8056 5704
rect 7980 5664 8056 5670
rect 8158 5704 8234 5710
rect 8158 5670 8170 5704
rect 8222 5670 8234 5704
rect 8158 5664 8234 5670
rect 8336 5704 8412 5710
rect 8336 5670 8348 5704
rect 8400 5670 8412 5704
rect 8336 5664 8412 5670
rect 8514 5704 8590 5710
rect 8514 5670 8526 5704
rect 8578 5670 8590 5704
rect 8514 5664 8590 5670
rect 8692 5704 8768 5710
rect 8692 5670 8704 5704
rect 8756 5670 8768 5704
rect 8692 5664 8768 5670
rect 8870 5704 8946 5710
rect 8870 5670 8882 5704
rect 8934 5670 8946 5704
rect 8870 5664 8946 5670
rect 9048 5704 9124 5710
rect 9048 5670 9060 5704
rect 9112 5670 9124 5704
rect 9048 5664 9124 5670
rect 9226 5704 9302 5710
rect 9226 5670 9238 5704
rect 9290 5670 9302 5704
rect 9226 5664 9302 5670
rect 9404 5704 9480 5710
rect 9404 5670 9416 5704
rect 9468 5670 9480 5704
rect 9404 5664 9480 5670
rect 9582 5704 9658 5710
rect 9582 5670 9594 5704
rect 9646 5670 9658 5704
rect 9582 5664 9658 5670
rect 9760 5704 9836 5710
rect 9760 5670 9772 5704
rect 9824 5670 9836 5704
rect 9760 5664 9836 5670
rect 10488 5705 10564 5711
rect 10488 5671 10500 5705
rect 10552 5671 10564 5705
rect 10488 5665 10564 5671
rect 10666 5705 10742 5711
rect 10666 5671 10678 5705
rect 10730 5671 10742 5705
rect 10666 5665 10742 5671
rect 10844 5705 10920 5711
rect 10844 5671 10856 5705
rect 10908 5671 10920 5705
rect 10844 5665 10920 5671
rect 11022 5705 11098 5711
rect 11022 5671 11034 5705
rect 11086 5671 11098 5705
rect 11022 5665 11098 5671
rect 11200 5705 11276 5711
rect 11200 5671 11212 5705
rect 11264 5671 11276 5705
rect 11200 5665 11276 5671
rect 11378 5705 11454 5711
rect 11378 5671 11390 5705
rect 11442 5671 11454 5705
rect 11378 5665 11454 5671
rect 11556 5705 11632 5711
rect 11556 5671 11568 5705
rect 11620 5671 11632 5705
rect 11556 5665 11632 5671
rect 11734 5705 11810 5711
rect 11734 5671 11746 5705
rect 11798 5671 11810 5705
rect 11734 5665 11810 5671
rect 11912 5705 11988 5711
rect 11912 5671 11924 5705
rect 11976 5671 11988 5705
rect 11912 5665 11988 5671
rect 12090 5705 12166 5711
rect 12090 5671 12102 5705
rect 12154 5671 12166 5705
rect 12090 5665 12166 5671
rect 12268 5705 12344 5711
rect 12268 5671 12280 5705
rect 12332 5671 12344 5705
rect 12268 5665 12344 5671
rect 12446 5705 12522 5711
rect 12446 5671 12458 5705
rect 12510 5671 12522 5705
rect 12446 5665 12522 5671
rect 14869 5643 14875 5841
rect 14909 5643 14915 5841
rect 15047 5701 15053 5899
rect 15087 5701 15093 5899
rect 15209 5841 15219 5899
rect 15277 5841 15287 5899
rect 15031 5643 15041 5701
rect 15099 5643 15109 5701
rect 15225 5643 15231 5841
rect 15265 5643 15271 5841
rect 15403 5701 15409 5899
rect 15443 5701 15449 5899
rect 15565 5841 15575 5899
rect 15633 5841 15643 5899
rect 15387 5643 15397 5701
rect 15455 5643 15465 5701
rect 15581 5643 15587 5841
rect 15621 5643 15627 5841
rect 15759 5701 15765 5899
rect 15799 5701 15805 5899
rect 15921 5841 15931 5899
rect 15989 5841 15999 5899
rect 17053 5841 17063 5899
rect 17121 5841 17131 5899
rect 15742 5643 15752 5701
rect 15810 5643 15820 5701
rect 15937 5643 15943 5841
rect 15977 5643 15983 5841
rect 14869 5631 14915 5643
rect 15047 5631 15093 5643
rect 15225 5631 15271 5643
rect 15403 5631 15449 5643
rect 15581 5631 15627 5643
rect 15759 5631 15805 5643
rect 15937 5631 15983 5643
rect 17069 5643 17075 5841
rect 17109 5643 17115 5841
rect 17247 5701 17253 5899
rect 17287 5701 17293 5899
rect 17409 5841 17419 5899
rect 17477 5841 17487 5899
rect 17232 5643 17242 5701
rect 17300 5643 17310 5701
rect 17425 5643 17431 5841
rect 17465 5643 17471 5841
rect 17603 5701 17609 5899
rect 17643 5701 17649 5899
rect 17765 5841 17775 5899
rect 17833 5841 17843 5899
rect 17587 5643 17597 5701
rect 17655 5643 17665 5701
rect 17781 5643 17787 5841
rect 17821 5643 17827 5841
rect 17959 5701 17965 5899
rect 17999 5701 18005 5899
rect 18121 5841 18131 5899
rect 18189 5841 18199 5899
rect 19254 5841 19264 5899
rect 19322 5841 19332 5899
rect 17943 5643 17953 5701
rect 18011 5643 18021 5701
rect 18137 5643 18143 5841
rect 18177 5643 18183 5841
rect 17069 5631 17115 5643
rect 17247 5631 17293 5643
rect 17425 5631 17471 5643
rect 17603 5631 17649 5643
rect 17781 5631 17827 5643
rect 17959 5631 18005 5643
rect 18137 5631 18183 5643
rect 19269 5643 19275 5841
rect 19309 5643 19315 5841
rect 19447 5701 19453 5899
rect 19487 5701 19493 5899
rect 19609 5841 19619 5899
rect 19677 5841 19687 5899
rect 19432 5643 19442 5701
rect 19500 5643 19510 5701
rect 19625 5643 19631 5841
rect 19665 5643 19671 5841
rect 19803 5701 19809 5899
rect 19843 5701 19849 5899
rect 19965 5841 19975 5899
rect 20033 5841 20043 5899
rect 19787 5643 19797 5701
rect 19855 5643 19865 5701
rect 19981 5643 19987 5841
rect 20021 5643 20027 5841
rect 20159 5701 20165 5899
rect 20199 5701 20205 5899
rect 20321 5841 20331 5899
rect 20462 5841 20472 5899
rect 20143 5643 20153 5701
rect 20211 5643 20221 5701
rect 20337 5643 20343 5841
rect 20377 5643 20383 5841
rect 19269 5631 19315 5643
rect 19447 5631 19493 5643
rect 19625 5631 19671 5643
rect 19803 5631 19849 5643
rect 19981 5631 20027 5643
rect 20159 5631 20205 5643
rect 20337 5631 20383 5643
rect 14943 5584 15019 5590
rect 15121 5584 15197 5590
rect 15299 5584 15375 5590
rect 15477 5584 15553 5590
rect 15655 5584 15731 5590
rect 15833 5584 15909 5590
rect 14863 5550 14955 5584
rect 15007 5550 15133 5584
rect 15185 5550 15311 5584
rect 15363 5550 15489 5584
rect 15541 5550 15667 5584
rect 15719 5550 15845 5584
rect 15897 5550 15909 5584
rect 14943 5544 15019 5550
rect 15121 5544 15197 5550
rect 15299 5544 15553 5550
rect 15655 5544 15731 5550
rect 15833 5544 15909 5550
rect 17143 5584 17219 5590
rect 17321 5584 17397 5590
rect 17499 5584 17575 5590
rect 17677 5584 17753 5590
rect 17855 5584 17931 5590
rect 18033 5584 18109 5590
rect 17143 5550 17155 5584
rect 17207 5550 17333 5584
rect 17385 5550 17511 5584
rect 17563 5550 17689 5584
rect 17741 5550 17867 5584
rect 17919 5550 18045 5584
rect 18097 5550 18109 5584
rect 17143 5544 17219 5550
rect 17321 5544 17397 5550
rect 17499 5544 17753 5550
rect 17855 5544 17931 5550
rect 18033 5544 18109 5550
rect 15368 5462 15485 5544
rect 17575 5462 17692 5544
rect 19343 5532 19353 5590
rect 19411 5584 19421 5590
rect 19521 5584 19597 5590
rect 19699 5584 19775 5590
rect 19877 5584 19953 5590
rect 20055 5584 20131 5590
rect 20233 5584 20309 5590
rect 19411 5550 19533 5584
rect 19585 5550 19711 5584
rect 19763 5550 19889 5584
rect 19941 5550 20067 5584
rect 20119 5550 20245 5584
rect 20297 5550 20309 5584
rect 19411 5532 19421 5550
rect 19521 5544 19597 5550
rect 19699 5544 19843 5550
rect 19877 5544 19953 5550
rect 20055 5544 20131 5550
rect 20233 5544 20309 5550
rect 19726 5462 19843 5544
rect 9760 5345 19843 5462
rect 8158 5232 8234 5238
rect 8336 5232 8412 5238
rect 8514 5232 8590 5238
rect 8692 5232 8768 5238
rect 8870 5232 8946 5238
rect 8158 5198 8170 5232
rect 8222 5198 8348 5232
rect 8400 5198 8526 5232
rect 8578 5198 8704 5232
rect 8756 5198 8882 5232
rect 8934 5198 8946 5232
rect 8158 5192 8234 5198
rect 8336 5192 8412 5198
rect 8514 5192 8590 5198
rect 8692 5192 8768 5198
rect 8870 5192 8946 5198
rect 9048 5232 9124 5238
rect 9226 5232 9302 5238
rect 9404 5232 9480 5238
rect 9582 5232 9658 5238
rect 9760 5232 9836 5345
rect 9048 5198 9060 5232
rect 9112 5198 9238 5232
rect 9290 5198 9416 5232
rect 9468 5198 9594 5232
rect 9646 5198 9772 5232
rect 9824 5198 9836 5232
rect 9048 5192 9124 5198
rect 9226 5192 9302 5198
rect 9404 5192 9480 5198
rect 9582 5192 9658 5198
rect 9760 5192 9836 5198
rect 10488 5232 10564 5345
rect 10666 5232 10742 5238
rect 10844 5232 10920 5238
rect 11022 5232 11098 5238
rect 11200 5232 11276 5238
rect 10488 5198 10500 5232
rect 10552 5198 10678 5232
rect 10730 5198 10856 5232
rect 10908 5198 11034 5232
rect 11086 5198 11212 5232
rect 11264 5198 11276 5232
rect 10488 5192 10564 5198
rect 10666 5192 10742 5198
rect 10844 5192 10920 5198
rect 11022 5192 11098 5198
rect 11200 5192 11276 5198
rect 11378 5232 11454 5238
rect 11556 5232 11632 5238
rect 11734 5232 11810 5238
rect 11912 5232 11988 5238
rect 12090 5232 12166 5238
rect 11378 5198 11390 5232
rect 11442 5198 11568 5232
rect 11620 5198 11746 5232
rect 11798 5198 11924 5232
rect 11976 5198 12102 5232
rect 12154 5198 12166 5232
rect 11378 5192 11454 5198
rect 11556 5192 11632 5198
rect 11734 5192 11810 5198
rect 11912 5192 11988 5198
rect 12090 5192 12166 5198
rect 2819 4319 2829 4321
rect 2083 4263 2149 4319
rect 2507 4303 2829 4319
rect 2507 4269 2524 4303
rect 2558 4269 2829 4303
rect 2507 4263 2829 4269
rect 2887 4319 2897 4321
rect 2937 4319 2993 5118
rect 4599 4319 4609 4321
rect 2887 4303 3421 4319
rect 2887 4269 2946 4303
rect 2980 4269 3370 4303
rect 3404 4269 3421 4303
rect 2887 4263 3421 4269
rect 3863 4263 3929 4319
rect 4287 4303 4609 4319
rect 4287 4269 4304 4303
rect 4338 4269 4609 4303
rect 4287 4263 4609 4269
rect 4667 4319 4677 4321
rect 4720 4319 4776 5118
rect 8068 5087 8078 5145
rect 8136 5139 9858 5145
rect 8136 5105 8446 5139
rect 8480 5105 8802 5139
rect 8836 5105 9158 5139
rect 9192 5105 9514 5139
rect 9548 5105 9858 5139
rect 8136 5099 9858 5105
rect 8136 5087 8146 5099
rect 9848 5087 9858 5099
rect 9916 5087 9926 5145
rect 10398 5087 10408 5145
rect 10466 5139 12188 5145
rect 10466 5105 10776 5139
rect 10810 5105 11132 5139
rect 11166 5105 11488 5139
rect 11522 5105 11844 5139
rect 11878 5105 12188 5139
rect 10466 5099 12188 5105
rect 10466 5087 10476 5099
rect 12178 5087 12188 5099
rect 12246 5087 12256 5145
rect 13796 5131 13872 5137
rect 13974 5131 14050 5137
rect 14152 5131 14228 5137
rect 14330 5131 14406 5137
rect 14508 5131 14584 5137
rect 14686 5131 14762 5137
rect 14864 5131 14940 5137
rect 15042 5131 15118 5137
rect 15220 5131 15296 5137
rect 15398 5131 15474 5137
rect 15576 5131 15652 5137
rect 15754 5131 15830 5137
rect 15932 5131 16008 5137
rect 16110 5131 16186 5137
rect 16288 5131 16364 5137
rect 16466 5131 16542 5137
rect 16644 5131 16720 5137
rect 16822 5131 16898 5137
rect 17000 5131 17076 5137
rect 17178 5131 17254 5137
rect 17356 5131 17432 5137
rect 17534 5131 17610 5137
rect 17712 5131 17788 5137
rect 17890 5131 17966 5137
rect 18068 5131 18144 5137
rect 13791 5097 13808 5131
rect 13860 5097 13986 5131
rect 14038 5097 14164 5131
rect 14216 5097 14342 5131
rect 14394 5097 14520 5131
rect 14572 5097 14698 5131
rect 14750 5097 14876 5131
rect 14928 5097 15054 5131
rect 15106 5097 15232 5131
rect 15284 5097 15410 5131
rect 15462 5097 15588 5131
rect 15640 5097 15766 5131
rect 15818 5097 15944 5131
rect 15996 5097 16122 5131
rect 16174 5097 16300 5131
rect 16352 5097 16478 5131
rect 16530 5097 16656 5131
rect 16708 5097 16834 5131
rect 16886 5097 17012 5131
rect 17064 5097 17190 5131
rect 17242 5097 17368 5131
rect 17420 5097 17546 5131
rect 17598 5097 17724 5131
rect 17776 5097 17902 5131
rect 17954 5097 18080 5131
rect 18132 5097 18212 5131
rect 13791 5057 18212 5097
rect 13791 5053 18131 5057
rect 13791 4995 13894 5053
rect 13952 5047 16030 5053
rect 16088 5047 18131 5053
rect 13952 5013 14262 5047
rect 14296 5013 14618 5047
rect 14652 5013 14974 5047
rect 15008 5013 15330 5047
rect 15364 5013 15686 5047
rect 15720 5013 16030 5047
rect 16088 5013 16398 5047
rect 16432 5013 16754 5047
rect 16788 5013 17110 5047
rect 17144 5013 17466 5047
rect 17500 5013 17822 5047
rect 17856 5013 18131 5047
rect 13952 4995 16030 5013
rect 16088 4995 18131 5013
rect 13791 4991 18131 4995
rect 13884 4985 18131 4991
rect 18121 4940 18131 4985
rect 18248 4940 18258 5057
rect 8246 4877 8256 4935
rect 8314 4923 8324 4935
rect 8780 4931 8790 4935
rect 8848 4931 8858 4935
rect 8715 4923 8725 4931
rect 8314 4917 8725 4923
rect 8314 4883 8624 4917
rect 8658 4883 8725 4917
rect 8314 4877 8725 4883
rect 8715 4873 8725 4877
rect 8917 4923 8927 4931
rect 9670 4923 9680 4935
rect 8917 4917 9680 4923
rect 8917 4883 8980 4917
rect 9014 4883 9336 4917
rect 9370 4883 9680 4917
rect 8917 4877 9680 4883
rect 9738 4877 9748 4935
rect 10576 4877 10586 4935
rect 10644 4923 10654 4935
rect 11466 4932 11476 4935
rect 11534 4932 11544 4935
rect 11394 4923 11404 4932
rect 10644 4917 11404 4923
rect 10644 4883 10954 4917
rect 10988 4883 11310 4917
rect 11344 4883 11404 4917
rect 10644 4877 11404 4883
rect 8917 4873 8927 4877
rect 11394 4874 11404 4877
rect 11596 4923 11606 4932
rect 12000 4923 12010 4935
rect 11596 4917 12010 4923
rect 11596 4883 11666 4917
rect 11700 4883 12010 4917
rect 11596 4877 12010 4883
rect 12068 4877 12078 4935
rect 11596 4874 11606 4877
rect 13706 4843 18056 4870
rect 8158 4824 8234 4830
rect 8158 4790 8170 4824
rect 8222 4790 8234 4824
rect 8158 4662 8234 4790
rect 8336 4824 8412 4830
rect 8336 4790 8348 4824
rect 8400 4790 8412 4824
rect 8336 4784 8412 4790
rect 8514 4824 8590 4830
rect 8514 4790 8526 4824
rect 8578 4790 8590 4824
rect 8514 4784 8590 4790
rect 8692 4824 8768 4830
rect 8692 4790 8704 4824
rect 8756 4790 8768 4824
rect 8692 4784 8768 4790
rect 8870 4824 8946 4830
rect 8870 4790 8882 4824
rect 8934 4790 8946 4824
rect 8870 4784 8946 4790
rect 9048 4824 9124 4830
rect 9048 4790 9060 4824
rect 9112 4790 9124 4824
rect 9048 4784 9124 4790
rect 9226 4824 9302 4830
rect 9226 4790 9238 4824
rect 9290 4790 9302 4824
rect 9226 4784 9302 4790
rect 9404 4824 9480 4830
rect 9404 4790 9416 4824
rect 9468 4790 9480 4824
rect 9404 4784 9480 4790
rect 9582 4824 9658 4830
rect 9582 4790 9594 4824
rect 9646 4790 9658 4824
rect 9582 4784 9658 4790
rect 9760 4824 9836 4830
rect 9760 4790 9772 4824
rect 9824 4790 9836 4824
rect 8336 4662 8412 4668
rect 8514 4662 8590 4668
rect 8692 4662 8768 4668
rect 8870 4662 8946 4668
rect 9048 4662 9124 4668
rect 9226 4662 9302 4668
rect 9404 4662 9480 4668
rect 9582 4662 9658 4668
rect 9760 4662 9836 4790
rect 8158 4628 8170 4662
rect 8222 4628 8348 4662
rect 8400 4628 8526 4662
rect 8578 4628 8704 4662
rect 8756 4628 8882 4662
rect 8934 4628 9060 4662
rect 9112 4628 9238 4662
rect 9290 4628 9416 4662
rect 9468 4628 9594 4662
rect 9646 4628 9772 4662
rect 9824 4628 9836 4662
rect 8158 4622 8234 4628
rect 8336 4622 8412 4628
rect 8514 4622 8590 4628
rect 8692 4622 8768 4628
rect 8870 4622 8946 4628
rect 9048 4622 9124 4628
rect 9226 4622 9302 4628
rect 9404 4622 9480 4628
rect 9582 4622 9658 4628
rect 9760 4622 9836 4628
rect 10488 4824 10564 4830
rect 10488 4790 10500 4824
rect 10552 4790 10564 4824
rect 10488 4662 10564 4790
rect 10666 4824 10742 4830
rect 10666 4790 10678 4824
rect 10730 4790 10742 4824
rect 10666 4784 10742 4790
rect 10844 4824 10920 4830
rect 10844 4790 10856 4824
rect 10908 4790 10920 4824
rect 10844 4784 10920 4790
rect 11022 4824 11098 4830
rect 11022 4790 11034 4824
rect 11086 4790 11098 4824
rect 11022 4784 11098 4790
rect 11200 4824 11276 4830
rect 11200 4790 11212 4824
rect 11264 4790 11276 4824
rect 11200 4784 11276 4790
rect 11378 4824 11454 4830
rect 11378 4790 11390 4824
rect 11442 4790 11454 4824
rect 11378 4784 11454 4790
rect 11556 4824 11632 4830
rect 11556 4790 11568 4824
rect 11620 4790 11632 4824
rect 11556 4784 11632 4790
rect 11734 4824 11810 4830
rect 11734 4790 11746 4824
rect 11798 4790 11810 4824
rect 11734 4784 11810 4790
rect 11912 4824 11988 4830
rect 11912 4790 11924 4824
rect 11976 4790 11988 4824
rect 11912 4784 11988 4790
rect 12090 4824 12166 4830
rect 12090 4790 12102 4824
rect 12154 4790 12166 4824
rect 10666 4662 10742 4668
rect 10844 4662 10920 4668
rect 11022 4662 11098 4668
rect 11200 4662 11276 4668
rect 11378 4662 11454 4668
rect 11556 4662 11632 4668
rect 11734 4662 11810 4668
rect 11912 4662 11988 4668
rect 12090 4662 12166 4790
rect 13706 4785 13716 4843
rect 13774 4825 15852 4843
rect 15910 4825 17988 4843
rect 13774 4791 14084 4825
rect 14118 4791 14440 4825
rect 14474 4791 14796 4825
rect 14830 4791 15152 4825
rect 15186 4791 15508 4825
rect 15542 4791 15852 4825
rect 15910 4791 16220 4825
rect 16254 4791 16576 4825
rect 16610 4791 16932 4825
rect 16966 4791 17288 4825
rect 17322 4791 17644 4825
rect 17678 4791 17988 4825
rect 13774 4785 15852 4791
rect 15910 4785 17988 4791
rect 18046 4785 18056 4843
rect 10488 4628 10500 4662
rect 10552 4628 10678 4662
rect 10730 4628 10856 4662
rect 10908 4628 11034 4662
rect 11086 4628 11212 4662
rect 11264 4628 11390 4662
rect 11442 4628 11568 4662
rect 11620 4628 11746 4662
rect 11798 4628 11924 4662
rect 11976 4628 12102 4662
rect 12154 4628 12166 4662
rect 10488 4622 10564 4628
rect 10666 4622 10742 4628
rect 10844 4622 10920 4628
rect 11022 4622 11098 4628
rect 11200 4622 11276 4628
rect 11378 4622 11454 4628
rect 11556 4622 11632 4628
rect 11734 4622 11810 4628
rect 11912 4622 11988 4628
rect 12090 4622 12166 4628
rect 13796 4742 13872 4747
rect 13974 4742 14050 4747
rect 14152 4742 14228 4747
rect 14330 4742 14406 4747
rect 14508 4742 14584 4747
rect 14686 4742 14762 4747
rect 14864 4742 14940 4747
rect 15042 4742 15118 4747
rect 15220 4742 15296 4747
rect 15398 4742 15474 4747
rect 15576 4742 15652 4747
rect 15754 4742 15830 4747
rect 15932 4742 16008 4747
rect 16110 4742 16186 4747
rect 16288 4742 16364 4747
rect 16466 4742 16542 4747
rect 16644 4742 16720 4747
rect 16822 4742 16898 4747
rect 17000 4742 17076 4747
rect 17178 4742 17254 4747
rect 17356 4742 17432 4747
rect 17534 4742 17610 4747
rect 17712 4742 17788 4747
rect 17890 4742 17966 4747
rect 18068 4742 18144 4747
rect 13796 4741 18213 4742
rect 13796 4707 13808 4741
rect 13860 4707 13986 4741
rect 14038 4707 14164 4741
rect 14216 4707 14342 4741
rect 14394 4707 14520 4741
rect 14572 4707 14698 4741
rect 14750 4707 14876 4741
rect 14928 4707 15054 4741
rect 15106 4707 15232 4741
rect 15284 4707 15410 4741
rect 15462 4707 15588 4741
rect 15640 4707 15766 4741
rect 15818 4707 15944 4741
rect 15996 4707 16122 4741
rect 16174 4707 16300 4741
rect 16352 4707 16478 4741
rect 16530 4707 16656 4741
rect 16708 4707 16834 4741
rect 16886 4707 17012 4741
rect 17064 4707 17190 4741
rect 17242 4707 17368 4741
rect 17420 4707 17546 4741
rect 17598 4707 17724 4741
rect 17776 4707 17902 4741
rect 17954 4707 18080 4741
rect 18132 4707 18213 4741
rect 13796 4631 18213 4707
rect 13796 4597 13808 4631
rect 13860 4597 13986 4631
rect 14038 4597 14164 4631
rect 14216 4597 14342 4631
rect 14394 4597 14520 4631
rect 14572 4597 14698 4631
rect 14750 4597 14876 4631
rect 14928 4597 15054 4631
rect 15106 4597 15232 4631
rect 15284 4597 15410 4631
rect 15462 4597 15588 4631
rect 15640 4597 15766 4631
rect 15818 4597 15944 4631
rect 15996 4597 16122 4631
rect 16174 4597 16300 4631
rect 16352 4597 16478 4631
rect 16530 4597 16656 4631
rect 16708 4597 16834 4631
rect 16886 4597 17012 4631
rect 17064 4597 17190 4631
rect 17242 4597 17368 4631
rect 17420 4597 17546 4631
rect 17598 4597 17724 4631
rect 17776 4597 17902 4631
rect 17954 4597 18080 4631
rect 18132 4597 18213 4631
rect 13796 4591 18213 4597
rect 8715 4575 8725 4577
rect 8068 4517 8078 4575
rect 8136 4569 8725 4575
rect 8917 4575 8927 4577
rect 11396 4575 11406 4576
rect 8917 4569 9858 4575
rect 8136 4535 8446 4569
rect 8480 4535 8725 4569
rect 8917 4535 9158 4569
rect 9192 4535 9514 4569
rect 9548 4535 9858 4569
rect 8136 4529 8725 4535
rect 8136 4517 8146 4529
rect 8715 4519 8725 4529
rect 8917 4529 9858 4535
rect 8917 4519 8927 4529
rect 8780 4517 8790 4519
rect 8848 4517 8858 4519
rect 9848 4517 9858 4529
rect 9916 4517 9926 4575
rect 10398 4517 10408 4575
rect 10466 4569 11406 4575
rect 11598 4575 11608 4576
rect 11598 4569 12188 4575
rect 10466 4535 10776 4569
rect 10810 4535 11132 4569
rect 11166 4535 11406 4569
rect 11598 4535 11844 4569
rect 11878 4535 12188 4569
rect 10466 4529 11406 4535
rect 10466 4517 10476 4529
rect 11396 4518 11406 4529
rect 11598 4529 12188 4535
rect 11598 4518 11608 4529
rect 11468 4517 11478 4518
rect 11536 4517 11546 4518
rect 12178 4517 12188 4529
rect 12246 4517 12256 4575
rect 13798 4553 18213 4591
rect 13798 4495 13894 4553
rect 13952 4547 16030 4553
rect 16088 4547 18132 4553
rect 13952 4513 14262 4547
rect 14296 4513 14618 4547
rect 14652 4513 14974 4547
rect 15008 4513 15330 4547
rect 15364 4513 15686 4547
rect 15720 4513 16030 4547
rect 16088 4513 16398 4547
rect 16432 4513 16754 4547
rect 16788 4513 17110 4547
rect 17144 4513 17466 4547
rect 17500 4513 17822 4547
rect 17856 4513 18132 4547
rect 13952 4495 16030 4513
rect 16088 4495 18132 4513
rect 13798 4472 18132 4495
rect 18122 4436 18132 4472
rect 18249 4436 18259 4553
rect 4667 4303 5201 4319
rect 8246 4307 8256 4365
rect 8314 4353 8324 4365
rect 9670 4353 9680 4365
rect 8314 4347 9680 4353
rect 8314 4313 8624 4347
rect 8658 4313 8980 4347
rect 9014 4313 9336 4347
rect 9370 4313 9680 4347
rect 8314 4307 9680 4313
rect 9738 4307 9748 4365
rect 10576 4307 10586 4365
rect 10644 4353 10654 4365
rect 12000 4353 12010 4365
rect 10644 4347 12010 4353
rect 10644 4313 10954 4347
rect 10988 4313 11310 4347
rect 11344 4313 11666 4347
rect 11700 4313 12010 4347
rect 10644 4307 12010 4313
rect 12068 4307 12078 4365
rect 4667 4269 4726 4303
rect 4760 4269 5150 4303
rect 5184 4269 5201 4303
rect 13706 4285 13716 4343
rect 13774 4331 13784 4343
rect 15842 4331 15852 4343
rect 13774 4325 15852 4331
rect 15910 4331 15920 4343
rect 17620 4331 17630 4387
rect 15910 4325 17630 4331
rect 17752 4331 17762 4387
rect 17978 4331 17988 4343
rect 13774 4291 14084 4325
rect 14118 4291 14440 4325
rect 14474 4291 14796 4325
rect 14830 4291 15152 4325
rect 15186 4291 15508 4325
rect 15542 4291 15852 4325
rect 15910 4291 16220 4325
rect 16254 4291 16576 4325
rect 16610 4291 16932 4325
rect 16966 4291 17288 4325
rect 17322 4291 17630 4325
rect 13774 4285 15852 4291
rect 15910 4285 17630 4291
rect 17752 4286 17988 4331
rect 17688 4285 17988 4286
rect 18046 4285 18056 4343
rect 4667 4263 5201 4269
rect 8158 4254 8234 4260
rect 3394 4225 3404 4227
rect 2348 4219 3404 4225
rect 2348 4185 2360 4219
rect 2394 4185 2572 4219
rect 2606 4185 2784 4219
rect 2818 4185 2996 4219
rect 3030 4185 3208 4219
rect 3242 4185 3404 4219
rect 2348 4179 3404 4185
rect 3394 4173 3404 4179
rect 3569 4173 3579 4227
rect 4118 4174 4128 4228
rect 4293 4225 4303 4228
rect 4293 4219 5246 4225
rect 4293 4185 4352 4219
rect 4386 4185 4564 4219
rect 4598 4185 4776 4219
rect 4810 4185 4988 4219
rect 5022 4185 5200 4219
rect 5234 4185 5246 4219
rect 8158 4220 8170 4254
rect 8222 4220 8234 4254
rect 8158 4214 8234 4220
rect 8336 4254 8412 4260
rect 8336 4220 8348 4254
rect 8400 4220 8412 4254
rect 8336 4214 8412 4220
rect 8514 4254 8590 4260
rect 8514 4220 8526 4254
rect 8578 4220 8590 4254
rect 8514 4214 8590 4220
rect 8692 4254 8768 4260
rect 8692 4220 8704 4254
rect 8756 4220 8768 4254
rect 8692 4214 8768 4220
rect 8870 4254 8946 4260
rect 8870 4220 8882 4254
rect 8934 4220 8946 4254
rect 8870 4214 8946 4220
rect 9048 4254 9124 4260
rect 9048 4220 9060 4254
rect 9112 4220 9124 4254
rect 9048 4214 9124 4220
rect 9226 4254 9302 4260
rect 9226 4220 9238 4254
rect 9290 4220 9302 4254
rect 9226 4214 9302 4220
rect 9404 4254 9480 4260
rect 9404 4220 9416 4254
rect 9468 4220 9480 4254
rect 9404 4214 9480 4220
rect 9582 4254 9658 4260
rect 9582 4220 9594 4254
rect 9646 4220 9658 4254
rect 9582 4214 9658 4220
rect 9760 4254 9836 4260
rect 9760 4220 9772 4254
rect 9824 4220 9836 4254
rect 9760 4214 9836 4220
rect 10488 4254 10564 4260
rect 10488 4220 10500 4254
rect 10552 4220 10564 4254
rect 10488 4214 10564 4220
rect 10666 4254 10742 4260
rect 10666 4220 10678 4254
rect 10730 4220 10742 4254
rect 10666 4214 10742 4220
rect 10844 4254 10920 4260
rect 10844 4220 10856 4254
rect 10908 4220 10920 4254
rect 10844 4214 10920 4220
rect 11022 4254 11098 4260
rect 11022 4220 11034 4254
rect 11086 4220 11098 4254
rect 11022 4214 11098 4220
rect 11200 4254 11276 4260
rect 11200 4220 11212 4254
rect 11264 4220 11276 4254
rect 11200 4214 11276 4220
rect 11378 4254 11454 4260
rect 11378 4220 11390 4254
rect 11442 4220 11454 4254
rect 11378 4214 11454 4220
rect 11556 4254 11632 4260
rect 11556 4220 11568 4254
rect 11620 4220 11632 4254
rect 11556 4214 11632 4220
rect 11734 4254 11810 4260
rect 11734 4220 11746 4254
rect 11798 4220 11810 4254
rect 11734 4214 11810 4220
rect 11912 4254 11988 4260
rect 11912 4220 11924 4254
rect 11976 4220 11988 4254
rect 11912 4214 11988 4220
rect 12090 4254 12166 4260
rect 12090 4220 12102 4254
rect 12154 4220 12166 4254
rect 12090 4214 12166 4220
rect 13796 4241 13872 4247
rect 13974 4241 14050 4247
rect 14152 4241 14228 4247
rect 14330 4241 14406 4247
rect 14508 4241 14584 4247
rect 14686 4241 14762 4247
rect 14864 4241 14940 4247
rect 15042 4241 15118 4247
rect 15220 4241 15296 4247
rect 15398 4241 15474 4247
rect 15576 4241 15652 4247
rect 15754 4241 15830 4247
rect 15932 4241 16008 4247
rect 16110 4241 16186 4247
rect 16288 4241 16364 4247
rect 16466 4241 16542 4247
rect 16644 4241 16720 4247
rect 16822 4241 16898 4247
rect 17000 4241 17076 4247
rect 17178 4241 17254 4247
rect 17356 4241 17610 4247
rect 17712 4241 17788 4247
rect 17890 4241 17966 4247
rect 18068 4241 18144 4247
rect 13796 4207 13808 4241
rect 13860 4207 13986 4241
rect 14038 4207 14164 4241
rect 14216 4207 14342 4241
rect 14394 4207 14520 4241
rect 14572 4207 14698 4241
rect 14750 4207 14876 4241
rect 14928 4207 15054 4241
rect 15106 4207 15232 4241
rect 15284 4207 15410 4241
rect 15462 4207 15588 4241
rect 15640 4207 15766 4241
rect 15818 4207 15944 4241
rect 15996 4207 16122 4241
rect 16174 4207 16300 4241
rect 16352 4207 16478 4241
rect 16530 4207 16656 4241
rect 16708 4207 16834 4241
rect 16886 4207 17012 4241
rect 17064 4207 17190 4241
rect 17242 4207 17368 4241
rect 17420 4207 17452 4241
rect 13796 4201 13872 4207
rect 13974 4201 14050 4207
rect 14152 4201 14228 4207
rect 14330 4201 14406 4207
rect 14508 4201 14584 4207
rect 14686 4201 14762 4207
rect 14864 4201 14940 4207
rect 15042 4201 15118 4207
rect 15220 4201 15296 4207
rect 15398 4201 15474 4207
rect 15576 4201 15652 4207
rect 15754 4201 15830 4207
rect 15932 4201 16008 4207
rect 16110 4201 16186 4207
rect 16288 4201 16364 4207
rect 16466 4201 16542 4207
rect 16644 4201 16720 4207
rect 16822 4201 16898 4207
rect 17000 4201 17076 4207
rect 17178 4201 17254 4207
rect 17356 4201 17452 4207
rect 4293 4179 5246 4185
rect 17442 4183 17452 4201
rect 17510 4207 17546 4241
rect 17598 4207 17724 4241
rect 17776 4207 17902 4241
rect 17954 4207 18080 4241
rect 18132 4207 18144 4241
rect 17510 4201 17610 4207
rect 17712 4201 17788 4207
rect 17890 4201 17966 4207
rect 18068 4201 18144 4207
rect 17510 4183 17520 4201
rect 4293 4174 4303 4179
rect 2246 3995 2256 4049
rect 2522 4043 2532 4049
rect 4874 4043 4884 4051
rect 2522 4037 3368 4043
rect 2522 4003 2686 4037
rect 2720 4003 2898 4037
rect 2932 4003 3110 4037
rect 3144 4003 3322 4037
rect 3356 4003 3368 4037
rect 2522 3997 3368 4003
rect 4030 4037 4884 4043
rect 4030 4003 4042 4037
rect 4076 4003 4254 4037
rect 4288 4003 4466 4037
rect 4500 4003 4678 4037
rect 4712 4003 4884 4037
rect 4030 3997 4884 4003
rect 5150 3997 5160 4051
rect 9761 4008 17630 4125
rect 2522 3995 2532 3997
rect 2819 3959 2829 3961
rect 2295 3953 2829 3959
rect 2295 3919 2312 3953
rect 2346 3919 2736 3953
rect 2770 3919 2829 3953
rect 2295 3903 2829 3919
rect 2887 3959 2897 3961
rect 4599 3959 4609 3961
rect 2887 3953 3209 3959
rect 2887 3919 3158 3953
rect 3192 3919 3209 3953
rect 2887 3903 3209 3919
rect 3567 3903 3633 3959
rect 4075 3953 4609 3959
rect 4075 3919 4092 3953
rect 4126 3919 4516 3953
rect 4550 3919 4609 3953
rect 4075 3903 4609 3919
rect 4667 3959 4677 3961
rect 4667 3953 4989 3959
rect 4667 3919 4938 3953
rect 4972 3919 4989 3953
rect 4667 3903 4989 3919
rect 5347 3903 5413 3959
rect 647 3692 657 3802
rect 767 3692 777 3802
rect 7803 3723 7879 3729
rect 7981 3723 8057 3729
rect 8159 3723 8235 3729
rect 8337 3723 8413 3729
rect 8515 3723 8591 3729
rect 8693 3723 8769 3729
rect 8871 3723 8947 3729
rect 9049 3723 9125 3729
rect 9227 3723 9303 3729
rect 9405 3723 9481 3729
rect 9583 3723 9659 3729
rect 9761 3723 9837 4008
rect 674 3523 750 3692
rect 7803 3689 7815 3723
rect 7867 3689 7993 3723
rect 8045 3689 8171 3723
rect 8223 3689 8349 3723
rect 8401 3689 8527 3723
rect 8579 3689 8705 3723
rect 8757 3689 8883 3723
rect 8935 3689 9061 3723
rect 9113 3689 9239 3723
rect 9291 3689 9417 3723
rect 9469 3689 9595 3723
rect 9647 3689 9773 3723
rect 9825 3689 9837 3723
rect 7803 3683 7879 3689
rect 7981 3683 8057 3689
rect 8159 3683 8235 3689
rect 8337 3683 8413 3689
rect 8515 3683 8591 3689
rect 8693 3683 8769 3689
rect 8871 3683 8947 3689
rect 9049 3683 9125 3689
rect 9227 3683 9303 3689
rect 9405 3683 9481 3689
rect 9583 3683 9659 3689
rect 9761 3683 9837 3689
rect 10490 3723 10566 4008
rect 17620 4007 17630 4008
rect 17752 4007 17762 4125
rect 10668 3723 10744 3729
rect 10846 3723 10922 3729
rect 11024 3723 11100 3729
rect 11202 3723 11278 3729
rect 11380 3723 11456 3729
rect 11558 3723 11634 3729
rect 11736 3723 11812 3729
rect 11914 3723 11990 3729
rect 12092 3723 12168 3729
rect 12270 3723 12346 3729
rect 12448 3723 12524 3729
rect 10490 3689 10502 3723
rect 10554 3689 10680 3723
rect 10732 3689 10858 3723
rect 10910 3689 11036 3723
rect 11088 3689 11214 3723
rect 11266 3689 11392 3723
rect 11444 3689 11570 3723
rect 11622 3689 11748 3723
rect 11800 3689 11926 3723
rect 11978 3689 12104 3723
rect 12156 3689 12282 3723
rect 12334 3689 12460 3723
rect 12512 3689 12524 3723
rect 10490 3683 10566 3689
rect 10668 3683 10744 3689
rect 10846 3683 10922 3689
rect 11024 3683 11100 3689
rect 11202 3683 11278 3689
rect 11380 3683 11456 3689
rect 11558 3683 11634 3689
rect 11736 3683 11812 3689
rect 11914 3683 11990 3689
rect 12092 3683 12168 3689
rect 12270 3683 12346 3689
rect 12448 3683 12524 3689
rect 11404 3645 11414 3646
rect 7713 3587 7723 3645
rect 7781 3639 8718 3645
rect 8910 3639 9859 3645
rect 7781 3605 8091 3639
rect 8125 3605 8447 3639
rect 8481 3605 8718 3639
rect 8910 3605 9159 3639
rect 9193 3605 9515 3639
rect 9549 3605 9859 3639
rect 7781 3599 8718 3605
rect 7781 3587 7791 3599
rect 8708 3587 8718 3599
rect 8910 3599 9859 3605
rect 8910 3587 8920 3599
rect 9849 3587 9859 3599
rect 9917 3587 9927 3645
rect 10400 3587 10410 3645
rect 10468 3639 11414 3645
rect 11606 3645 11616 3646
rect 11606 3639 12546 3645
rect 10468 3605 10778 3639
rect 10812 3605 11134 3639
rect 11168 3605 11414 3639
rect 11606 3605 11846 3639
rect 11880 3605 12202 3639
rect 12236 3605 12546 3639
rect 10468 3599 11414 3605
rect 10468 3587 10478 3599
rect 11404 3588 11414 3599
rect 11606 3599 12546 3605
rect 11606 3588 11616 3599
rect 11468 3587 11478 3588
rect 11536 3587 11546 3588
rect 12536 3587 12546 3599
rect 12604 3587 12614 3645
rect 17442 3633 17452 3651
rect 17354 3627 17452 3633
rect 17199 3593 17366 3627
rect 17418 3593 17452 3627
rect 17510 3633 17520 3651
rect 17510 3627 17608 3633
rect 17510 3593 17544 3627
rect 17596 3593 17762 3627
rect 17354 3587 17608 3593
rect 17280 3549 17326 3555
rect 17636 3550 17682 3555
rect 17621 3549 17631 3550
rect 17268 3543 17630 3549
rect 17268 3530 17286 3543
rect 17320 3530 17630 3543
rect 852 3523 928 3529
rect 1030 3523 1106 3529
rect 1208 3523 1284 3529
rect 1386 3523 1462 3529
rect 1564 3523 1640 3529
rect 1742 3523 1818 3529
rect 1920 3523 1996 3529
rect 2098 3523 2174 3529
rect 2276 3523 2352 3529
rect 2454 3523 2530 3529
rect 2632 3523 2708 3529
rect 2810 3523 2886 3529
rect 2988 3523 3064 3529
rect 3166 3523 3242 3529
rect 3344 3523 3420 3529
rect 674 3489 686 3523
rect 738 3489 864 3523
rect 916 3489 1042 3523
rect 1094 3489 1220 3523
rect 1272 3489 1398 3523
rect 1450 3489 1576 3523
rect 1628 3489 1754 3523
rect 1806 3489 1932 3523
rect 1984 3489 2110 3523
rect 2162 3489 2288 3523
rect 2340 3489 2466 3523
rect 2518 3489 2644 3523
rect 2696 3489 2822 3523
rect 2874 3489 3000 3523
rect 3052 3489 3178 3523
rect 3230 3489 3356 3523
rect 3408 3489 3420 3523
rect 674 3483 750 3489
rect 852 3483 928 3489
rect 1030 3483 1106 3489
rect 1208 3483 1284 3489
rect 1386 3483 1462 3489
rect 1564 3483 1640 3489
rect 1742 3483 1818 3489
rect 1920 3483 1996 3489
rect 2098 3483 2174 3489
rect 2276 3483 2352 3489
rect 2454 3483 2530 3489
rect 2632 3483 2708 3489
rect 2810 3483 2886 3489
rect 2988 3483 3064 3489
rect 3166 3483 3242 3489
rect 3344 3483 3420 3489
rect 4074 3523 4150 3529
rect 4252 3523 4328 3529
rect 4430 3523 4506 3529
rect 4608 3523 4684 3529
rect 4786 3523 4862 3529
rect 4964 3523 5040 3529
rect 5142 3523 5218 3529
rect 5320 3523 5396 3529
rect 5498 3523 5574 3529
rect 5676 3523 5752 3529
rect 5854 3523 5930 3529
rect 6032 3523 6108 3529
rect 6210 3523 6286 3529
rect 6388 3523 6464 3529
rect 6566 3523 6642 3529
rect 6744 3523 6820 3529
rect 4074 3489 4086 3523
rect 4138 3489 4264 3523
rect 4316 3489 4442 3523
rect 4494 3489 4620 3523
rect 4672 3489 4798 3523
rect 4850 3489 4976 3523
rect 5028 3489 5154 3523
rect 5206 3489 5332 3523
rect 5384 3489 5510 3523
rect 5562 3489 5688 3523
rect 5740 3489 5866 3523
rect 5918 3489 6044 3523
rect 6096 3489 6222 3523
rect 6274 3489 6400 3523
rect 6452 3489 6578 3523
rect 6630 3489 6756 3523
rect 6808 3489 6820 3523
rect 4074 3483 4150 3489
rect 4252 3483 4328 3489
rect 4430 3483 4506 3489
rect 4608 3483 4684 3489
rect 4786 3483 4862 3489
rect 4964 3483 5040 3489
rect 5142 3483 5218 3489
rect 5320 3483 5396 3489
rect 5498 3483 5574 3489
rect 5676 3483 5752 3489
rect 5854 3483 5930 3489
rect 6032 3483 6108 3489
rect 6210 3483 6286 3489
rect 6388 3483 6464 3489
rect 6566 3483 6642 3489
rect 6744 3483 6820 3489
rect 4876 3445 4886 3448
rect 584 3387 594 3445
rect 652 3439 2018 3445
rect 652 3405 962 3439
rect 996 3405 1318 3439
rect 1352 3405 1674 3439
rect 1708 3405 2018 3439
rect 652 3399 2018 3405
rect 652 3387 662 3399
rect 2008 3387 2018 3399
rect 2076 3399 2256 3445
rect 2522 3439 3442 3445
rect 2522 3405 2742 3439
rect 2776 3405 3098 3439
rect 3132 3405 3442 3439
rect 2076 3387 2086 3399
rect 2246 3391 2256 3399
rect 2522 3399 3442 3405
rect 2522 3391 2532 3399
rect 3432 3387 3442 3399
rect 3500 3399 3994 3445
rect 4052 3439 4886 3445
rect 5152 3445 5162 3448
rect 4052 3405 4362 3439
rect 4396 3405 4718 3439
rect 4752 3405 4886 3439
rect 3500 3387 3510 3399
rect 3984 3387 3994 3399
rect 4052 3399 4886 3405
rect 4052 3387 4062 3399
rect 4876 3394 4886 3399
rect 5152 3399 5418 3445
rect 5476 3439 6842 3445
rect 5476 3405 5786 3439
rect 5820 3405 6142 3439
rect 6176 3405 6498 3439
rect 6532 3405 6842 3439
rect 5152 3394 5162 3399
rect 5408 3387 5418 3399
rect 5476 3399 6842 3405
rect 5476 3387 5486 3399
rect 6832 3387 6842 3399
rect 6900 3387 6910 3445
rect 8247 3423 8257 3435
rect 7901 3417 8257 3423
rect 8315 3423 8325 3435
rect 9315 3423 9325 3435
rect 8315 3417 9325 3423
rect 9383 3423 9393 3435
rect 10934 3423 10944 3435
rect 9383 3417 9739 3423
rect 7901 3383 7913 3417
rect 7947 3383 8257 3417
rect 8315 3383 8625 3417
rect 8659 3383 8981 3417
rect 9015 3383 9325 3417
rect 9383 3383 9693 3417
rect 9727 3383 9739 3417
rect 7901 3377 8257 3383
rect 8315 3377 9325 3383
rect 9383 3377 9739 3383
rect 10588 3417 10944 3423
rect 11002 3423 11012 3435
rect 12002 3423 12012 3435
rect 11002 3417 12012 3423
rect 12070 3423 12080 3435
rect 12070 3417 12426 3423
rect 10588 3383 10600 3417
rect 10634 3383 10944 3417
rect 11002 3383 11312 3417
rect 11346 3383 11668 3417
rect 11702 3383 12012 3417
rect 12070 3383 12380 3417
rect 12414 3383 12426 3417
rect 10588 3377 10944 3383
rect 11002 3377 12012 3383
rect 12070 3377 12426 3383
rect 7803 3333 7879 3339
rect 7803 3299 7815 3333
rect 7867 3299 7879 3333
rect 1474 3223 1484 3235
rect 772 3217 1484 3223
rect 1542 3223 1552 3235
rect 2542 3223 2552 3235
rect 1542 3217 2552 3223
rect 2610 3223 2620 3235
rect 4874 3223 4884 3235
rect 2610 3217 3322 3223
rect 772 3183 784 3217
rect 818 3183 1140 3217
rect 1174 3183 1484 3217
rect 1542 3183 1852 3217
rect 1886 3183 2208 3217
rect 2242 3183 2552 3217
rect 2610 3183 2920 3217
rect 2954 3183 3276 3217
rect 3310 3183 3322 3217
rect 772 3177 1484 3183
rect 1542 3177 2552 3183
rect 2610 3177 3322 3183
rect 4172 3217 4884 3223
rect 4942 3223 4952 3235
rect 5942 3223 5952 3235
rect 4942 3217 5952 3223
rect 6010 3223 6020 3235
rect 7803 3223 7879 3299
rect 7981 3333 8057 3339
rect 7981 3299 7993 3333
rect 8045 3299 8057 3333
rect 7981 3293 8057 3299
rect 8159 3333 8235 3339
rect 8159 3299 8171 3333
rect 8223 3299 8235 3333
rect 8159 3293 8235 3299
rect 8337 3333 8413 3339
rect 8337 3299 8349 3333
rect 8401 3299 8413 3333
rect 8337 3293 8413 3299
rect 8515 3333 8591 3339
rect 8515 3299 8527 3333
rect 8579 3299 8591 3333
rect 8515 3293 8591 3299
rect 8693 3333 8769 3339
rect 8693 3299 8705 3333
rect 8757 3299 8769 3333
rect 8693 3293 8769 3299
rect 8871 3333 8947 3339
rect 8871 3299 8883 3333
rect 8935 3299 8947 3333
rect 8871 3293 8947 3299
rect 9049 3333 9125 3339
rect 9049 3299 9061 3333
rect 9113 3299 9125 3333
rect 9049 3293 9125 3299
rect 9227 3333 9303 3339
rect 9227 3299 9239 3333
rect 9291 3299 9303 3333
rect 9227 3293 9303 3299
rect 9405 3333 9481 3339
rect 9405 3299 9417 3333
rect 9469 3299 9481 3333
rect 9405 3293 9481 3299
rect 9583 3333 9659 3339
rect 9583 3299 9595 3333
rect 9647 3299 9659 3333
rect 9583 3293 9659 3299
rect 9761 3333 9837 3339
rect 9761 3299 9773 3333
rect 9825 3299 9837 3333
rect 7981 3223 8057 3229
rect 8159 3223 8235 3229
rect 8337 3223 8413 3229
rect 8515 3223 8591 3229
rect 8693 3223 8769 3229
rect 8871 3223 8947 3229
rect 9049 3223 9125 3229
rect 9227 3223 9303 3229
rect 9405 3223 9481 3229
rect 9583 3223 9659 3229
rect 9761 3223 9837 3299
rect 6010 3217 6722 3223
rect 4172 3183 4184 3217
rect 4218 3183 4540 3217
rect 4574 3183 4884 3217
rect 4942 3183 5252 3217
rect 5286 3183 5608 3217
rect 5642 3183 5952 3217
rect 6010 3183 6320 3217
rect 6354 3183 6676 3217
rect 6710 3183 6722 3217
rect 7803 3189 7815 3223
rect 7867 3189 7993 3223
rect 8045 3189 8171 3223
rect 8223 3189 8349 3223
rect 8401 3189 8527 3223
rect 8579 3189 8705 3223
rect 8757 3189 8883 3223
rect 8935 3189 9061 3223
rect 9113 3189 9239 3223
rect 9291 3189 9417 3223
rect 9469 3189 9595 3223
rect 9647 3189 9773 3223
rect 9825 3189 9837 3223
rect 7803 3183 7879 3189
rect 7981 3183 8057 3189
rect 8159 3183 8235 3189
rect 8337 3183 8413 3189
rect 8515 3183 8591 3189
rect 8693 3183 8769 3189
rect 8871 3183 8947 3189
rect 9049 3183 9125 3189
rect 9227 3183 9303 3189
rect 9405 3183 9481 3189
rect 9583 3183 9659 3189
rect 9761 3183 9837 3189
rect 10490 3333 10566 3339
rect 10490 3299 10502 3333
rect 10554 3299 10566 3333
rect 10490 3223 10566 3299
rect 10668 3333 10744 3339
rect 10668 3299 10680 3333
rect 10732 3299 10744 3333
rect 10668 3293 10744 3299
rect 10846 3333 10922 3339
rect 10846 3299 10858 3333
rect 10910 3299 10922 3333
rect 10846 3293 10922 3299
rect 11024 3333 11100 3339
rect 11024 3299 11036 3333
rect 11088 3299 11100 3333
rect 11024 3293 11100 3299
rect 11202 3333 11278 3339
rect 11202 3299 11214 3333
rect 11266 3299 11278 3333
rect 11202 3293 11278 3299
rect 11380 3333 11456 3339
rect 11380 3299 11392 3333
rect 11444 3299 11456 3333
rect 11380 3293 11456 3299
rect 11558 3333 11634 3339
rect 11558 3299 11570 3333
rect 11622 3299 11634 3333
rect 11558 3293 11634 3299
rect 11736 3333 11812 3339
rect 11736 3299 11748 3333
rect 11800 3299 11812 3333
rect 11736 3293 11812 3299
rect 11914 3333 11990 3339
rect 11914 3299 11926 3333
rect 11978 3299 11990 3333
rect 11914 3293 11990 3299
rect 12092 3333 12168 3339
rect 12092 3299 12104 3333
rect 12156 3299 12168 3333
rect 12092 3293 12168 3299
rect 12270 3333 12346 3339
rect 12270 3299 12282 3333
rect 12334 3299 12346 3333
rect 12270 3293 12346 3299
rect 12448 3333 12524 3339
rect 12448 3299 12460 3333
rect 12512 3299 12524 3333
rect 10668 3223 10744 3229
rect 10846 3223 10922 3229
rect 11024 3223 11100 3229
rect 11202 3223 11278 3229
rect 11380 3223 11456 3229
rect 11558 3223 11634 3229
rect 11736 3223 11812 3229
rect 11914 3223 11990 3229
rect 12092 3223 12168 3229
rect 12270 3223 12346 3229
rect 12448 3223 12524 3299
rect 17264 3278 17274 3530
rect 17332 3493 17630 3530
rect 17332 3492 17350 3493
rect 17332 3278 17342 3492
rect 17615 3491 17630 3493
rect 17615 3433 17631 3491
rect 17752 3433 17762 3550
rect 17442 3279 17452 3416
rect 17510 3279 17520 3416
rect 17280 3275 17326 3278
rect 17442 3275 17520 3279
rect 10490 3189 10502 3223
rect 10554 3189 10680 3223
rect 10732 3189 10858 3223
rect 10910 3189 11036 3223
rect 11088 3189 11214 3223
rect 11266 3189 11392 3223
rect 11444 3189 11570 3223
rect 11622 3189 11748 3223
rect 11800 3189 11926 3223
rect 11978 3189 12104 3223
rect 12156 3189 12282 3223
rect 12334 3189 12460 3223
rect 12512 3189 12524 3223
rect 17354 3237 17430 3243
rect 17354 3203 17366 3237
rect 17418 3203 17430 3237
rect 17354 3197 17430 3203
rect 17532 3237 17608 3243
rect 17532 3203 17544 3237
rect 17596 3203 17608 3237
rect 17532 3197 17608 3203
rect 10490 3183 10566 3189
rect 10668 3183 10744 3189
rect 10846 3183 10922 3189
rect 11024 3183 11100 3189
rect 11202 3183 11278 3189
rect 11380 3183 11456 3189
rect 11558 3183 11634 3189
rect 11736 3183 11812 3189
rect 11914 3183 11990 3189
rect 12092 3183 12168 3189
rect 12270 3183 12346 3189
rect 12448 3183 12524 3189
rect 4172 3177 4884 3183
rect 4942 3177 5952 3183
rect 6010 3177 6722 3183
rect 18888 3154 19016 5228
rect 19255 5122 19331 5128
rect 19433 5122 19509 5128
rect 19611 5122 19687 5128
rect 19789 5122 19865 5128
rect 19967 5122 20043 5128
rect 20145 5122 20221 5128
rect 20321 5122 20331 5141
rect 20477 5128 20525 5141
rect 20477 5122 20577 5128
rect 20679 5122 20755 5128
rect 20857 5122 20933 5128
rect 21035 5122 21111 5128
rect 21213 5122 21289 5128
rect 21391 5122 21467 5128
rect 21569 5122 21645 5128
rect 19166 5106 19267 5122
rect 19165 4986 19175 5106
rect 19233 5088 19267 5106
rect 19319 5088 19445 5122
rect 19497 5088 19623 5122
rect 19675 5110 19801 5122
rect 19675 5088 19709 5110
rect 19233 5038 19709 5088
rect 19233 5004 19543 5038
rect 19577 5021 19709 5038
rect 19767 5088 19801 5110
rect 19853 5088 19979 5122
rect 20031 5088 20157 5122
rect 20209 5088 20331 5122
rect 20477 5088 20513 5122
rect 20565 5088 20691 5122
rect 20743 5088 20869 5122
rect 20921 5088 21047 5122
rect 21099 5115 21225 5122
rect 21099 5088 21132 5115
rect 19767 5038 20331 5088
rect 19767 5021 19899 5038
rect 19577 5004 19899 5021
rect 19933 5004 20255 5038
rect 20289 5004 20331 5038
rect 19233 5001 20331 5004
rect 20477 5038 21132 5088
rect 20477 5004 20611 5038
rect 20645 5004 20967 5038
rect 21001 5026 21132 5038
rect 21190 5088 21225 5115
rect 21277 5088 21403 5122
rect 21455 5088 21581 5122
rect 21633 5106 21736 5122
rect 21633 5088 21667 5106
rect 21190 5038 21667 5088
rect 21190 5026 21323 5038
rect 21001 5004 21323 5026
rect 21357 5004 21667 5038
rect 21725 5022 21736 5106
rect 20477 5001 21667 5004
rect 19233 4998 21667 5001
rect 19233 4986 19243 4998
rect 21657 4986 21667 4998
rect 21725 4986 21735 5022
rect 19343 4776 19353 4834
rect 19411 4822 19421 4834
rect 20055 4822 20065 4831
rect 19411 4816 20065 4822
rect 20123 4822 20133 4831
rect 20769 4822 20779 4835
rect 20123 4816 20779 4822
rect 20837 4822 20847 4835
rect 21479 4822 21489 4834
rect 20837 4816 21489 4822
rect 19411 4782 19721 4816
rect 19755 4782 20065 4816
rect 20123 4782 20433 4816
rect 20467 4782 20779 4816
rect 20837 4782 21145 4816
rect 21179 4782 21489 4816
rect 19411 4776 20065 4782
rect 20055 4773 20065 4776
rect 20123 4777 20779 4782
rect 20837 4777 21489 4782
rect 20123 4776 21489 4777
rect 21547 4776 21557 4834
rect 20123 4773 20133 4776
rect 19255 4733 19331 4738
rect 19433 4733 19509 4738
rect 19611 4733 19687 4738
rect 19789 4733 19865 4738
rect 19967 4733 20043 4738
rect 20145 4733 20221 4738
rect 20323 4733 20399 4738
rect 20501 4733 20577 4738
rect 20679 4733 20755 4738
rect 20857 4733 20933 4738
rect 21035 4733 21111 4738
rect 21213 4733 21289 4738
rect 21391 4733 21467 4738
rect 21569 4733 21645 4738
rect 19168 4732 21736 4733
rect 19168 4725 19267 4732
rect 19166 4546 19176 4725
rect 19234 4698 19267 4725
rect 19319 4698 19445 4732
rect 19497 4698 19623 4732
rect 19675 4719 19801 4732
rect 19675 4698 19710 4719
rect 19234 4624 19710 4698
rect 19234 4590 19267 4624
rect 19319 4590 19445 4624
rect 19497 4590 19623 4624
rect 19675 4590 19710 4624
rect 19165 4488 19175 4546
rect 19234 4540 19710 4590
rect 19234 4517 19543 4540
rect 19233 4506 19543 4517
rect 19577 4511 19710 4540
rect 19768 4698 19801 4719
rect 19853 4698 19979 4732
rect 20031 4698 20157 4732
rect 20209 4698 20335 4732
rect 20387 4730 20513 4732
rect 20387 4698 20420 4730
rect 19768 4624 20420 4698
rect 19768 4590 19801 4624
rect 19853 4590 19979 4624
rect 20031 4590 20157 4624
rect 20209 4590 20335 4624
rect 20387 4590 20420 4624
rect 19768 4540 20420 4590
rect 19768 4511 19899 4540
rect 19577 4506 19899 4511
rect 19933 4506 20255 4540
rect 20289 4522 20420 4540
rect 20478 4698 20513 4730
rect 20565 4698 20691 4732
rect 20743 4698 20869 4732
rect 20921 4698 21047 4732
rect 21099 4723 21225 4732
rect 21099 4698 21133 4723
rect 20478 4624 21133 4698
rect 20478 4590 20513 4624
rect 20565 4590 20691 4624
rect 20743 4590 20869 4624
rect 20921 4590 21047 4624
rect 21099 4590 21133 4624
rect 20478 4540 21133 4590
rect 20478 4522 20611 4540
rect 20289 4506 20611 4522
rect 20645 4506 20967 4540
rect 21001 4515 21133 4540
rect 21191 4698 21225 4723
rect 21277 4698 21403 4732
rect 21455 4698 21581 4732
rect 21633 4716 21736 4732
rect 21633 4698 21667 4716
rect 21191 4624 21667 4698
rect 21191 4590 21225 4624
rect 21277 4590 21403 4624
rect 21455 4590 21581 4624
rect 21633 4590 21667 4624
rect 21191 4540 21667 4590
rect 21191 4515 21323 4540
rect 21001 4506 21323 4515
rect 21357 4506 21667 4540
rect 21725 4521 21736 4716
rect 19233 4500 21667 4506
rect 19233 4488 19243 4500
rect 21657 4488 21667 4500
rect 21725 4488 21735 4521
rect 19343 4278 19353 4336
rect 19411 4324 19421 4336
rect 20055 4324 20065 4331
rect 19411 4318 20065 4324
rect 20123 4324 20133 4331
rect 20768 4324 20778 4334
rect 20123 4318 20778 4324
rect 20836 4324 20846 4334
rect 21479 4324 21489 4336
rect 20836 4318 21489 4324
rect 19411 4284 19721 4318
rect 19755 4284 20065 4318
rect 20123 4284 20433 4318
rect 20467 4284 20778 4318
rect 20836 4284 21145 4318
rect 21179 4284 21489 4318
rect 19411 4278 20065 4284
rect 20055 4273 20065 4278
rect 20123 4278 20778 4284
rect 20123 4273 20133 4278
rect 20768 4276 20778 4278
rect 20836 4278 21489 4284
rect 21547 4278 21557 4336
rect 20836 4276 20846 4278
rect 19255 4234 19331 4240
rect 19433 4234 19509 4240
rect 19611 4234 19687 4240
rect 19789 4234 19865 4240
rect 19967 4234 20043 4240
rect 20145 4234 20221 4240
rect 20323 4234 20399 4240
rect 20501 4234 20577 4240
rect 20679 4234 20755 4240
rect 20857 4234 20933 4240
rect 21035 4234 21111 4240
rect 21213 4234 21289 4240
rect 21391 4234 21467 4240
rect 21569 4234 21645 4240
rect 19167 4224 19267 4234
rect 19165 3990 19175 4224
rect 19233 4200 19267 4224
rect 19319 4200 19445 4234
rect 19497 4200 19623 4234
rect 19675 4223 19801 4234
rect 19675 4200 19709 4223
rect 19233 4126 19709 4200
rect 19233 4092 19267 4126
rect 19319 4092 19445 4126
rect 19497 4092 19623 4126
rect 19675 4092 19709 4126
rect 19233 4042 19709 4092
rect 19233 4008 19543 4042
rect 19577 4015 19709 4042
rect 19767 4200 19801 4223
rect 19853 4200 19979 4234
rect 20031 4200 20157 4234
rect 20209 4200 20335 4234
rect 20387 4223 20513 4234
rect 20387 4200 20422 4223
rect 19767 4126 20422 4200
rect 19767 4092 19801 4126
rect 19853 4092 19979 4126
rect 20031 4092 20157 4126
rect 20209 4092 20335 4126
rect 20387 4092 20422 4126
rect 19767 4042 20422 4092
rect 19767 4015 19899 4042
rect 19577 4008 19899 4015
rect 19933 4008 20255 4042
rect 20289 4015 20422 4042
rect 20480 4200 20513 4223
rect 20565 4200 20691 4234
rect 20743 4200 20869 4234
rect 20921 4200 21047 4234
rect 21099 4230 21225 4234
rect 21099 4200 21133 4230
rect 20480 4126 21133 4200
rect 20480 4092 20513 4126
rect 20565 4092 20691 4126
rect 20743 4092 20869 4126
rect 20921 4092 21047 4126
rect 21099 4092 21133 4126
rect 20480 4042 21133 4092
rect 20480 4015 20611 4042
rect 20289 4008 20611 4015
rect 20645 4008 20967 4042
rect 21001 4022 21133 4042
rect 21191 4200 21225 4230
rect 21277 4200 21403 4234
rect 21455 4200 21581 4234
rect 21633 4218 21735 4234
rect 21633 4200 21666 4218
rect 21191 4126 21666 4200
rect 21191 4092 21225 4126
rect 21277 4092 21403 4126
rect 21455 4092 21581 4126
rect 21633 4092 21666 4126
rect 21191 4042 21666 4092
rect 21724 4048 21735 4218
rect 21191 4022 21323 4042
rect 21001 4008 21323 4022
rect 21357 4010 21666 4042
rect 21357 4008 21667 4010
rect 19233 4002 21667 4008
rect 19233 3990 19243 4002
rect 21657 3990 21667 4002
rect 21725 3990 21735 4048
rect 19343 3780 19353 3838
rect 19411 3826 19421 3838
rect 20055 3826 20065 3837
rect 19411 3820 20065 3826
rect 20123 3826 20133 3837
rect 20764 3826 20774 3841
rect 20123 3820 20774 3826
rect 20832 3826 20842 3841
rect 21479 3826 21489 3838
rect 20832 3820 21489 3826
rect 19411 3786 19721 3820
rect 19755 3786 20065 3820
rect 20123 3786 20433 3820
rect 20467 3786 20774 3820
rect 20832 3786 21145 3820
rect 21179 3786 21489 3820
rect 19411 3780 20065 3786
rect 20055 3779 20065 3780
rect 20123 3783 20774 3786
rect 20832 3783 21489 3786
rect 20123 3780 21489 3783
rect 21547 3780 21557 3838
rect 20123 3779 20133 3780
rect 19255 3736 19331 3742
rect 19433 3736 19509 3742
rect 19611 3736 19687 3742
rect 19789 3736 19865 3742
rect 19967 3736 20043 3742
rect 20145 3736 20221 3742
rect 20323 3736 20399 3742
rect 20501 3736 20577 3742
rect 20679 3736 20755 3742
rect 20857 3736 20933 3742
rect 21035 3736 21111 3742
rect 21213 3736 21289 3742
rect 21391 3736 21467 3742
rect 21569 3736 21645 3742
rect 19165 3492 19175 3736
rect 19233 3702 19267 3736
rect 19319 3702 19445 3736
rect 19497 3702 19623 3736
rect 19675 3726 19801 3736
rect 19675 3702 19708 3726
rect 19233 3628 19708 3702
rect 19233 3594 19267 3628
rect 19319 3594 19445 3628
rect 19497 3594 19623 3628
rect 19675 3594 19708 3628
rect 19233 3544 19708 3594
rect 19233 3510 19543 3544
rect 19577 3518 19708 3544
rect 19766 3702 19801 3726
rect 19853 3702 19979 3736
rect 20031 3702 20157 3736
rect 20209 3702 20335 3736
rect 20387 3723 20513 3736
rect 20387 3702 20420 3723
rect 19766 3628 20420 3702
rect 19766 3594 19801 3628
rect 19853 3594 19979 3628
rect 20031 3594 20157 3628
rect 20209 3594 20335 3628
rect 20387 3594 20420 3628
rect 19766 3544 20420 3594
rect 19766 3518 19899 3544
rect 19577 3510 19899 3518
rect 19933 3510 20255 3544
rect 20289 3515 20420 3544
rect 20478 3702 20513 3723
rect 20565 3702 20691 3736
rect 20743 3702 20869 3736
rect 20921 3702 21047 3736
rect 21099 3721 21225 3736
rect 21099 3702 21133 3721
rect 20478 3628 21133 3702
rect 20478 3594 20513 3628
rect 20565 3594 20691 3628
rect 20743 3594 20869 3628
rect 20921 3594 21047 3628
rect 21099 3594 21133 3628
rect 20478 3544 21133 3594
rect 20478 3515 20611 3544
rect 20289 3510 20611 3515
rect 20645 3510 20967 3544
rect 21001 3513 21133 3544
rect 21191 3702 21225 3721
rect 21277 3702 21403 3736
rect 21455 3702 21581 3736
rect 21633 3702 21667 3736
rect 21191 3628 21667 3702
rect 21191 3594 21225 3628
rect 21277 3594 21403 3628
rect 21455 3594 21581 3628
rect 21633 3594 21667 3628
rect 21191 3544 21667 3594
rect 21191 3513 21323 3544
rect 21001 3510 21323 3513
rect 21357 3510 21667 3544
rect 19233 3504 21667 3510
rect 19233 3492 19243 3504
rect 21657 3492 21667 3504
rect 21725 3492 21735 3736
rect 19343 3282 19353 3340
rect 19411 3328 19421 3340
rect 19700 3328 19710 3339
rect 19411 3282 19710 3328
rect 19768 3328 19778 3339
rect 20056 3328 20066 3339
rect 19700 3281 19710 3282
rect 19768 3282 20066 3328
rect 20124 3328 20134 3339
rect 20413 3328 20423 3340
rect 19768 3281 19778 3282
rect 20056 3281 20066 3282
rect 20124 3282 20423 3328
rect 20481 3328 20491 3340
rect 20769 3328 20779 3337
rect 20481 3282 20779 3328
rect 20837 3328 20847 3337
rect 21125 3328 21135 3338
rect 20124 3281 20134 3282
rect 20769 3279 20779 3282
rect 20837 3282 21135 3328
rect 21193 3328 21203 3338
rect 21479 3328 21489 3340
rect 20837 3279 20847 3282
rect 21125 3280 21135 3282
rect 21193 3282 21489 3328
rect 21547 3282 21557 3340
rect 21193 3280 21203 3282
rect 19255 3238 19331 3244
rect 19255 3204 19267 3238
rect 19319 3204 19331 3238
rect 19255 3198 19331 3204
rect 19433 3238 19509 3244
rect 19433 3204 19445 3238
rect 19497 3204 19509 3238
rect 19433 3198 19509 3204
rect 19611 3238 19687 3244
rect 19611 3204 19623 3238
rect 19675 3204 19687 3238
rect 19611 3198 19687 3204
rect 19789 3238 19865 3244
rect 19789 3204 19801 3238
rect 19853 3204 19865 3238
rect 19789 3198 19865 3204
rect 19967 3238 20043 3244
rect 19967 3204 19979 3238
rect 20031 3204 20043 3238
rect 19967 3198 20043 3204
rect 20145 3238 20221 3244
rect 20145 3204 20157 3238
rect 20209 3204 20221 3238
rect 20145 3198 20221 3204
rect 20323 3238 20399 3244
rect 20323 3204 20335 3238
rect 20387 3204 20399 3238
rect 20323 3198 20399 3204
rect 20501 3238 20577 3244
rect 20501 3204 20513 3238
rect 20565 3204 20577 3238
rect 20501 3198 20577 3204
rect 20679 3238 20755 3244
rect 20679 3204 20691 3238
rect 20743 3204 20755 3238
rect 20679 3198 20755 3204
rect 20857 3238 20933 3244
rect 20857 3204 20869 3238
rect 20921 3204 20933 3238
rect 20857 3198 20933 3204
rect 21035 3238 21111 3244
rect 21035 3204 21047 3238
rect 21099 3204 21111 3238
rect 21035 3198 21111 3204
rect 21213 3238 21289 3244
rect 21213 3204 21225 3238
rect 21277 3204 21289 3238
rect 21213 3198 21289 3204
rect 21391 3238 21467 3244
rect 21391 3204 21403 3238
rect 21455 3204 21467 3238
rect 21391 3198 21467 3204
rect 21569 3238 21645 3244
rect 21569 3204 21581 3238
rect 21633 3204 21645 3238
rect 21569 3198 21645 3204
rect 21891 3180 22019 5236
rect 674 3133 750 3139
rect 674 3099 686 3133
rect 738 3099 750 3133
rect 674 3023 750 3099
rect 852 3133 928 3139
rect 852 3099 864 3133
rect 916 3099 928 3133
rect 852 3093 928 3099
rect 1030 3133 1106 3139
rect 1030 3099 1042 3133
rect 1094 3099 1106 3133
rect 1030 3093 1106 3099
rect 1208 3133 1284 3139
rect 1208 3099 1220 3133
rect 1272 3099 1284 3133
rect 1208 3093 1284 3099
rect 1386 3133 1462 3139
rect 1386 3099 1398 3133
rect 1450 3099 1462 3133
rect 1386 3093 1462 3099
rect 1564 3133 1640 3139
rect 1564 3099 1576 3133
rect 1628 3099 1640 3133
rect 1564 3093 1640 3099
rect 1742 3133 1818 3139
rect 1742 3099 1754 3133
rect 1806 3099 1818 3133
rect 1742 3093 1818 3099
rect 1920 3133 1996 3139
rect 1920 3099 1932 3133
rect 1984 3099 1996 3133
rect 1920 3093 1996 3099
rect 2098 3133 2174 3139
rect 2098 3099 2110 3133
rect 2162 3099 2174 3133
rect 2098 3093 2174 3099
rect 2276 3133 2352 3139
rect 2276 3099 2288 3133
rect 2340 3099 2352 3133
rect 2276 3093 2352 3099
rect 2454 3133 2530 3139
rect 2454 3099 2466 3133
rect 2518 3099 2530 3133
rect 2454 3093 2530 3099
rect 2632 3133 2708 3139
rect 2632 3099 2644 3133
rect 2696 3099 2708 3133
rect 2632 3093 2708 3099
rect 2810 3133 2886 3139
rect 2810 3099 2822 3133
rect 2874 3099 2886 3133
rect 2810 3093 2886 3099
rect 2988 3133 3064 3139
rect 2988 3099 3000 3133
rect 3052 3099 3064 3133
rect 2988 3093 3064 3099
rect 3166 3133 3242 3139
rect 3166 3099 3178 3133
rect 3230 3099 3242 3133
rect 3166 3093 3242 3099
rect 3344 3133 3420 3139
rect 3344 3099 3356 3133
rect 3408 3099 3420 3133
rect 852 3023 928 3029
rect 1030 3023 1106 3029
rect 1208 3023 1284 3029
rect 1386 3023 1462 3029
rect 1564 3023 1640 3029
rect 1742 3023 1818 3029
rect 1920 3023 1996 3029
rect 2098 3023 2174 3029
rect 2276 3023 2352 3029
rect 2454 3023 2530 3029
rect 2632 3023 2708 3029
rect 2810 3023 2886 3029
rect 2988 3023 3064 3029
rect 3166 3023 3242 3029
rect 3344 3023 3420 3099
rect 674 2989 686 3023
rect 738 2989 864 3023
rect 916 2989 1042 3023
rect 1094 2989 1220 3023
rect 1272 2989 1398 3023
rect 1450 2989 1576 3023
rect 1628 2989 1754 3023
rect 1806 2989 1932 3023
rect 1984 2989 2110 3023
rect 2162 2989 2288 3023
rect 2340 2989 2466 3023
rect 2518 2989 2644 3023
rect 2696 2989 2822 3023
rect 2874 2989 3000 3023
rect 3052 2989 3178 3023
rect 3230 2989 3356 3023
rect 3408 2989 3420 3023
rect 674 2983 750 2989
rect 852 2983 928 2989
rect 1030 2983 1106 2989
rect 1208 2983 1284 2989
rect 1386 2983 1462 2989
rect 1564 2983 1640 2989
rect 1742 2983 1818 2989
rect 1920 2983 1996 2989
rect 2098 2983 2174 2989
rect 2276 2983 2352 2989
rect 2454 2983 2530 2989
rect 2632 2983 2708 2989
rect 2810 2983 2886 2989
rect 2988 2983 3064 2989
rect 3166 2983 3242 2989
rect 3344 2983 3420 2989
rect 4074 3133 4150 3139
rect 4074 3099 4086 3133
rect 4138 3099 4150 3133
rect 4074 3023 4150 3099
rect 4252 3133 4328 3139
rect 4252 3099 4264 3133
rect 4316 3099 4328 3133
rect 4252 3093 4328 3099
rect 4430 3133 4506 3139
rect 4430 3099 4442 3133
rect 4494 3099 4506 3133
rect 4430 3093 4506 3099
rect 4608 3133 4684 3139
rect 4608 3099 4620 3133
rect 4672 3099 4684 3133
rect 4608 3093 4684 3099
rect 4786 3133 4862 3139
rect 4786 3099 4798 3133
rect 4850 3099 4862 3133
rect 4786 3093 4862 3099
rect 4964 3133 5040 3139
rect 4964 3099 4976 3133
rect 5028 3099 5040 3133
rect 4964 3093 5040 3099
rect 5142 3133 5218 3139
rect 5142 3099 5154 3133
rect 5206 3099 5218 3133
rect 5142 3093 5218 3099
rect 5320 3133 5396 3139
rect 5320 3099 5332 3133
rect 5384 3099 5396 3133
rect 5320 3093 5396 3099
rect 5498 3133 5574 3139
rect 5498 3099 5510 3133
rect 5562 3099 5574 3133
rect 5498 3093 5574 3099
rect 5676 3133 5752 3139
rect 5676 3099 5688 3133
rect 5740 3099 5752 3133
rect 5676 3093 5752 3099
rect 5854 3133 5930 3139
rect 5854 3099 5866 3133
rect 5918 3099 5930 3133
rect 5854 3093 5930 3099
rect 6032 3133 6108 3139
rect 6032 3099 6044 3133
rect 6096 3099 6108 3133
rect 6032 3093 6108 3099
rect 6210 3133 6286 3139
rect 6210 3099 6222 3133
rect 6274 3099 6286 3133
rect 6210 3093 6286 3099
rect 6388 3133 6464 3139
rect 6388 3099 6400 3133
rect 6452 3099 6464 3133
rect 6388 3093 6464 3099
rect 6566 3133 6642 3139
rect 6566 3099 6578 3133
rect 6630 3099 6642 3133
rect 6566 3093 6642 3099
rect 6744 3133 6820 3139
rect 6744 3099 6756 3133
rect 6808 3099 6820 3133
rect 4252 3023 4328 3029
rect 4430 3023 4506 3029
rect 4608 3023 4684 3029
rect 4786 3023 4862 3029
rect 4964 3023 5040 3029
rect 5142 3023 5218 3029
rect 5320 3023 5396 3029
rect 5498 3023 5574 3029
rect 5676 3023 5752 3029
rect 5854 3023 5930 3029
rect 6032 3023 6108 3029
rect 6210 3023 6286 3029
rect 6388 3023 6464 3029
rect 6566 3023 6642 3029
rect 6744 3023 6820 3099
rect 7713 3087 7723 3145
rect 7781 3139 8791 3145
rect 8849 3139 9859 3145
rect 7781 3105 8091 3139
rect 8125 3105 8447 3139
rect 8481 3105 8791 3139
rect 8849 3105 9159 3139
rect 9193 3105 9515 3139
rect 9549 3105 9859 3139
rect 7781 3099 8791 3105
rect 7781 3087 7791 3099
rect 8781 3087 8791 3099
rect 8849 3099 9859 3105
rect 8849 3087 8859 3099
rect 9849 3087 9859 3099
rect 9917 3087 9927 3145
rect 10400 3087 10410 3145
rect 10468 3139 11478 3145
rect 11536 3139 12546 3145
rect 10468 3105 10778 3139
rect 10812 3105 11134 3139
rect 11168 3105 11478 3139
rect 11536 3105 11846 3139
rect 11880 3105 12202 3139
rect 12236 3105 12546 3139
rect 10468 3099 11478 3105
rect 10468 3087 10478 3099
rect 11468 3087 11478 3099
rect 11536 3099 12546 3105
rect 11536 3087 11546 3099
rect 12536 3087 12546 3099
rect 12604 3087 12614 3145
rect 18888 3136 21891 3154
rect 18888 3102 19053 3136
rect 21864 3102 21891 3136
rect 14853 3039 14863 3097
rect 14921 3039 14931 3097
rect 18888 3052 21891 3102
rect 22019 3052 22027 3154
rect 4074 2989 4086 3023
rect 4138 2989 4264 3023
rect 4316 2989 4442 3023
rect 4494 2989 4620 3023
rect 4672 2989 4798 3023
rect 4850 2989 4976 3023
rect 5028 2989 5154 3023
rect 5206 2989 5332 3023
rect 5384 2989 5510 3023
rect 5562 2989 5688 3023
rect 5740 2989 5866 3023
rect 5918 2989 6044 3023
rect 6096 2989 6222 3023
rect 6274 2989 6400 3023
rect 6452 2989 6578 3023
rect 6630 2989 6756 3023
rect 6808 2989 6820 3023
rect 4074 2983 4150 2989
rect 4252 2983 4328 2989
rect 4430 2983 4506 2989
rect 4608 2983 4684 2989
rect 4786 2983 4862 2989
rect 4964 2983 5040 2989
rect 5142 2983 5218 2989
rect 5320 2983 5396 2989
rect 5498 2983 5574 2989
rect 5676 2983 5752 2989
rect 5854 2983 5930 2989
rect 6032 2983 6108 2989
rect 6210 2983 6286 2989
rect 6388 2983 6464 2989
rect 6566 2983 6642 2989
rect 6744 2983 6820 2989
rect 584 2887 594 2945
rect 652 2939 2018 2945
rect 2076 2939 3442 2945
rect 652 2905 962 2939
rect 996 2905 1318 2939
rect 1352 2905 1674 2939
rect 1708 2905 2018 2939
rect 2076 2905 2386 2939
rect 2420 2905 2742 2939
rect 2776 2905 3098 2939
rect 3132 2905 3442 2939
rect 652 2899 2018 2905
rect 652 2887 662 2899
rect 2008 2887 2018 2899
rect 2076 2899 3442 2905
rect 2076 2887 2086 2899
rect 3432 2887 3442 2899
rect 3500 2887 3510 2945
rect 3984 2887 3994 2945
rect 4052 2939 5418 2945
rect 5476 2939 6842 2945
rect 4052 2905 4362 2939
rect 4396 2905 4718 2939
rect 4752 2905 5074 2939
rect 5108 2905 5418 2939
rect 5476 2905 5786 2939
rect 5820 2905 6142 2939
rect 6176 2905 6498 2939
rect 6532 2905 6842 2939
rect 4052 2899 5418 2905
rect 4052 2887 4062 2899
rect 5408 2887 5418 2899
rect 5476 2899 6842 2905
rect 5476 2887 5486 2899
rect 6832 2887 6842 2899
rect 6900 2887 6910 2945
rect 8247 2923 8257 2935
rect 7901 2917 8257 2923
rect 8315 2923 8325 2935
rect 9315 2923 9325 2935
rect 8315 2917 9325 2923
rect 9383 2923 9393 2935
rect 10934 2923 10944 2935
rect 9383 2917 9739 2923
rect 7901 2883 7913 2917
rect 7947 2883 8257 2917
rect 8315 2883 8625 2917
rect 8659 2883 8981 2917
rect 9015 2883 9325 2917
rect 9383 2883 9693 2917
rect 9727 2883 9739 2917
rect 7901 2877 8257 2883
rect 8315 2877 9325 2883
rect 9383 2877 9739 2883
rect 10588 2917 10944 2923
rect 11002 2923 11012 2935
rect 12002 2923 12012 2935
rect 11002 2917 12012 2923
rect 12070 2923 12080 2935
rect 12070 2917 12426 2923
rect 10588 2883 10600 2917
rect 10634 2883 10944 2917
rect 11002 2883 11312 2917
rect 11346 2883 11668 2917
rect 11702 2883 12012 2917
rect 12070 2883 12380 2917
rect 12414 2883 12426 2917
rect 10588 2877 10944 2883
rect 11002 2877 12012 2883
rect 12070 2877 12426 2883
rect 7803 2833 7879 2839
rect 7803 2799 7815 2833
rect 7867 2799 7879 2833
rect 1474 2723 1484 2735
rect 772 2717 1484 2723
rect 1542 2723 1552 2735
rect 2542 2723 2552 2735
rect 1542 2717 2552 2723
rect 2610 2723 2620 2735
rect 4874 2723 4884 2735
rect 2610 2717 3322 2723
rect 772 2683 784 2717
rect 818 2683 1140 2717
rect 1174 2683 1484 2717
rect 1542 2683 1852 2717
rect 1886 2683 2208 2717
rect 2242 2683 2552 2717
rect 2610 2683 2920 2717
rect 2954 2683 3276 2717
rect 3310 2683 3322 2717
rect 772 2677 1484 2683
rect 1542 2677 2552 2683
rect 2610 2677 3322 2683
rect 4172 2717 4884 2723
rect 4942 2723 4952 2735
rect 5942 2723 5952 2736
rect 4942 2717 5952 2723
rect 6010 2723 6020 2736
rect 7803 2723 7879 2799
rect 7981 2833 8057 2839
rect 7981 2799 7993 2833
rect 8045 2799 8057 2833
rect 7981 2793 8057 2799
rect 8159 2833 8235 2839
rect 8159 2799 8171 2833
rect 8223 2799 8235 2833
rect 8159 2793 8235 2799
rect 8337 2833 8413 2839
rect 8337 2799 8349 2833
rect 8401 2799 8413 2833
rect 8337 2793 8413 2799
rect 8515 2833 8591 2839
rect 8515 2799 8527 2833
rect 8579 2799 8591 2833
rect 8515 2793 8591 2799
rect 8693 2833 8769 2839
rect 8693 2799 8705 2833
rect 8757 2799 8769 2833
rect 8693 2793 8769 2799
rect 8871 2833 8947 2839
rect 8871 2799 8883 2833
rect 8935 2799 8947 2833
rect 8871 2793 8947 2799
rect 9049 2833 9125 2839
rect 9049 2799 9061 2833
rect 9113 2799 9125 2833
rect 9049 2793 9125 2799
rect 9227 2833 9303 2839
rect 9227 2799 9239 2833
rect 9291 2799 9303 2833
rect 9227 2793 9303 2799
rect 9405 2833 9481 2839
rect 9405 2799 9417 2833
rect 9469 2799 9481 2833
rect 9405 2793 9481 2799
rect 9583 2833 9659 2839
rect 9583 2799 9595 2833
rect 9647 2799 9659 2833
rect 9583 2793 9659 2799
rect 9761 2833 9837 2839
rect 9761 2799 9773 2833
rect 9825 2799 9837 2833
rect 7981 2723 8057 2729
rect 8159 2723 8235 2729
rect 8337 2723 8413 2729
rect 8515 2723 8591 2729
rect 8693 2723 8769 2729
rect 8871 2723 8947 2729
rect 9049 2723 9125 2729
rect 9227 2723 9303 2729
rect 9405 2723 9481 2729
rect 9583 2723 9659 2729
rect 9761 2723 9837 2799
rect 6010 2717 6722 2723
rect 4172 2683 4184 2717
rect 4218 2683 4540 2717
rect 4574 2683 4884 2717
rect 4942 2683 5252 2717
rect 5286 2683 5608 2717
rect 5642 2683 5952 2717
rect 6010 2683 6320 2717
rect 6354 2683 6676 2717
rect 6710 2683 6722 2717
rect 7803 2689 7815 2723
rect 7867 2689 7993 2723
rect 8045 2689 8171 2723
rect 8223 2689 8349 2723
rect 8401 2689 8527 2723
rect 8579 2689 8705 2723
rect 8757 2689 8883 2723
rect 8935 2689 9061 2723
rect 9113 2689 9239 2723
rect 9291 2689 9417 2723
rect 9469 2689 9595 2723
rect 9647 2689 9773 2723
rect 9825 2689 9837 2723
rect 7803 2683 7879 2689
rect 7981 2683 8057 2689
rect 8159 2683 8235 2689
rect 8337 2683 8413 2689
rect 8515 2683 8591 2689
rect 8693 2683 8769 2689
rect 8871 2683 8947 2689
rect 9049 2683 9125 2689
rect 9227 2683 9303 2689
rect 9405 2683 9481 2689
rect 9583 2683 9659 2689
rect 9761 2683 9837 2689
rect 10490 2833 10566 2839
rect 10490 2799 10502 2833
rect 10554 2799 10566 2833
rect 10490 2723 10566 2799
rect 10668 2833 10744 2839
rect 10668 2799 10680 2833
rect 10732 2799 10744 2833
rect 10668 2793 10744 2799
rect 10846 2833 10922 2839
rect 10846 2799 10858 2833
rect 10910 2799 10922 2833
rect 10846 2793 10922 2799
rect 11024 2833 11100 2839
rect 11024 2799 11036 2833
rect 11088 2799 11100 2833
rect 11024 2793 11100 2799
rect 11202 2833 11278 2839
rect 11202 2799 11214 2833
rect 11266 2799 11278 2833
rect 11202 2793 11278 2799
rect 11380 2833 11456 2839
rect 11380 2799 11392 2833
rect 11444 2799 11456 2833
rect 11380 2793 11456 2799
rect 11558 2833 11634 2839
rect 11558 2799 11570 2833
rect 11622 2799 11634 2833
rect 11558 2793 11634 2799
rect 11736 2833 11812 2839
rect 11736 2799 11748 2833
rect 11800 2799 11812 2833
rect 11736 2793 11812 2799
rect 11914 2833 11990 2839
rect 11914 2799 11926 2833
rect 11978 2799 11990 2833
rect 11914 2793 11990 2799
rect 12092 2833 12168 2839
rect 12092 2799 12104 2833
rect 12156 2799 12168 2833
rect 12092 2793 12168 2799
rect 12270 2833 12346 2839
rect 12270 2799 12282 2833
rect 12334 2799 12346 2833
rect 12270 2793 12346 2799
rect 12448 2833 12524 2839
rect 12448 2799 12460 2833
rect 12512 2799 12524 2833
rect 10668 2723 10744 2729
rect 10846 2723 10922 2729
rect 11024 2723 11100 2729
rect 11202 2723 11278 2729
rect 11380 2723 11456 2729
rect 11558 2723 11634 2729
rect 11736 2723 11812 2729
rect 11914 2723 11990 2729
rect 12092 2723 12168 2729
rect 12270 2723 12346 2729
rect 12448 2723 12524 2799
rect 10490 2689 10502 2723
rect 10554 2689 10680 2723
rect 10732 2689 10858 2723
rect 10910 2689 11036 2723
rect 11088 2689 11214 2723
rect 11266 2689 11392 2723
rect 11444 2689 11570 2723
rect 11622 2689 11748 2723
rect 11800 2689 11926 2723
rect 11978 2689 12104 2723
rect 12156 2689 12282 2723
rect 12334 2689 12460 2723
rect 12512 2689 12524 2723
rect 10490 2683 10566 2689
rect 10668 2683 10744 2689
rect 10846 2683 10922 2689
rect 11024 2683 11100 2689
rect 11202 2683 11278 2689
rect 11380 2683 11456 2689
rect 11558 2683 11634 2689
rect 11736 2683 11812 2689
rect 11914 2683 11990 2689
rect 12092 2683 12168 2689
rect 12270 2683 12346 2689
rect 12448 2683 12524 2689
rect 4172 2677 4884 2683
rect 4942 2678 5952 2683
rect 6010 2678 6722 2683
rect 4942 2677 6722 2678
rect 674 2633 750 2639
rect 674 2599 686 2633
rect 738 2599 750 2633
rect 674 2523 750 2599
rect 852 2633 928 2639
rect 852 2599 864 2633
rect 916 2599 928 2633
rect 852 2593 928 2599
rect 1030 2633 1106 2639
rect 1030 2599 1042 2633
rect 1094 2599 1106 2633
rect 1030 2593 1106 2599
rect 1208 2633 1284 2639
rect 1208 2599 1220 2633
rect 1272 2599 1284 2633
rect 1208 2593 1284 2599
rect 1386 2633 1462 2639
rect 1386 2599 1398 2633
rect 1450 2599 1462 2633
rect 1386 2593 1462 2599
rect 1564 2633 1640 2639
rect 1564 2599 1576 2633
rect 1628 2599 1640 2633
rect 1564 2593 1640 2599
rect 1742 2633 1818 2639
rect 1742 2599 1754 2633
rect 1806 2599 1818 2633
rect 1742 2593 1818 2599
rect 1920 2633 1996 2639
rect 1920 2599 1932 2633
rect 1984 2599 1996 2633
rect 1920 2593 1996 2599
rect 2098 2633 2174 2639
rect 2098 2599 2110 2633
rect 2162 2599 2174 2633
rect 2098 2593 2174 2599
rect 2276 2633 2352 2639
rect 2276 2599 2288 2633
rect 2340 2599 2352 2633
rect 2276 2593 2352 2599
rect 2454 2633 2530 2639
rect 2454 2599 2466 2633
rect 2518 2599 2530 2633
rect 2454 2593 2530 2599
rect 2632 2633 2708 2639
rect 2632 2599 2644 2633
rect 2696 2599 2708 2633
rect 2632 2593 2708 2599
rect 2810 2633 2886 2639
rect 2810 2599 2822 2633
rect 2874 2599 2886 2633
rect 2810 2593 2886 2599
rect 2988 2633 3064 2639
rect 2988 2599 3000 2633
rect 3052 2599 3064 2633
rect 2988 2593 3064 2599
rect 3166 2633 3242 2639
rect 3166 2599 3178 2633
rect 3230 2599 3242 2633
rect 3166 2593 3242 2599
rect 3344 2633 3420 2639
rect 3344 2599 3356 2633
rect 3408 2599 3420 2633
rect 852 2523 928 2529
rect 1030 2523 1106 2529
rect 1208 2523 1284 2529
rect 1386 2523 1462 2529
rect 1564 2523 1640 2529
rect 1742 2523 1818 2529
rect 1920 2523 1996 2529
rect 2098 2523 2174 2529
rect 2276 2523 2352 2529
rect 2454 2523 2530 2529
rect 2632 2523 2708 2529
rect 2810 2523 2886 2529
rect 2988 2523 3064 2529
rect 3166 2523 3242 2529
rect 3344 2523 3420 2599
rect 674 2489 686 2523
rect 738 2489 864 2523
rect 916 2489 1042 2523
rect 1094 2489 1220 2523
rect 1272 2489 1398 2523
rect 1450 2489 1576 2523
rect 1628 2489 1754 2523
rect 1806 2489 1932 2523
rect 1984 2489 2110 2523
rect 2162 2489 2288 2523
rect 2340 2489 2466 2523
rect 2518 2489 2644 2523
rect 2696 2489 2822 2523
rect 2874 2489 3000 2523
rect 3052 2489 3178 2523
rect 3230 2489 3356 2523
rect 3408 2489 3420 2523
rect 674 2483 750 2489
rect 852 2483 928 2489
rect 1030 2483 1106 2489
rect 1208 2483 1284 2489
rect 1386 2483 1462 2489
rect 1564 2483 1640 2489
rect 1742 2483 1818 2489
rect 1920 2483 1996 2489
rect 2098 2483 2174 2489
rect 2276 2483 2352 2489
rect 2454 2483 2530 2489
rect 2632 2483 2708 2489
rect 2810 2483 2886 2489
rect 2988 2483 3064 2489
rect 3166 2483 3242 2489
rect 3344 2483 3420 2489
rect 4074 2633 4150 2639
rect 4074 2599 4086 2633
rect 4138 2599 4150 2633
rect 4074 2523 4150 2599
rect 4252 2633 4328 2639
rect 4252 2599 4264 2633
rect 4316 2599 4328 2633
rect 4252 2593 4328 2599
rect 4430 2633 4506 2639
rect 4430 2599 4442 2633
rect 4494 2599 4506 2633
rect 4430 2593 4506 2599
rect 4608 2633 4684 2639
rect 4608 2599 4620 2633
rect 4672 2599 4684 2633
rect 4608 2593 4684 2599
rect 4786 2633 4862 2639
rect 4786 2599 4798 2633
rect 4850 2599 4862 2633
rect 4786 2593 4862 2599
rect 4964 2633 5040 2639
rect 4964 2599 4976 2633
rect 5028 2599 5040 2633
rect 4964 2593 5040 2599
rect 5142 2633 5218 2639
rect 5142 2599 5154 2633
rect 5206 2599 5218 2633
rect 5142 2593 5218 2599
rect 5320 2633 5396 2639
rect 5320 2599 5332 2633
rect 5384 2599 5396 2633
rect 5320 2593 5396 2599
rect 5498 2633 5574 2639
rect 5498 2599 5510 2633
rect 5562 2599 5574 2633
rect 5498 2593 5574 2599
rect 5676 2633 5752 2639
rect 5676 2599 5688 2633
rect 5740 2599 5752 2633
rect 5676 2593 5752 2599
rect 5854 2633 5930 2639
rect 5854 2599 5866 2633
rect 5918 2599 5930 2633
rect 5854 2593 5930 2599
rect 6032 2633 6108 2639
rect 6032 2599 6044 2633
rect 6096 2599 6108 2633
rect 6032 2593 6108 2599
rect 6210 2633 6286 2639
rect 6210 2599 6222 2633
rect 6274 2599 6286 2633
rect 6210 2593 6286 2599
rect 6388 2633 6464 2639
rect 6388 2599 6400 2633
rect 6452 2599 6464 2633
rect 6388 2593 6464 2599
rect 6566 2633 6642 2639
rect 6566 2599 6578 2633
rect 6630 2599 6642 2633
rect 6566 2593 6642 2599
rect 6744 2633 6820 2639
rect 6744 2599 6756 2633
rect 6808 2599 6820 2633
rect 4252 2523 4328 2529
rect 4430 2523 4506 2529
rect 4608 2523 4684 2529
rect 4786 2523 4862 2529
rect 4964 2523 5040 2529
rect 5142 2523 5218 2529
rect 5320 2523 5396 2529
rect 5498 2523 5574 2529
rect 5676 2523 5752 2529
rect 5854 2523 5930 2529
rect 6032 2523 6108 2529
rect 6210 2523 6286 2529
rect 6388 2523 6464 2529
rect 6566 2523 6642 2529
rect 6744 2523 6820 2599
rect 7713 2587 7723 2645
rect 7781 2639 8791 2645
rect 8849 2639 9859 2645
rect 7781 2605 8091 2639
rect 8125 2605 8447 2639
rect 8481 2605 8791 2639
rect 8849 2605 9159 2639
rect 9193 2605 9515 2639
rect 9549 2605 9859 2639
rect 7781 2599 8791 2605
rect 7781 2587 7791 2599
rect 8781 2587 8791 2599
rect 8849 2599 9859 2605
rect 8849 2587 8859 2599
rect 9849 2587 9859 2599
rect 9917 2587 9927 2645
rect 10400 2587 10410 2645
rect 10468 2639 11478 2645
rect 11536 2639 12546 2645
rect 10468 2605 10778 2639
rect 10812 2605 11134 2639
rect 11168 2605 11478 2639
rect 11536 2605 11846 2639
rect 11880 2605 12202 2639
rect 12236 2605 12546 2639
rect 10468 2599 11478 2605
rect 10468 2587 10478 2599
rect 11468 2587 11478 2599
rect 11536 2599 12546 2605
rect 11536 2587 11546 2599
rect 12536 2587 12546 2599
rect 12604 2587 12614 2645
rect 14863 2628 14921 3039
rect 17238 2694 17272 2712
rect 16640 2688 16716 2694
rect 16818 2688 16894 2694
rect 16996 2688 17072 2694
rect 17174 2688 17272 2694
rect 16640 2654 16652 2688
rect 16704 2654 16830 2688
rect 16882 2654 17008 2688
rect 17060 2654 17186 2688
rect 17238 2654 17272 2688
rect 17330 2694 17364 2712
rect 17330 2688 17428 2694
rect 17530 2688 17606 2694
rect 17708 2688 17784 2694
rect 17886 2688 17962 2694
rect 18064 2688 18140 2694
rect 17330 2654 17364 2688
rect 17416 2654 17542 2688
rect 17594 2654 17720 2688
rect 17772 2654 17898 2688
rect 17950 2654 18076 2688
rect 18128 2654 18140 2688
rect 16640 2648 16716 2654
rect 16818 2648 16894 2654
rect 16996 2648 17072 2654
rect 17174 2648 17250 2654
rect 17352 2648 17428 2654
rect 17530 2648 17606 2654
rect 17708 2648 17784 2654
rect 17886 2648 17962 2654
rect 18064 2648 18140 2654
rect 13670 2622 13894 2628
rect 13670 2596 13756 2622
rect 13666 2588 13756 2596
rect 13808 2588 13894 2622
rect 4074 2489 4086 2523
rect 4138 2489 4264 2523
rect 4316 2489 4442 2523
rect 4494 2489 4620 2523
rect 4672 2489 4798 2523
rect 4850 2489 4976 2523
rect 5028 2489 5154 2523
rect 5206 2489 5332 2523
rect 5384 2489 5510 2523
rect 5562 2489 5688 2523
rect 5740 2489 5866 2523
rect 5918 2489 6044 2523
rect 6096 2489 6222 2523
rect 6274 2489 6400 2523
rect 6452 2489 6578 2523
rect 6630 2489 6756 2523
rect 6808 2489 6820 2523
rect 4074 2483 4150 2489
rect 4252 2483 4328 2489
rect 4430 2483 4506 2489
rect 4608 2483 4684 2489
rect 4786 2483 4862 2489
rect 4964 2483 5040 2489
rect 5142 2483 5218 2489
rect 5320 2483 5396 2489
rect 5498 2483 5574 2489
rect 5676 2483 5752 2489
rect 5854 2483 5930 2489
rect 6032 2483 6108 2489
rect 6210 2483 6286 2489
rect 6388 2483 6464 2489
rect 6566 2483 6642 2489
rect 6744 2483 6820 2489
rect 13666 2582 13894 2588
rect 14036 2622 14112 2628
rect 14328 2622 14404 2628
rect 14620 2622 14696 2628
rect 14863 2622 14988 2628
rect 15204 2622 15280 2628
rect 15496 2626 15572 2628
rect 15422 2622 15646 2626
rect 14036 2588 14048 2622
rect 14100 2588 14340 2622
rect 14392 2588 14632 2622
rect 14684 2588 14924 2622
rect 14976 2588 15216 2622
rect 15268 2588 15348 2622
rect 14036 2582 14112 2588
rect 13666 2538 13716 2582
rect 584 2387 594 2445
rect 652 2439 2018 2445
rect 2076 2439 3442 2445
rect 652 2405 962 2439
rect 996 2405 1318 2439
rect 1352 2405 1674 2439
rect 1708 2405 2018 2439
rect 2076 2405 2386 2439
rect 2420 2405 2742 2439
rect 2776 2405 3098 2439
rect 3132 2405 3442 2439
rect 652 2399 2018 2405
rect 652 2387 662 2399
rect 2008 2387 2018 2399
rect 2076 2399 3442 2405
rect 2076 2387 2086 2399
rect 3432 2387 3442 2399
rect 3500 2387 3510 2445
rect 3984 2387 3994 2445
rect 4052 2439 5418 2445
rect 5476 2439 6842 2445
rect 4052 2405 4362 2439
rect 4396 2405 4718 2439
rect 4752 2405 5074 2439
rect 5108 2405 5418 2439
rect 5476 2405 5786 2439
rect 5820 2405 6142 2439
rect 6176 2405 6498 2439
rect 6532 2405 6842 2439
rect 4052 2399 5418 2405
rect 4052 2387 4062 2399
rect 5408 2387 5418 2399
rect 5476 2399 6842 2405
rect 5476 2387 5486 2399
rect 6832 2387 6842 2399
rect 6900 2387 6910 2445
rect 8247 2423 8257 2435
rect 7901 2417 8257 2423
rect 8315 2423 8325 2435
rect 8588 2426 8800 2431
rect 8588 2423 8609 2426
rect 7901 2383 7913 2417
rect 7947 2383 8257 2417
rect 7901 2377 8257 2383
rect 8315 2377 8609 2423
rect 8800 2423 8810 2426
rect 9315 2423 9325 2435
rect 8800 2417 9325 2423
rect 9383 2423 9393 2435
rect 10934 2423 10944 2435
rect 9383 2417 9739 2423
rect 8800 2383 8981 2417
rect 9015 2383 9325 2417
rect 9383 2383 9693 2417
rect 9727 2383 9739 2417
rect 8588 2373 8609 2377
rect 8800 2377 9325 2383
rect 9383 2377 9739 2383
rect 10588 2417 10944 2423
rect 11002 2423 11012 2435
rect 11646 2427 11724 2435
rect 11544 2426 11756 2427
rect 11536 2423 11546 2426
rect 11002 2417 11546 2423
rect 11752 2423 11762 2426
rect 12002 2423 12012 2435
rect 10588 2383 10600 2417
rect 10634 2383 10944 2417
rect 11002 2383 11312 2417
rect 11346 2383 11546 2417
rect 10588 2377 10944 2383
rect 11002 2377 11546 2383
rect 8800 2373 8810 2377
rect 11536 2368 11546 2377
rect 11752 2377 12012 2423
rect 12070 2423 12080 2435
rect 12070 2417 12426 2423
rect 12070 2383 12380 2417
rect 12414 2383 12426 2417
rect 12070 2377 12426 2383
rect 11752 2368 11762 2377
rect 7803 2333 7879 2339
rect 7803 2299 7815 2333
rect 7867 2299 7879 2333
rect 7803 2293 7879 2299
rect 7981 2333 8057 2339
rect 7981 2299 7993 2333
rect 8045 2299 8057 2333
rect 7981 2293 8057 2299
rect 8159 2333 8235 2339
rect 8159 2299 8171 2333
rect 8223 2299 8235 2333
rect 8159 2293 8235 2299
rect 8337 2333 8413 2339
rect 8337 2299 8349 2333
rect 8401 2299 8413 2333
rect 8337 2293 8413 2299
rect 8515 2333 8591 2339
rect 8515 2299 8527 2333
rect 8579 2299 8591 2333
rect 8515 2293 8591 2299
rect 8693 2333 8769 2339
rect 8693 2299 8705 2333
rect 8757 2299 8769 2333
rect 8693 2293 8769 2299
rect 8871 2333 8947 2339
rect 8871 2299 8883 2333
rect 8935 2299 8947 2333
rect 8871 2293 8947 2299
rect 9049 2333 9125 2339
rect 9049 2299 9061 2333
rect 9113 2299 9125 2333
rect 9049 2293 9125 2299
rect 9227 2333 9303 2339
rect 9227 2299 9239 2333
rect 9291 2299 9303 2333
rect 9227 2293 9303 2299
rect 9405 2333 9481 2339
rect 9405 2299 9417 2333
rect 9469 2299 9481 2333
rect 9405 2293 9481 2299
rect 9583 2333 9659 2339
rect 9583 2299 9595 2333
rect 9647 2299 9659 2333
rect 9583 2293 9659 2299
rect 9761 2333 9837 2339
rect 9761 2299 9773 2333
rect 9825 2299 9837 2333
rect 9761 2293 9837 2299
rect 10490 2333 10566 2339
rect 10490 2299 10502 2333
rect 10554 2299 10566 2333
rect 10490 2293 10566 2299
rect 10668 2333 10744 2339
rect 10668 2299 10680 2333
rect 10732 2299 10744 2333
rect 10668 2293 10744 2299
rect 10846 2333 10922 2339
rect 10846 2299 10858 2333
rect 10910 2299 10922 2333
rect 10846 2293 10922 2299
rect 11024 2333 11100 2339
rect 11024 2299 11036 2333
rect 11088 2299 11100 2333
rect 11024 2293 11100 2299
rect 11202 2333 11278 2339
rect 11202 2299 11214 2333
rect 11266 2299 11278 2333
rect 11202 2293 11278 2299
rect 11380 2333 11456 2339
rect 11380 2299 11392 2333
rect 11444 2299 11456 2333
rect 11380 2293 11456 2299
rect 11558 2333 11634 2339
rect 11558 2299 11570 2333
rect 11622 2299 11634 2333
rect 11558 2293 11634 2299
rect 11736 2333 11812 2339
rect 11736 2299 11748 2333
rect 11800 2299 11812 2333
rect 11736 2293 11812 2299
rect 11914 2333 11990 2339
rect 11914 2299 11926 2333
rect 11978 2299 11990 2333
rect 11914 2293 11990 2299
rect 12092 2333 12168 2339
rect 12092 2299 12104 2333
rect 12156 2299 12168 2333
rect 12092 2293 12168 2299
rect 12270 2333 12346 2339
rect 12270 2299 12282 2333
rect 12334 2299 12346 2333
rect 12270 2293 12346 2299
rect 12448 2333 12524 2339
rect 12448 2299 12460 2333
rect 12512 2299 12524 2333
rect 12448 2293 12524 2299
rect 13666 2282 13676 2538
rect 13710 2282 13716 2538
rect 13666 2238 13716 2282
rect 13848 2538 13894 2582
rect 14146 2550 14180 2588
rect 14328 2582 14404 2588
rect 14620 2582 14696 2588
rect 14912 2582 14988 2588
rect 15204 2582 15280 2588
rect 15314 2550 15348 2588
rect 15422 2588 15508 2622
rect 15560 2588 15646 2622
rect 16738 2608 17420 2610
rect 15422 2580 15646 2588
rect 13848 2282 13854 2538
rect 13888 2282 13894 2538
rect 13848 2238 13894 2282
rect 13962 2538 14008 2550
rect 14140 2538 14186 2550
rect 14254 2538 14300 2550
rect 14432 2538 14478 2550
rect 14546 2538 14592 2550
rect 14724 2538 14770 2550
rect 14838 2538 14884 2550
rect 15016 2538 15062 2550
rect 15130 2538 15176 2550
rect 15308 2538 15354 2550
rect 15422 2538 15468 2580
rect 13962 2282 13968 2538
rect 14002 2282 14008 2538
rect 14124 2480 14134 2538
rect 14192 2480 14202 2538
rect 13962 2270 14008 2282
rect 14140 2282 14146 2480
rect 14180 2282 14186 2480
rect 14140 2270 14186 2282
rect 14254 2282 14260 2538
rect 14294 2282 14300 2538
rect 14416 2480 14426 2538
rect 14484 2480 14494 2538
rect 14254 2270 14300 2282
rect 14432 2282 14438 2480
rect 14472 2282 14478 2480
rect 14432 2270 14478 2282
rect 14546 2282 14552 2538
rect 14586 2282 14592 2538
rect 14708 2480 14718 2538
rect 14776 2480 14786 2538
rect 14546 2270 14592 2282
rect 14724 2282 14730 2480
rect 14764 2282 14770 2480
rect 14724 2270 14770 2282
rect 14838 2282 14844 2538
rect 14878 2282 14884 2538
rect 15000 2480 15010 2538
rect 15068 2480 15078 2538
rect 14838 2270 14884 2282
rect 15016 2282 15022 2480
rect 15056 2282 15062 2480
rect 15016 2270 15062 2282
rect 15130 2282 15136 2538
rect 15170 2282 15176 2538
rect 15292 2480 15302 2538
rect 15360 2480 15370 2538
rect 15130 2270 15176 2282
rect 15308 2282 15314 2480
rect 15348 2282 15354 2480
rect 15308 2270 15354 2282
rect 15422 2282 15428 2538
rect 15462 2282 15468 2538
rect 1474 2223 1484 2235
rect 772 2217 1484 2223
rect 1542 2223 1552 2235
rect 2542 2223 2552 2235
rect 1542 2217 2552 2223
rect 2610 2223 2620 2235
rect 4874 2223 4884 2235
rect 2610 2217 3322 2223
rect 772 2183 784 2217
rect 818 2183 1140 2217
rect 1174 2183 1484 2217
rect 1542 2183 1852 2217
rect 1886 2183 2208 2217
rect 2242 2183 2552 2217
rect 2610 2183 2920 2217
rect 2954 2183 3276 2217
rect 3310 2183 3322 2217
rect 772 2177 1484 2183
rect 1542 2177 2552 2183
rect 2610 2177 3322 2183
rect 4172 2217 4884 2223
rect 4942 2223 4952 2235
rect 5942 2223 5952 2235
rect 4942 2217 5952 2223
rect 6010 2223 6020 2235
rect 13666 2232 13894 2238
rect 6010 2217 6722 2223
rect 4172 2183 4184 2217
rect 4218 2183 4540 2217
rect 4574 2183 4884 2217
rect 4942 2183 5252 2217
rect 5286 2183 5608 2217
rect 5642 2183 5952 2217
rect 6010 2183 6320 2217
rect 6354 2183 6676 2217
rect 6710 2183 6722 2217
rect 4172 2177 4884 2183
rect 4942 2177 5952 2183
rect 6010 2177 6722 2183
rect 13666 2198 13756 2232
rect 13808 2198 13894 2232
rect 13666 2192 13894 2198
rect 674 2133 750 2139
rect 674 2099 686 2133
rect 738 2099 750 2133
rect 674 2023 750 2099
rect 852 2133 928 2139
rect 852 2099 864 2133
rect 916 2099 928 2133
rect 852 2093 928 2099
rect 1030 2133 1106 2139
rect 1030 2099 1042 2133
rect 1094 2099 1106 2133
rect 1030 2093 1106 2099
rect 1208 2133 1284 2139
rect 1208 2099 1220 2133
rect 1272 2099 1284 2133
rect 1208 2093 1284 2099
rect 1386 2133 1462 2139
rect 1386 2099 1398 2133
rect 1450 2099 1462 2133
rect 1386 2093 1462 2099
rect 1564 2133 1640 2139
rect 1564 2099 1576 2133
rect 1628 2099 1640 2133
rect 1564 2093 1640 2099
rect 1742 2133 1818 2139
rect 1742 2099 1754 2133
rect 1806 2099 1818 2133
rect 1742 2093 1818 2099
rect 1920 2133 1996 2139
rect 1920 2099 1932 2133
rect 1984 2099 1996 2133
rect 1920 2093 1996 2099
rect 2098 2133 2174 2139
rect 2098 2099 2110 2133
rect 2162 2099 2174 2133
rect 2098 2093 2174 2099
rect 2276 2133 2352 2139
rect 2276 2099 2288 2133
rect 2340 2099 2352 2133
rect 2276 2093 2352 2099
rect 2454 2133 2530 2139
rect 2454 2099 2466 2133
rect 2518 2099 2530 2133
rect 2454 2093 2530 2099
rect 2632 2133 2708 2139
rect 2632 2099 2644 2133
rect 2696 2099 2708 2133
rect 2632 2093 2708 2099
rect 2810 2133 2886 2139
rect 2810 2099 2822 2133
rect 2874 2099 2886 2133
rect 2810 2093 2886 2099
rect 2988 2133 3064 2139
rect 2988 2099 3000 2133
rect 3052 2099 3064 2133
rect 2988 2093 3064 2099
rect 3166 2133 3242 2139
rect 3166 2099 3178 2133
rect 3230 2099 3242 2133
rect 3166 2093 3242 2099
rect 3344 2133 3420 2139
rect 3344 2099 3356 2133
rect 3408 2099 3420 2133
rect 852 2023 928 2029
rect 1030 2023 1106 2029
rect 1208 2023 1284 2029
rect 1386 2023 1462 2029
rect 1564 2023 1640 2029
rect 1742 2023 1818 2029
rect 1920 2023 1996 2029
rect 2098 2023 2174 2029
rect 2276 2023 2352 2029
rect 2454 2023 2530 2029
rect 2632 2023 2708 2029
rect 2810 2023 2886 2029
rect 2988 2023 3064 2029
rect 3166 2023 3242 2029
rect 3344 2023 3420 2099
rect 674 1989 686 2023
rect 738 1989 864 2023
rect 916 1989 1042 2023
rect 1094 1989 1220 2023
rect 1272 1989 1398 2023
rect 1450 1989 1576 2023
rect 1628 1989 1754 2023
rect 1806 1989 1932 2023
rect 1984 1989 2110 2023
rect 2162 1989 2288 2023
rect 2340 1989 2466 2023
rect 2518 1989 2644 2023
rect 2696 1989 2822 2023
rect 2874 1989 3000 2023
rect 3052 1989 3178 2023
rect 3230 1989 3356 2023
rect 3408 1989 3420 2023
rect 674 1983 750 1989
rect 852 1983 928 1989
rect 1030 1983 1106 1989
rect 1208 1983 1284 1989
rect 1386 1983 1462 1989
rect 1564 1983 1640 1989
rect 1742 1983 1818 1989
rect 1920 1983 1996 1989
rect 2098 1983 2174 1989
rect 2276 1983 2352 1989
rect 2454 1983 2530 1989
rect 2632 1983 2708 1989
rect 2810 1983 2886 1989
rect 2988 1983 3064 1989
rect 3166 1983 3242 1989
rect 3344 1983 3420 1989
rect 4074 2133 4150 2139
rect 4074 2099 4086 2133
rect 4138 2099 4150 2133
rect 4074 2023 4150 2099
rect 4252 2133 4328 2139
rect 4252 2099 4264 2133
rect 4316 2099 4328 2133
rect 4252 2093 4328 2099
rect 4430 2133 4506 2139
rect 4430 2099 4442 2133
rect 4494 2099 4506 2133
rect 4430 2093 4506 2099
rect 4608 2133 4684 2139
rect 4608 2099 4620 2133
rect 4672 2099 4684 2133
rect 4608 2093 4684 2099
rect 4786 2133 4862 2139
rect 4786 2099 4798 2133
rect 4850 2099 4862 2133
rect 4786 2093 4862 2099
rect 4964 2133 5040 2139
rect 4964 2099 4976 2133
rect 5028 2099 5040 2133
rect 4964 2093 5040 2099
rect 5142 2133 5218 2139
rect 5142 2099 5154 2133
rect 5206 2099 5218 2133
rect 5142 2093 5218 2099
rect 5320 2133 5396 2139
rect 5320 2099 5332 2133
rect 5384 2099 5396 2133
rect 5320 2093 5396 2099
rect 5498 2133 5574 2139
rect 5498 2099 5510 2133
rect 5562 2099 5574 2133
rect 5498 2093 5574 2099
rect 5676 2133 5752 2139
rect 5676 2099 5688 2133
rect 5740 2099 5752 2133
rect 5676 2093 5752 2099
rect 5854 2133 5930 2139
rect 5854 2099 5866 2133
rect 5918 2099 5930 2133
rect 5854 2093 5930 2099
rect 6032 2133 6108 2139
rect 6032 2099 6044 2133
rect 6096 2099 6108 2133
rect 6032 2093 6108 2099
rect 6210 2133 6286 2139
rect 6210 2099 6222 2133
rect 6274 2099 6286 2133
rect 6210 2093 6286 2099
rect 6388 2133 6464 2139
rect 6388 2099 6400 2133
rect 6452 2099 6464 2133
rect 6388 2093 6464 2099
rect 6566 2133 6642 2139
rect 6566 2099 6578 2133
rect 6630 2099 6642 2133
rect 6566 2093 6642 2099
rect 6744 2133 6820 2139
rect 6744 2099 6756 2133
rect 6808 2099 6820 2133
rect 4252 2023 4328 2029
rect 4430 2023 4506 2029
rect 4608 2023 4684 2029
rect 4786 2023 4862 2029
rect 4964 2023 5040 2029
rect 5142 2023 5218 2029
rect 5320 2023 5396 2029
rect 5498 2023 5574 2029
rect 5676 2023 5752 2029
rect 5854 2023 5930 2029
rect 6032 2023 6108 2029
rect 6210 2023 6286 2029
rect 6388 2023 6464 2029
rect 6566 2023 6642 2029
rect 6744 2023 6820 2099
rect 13666 2132 13712 2192
rect 13848 2132 13894 2192
rect 13666 2124 13894 2132
rect 13666 2090 13756 2124
rect 13808 2090 13894 2124
rect 13666 2086 13894 2090
rect 13666 2052 13712 2086
rect 13744 2084 13820 2086
rect 13666 2040 13716 2052
rect 4074 1989 4086 2023
rect 4138 1989 4264 2023
rect 4316 1989 4442 2023
rect 4494 1989 4620 2023
rect 4672 1989 4798 2023
rect 4850 1989 4976 2023
rect 5028 1989 5154 2023
rect 5206 1989 5332 2023
rect 5384 1989 5510 2023
rect 5562 1989 5688 2023
rect 5740 1989 5866 2023
rect 5918 1989 6044 2023
rect 6096 1989 6222 2023
rect 6274 1989 6400 2023
rect 6452 1989 6578 2023
rect 6630 1989 6756 2023
rect 6808 1989 6820 2023
rect 4074 1983 4150 1989
rect 4252 1983 4328 1989
rect 4430 1983 4506 1989
rect 4608 1983 4684 1989
rect 4786 1983 4862 1989
rect 4964 1983 5040 1989
rect 5142 1983 5218 1989
rect 5320 1983 5396 1989
rect 5498 1983 5574 1989
rect 5676 1983 5752 1989
rect 5854 1983 5930 1989
rect 6032 1983 6108 1989
rect 6210 1983 6286 1989
rect 6388 1983 6464 1989
rect 6566 1983 6642 1989
rect 6744 1983 6820 1989
rect 7803 2023 7879 2029
rect 7981 2023 8057 2029
rect 8159 2023 8235 2029
rect 8337 2023 8413 2029
rect 8515 2023 8591 2029
rect 8693 2023 8769 2029
rect 8871 2023 8947 2029
rect 9049 2023 9125 2029
rect 9227 2023 9303 2029
rect 9405 2023 9481 2029
rect 9583 2023 9659 2029
rect 9761 2023 9837 2029
rect 7803 1989 7815 2023
rect 7867 1989 7993 2023
rect 8045 1989 8171 2023
rect 8223 1989 8349 2023
rect 8401 1989 8527 2023
rect 8579 1989 8705 2023
rect 8757 1989 8883 2023
rect 8935 1989 9061 2023
rect 9113 1989 9239 2023
rect 9291 1989 9417 2023
rect 9469 1989 9595 2023
rect 9647 1989 9773 2023
rect 9825 1989 9837 2023
rect 7803 1983 7879 1989
rect 7981 1983 8057 1989
rect 8159 1983 8235 1989
rect 8337 1983 8413 1989
rect 8515 1983 8591 1989
rect 8693 1983 8769 1989
rect 8871 1983 8947 1989
rect 9049 1983 9125 1989
rect 9227 1983 9303 1989
rect 9405 1983 9481 1989
rect 9583 1983 9659 1989
rect 9761 1983 9837 1989
rect 10490 2023 10566 2029
rect 10668 2023 10744 2029
rect 10846 2023 10922 2029
rect 11024 2023 11100 2029
rect 11202 2023 11278 2029
rect 11380 2023 11456 2029
rect 11558 2023 11634 2029
rect 11736 2023 11812 2029
rect 11914 2023 11990 2029
rect 12092 2023 12168 2029
rect 12270 2023 12346 2029
rect 12448 2023 12524 2029
rect 10490 1989 10502 2023
rect 10554 1989 10680 2023
rect 10732 1989 10858 2023
rect 10910 1989 11036 2023
rect 11088 1989 11214 2023
rect 11266 1989 11392 2023
rect 11444 1989 11570 2023
rect 11622 1989 11748 2023
rect 11800 1989 11926 2023
rect 11978 1989 12104 2023
rect 12156 1989 12282 2023
rect 12334 1989 12460 2023
rect 12512 1989 12524 2023
rect 10490 1983 10566 1989
rect 10668 1983 10744 1989
rect 10846 1983 10922 1989
rect 11024 1983 11100 1989
rect 11202 1983 11278 1989
rect 11380 1983 11456 1989
rect 11558 1983 11634 1989
rect 11736 1983 11812 1989
rect 11914 1983 11990 1989
rect 12092 1983 12168 1989
rect 12270 1983 12346 1989
rect 12448 1983 12524 1989
rect 8583 1945 8593 1946
rect 584 1887 594 1945
rect 652 1939 2018 1945
rect 2076 1939 3442 1945
rect 652 1905 962 1939
rect 996 1905 1318 1939
rect 1352 1905 1674 1939
rect 1708 1905 2018 1939
rect 2076 1905 2386 1939
rect 2420 1905 2742 1939
rect 2776 1905 3098 1939
rect 3132 1905 3442 1939
rect 652 1899 2018 1905
rect 652 1887 662 1899
rect 2008 1887 2018 1899
rect 2076 1899 3442 1905
rect 2076 1887 2086 1899
rect 3432 1887 3442 1899
rect 3500 1887 3510 1945
rect 3984 1887 3994 1945
rect 4052 1939 5418 1945
rect 5476 1939 6842 1945
rect 4052 1905 4362 1939
rect 4396 1905 4718 1939
rect 4752 1905 5074 1939
rect 5108 1905 5418 1939
rect 5476 1905 5786 1939
rect 5820 1905 6142 1939
rect 6176 1905 6498 1939
rect 6532 1905 6842 1939
rect 4052 1899 5418 1905
rect 4052 1887 4062 1899
rect 5408 1887 5418 1899
rect 5476 1899 6842 1905
rect 5476 1887 5486 1899
rect 6832 1887 6842 1899
rect 6900 1887 6910 1945
rect 7713 1887 7723 1945
rect 7781 1939 8593 1945
rect 8857 1945 8867 1946
rect 11492 1945 11502 1946
rect 11708 1945 11718 1946
rect 8857 1939 9859 1945
rect 7781 1905 8091 1939
rect 8125 1905 8447 1939
rect 8481 1905 8593 1939
rect 8857 1905 9159 1939
rect 9193 1905 9515 1939
rect 9549 1905 9859 1939
rect 7781 1899 8593 1905
rect 7781 1887 7791 1899
rect 8583 1887 8593 1899
rect 8857 1899 9859 1905
rect 8857 1887 8867 1899
rect 9849 1887 9859 1899
rect 9917 1887 9927 1945
rect 10400 1887 10410 1945
rect 10468 1939 11478 1945
rect 11708 1939 12546 1945
rect 10468 1905 10778 1939
rect 10812 1905 11134 1939
rect 11168 1905 11478 1939
rect 11708 1905 11846 1939
rect 11880 1905 12202 1939
rect 12236 1905 12546 1939
rect 10468 1899 11478 1905
rect 10468 1887 10478 1899
rect 11468 1887 11478 1899
rect 11708 1899 12546 1905
rect 11708 1887 11745 1899
rect 12536 1887 12546 1899
rect 12604 1887 12614 1945
rect 11492 1886 11502 1887
rect 11708 1886 11718 1887
rect 13666 1784 13676 2040
rect 13710 1784 13716 2040
rect 13666 1772 13716 1784
rect 13848 2040 13894 2086
rect 13968 2052 14002 2270
rect 14036 2232 14112 2238
rect 14036 2198 14048 2232
rect 14100 2198 14112 2232
rect 14036 2192 14112 2198
rect 14057 2130 14091 2192
rect 14036 2124 14112 2130
rect 14036 2090 14048 2124
rect 14100 2090 14112 2124
rect 14036 2084 14112 2090
rect 14260 2052 14294 2270
rect 14328 2232 14404 2238
rect 14328 2198 14340 2232
rect 14392 2198 14404 2232
rect 14328 2192 14404 2198
rect 14348 2130 14382 2192
rect 14328 2124 14404 2130
rect 14328 2090 14340 2124
rect 14392 2090 14404 2124
rect 14328 2084 14404 2090
rect 14552 2052 14586 2270
rect 14620 2232 14696 2238
rect 14620 2198 14632 2232
rect 14684 2198 14696 2232
rect 14620 2192 14696 2198
rect 14641 2130 14675 2192
rect 14620 2124 14696 2130
rect 14620 2090 14632 2124
rect 14684 2090 14696 2124
rect 14620 2084 14696 2090
rect 14844 2052 14878 2270
rect 14912 2232 14988 2238
rect 14912 2198 14924 2232
rect 14976 2198 14988 2232
rect 14912 2192 14988 2198
rect 14933 2130 14967 2192
rect 14912 2124 14988 2130
rect 14912 2090 14924 2124
rect 14976 2090 14988 2124
rect 14912 2084 14988 2090
rect 15136 2052 15170 2270
rect 15422 2238 15468 2282
rect 15600 2538 15646 2580
rect 16728 2550 16738 2608
rect 16796 2604 17420 2608
rect 17535 2604 18162 2610
rect 16796 2570 17106 2604
rect 17140 2570 17420 2604
rect 17535 2570 17818 2604
rect 17852 2570 18162 2604
rect 16796 2564 17420 2570
rect 16796 2550 16806 2564
rect 15600 2282 15606 2538
rect 15640 2282 15646 2538
rect 17410 2514 17420 2564
rect 17535 2564 18162 2570
rect 17535 2514 17545 2564
rect 18152 2552 18162 2564
rect 18220 2552 18230 2610
rect 16550 2342 16560 2400
rect 16618 2388 16628 2400
rect 17974 2388 17984 2400
rect 16618 2382 17984 2388
rect 16618 2348 16928 2382
rect 16962 2348 17284 2382
rect 17318 2348 17640 2382
rect 17674 2348 17984 2382
rect 16618 2342 17984 2348
rect 18042 2342 18052 2400
rect 15600 2238 15646 2282
rect 15204 2232 15280 2238
rect 15204 2198 15216 2232
rect 15268 2198 15280 2232
rect 15204 2192 15280 2198
rect 15422 2232 15646 2238
rect 15422 2198 15508 2232
rect 15560 2198 15646 2232
rect 15422 2192 15646 2198
rect 15225 2130 15259 2192
rect 15422 2130 15468 2192
rect 15600 2130 15646 2192
rect 16640 2299 16716 2304
rect 16640 2298 16722 2299
rect 16818 2298 16894 2304
rect 16996 2298 17072 2304
rect 17174 2298 17250 2304
rect 17352 2298 17428 2304
rect 17530 2298 17606 2304
rect 17708 2298 17784 2304
rect 17886 2298 17962 2304
rect 18064 2298 18140 2304
rect 16640 2264 16652 2298
rect 16704 2264 16830 2298
rect 16882 2264 17008 2298
rect 17060 2264 17186 2298
rect 17238 2283 17364 2298
rect 17238 2264 17243 2283
rect 16640 2188 16722 2264
rect 16818 2258 16894 2264
rect 16996 2258 17072 2264
rect 17174 2258 17243 2264
rect 17233 2194 17243 2258
rect 16818 2188 16894 2194
rect 16996 2188 17072 2194
rect 17174 2188 17243 2194
rect 16640 2154 16652 2188
rect 16704 2154 16830 2188
rect 16882 2154 17008 2188
rect 17060 2154 17186 2188
rect 17238 2166 17243 2188
rect 17361 2264 17364 2283
rect 17416 2264 17542 2298
rect 17594 2264 17720 2298
rect 17772 2264 17898 2298
rect 17950 2264 18076 2298
rect 18128 2264 18140 2298
rect 17361 2258 17428 2264
rect 17530 2258 17606 2264
rect 17708 2258 17784 2264
rect 17886 2258 17962 2264
rect 17361 2194 17371 2258
rect 17361 2188 17428 2194
rect 17530 2188 17606 2194
rect 17708 2188 17784 2194
rect 17886 2188 17962 2194
rect 18064 2188 18140 2264
rect 17361 2166 17364 2188
rect 17238 2154 17364 2166
rect 17416 2154 17542 2188
rect 17594 2154 17720 2188
rect 17772 2154 17898 2188
rect 17950 2154 18076 2188
rect 18128 2154 18140 2188
rect 16640 2148 16716 2154
rect 16818 2148 16894 2154
rect 16996 2148 17072 2154
rect 17174 2148 17250 2154
rect 17352 2148 17428 2154
rect 17530 2148 17606 2154
rect 17708 2148 17784 2154
rect 17886 2148 17962 2154
rect 18064 2148 18140 2154
rect 15204 2124 15280 2130
rect 15204 2090 15216 2124
rect 15268 2090 15280 2124
rect 15204 2084 15280 2090
rect 15422 2124 15646 2130
rect 15422 2090 15508 2124
rect 15560 2090 15646 2124
rect 15422 2084 15646 2090
rect 13848 1784 13854 2040
rect 13888 1784 13894 2040
rect 1474 1723 1484 1735
rect 772 1717 1484 1723
rect 1542 1723 1552 1735
rect 2542 1723 2552 1735
rect 1542 1717 2552 1723
rect 2610 1723 2620 1735
rect 4874 1723 4884 1735
rect 2610 1717 3322 1723
rect 772 1683 784 1717
rect 818 1683 1140 1717
rect 1174 1683 1484 1717
rect 1542 1683 1852 1717
rect 1886 1683 2208 1717
rect 2242 1683 2552 1717
rect 2610 1683 2920 1717
rect 2954 1683 3276 1717
rect 3310 1683 3322 1717
rect 772 1677 1484 1683
rect 1542 1677 2552 1683
rect 2610 1677 3322 1683
rect 4172 1717 4884 1723
rect 4942 1723 4952 1735
rect 5942 1723 5952 1735
rect 4942 1717 5952 1723
rect 6010 1723 6020 1735
rect 8247 1723 8257 1735
rect 6010 1717 6722 1723
rect 4172 1683 4184 1717
rect 4218 1683 4540 1717
rect 4574 1683 4884 1717
rect 4942 1683 5252 1717
rect 5286 1683 5608 1717
rect 5642 1683 5952 1717
rect 6010 1683 6320 1717
rect 6354 1683 6676 1717
rect 6710 1683 6722 1717
rect 4172 1677 4884 1683
rect 4942 1677 5952 1683
rect 6010 1677 6722 1683
rect 7901 1717 8257 1723
rect 8315 1723 8325 1735
rect 9315 1723 9325 1735
rect 8315 1717 9325 1723
rect 9383 1723 9393 1735
rect 10934 1723 10944 1735
rect 9383 1717 9739 1723
rect 7901 1683 7913 1717
rect 7947 1683 8257 1717
rect 8315 1683 8625 1717
rect 8659 1683 8981 1717
rect 9015 1683 9325 1717
rect 9383 1683 9693 1717
rect 9727 1683 9739 1717
rect 7901 1677 8257 1683
rect 8315 1677 9325 1683
rect 9383 1677 9739 1683
rect 10588 1717 10944 1723
rect 11002 1723 11012 1735
rect 12002 1723 12012 1735
rect 11002 1717 12012 1723
rect 12070 1723 12080 1735
rect 13666 1726 13712 1772
rect 13744 1734 13820 1740
rect 13744 1726 13756 1734
rect 12070 1717 12426 1723
rect 10588 1683 10600 1717
rect 10634 1683 10944 1717
rect 11002 1683 11312 1717
rect 11346 1683 11668 1717
rect 11702 1683 12012 1717
rect 12070 1683 12380 1717
rect 12414 1683 12426 1717
rect 10588 1677 10944 1683
rect 11002 1677 12012 1683
rect 12070 1677 12426 1683
rect 13666 1700 13756 1726
rect 13808 1726 13820 1734
rect 13848 1726 13894 1784
rect 13962 2040 14008 2052
rect 13962 1784 13968 2040
rect 14002 1784 14008 2040
rect 13962 1772 14008 1784
rect 14140 2040 14186 2052
rect 14140 1784 14146 2040
rect 14180 1784 14186 2040
rect 14140 1772 14186 1784
rect 14254 2040 14300 2052
rect 14254 1784 14260 2040
rect 14294 1784 14300 2040
rect 14254 1772 14300 1784
rect 14432 2040 14478 2052
rect 14432 1784 14438 2040
rect 14472 1784 14478 2040
rect 14432 1772 14478 1784
rect 14546 2040 14592 2052
rect 14546 1784 14552 2040
rect 14586 1784 14592 2040
rect 14546 1772 14592 1784
rect 14724 2040 14770 2052
rect 14724 1784 14730 2040
rect 14764 1784 14770 2040
rect 14724 1772 14770 1784
rect 14838 2040 14884 2052
rect 14838 1784 14844 2040
rect 14878 1784 14884 2040
rect 14838 1772 14884 1784
rect 15016 2040 15062 2052
rect 15016 1784 15022 2040
rect 15056 1784 15062 2040
rect 15016 1772 15062 1784
rect 15130 2040 15176 2052
rect 15130 1784 15136 2040
rect 15170 1784 15176 2040
rect 15130 1772 15176 1784
rect 15308 2040 15354 2052
rect 15308 1784 15314 2040
rect 15348 1784 15354 2040
rect 15308 1772 15354 1784
rect 15422 2040 15468 2084
rect 15422 1784 15428 2040
rect 15462 1784 15468 2040
rect 13808 1700 13894 1726
rect 13666 1680 13894 1700
rect 14036 1734 14112 1740
rect 14036 1700 14048 1734
rect 14100 1700 14112 1734
rect 14036 1694 14112 1700
rect 674 1633 750 1639
rect 674 1599 686 1633
rect 738 1599 750 1633
rect 674 1523 750 1599
rect 852 1633 928 1639
rect 852 1599 864 1633
rect 916 1599 928 1633
rect 852 1593 928 1599
rect 1030 1633 1106 1639
rect 1030 1599 1042 1633
rect 1094 1599 1106 1633
rect 1030 1593 1106 1599
rect 1208 1633 1284 1639
rect 1208 1599 1220 1633
rect 1272 1599 1284 1633
rect 1208 1593 1284 1599
rect 1386 1633 1462 1639
rect 1386 1599 1398 1633
rect 1450 1599 1462 1633
rect 1386 1593 1462 1599
rect 1564 1633 1640 1639
rect 1564 1599 1576 1633
rect 1628 1599 1640 1633
rect 1564 1593 1640 1599
rect 1742 1633 1818 1639
rect 1742 1599 1754 1633
rect 1806 1599 1818 1633
rect 1742 1593 1818 1599
rect 1920 1633 1996 1639
rect 1920 1599 1932 1633
rect 1984 1599 1996 1633
rect 1920 1593 1996 1599
rect 2098 1633 2174 1639
rect 2098 1599 2110 1633
rect 2162 1599 2174 1633
rect 2098 1593 2174 1599
rect 2276 1633 2352 1639
rect 2276 1599 2288 1633
rect 2340 1599 2352 1633
rect 2276 1593 2352 1599
rect 2454 1633 2530 1639
rect 2454 1599 2466 1633
rect 2518 1599 2530 1633
rect 2454 1593 2530 1599
rect 2632 1633 2708 1639
rect 2632 1599 2644 1633
rect 2696 1599 2708 1633
rect 2632 1593 2708 1599
rect 2810 1633 2886 1639
rect 2810 1599 2822 1633
rect 2874 1599 2886 1633
rect 2810 1593 2886 1599
rect 2988 1633 3064 1639
rect 2988 1599 3000 1633
rect 3052 1599 3064 1633
rect 2988 1593 3064 1599
rect 3166 1633 3242 1639
rect 3166 1599 3178 1633
rect 3230 1599 3242 1633
rect 3166 1593 3242 1599
rect 3344 1633 3420 1639
rect 3344 1599 3356 1633
rect 3408 1599 3420 1633
rect 852 1523 928 1529
rect 1030 1523 1106 1529
rect 1208 1523 1284 1529
rect 1386 1523 1462 1529
rect 1564 1523 1640 1529
rect 1742 1523 1818 1529
rect 1920 1523 1996 1529
rect 2098 1523 2174 1529
rect 2276 1523 2352 1529
rect 2454 1523 2530 1529
rect 2632 1523 2708 1529
rect 2810 1523 2886 1529
rect 2988 1523 3064 1529
rect 3166 1523 3242 1529
rect 3344 1523 3420 1599
rect 674 1489 686 1523
rect 738 1489 864 1523
rect 916 1489 1042 1523
rect 1094 1489 1220 1523
rect 1272 1489 1398 1523
rect 1450 1489 1576 1523
rect 1628 1489 1754 1523
rect 1806 1489 1932 1523
rect 1984 1489 2110 1523
rect 2162 1489 2288 1523
rect 2340 1489 2466 1523
rect 2518 1489 2644 1523
rect 2696 1489 2822 1523
rect 2874 1489 3000 1523
rect 3052 1489 3178 1523
rect 3230 1489 3356 1523
rect 3408 1489 3420 1523
rect 674 1483 750 1489
rect 852 1483 928 1489
rect 1030 1483 1106 1489
rect 1208 1483 1284 1489
rect 1386 1483 1462 1489
rect 1564 1483 1640 1489
rect 1742 1483 1818 1489
rect 1920 1483 1996 1489
rect 2098 1483 2174 1489
rect 2276 1483 2352 1489
rect 2454 1483 2530 1489
rect 2632 1483 2708 1489
rect 2810 1483 2886 1489
rect 2988 1483 3064 1489
rect 3166 1483 3242 1489
rect 3344 1483 3420 1489
rect 4074 1633 4150 1639
rect 4074 1599 4086 1633
rect 4138 1599 4150 1633
rect 4074 1523 4150 1599
rect 4252 1633 4328 1639
rect 4252 1599 4264 1633
rect 4316 1599 4328 1633
rect 4252 1593 4328 1599
rect 4430 1633 4506 1639
rect 4430 1599 4442 1633
rect 4494 1599 4506 1633
rect 4430 1593 4506 1599
rect 4608 1633 4684 1639
rect 4608 1599 4620 1633
rect 4672 1599 4684 1633
rect 4608 1593 4684 1599
rect 4786 1633 4862 1639
rect 4786 1599 4798 1633
rect 4850 1599 4862 1633
rect 4786 1593 4862 1599
rect 4964 1633 5040 1639
rect 4964 1599 4976 1633
rect 5028 1599 5040 1633
rect 4964 1593 5040 1599
rect 5142 1633 5218 1639
rect 5142 1599 5154 1633
rect 5206 1599 5218 1633
rect 5142 1593 5218 1599
rect 5320 1633 5396 1639
rect 5320 1599 5332 1633
rect 5384 1599 5396 1633
rect 5320 1593 5396 1599
rect 5498 1633 5574 1639
rect 5498 1599 5510 1633
rect 5562 1599 5574 1633
rect 5498 1593 5574 1599
rect 5676 1633 5752 1639
rect 5676 1599 5688 1633
rect 5740 1599 5752 1633
rect 5676 1593 5752 1599
rect 5854 1633 5930 1639
rect 5854 1599 5866 1633
rect 5918 1599 5930 1633
rect 5854 1593 5930 1599
rect 6032 1633 6108 1639
rect 6032 1599 6044 1633
rect 6096 1599 6108 1633
rect 6032 1593 6108 1599
rect 6210 1633 6286 1639
rect 6210 1599 6222 1633
rect 6274 1599 6286 1633
rect 6210 1593 6286 1599
rect 6388 1633 6464 1639
rect 6388 1599 6400 1633
rect 6452 1599 6464 1633
rect 6388 1593 6464 1599
rect 6566 1633 6642 1639
rect 6566 1599 6578 1633
rect 6630 1599 6642 1633
rect 6566 1593 6642 1599
rect 6744 1633 6820 1639
rect 6744 1599 6756 1633
rect 6808 1599 6820 1633
rect 4252 1523 4328 1529
rect 4430 1523 4506 1529
rect 4608 1523 4684 1529
rect 4786 1523 4862 1529
rect 4964 1523 5040 1529
rect 5142 1523 5218 1529
rect 5320 1523 5396 1529
rect 5498 1523 5574 1529
rect 5676 1523 5752 1529
rect 5854 1523 5930 1529
rect 6032 1523 6108 1529
rect 6210 1523 6286 1529
rect 6388 1523 6464 1529
rect 6566 1523 6642 1529
rect 6744 1523 6820 1599
rect 4074 1489 4086 1523
rect 4138 1489 4264 1523
rect 4316 1489 4442 1523
rect 4494 1489 4620 1523
rect 4672 1489 4798 1523
rect 4850 1489 4976 1523
rect 5028 1489 5154 1523
rect 5206 1489 5332 1523
rect 5384 1489 5510 1523
rect 5562 1489 5688 1523
rect 5740 1489 5866 1523
rect 5918 1489 6044 1523
rect 6096 1489 6222 1523
rect 6274 1489 6400 1523
rect 6452 1489 6578 1523
rect 6630 1489 6756 1523
rect 6808 1489 6820 1523
rect 4074 1483 4150 1489
rect 4252 1483 4328 1489
rect 4430 1483 4506 1489
rect 4608 1483 4684 1489
rect 4786 1483 4862 1489
rect 4964 1483 5040 1489
rect 5142 1483 5218 1489
rect 5320 1483 5396 1489
rect 5498 1483 5574 1489
rect 5676 1483 5752 1489
rect 5854 1483 5930 1489
rect 6032 1483 6108 1489
rect 6210 1483 6286 1489
rect 6388 1483 6464 1489
rect 6566 1483 6642 1489
rect 6744 1483 6820 1489
rect 7803 1633 7879 1639
rect 7803 1599 7815 1633
rect 7867 1599 7879 1633
rect 7803 1523 7879 1599
rect 7981 1633 8057 1639
rect 7981 1599 7993 1633
rect 8045 1599 8057 1633
rect 7981 1593 8057 1599
rect 8159 1633 8235 1639
rect 8159 1599 8171 1633
rect 8223 1599 8235 1633
rect 8159 1593 8235 1599
rect 8337 1633 8413 1639
rect 8337 1599 8349 1633
rect 8401 1599 8413 1633
rect 8337 1593 8413 1599
rect 8515 1633 8591 1639
rect 8515 1599 8527 1633
rect 8579 1599 8591 1633
rect 8515 1593 8591 1599
rect 8693 1633 8769 1639
rect 8693 1599 8705 1633
rect 8757 1599 8769 1633
rect 8693 1593 8769 1599
rect 8871 1633 8947 1639
rect 8871 1599 8883 1633
rect 8935 1599 8947 1633
rect 8871 1593 8947 1599
rect 9049 1633 9125 1639
rect 9049 1599 9061 1633
rect 9113 1599 9125 1633
rect 9049 1593 9125 1599
rect 9227 1633 9303 1639
rect 9227 1599 9239 1633
rect 9291 1599 9303 1633
rect 9227 1593 9303 1599
rect 9405 1633 9481 1639
rect 9405 1599 9417 1633
rect 9469 1599 9481 1633
rect 9405 1593 9481 1599
rect 9583 1633 9659 1639
rect 9583 1599 9595 1633
rect 9647 1599 9659 1633
rect 9583 1593 9659 1599
rect 9761 1633 9837 1639
rect 9761 1599 9773 1633
rect 9825 1599 9837 1633
rect 7981 1523 8057 1529
rect 8159 1523 8235 1529
rect 8337 1523 8413 1529
rect 8515 1523 8591 1529
rect 8693 1523 8769 1529
rect 8871 1523 8947 1529
rect 9049 1523 9125 1529
rect 9227 1523 9303 1529
rect 9405 1523 9481 1529
rect 9583 1523 9659 1529
rect 9761 1523 9837 1599
rect 7803 1489 7815 1523
rect 7867 1489 7993 1523
rect 8045 1489 8171 1523
rect 8223 1489 8349 1523
rect 8401 1489 8527 1523
rect 8579 1489 8705 1523
rect 8757 1489 8883 1523
rect 8935 1489 9061 1523
rect 9113 1489 9239 1523
rect 9291 1489 9417 1523
rect 9469 1489 9595 1523
rect 9647 1489 9773 1523
rect 9825 1489 9837 1523
rect 7803 1483 7879 1489
rect 7981 1483 8057 1489
rect 8159 1483 8235 1489
rect 8337 1483 8413 1489
rect 8515 1483 8591 1489
rect 8693 1483 8769 1489
rect 8871 1483 8947 1489
rect 9049 1483 9125 1489
rect 9227 1483 9303 1489
rect 9405 1483 9481 1489
rect 9583 1483 9659 1489
rect 9761 1483 9837 1489
rect 10490 1633 10566 1639
rect 10490 1599 10502 1633
rect 10554 1599 10566 1633
rect 10490 1523 10566 1599
rect 10668 1633 10744 1639
rect 10668 1599 10680 1633
rect 10732 1599 10744 1633
rect 10668 1593 10744 1599
rect 10846 1633 10922 1639
rect 10846 1599 10858 1633
rect 10910 1599 10922 1633
rect 10846 1593 10922 1599
rect 11024 1633 11100 1639
rect 11024 1599 11036 1633
rect 11088 1599 11100 1633
rect 11024 1593 11100 1599
rect 11202 1633 11278 1639
rect 11202 1599 11214 1633
rect 11266 1599 11278 1633
rect 11202 1593 11278 1599
rect 11380 1633 11456 1639
rect 11380 1599 11392 1633
rect 11444 1599 11456 1633
rect 11380 1593 11456 1599
rect 11558 1633 11634 1639
rect 11558 1599 11570 1633
rect 11622 1599 11634 1633
rect 11558 1593 11634 1599
rect 11736 1633 11812 1639
rect 11736 1599 11748 1633
rect 11800 1599 11812 1633
rect 11736 1593 11812 1599
rect 11914 1633 11990 1639
rect 11914 1599 11926 1633
rect 11978 1599 11990 1633
rect 11914 1593 11990 1599
rect 12092 1633 12168 1639
rect 12092 1599 12104 1633
rect 12156 1599 12168 1633
rect 12092 1593 12168 1599
rect 12270 1633 12346 1639
rect 12270 1599 12282 1633
rect 12334 1599 12346 1633
rect 12270 1593 12346 1599
rect 12448 1633 12524 1639
rect 12448 1599 12460 1633
rect 12512 1599 12524 1633
rect 10668 1523 10744 1529
rect 10846 1523 10922 1529
rect 11024 1523 11100 1529
rect 11202 1523 11278 1529
rect 11380 1523 11456 1529
rect 11558 1523 11634 1529
rect 11736 1523 11812 1529
rect 11914 1523 11990 1529
rect 12092 1523 12168 1529
rect 12270 1523 12346 1529
rect 12448 1523 12524 1599
rect 10490 1489 10502 1523
rect 10554 1489 10680 1523
rect 10732 1489 10858 1523
rect 10910 1489 11036 1523
rect 11088 1489 11214 1523
rect 11266 1489 11392 1523
rect 11444 1489 11570 1523
rect 11622 1489 11748 1523
rect 11800 1489 11926 1523
rect 11978 1489 12104 1523
rect 12156 1489 12282 1523
rect 12334 1489 12460 1523
rect 12512 1489 12524 1523
rect 10490 1483 10566 1489
rect 10668 1483 10744 1489
rect 10846 1483 10922 1489
rect 11024 1483 11100 1489
rect 11202 1483 11278 1489
rect 11380 1483 11456 1489
rect 11558 1483 11634 1489
rect 11736 1483 11812 1489
rect 11914 1483 11990 1489
rect 12092 1483 12168 1489
rect 12270 1483 12346 1489
rect 12448 1483 12524 1489
rect 13666 1634 13712 1680
rect 13848 1634 13894 1680
rect 13666 1626 13894 1634
rect 14057 1632 14091 1694
rect 13666 1592 13756 1626
rect 13808 1592 13894 1626
rect 13666 1588 13894 1592
rect 13666 1554 13712 1588
rect 13744 1586 13820 1588
rect 13666 1542 13716 1554
rect 584 1387 594 1445
rect 652 1439 2018 1445
rect 2076 1439 3442 1445
rect 652 1405 962 1439
rect 996 1405 1318 1439
rect 1352 1405 1674 1439
rect 1708 1405 2018 1439
rect 2076 1405 2386 1439
rect 2420 1405 2742 1439
rect 2776 1405 3098 1439
rect 3132 1405 3442 1439
rect 652 1399 2018 1405
rect 652 1387 662 1399
rect 2008 1387 2018 1399
rect 2076 1399 3442 1405
rect 2076 1387 2086 1399
rect 3432 1387 3442 1399
rect 3500 1387 3510 1445
rect 3984 1387 3994 1445
rect 4052 1439 5418 1445
rect 5476 1439 6842 1445
rect 4052 1405 4362 1439
rect 4396 1405 4718 1439
rect 4752 1405 5074 1439
rect 5108 1405 5418 1439
rect 5476 1405 5786 1439
rect 5820 1405 6142 1439
rect 6176 1405 6498 1439
rect 6532 1405 6842 1439
rect 4052 1399 5418 1405
rect 4052 1387 4062 1399
rect 5408 1387 5418 1399
rect 5476 1399 6842 1405
rect 5476 1387 5486 1399
rect 6832 1387 6842 1399
rect 6900 1387 6910 1445
rect 7713 1387 7723 1445
rect 7781 1439 8791 1445
rect 8849 1439 9859 1445
rect 7781 1405 8091 1439
rect 8125 1405 8447 1439
rect 8481 1405 8791 1439
rect 8849 1405 9159 1439
rect 9193 1405 9515 1439
rect 9549 1405 9859 1439
rect 7781 1399 8791 1405
rect 7781 1387 7791 1399
rect 8781 1387 8791 1399
rect 8849 1399 9859 1405
rect 8849 1387 8859 1399
rect 9849 1387 9859 1399
rect 9917 1387 9927 1445
rect 10400 1387 10410 1445
rect 10468 1439 11478 1445
rect 11536 1439 12546 1445
rect 10468 1405 10778 1439
rect 10812 1405 11134 1439
rect 11168 1405 11478 1439
rect 11536 1405 11846 1439
rect 11880 1405 12202 1439
rect 12236 1405 12546 1439
rect 10468 1399 11478 1405
rect 10468 1387 10478 1399
rect 11468 1387 11478 1399
rect 11536 1399 12546 1405
rect 11536 1387 11546 1399
rect 12536 1387 12546 1399
rect 12604 1387 12614 1445
rect 13666 1286 13676 1542
rect 13710 1286 13716 1542
rect 13666 1274 13716 1286
rect 13848 1542 13894 1588
rect 14036 1626 14112 1632
rect 14036 1592 14048 1626
rect 14100 1592 14112 1626
rect 14036 1586 14112 1592
rect 14146 1554 14180 1772
rect 14328 1734 14404 1740
rect 14328 1700 14340 1734
rect 14392 1700 14404 1734
rect 14328 1694 14404 1700
rect 14349 1632 14383 1694
rect 14328 1626 14404 1632
rect 14328 1592 14340 1626
rect 14392 1592 14404 1626
rect 14328 1586 14404 1592
rect 14438 1554 14472 1772
rect 14620 1734 14696 1740
rect 14620 1700 14632 1734
rect 14684 1700 14696 1734
rect 14620 1694 14696 1700
rect 14641 1632 14675 1694
rect 14620 1626 14696 1632
rect 14620 1592 14632 1626
rect 14684 1592 14696 1626
rect 14620 1586 14696 1592
rect 14730 1554 14764 1772
rect 14912 1734 14988 1740
rect 14912 1700 14924 1734
rect 14976 1700 14988 1734
rect 14912 1694 14988 1700
rect 14933 1632 14967 1694
rect 14912 1626 14988 1632
rect 14912 1592 14924 1626
rect 14976 1592 14988 1626
rect 14912 1586 14988 1592
rect 15022 1554 15056 1772
rect 15204 1734 15280 1740
rect 15204 1700 15216 1734
rect 15268 1700 15280 1734
rect 15204 1694 15280 1700
rect 15224 1632 15258 1694
rect 15204 1626 15280 1632
rect 15204 1592 15216 1626
rect 15268 1592 15280 1626
rect 15204 1586 15280 1592
rect 15314 1554 15348 1772
rect 15422 1740 15468 1784
rect 15600 2040 15646 2084
rect 16728 2057 16738 2115
rect 16796 2110 16806 2115
rect 16796 2104 17183 2110
rect 16796 2070 17106 2104
rect 17140 2070 17183 2104
rect 16796 2064 17183 2070
rect 16796 2057 16806 2064
rect 17173 2052 17183 2064
rect 17241 2104 17539 2110
rect 17241 2070 17462 2104
rect 17496 2070 17539 2104
rect 17241 2064 17539 2070
rect 17241 2052 17251 2064
rect 17529 2052 17539 2064
rect 17597 2104 18162 2110
rect 17597 2070 17818 2104
rect 17852 2070 18162 2104
rect 17597 2064 18162 2070
rect 17597 2052 17607 2064
rect 18152 2052 18162 2064
rect 18220 2052 18230 2110
rect 15600 1784 15606 2040
rect 15640 1784 15646 2040
rect 16550 1842 16560 1900
rect 16618 1888 16628 1900
rect 16905 1888 16915 1901
rect 16618 1843 16915 1888
rect 16973 1888 16983 1901
rect 17796 1888 17806 1900
rect 16973 1882 17806 1888
rect 16973 1848 17284 1882
rect 17318 1848 17640 1882
rect 17674 1848 17806 1882
rect 16973 1843 17806 1848
rect 16618 1842 17806 1843
rect 17864 1888 17874 1900
rect 17974 1888 17984 1900
rect 17864 1842 17984 1888
rect 18042 1842 18052 1900
rect 15600 1740 15646 1784
rect 16636 1798 18143 1804
rect 16636 1764 16652 1798
rect 16704 1764 16830 1798
rect 16882 1764 17008 1798
rect 17060 1764 17186 1798
rect 17238 1764 17364 1798
rect 17416 1764 17542 1798
rect 17594 1764 17720 1798
rect 17772 1764 17898 1798
rect 17950 1764 18076 1798
rect 18128 1764 18143 1798
rect 16636 1756 18143 1764
rect 15422 1734 15646 1740
rect 15422 1700 15508 1734
rect 15560 1700 15646 1734
rect 15422 1694 15646 1700
rect 15422 1632 15468 1694
rect 15600 1632 15646 1694
rect 15422 1626 15646 1632
rect 15422 1592 15508 1626
rect 15560 1592 15646 1626
rect 15422 1586 15646 1592
rect 16640 1628 16716 1634
rect 16818 1628 16894 1634
rect 16996 1628 17072 1634
rect 17173 1628 17183 1646
rect 17241 1628 17251 1646
rect 17352 1628 17428 1634
rect 17529 1628 17539 1646
rect 17597 1628 17607 1646
rect 17708 1628 17784 1634
rect 17886 1628 17962 1634
rect 18064 1628 18140 1634
rect 16640 1594 16652 1628
rect 16704 1594 16830 1628
rect 16882 1594 17008 1628
rect 17060 1594 17183 1628
rect 17241 1594 17364 1628
rect 17416 1594 17539 1628
rect 17597 1594 17720 1628
rect 17772 1594 17898 1628
rect 17950 1594 18076 1628
rect 18128 1594 18140 1628
rect 16640 1588 16716 1594
rect 16818 1588 16894 1594
rect 16996 1588 17072 1594
rect 17173 1588 17183 1594
rect 17241 1588 17251 1594
rect 17352 1588 17428 1594
rect 17529 1588 17539 1594
rect 17597 1588 17607 1594
rect 17708 1588 17784 1594
rect 17886 1588 17962 1594
rect 18064 1588 18140 1594
rect 13848 1286 13854 1542
rect 13888 1286 13894 1542
rect 1474 1223 1484 1235
rect 772 1217 1484 1223
rect 1542 1223 1552 1235
rect 2542 1223 2552 1235
rect 1542 1217 2552 1223
rect 2610 1223 2620 1235
rect 4874 1223 4884 1235
rect 2610 1217 3322 1223
rect 772 1183 784 1217
rect 818 1183 1140 1217
rect 1174 1183 1484 1217
rect 1542 1183 1852 1217
rect 1886 1183 2208 1217
rect 2242 1183 2552 1217
rect 2610 1183 2920 1217
rect 2954 1183 3276 1217
rect 3310 1183 3322 1217
rect 772 1177 1484 1183
rect 1542 1177 2552 1183
rect 2610 1177 3322 1183
rect 4172 1217 4884 1223
rect 4942 1223 4952 1235
rect 5942 1223 5952 1235
rect 4942 1217 5952 1223
rect 6010 1223 6020 1235
rect 8247 1223 8257 1235
rect 6010 1217 6722 1223
rect 4172 1183 4184 1217
rect 4218 1183 4540 1217
rect 4574 1183 4884 1217
rect 4942 1183 5252 1217
rect 5286 1183 5608 1217
rect 5642 1183 5952 1217
rect 6010 1183 6320 1217
rect 6354 1183 6676 1217
rect 6710 1183 6722 1217
rect 4172 1177 4884 1183
rect 4942 1177 5952 1183
rect 6010 1177 6722 1183
rect 7901 1217 8257 1223
rect 8315 1223 8325 1235
rect 9315 1223 9325 1235
rect 8315 1217 9325 1223
rect 9383 1223 9393 1235
rect 10934 1223 10944 1235
rect 9383 1217 9739 1223
rect 7901 1183 7913 1217
rect 7947 1183 8257 1217
rect 8315 1183 8625 1217
rect 8659 1183 8981 1217
rect 9015 1183 9325 1217
rect 9383 1183 9693 1217
rect 9727 1183 9739 1217
rect 7901 1177 8257 1183
rect 8315 1177 9325 1183
rect 9383 1177 9739 1183
rect 10588 1217 10944 1223
rect 11002 1223 11012 1235
rect 12002 1223 12012 1235
rect 11002 1217 12012 1223
rect 12070 1223 12080 1235
rect 13666 1224 13712 1274
rect 13744 1236 13820 1242
rect 13744 1224 13756 1236
rect 12070 1217 12426 1223
rect 10588 1183 10600 1217
rect 10634 1183 10944 1217
rect 11002 1183 11312 1217
rect 11346 1183 11668 1217
rect 11702 1183 12012 1217
rect 12070 1183 12380 1217
rect 12414 1183 12426 1217
rect 10588 1177 10944 1183
rect 11002 1177 12012 1183
rect 12070 1177 12426 1183
rect 13666 1202 13756 1224
rect 13808 1224 13820 1236
rect 13848 1224 13894 1286
rect 13962 1542 14008 1554
rect 13962 1286 13968 1542
rect 14002 1286 14008 1542
rect 13962 1274 14008 1286
rect 14140 1542 14186 1554
rect 14140 1286 14146 1542
rect 14180 1286 14186 1542
rect 14140 1274 14186 1286
rect 14254 1542 14300 1554
rect 14254 1286 14260 1542
rect 14294 1286 14300 1542
rect 14254 1274 14300 1286
rect 14432 1542 14478 1554
rect 14432 1286 14438 1542
rect 14472 1286 14478 1542
rect 14432 1274 14478 1286
rect 14546 1542 14592 1554
rect 14546 1286 14552 1542
rect 14586 1286 14592 1542
rect 14546 1274 14592 1286
rect 14724 1542 14770 1554
rect 14724 1286 14730 1542
rect 14764 1286 14770 1542
rect 14724 1274 14770 1286
rect 14838 1542 14884 1554
rect 14838 1286 14844 1542
rect 14878 1286 14884 1542
rect 14838 1274 14884 1286
rect 15016 1542 15062 1554
rect 15016 1286 15022 1542
rect 15056 1286 15062 1542
rect 15016 1274 15062 1286
rect 15130 1542 15176 1554
rect 15130 1286 15136 1542
rect 15170 1286 15176 1542
rect 15130 1274 15176 1286
rect 15308 1542 15354 1554
rect 15308 1286 15314 1542
rect 15348 1286 15354 1542
rect 15308 1274 15354 1286
rect 15422 1542 15468 1586
rect 15422 1286 15428 1542
rect 15462 1286 15468 1542
rect 13808 1202 13894 1224
rect 13666 1178 13894 1202
rect 13666 1142 13712 1178
rect 13848 1142 13894 1178
rect 674 1133 750 1139
rect 674 1099 686 1133
rect 738 1099 750 1133
rect 674 1023 750 1099
rect 852 1133 928 1139
rect 852 1099 864 1133
rect 916 1099 928 1133
rect 852 1093 928 1099
rect 1030 1133 1106 1139
rect 1030 1099 1042 1133
rect 1094 1099 1106 1133
rect 1030 1093 1106 1099
rect 1208 1133 1284 1139
rect 1208 1099 1220 1133
rect 1272 1099 1284 1133
rect 1208 1093 1284 1099
rect 1386 1133 1462 1139
rect 1386 1099 1398 1133
rect 1450 1099 1462 1133
rect 1386 1093 1462 1099
rect 1564 1133 1640 1139
rect 1564 1099 1576 1133
rect 1628 1099 1640 1133
rect 1564 1093 1640 1099
rect 1742 1133 1818 1139
rect 1742 1099 1754 1133
rect 1806 1099 1818 1133
rect 1742 1093 1818 1099
rect 1920 1133 1996 1139
rect 1920 1099 1932 1133
rect 1984 1099 1996 1133
rect 1920 1093 1996 1099
rect 2098 1133 2174 1139
rect 2098 1099 2110 1133
rect 2162 1099 2174 1133
rect 2098 1093 2174 1099
rect 2276 1133 2352 1139
rect 2276 1099 2288 1133
rect 2340 1099 2352 1133
rect 2276 1093 2352 1099
rect 2454 1133 2530 1139
rect 2454 1099 2466 1133
rect 2518 1099 2530 1133
rect 2454 1093 2530 1099
rect 2632 1133 2708 1139
rect 2632 1099 2644 1133
rect 2696 1099 2708 1133
rect 2632 1093 2708 1099
rect 2810 1133 2886 1139
rect 2810 1099 2822 1133
rect 2874 1099 2886 1133
rect 2810 1093 2886 1099
rect 2988 1133 3064 1139
rect 2988 1099 3000 1133
rect 3052 1099 3064 1133
rect 2988 1093 3064 1099
rect 3166 1133 3242 1139
rect 3166 1099 3178 1133
rect 3230 1099 3242 1133
rect 3166 1093 3242 1099
rect 3344 1133 3420 1139
rect 3344 1099 3356 1133
rect 3408 1099 3420 1133
rect 852 1023 928 1029
rect 1030 1023 1106 1029
rect 1208 1023 1284 1029
rect 1386 1023 1462 1029
rect 1564 1023 1640 1029
rect 1742 1023 1818 1029
rect 1920 1023 1996 1029
rect 2098 1023 2174 1029
rect 2276 1023 2352 1029
rect 2454 1023 2530 1029
rect 2632 1023 2708 1029
rect 2810 1023 2886 1029
rect 2988 1023 3064 1029
rect 3166 1023 3242 1029
rect 3344 1023 3420 1099
rect 674 989 686 1023
rect 738 989 864 1023
rect 916 989 1042 1023
rect 1094 989 1220 1023
rect 1272 989 1398 1023
rect 1450 989 1576 1023
rect 1628 989 1754 1023
rect 1806 989 1932 1023
rect 1984 989 2110 1023
rect 2162 989 2288 1023
rect 2340 989 2466 1023
rect 2518 989 2644 1023
rect 2696 989 2822 1023
rect 2874 989 3000 1023
rect 3052 989 3178 1023
rect 3230 989 3356 1023
rect 3408 989 3420 1023
rect 674 983 750 989
rect 852 983 928 989
rect 1030 983 1106 989
rect 1208 983 1284 989
rect 1386 983 1462 989
rect 1564 983 1640 989
rect 1742 983 1818 989
rect 1920 983 1996 989
rect 2098 983 2174 989
rect 2276 983 2352 989
rect 2454 983 2530 989
rect 2632 983 2708 989
rect 2810 983 2886 989
rect 2988 983 3064 989
rect 3166 983 3242 989
rect 3344 983 3420 989
rect 4074 1133 4150 1139
rect 4074 1099 4086 1133
rect 4138 1099 4150 1133
rect 4074 1023 4150 1099
rect 4252 1133 4328 1139
rect 4252 1099 4264 1133
rect 4316 1099 4328 1133
rect 4252 1093 4328 1099
rect 4430 1133 4506 1139
rect 4430 1099 4442 1133
rect 4494 1099 4506 1133
rect 4430 1093 4506 1099
rect 4608 1133 4684 1139
rect 4608 1099 4620 1133
rect 4672 1099 4684 1133
rect 4608 1093 4684 1099
rect 4786 1133 4862 1139
rect 4786 1099 4798 1133
rect 4850 1099 4862 1133
rect 4786 1093 4862 1099
rect 4964 1133 5040 1139
rect 4964 1099 4976 1133
rect 5028 1099 5040 1133
rect 4964 1093 5040 1099
rect 5142 1133 5218 1139
rect 5142 1099 5154 1133
rect 5206 1099 5218 1133
rect 5142 1093 5218 1099
rect 5320 1133 5396 1139
rect 5320 1099 5332 1133
rect 5384 1099 5396 1133
rect 5320 1093 5396 1099
rect 5498 1133 5574 1139
rect 5498 1099 5510 1133
rect 5562 1099 5574 1133
rect 5498 1093 5574 1099
rect 5676 1133 5752 1139
rect 5676 1099 5688 1133
rect 5740 1099 5752 1133
rect 5676 1093 5752 1099
rect 5854 1133 5930 1139
rect 5854 1099 5866 1133
rect 5918 1099 5930 1133
rect 5854 1093 5930 1099
rect 6032 1133 6108 1139
rect 6032 1099 6044 1133
rect 6096 1099 6108 1133
rect 6032 1093 6108 1099
rect 6210 1133 6286 1139
rect 6210 1099 6222 1133
rect 6274 1099 6286 1133
rect 6210 1093 6286 1099
rect 6388 1133 6464 1139
rect 6388 1099 6400 1133
rect 6452 1099 6464 1133
rect 6388 1093 6464 1099
rect 6566 1133 6642 1139
rect 6566 1099 6578 1133
rect 6630 1099 6642 1133
rect 6566 1093 6642 1099
rect 6744 1133 6820 1139
rect 6744 1099 6756 1133
rect 6808 1099 6820 1133
rect 4252 1023 4328 1029
rect 4430 1023 4506 1029
rect 4608 1023 4684 1029
rect 4786 1023 4862 1029
rect 4964 1023 5040 1029
rect 5142 1023 5218 1029
rect 5320 1023 5396 1029
rect 5498 1023 5574 1029
rect 5676 1023 5752 1029
rect 5854 1023 5930 1029
rect 6032 1023 6108 1029
rect 6210 1023 6286 1029
rect 6388 1023 6464 1029
rect 6566 1023 6642 1029
rect 6744 1023 6820 1099
rect 4074 989 4086 1023
rect 4138 989 4264 1023
rect 4316 989 4442 1023
rect 4494 989 4620 1023
rect 4672 989 4798 1023
rect 4850 989 4976 1023
rect 5028 989 5154 1023
rect 5206 989 5332 1023
rect 5384 989 5510 1023
rect 5562 989 5688 1023
rect 5740 989 5866 1023
rect 5918 989 6044 1023
rect 6096 989 6222 1023
rect 6274 989 6400 1023
rect 6452 989 6578 1023
rect 6630 989 6756 1023
rect 6808 989 6820 1023
rect 4074 983 4150 989
rect 4252 983 4328 989
rect 4430 983 4506 989
rect 4608 983 4684 989
rect 4786 983 4862 989
rect 4964 983 5040 989
rect 5142 983 5218 989
rect 5320 983 5396 989
rect 5498 983 5574 989
rect 5676 983 5752 989
rect 5854 983 5930 989
rect 6032 983 6108 989
rect 6210 983 6286 989
rect 6388 983 6464 989
rect 6566 983 6642 989
rect 6744 983 6820 989
rect 7803 1133 7879 1139
rect 7803 1099 7815 1133
rect 7867 1099 7879 1133
rect 7803 1023 7879 1099
rect 7981 1133 8057 1139
rect 7981 1099 7993 1133
rect 8045 1099 8057 1133
rect 7981 1093 8057 1099
rect 8159 1133 8235 1139
rect 8159 1099 8171 1133
rect 8223 1099 8235 1133
rect 8159 1093 8235 1099
rect 8337 1133 8413 1139
rect 8337 1099 8349 1133
rect 8401 1099 8413 1133
rect 8337 1093 8413 1099
rect 8515 1133 8591 1139
rect 8515 1099 8527 1133
rect 8579 1099 8591 1133
rect 8515 1093 8591 1099
rect 8693 1133 8769 1139
rect 8693 1099 8705 1133
rect 8757 1099 8769 1133
rect 8693 1093 8769 1099
rect 8871 1133 8947 1139
rect 8871 1099 8883 1133
rect 8935 1099 8947 1133
rect 8871 1093 8947 1099
rect 9049 1133 9125 1139
rect 9049 1099 9061 1133
rect 9113 1099 9125 1133
rect 9049 1093 9125 1099
rect 9227 1133 9303 1139
rect 9227 1099 9239 1133
rect 9291 1099 9303 1133
rect 9227 1093 9303 1099
rect 9405 1133 9481 1139
rect 9405 1099 9417 1133
rect 9469 1099 9481 1133
rect 9405 1093 9481 1099
rect 9583 1133 9659 1139
rect 9583 1099 9595 1133
rect 9647 1099 9659 1133
rect 9583 1093 9659 1099
rect 9761 1133 9837 1139
rect 9761 1099 9773 1133
rect 9825 1099 9837 1133
rect 7981 1023 8057 1029
rect 8159 1023 8235 1029
rect 8337 1023 8413 1029
rect 8515 1023 8591 1029
rect 8693 1023 8769 1029
rect 8871 1023 8947 1029
rect 9049 1023 9125 1029
rect 9227 1023 9303 1029
rect 9405 1023 9481 1029
rect 9583 1023 9659 1029
rect 9761 1023 9837 1099
rect 7803 989 7815 1023
rect 7867 989 7993 1023
rect 8045 989 8171 1023
rect 8223 989 8349 1023
rect 8401 989 8527 1023
rect 8579 989 8705 1023
rect 8757 989 8883 1023
rect 8935 989 9061 1023
rect 9113 989 9239 1023
rect 9291 989 9417 1023
rect 9469 989 9595 1023
rect 9647 989 9773 1023
rect 9825 989 9837 1023
rect 7803 983 7879 989
rect 7981 983 8057 989
rect 8159 983 8235 989
rect 8337 983 8413 989
rect 8515 983 8591 989
rect 8693 983 8769 989
rect 8871 983 8947 989
rect 9049 983 9125 989
rect 9227 983 9303 989
rect 9405 983 9481 989
rect 9583 983 9659 989
rect 9761 983 9837 989
rect 10490 1133 10566 1139
rect 10490 1099 10502 1133
rect 10554 1099 10566 1133
rect 10490 1023 10566 1099
rect 10668 1133 10744 1139
rect 10668 1099 10680 1133
rect 10732 1099 10744 1133
rect 10668 1093 10744 1099
rect 10846 1133 10922 1139
rect 10846 1099 10858 1133
rect 10910 1099 10922 1133
rect 10846 1093 10922 1099
rect 11024 1133 11100 1139
rect 11024 1099 11036 1133
rect 11088 1099 11100 1133
rect 11024 1093 11100 1099
rect 11202 1133 11278 1139
rect 11202 1099 11214 1133
rect 11266 1099 11278 1133
rect 11202 1093 11278 1099
rect 11380 1133 11456 1139
rect 11380 1099 11392 1133
rect 11444 1099 11456 1133
rect 11380 1093 11456 1099
rect 11558 1133 11634 1139
rect 11558 1099 11570 1133
rect 11622 1099 11634 1133
rect 11558 1093 11634 1099
rect 11736 1133 11812 1139
rect 11736 1099 11748 1133
rect 11800 1099 11812 1133
rect 11736 1093 11812 1099
rect 11914 1133 11990 1139
rect 11914 1099 11926 1133
rect 11978 1099 11990 1133
rect 11914 1093 11990 1099
rect 12092 1133 12168 1139
rect 12092 1099 12104 1133
rect 12156 1099 12168 1133
rect 12092 1093 12168 1099
rect 12270 1133 12346 1139
rect 12270 1099 12282 1133
rect 12334 1099 12346 1133
rect 12270 1093 12346 1099
rect 12448 1133 12524 1139
rect 12448 1099 12460 1133
rect 12512 1099 12524 1133
rect 10668 1023 10744 1029
rect 10846 1023 10922 1029
rect 11024 1023 11100 1029
rect 11202 1023 11278 1029
rect 11380 1023 11456 1029
rect 11558 1023 11634 1029
rect 11736 1023 11812 1029
rect 11914 1023 11990 1029
rect 12092 1023 12168 1029
rect 12270 1023 12346 1029
rect 12448 1023 12524 1099
rect 10490 989 10502 1023
rect 10554 989 10680 1023
rect 10732 989 10858 1023
rect 10910 989 11036 1023
rect 11088 989 11214 1023
rect 11266 989 11392 1023
rect 11444 989 11570 1023
rect 11622 989 11748 1023
rect 11800 989 11926 1023
rect 11978 989 12104 1023
rect 12156 989 12282 1023
rect 12334 989 12460 1023
rect 12512 989 12524 1023
rect 10490 983 10566 989
rect 10668 983 10744 989
rect 10846 983 10922 989
rect 11024 983 11100 989
rect 11202 983 11278 989
rect 11380 983 11456 989
rect 11558 983 11634 989
rect 11736 983 11812 989
rect 11914 983 11990 989
rect 12092 983 12168 989
rect 12270 983 12346 989
rect 12448 983 12524 989
rect 13666 1128 13894 1142
rect 13666 1096 13756 1128
rect 13666 1056 13712 1096
rect 13744 1094 13756 1096
rect 13808 1096 13894 1128
rect 13808 1094 13820 1096
rect 13744 1088 13820 1094
rect 13666 1044 13716 1056
rect 584 887 594 945
rect 652 939 2018 945
rect 2076 939 3442 945
rect 652 905 962 939
rect 996 905 1318 939
rect 1352 905 1674 939
rect 1708 905 2018 939
rect 2076 905 2386 939
rect 2420 905 2742 939
rect 2776 905 3098 939
rect 3132 905 3442 939
rect 652 899 2018 905
rect 652 887 662 899
rect 2008 887 2018 899
rect 2076 899 3442 905
rect 2076 887 2086 899
rect 3432 887 3442 899
rect 3500 899 3994 945
rect 4052 939 5418 945
rect 5476 939 6842 945
rect 4052 905 4362 939
rect 4396 905 4718 939
rect 4752 905 5074 939
rect 5108 905 5418 939
rect 5476 905 5786 939
rect 5820 905 6142 939
rect 6176 905 6498 939
rect 6532 905 6842 939
rect 3500 887 3510 899
rect 3984 887 3994 899
rect 4052 899 5418 905
rect 4052 887 4062 899
rect 5408 887 5418 899
rect 5476 899 6842 905
rect 5476 887 5486 899
rect 6832 887 6842 899
rect 6900 887 6910 945
rect 7713 887 7723 945
rect 7781 939 8791 945
rect 8849 939 9859 945
rect 7781 905 8091 939
rect 8125 905 8447 939
rect 8481 905 8791 939
rect 8849 905 9159 939
rect 9193 905 9515 939
rect 9549 905 9859 939
rect 7781 899 8791 905
rect 7781 887 7791 899
rect 8781 887 8791 899
rect 8849 899 9859 905
rect 8849 887 8859 899
rect 9849 887 9859 899
rect 9917 887 9927 945
rect 10400 887 10410 945
rect 10468 939 11478 945
rect 11536 939 12546 945
rect 10468 905 10778 939
rect 10812 905 11134 939
rect 11168 905 11478 939
rect 11536 905 11846 939
rect 11880 905 12202 939
rect 12236 905 12546 939
rect 10468 899 11478 905
rect 10468 887 10478 899
rect 11468 887 11478 899
rect 11536 899 12546 905
rect 11536 887 11546 899
rect 12536 887 12546 899
rect 12604 887 12614 945
rect 13666 788 13676 1044
rect 13710 788 13716 1044
rect 13666 776 13716 788
rect 13848 1044 13894 1096
rect 13968 1056 14002 1274
rect 14036 1236 14112 1242
rect 14036 1202 14048 1236
rect 14100 1202 14112 1236
rect 14036 1196 14112 1202
rect 14056 1134 14090 1196
rect 14036 1128 14112 1134
rect 14036 1094 14048 1128
rect 14100 1094 14112 1128
rect 14036 1088 14112 1094
rect 14260 1056 14294 1274
rect 14328 1236 14404 1242
rect 14328 1202 14340 1236
rect 14392 1202 14404 1236
rect 14328 1196 14404 1202
rect 14348 1134 14382 1196
rect 14328 1128 14404 1134
rect 14328 1094 14340 1128
rect 14392 1094 14404 1128
rect 14328 1088 14404 1094
rect 14552 1056 14586 1274
rect 14620 1236 14696 1242
rect 14620 1202 14632 1236
rect 14684 1202 14696 1236
rect 14620 1196 14696 1202
rect 14642 1134 14676 1196
rect 14620 1128 14696 1134
rect 14620 1094 14632 1128
rect 14684 1094 14696 1128
rect 14620 1088 14696 1094
rect 14844 1056 14878 1274
rect 14912 1236 14988 1242
rect 14912 1202 14924 1236
rect 14976 1202 14988 1236
rect 14912 1196 14988 1202
rect 14934 1134 14968 1196
rect 14912 1128 14988 1134
rect 14912 1094 14924 1128
rect 14976 1094 14988 1128
rect 14912 1088 14988 1094
rect 15136 1056 15170 1274
rect 15422 1272 15468 1286
rect 15600 1542 15646 1586
rect 15600 1286 15606 1542
rect 15640 1286 15646 1542
rect 16728 1492 16738 1550
rect 16796 1504 16916 1550
rect 16796 1492 16806 1504
rect 16906 1492 16916 1504
rect 16974 1544 17806 1550
rect 16974 1510 17106 1544
rect 17140 1510 17462 1544
rect 17496 1510 17806 1544
rect 16974 1504 17806 1510
rect 16974 1492 16984 1504
rect 17796 1492 17806 1504
rect 17864 1504 18162 1550
rect 17864 1492 17874 1504
rect 18152 1492 18162 1504
rect 18220 1492 18230 1550
rect 15600 1272 15646 1286
rect 16550 1282 16560 1340
rect 16618 1328 16628 1340
rect 17974 1328 17984 1340
rect 16618 1322 17984 1328
rect 16618 1288 16928 1322
rect 16962 1288 17284 1322
rect 17318 1288 17640 1322
rect 17674 1288 17984 1322
rect 16618 1282 17984 1288
rect 18042 1282 18052 1340
rect 15204 1236 15280 1242
rect 15204 1202 15216 1236
rect 15268 1202 15280 1236
rect 15204 1196 15280 1202
rect 15422 1236 15646 1272
rect 15422 1202 15508 1236
rect 15560 1202 15646 1236
rect 15224 1134 15258 1196
rect 15422 1190 15646 1202
rect 15422 1136 15468 1190
rect 15600 1136 15646 1190
rect 15204 1128 15280 1134
rect 15204 1094 15216 1128
rect 15268 1094 15280 1128
rect 15204 1088 15280 1094
rect 15422 1128 15646 1136
rect 15422 1094 15508 1128
rect 15560 1094 15646 1128
rect 15422 1062 15646 1094
rect 16640 1238 16716 1244
rect 16818 1238 16894 1244
rect 16996 1238 17072 1244
rect 17174 1238 17250 1244
rect 17352 1238 17428 1244
rect 17530 1238 17606 1244
rect 17708 1238 17784 1244
rect 17886 1238 17962 1244
rect 18064 1238 18140 1244
rect 16640 1204 16652 1238
rect 16704 1204 16830 1238
rect 16882 1204 17008 1238
rect 17060 1204 17186 1238
rect 17238 1204 17364 1238
rect 17416 1204 17542 1238
rect 17594 1204 17720 1238
rect 17772 1204 17898 1238
rect 17950 1204 18076 1238
rect 18128 1204 18140 1238
rect 16640 1128 16716 1204
rect 16818 1198 16894 1204
rect 16996 1198 17072 1204
rect 17174 1198 17250 1204
rect 17352 1198 17428 1204
rect 17530 1198 17606 1204
rect 17708 1198 17784 1204
rect 17886 1198 17962 1204
rect 16818 1128 16894 1134
rect 16996 1128 17072 1134
rect 17174 1128 17250 1134
rect 17352 1128 17428 1134
rect 17530 1128 17606 1134
rect 17708 1128 17784 1134
rect 17886 1128 17962 1134
rect 18064 1128 18140 1204
rect 16640 1094 16652 1128
rect 16704 1094 16830 1128
rect 16882 1094 17008 1128
rect 17060 1094 17186 1128
rect 17238 1094 17364 1128
rect 17416 1094 17542 1128
rect 17594 1094 17720 1128
rect 17772 1094 17898 1128
rect 17950 1094 18076 1128
rect 18128 1094 18140 1128
rect 16640 1088 16716 1094
rect 16818 1088 16894 1094
rect 16996 1088 17072 1094
rect 17174 1088 17250 1094
rect 17352 1088 17428 1094
rect 17530 1088 17606 1094
rect 17708 1088 17784 1094
rect 17886 1088 17962 1094
rect 18064 1088 18140 1094
rect 13848 788 13854 1044
rect 13888 788 13894 1044
rect 13666 744 13712 776
rect 13848 744 13894 788
rect 13962 1044 14008 1056
rect 13962 788 13968 1044
rect 14002 788 14008 1044
rect 14140 1044 14186 1056
rect 14140 846 14146 1044
rect 14180 846 14186 1044
rect 14254 1044 14300 1056
rect 14124 788 14134 846
rect 14192 788 14202 846
rect 14254 788 14260 1044
rect 14294 788 14300 1044
rect 14432 1044 14478 1056
rect 14432 846 14438 1044
rect 14472 846 14478 1044
rect 14546 1044 14592 1056
rect 14416 788 14426 846
rect 14484 788 14494 846
rect 14546 788 14552 1044
rect 14586 788 14592 1044
rect 14724 1044 14770 1056
rect 14724 846 14730 1044
rect 14764 846 14770 1044
rect 14838 1044 14884 1056
rect 14708 788 14718 846
rect 14776 788 14786 846
rect 14838 788 14844 1044
rect 14878 788 14884 1044
rect 15016 1044 15062 1056
rect 15016 846 15022 1044
rect 15056 846 15062 1044
rect 15130 1044 15176 1056
rect 15000 788 15010 846
rect 15068 788 15078 846
rect 15130 788 15136 1044
rect 15170 788 15176 1044
rect 15308 1044 15354 1056
rect 15308 846 15314 1044
rect 15348 846 15354 1044
rect 15422 1044 15468 1062
rect 15292 788 15302 846
rect 15360 788 15370 846
rect 15422 788 15428 1044
rect 15462 788 15468 1044
rect 13962 776 14008 788
rect 14140 776 14186 788
rect 14254 776 14300 788
rect 14432 776 14478 788
rect 14546 776 14592 788
rect 14724 776 14770 788
rect 14838 776 14884 788
rect 15016 776 15062 788
rect 15130 776 15176 788
rect 15308 776 15354 788
rect 15422 748 15468 788
rect 15600 1044 15646 1062
rect 15600 788 15606 1044
rect 15640 788 15646 1044
rect 16728 992 16738 1050
rect 16796 1044 18162 1050
rect 16796 1010 17106 1044
rect 17140 1010 17462 1044
rect 17496 1010 17818 1044
rect 17852 1010 18162 1044
rect 16796 1004 18162 1010
rect 16796 992 16806 1004
rect 18152 992 18162 1004
rect 18220 992 18230 1050
rect 15600 748 15646 788
rect 16550 782 16560 840
rect 16618 828 16628 840
rect 17974 828 17984 840
rect 16618 822 17984 828
rect 16618 788 16928 822
rect 16962 788 17284 822
rect 17318 788 17640 822
rect 17674 788 17984 822
rect 16618 782 17984 788
rect 18042 782 18052 840
rect 13666 738 13894 744
rect 1474 723 1484 735
rect 772 717 1484 723
rect 1542 723 1552 735
rect 2542 723 2552 735
rect 1542 717 2552 723
rect 2610 723 2620 735
rect 4874 723 4884 735
rect 2610 717 3322 723
rect 772 683 784 717
rect 818 683 1140 717
rect 1174 683 1484 717
rect 1542 683 1852 717
rect 1886 683 2208 717
rect 2242 683 2552 717
rect 2610 683 2920 717
rect 2954 683 3276 717
rect 3310 683 3322 717
rect 772 677 1484 683
rect 1542 677 2552 683
rect 2610 677 3322 683
rect 4172 717 4884 723
rect 4942 723 4952 735
rect 5942 723 5952 735
rect 4942 717 5952 723
rect 6010 723 6020 735
rect 8247 723 8257 735
rect 6010 717 6722 723
rect 4172 683 4184 717
rect 4218 683 4540 717
rect 4574 683 4884 717
rect 4942 683 5252 717
rect 5286 683 5608 717
rect 5642 683 5952 717
rect 6010 683 6320 717
rect 6354 683 6676 717
rect 6710 683 6722 717
rect 4172 677 4884 683
rect 4942 677 5952 683
rect 6010 677 6722 683
rect 7901 717 8257 723
rect 8315 723 8325 735
rect 9315 723 9325 735
rect 8315 717 9325 723
rect 9383 723 9393 735
rect 10934 723 10944 735
rect 9383 717 9739 723
rect 7901 683 7913 717
rect 7947 683 8257 717
rect 8315 683 8625 717
rect 8659 683 8981 717
rect 9015 683 9325 717
rect 9383 683 9693 717
rect 9727 683 9739 717
rect 7901 677 8257 683
rect 8315 677 9325 683
rect 9383 677 9739 683
rect 10588 717 10944 723
rect 11002 723 11012 735
rect 12002 723 12012 735
rect 11002 717 12012 723
rect 12070 723 12080 735
rect 12070 717 12426 723
rect 10588 683 10600 717
rect 10634 683 10944 717
rect 11002 683 11312 717
rect 11346 683 11668 717
rect 11702 683 12012 717
rect 12070 683 12380 717
rect 12414 683 12426 717
rect 13666 704 13756 738
rect 13808 704 13894 738
rect 13666 698 13894 704
rect 14036 738 14112 744
rect 14328 738 14404 744
rect 14620 738 14696 744
rect 14912 738 14988 744
rect 15204 738 15280 744
rect 14036 704 14048 738
rect 14100 704 14340 738
rect 14392 704 14632 738
rect 14684 704 14924 738
rect 14976 704 15216 738
rect 15268 704 15280 738
rect 14036 698 14112 704
rect 14328 698 14404 704
rect 14620 698 14696 704
rect 14912 698 14988 704
rect 15204 698 15280 704
rect 15422 738 15646 748
rect 15422 704 15508 738
rect 15560 704 15646 738
rect 15422 702 15646 704
rect 15496 698 15572 702
rect 15600 696 15646 702
rect 16640 738 16716 744
rect 16818 738 16894 744
rect 16996 738 17072 744
rect 17174 738 17250 744
rect 17352 739 17428 744
rect 17351 738 17361 739
rect 17419 738 17429 739
rect 17530 738 17606 744
rect 17708 738 17784 744
rect 17886 738 17962 744
rect 18064 738 18140 744
rect 16640 704 16652 738
rect 16704 704 16830 738
rect 16882 704 17008 738
rect 17060 704 17186 738
rect 17238 704 17361 738
rect 17419 704 17542 738
rect 17594 704 17720 738
rect 17772 704 17898 738
rect 17950 704 18076 738
rect 18128 704 18140 738
rect 16640 698 16716 704
rect 16818 698 16894 704
rect 16996 698 17072 704
rect 17174 698 17250 704
rect 10588 677 10944 683
rect 11002 677 12012 683
rect 12070 677 12426 683
rect 17351 681 17361 704
rect 17419 681 17429 704
rect 17530 698 17606 704
rect 17708 698 17784 704
rect 17886 698 17962 704
rect 18064 698 18140 704
rect 674 633 750 639
rect 674 599 686 633
rect 738 599 750 633
rect 674 593 750 599
rect 852 633 928 639
rect 852 599 864 633
rect 916 599 928 633
rect 852 593 928 599
rect 1030 633 1106 639
rect 1030 599 1042 633
rect 1094 599 1106 633
rect 1030 593 1106 599
rect 1208 633 1284 639
rect 1208 599 1220 633
rect 1272 599 1284 633
rect 1208 593 1284 599
rect 1386 633 1462 639
rect 1386 599 1398 633
rect 1450 599 1462 633
rect 1386 593 1462 599
rect 1564 633 1640 639
rect 1564 599 1576 633
rect 1628 599 1640 633
rect 1564 593 1640 599
rect 1742 633 1818 639
rect 1742 599 1754 633
rect 1806 599 1818 633
rect 1742 593 1818 599
rect 1920 633 1996 639
rect 1920 599 1932 633
rect 1984 599 1996 633
rect 1920 593 1996 599
rect 2098 633 2174 639
rect 2098 599 2110 633
rect 2162 599 2174 633
rect 2098 593 2174 599
rect 2276 633 2352 639
rect 2276 599 2288 633
rect 2340 599 2352 633
rect 2276 593 2352 599
rect 2454 633 2530 639
rect 2454 599 2466 633
rect 2518 599 2530 633
rect 2454 593 2530 599
rect 2632 633 2708 639
rect 2632 599 2644 633
rect 2696 599 2708 633
rect 2632 593 2708 599
rect 2810 633 2886 639
rect 2810 599 2822 633
rect 2874 599 2886 633
rect 2810 593 2886 599
rect 2988 633 3064 639
rect 2988 599 3000 633
rect 3052 599 3064 633
rect 2988 593 3064 599
rect 3166 633 3242 639
rect 3166 599 3178 633
rect 3230 599 3242 633
rect 3166 593 3242 599
rect 3344 633 3420 639
rect 3344 599 3356 633
rect 3408 599 3420 633
rect 3344 593 3420 599
rect 4074 633 4150 639
rect 4252 633 4328 639
rect 4430 633 4506 639
rect 4608 633 4684 639
rect 4786 633 4862 639
rect 4964 633 5040 639
rect 5142 633 5218 639
rect 5320 633 5396 639
rect 5498 633 5574 639
rect 5676 633 5752 639
rect 5854 633 5930 639
rect 6032 633 6108 639
rect 6210 633 6286 639
rect 6388 633 6464 639
rect 6566 633 6642 639
rect 6744 633 6820 639
rect 4074 599 4086 633
rect 4138 599 4264 633
rect 4316 599 4442 633
rect 4494 599 4620 633
rect 4672 599 4798 633
rect 4850 599 4976 633
rect 5028 599 5154 633
rect 5206 599 5332 633
rect 5384 599 5510 633
rect 5562 599 5688 633
rect 5740 599 5866 633
rect 5918 599 6044 633
rect 6096 599 6222 633
rect 6274 599 6400 633
rect 6452 599 6578 633
rect 6630 599 6756 633
rect 6808 599 6820 633
rect 4074 593 4150 599
rect 4252 593 4328 599
rect 4430 593 4506 599
rect 4608 593 4684 599
rect 4786 593 4862 599
rect 4964 593 5040 599
rect 5142 593 5218 599
rect 5320 410 5396 599
rect 5498 593 5574 599
rect 5676 593 5752 599
rect 5854 593 5930 599
rect 6032 593 6108 599
rect 6210 593 6286 599
rect 6388 593 6464 599
rect 6566 593 6642 599
rect 6744 593 6820 599
rect 7803 633 7879 639
rect 7981 633 8057 639
rect 8159 633 8235 639
rect 8337 633 8413 639
rect 8515 633 8591 639
rect 8693 633 8769 639
rect 8871 633 8947 639
rect 9049 633 9125 639
rect 9227 633 9303 639
rect 9405 633 9481 639
rect 9583 633 9659 639
rect 9761 633 9837 639
rect 7803 599 7815 633
rect 7867 599 7993 633
rect 8045 599 8171 633
rect 8223 599 8349 633
rect 8401 599 8527 633
rect 8579 599 8705 633
rect 8757 599 8883 633
rect 8935 599 9061 633
rect 9113 599 9239 633
rect 9291 599 9417 633
rect 9469 599 9595 633
rect 9647 599 9773 633
rect 9825 609 9837 633
rect 10490 633 10566 639
rect 10668 633 10744 639
rect 10846 633 10922 639
rect 11024 633 11100 639
rect 11202 633 11278 639
rect 11380 633 11456 639
rect 11558 633 11634 639
rect 11736 633 11812 639
rect 11914 633 11990 639
rect 12092 633 12168 639
rect 12270 633 12346 639
rect 12448 633 12524 639
rect 9825 599 9838 609
rect 7803 593 7879 599
rect 7981 593 8057 599
rect 8159 593 8235 599
rect 8337 593 8413 599
rect 8515 593 8591 599
rect 8693 593 8769 599
rect 8871 593 8947 599
rect 9049 593 9125 599
rect 9227 593 9303 599
rect 9405 593 9481 599
rect 9583 593 9659 599
rect 9761 593 9838 599
rect 9762 410 9838 593
rect 10490 599 10502 633
rect 10554 599 10680 633
rect 10732 599 10858 633
rect 10910 599 11036 633
rect 11088 599 11214 633
rect 11266 599 11392 633
rect 11444 599 11570 633
rect 11622 599 11748 633
rect 11800 599 11926 633
rect 11978 599 12104 633
rect 12156 599 12282 633
rect 12334 599 12460 633
rect 12512 599 12524 633
rect 10490 410 10566 599
rect 10668 593 10744 599
rect 10846 593 10922 599
rect 11024 593 11100 599
rect 11202 593 11278 599
rect 11380 593 11456 599
rect 11558 593 11634 599
rect 11736 593 11812 599
rect 11914 593 11990 599
rect 12092 593 12168 599
rect 12270 593 12346 599
rect 12448 593 12524 599
rect 14097 613 14224 619
rect 14097 516 14109 613
rect 14212 516 14224 613
rect 14097 510 14224 516
rect 15267 614 15394 620
rect 15267 517 15279 614
rect 15382 517 15394 614
rect 16535 611 16652 617
rect 16535 524 16547 611
rect 16640 524 16652 611
rect 16535 518 16652 524
rect 17957 600 18074 606
rect 15267 511 15394 517
rect 17957 513 17969 600
rect 18062 513 18074 600
rect 17957 507 18074 513
rect 5320 380 17429 410
rect 5320 322 17361 380
rect 17419 322 17429 380
rect 5320 293 17429 322
rect 18888 149 19016 3052
rect 19613 2614 19689 2620
rect 19791 2614 19867 2620
rect 19969 2614 20045 2620
rect 20147 2614 20223 2620
rect 20325 2614 20401 2620
rect 20503 2614 20579 2620
rect 20681 2614 20757 2620
rect 20859 2614 20935 2620
rect 21037 2614 21113 2620
rect 19611 2580 19625 2614
rect 19677 2580 19803 2614
rect 19855 2580 19981 2614
rect 20033 2580 20159 2614
rect 20211 2580 20337 2614
rect 20389 2580 20515 2614
rect 20567 2580 20693 2614
rect 20745 2580 20871 2614
rect 20923 2580 21049 2614
rect 21101 2580 21488 2614
rect 19613 2574 19689 2580
rect 19791 2574 19867 2580
rect 19969 2574 20045 2580
rect 20147 2574 20223 2580
rect 20325 2574 20401 2580
rect 20503 2574 20579 2580
rect 20681 2574 20757 2580
rect 20859 2574 20935 2580
rect 21037 2574 21113 2580
rect 20056 2536 20066 2537
rect 19701 2478 19711 2536
rect 19769 2490 20066 2536
rect 20124 2536 20134 2537
rect 20769 2536 20779 2539
rect 19769 2478 19779 2490
rect 20056 2479 20066 2490
rect 20124 2490 20423 2536
rect 20124 2479 20134 2490
rect 20413 2478 20423 2490
rect 20481 2490 20779 2536
rect 20837 2536 20847 2539
rect 20481 2478 20491 2490
rect 20769 2481 20779 2490
rect 20837 2490 21135 2536
rect 20837 2481 20847 2490
rect 21125 2478 21135 2490
rect 21193 2478 21203 2536
rect 19523 2268 19533 2326
rect 19591 2314 19601 2326
rect 20235 2314 20245 2321
rect 19591 2308 20245 2314
rect 20303 2314 20313 2321
rect 20947 2314 20957 2326
rect 20303 2308 20957 2314
rect 19591 2274 19901 2308
rect 19935 2274 20245 2308
rect 20303 2274 20613 2308
rect 20647 2274 20957 2308
rect 19591 2268 20245 2274
rect 20235 2263 20245 2268
rect 20303 2268 20957 2274
rect 21015 2268 21025 2326
rect 20303 2263 20313 2268
rect 19613 2224 19689 2230
rect 19791 2224 19867 2230
rect 19969 2224 20045 2230
rect 20147 2224 20223 2230
rect 20325 2224 20401 2230
rect 20503 2224 20579 2230
rect 20681 2224 20757 2230
rect 20859 2224 20935 2230
rect 21037 2224 21113 2230
rect 19613 2218 19625 2224
rect 19603 2190 19625 2218
rect 19677 2190 19803 2224
rect 19855 2190 19981 2224
rect 20033 2190 20159 2224
rect 20211 2190 20337 2224
rect 20389 2190 20515 2224
rect 20567 2190 20693 2224
rect 20745 2190 20871 2224
rect 20923 2190 21049 2224
rect 21101 2218 21113 2224
rect 21360 2218 21488 2580
rect 21101 2190 21488 2218
rect 19603 2116 21488 2190
rect 19603 2090 19625 2116
rect 19613 2082 19625 2090
rect 19677 2082 19803 2116
rect 19855 2082 19981 2116
rect 20033 2082 20159 2116
rect 20211 2082 20337 2116
rect 20389 2082 20515 2116
rect 20567 2082 20693 2116
rect 20745 2082 20871 2116
rect 20923 2082 21049 2116
rect 21101 2090 21488 2116
rect 21101 2082 21113 2090
rect 19613 2076 19689 2082
rect 19791 2076 19867 2082
rect 19969 2076 20045 2082
rect 20147 2076 20223 2082
rect 20325 2076 20401 2082
rect 20503 2076 20579 2082
rect 20681 2076 20757 2082
rect 20859 2076 20935 2082
rect 21037 2076 21113 2082
rect 20056 2038 20066 2040
rect 19701 1980 19711 2038
rect 19769 1992 20066 2038
rect 20124 2038 20134 2040
rect 20414 2038 20424 2041
rect 19769 1980 19779 1992
rect 20056 1982 20066 1992
rect 20124 1992 20424 2038
rect 20482 2038 20492 2041
rect 20124 1982 20134 1992
rect 20414 1983 20424 1992
rect 20482 1992 20779 2038
rect 20482 1983 20492 1992
rect 20769 1980 20779 1992
rect 20837 1992 21135 2038
rect 20837 1980 20847 1992
rect 21125 1980 21135 1992
rect 21193 1980 21203 2038
rect 19523 1769 19533 1827
rect 19591 1816 19601 1827
rect 20235 1816 20245 1827
rect 19591 1810 20245 1816
rect 20303 1816 20313 1827
rect 20947 1816 20957 1829
rect 20303 1810 20957 1816
rect 19591 1776 19901 1810
rect 19935 1776 20245 1810
rect 20303 1776 20613 1810
rect 20647 1776 20957 1810
rect 19591 1770 20245 1776
rect 19591 1769 19601 1770
rect 20235 1769 20245 1770
rect 20303 1771 20957 1776
rect 21015 1771 21025 1829
rect 20303 1770 21015 1771
rect 20303 1769 20313 1770
rect 19613 1726 19689 1732
rect 19791 1726 19867 1732
rect 19969 1726 20045 1732
rect 20147 1726 20223 1732
rect 20325 1726 20401 1732
rect 20503 1726 20579 1732
rect 20681 1726 20757 1732
rect 20859 1726 20935 1732
rect 21037 1726 21113 1732
rect 19613 1720 19625 1726
rect 19603 1692 19625 1720
rect 19677 1692 19803 1726
rect 19855 1692 19981 1726
rect 20033 1692 20159 1726
rect 20211 1692 20337 1726
rect 20389 1692 20515 1726
rect 20567 1692 20693 1726
rect 20745 1692 20871 1726
rect 20923 1692 21049 1726
rect 21101 1720 21113 1726
rect 21360 1720 21488 2090
rect 21101 1692 21488 1720
rect 19603 1618 21488 1692
rect 19603 1592 19625 1618
rect 19613 1584 19625 1592
rect 19677 1584 19803 1618
rect 19855 1584 19981 1618
rect 20033 1584 20159 1618
rect 20211 1584 20337 1618
rect 20389 1584 20515 1618
rect 20567 1584 20693 1618
rect 20745 1584 20871 1618
rect 20923 1584 21049 1618
rect 21101 1592 21488 1618
rect 21101 1584 21181 1592
rect 19613 1578 19689 1584
rect 19723 1510 19757 1584
rect 19791 1578 19867 1584
rect 19969 1578 20045 1584
rect 20079 1510 20113 1584
rect 20147 1578 20223 1584
rect 20325 1578 20401 1584
rect 20435 1518 20469 1584
rect 20503 1578 20579 1584
rect 20681 1578 20757 1584
rect 20413 1510 20423 1518
rect 19701 1452 19711 1510
rect 19769 1504 20423 1510
rect 20481 1510 20491 1518
rect 20791 1510 20825 1584
rect 20859 1578 20935 1584
rect 21037 1578 21113 1584
rect 21147 1510 21181 1584
rect 20481 1504 21135 1510
rect 19769 1470 20079 1504
rect 20113 1470 20423 1504
rect 20481 1470 20791 1504
rect 20825 1470 21135 1504
rect 19769 1464 20423 1470
rect 19769 1452 19779 1464
rect 20413 1460 20423 1464
rect 20481 1464 21135 1470
rect 20481 1460 20491 1464
rect 21125 1452 21135 1464
rect 21193 1452 21203 1510
rect 19523 1301 19533 1359
rect 19591 1348 19601 1359
rect 20234 1348 20244 1359
rect 19591 1342 20244 1348
rect 20302 1348 20312 1359
rect 20947 1348 20957 1360
rect 20302 1342 20957 1348
rect 19591 1308 19901 1342
rect 19935 1308 20244 1342
rect 20302 1308 20613 1342
rect 20647 1308 20957 1342
rect 19591 1302 20244 1308
rect 19591 1301 19601 1302
rect 20234 1301 20244 1302
rect 20302 1302 20957 1308
rect 21015 1302 21025 1360
rect 20302 1301 20312 1302
rect 19613 1228 19689 1234
rect 19791 1228 19867 1234
rect 19969 1228 20045 1234
rect 20147 1228 20223 1234
rect 20325 1228 20401 1234
rect 20503 1228 20579 1234
rect 20681 1228 20757 1234
rect 20859 1228 20935 1234
rect 21037 1228 21113 1234
rect 19613 1220 19625 1228
rect 19609 1194 19625 1220
rect 19677 1194 19803 1228
rect 19855 1194 19981 1228
rect 20033 1194 20159 1228
rect 20211 1194 20337 1228
rect 20389 1194 20515 1228
rect 20567 1194 20693 1228
rect 20745 1194 20871 1228
rect 20923 1194 21049 1228
rect 21101 1220 21196 1228
rect 21360 1220 21488 1592
rect 21101 1194 22312 1220
rect 19609 1120 22312 1194
rect 19609 1092 19625 1120
rect 19613 1086 19625 1092
rect 19677 1086 19803 1120
rect 19855 1086 19981 1120
rect 20033 1086 20159 1120
rect 20211 1086 20337 1120
rect 20389 1086 20515 1120
rect 20567 1086 20693 1120
rect 20745 1086 20871 1120
rect 20923 1086 21049 1120
rect 21101 1092 22312 1120
rect 21101 1086 21196 1092
rect 19613 1080 19689 1086
rect 19723 1012 19757 1086
rect 19791 1080 19867 1086
rect 19969 1080 20045 1086
rect 20079 1012 20113 1086
rect 20147 1080 20223 1086
rect 20325 1080 20401 1086
rect 20435 1020 20469 1086
rect 20503 1080 20579 1086
rect 20681 1080 20757 1086
rect 20413 1012 20423 1020
rect 19701 954 19711 1012
rect 19769 1006 20423 1012
rect 20481 1012 20491 1020
rect 20791 1012 20825 1086
rect 20859 1080 20935 1086
rect 21037 1080 21113 1086
rect 21147 1012 21181 1086
rect 20481 1006 21135 1012
rect 19769 972 20079 1006
rect 20113 972 20423 1006
rect 20481 972 20791 1006
rect 20825 972 21135 1006
rect 19769 966 20423 972
rect 19769 954 19779 966
rect 20413 962 20423 966
rect 20481 966 21135 972
rect 20481 962 20491 966
rect 21125 954 21135 966
rect 21193 954 21203 1012
rect 19523 804 19533 862
rect 19591 850 19601 862
rect 19879 850 19889 857
rect 19591 804 19889 850
rect 19947 850 19957 857
rect 20235 850 20245 855
rect 19879 799 19889 804
rect 19947 804 20245 850
rect 20303 850 20313 855
rect 20591 850 20601 858
rect 19947 799 19957 804
rect 20235 797 20245 804
rect 20303 804 20601 850
rect 20659 850 20669 858
rect 20947 850 20957 862
rect 20303 797 20313 804
rect 20591 800 20601 804
rect 20659 804 20957 850
rect 21015 804 21025 862
rect 20659 800 20669 804
rect 19613 730 19689 736
rect 19791 730 19867 736
rect 19969 730 20045 736
rect 20147 730 20223 736
rect 20325 730 20401 736
rect 20503 730 20579 736
rect 20681 730 20757 736
rect 20859 730 20935 736
rect 21037 730 21113 736
rect 21360 730 21488 1092
rect 19613 696 19625 730
rect 19677 696 19803 730
rect 19855 696 19981 730
rect 20033 696 20159 730
rect 20211 696 20337 730
rect 20389 696 20515 730
rect 20567 696 20693 730
rect 20745 696 20871 730
rect 20923 696 21049 730
rect 21101 696 21488 730
rect 19613 690 19689 696
rect 19791 690 19867 696
rect 19969 690 20045 696
rect 20147 690 20223 696
rect 20325 690 20401 696
rect 20503 690 20579 696
rect 20681 690 20757 696
rect 20859 690 20935 696
rect 21037 690 21113 696
rect 19523 634 19533 640
rect 19337 628 19533 634
rect 19591 634 19601 640
rect 19879 634 19889 639
rect 19591 628 19889 634
rect 19947 634 19957 639
rect 20235 634 20245 642
rect 19947 628 20245 634
rect 20303 634 20313 642
rect 20591 634 20601 640
rect 20303 628 20601 634
rect 20659 634 20669 640
rect 20947 634 20957 639
rect 20659 628 20957 634
rect 21015 635 21025 639
rect 21015 634 21146 635
rect 21015 628 21389 634
rect 19337 594 19349 628
rect 21377 594 21389 628
rect 19337 588 19533 594
rect 19489 582 19533 588
rect 19591 582 19889 594
rect 19489 581 19889 582
rect 19947 584 20245 594
rect 20303 584 20601 594
rect 19947 582 20601 584
rect 20659 582 20957 594
rect 19947 581 20957 582
rect 21015 588 21389 594
rect 21015 581 21146 588
rect 19489 149 19617 581
rect 20212 149 20340 581
rect 20918 149 21046 581
rect 87 148 22071 149
rect 87 141 21891 148
rect 87 139 4818 141
rect 87 134 2500 139
rect 87 71 1419 134
rect 1609 71 2500 134
rect 2690 71 4818 139
rect 5008 139 8217 141
rect 5008 71 5891 139
rect 6071 71 8217 139
rect 8355 139 21891 141
rect 8355 129 10910 139
rect 8355 71 9273 129
rect 9440 71 10910 129
rect 11036 129 21891 139
rect 11036 122 14118 129
rect 11036 71 11978 122
rect 12097 71 14118 122
rect 87 22 304 71
rect 13205 70 14118 71
rect 13205 22 13476 70
rect 14211 127 21891 129
rect 14211 123 16542 127
rect 14211 70 15279 123
rect 15372 70 16542 123
rect 16635 122 21891 127
rect 16635 70 17969 122
rect 18062 70 21891 122
rect 87 21 8217 22
rect 292 20 8217 21
rect 8355 20 9273 22
rect 292 16 9273 20
rect 9263 13 9273 16
rect 9440 21 13476 22
rect 18366 21 21891 70
rect 9440 16 13217 21
rect 9440 13 9450 16
rect 13464 15 18378 21
rect 21885 20 21891 21
rect 22019 21 22071 148
rect 22019 20 22025 21
<< via1 >>
rect 7286 18835 7350 18847
rect 7286 18801 7303 18835
rect 7303 18801 7337 18835
rect 7337 18801 7350 18835
rect 7286 18783 7350 18801
rect 8246 18835 8310 18847
rect 8246 18801 8262 18835
rect 8262 18801 8296 18835
rect 8296 18801 8310 18835
rect 8246 18783 8310 18801
rect 20216 18837 20280 18851
rect 20216 18803 20224 18837
rect 20224 18803 20258 18837
rect 20258 18803 20280 18837
rect 20216 18787 20280 18803
rect 21180 18835 21244 18854
rect 21180 18801 21192 18835
rect 21192 18801 21226 18835
rect 21226 18801 21244 18835
rect 21180 18790 21244 18801
rect 8229 18290 8293 18354
rect 7292 18023 7356 18041
rect 7292 17989 7303 18023
rect 7303 17989 7337 18023
rect 7337 17989 7356 18023
rect 7292 17977 7356 17989
rect 8247 18024 8311 18037
rect 8247 17990 8264 18024
rect 8264 17990 8298 18024
rect 8298 17990 8311 18024
rect 8247 17973 8311 17990
rect 17762 18292 17826 18356
rect 7287 17036 7351 17051
rect 7287 17002 7303 17036
rect 7303 17002 7337 17036
rect 7337 17002 7351 17036
rect 7287 16987 7351 17002
rect 8249 17035 8313 17054
rect 8249 17001 8263 17035
rect 8263 17001 8297 17035
rect 8297 17001 8313 17035
rect 8249 16990 8313 17001
rect 5457 13073 5869 13485
rect 8223 16490 8287 16554
rect 12699 17071 12763 17135
rect 7290 16223 7354 16240
rect 7290 16189 7304 16223
rect 7304 16189 7338 16223
rect 7338 16189 7354 16223
rect 7290 16176 7354 16189
rect 8248 16223 8312 16240
rect 8248 16189 8261 16223
rect 8261 16189 8295 16223
rect 8295 16189 8312 16223
rect 8248 16176 8312 16189
rect 10594 16488 10658 16552
rect 7286 15235 7350 15250
rect 7286 15201 7301 15235
rect 7301 15201 7335 15235
rect 7335 15201 7350 15235
rect 7286 15186 7350 15201
rect 8247 15235 8311 15250
rect 8247 15201 8265 15235
rect 8265 15201 8299 15235
rect 8299 15201 8311 15235
rect 8247 15186 8311 15201
rect 6815 14170 6910 14689
rect 8227 14690 8291 14754
rect 7288 14423 7352 14437
rect 7288 14389 7304 14423
rect 7304 14389 7338 14423
rect 7338 14389 7352 14423
rect 7288 14373 7352 14389
rect 8250 14424 8314 14440
rect 8250 14390 8263 14424
rect 8263 14390 8297 14424
rect 8297 14390 8314 14424
rect 8250 14376 8314 14390
rect 10637 14689 10701 14753
rect 20215 18024 20279 18035
rect 20215 17990 20233 18024
rect 20233 17990 20267 18024
rect 20267 17990 20279 18024
rect 20215 17971 20279 17990
rect 21182 18026 21246 18038
rect 21182 17992 21196 18026
rect 21196 17992 21230 18026
rect 21230 17992 21246 18026
rect 21182 17974 21246 17992
rect 20219 17039 20283 17055
rect 20219 17005 20229 17039
rect 20229 17005 20263 17039
rect 20263 17005 20283 17039
rect 20219 16991 20283 17005
rect 21179 17035 21243 17053
rect 21179 17001 21194 17035
rect 21194 17001 21228 17035
rect 21228 17001 21243 17035
rect 21179 16989 21243 17001
rect 17775 16490 17839 16554
rect 14228 16153 14292 16217
rect 20218 16226 20282 16239
rect 20218 16192 20229 16226
rect 20229 16192 20263 16226
rect 20263 16192 20282 16226
rect 20218 16175 20282 16192
rect 21177 16228 21241 16238
rect 21177 16194 21194 16228
rect 21194 16194 21228 16228
rect 21228 16194 21241 16228
rect 21177 16174 21241 16194
rect 14228 15679 14292 15743
rect 14839 15523 14903 15587
rect 17237 15527 17301 15591
rect 14177 15158 14241 15222
rect 20218 15235 20282 15253
rect 20218 15201 20235 15235
rect 20235 15201 20269 15235
rect 20269 15201 20282 15235
rect 20218 15189 20282 15201
rect 21179 15235 21243 15252
rect 21179 15201 21196 15235
rect 21196 15201 21230 15235
rect 21230 15201 21243 15235
rect 21179 15188 21243 15201
rect 16278 14985 16342 15049
rect 14379 14807 14443 14871
rect 11404 14078 11468 14142
rect 12702 14078 12766 14142
rect 11404 13749 11468 13813
rect 7285 13436 7349 13448
rect 7285 13402 7304 13436
rect 7304 13402 7338 13436
rect 7338 13402 7349 13436
rect 7285 13384 7349 13402
rect 8252 13436 8316 13450
rect 8252 13402 8262 13436
rect 8262 13402 8296 13436
rect 8296 13402 8316 13436
rect 8252 13386 8316 13402
rect 8224 12890 8288 12954
rect 7287 12623 7351 12640
rect 7287 12589 7301 12623
rect 7301 12589 7335 12623
rect 7335 12589 7351 12623
rect 7287 12576 7351 12589
rect 8253 12623 8317 12642
rect 8253 12589 8264 12623
rect 8264 12589 8298 12623
rect 8298 12589 8317 12623
rect 8253 12578 8317 12589
rect 10637 12886 10701 12950
rect 17830 14690 17894 14754
rect 20217 14422 20281 14437
rect 20217 14388 20231 14422
rect 20231 14388 20265 14422
rect 20265 14388 20281 14422
rect 20217 14373 20281 14388
rect 21180 14426 21244 14442
rect 21180 14392 21200 14426
rect 21200 14392 21234 14426
rect 21234 14392 21244 14426
rect 21180 14378 21244 14392
rect 15945 14237 16009 14301
rect 20218 13439 20282 13450
rect 20218 13405 20231 13439
rect 20231 13405 20265 13439
rect 20265 13405 20282 13439
rect 20218 13386 20282 13405
rect 21178 13439 21242 13450
rect 21178 13405 21192 13439
rect 21192 13405 21226 13439
rect 21226 13405 21242 13439
rect 21178 13386 21242 13405
rect 17835 12892 17899 12956
rect 14379 12818 14443 12882
rect 20215 12624 20279 12636
rect 20215 12590 20229 12624
rect 20229 12590 20263 12624
rect 20263 12590 20279 12624
rect 20215 12572 20279 12590
rect 21180 12620 21244 12638
rect 21180 12586 21196 12620
rect 21196 12586 21230 12620
rect 21230 12586 21244 12620
rect 21180 12574 21244 12586
rect 13401 12235 13465 12299
rect 6348 11514 6458 11637
rect 7287 11635 7351 11651
rect 7287 11601 7301 11635
rect 7301 11601 7335 11635
rect 7335 11601 7351 11635
rect 7287 11587 7351 11601
rect 8250 11636 8314 11651
rect 8250 11602 8262 11636
rect 8262 11602 8296 11636
rect 8296 11602 8314 11636
rect 8250 11587 8314 11602
rect 6335 11102 6747 11514
rect 6348 11097 6458 11102
rect 8231 11092 8295 11156
rect 14673 12121 14737 12185
rect 17223 12121 17287 12185
rect 11241 11936 11305 12000
rect 15397 11936 15461 12000
rect 20217 11639 20281 11649
rect 20217 11605 20231 11639
rect 20231 11605 20265 11639
rect 20265 11605 20281 11639
rect 20217 11585 20281 11605
rect 21182 11633 21246 11650
rect 21182 11599 21196 11633
rect 21196 11599 21230 11633
rect 21230 11599 21246 11633
rect 21182 11586 21246 11599
rect 7287 10823 7351 10837
rect 7287 10789 7300 10823
rect 7300 10789 7334 10823
rect 7334 10789 7351 10823
rect 7287 10773 7351 10789
rect 8250 10823 8314 10841
rect 8250 10789 8262 10823
rect 8262 10789 8296 10823
rect 8296 10789 8314 10823
rect 8250 10777 8314 10789
rect 17771 11088 17835 11152
rect 21885 11539 21996 11732
rect 21885 11429 21997 11539
rect 21885 11225 21996 11429
rect 20217 10819 20281 10838
rect 20217 10785 20231 10819
rect 20231 10785 20265 10819
rect 20265 10785 20281 10819
rect 20217 10774 20281 10785
rect 21179 10824 21243 10839
rect 21179 10790 21190 10824
rect 21190 10790 21224 10824
rect 21224 10790 21243 10824
rect 21179 10775 21243 10790
rect 7287 9834 7351 9851
rect 7287 9800 7302 9834
rect 7302 9800 7336 9834
rect 7336 9800 7351 9834
rect 7287 9787 7351 9800
rect 8248 9837 8312 9852
rect 8248 9803 8262 9837
rect 8262 9803 8296 9837
rect 8296 9803 8312 9837
rect 8248 9788 8312 9803
rect 20219 9835 20283 9850
rect 20219 9801 20233 9835
rect 20233 9801 20267 9835
rect 20267 9801 20283 9835
rect 20219 9786 20283 9801
rect 21179 9839 21243 9850
rect 21179 9805 21194 9839
rect 21194 9805 21228 9839
rect 21228 9805 21243 9839
rect 21179 9786 21243 9805
rect 8232 9291 8296 9355
rect 10569 9294 10633 9358
rect 17789 9296 17853 9360
rect 7290 9026 7354 9037
rect 7290 8992 7303 9026
rect 7303 8992 7337 9026
rect 7337 8992 7354 9026
rect 7290 8973 7354 8992
rect 8247 9026 8311 9039
rect 8247 8992 8260 9026
rect 8260 8992 8294 9026
rect 8294 8992 8311 9026
rect 8247 8975 8311 8992
rect 22399 9295 22509 9835
rect 20216 9023 20280 9040
rect 20216 8989 20237 9023
rect 20237 8989 20271 9023
rect 20271 8989 20280 9023
rect 20216 8976 20280 8989
rect 21181 9021 21245 9039
rect 21181 8987 21196 9021
rect 21196 8987 21230 9021
rect 21230 8987 21245 9021
rect 21181 8975 21245 8987
rect 8256 6991 8314 7002
rect 9324 6991 9382 7005
rect 10942 6991 11000 7002
rect 12010 6991 12068 7007
rect 8256 6957 8314 6991
rect 9324 6957 9382 6991
rect 10942 6957 11000 6991
rect 12010 6957 12068 6991
rect 8256 6944 8314 6957
rect 9324 6947 9382 6957
rect 10942 6944 11000 6957
rect 12010 6949 12068 6957
rect 14862 6608 14874 6666
rect 14874 6608 14908 6666
rect 14908 6608 14920 6666
rect 8078 6597 8136 6598
rect 9502 6597 9560 6603
rect 8078 6563 8090 6597
rect 8090 6563 8124 6597
rect 8124 6563 8136 6597
rect 9502 6563 9514 6597
rect 9514 6563 9548 6597
rect 9548 6563 9560 6597
rect 8078 6540 8136 6563
rect 9502 6545 9560 6563
rect 12188 6597 12246 6604
rect 10764 6563 10776 6597
rect 10776 6563 10810 6597
rect 10810 6563 10822 6597
rect 12188 6563 12200 6597
rect 12200 6563 12234 6597
rect 12234 6563 12246 6597
rect 10764 6539 10822 6563
rect 12188 6546 12246 6563
rect 15218 6608 15230 6666
rect 15230 6608 15264 6666
rect 15264 6608 15276 6666
rect 15040 6410 15052 6468
rect 15052 6410 15086 6468
rect 15086 6410 15098 6468
rect 15574 6608 15586 6666
rect 15586 6608 15620 6666
rect 15620 6608 15632 6666
rect 15396 6410 15408 6468
rect 15408 6410 15442 6468
rect 15442 6410 15454 6468
rect 15930 6608 15942 6666
rect 15942 6608 15976 6666
rect 15976 6608 15988 6666
rect 17063 6608 17074 6666
rect 17074 6608 17108 6666
rect 17108 6608 17121 6666
rect 15752 6410 15764 6468
rect 15764 6410 15798 6468
rect 15798 6410 15810 6468
rect 17418 6608 17430 6666
rect 17430 6608 17464 6666
rect 17464 6608 17476 6666
rect 17240 6410 17252 6468
rect 17252 6410 17286 6468
rect 17286 6410 17298 6468
rect 17774 6608 17786 6666
rect 17786 6608 17820 6666
rect 17820 6608 17832 6666
rect 17596 6410 17608 6467
rect 17608 6410 17642 6467
rect 17642 6410 17654 6467
rect 17596 6409 17654 6410
rect 18130 6608 18142 6666
rect 18142 6608 18176 6666
rect 18176 6608 18188 6666
rect 19262 6608 19274 6666
rect 19274 6608 19308 6666
rect 19308 6608 19320 6666
rect 17952 6410 17964 6468
rect 17964 6410 17998 6468
rect 17998 6410 18010 6468
rect 19618 6608 19630 6666
rect 19630 6608 19664 6666
rect 19664 6608 19676 6666
rect 19440 6410 19452 6468
rect 19452 6410 19486 6468
rect 19486 6410 19498 6468
rect 19974 6608 19986 6666
rect 19986 6608 20020 6666
rect 20020 6608 20032 6666
rect 19796 6410 19808 6468
rect 19808 6410 19842 6468
rect 19842 6410 19854 6468
rect 20330 6608 20342 6666
rect 20342 6608 20376 6666
rect 20376 6608 20388 6666
rect 20152 6410 20164 6468
rect 20164 6410 20198 6468
rect 20198 6410 20210 6468
rect 8256 6375 8314 6393
rect 9324 6375 9382 6393
rect 8256 6341 8268 6375
rect 8268 6341 8302 6375
rect 8302 6341 8314 6375
rect 9324 6341 9336 6375
rect 9336 6341 9370 6375
rect 9370 6341 9382 6375
rect 8256 6335 8314 6341
rect 9324 6335 9382 6341
rect 10942 6375 11000 6393
rect 12010 6375 12068 6393
rect 10942 6341 10954 6375
rect 10954 6341 10988 6375
rect 10988 6341 11000 6375
rect 12010 6341 12022 6375
rect 12022 6341 12056 6375
rect 12056 6341 12068 6375
rect 10942 6335 11000 6341
rect 12010 6335 12068 6341
rect 20241 6351 20299 6357
rect 20241 6317 20244 6351
rect 20244 6317 20296 6351
rect 20296 6317 20299 6351
rect 12446 6248 12458 6280
rect 12458 6248 12510 6280
rect 12510 6248 12525 6280
rect 9768 6151 9826 6209
rect 10497 6151 10555 6209
rect 12446 6113 12525 6248
rect 12446 6080 12458 6113
rect 12458 6080 12510 6113
rect 12510 6080 12525 6113
rect 20241 6299 20299 6317
rect 12844 6111 12957 6228
rect 8078 6019 8136 6025
rect 8722 6019 8914 6032
rect 9502 6019 9560 6025
rect 8078 5985 8090 6019
rect 8090 5985 8124 6019
rect 8124 5985 8136 6019
rect 8722 5985 8802 6019
rect 8802 5985 8836 6019
rect 8836 5985 8914 6019
rect 9502 5985 9514 6019
rect 9514 5985 9548 6019
rect 9548 5985 9560 6019
rect 8078 5967 8136 5985
rect 8722 5974 8914 5985
rect 8790 5967 8848 5974
rect 9502 5967 9560 5985
rect 10764 6020 10822 6026
rect 11408 6020 11600 6030
rect 12188 6020 12246 6026
rect 10764 5986 10776 6020
rect 10776 5986 10810 6020
rect 10810 5986 10822 6020
rect 11408 5986 11488 6020
rect 11488 5986 11522 6020
rect 11522 5986 11600 6020
rect 12188 5986 12200 6020
rect 12200 5986 12234 6020
rect 12234 5986 12246 6020
rect 10764 5968 10822 5986
rect 11408 5972 11600 5986
rect 11476 5968 11534 5972
rect 12188 5968 12246 5986
rect 14863 5841 14875 5899
rect 14875 5841 14909 5899
rect 14909 5841 14921 5899
rect 8256 5797 8314 5815
rect 9324 5797 9382 5815
rect 8256 5763 8268 5797
rect 8268 5763 8302 5797
rect 8302 5763 8314 5797
rect 9324 5763 9336 5797
rect 9336 5763 9370 5797
rect 9370 5763 9382 5797
rect 8256 5757 8314 5763
rect 9324 5757 9382 5763
rect 10942 5798 11000 5816
rect 12010 5798 12068 5816
rect 10942 5764 10954 5798
rect 10954 5764 10988 5798
rect 10988 5764 11000 5798
rect 12010 5764 12022 5798
rect 12022 5764 12056 5798
rect 12056 5764 12068 5798
rect 10942 5758 11000 5764
rect 12010 5758 12068 5764
rect 15219 5841 15231 5899
rect 15231 5841 15265 5899
rect 15265 5841 15277 5899
rect 15041 5643 15053 5701
rect 15053 5643 15087 5701
rect 15087 5643 15099 5701
rect 15575 5841 15587 5899
rect 15587 5841 15621 5899
rect 15621 5841 15633 5899
rect 15397 5643 15409 5701
rect 15409 5643 15443 5701
rect 15443 5643 15455 5701
rect 15931 5841 15943 5899
rect 15943 5841 15977 5899
rect 15977 5841 15989 5899
rect 17063 5841 17075 5899
rect 17075 5841 17109 5899
rect 17109 5841 17121 5899
rect 15752 5643 15765 5701
rect 15765 5643 15799 5701
rect 15799 5643 15810 5701
rect 17419 5841 17431 5899
rect 17431 5841 17465 5899
rect 17465 5841 17477 5899
rect 17242 5643 17253 5701
rect 17253 5643 17287 5701
rect 17287 5643 17300 5701
rect 17775 5841 17787 5899
rect 17787 5841 17821 5899
rect 17821 5841 17833 5899
rect 17597 5643 17609 5701
rect 17609 5643 17643 5701
rect 17643 5643 17655 5701
rect 18131 5841 18143 5899
rect 18143 5841 18177 5899
rect 18177 5841 18189 5899
rect 19264 5841 19275 5899
rect 19275 5841 19309 5899
rect 19309 5841 19322 5899
rect 17953 5643 17965 5701
rect 17965 5643 17999 5701
rect 17999 5643 18011 5701
rect 19619 5841 19631 5899
rect 19631 5841 19665 5899
rect 19665 5841 19677 5899
rect 19442 5643 19453 5701
rect 19453 5643 19487 5701
rect 19487 5643 19500 5701
rect 19975 5841 19987 5899
rect 19987 5841 20021 5899
rect 20021 5841 20033 5899
rect 19797 5643 19809 5701
rect 19809 5643 19843 5701
rect 19843 5643 19855 5701
rect 20331 5841 20343 5899
rect 20343 5841 20377 5899
rect 20377 5841 20462 5899
rect 20153 5643 20165 5701
rect 20165 5643 20199 5701
rect 20199 5643 20211 5701
rect 19353 5584 19411 5590
rect 19353 5550 19355 5584
rect 19355 5550 19407 5584
rect 19407 5550 19411 5584
rect 19353 5532 19411 5550
rect 2829 4263 2887 4321
rect 4609 4263 4667 4321
rect 8078 5139 8136 5145
rect 9858 5139 9916 5145
rect 8078 5105 8090 5139
rect 8090 5105 8124 5139
rect 8124 5105 8136 5139
rect 9858 5105 9870 5139
rect 9870 5105 9904 5139
rect 9904 5105 9916 5139
rect 8078 5087 8136 5105
rect 9858 5087 9916 5105
rect 10408 5139 10466 5145
rect 12188 5139 12246 5145
rect 10408 5105 10420 5139
rect 10420 5105 10454 5139
rect 10454 5105 10466 5139
rect 12188 5105 12200 5139
rect 12200 5105 12234 5139
rect 12234 5105 12246 5139
rect 10408 5087 10466 5105
rect 12188 5087 12246 5105
rect 13894 5047 13952 5053
rect 16030 5047 16088 5053
rect 18131 5047 18248 5057
rect 13894 5013 13906 5047
rect 13906 5013 13940 5047
rect 13940 5013 13952 5047
rect 16030 5013 16042 5047
rect 16042 5013 16076 5047
rect 16076 5013 16088 5047
rect 18131 5013 18178 5047
rect 18178 5013 18212 5047
rect 18212 5013 18248 5047
rect 13894 4995 13952 5013
rect 16030 4995 16088 5013
rect 18131 4940 18248 5013
rect 8256 4917 8314 4935
rect 8790 4931 8848 4935
rect 8256 4883 8268 4917
rect 8268 4883 8302 4917
rect 8302 4883 8314 4917
rect 8256 4877 8314 4883
rect 8725 4873 8917 4931
rect 9680 4917 9738 4935
rect 9680 4883 9692 4917
rect 9692 4883 9726 4917
rect 9726 4883 9738 4917
rect 9680 4877 9738 4883
rect 10586 4917 10644 4935
rect 11476 4932 11534 4935
rect 10586 4883 10598 4917
rect 10598 4883 10632 4917
rect 10632 4883 10644 4917
rect 10586 4877 10644 4883
rect 11404 4874 11596 4932
rect 12010 4917 12068 4935
rect 12010 4883 12022 4917
rect 12022 4883 12056 4917
rect 12056 4883 12068 4917
rect 12010 4877 12068 4883
rect 13716 4825 13774 4843
rect 15852 4825 15910 4843
rect 17988 4825 18046 4843
rect 13716 4791 13728 4825
rect 13728 4791 13762 4825
rect 13762 4791 13774 4825
rect 15852 4791 15864 4825
rect 15864 4791 15898 4825
rect 15898 4791 15910 4825
rect 17988 4791 18000 4825
rect 18000 4791 18034 4825
rect 18034 4791 18046 4825
rect 13716 4785 13774 4791
rect 15852 4785 15910 4791
rect 17988 4785 18046 4791
rect 8078 4569 8136 4575
rect 8725 4569 8917 4577
rect 9858 4569 9916 4575
rect 8078 4535 8090 4569
rect 8090 4535 8124 4569
rect 8124 4535 8136 4569
rect 8725 4535 8802 4569
rect 8802 4535 8836 4569
rect 8836 4535 8917 4569
rect 9858 4535 9870 4569
rect 9870 4535 9904 4569
rect 9904 4535 9916 4569
rect 8078 4517 8136 4535
rect 8725 4519 8917 4535
rect 8790 4517 8848 4519
rect 9858 4517 9916 4535
rect 10408 4569 10466 4575
rect 11406 4569 11598 4576
rect 12188 4569 12246 4575
rect 10408 4535 10420 4569
rect 10420 4535 10454 4569
rect 10454 4535 10466 4569
rect 11406 4535 11488 4569
rect 11488 4535 11522 4569
rect 11522 4535 11598 4569
rect 12188 4535 12200 4569
rect 12200 4535 12234 4569
rect 12234 4535 12246 4569
rect 10408 4517 10466 4535
rect 11406 4518 11598 4535
rect 11478 4517 11536 4518
rect 12188 4517 12246 4535
rect 13894 4547 13952 4553
rect 16030 4547 16088 4553
rect 18132 4547 18249 4553
rect 13894 4513 13906 4547
rect 13906 4513 13940 4547
rect 13940 4513 13952 4547
rect 16030 4513 16042 4547
rect 16042 4513 16076 4547
rect 16076 4513 16088 4547
rect 18132 4513 18178 4547
rect 18178 4513 18212 4547
rect 18212 4513 18249 4547
rect 13894 4495 13952 4513
rect 16030 4495 16088 4513
rect 18132 4436 18249 4513
rect 8256 4347 8314 4365
rect 9680 4347 9738 4365
rect 8256 4313 8268 4347
rect 8268 4313 8302 4347
rect 8302 4313 8314 4347
rect 9680 4313 9692 4347
rect 9692 4313 9726 4347
rect 9726 4313 9738 4347
rect 8256 4307 8314 4313
rect 9680 4307 9738 4313
rect 10586 4347 10644 4365
rect 12010 4347 12068 4365
rect 10586 4313 10598 4347
rect 10598 4313 10632 4347
rect 10632 4313 10644 4347
rect 12010 4313 12022 4347
rect 12022 4313 12056 4347
rect 12056 4313 12068 4347
rect 10586 4307 10644 4313
rect 12010 4307 12068 4313
rect 13716 4325 13774 4343
rect 15852 4325 15910 4343
rect 17630 4325 17752 4387
rect 13716 4291 13728 4325
rect 13728 4291 13762 4325
rect 13762 4291 13774 4325
rect 15852 4291 15864 4325
rect 15864 4291 15898 4325
rect 15898 4291 15910 4325
rect 17630 4291 17644 4325
rect 17644 4291 17678 4325
rect 17678 4291 17752 4325
rect 13716 4285 13774 4291
rect 15852 4285 15910 4291
rect 17630 4286 17752 4291
rect 17988 4325 18046 4343
rect 17988 4291 18000 4325
rect 18000 4291 18034 4325
rect 18034 4291 18046 4325
rect 17630 4285 17688 4286
rect 17988 4285 18046 4291
rect 3404 4219 3569 4227
rect 3404 4185 3420 4219
rect 3420 4185 3454 4219
rect 3454 4185 3569 4219
rect 3404 4173 3569 4185
rect 4128 4219 4293 4228
rect 4128 4185 4140 4219
rect 4140 4185 4174 4219
rect 4174 4185 4293 4219
rect 4128 4174 4293 4185
rect 17452 4183 17510 4241
rect 2256 4037 2522 4049
rect 2256 4003 2262 4037
rect 2262 4003 2296 4037
rect 2296 4003 2474 4037
rect 2474 4003 2508 4037
rect 2508 4003 2522 4037
rect 2256 3995 2522 4003
rect 4884 4037 5150 4051
rect 4884 4003 4890 4037
rect 4890 4003 4924 4037
rect 4924 4003 5102 4037
rect 5102 4003 5136 4037
rect 5136 4003 5150 4037
rect 4884 3997 5150 4003
rect 2829 3903 2887 3961
rect 4609 3903 4667 3961
rect 657 3692 767 3802
rect 17630 4007 17752 4125
rect 7723 3639 7781 3645
rect 8718 3639 8910 3645
rect 9859 3639 9917 3645
rect 7723 3605 7735 3639
rect 7735 3605 7769 3639
rect 7769 3605 7781 3639
rect 8718 3605 8803 3639
rect 8803 3605 8837 3639
rect 8837 3605 8910 3639
rect 9859 3605 9871 3639
rect 9871 3605 9905 3639
rect 9905 3605 9917 3639
rect 7723 3587 7781 3605
rect 8718 3587 8910 3605
rect 9859 3587 9917 3605
rect 10410 3639 10468 3645
rect 11414 3639 11606 3646
rect 12546 3639 12604 3645
rect 10410 3605 10422 3639
rect 10422 3605 10456 3639
rect 10456 3605 10468 3639
rect 11414 3605 11490 3639
rect 11490 3605 11524 3639
rect 11524 3605 11606 3639
rect 12546 3605 12558 3639
rect 12558 3605 12592 3639
rect 12592 3605 12604 3639
rect 10410 3587 10468 3605
rect 11414 3588 11606 3605
rect 11478 3587 11536 3588
rect 12546 3587 12604 3605
rect 17452 3593 17510 3651
rect 17631 3549 17752 3550
rect 17630 3543 17752 3549
rect 594 3439 652 3445
rect 2018 3439 2076 3445
rect 594 3405 606 3439
rect 606 3405 640 3439
rect 640 3405 652 3439
rect 2018 3405 2030 3439
rect 2030 3405 2064 3439
rect 2064 3405 2076 3439
rect 594 3387 652 3405
rect 2018 3387 2076 3405
rect 2256 3439 2522 3445
rect 3442 3439 3500 3445
rect 2256 3405 2386 3439
rect 2386 3405 2420 3439
rect 2420 3405 2522 3439
rect 3442 3405 3454 3439
rect 3454 3405 3488 3439
rect 3488 3405 3500 3439
rect 2256 3391 2522 3405
rect 3442 3387 3500 3405
rect 3994 3439 4052 3445
rect 4886 3439 5152 3448
rect 3994 3405 4006 3439
rect 4006 3405 4040 3439
rect 4040 3405 4052 3439
rect 4886 3405 5074 3439
rect 5074 3405 5108 3439
rect 5108 3405 5152 3439
rect 3994 3387 4052 3405
rect 4886 3394 5152 3405
rect 5418 3439 5476 3445
rect 6842 3439 6900 3445
rect 5418 3405 5430 3439
rect 5430 3405 5464 3439
rect 5464 3405 5476 3439
rect 6842 3405 6854 3439
rect 6854 3405 6888 3439
rect 6888 3405 6900 3439
rect 5418 3387 5476 3405
rect 6842 3387 6900 3405
rect 8257 3417 8315 3435
rect 9325 3417 9383 3435
rect 8257 3383 8269 3417
rect 8269 3383 8303 3417
rect 8303 3383 8315 3417
rect 9325 3383 9337 3417
rect 9337 3383 9371 3417
rect 9371 3383 9383 3417
rect 8257 3377 8315 3383
rect 9325 3377 9383 3383
rect 10944 3417 11002 3435
rect 12012 3417 12070 3435
rect 10944 3383 10956 3417
rect 10956 3383 10990 3417
rect 10990 3383 11002 3417
rect 12012 3383 12024 3417
rect 12024 3383 12058 3417
rect 12058 3383 12070 3417
rect 10944 3377 11002 3383
rect 12012 3377 12070 3383
rect 1484 3217 1542 3235
rect 2552 3217 2610 3235
rect 1484 3183 1496 3217
rect 1496 3183 1530 3217
rect 1530 3183 1542 3217
rect 2552 3183 2564 3217
rect 2564 3183 2598 3217
rect 2598 3183 2610 3217
rect 1484 3177 1542 3183
rect 2552 3177 2610 3183
rect 4884 3217 4942 3235
rect 5952 3217 6010 3235
rect 4884 3183 4896 3217
rect 4896 3183 4930 3217
rect 4930 3183 4942 3217
rect 5952 3183 5964 3217
rect 5964 3183 5998 3217
rect 5998 3183 6010 3217
rect 17274 3287 17286 3530
rect 17286 3287 17320 3530
rect 17320 3287 17332 3530
rect 17274 3278 17332 3287
rect 17630 3491 17642 3543
rect 17631 3447 17642 3491
rect 17642 3447 17676 3543
rect 17676 3447 17752 3543
rect 17631 3433 17752 3447
rect 17452 3404 17510 3416
rect 17452 3287 17464 3404
rect 17464 3287 17498 3404
rect 17498 3287 17510 3404
rect 17452 3279 17510 3287
rect 4884 3177 4942 3183
rect 5952 3177 6010 3183
rect 20331 5122 20477 5141
rect 19175 5038 19233 5106
rect 19175 5004 19187 5038
rect 19187 5004 19221 5038
rect 19221 5004 19233 5038
rect 19709 5021 19767 5110
rect 20331 5088 20335 5122
rect 20335 5088 20387 5122
rect 20387 5088 20477 5122
rect 19175 4986 19233 5004
rect 20331 5001 20477 5088
rect 21132 5026 21190 5115
rect 21667 5038 21725 5106
rect 21667 5004 21679 5038
rect 21679 5004 21713 5038
rect 21713 5004 21725 5038
rect 21667 4986 21725 5004
rect 19353 4816 19411 4834
rect 20065 4816 20123 4831
rect 20779 4816 20837 4835
rect 21489 4816 21547 4834
rect 19353 4782 19365 4816
rect 19365 4782 19399 4816
rect 19399 4782 19411 4816
rect 20065 4782 20077 4816
rect 20077 4782 20111 4816
rect 20111 4782 20123 4816
rect 20779 4782 20789 4816
rect 20789 4782 20823 4816
rect 20823 4782 20837 4816
rect 21489 4782 21501 4816
rect 21501 4782 21535 4816
rect 21535 4782 21547 4816
rect 19353 4776 19411 4782
rect 20065 4773 20123 4782
rect 20779 4777 20837 4782
rect 21489 4776 21547 4782
rect 19176 4546 19234 4725
rect 19175 4540 19234 4546
rect 19175 4506 19187 4540
rect 19187 4506 19221 4540
rect 19221 4517 19234 4540
rect 19221 4506 19233 4517
rect 19710 4511 19768 4719
rect 20420 4522 20478 4730
rect 21133 4515 21191 4723
rect 21667 4540 21725 4716
rect 21667 4506 21679 4540
rect 21679 4506 21713 4540
rect 21713 4506 21725 4540
rect 19175 4488 19233 4506
rect 21667 4488 21725 4506
rect 19353 4318 19411 4336
rect 20065 4318 20123 4331
rect 20778 4318 20836 4334
rect 21489 4318 21547 4336
rect 19353 4284 19365 4318
rect 19365 4284 19399 4318
rect 19399 4284 19411 4318
rect 20065 4284 20077 4318
rect 20077 4284 20111 4318
rect 20111 4284 20123 4318
rect 20778 4284 20789 4318
rect 20789 4284 20823 4318
rect 20823 4284 20836 4318
rect 21489 4284 21501 4318
rect 21501 4284 21535 4318
rect 21535 4284 21547 4318
rect 19353 4278 19411 4284
rect 20065 4273 20123 4284
rect 20778 4276 20836 4284
rect 21489 4278 21547 4284
rect 19175 4042 19233 4224
rect 19175 4008 19187 4042
rect 19187 4008 19221 4042
rect 19221 4008 19233 4042
rect 19709 4015 19767 4223
rect 20422 4015 20480 4223
rect 21133 4022 21191 4230
rect 21666 4048 21724 4218
rect 21666 4042 21725 4048
rect 21666 4010 21679 4042
rect 21667 4008 21679 4010
rect 21679 4008 21713 4042
rect 21713 4008 21725 4042
rect 19175 3990 19233 4008
rect 21667 3990 21725 4008
rect 19353 3820 19411 3838
rect 20065 3820 20123 3837
rect 20774 3820 20832 3841
rect 21489 3820 21547 3838
rect 19353 3786 19365 3820
rect 19365 3786 19399 3820
rect 19399 3786 19411 3820
rect 20065 3786 20077 3820
rect 20077 3786 20111 3820
rect 20111 3786 20123 3820
rect 20774 3786 20789 3820
rect 20789 3786 20823 3820
rect 20823 3786 20832 3820
rect 21489 3786 21501 3820
rect 21501 3786 21535 3820
rect 21535 3786 21547 3820
rect 19353 3780 19411 3786
rect 20065 3779 20123 3786
rect 20774 3783 20832 3786
rect 21489 3780 21547 3786
rect 19175 3544 19233 3736
rect 19175 3510 19187 3544
rect 19187 3510 19221 3544
rect 19221 3510 19233 3544
rect 19708 3518 19766 3726
rect 20420 3515 20478 3723
rect 21133 3513 21191 3721
rect 21667 3544 21725 3736
rect 21667 3510 21679 3544
rect 21679 3510 21713 3544
rect 21713 3510 21725 3544
rect 19175 3492 19233 3510
rect 21667 3492 21725 3510
rect 19353 3322 19411 3340
rect 19353 3288 19365 3322
rect 19365 3288 19399 3322
rect 19399 3288 19411 3322
rect 19353 3282 19411 3288
rect 19710 3322 19768 3339
rect 19710 3288 19721 3322
rect 19721 3288 19755 3322
rect 19755 3288 19768 3322
rect 19710 3281 19768 3288
rect 20066 3322 20124 3339
rect 20066 3288 20077 3322
rect 20077 3288 20111 3322
rect 20111 3288 20124 3322
rect 20066 3281 20124 3288
rect 20423 3322 20481 3340
rect 20423 3288 20433 3322
rect 20433 3288 20467 3322
rect 20467 3288 20481 3322
rect 20423 3282 20481 3288
rect 20779 3322 20837 3337
rect 20779 3288 20789 3322
rect 20789 3288 20823 3322
rect 20823 3288 20837 3322
rect 20779 3279 20837 3288
rect 21135 3322 21193 3338
rect 21135 3288 21145 3322
rect 21145 3288 21179 3322
rect 21179 3288 21193 3322
rect 21135 3280 21193 3288
rect 21489 3322 21547 3340
rect 21489 3288 21501 3322
rect 21501 3288 21535 3322
rect 21535 3288 21547 3322
rect 21489 3282 21547 3288
rect 7723 3139 7781 3145
rect 8791 3139 8849 3145
rect 9859 3139 9917 3145
rect 7723 3105 7735 3139
rect 7735 3105 7769 3139
rect 7769 3105 7781 3139
rect 8791 3105 8803 3139
rect 8803 3105 8837 3139
rect 8837 3105 8849 3139
rect 9859 3105 9871 3139
rect 9871 3105 9905 3139
rect 9905 3105 9917 3139
rect 7723 3087 7781 3105
rect 8791 3087 8849 3105
rect 9859 3087 9917 3105
rect 10410 3139 10468 3145
rect 11478 3139 11536 3145
rect 12546 3139 12604 3145
rect 10410 3105 10422 3139
rect 10422 3105 10456 3139
rect 10456 3105 10468 3139
rect 11478 3105 11490 3139
rect 11490 3105 11524 3139
rect 11524 3105 11536 3139
rect 12546 3105 12558 3139
rect 12558 3105 12592 3139
rect 12592 3105 12604 3139
rect 10410 3087 10468 3105
rect 11478 3087 11536 3105
rect 12546 3087 12604 3105
rect 14863 3039 14921 3097
rect 21891 3052 22019 3180
rect 594 2939 652 2945
rect 2018 2939 2076 2945
rect 3442 2939 3500 2945
rect 594 2905 606 2939
rect 606 2905 640 2939
rect 640 2905 652 2939
rect 2018 2905 2030 2939
rect 2030 2905 2064 2939
rect 2064 2905 2076 2939
rect 3442 2905 3454 2939
rect 3454 2905 3488 2939
rect 3488 2905 3500 2939
rect 594 2887 652 2905
rect 2018 2887 2076 2905
rect 3442 2887 3500 2905
rect 3994 2939 4052 2945
rect 5418 2939 5476 2945
rect 6842 2939 6900 2945
rect 3994 2905 4006 2939
rect 4006 2905 4040 2939
rect 4040 2905 4052 2939
rect 5418 2905 5430 2939
rect 5430 2905 5464 2939
rect 5464 2905 5476 2939
rect 6842 2905 6854 2939
rect 6854 2905 6888 2939
rect 6888 2905 6900 2939
rect 3994 2887 4052 2905
rect 5418 2887 5476 2905
rect 6842 2887 6900 2905
rect 8257 2917 8315 2935
rect 9325 2917 9383 2935
rect 8257 2883 8269 2917
rect 8269 2883 8303 2917
rect 8303 2883 8315 2917
rect 9325 2883 9337 2917
rect 9337 2883 9371 2917
rect 9371 2883 9383 2917
rect 8257 2877 8315 2883
rect 9325 2877 9383 2883
rect 10944 2917 11002 2935
rect 12012 2917 12070 2935
rect 10944 2883 10956 2917
rect 10956 2883 10990 2917
rect 10990 2883 11002 2917
rect 12012 2883 12024 2917
rect 12024 2883 12058 2917
rect 12058 2883 12070 2917
rect 10944 2877 11002 2883
rect 12012 2877 12070 2883
rect 1484 2717 1542 2735
rect 2552 2717 2610 2735
rect 1484 2683 1496 2717
rect 1496 2683 1530 2717
rect 1530 2683 1542 2717
rect 2552 2683 2564 2717
rect 2564 2683 2598 2717
rect 2598 2683 2610 2717
rect 1484 2677 1542 2683
rect 2552 2677 2610 2683
rect 4884 2717 4942 2735
rect 5952 2717 6010 2736
rect 4884 2683 4896 2717
rect 4896 2683 4930 2717
rect 4930 2683 4942 2717
rect 5952 2683 5964 2717
rect 5964 2683 5998 2717
rect 5998 2683 6010 2717
rect 4884 2677 4942 2683
rect 5952 2678 6010 2683
rect 7723 2639 7781 2645
rect 8791 2639 8849 2645
rect 9859 2639 9917 2645
rect 7723 2605 7735 2639
rect 7735 2605 7769 2639
rect 7769 2605 7781 2639
rect 8791 2605 8803 2639
rect 8803 2605 8837 2639
rect 8837 2605 8849 2639
rect 9859 2605 9871 2639
rect 9871 2605 9905 2639
rect 9905 2605 9917 2639
rect 7723 2587 7781 2605
rect 8791 2587 8849 2605
rect 9859 2587 9917 2605
rect 10410 2639 10468 2645
rect 11478 2639 11536 2645
rect 12546 2639 12604 2645
rect 10410 2605 10422 2639
rect 10422 2605 10456 2639
rect 10456 2605 10468 2639
rect 11478 2605 11490 2639
rect 11490 2605 11524 2639
rect 11524 2605 11536 2639
rect 12546 2605 12558 2639
rect 12558 2605 12592 2639
rect 12592 2605 12604 2639
rect 10410 2587 10468 2605
rect 11478 2587 11536 2605
rect 12546 2587 12604 2605
rect 17272 2654 17330 2712
rect 594 2439 652 2445
rect 2018 2439 2076 2445
rect 3442 2439 3500 2445
rect 594 2405 606 2439
rect 606 2405 640 2439
rect 640 2405 652 2439
rect 2018 2405 2030 2439
rect 2030 2405 2064 2439
rect 2064 2405 2076 2439
rect 3442 2405 3454 2439
rect 3454 2405 3488 2439
rect 3488 2405 3500 2439
rect 594 2387 652 2405
rect 2018 2387 2076 2405
rect 3442 2387 3500 2405
rect 3994 2439 4052 2445
rect 5418 2439 5476 2445
rect 6842 2439 6900 2445
rect 3994 2405 4006 2439
rect 4006 2405 4040 2439
rect 4040 2405 4052 2439
rect 5418 2405 5430 2439
rect 5430 2405 5464 2439
rect 5464 2405 5476 2439
rect 6842 2405 6854 2439
rect 6854 2405 6888 2439
rect 6888 2405 6900 2439
rect 3994 2387 4052 2405
rect 5418 2387 5476 2405
rect 6842 2387 6900 2405
rect 8257 2417 8315 2435
rect 8257 2383 8269 2417
rect 8269 2383 8303 2417
rect 8303 2383 8315 2417
rect 8257 2377 8315 2383
rect 8609 2417 8800 2426
rect 9325 2417 9383 2435
rect 8609 2383 8625 2417
rect 8625 2383 8659 2417
rect 8659 2383 8800 2417
rect 9325 2383 9337 2417
rect 9337 2383 9371 2417
rect 9371 2383 9383 2417
rect 8609 2373 8800 2383
rect 9325 2377 9383 2383
rect 10944 2417 11002 2435
rect 11546 2417 11752 2426
rect 10944 2383 10956 2417
rect 10956 2383 10990 2417
rect 10990 2383 11002 2417
rect 11546 2383 11668 2417
rect 11668 2383 11702 2417
rect 11702 2383 11752 2417
rect 10944 2377 11002 2383
rect 11546 2368 11752 2383
rect 12012 2417 12070 2435
rect 12012 2383 12024 2417
rect 12024 2383 12058 2417
rect 12058 2383 12070 2417
rect 12012 2377 12070 2383
rect 14134 2480 14146 2538
rect 14146 2480 14180 2538
rect 14180 2480 14192 2538
rect 14426 2480 14438 2538
rect 14438 2480 14472 2538
rect 14472 2480 14484 2538
rect 14718 2480 14730 2538
rect 14730 2480 14764 2538
rect 14764 2480 14776 2538
rect 15010 2480 15022 2538
rect 15022 2480 15056 2538
rect 15056 2480 15068 2538
rect 15302 2480 15314 2538
rect 15314 2480 15348 2538
rect 15348 2480 15360 2538
rect 1484 2217 1542 2235
rect 2552 2217 2610 2235
rect 1484 2183 1496 2217
rect 1496 2183 1530 2217
rect 1530 2183 1542 2217
rect 2552 2183 2564 2217
rect 2564 2183 2598 2217
rect 2598 2183 2610 2217
rect 1484 2177 1542 2183
rect 2552 2177 2610 2183
rect 4884 2217 4942 2235
rect 5952 2217 6010 2235
rect 4884 2183 4896 2217
rect 4896 2183 4930 2217
rect 4930 2183 4942 2217
rect 5952 2183 5964 2217
rect 5964 2183 5998 2217
rect 5998 2183 6010 2217
rect 4884 2177 4942 2183
rect 5952 2177 6010 2183
rect 594 1939 652 1945
rect 2018 1939 2076 1945
rect 3442 1939 3500 1945
rect 594 1905 606 1939
rect 606 1905 640 1939
rect 640 1905 652 1939
rect 2018 1905 2030 1939
rect 2030 1905 2064 1939
rect 2064 1905 2076 1939
rect 3442 1905 3454 1939
rect 3454 1905 3488 1939
rect 3488 1905 3500 1939
rect 594 1887 652 1905
rect 2018 1887 2076 1905
rect 3442 1887 3500 1905
rect 3994 1939 4052 1945
rect 5418 1939 5476 1945
rect 6842 1939 6900 1945
rect 3994 1905 4006 1939
rect 4006 1905 4040 1939
rect 4040 1905 4052 1939
rect 5418 1905 5430 1939
rect 5430 1905 5464 1939
rect 5464 1905 5476 1939
rect 6842 1905 6854 1939
rect 6854 1905 6888 1939
rect 6888 1905 6900 1939
rect 3994 1887 4052 1905
rect 5418 1887 5476 1905
rect 6842 1887 6900 1905
rect 7723 1939 7781 1945
rect 8593 1939 8857 1946
rect 11502 1945 11708 1946
rect 9859 1939 9917 1945
rect 7723 1905 7735 1939
rect 7735 1905 7769 1939
rect 7769 1905 7781 1939
rect 8593 1905 8803 1939
rect 8803 1905 8837 1939
rect 8837 1905 8857 1939
rect 9859 1905 9871 1939
rect 9871 1905 9905 1939
rect 9905 1905 9917 1939
rect 7723 1887 7781 1905
rect 8593 1887 8857 1905
rect 9859 1887 9917 1905
rect 10410 1939 10468 1945
rect 11478 1939 11708 1945
rect 12546 1939 12604 1945
rect 10410 1905 10422 1939
rect 10422 1905 10456 1939
rect 10456 1905 10468 1939
rect 11478 1905 11490 1939
rect 11490 1905 11524 1939
rect 11524 1905 11708 1939
rect 12546 1905 12558 1939
rect 12558 1905 12592 1939
rect 12592 1905 12604 1939
rect 10410 1887 10468 1905
rect 11478 1887 11708 1905
rect 12546 1887 12604 1905
rect 11502 1886 11708 1887
rect 16738 2604 16796 2608
rect 17420 2604 17535 2610
rect 18162 2604 18220 2610
rect 16738 2570 16750 2604
rect 16750 2570 16784 2604
rect 16784 2570 16796 2604
rect 17420 2570 17462 2604
rect 17462 2570 17496 2604
rect 17496 2570 17535 2604
rect 18162 2570 18174 2604
rect 18174 2570 18208 2604
rect 18208 2570 18220 2604
rect 16738 2550 16796 2570
rect 17420 2514 17535 2570
rect 18162 2552 18220 2570
rect 16560 2382 16618 2400
rect 17984 2382 18042 2400
rect 16560 2348 16572 2382
rect 16572 2348 16606 2382
rect 16606 2348 16618 2382
rect 17984 2348 17996 2382
rect 17996 2348 18030 2382
rect 18030 2348 18042 2382
rect 16560 2342 16618 2348
rect 17984 2342 18042 2348
rect 17243 2166 17361 2283
rect 1484 1717 1542 1735
rect 2552 1717 2610 1735
rect 1484 1683 1496 1717
rect 1496 1683 1530 1717
rect 1530 1683 1542 1717
rect 2552 1683 2564 1717
rect 2564 1683 2598 1717
rect 2598 1683 2610 1717
rect 1484 1677 1542 1683
rect 2552 1677 2610 1683
rect 4884 1717 4942 1735
rect 5952 1717 6010 1735
rect 4884 1683 4896 1717
rect 4896 1683 4930 1717
rect 4930 1683 4942 1717
rect 5952 1683 5964 1717
rect 5964 1683 5998 1717
rect 5998 1683 6010 1717
rect 4884 1677 4942 1683
rect 5952 1677 6010 1683
rect 8257 1717 8315 1735
rect 9325 1717 9383 1735
rect 8257 1683 8269 1717
rect 8269 1683 8303 1717
rect 8303 1683 8315 1717
rect 9325 1683 9337 1717
rect 9337 1683 9371 1717
rect 9371 1683 9383 1717
rect 8257 1677 8315 1683
rect 9325 1677 9383 1683
rect 10944 1717 11002 1735
rect 12012 1717 12070 1735
rect 10944 1683 10956 1717
rect 10956 1683 10990 1717
rect 10990 1683 11002 1717
rect 12012 1683 12024 1717
rect 12024 1683 12058 1717
rect 12058 1683 12070 1717
rect 10944 1677 11002 1683
rect 12012 1677 12070 1683
rect 594 1439 652 1445
rect 2018 1439 2076 1445
rect 3442 1439 3500 1445
rect 594 1405 606 1439
rect 606 1405 640 1439
rect 640 1405 652 1439
rect 2018 1405 2030 1439
rect 2030 1405 2064 1439
rect 2064 1405 2076 1439
rect 3442 1405 3454 1439
rect 3454 1405 3488 1439
rect 3488 1405 3500 1439
rect 594 1387 652 1405
rect 2018 1387 2076 1405
rect 3442 1387 3500 1405
rect 3994 1439 4052 1445
rect 5418 1439 5476 1445
rect 6842 1439 6900 1445
rect 3994 1405 4006 1439
rect 4006 1405 4040 1439
rect 4040 1405 4052 1439
rect 5418 1405 5430 1439
rect 5430 1405 5464 1439
rect 5464 1405 5476 1439
rect 6842 1405 6854 1439
rect 6854 1405 6888 1439
rect 6888 1405 6900 1439
rect 3994 1387 4052 1405
rect 5418 1387 5476 1405
rect 6842 1387 6900 1405
rect 7723 1439 7781 1445
rect 8791 1439 8849 1445
rect 9859 1439 9917 1445
rect 7723 1405 7735 1439
rect 7735 1405 7769 1439
rect 7769 1405 7781 1439
rect 8791 1405 8803 1439
rect 8803 1405 8837 1439
rect 8837 1405 8849 1439
rect 9859 1405 9871 1439
rect 9871 1405 9905 1439
rect 9905 1405 9917 1439
rect 7723 1387 7781 1405
rect 8791 1387 8849 1405
rect 9859 1387 9917 1405
rect 10410 1439 10468 1445
rect 11478 1439 11536 1445
rect 12546 1439 12604 1445
rect 10410 1405 10422 1439
rect 10422 1405 10456 1439
rect 10456 1405 10468 1439
rect 11478 1405 11490 1439
rect 11490 1405 11524 1439
rect 11524 1405 11536 1439
rect 12546 1405 12558 1439
rect 12558 1405 12592 1439
rect 12592 1405 12604 1439
rect 10410 1387 10468 1405
rect 11478 1387 11536 1405
rect 12546 1387 12604 1405
rect 16738 2104 16796 2115
rect 16738 2070 16750 2104
rect 16750 2070 16784 2104
rect 16784 2070 16796 2104
rect 16738 2057 16796 2070
rect 17183 2052 17241 2110
rect 17539 2052 17597 2110
rect 18162 2104 18220 2110
rect 18162 2070 18174 2104
rect 18174 2070 18208 2104
rect 18208 2070 18220 2104
rect 18162 2052 18220 2070
rect 16560 1882 16618 1900
rect 16560 1848 16572 1882
rect 16572 1848 16606 1882
rect 16606 1848 16618 1882
rect 16560 1842 16618 1848
rect 16915 1882 16973 1901
rect 16915 1848 16928 1882
rect 16928 1848 16962 1882
rect 16962 1848 16973 1882
rect 16915 1843 16973 1848
rect 17806 1842 17864 1900
rect 17984 1882 18042 1900
rect 17984 1848 17996 1882
rect 17996 1848 18030 1882
rect 18030 1848 18042 1882
rect 17984 1842 18042 1848
rect 17183 1628 17241 1646
rect 17539 1628 17597 1646
rect 17183 1594 17186 1628
rect 17186 1594 17238 1628
rect 17238 1594 17241 1628
rect 17539 1594 17542 1628
rect 17542 1594 17594 1628
rect 17594 1594 17597 1628
rect 17183 1588 17241 1594
rect 17539 1588 17597 1594
rect 1484 1217 1542 1235
rect 2552 1217 2610 1235
rect 1484 1183 1496 1217
rect 1496 1183 1530 1217
rect 1530 1183 1542 1217
rect 2552 1183 2564 1217
rect 2564 1183 2598 1217
rect 2598 1183 2610 1217
rect 1484 1177 1542 1183
rect 2552 1177 2610 1183
rect 4884 1217 4942 1235
rect 5952 1217 6010 1235
rect 4884 1183 4896 1217
rect 4896 1183 4930 1217
rect 4930 1183 4942 1217
rect 5952 1183 5964 1217
rect 5964 1183 5998 1217
rect 5998 1183 6010 1217
rect 4884 1177 4942 1183
rect 5952 1177 6010 1183
rect 8257 1217 8315 1235
rect 9325 1217 9383 1235
rect 8257 1183 8269 1217
rect 8269 1183 8303 1217
rect 8303 1183 8315 1217
rect 9325 1183 9337 1217
rect 9337 1183 9371 1217
rect 9371 1183 9383 1217
rect 8257 1177 8315 1183
rect 9325 1177 9383 1183
rect 10944 1217 11002 1235
rect 12012 1217 12070 1235
rect 10944 1183 10956 1217
rect 10956 1183 10990 1217
rect 10990 1183 11002 1217
rect 12012 1183 12024 1217
rect 12024 1183 12058 1217
rect 12058 1183 12070 1217
rect 10944 1177 11002 1183
rect 12012 1177 12070 1183
rect 594 939 652 945
rect 2018 939 2076 945
rect 3442 939 3500 945
rect 594 905 606 939
rect 606 905 640 939
rect 640 905 652 939
rect 2018 905 2030 939
rect 2030 905 2064 939
rect 2064 905 2076 939
rect 3442 905 3454 939
rect 3454 905 3488 939
rect 3488 905 3500 939
rect 594 887 652 905
rect 2018 887 2076 905
rect 3442 887 3500 905
rect 3994 939 4052 945
rect 5418 939 5476 945
rect 6842 939 6900 945
rect 3994 905 4006 939
rect 4006 905 4040 939
rect 4040 905 4052 939
rect 5418 905 5430 939
rect 5430 905 5464 939
rect 5464 905 5476 939
rect 6842 905 6854 939
rect 6854 905 6888 939
rect 6888 905 6900 939
rect 3994 887 4052 905
rect 5418 887 5476 905
rect 6842 887 6900 905
rect 7723 939 7781 945
rect 8791 939 8849 945
rect 9859 939 9917 945
rect 7723 905 7735 939
rect 7735 905 7769 939
rect 7769 905 7781 939
rect 8791 905 8803 939
rect 8803 905 8837 939
rect 8837 905 8849 939
rect 9859 905 9871 939
rect 9871 905 9905 939
rect 9905 905 9917 939
rect 7723 887 7781 905
rect 8791 887 8849 905
rect 9859 887 9917 905
rect 10410 939 10468 945
rect 11478 939 11536 945
rect 12546 939 12604 945
rect 10410 905 10422 939
rect 10422 905 10456 939
rect 10456 905 10468 939
rect 11478 905 11490 939
rect 11490 905 11524 939
rect 11524 905 11536 939
rect 12546 905 12558 939
rect 12558 905 12592 939
rect 12592 905 12604 939
rect 10410 887 10468 905
rect 11478 887 11536 905
rect 12546 887 12604 905
rect 16738 1544 16796 1550
rect 16738 1510 16750 1544
rect 16750 1510 16784 1544
rect 16784 1510 16796 1544
rect 16738 1492 16796 1510
rect 16916 1492 16974 1550
rect 17806 1544 17864 1550
rect 17806 1510 17818 1544
rect 17818 1510 17852 1544
rect 17852 1510 17864 1544
rect 17806 1492 17864 1510
rect 18162 1544 18220 1550
rect 18162 1510 18174 1544
rect 18174 1510 18208 1544
rect 18208 1510 18220 1544
rect 18162 1492 18220 1510
rect 16560 1322 16618 1340
rect 17984 1322 18042 1340
rect 16560 1288 16572 1322
rect 16572 1288 16606 1322
rect 16606 1288 16618 1322
rect 17984 1288 17996 1322
rect 17996 1288 18030 1322
rect 18030 1288 18042 1322
rect 16560 1282 16618 1288
rect 17984 1282 18042 1288
rect 14134 788 14146 846
rect 14146 788 14180 846
rect 14180 788 14192 846
rect 14426 788 14438 846
rect 14438 788 14472 846
rect 14472 788 14484 846
rect 14718 788 14730 846
rect 14730 788 14764 846
rect 14764 788 14776 846
rect 15010 788 15022 846
rect 15022 788 15056 846
rect 15056 788 15068 846
rect 15302 788 15314 846
rect 15314 788 15348 846
rect 15348 788 15360 846
rect 16738 1044 16796 1050
rect 18162 1044 18220 1050
rect 16738 1010 16750 1044
rect 16750 1010 16784 1044
rect 16784 1010 16796 1044
rect 18162 1010 18174 1044
rect 18174 1010 18208 1044
rect 18208 1010 18220 1044
rect 16738 992 16796 1010
rect 18162 992 18220 1010
rect 16560 822 16618 840
rect 17984 822 18042 840
rect 16560 788 16572 822
rect 16572 788 16606 822
rect 16606 788 16618 822
rect 17984 788 17996 822
rect 17996 788 18030 822
rect 18030 788 18042 822
rect 16560 782 16618 788
rect 17984 782 18042 788
rect 1484 717 1542 735
rect 2552 717 2610 735
rect 1484 683 1496 717
rect 1496 683 1530 717
rect 1530 683 1542 717
rect 2552 683 2564 717
rect 2564 683 2598 717
rect 2598 683 2610 717
rect 1484 677 1542 683
rect 2552 677 2610 683
rect 4884 717 4942 735
rect 5952 717 6010 735
rect 4884 683 4896 717
rect 4896 683 4930 717
rect 4930 683 4942 717
rect 5952 683 5964 717
rect 5964 683 5998 717
rect 5998 683 6010 717
rect 4884 677 4942 683
rect 5952 677 6010 683
rect 8257 717 8315 735
rect 9325 717 9383 735
rect 8257 683 8269 717
rect 8269 683 8303 717
rect 8303 683 8315 717
rect 9325 683 9337 717
rect 9337 683 9371 717
rect 9371 683 9383 717
rect 8257 677 8315 683
rect 9325 677 9383 683
rect 10944 717 11002 735
rect 12012 717 12070 735
rect 10944 683 10956 717
rect 10956 683 10990 717
rect 10990 683 11002 717
rect 12012 683 12024 717
rect 12024 683 12058 717
rect 12058 683 12070 717
rect 17361 738 17419 739
rect 17361 704 17364 738
rect 17364 704 17416 738
rect 17416 704 17419 738
rect 10944 677 11002 683
rect 12012 677 12070 683
rect 17361 681 17419 704
rect 14109 516 14212 613
rect 15279 517 15382 614
rect 16547 524 16640 611
rect 17969 513 18062 600
rect 17361 322 17419 380
rect 19711 2530 19769 2536
rect 19711 2496 19723 2530
rect 19723 2496 19757 2530
rect 19757 2496 19769 2530
rect 19711 2478 19769 2496
rect 20066 2530 20124 2537
rect 20066 2496 20079 2530
rect 20079 2496 20113 2530
rect 20113 2496 20124 2530
rect 20066 2479 20124 2496
rect 20423 2530 20481 2536
rect 20423 2496 20435 2530
rect 20435 2496 20469 2530
rect 20469 2496 20481 2530
rect 20423 2478 20481 2496
rect 20779 2530 20837 2539
rect 20779 2496 20791 2530
rect 20791 2496 20825 2530
rect 20825 2496 20837 2530
rect 20779 2481 20837 2496
rect 21135 2530 21193 2536
rect 21135 2496 21147 2530
rect 21147 2496 21181 2530
rect 21181 2496 21193 2530
rect 21135 2478 21193 2496
rect 19533 2308 19591 2326
rect 20245 2308 20303 2321
rect 20957 2308 21015 2326
rect 19533 2274 19545 2308
rect 19545 2274 19579 2308
rect 19579 2274 19591 2308
rect 20245 2274 20257 2308
rect 20257 2274 20291 2308
rect 20291 2274 20303 2308
rect 20957 2274 20969 2308
rect 20969 2274 21003 2308
rect 21003 2274 21015 2308
rect 19533 2268 19591 2274
rect 20245 2263 20303 2274
rect 20957 2268 21015 2274
rect 19711 2032 19769 2038
rect 19711 1998 19723 2032
rect 19723 1998 19757 2032
rect 19757 1998 19769 2032
rect 19711 1980 19769 1998
rect 20066 2032 20124 2040
rect 20066 1998 20079 2032
rect 20079 1998 20113 2032
rect 20113 1998 20124 2032
rect 20066 1982 20124 1998
rect 20424 2032 20482 2041
rect 20424 1998 20435 2032
rect 20435 1998 20469 2032
rect 20469 1998 20482 2032
rect 20424 1983 20482 1998
rect 20779 2032 20837 2038
rect 20779 1998 20791 2032
rect 20791 1998 20825 2032
rect 20825 1998 20837 2032
rect 20779 1980 20837 1998
rect 21135 2032 21193 2038
rect 21135 1998 21147 2032
rect 21147 1998 21181 2032
rect 21181 1998 21193 2032
rect 21135 1980 21193 1998
rect 19533 1810 19591 1827
rect 20245 1810 20303 1827
rect 20957 1810 21015 1829
rect 19533 1776 19545 1810
rect 19545 1776 19579 1810
rect 19579 1776 19591 1810
rect 20245 1776 20257 1810
rect 20257 1776 20291 1810
rect 20291 1776 20303 1810
rect 20957 1776 20969 1810
rect 20969 1776 21003 1810
rect 21003 1776 21015 1810
rect 19533 1769 19591 1776
rect 20245 1769 20303 1776
rect 20957 1771 21015 1776
rect 19711 1504 19769 1510
rect 20423 1504 20481 1518
rect 21135 1504 21193 1510
rect 19711 1470 19723 1504
rect 19723 1470 19757 1504
rect 19757 1470 19769 1504
rect 20423 1470 20435 1504
rect 20435 1470 20469 1504
rect 20469 1470 20481 1504
rect 21135 1470 21147 1504
rect 21147 1470 21181 1504
rect 21181 1470 21193 1504
rect 19711 1452 19769 1470
rect 20423 1460 20481 1470
rect 21135 1452 21193 1470
rect 19533 1342 19591 1359
rect 20244 1342 20302 1359
rect 20957 1342 21015 1360
rect 19533 1308 19545 1342
rect 19545 1308 19579 1342
rect 19579 1308 19591 1342
rect 20244 1308 20257 1342
rect 20257 1308 20291 1342
rect 20291 1308 20302 1342
rect 20957 1308 20969 1342
rect 20969 1308 21003 1342
rect 21003 1308 21015 1342
rect 19533 1301 19591 1308
rect 20244 1301 20302 1308
rect 20957 1302 21015 1308
rect 19711 1006 19769 1012
rect 20423 1006 20481 1020
rect 21135 1006 21193 1012
rect 19711 972 19723 1006
rect 19723 972 19757 1006
rect 19757 972 19769 1006
rect 20423 972 20435 1006
rect 20435 972 20469 1006
rect 20469 972 20481 1006
rect 21135 972 21147 1006
rect 21147 972 21181 1006
rect 21181 972 21193 1006
rect 19711 954 19769 972
rect 20423 962 20481 972
rect 21135 954 21193 972
rect 19533 844 19591 862
rect 19533 810 19545 844
rect 19545 810 19579 844
rect 19579 810 19591 844
rect 19533 804 19591 810
rect 19889 844 19947 857
rect 19889 810 19901 844
rect 19901 810 19935 844
rect 19935 810 19947 844
rect 19889 799 19947 810
rect 20245 844 20303 855
rect 20245 810 20257 844
rect 20257 810 20291 844
rect 20291 810 20303 844
rect 20245 797 20303 810
rect 20601 844 20659 858
rect 20601 810 20613 844
rect 20613 810 20647 844
rect 20647 810 20659 844
rect 20601 800 20659 810
rect 20957 844 21015 862
rect 20957 810 20969 844
rect 20969 810 21003 844
rect 21003 810 21015 844
rect 20957 804 21015 810
rect 19533 628 19591 640
rect 19889 628 19947 639
rect 20245 628 20303 642
rect 20601 628 20659 640
rect 20957 628 21015 639
rect 19533 594 19591 628
rect 19889 594 19947 628
rect 20245 594 20303 628
rect 20601 594 20659 628
rect 20957 594 21015 628
rect 19533 582 19591 594
rect 19889 581 19947 594
rect 20245 584 20303 594
rect 20601 582 20659 594
rect 20957 581 21015 594
rect 1419 71 1609 134
rect 2500 71 2690 139
rect 4818 71 5008 141
rect 5891 71 6071 139
rect 8217 71 8355 141
rect 9273 71 9440 129
rect 10910 71 11036 139
rect 11978 71 12097 122
rect 1419 23 1609 71
rect 2500 28 2690 71
rect 4818 30 5008 71
rect 5891 23 6071 71
rect 8217 22 8355 71
rect 9273 22 9440 71
rect 10910 25 11036 71
rect 11978 25 12097 71
rect 14118 42 14211 129
rect 15279 36 15372 123
rect 16542 40 16635 127
rect 17969 35 18062 122
rect 8217 20 8355 22
rect 9273 13 9440 22
rect 21891 20 22019 148
<< metal2 >>
rect 21192 18864 21256 18865
rect 7286 18847 7350 18857
rect 8246 18847 8310 18857
rect 7284 18845 7286 18846
rect 7277 18793 7286 18845
rect 7284 18790 7286 18793
rect 7350 18845 7358 18846
rect 7350 18793 8246 18845
rect 7350 18790 7358 18793
rect 7286 18773 7350 18783
rect 20216 18851 20280 18861
rect 8310 18793 8313 18845
rect 8246 18773 8310 18783
rect 21180 18855 21256 18864
rect 21180 18854 21192 18855
rect 20280 18793 21180 18845
rect 20216 18777 20280 18787
rect 21256 18793 21272 18845
rect 21244 18790 21256 18791
rect 21180 18781 21256 18790
rect 21180 18780 21244 18781
rect 8229 18514 13131 18578
rect 8229 18354 8293 18514
rect 8229 18280 8293 18290
rect 7292 18041 7356 18051
rect 7277 17985 7292 18037
rect 7587 18037 7643 18046
rect 8247 18037 8311 18047
rect 7356 18036 8247 18037
rect 7356 17985 7587 18036
rect 7292 17967 7356 17977
rect 7643 17985 8247 18036
rect 7587 17970 7643 17980
rect 8247 17963 8311 17973
rect 13067 17415 13131 18514
rect 17762 18356 17826 18366
rect 17762 18282 17826 18292
rect 20867 18046 20931 18056
rect 20215 18038 20279 18045
rect 20215 18035 20867 18038
rect 20279 17986 20867 18035
rect 21182 18038 21246 18048
rect 20931 17986 21182 18038
rect 20867 17972 20931 17982
rect 21246 17986 21272 18038
rect 20215 17961 20279 17971
rect 21182 17964 21246 17974
rect 13067 17341 13131 17351
rect 12699 17135 12763 17145
rect 7287 17051 7351 17061
rect 8249 17054 8313 17064
rect 12699 17061 12763 17071
rect 7277 16993 7287 17045
rect 7351 16993 8249 17045
rect 7287 16977 7351 16987
rect 20219 17055 20283 17065
rect 8313 16993 8315 17045
rect 20204 16993 20219 17045
rect 8249 16980 8313 16990
rect 21179 17061 21243 17063
rect 21179 17053 21255 17061
rect 21243 17051 21255 17053
rect 20283 16993 21179 17045
rect 20219 16981 20283 16991
rect 21255 16993 21272 17045
rect 21179 16987 21191 16989
rect 21179 16979 21255 16987
rect 21191 16977 21255 16979
rect 8223 16554 8287 16564
rect 8223 16385 8287 16490
rect 10594 16552 10658 16562
rect 10594 16478 10658 16488
rect 17775 16554 17839 16564
rect 17775 16480 17839 16490
rect 14481 16440 14545 16450
rect 8223 16321 10938 16385
rect 7290 16240 7354 16250
rect 7277 16185 7290 16237
rect 7589 16237 7645 16247
rect 8248 16240 8312 16250
rect 7354 16185 7589 16237
rect 7290 16166 7354 16176
rect 7645 16185 8248 16237
rect 7589 16171 7645 16181
rect 8312 16185 8324 16237
rect 8248 16166 8312 16176
rect 10874 15829 10938 16321
rect 10874 15755 10938 15765
rect 12353 16271 12417 16281
rect 7286 15250 7350 15260
rect 7277 15193 7286 15245
rect 8247 15250 8311 15260
rect 7350 15193 8247 15245
rect 7286 15176 7350 15186
rect 8311 15193 8315 15245
rect 8247 15176 8311 15186
rect 12353 14878 12417 16207
rect 12701 16272 12765 16282
rect 12499 14878 12563 14888
rect 10637 14814 12499 14878
rect 8227 14754 8291 14764
rect 6815 14689 6910 14699
rect 613 14302 6815 14508
rect 613 3802 819 14302
rect 8227 14582 8291 14690
rect 10637 14753 10701 14814
rect 12499 14804 12563 14814
rect 10637 14679 10701 14689
rect 8227 14518 10702 14582
rect 6910 14302 6912 14508
rect 7288 14437 7352 14447
rect 7584 14438 7640 14448
rect 7277 14385 7288 14437
rect 7352 14385 7584 14437
rect 7288 14363 7352 14373
rect 8250 14440 8314 14450
rect 7640 14385 8250 14437
rect 7584 14372 7640 14382
rect 8314 14385 8319 14437
rect 8250 14366 8314 14376
rect 6815 14160 6910 14170
rect 10638 13986 10702 14518
rect 12701 14502 12765 16208
rect 14228 16217 14292 16227
rect 14228 16143 14292 16153
rect 14481 15828 14545 16376
rect 20218 16239 20282 16249
rect 20201 16186 20218 16238
rect 20863 16241 20927 16251
rect 20282 16186 20863 16238
rect 20218 16165 20282 16175
rect 21177 16238 21241 16248
rect 20927 16186 21177 16238
rect 20863 16167 20927 16177
rect 21241 16186 21272 16238
rect 21177 16164 21241 16174
rect 14481 15754 14545 15764
rect 15729 15765 15793 15775
rect 16489 15765 16553 15775
rect 14228 15743 14292 15753
rect 15793 15701 16489 15765
rect 15729 15691 15793 15701
rect 16489 15691 16553 15701
rect 14228 15669 14292 15679
rect 14839 15587 14903 15597
rect 14839 15513 14903 15523
rect 15155 15587 15219 15597
rect 16777 15587 16841 15597
rect 15219 15523 16777 15587
rect 15155 15513 15219 15523
rect 16777 15513 16841 15523
rect 17237 15591 17301 15601
rect 17237 15517 17301 15527
rect 20218 15253 20282 15263
rect 21191 15262 21255 15266
rect 14177 15222 14241 15232
rect 20215 15193 20218 15245
rect 21179 15256 21255 15262
rect 21179 15252 21191 15256
rect 20282 15193 21179 15245
rect 20218 15179 20282 15189
rect 21255 15193 21272 15245
rect 21243 15188 21255 15192
rect 21179 15182 21255 15188
rect 21179 15178 21243 15182
rect 14177 15148 14241 15158
rect 16278 15049 16342 15059
rect 16278 14975 16342 14985
rect 14379 14871 14443 14881
rect 14379 14797 14443 14807
rect 17830 14754 17894 14764
rect 17023 14690 17830 14754
rect 15947 14639 16011 14649
rect 16277 14639 16341 14649
rect 16011 14575 16277 14639
rect 15947 14565 16011 14575
rect 16277 14565 16341 14575
rect 14377 14521 14441 14531
rect 12701 14438 12937 14502
rect 11404 14142 11468 14152
rect 11404 14068 11468 14078
rect 11836 14142 11900 14152
rect 12479 14142 12543 14152
rect 11900 14078 12479 14142
rect 11836 14068 11900 14078
rect 12479 14068 12543 14078
rect 12702 14142 12766 14152
rect 12702 14068 12766 14078
rect 11404 13986 11468 13996
rect 10638 13966 11404 13986
rect 10637 13922 11404 13966
rect 11468 13922 11473 13986
rect 5457 13485 5869 13491
rect 7285 13448 7349 13458
rect 7277 13393 7285 13445
rect 7879 13446 7935 13456
rect 7349 13393 7879 13445
rect 7285 13374 7349 13384
rect 8252 13450 8316 13460
rect 7935 13393 8252 13445
rect 7879 13380 7935 13390
rect 8316 13393 8328 13445
rect 8252 13376 8316 13386
rect 10637 13195 10701 13922
rect 11404 13912 11468 13922
rect 11404 13813 11468 13823
rect 11404 13739 11468 13749
rect 11835 13812 11899 13822
rect 12873 13812 12937 14438
rect 11899 13748 12937 13812
rect 11835 13738 11899 13748
rect 14377 13282 14441 14457
rect 15945 14301 16009 14311
rect 15945 14227 16009 14237
rect 15581 14121 15645 14131
rect 17023 14121 17087 14690
rect 17830 14680 17894 14690
rect 20217 14438 20281 14447
rect 20864 14442 20928 14452
rect 20217 14437 20864 14438
rect 20281 14386 20864 14437
rect 20217 14363 20281 14373
rect 21180 14442 21244 14452
rect 20928 14386 21180 14438
rect 20864 14368 20928 14378
rect 21244 14386 21272 14438
rect 21180 14368 21244 14378
rect 15645 14057 17087 14121
rect 15581 14047 15645 14057
rect 15579 13810 15643 13820
rect 15643 13746 17082 13810
rect 15579 13736 15643 13746
rect 14377 13208 14441 13218
rect 5457 10415 5869 13073
rect 8224 13131 10701 13195
rect 8224 12954 8288 13131
rect 8224 12880 8288 12890
rect 10637 12950 10701 12960
rect 17018 12956 17082 13746
rect 20218 13450 20282 13460
rect 20215 13393 20218 13445
rect 20575 13451 20639 13461
rect 20282 13393 20575 13445
rect 20218 13376 20282 13386
rect 21178 13450 21242 13460
rect 20639 13393 21178 13445
rect 20575 13377 20639 13387
rect 21242 13393 21272 13445
rect 21178 13376 21242 13386
rect 17835 12956 17899 12966
rect 17018 12892 17835 12956
rect 7287 12640 7351 12650
rect 7277 12585 7287 12637
rect 8180 12642 8317 12652
rect 8180 12638 8253 12642
rect 8180 12637 8187 12638
rect 7351 12585 8187 12637
rect 7287 12566 7351 12576
rect 8180 12582 8187 12585
rect 8243 12582 8253 12638
rect 8180 12578 8253 12582
rect 8317 12585 8346 12637
rect 8180 12568 8317 12578
rect 10637 12333 10701 12886
rect 14379 12882 14443 12892
rect 17835 12882 17899 12892
rect 14379 12808 14443 12818
rect 20264 12646 20328 12651
rect 20215 12641 20328 12646
rect 20215 12638 20264 12641
rect 20204 12636 20264 12638
rect 21180 12638 21244 12648
rect 20204 12586 20215 12636
rect 20328 12586 21180 12638
rect 20279 12572 20328 12577
rect 20215 12567 20328 12572
rect 21244 12586 21272 12638
rect 20215 12562 20279 12567
rect 21180 12564 21244 12574
rect 15508 12363 15572 12373
rect 16497 12363 16561 12373
rect 11611 12333 11675 12343
rect 12901 12333 12965 12343
rect 10637 12269 11611 12333
rect 11675 12269 12901 12333
rect 11611 12259 11675 12269
rect 12901 12259 12965 12269
rect 13401 12299 13465 12309
rect 15572 12299 16497 12363
rect 15508 12289 15572 12299
rect 16497 12289 16561 12299
rect 13401 12225 13465 12235
rect 14673 12185 14737 12195
rect 14673 12111 14737 12121
rect 14965 12181 15029 12191
rect 16807 12181 16871 12191
rect 15029 12117 16807 12181
rect 14965 12107 15029 12117
rect 16807 12107 16871 12117
rect 17223 12185 17287 12195
rect 17223 12111 17287 12121
rect 11241 12000 11305 12010
rect 11241 11926 11305 11936
rect 12001 12000 12065 12010
rect 15014 12000 15078 12010
rect 12065 11936 15014 12000
rect 12001 11926 12065 11936
rect 15014 11926 15078 11936
rect 15397 12000 15461 12010
rect 15397 11926 15461 11936
rect 21885 11732 21996 11742
rect 6335 11649 6747 11670
rect 6331 11637 6747 11649
rect 7287 11651 7351 11661
rect 6331 11514 6348 11637
rect 6458 11514 6747 11637
rect 7277 11593 7287 11645
rect 7878 11647 7934 11657
rect 7351 11593 7878 11645
rect 7287 11577 7351 11587
rect 8250 11651 8314 11661
rect 7934 11593 8250 11645
rect 7878 11581 7934 11591
rect 20217 11649 20281 11659
rect 8314 11593 8316 11645
rect 20215 11593 20217 11645
rect 8250 11577 8314 11587
rect 20574 11652 20638 11662
rect 20281 11593 20574 11645
rect 20217 11575 20281 11585
rect 21182 11650 21246 11660
rect 20638 11593 21182 11645
rect 20574 11578 20638 11588
rect 21246 11593 21272 11645
rect 21182 11576 21246 11586
rect 23475 11592 23656 11602
rect 6331 11443 6335 11514
rect 6334 11102 6335 11105
rect 21881 11429 21885 11539
rect 21997 11429 23475 11539
rect 23475 11363 23656 11373
rect 21885 11215 21996 11225
rect 6334 11097 6348 11102
rect 6458 11097 6747 11102
rect 6334 10899 6747 11097
rect 8231 11156 8295 11166
rect 8231 11007 8295 11092
rect 17771 11152 17835 11162
rect 17771 11078 17835 11088
rect 12494 11008 12558 11018
rect 8231 10944 12494 11007
rect 8231 10943 12558 10944
rect 12494 10934 12558 10943
rect 3439 5643 3448 5735
rect 3540 5643 3549 5735
rect 3448 4676 3540 5643
rect 4166 5350 4258 5365
rect 3448 4564 3541 4676
rect 2829 4321 2887 4331
rect 2256 4049 2522 4059
rect 2256 3985 2522 3995
rect 613 3692 657 3802
rect 767 3692 819 3802
rect 613 3682 819 3692
rect 2338 3455 2430 3985
rect 2829 3961 2887 4263
rect 3448 4237 3540 4564
rect 4166 4238 4258 5258
rect 5457 4656 5870 10415
rect 4609 4321 4667 4331
rect 3404 4227 3569 4237
rect 3404 4163 3569 4173
rect 4128 4228 4293 4238
rect 4128 4164 4293 4174
rect 2829 3892 2887 3903
rect 4609 3961 4667 4263
rect 5457 4254 5462 4656
rect 5864 4455 5870 4656
rect 5457 4249 5664 4254
rect 5462 4245 5870 4249
rect 5664 4210 5870 4245
rect 4884 4051 5150 4061
rect 4884 3987 5150 3997
rect 4609 3895 4667 3903
rect 4961 3458 5053 3987
rect 6335 3586 6747 10899
rect 8195 10849 8320 10852
rect 7287 10837 7351 10847
rect 8192 10841 8320 10849
rect 8192 10839 8250 10841
rect 7277 10785 7287 10837
rect 7351 10785 8192 10837
rect 8248 10783 8250 10839
rect 8192 10777 8250 10783
rect 8314 10777 8320 10841
rect 8192 10773 8320 10777
rect 7287 10763 7351 10773
rect 8195 10765 8320 10773
rect 20217 10844 20281 10848
rect 20217 10838 20333 10844
rect 21179 10839 21243 10849
rect 20281 10834 21179 10838
rect 20333 10786 21179 10834
rect 20217 10770 20269 10774
rect 20217 10764 20333 10770
rect 21243 10786 21272 10838
rect 21179 10765 21243 10775
rect 20269 10760 20333 10764
rect 11231 10441 11295 10451
rect 7287 9851 7351 9861
rect 7277 9793 7287 9845
rect 7871 9858 7935 9868
rect 7351 9794 7871 9845
rect 8248 9852 8312 9862
rect 7935 9794 8248 9845
rect 7351 9793 8248 9794
rect 7287 9777 7351 9787
rect 7871 9784 7935 9793
rect 8312 9793 8318 9845
rect 8248 9778 8312 9788
rect 10707 9585 10771 9595
rect 8232 9521 10707 9585
rect 8232 9355 8296 9521
rect 10707 9511 10771 9521
rect 8232 9281 8296 9291
rect 10569 9358 10633 9368
rect 11231 9358 11295 10377
rect 20219 9850 20283 9860
rect 20216 9793 20219 9845
rect 20574 9848 20638 9858
rect 20283 9793 20574 9845
rect 20219 9776 20283 9786
rect 21179 9850 21243 9860
rect 20638 9793 21179 9845
rect 20574 9774 20638 9784
rect 21243 9793 21272 9845
rect 22387 9835 22593 9877
rect 21179 9776 21243 9786
rect 10633 9294 11295 9358
rect 17789 9360 17853 9370
rect 10569 9284 10633 9294
rect 17789 9286 17853 9296
rect 22387 9295 22399 9835
rect 22509 9295 22593 9835
rect 7290 9037 7354 9047
rect 8186 9039 8311 9049
rect 7277 8985 7290 9037
rect 7354 8985 8186 9037
rect 7290 8963 7354 8973
rect 20216 9047 20280 9050
rect 20216 9040 20332 9047
rect 20280 9038 20332 9040
rect 21181 9039 21245 9049
rect 20280 9037 21181 9038
rect 8311 8985 8312 9037
rect 8186 8965 8311 8975
rect 20332 8986 21181 9037
rect 20216 8973 20268 8976
rect 20216 8966 20332 8973
rect 20268 8963 20332 8966
rect 21245 8986 21272 9038
rect 21181 8965 21245 8975
rect 8256 7002 8314 7012
rect 8078 6598 8136 6608
rect 8078 6025 8136 6540
rect 8078 5957 8136 5967
rect 8256 6393 8314 6944
rect 8256 5815 8314 6335
rect 9324 7005 9382 7015
rect 9324 6393 9382 6947
rect 10942 7002 11000 7012
rect 8722 6032 8914 6042
rect 8722 5967 8790 5974
rect 8848 5967 8914 5974
rect 8722 5964 8914 5967
rect 8256 5747 8314 5757
rect 8765 5730 8875 5964
rect 9324 5815 9382 6335
rect 9502 6603 9560 6613
rect 9502 6025 9560 6545
rect 10764 6597 10822 6607
rect 9768 6209 9826 6219
rect 10497 6209 10555 6219
rect 9826 6151 10497 6209
rect 9768 6141 9826 6151
rect 10497 6141 10555 6151
rect 9502 5957 9560 5967
rect 10764 6026 10822 6539
rect 10764 5958 10822 5968
rect 10942 6393 11000 6944
rect 9324 5747 9382 5757
rect 10942 5816 11000 6335
rect 12010 7007 12068 7017
rect 12010 6393 12068 6949
rect 14862 6666 14920 6676
rect 15218 6666 15276 6676
rect 15574 6666 15632 6676
rect 15930 6666 15988 6676
rect 17063 6666 17121 6676
rect 17418 6666 17476 6676
rect 17774 6666 17832 6676
rect 18130 6666 18188 6676
rect 19262 6666 19320 6676
rect 19618 6666 19676 6676
rect 19974 6666 20032 6676
rect 20330 6666 20388 6676
rect 11408 6030 11600 6040
rect 11408 5968 11476 5972
rect 11534 5968 11600 5972
rect 11408 5962 11600 5968
rect 10942 5748 11000 5758
rect 8765 5648 8789 5730
rect 8871 5648 8875 5730
rect 8078 5145 8136 5155
rect 8078 4575 8136 5087
rect 8078 4507 8136 4517
rect 8256 4935 8314 4945
rect 8765 4941 8875 5648
rect 11445 5345 11555 5962
rect 12010 5816 12068 6335
rect 12188 6604 12246 6614
rect 14920 6608 15218 6666
rect 15276 6608 15574 6666
rect 15632 6608 15930 6666
rect 15988 6608 16109 6666
rect 14862 6598 14920 6608
rect 15218 6598 15276 6608
rect 15574 6598 15632 6608
rect 15930 6598 15988 6608
rect 12188 6026 12246 6546
rect 15040 6468 15098 6478
rect 15396 6468 15454 6478
rect 15752 6468 15810 6478
rect 15098 6410 15396 6468
rect 15454 6410 15752 6468
rect 15040 6400 15098 6410
rect 15396 6400 15454 6410
rect 15752 6400 15810 6410
rect 12446 6280 12525 6290
rect 12844 6228 12957 6238
rect 12525 6111 12844 6228
rect 12844 6101 12957 6111
rect 12446 6070 12525 6080
rect 12188 5958 12246 5968
rect 12010 5748 12068 5758
rect 14863 5899 14921 5909
rect 15219 5899 15277 5909
rect 15575 5899 15633 5909
rect 15931 5899 15989 5909
rect 14921 5841 15219 5899
rect 15277 5841 15575 5899
rect 15633 5841 15931 5899
rect 14863 5450 14921 5841
rect 15219 5831 15277 5841
rect 15575 5831 15633 5841
rect 15931 5831 15989 5841
rect 15041 5701 15099 5711
rect 15397 5701 15455 5711
rect 15752 5701 15810 5711
rect 16051 5701 16109 6608
rect 15099 5643 15397 5701
rect 15455 5643 15752 5701
rect 15810 5643 16109 5701
rect 16893 6608 17063 6666
rect 17121 6608 17418 6666
rect 17476 6608 17774 6666
rect 17832 6608 18130 6666
rect 18188 6608 18189 6666
rect 16893 6568 18189 6608
rect 19074 6608 19262 6666
rect 19320 6608 19618 6666
rect 19676 6608 19974 6666
rect 20032 6608 20330 6666
rect 19074 6568 20388 6608
rect 16893 5738 17000 6568
rect 17240 6468 17298 6478
rect 17596 6468 17654 6477
rect 17952 6468 18010 6478
rect 17298 6467 17952 6468
rect 17298 6410 17596 6467
rect 17240 6400 17298 6410
rect 17654 6410 17952 6467
rect 17596 6399 17654 6409
rect 17952 6400 18010 6410
rect 17064 5909 18248 5930
rect 17063 5899 18248 5909
rect 17121 5841 17419 5899
rect 17477 5841 17775 5899
rect 17833 5841 18131 5899
rect 18189 5841 18248 5899
rect 17063 5832 18248 5841
rect 17063 5831 17121 5832
rect 17419 5831 17477 5832
rect 17775 5831 17833 5832
rect 16893 5701 18022 5738
rect 16893 5643 17242 5701
rect 17300 5643 17597 5701
rect 17655 5643 17953 5701
rect 18011 5643 18022 5701
rect 15041 5633 15099 5643
rect 15397 5633 15455 5643
rect 15752 5633 15810 5643
rect 16893 5640 18022 5643
rect 17242 5633 17300 5640
rect 17597 5633 17655 5640
rect 17953 5633 18011 5640
rect 14863 5382 14921 5392
rect 11445 5263 11473 5345
rect 9858 5145 9916 5155
rect 8256 4365 8314 4877
rect 8725 4935 8917 4941
rect 8725 4931 8790 4935
rect 8848 4931 8917 4935
rect 8725 4863 8917 4873
rect 9680 4935 9738 4945
rect 9680 4681 9738 4877
rect 8725 4577 8917 4587
rect 9660 4569 9752 4681
rect 9858 4575 9916 5087
rect 8725 4517 8790 4519
rect 8848 4517 8917 4519
rect 8725 4509 8917 4517
rect 8763 4464 8873 4509
rect 8256 4297 8314 4307
rect 8757 4454 8881 4464
rect 9680 4365 9738 4569
rect 9858 4507 9916 4517
rect 10408 5145 10466 5155
rect 10408 4575 10466 5087
rect 10408 4507 10466 4517
rect 10586 4935 10644 4945
rect 11445 4942 11555 5263
rect 12188 5145 12246 5155
rect 10586 4455 10644 4877
rect 11404 4935 11596 4942
rect 11404 4932 11476 4935
rect 11534 4932 11596 4935
rect 11404 4864 11596 4874
rect 12010 4935 12068 4945
rect 11406 4576 11598 4586
rect 11406 4517 11478 4518
rect 11536 4517 11598 4518
rect 11406 4508 11598 4517
rect 10570 4365 10662 4455
rect 10570 4343 10586 4365
rect 9680 4297 9738 4307
rect 10644 4343 10662 4365
rect 10586 4297 10644 4307
rect 8757 4239 8881 4249
rect 8763 3655 8873 4239
rect 11450 3656 11560 4508
rect 12010 4365 12068 4877
rect 12188 4575 12246 5087
rect 13894 5053 13952 5063
rect 12188 4507 12246 4517
rect 13716 4843 13774 4853
rect 12010 4297 12068 4307
rect 13716 4343 13774 4785
rect 13894 4553 13952 4995
rect 16030 5053 16088 5063
rect 13894 4485 13952 4495
rect 15852 4843 15910 4853
rect 13716 4275 13774 4285
rect 15852 4343 15910 4785
rect 16030 4553 16088 4995
rect 18131 5057 18248 5832
rect 19074 5731 19200 6568
rect 19440 6468 19498 6478
rect 19796 6468 19854 6478
rect 20152 6468 20210 6478
rect 19498 6410 19796 6468
rect 19854 6410 20152 6468
rect 19440 6400 19498 6410
rect 19796 6400 19854 6410
rect 20152 6400 20210 6410
rect 20241 6357 20299 6367
rect 19264 5899 19322 5909
rect 19619 5899 19677 5909
rect 19975 5899 20033 5909
rect 20241 5899 20299 6299
rect 20331 5899 20462 5909
rect 19322 5841 19619 5899
rect 19677 5841 19975 5899
rect 20033 5841 20331 5899
rect 19264 5831 19322 5841
rect 19619 5831 19677 5841
rect 19975 5831 20033 5841
rect 19074 5701 20211 5731
rect 19074 5643 19442 5701
rect 19500 5643 19797 5701
rect 19855 5643 20153 5701
rect 19074 5633 20211 5643
rect 19353 5590 19411 5600
rect 16030 4485 16088 4495
rect 17988 4843 18046 4853
rect 15852 4275 15910 4285
rect 17630 4387 17752 4397
rect 17688 4285 17752 4286
rect 17452 4241 17510 4251
rect 7723 3645 7781 3655
rect 594 3445 652 3455
rect 594 2945 652 3387
rect 2018 3445 2076 3455
rect 594 2445 652 2887
rect 594 1945 652 2387
rect 594 1445 652 1887
rect 594 945 652 1387
rect 594 877 652 887
rect 1484 3235 1542 3245
rect 1484 2735 1542 3177
rect 1484 2235 1542 2677
rect 1484 1735 1542 2177
rect 1484 1235 1542 1677
rect 1484 735 1542 1177
rect 2018 2945 2076 3387
rect 2256 3445 2522 3455
rect 2256 3381 2522 3391
rect 3442 3445 3500 3455
rect 2018 2445 2076 2887
rect 2018 1945 2076 2387
rect 2018 1445 2076 1887
rect 2018 945 2076 1387
rect 2018 877 2076 887
rect 2552 3235 2610 3245
rect 2552 2735 2610 3177
rect 2552 2235 2610 2677
rect 2552 1735 2610 2177
rect 2552 1235 2610 1677
rect 1484 144 1542 677
rect 2552 735 2610 1177
rect 3442 2945 3500 3387
rect 3442 2445 3500 2887
rect 3442 1945 3500 2387
rect 3442 1445 3500 1887
rect 3442 945 3500 1387
rect 3442 877 3500 887
rect 3994 3445 4052 3455
rect 3994 2945 4052 3387
rect 4886 3448 5152 3458
rect 4886 3384 5152 3394
rect 5418 3445 5476 3455
rect 3994 2445 4052 2887
rect 3994 1945 4052 2387
rect 3994 1445 4052 1887
rect 3994 945 4052 1387
rect 3994 877 4052 887
rect 4884 3235 4942 3245
rect 4884 2735 4942 3177
rect 4884 2235 4942 2677
rect 4884 1735 4942 2177
rect 4884 1235 4942 1677
rect 2552 149 2610 677
rect 4884 735 4942 1177
rect 5418 2945 5476 3387
rect 5418 2445 5476 2887
rect 5418 1945 5476 2387
rect 5418 1445 5476 1887
rect 5418 945 5476 1387
rect 5418 877 5476 887
rect 5952 3235 6010 3245
rect 6331 3184 6340 3586
rect 6742 3184 6751 3586
rect 6842 3445 6900 3455
rect 6335 3179 6747 3184
rect 5952 2736 6010 3177
rect 5952 2235 6010 2678
rect 5952 1735 6010 2177
rect 5952 1235 6010 1677
rect 4884 151 4942 677
rect 5952 735 6010 1177
rect 6842 2945 6900 3387
rect 6842 2445 6900 2887
rect 7723 3145 7781 3587
rect 8718 3645 8910 3655
rect 8718 3577 8910 3587
rect 9859 3645 9917 3655
rect 8790 3536 8849 3577
rect 7723 2645 7781 3087
rect 7723 2577 7781 2587
rect 8257 3435 8315 3445
rect 8257 2935 8315 3377
rect 6842 1945 6900 2387
rect 8257 2435 8315 2877
rect 8791 3145 8849 3536
rect 8791 2645 8849 3087
rect 8791 2577 8849 2587
rect 9325 3435 9383 3445
rect 9325 2935 9383 3377
rect 8257 2367 8315 2377
rect 8609 2426 8800 2436
rect 8609 2363 8800 2373
rect 9325 2435 9383 2877
rect 9859 3145 9917 3587
rect 9859 2645 9917 3087
rect 9859 2577 9917 2587
rect 10410 3645 10468 3655
rect 10410 3145 10468 3587
rect 11414 3646 11606 3656
rect 11414 3578 11452 3588
rect 10410 2645 10468 3087
rect 10410 2577 10468 2587
rect 10944 3435 11002 3445
rect 10944 2935 11002 3377
rect 11558 3578 11606 3588
rect 12546 3645 12604 3655
rect 12012 3435 12070 3445
rect 11558 3379 11561 3388
rect 11558 3270 11561 3279
rect 11452 3172 11558 3182
rect 9325 2367 9383 2377
rect 10944 2435 11002 2877
rect 11478 3145 11536 3172
rect 11478 2645 11536 3087
rect 11478 2577 11536 2587
rect 12012 2935 12070 3377
rect 11591 2436 11701 2439
rect 10944 2367 11002 2377
rect 11546 2426 11752 2436
rect 8670 1956 8780 2363
rect 11546 2358 11752 2368
rect 12012 2435 12070 2877
rect 12546 3145 12604 3587
rect 17452 3651 17510 4183
rect 17452 3583 17510 3593
rect 17630 4125 17752 4285
rect 17988 4343 18046 4785
rect 18131 4563 18248 4940
rect 19175 5106 19233 5116
rect 19175 4735 19233 4986
rect 19353 4834 19411 5532
rect 20331 5151 20462 5841
rect 20331 5141 20477 5151
rect 19175 4725 19234 4735
rect 18131 4553 18249 4563
rect 18131 4444 18132 4553
rect 18132 4426 18249 4436
rect 19175 4546 19176 4725
rect 19233 4507 19234 4517
rect 17988 4275 18046 4285
rect 17630 3550 17752 4007
rect 17630 3549 17631 3550
rect 17274 3530 17332 3540
rect 17272 3278 17274 3334
rect 17630 3481 17631 3491
rect 19175 4224 19233 4488
rect 19175 3736 19233 3990
rect 19175 3482 19233 3492
rect 19353 4336 19411 4776
rect 19353 3838 19411 4278
rect 17272 3268 17332 3278
rect 17433 3416 17535 3426
rect 17631 3423 17752 3433
rect 17433 3279 17452 3416
rect 17510 3279 17535 3416
rect 12546 2645 12604 3087
rect 14863 3097 14921 3107
rect 14863 3029 14921 3039
rect 17272 2712 17330 3268
rect 17433 3017 17535 3279
rect 19353 3340 19411 3780
rect 19709 5110 19767 5120
rect 19709 4729 19767 5021
rect 21132 5115 21190 5125
rect 20477 5001 20478 5113
rect 21190 5026 21191 5109
rect 21132 5016 21191 5026
rect 20331 4991 20478 5001
rect 20066 4841 20124 4843
rect 20065 4831 20124 4841
rect 20123 4773 20124 4831
rect 20065 4763 20124 4773
rect 19709 4719 19768 4729
rect 19709 4511 19710 4719
rect 19709 4501 19768 4511
rect 19709 4223 19767 4501
rect 20066 4341 20124 4763
rect 20065 4331 20124 4341
rect 20123 4273 20124 4331
rect 20065 4263 20124 4273
rect 19709 3736 19767 4015
rect 20066 3847 20124 4263
rect 20065 3837 20124 3847
rect 20123 3779 20124 3837
rect 20065 3769 20124 3779
rect 19708 3726 19767 3736
rect 19766 3680 19767 3726
rect 19708 3508 19766 3518
rect 19353 3272 19411 3282
rect 19710 3339 19768 3349
rect 20066 3339 20124 3769
rect 20420 4730 20478 4991
rect 20420 4233 20478 4522
rect 20779 4835 20837 4845
rect 20779 4344 20837 4777
rect 20778 4334 20837 4344
rect 20836 4276 20837 4334
rect 20778 4266 20837 4276
rect 20420 4223 20480 4233
rect 20420 4015 20422 4223
rect 20420 4005 20480 4015
rect 20420 3723 20478 4005
rect 20779 3851 20837 4266
rect 20774 3841 20837 3851
rect 20832 3783 20837 3841
rect 20774 3773 20837 3783
rect 20420 3505 20478 3515
rect 19768 3281 19769 3335
rect 19710 3271 19769 3281
rect 17432 3008 17542 3017
rect 17432 3007 17433 3008
rect 17535 3007 17542 3008
rect 17432 2887 17433 2897
rect 12546 2577 12604 2587
rect 16738 2608 16796 2618
rect 14134 2538 14192 2548
rect 14426 2538 14484 2548
rect 14718 2538 14776 2548
rect 15010 2538 15068 2548
rect 15302 2538 15360 2548
rect 14192 2480 14426 2538
rect 14484 2480 14718 2538
rect 14776 2480 15010 2538
rect 15068 2480 15302 2538
rect 14134 2470 14192 2480
rect 14426 2470 14484 2480
rect 14718 2470 14776 2480
rect 15010 2470 15068 2480
rect 15302 2470 15360 2480
rect 12012 2367 12070 2377
rect 16560 2400 16618 2410
rect 11591 1956 11701 2358
rect 6842 1445 6900 1887
rect 6842 945 6900 1387
rect 6842 877 6900 887
rect 7723 1945 7781 1955
rect 7723 1445 7781 1887
rect 8593 1946 8857 1956
rect 11500 1955 11708 1956
rect 8593 1877 8857 1887
rect 9859 1945 9917 1955
rect 7723 945 7781 1387
rect 7723 877 7781 887
rect 8257 1735 8315 1745
rect 8257 1235 8315 1677
rect 1419 134 1609 144
rect 1419 13 1609 23
rect 2500 139 2690 149
rect 2500 18 2690 28
rect 4818 141 5008 151
rect 5952 149 6010 677
rect 8257 735 8315 1177
rect 8791 1445 8849 1877
rect 8791 945 8849 1387
rect 8791 877 8849 887
rect 9325 1735 9383 1745
rect 9325 1235 9383 1677
rect 8257 151 8315 677
rect 9325 735 9383 1177
rect 9859 1445 9917 1887
rect 9859 945 9917 1387
rect 9859 877 9917 887
rect 10410 1945 10468 1955
rect 10410 1445 10468 1887
rect 11478 1946 11708 1955
rect 11478 1945 11502 1946
rect 11478 1886 11502 1887
rect 11478 1876 11708 1886
rect 12546 1945 12604 1955
rect 10410 945 10468 1387
rect 10410 877 10468 887
rect 10944 1735 11002 1745
rect 10944 1235 11002 1677
rect 4818 20 5008 30
rect 5891 139 6071 149
rect 5891 13 6071 23
rect 8217 141 8355 151
rect 9325 139 9383 677
rect 10944 735 11002 1177
rect 11478 1445 11536 1876
rect 11478 945 11536 1387
rect 11478 877 11536 887
rect 12012 1735 12070 1745
rect 12012 1235 12070 1677
rect 10944 149 11002 677
rect 12012 735 12070 1177
rect 12546 1445 12604 1887
rect 16560 1900 16618 2342
rect 16738 2115 16796 2550
rect 17272 2293 17330 2654
rect 17535 2887 17542 2897
rect 17433 2620 17535 2803
rect 17420 2610 17535 2620
rect 17420 2504 17535 2514
rect 18162 2610 18220 2620
rect 17984 2400 18042 2410
rect 17243 2283 17361 2293
rect 17243 2156 17361 2166
rect 16738 2047 16796 2057
rect 17183 2110 17241 2120
rect 16560 1832 16618 1842
rect 16915 1901 16973 1911
rect 16973 1843 16974 1880
rect 16915 1833 16974 1843
rect 12546 945 12604 1387
rect 16738 1550 16796 1560
rect 12546 877 12604 887
rect 16560 1340 16618 1350
rect 14134 846 14192 856
rect 14426 846 14484 856
rect 14718 846 14776 856
rect 15010 846 15068 856
rect 15302 846 15360 856
rect 10910 139 11036 149
rect 8217 10 8355 20
rect 9273 129 9440 139
rect 12012 132 12070 677
rect 14133 788 14134 801
rect 14192 788 14426 846
rect 14484 788 14718 846
rect 14776 788 15010 846
rect 15068 788 15302 846
rect 14133 778 14192 788
rect 14426 778 14484 788
rect 14718 778 14776 788
rect 15010 778 15068 788
rect 14133 623 14191 778
rect 15302 624 15360 788
rect 16560 840 16618 1282
rect 16738 1050 16796 1492
rect 16916 1550 16974 1833
rect 17183 1646 17241 2052
rect 17183 1578 17241 1588
rect 17539 2110 17597 2120
rect 17539 1646 17597 2052
rect 17539 1578 17597 1588
rect 17806 1900 17864 1910
rect 16916 1482 16974 1492
rect 17806 1550 17864 1842
rect 17984 1900 18042 2342
rect 18162 2110 18220 2552
rect 19711 2536 19769 3271
rect 18162 2042 18220 2052
rect 19533 2326 19591 2336
rect 17984 1832 18042 1842
rect 19533 1827 19591 2268
rect 19711 2038 19769 2478
rect 19711 1970 19769 1980
rect 20066 2537 20124 3281
rect 20066 2040 20124 2479
rect 20423 3340 20481 3350
rect 20423 2536 20481 3282
rect 20066 1972 20124 1982
rect 20245 2321 20303 2331
rect 17806 1482 17864 1492
rect 18162 1550 18220 1560
rect 16738 982 16796 992
rect 17984 1340 18042 1350
rect 14109 613 14212 623
rect 14109 506 14212 516
rect 15279 614 15382 624
rect 16560 621 16618 782
rect 17984 840 18042 1282
rect 18162 1050 18220 1492
rect 18162 982 18220 992
rect 19533 1359 19591 1769
rect 20245 1827 20303 2263
rect 20423 2051 20481 2478
rect 20779 3337 20837 3773
rect 21133 4723 21191 5016
rect 21667 5106 21725 5116
rect 21133 4230 21191 4515
rect 21133 3721 21191 4022
rect 21133 3503 21191 3513
rect 21489 4834 21547 4844
rect 21489 4336 21547 4776
rect 21489 3838 21547 4278
rect 21667 4716 21725 4986
rect 21667 4228 21725 4488
rect 21666 4218 21725 4228
rect 21724 4048 21725 4218
rect 21666 4000 21667 4010
rect 20779 2539 20837 3279
rect 20423 2041 20482 2051
rect 20423 1983 20424 2041
rect 20423 1973 20482 1983
rect 20779 2038 20837 2481
rect 21135 3338 21193 3348
rect 21135 2536 21193 3280
rect 21489 3340 21547 3780
rect 21667 3736 21725 3990
rect 21667 3482 21725 3492
rect 21489 3272 21547 3282
rect 21880 3180 22031 3192
rect 21880 3052 21891 3180
rect 22019 3052 22031 3180
rect 21880 3042 22031 3052
rect 20779 1970 20837 1980
rect 20957 2326 21015 2336
rect 17361 739 17419 749
rect 15279 507 15382 517
rect 16547 611 16640 621
rect 16547 514 16640 524
rect 14133 139 14191 506
rect 10910 15 11036 25
rect 11978 122 12097 132
rect 14118 129 14211 139
rect 15302 133 15360 507
rect 16560 137 16618 514
rect 17361 380 17419 681
rect 17984 610 18042 782
rect 19533 862 19591 1301
rect 19711 1510 19769 1520
rect 19711 1012 19769 1452
rect 20245 1369 20303 1769
rect 20957 1829 21015 2268
rect 21135 2038 21193 2478
rect 21135 1970 21193 1980
rect 20244 1359 20303 1369
rect 20302 1301 20303 1359
rect 20244 1291 20303 1301
rect 19711 944 19769 954
rect 19533 640 19591 804
rect 17969 600 18062 610
rect 19533 572 19591 582
rect 19889 857 19947 867
rect 19889 639 19947 799
rect 19889 571 19947 581
rect 20245 855 20303 1291
rect 20423 1518 20481 1528
rect 20423 1020 20481 1460
rect 20423 952 20481 962
rect 20957 1360 21015 1771
rect 20245 642 20303 797
rect 20245 574 20303 584
rect 20601 858 20659 868
rect 20601 640 20659 800
rect 20601 572 20659 582
rect 20957 862 21015 1302
rect 21135 1510 21193 1520
rect 21135 1012 21193 1452
rect 21135 944 21193 954
rect 20957 639 21015 804
rect 20957 571 21015 581
rect 17969 503 18062 513
rect 17361 312 17419 322
rect 14118 32 14211 42
rect 15279 123 15372 133
rect 15279 26 15372 36
rect 16542 127 16635 137
rect 17984 132 18042 503
rect 21891 148 22019 3042
rect 22387 3004 22593 9295
rect 22387 2788 22593 2798
rect 16542 30 16635 40
rect 17969 122 18062 132
rect 17969 25 18062 35
rect 11978 15 12097 25
rect 21891 14 22019 20
rect 9273 3 9440 13
<< via2 >>
rect 7293 18790 7349 18846
rect 21192 18854 21256 18855
rect 21192 18791 21244 18854
rect 21244 18791 21256 18854
rect 7587 17980 7643 18036
rect 17762 18292 17826 18356
rect 20867 17982 20931 18046
rect 13067 17351 13131 17415
rect 12699 17071 12763 17135
rect 7291 16989 7347 17045
rect 21191 16989 21243 17051
rect 21243 16989 21255 17051
rect 21191 16987 21255 16989
rect 10594 16488 10658 16552
rect 17775 16490 17839 16554
rect 7589 16181 7645 16237
rect 14481 16376 14545 16440
rect 10874 15765 10938 15829
rect 12353 16207 12417 16271
rect 7291 15190 7347 15246
rect 12701 16208 12765 16272
rect 12499 14814 12563 14878
rect 7584 14382 7640 14438
rect 14228 16153 14292 16217
rect 20863 16177 20927 16241
rect 14481 15764 14545 15828
rect 14228 15679 14292 15743
rect 15729 15701 15793 15765
rect 16489 15701 16553 15765
rect 14839 15523 14903 15587
rect 15155 15523 15219 15587
rect 16777 15523 16841 15587
rect 17237 15527 17301 15591
rect 14177 15158 14241 15222
rect 21191 15252 21255 15256
rect 21191 15192 21243 15252
rect 21243 15192 21255 15252
rect 16278 14985 16342 15049
rect 14379 14807 14443 14871
rect 15947 14575 16011 14639
rect 16277 14575 16341 14639
rect 11404 14078 11468 14142
rect 11836 14078 11900 14142
rect 12479 14078 12543 14142
rect 12702 14078 12766 14142
rect 11404 13922 11468 13986
rect 7879 13390 7935 13446
rect 11404 13749 11468 13813
rect 11835 13748 11899 13812
rect 14377 14457 14441 14521
rect 15945 14237 16009 14301
rect 20864 14378 20928 14442
rect 15581 14057 15645 14121
rect 15579 13746 15643 13810
rect 14377 13218 14441 13282
rect 20575 13387 20639 13451
rect 8187 12582 8243 12638
rect 14379 12818 14443 12882
rect 20264 12636 20328 12641
rect 20264 12577 20279 12636
rect 20279 12577 20328 12636
rect 11611 12269 11675 12333
rect 12901 12269 12965 12333
rect 13401 12235 13465 12299
rect 15508 12299 15572 12363
rect 16497 12299 16561 12363
rect 14673 12121 14737 12185
rect 14965 12117 15029 12181
rect 16807 12117 16871 12181
rect 17223 12121 17287 12185
rect 11241 11936 11305 12000
rect 12001 11936 12065 12000
rect 15014 11936 15078 12000
rect 15397 11936 15461 12000
rect 7878 11591 7934 11647
rect 20574 11588 20638 11652
rect 23475 11373 23656 11592
rect 17771 11088 17835 11152
rect 12494 10944 12558 11008
rect 3448 5643 3540 5735
rect 4166 5258 4258 5350
rect 5462 4455 5864 4656
rect 5462 4254 5870 4455
rect 5664 4249 5870 4254
rect 8192 10783 8248 10839
rect 20269 10774 20281 10834
rect 20281 10774 20333 10834
rect 20269 10770 20333 10774
rect 11231 10377 11295 10441
rect 7871 9794 7935 9858
rect 10707 9521 10771 9585
rect 20574 9784 20638 9848
rect 17789 9296 17853 9360
rect 8186 8975 8247 9039
rect 8247 8975 8250 9039
rect 20268 8976 20280 9037
rect 20280 8976 20332 9037
rect 20268 8973 20332 8976
rect 8789 5648 8871 5730
rect 14863 5392 14921 5450
rect 11473 5263 11555 5345
rect 8757 4249 8881 4454
rect 6340 3184 6742 3586
rect 11452 3587 11478 3588
rect 11478 3587 11536 3588
rect 11536 3587 11558 3588
rect 11452 3379 11558 3587
rect 11452 3279 11561 3379
rect 11452 3182 11558 3279
rect 14863 3039 14921 3097
rect 17433 3007 17535 3008
rect 17432 2897 17542 3007
rect 17433 2803 17535 2897
rect 22387 2798 22593 3004
<< metal3 >>
rect 7289 20620 7353 20626
rect 7289 18851 7353 20556
rect 21191 20620 21255 20628
rect 7581 20222 7645 20228
rect 7288 18846 7354 18851
rect 7288 18790 7293 18846
rect 7349 18790 7354 18846
rect 7288 18785 7354 18790
rect 7289 17050 7353 18785
rect 7581 18041 7645 20158
rect 20857 20156 20867 20220
rect 20931 20156 20941 20220
rect 7872 19819 7936 19825
rect 20567 19756 20577 19820
rect 20641 19756 20651 19820
rect 7577 18036 7653 18041
rect 7577 17980 7587 18036
rect 7643 17980 7653 18036
rect 7577 17975 7653 17980
rect 7281 17045 7357 17050
rect 7281 16989 7291 17045
rect 7347 16989 7357 17045
rect 7281 16984 7357 16989
rect 7289 15251 7353 16984
rect 7581 16242 7645 17975
rect 7579 16237 7655 16242
rect 7579 16181 7589 16237
rect 7645 16181 7655 16237
rect 7579 16176 7655 16181
rect 7281 15246 7357 15251
rect 7281 15190 7291 15246
rect 7347 15190 7357 15246
rect 7281 15185 7357 15190
rect 7289 15183 7353 15185
rect 7581 14443 7645 16176
rect 7574 14438 7650 14443
rect 7574 14382 7584 14438
rect 7640 14382 7650 14438
rect 7574 14377 7650 14382
rect 7581 14374 7645 14377
rect 7872 13451 7936 19755
rect 8182 19421 8246 19427
rect 7869 13446 7945 13451
rect 7869 13390 7879 13446
rect 7935 13390 7945 13446
rect 7869 13385 7945 13390
rect 7872 11652 7936 13385
rect 8182 12643 8246 19357
rect 20259 19356 20269 19420
rect 20333 19356 20343 19420
rect 9271 17859 10429 19019
rect 11071 17859 12229 19019
rect 12871 17859 14029 19019
rect 14671 17859 15829 19019
rect 16471 17859 17629 19019
rect 17752 18356 17836 18361
rect 17752 18292 17762 18356
rect 17826 18292 17836 18356
rect 17752 18287 17836 18292
rect 13046 17415 13151 17439
rect 17762 17438 17826 18287
rect 18271 17859 19429 19019
rect 13046 17351 13067 17415
rect 13131 17351 13151 17415
rect 13046 17328 13151 17351
rect 17262 17374 17826 17438
rect 17262 17219 17326 17374
rect 9271 16059 10429 17219
rect 10574 16552 10680 16574
rect 10574 16488 10594 16552
rect 10658 16488 10680 16552
rect 10574 16467 10680 16488
rect 11071 16271 12229 17219
rect 12689 17135 12773 17140
rect 12871 17135 14029 17219
rect 12689 17071 12699 17135
rect 12763 17071 14029 17135
rect 12689 17066 12773 17071
rect 12343 16271 12427 16276
rect 11071 16207 12353 16271
rect 12417 16207 12427 16271
rect 11071 16059 12229 16207
rect 12343 16202 12427 16207
rect 12687 16272 12779 16305
rect 12687 16208 12701 16272
rect 12765 16208 12779 16272
rect 12687 16183 12779 16208
rect 12871 16059 14029 17071
rect 14671 16856 15829 17219
rect 14228 16792 15829 16856
rect 14228 16222 14292 16792
rect 14471 16440 14555 16469
rect 14471 16376 14481 16440
rect 14545 16376 14555 16440
rect 14471 16352 14555 16376
rect 14218 16217 14302 16222
rect 14218 16153 14228 16217
rect 14292 16153 14302 16217
rect 14218 16148 14302 16153
rect 14671 16059 15829 16792
rect 16471 16059 17629 17219
rect 17757 16554 17855 16573
rect 17757 16490 17775 16554
rect 17839 16490 17855 16554
rect 17757 16473 17855 16490
rect 18271 16059 19429 17219
rect 11615 15970 11679 16059
rect 11615 15906 16176 15970
rect 10833 15829 10973 15860
rect 10833 15765 10874 15829
rect 10938 15765 10973 15829
rect 10833 15731 10973 15765
rect 14450 15828 14579 15836
rect 14450 15764 14481 15828
rect 14545 15764 14579 15828
rect 14450 15756 14579 15764
rect 15719 15765 15803 15770
rect 14218 15743 14302 15748
rect 11825 15679 14228 15743
rect 14292 15679 14302 15743
rect 15719 15701 15729 15765
rect 15793 15701 15803 15765
rect 15719 15696 15803 15701
rect 11825 15419 11889 15679
rect 14218 15674 14302 15679
rect 14829 15587 14913 15592
rect 12312 15523 14839 15587
rect 14903 15523 14913 15587
rect 9271 14259 10429 15419
rect 11071 14259 12229 15419
rect 11404 14147 11468 14259
rect 11394 14142 11478 14147
rect 11394 14078 11404 14142
rect 11468 14078 11478 14142
rect 11394 14073 11478 14078
rect 11814 14142 11920 14160
rect 11814 14078 11836 14142
rect 11900 14078 11920 14142
rect 11404 13991 11468 14073
rect 11814 14063 11920 14078
rect 11394 13986 11478 13991
rect 11394 13922 11404 13986
rect 11468 13922 11478 13986
rect 11394 13917 11478 13922
rect 11404 13818 11468 13917
rect 11394 13813 11478 13818
rect 11394 13749 11404 13813
rect 11468 13749 11478 13813
rect 11394 13744 11478 13749
rect 11816 13817 11908 13842
rect 11816 13812 11909 13817
rect 11816 13748 11835 13812
rect 11899 13748 11909 13812
rect 11404 13619 11468 13744
rect 11816 13743 11909 13748
rect 11816 13720 11908 13743
rect 8177 12638 8253 12643
rect 8177 12582 8187 12638
rect 8243 12582 8253 12638
rect 8177 12577 8253 12582
rect 7868 11647 7944 11652
rect 7868 11591 7878 11647
rect 7934 11591 7944 11647
rect 7868 11586 7944 11591
rect 7872 9863 7936 11586
rect 8182 10844 8246 12577
rect 9271 12459 10429 13619
rect 11071 12459 12229 13619
rect 11241 12005 11305 12459
rect 11601 12333 11685 12338
rect 11601 12269 11611 12333
rect 11675 12269 11685 12333
rect 11601 12264 11685 12269
rect 11231 12000 11315 12005
rect 11231 11936 11241 12000
rect 11305 11936 11315 12000
rect 11231 11931 11315 11936
rect 11611 11819 11675 12264
rect 11981 12000 12082 12016
rect 11981 11936 12001 12000
rect 12065 11936 12082 12000
rect 11981 11918 12082 11936
rect 8182 10839 8258 10844
rect 8182 10783 8192 10839
rect 8248 10783 8258 10839
rect 8182 10778 8258 10783
rect 7861 9858 7945 9863
rect 7861 9794 7871 9858
rect 7935 9794 7945 9858
rect 7861 9789 7945 9794
rect 7872 9782 7936 9789
rect 8182 9044 8246 10778
rect 9271 10659 10429 11819
rect 11071 11013 12229 11819
rect 12312 11013 12376 15523
rect 14829 15518 14913 15523
rect 15132 15587 15242 15603
rect 15132 15523 15155 15587
rect 15219 15523 15242 15587
rect 15132 15509 15242 15523
rect 15729 15419 15793 15696
rect 12489 14878 12573 14883
rect 12871 14878 14029 15419
rect 14152 15222 14261 15245
rect 14152 15158 14177 15222
rect 14241 15158 14261 15222
rect 14152 15138 14261 15158
rect 12489 14814 12499 14878
rect 12563 14814 14029 14878
rect 12489 14809 12573 14814
rect 12871 14259 14029 14814
rect 14369 14871 14453 14876
rect 14671 14871 15829 15419
rect 14369 14807 14379 14871
rect 14443 14807 15829 14871
rect 14369 14802 14453 14807
rect 14354 14521 14460 14544
rect 14354 14457 14377 14521
rect 14441 14457 14460 14521
rect 14354 14437 14460 14457
rect 14671 14259 15829 14807
rect 15933 14639 16024 14678
rect 15933 14575 15947 14639
rect 16011 14575 16024 14639
rect 15933 14538 16024 14575
rect 15935 14301 16019 14306
rect 12468 14142 12555 14176
rect 12468 14078 12479 14142
rect 12543 14078 12555 14142
rect 12468 14047 12555 14078
rect 12692 14142 12776 14147
rect 12692 14078 12702 14142
rect 12766 14078 12776 14142
rect 12692 14073 12776 14078
rect 13419 14091 13483 14259
rect 15935 14237 15945 14301
rect 16009 14237 16019 14301
rect 15935 14232 16019 14237
rect 15550 14121 15675 14151
rect 11071 10949 12376 11013
rect 12476 11008 12574 11039
rect 11071 10659 12229 10949
rect 12476 10944 12494 11008
rect 12558 10944 12574 11008
rect 12702 11024 12766 14073
rect 13419 14027 14983 14091
rect 15550 14057 15581 14121
rect 15645 14057 15675 14121
rect 15550 14030 15675 14057
rect 14919 13619 14983 14027
rect 15557 13810 15661 13830
rect 15557 13746 15579 13810
rect 15643 13746 15661 13810
rect 15557 13730 15661 13746
rect 12871 12882 14029 13619
rect 14355 13282 14461 13304
rect 14355 13218 14377 13282
rect 14441 13218 14461 13282
rect 14355 13197 14461 13218
rect 14369 12882 14453 12887
rect 12871 12818 14379 12882
rect 14443 12818 14453 12882
rect 12871 12459 14029 12818
rect 14369 12813 14453 12818
rect 14671 12459 15829 13619
rect 12901 12338 12965 12459
rect 15508 12368 15572 12459
rect 15498 12363 15582 12368
rect 12891 12333 12975 12338
rect 12891 12269 12901 12333
rect 12965 12269 12975 12333
rect 12891 12264 12975 12269
rect 13378 12299 13486 12325
rect 13378 12235 13401 12299
rect 13465 12235 13486 12299
rect 15498 12299 15508 12363
rect 15572 12299 15582 12363
rect 15498 12294 15582 12299
rect 13378 12212 13486 12235
rect 14663 12185 14747 12190
rect 14154 12121 14673 12185
rect 14737 12121 14747 12185
rect 12871 11024 14029 11819
rect 12702 11022 14029 11024
rect 14154 11022 14218 12121
rect 14663 12116 14747 12121
rect 14944 12181 15049 12205
rect 14944 12117 14965 12181
rect 15029 12117 15049 12181
rect 14944 12096 15049 12117
rect 14994 12000 15095 12019
rect 14994 11936 15014 12000
rect 15078 11936 15095 12000
rect 14994 11921 15095 11936
rect 15387 12000 15471 12005
rect 15387 11936 15397 12000
rect 15461 11936 15471 12000
rect 15387 11931 15471 11936
rect 15397 11819 15461 11931
rect 12702 10960 14218 11022
rect 12476 10919 12574 10944
rect 12871 10958 14218 10960
rect 14671 11107 15829 11819
rect 15945 11107 16009 14232
rect 16112 11275 16176 15906
rect 16489 15770 16553 16059
rect 16479 15765 16563 15770
rect 16479 15701 16489 15765
rect 16553 15701 16563 15765
rect 16479 15696 16563 15701
rect 16754 15587 16864 15602
rect 17237 15596 17301 16059
rect 16754 15523 16777 15587
rect 16841 15523 16864 15587
rect 16754 15508 16864 15523
rect 17227 15591 17311 15596
rect 17227 15527 17237 15591
rect 17301 15527 17311 15591
rect 17227 15522 17311 15527
rect 16268 15049 16352 15054
rect 16471 15049 17629 15419
rect 16268 14985 16278 15049
rect 16342 14985 17629 15049
rect 16268 14980 16352 14985
rect 16264 14639 16355 14677
rect 16264 14575 16277 14639
rect 16341 14575 16355 14639
rect 16264 14537 16355 14575
rect 16471 14259 17629 14985
rect 18271 14259 19429 15419
rect 16471 12459 17629 13619
rect 18271 12459 19429 13619
rect 20270 12646 20334 19356
rect 20577 13456 20641 19756
rect 20867 18051 20931 20156
rect 21191 18860 21255 20556
rect 21182 18855 21266 18860
rect 21182 18791 21192 18855
rect 21256 18791 21266 18855
rect 21182 18786 21266 18791
rect 20857 18046 20941 18051
rect 20857 17982 20867 18046
rect 20931 17982 20941 18046
rect 20857 17977 20941 17982
rect 20867 16246 20931 17977
rect 21191 17056 21255 18786
rect 21181 17051 21265 17056
rect 21181 16987 21191 17051
rect 21255 16987 21265 17051
rect 21181 16982 21265 16987
rect 20853 16241 20937 16246
rect 20853 16177 20863 16241
rect 20927 16177 20937 16241
rect 20853 16172 20937 16177
rect 20867 14447 20931 16172
rect 21191 15261 21255 16982
rect 21181 15256 21265 15261
rect 21181 15192 21191 15256
rect 21255 15192 21265 15256
rect 21181 15187 21265 15192
rect 21191 15185 21255 15187
rect 20854 14442 20938 14447
rect 20854 14378 20864 14442
rect 20928 14378 20938 14442
rect 20854 14373 20938 14378
rect 20565 13451 20649 13456
rect 20565 13387 20575 13451
rect 20639 13387 20649 13451
rect 20565 13382 20649 13387
rect 20254 12641 20338 12646
rect 20254 12577 20264 12641
rect 20328 12577 20338 12641
rect 20254 12572 20338 12577
rect 16487 12363 16571 12368
rect 16487 12299 16497 12363
rect 16561 12299 16571 12363
rect 16487 12294 16571 12299
rect 16497 11819 16561 12294
rect 16786 12181 16891 12203
rect 17223 12190 17287 12459
rect 16786 12117 16807 12181
rect 16871 12117 16891 12181
rect 16786 12094 16891 12117
rect 17213 12185 17297 12190
rect 17213 12121 17223 12185
rect 17287 12121 17297 12185
rect 17213 12116 17297 12121
rect 16471 11275 17629 11819
rect 16112 11211 17629 11275
rect 14671 11043 16012 11107
rect 12871 10659 14029 10958
rect 14671 10659 15829 11043
rect 16471 10659 17629 11211
rect 17754 11152 17856 11173
rect 17754 11088 17771 11152
rect 17835 11088 17856 11152
rect 17754 11070 17856 11088
rect 18271 10659 19429 11819
rect 20270 10839 20334 12572
rect 20577 11657 20641 13382
rect 20564 11652 20648 11657
rect 20564 11588 20574 11652
rect 20638 11588 20648 11652
rect 20564 11583 20648 11588
rect 23462 11592 23668 11618
rect 20259 10834 20343 10839
rect 20259 10770 20269 10834
rect 20333 10770 20343 10834
rect 20259 10765 20343 10770
rect 11210 10441 11316 10464
rect 11210 10377 11231 10441
rect 11295 10377 11316 10441
rect 11210 10360 11316 10377
rect 17250 10217 17314 10659
rect 17250 10153 17853 10217
rect 8176 9039 8260 9044
rect 8176 8975 8186 9039
rect 8250 8975 8260 9039
rect 8176 8970 8260 8975
rect 9271 8859 10429 10019
rect 10693 9585 10791 9603
rect 10693 9521 10707 9585
rect 10771 9521 10791 9585
rect 10693 9500 10791 9521
rect 11071 8859 12229 10019
rect 12871 8859 14029 10019
rect 14671 8859 15829 10019
rect 16471 8859 17629 10019
rect 17789 9365 17853 10153
rect 17779 9360 17863 9365
rect 17779 9296 17789 9360
rect 17853 9296 17863 9360
rect 17779 9291 17863 9296
rect 17789 9287 17853 9291
rect 18271 8859 19429 10019
rect 20270 9042 20334 10765
rect 20577 9853 20641 11583
rect 23462 11373 23475 11592
rect 23656 11373 23668 11592
rect 20564 9848 20648 9853
rect 20564 9784 20574 9848
rect 20638 9784 20648 9848
rect 20564 9779 20648 9784
rect 20577 9770 20641 9779
rect 20258 9037 20342 9042
rect 20258 8973 20268 9037
rect 20332 8973 20342 9037
rect 20258 8968 20342 8973
rect 20270 8967 20334 8968
rect 3443 5735 3545 5740
rect 3443 5643 3448 5735
rect 3540 5730 8876 5735
rect 3540 5648 8789 5730
rect 8871 5648 8876 5730
rect 3540 5643 8876 5648
rect 3443 5638 3545 5643
rect 14853 5450 14931 5455
rect 14853 5392 14863 5450
rect 14921 5392 14931 5450
rect 4161 5350 4263 5355
rect 4161 5258 4166 5350
rect 4258 5345 11560 5350
rect 4258 5263 11473 5345
rect 11555 5263 11560 5345
rect 4258 5258 11560 5263
rect 4161 5253 4263 5258
rect 5457 4656 8891 4661
rect 5457 4254 5462 4656
rect 5864 4455 8891 4656
rect 5870 4454 8891 4455
rect 5457 4249 5664 4254
rect 5870 4249 8757 4454
rect 8881 4249 8891 4454
rect 5654 4244 5880 4249
rect 8747 4244 8891 4249
rect 14853 3833 14931 5392
rect 23462 3833 23668 11373
rect 13209 3627 23668 3833
rect 11442 3591 11568 3593
rect 6335 3588 11579 3591
rect 6335 3586 11452 3588
rect 6335 3394 6340 3586
rect 6333 3210 6340 3394
rect 6335 3184 6340 3210
rect 6742 3184 11452 3586
rect 11558 3379 11579 3588
rect 11561 3279 11579 3379
rect 6335 3182 11452 3184
rect 11558 3182 11579 3279
rect 6335 3179 11579 3182
rect 11442 3177 11568 3179
rect 13209 2681 13415 3627
rect 14853 3097 14931 3627
rect 14853 3039 14863 3097
rect 14921 3039 14931 3097
rect 14853 3030 14931 3039
rect 17423 3012 17545 3013
rect 17422 3008 17552 3012
rect 17422 3007 17433 3008
rect 17535 3007 17552 3008
rect 17422 2897 17432 3007
rect 17542 3006 17552 3007
rect 22377 3006 22603 3009
rect 17542 3004 22603 3006
rect 17542 2897 22387 3004
rect 17422 2892 17433 2897
rect 17423 2803 17433 2892
rect 17535 2803 22387 2897
rect 17423 2800 22387 2803
rect 17423 2798 17545 2800
rect 22377 2798 22387 2800
rect 22593 2798 22603 3004
rect 22377 2793 22603 2798
rect -170 2475 13415 2681
<< via3 >>
rect 7289 20556 7353 20620
rect 21191 20556 21255 20620
rect 7581 20158 7645 20222
rect 20867 20156 20931 20220
rect 7872 19755 7936 19819
rect 20577 19756 20641 19820
rect 8182 19357 8246 19421
rect 20269 19356 20333 19420
rect 13067 17351 13131 17415
rect 10594 16488 10658 16552
rect 12701 16208 12765 16272
rect 14481 16376 14545 16440
rect 17775 16490 17839 16554
rect 10874 15765 10938 15829
rect 14481 15764 14545 15828
rect 11836 14078 11900 14142
rect 11835 13748 11899 13812
rect 12001 11936 12065 12000
rect 15155 15523 15219 15587
rect 14177 15158 14241 15222
rect 14377 14457 14441 14521
rect 15947 14575 16011 14639
rect 12479 14078 12543 14142
rect 12494 10944 12558 11008
rect 15581 14057 15645 14121
rect 15579 13746 15643 13810
rect 14377 13218 14441 13282
rect 13401 12235 13465 12299
rect 14965 12117 15029 12181
rect 15014 11936 15078 12000
rect 16777 15523 16841 15587
rect 16277 14575 16341 14639
rect 16807 12117 16871 12181
rect 17771 11088 17835 11152
rect 11231 10377 11295 10441
rect 10707 9521 10771 9585
<< mimcap >>
rect 9371 18879 10331 18919
rect 9371 17999 9411 18879
rect 10291 17999 10331 18879
rect 9371 17959 10331 17999
rect 11171 18879 12131 18919
rect 11171 17999 11211 18879
rect 12091 17999 12131 18879
rect 11171 17959 12131 17999
rect 12971 18879 13931 18919
rect 12971 17999 13011 18879
rect 13891 17999 13931 18879
rect 12971 17959 13931 17999
rect 14771 18879 15731 18919
rect 14771 17999 14811 18879
rect 15691 17999 15731 18879
rect 14771 17959 15731 17999
rect 16571 18879 17531 18919
rect 16571 17999 16611 18879
rect 17491 17999 17531 18879
rect 16571 17959 17531 17999
rect 18371 18879 19331 18919
rect 18371 17999 18411 18879
rect 19291 17999 19331 18879
rect 18371 17959 19331 17999
rect 9371 17079 10331 17119
rect 9371 16199 9411 17079
rect 10291 16199 10331 17079
rect 9371 16159 10331 16199
rect 11171 17079 12131 17119
rect 11171 16199 11211 17079
rect 12091 16199 12131 17079
rect 11171 16159 12131 16199
rect 12971 17079 13931 17119
rect 12971 16199 13011 17079
rect 13891 16199 13931 17079
rect 12971 16159 13931 16199
rect 14771 17079 15731 17119
rect 14771 16199 14811 17079
rect 15691 16199 15731 17079
rect 14771 16159 15731 16199
rect 16571 17079 17531 17119
rect 16571 16199 16611 17079
rect 17491 16199 17531 17079
rect 16571 16159 17531 16199
rect 18371 17079 19331 17119
rect 18371 16199 18411 17079
rect 19291 16199 19331 17079
rect 18371 16159 19331 16199
rect 9371 15279 10331 15319
rect 9371 14399 9411 15279
rect 10291 14399 10331 15279
rect 9371 14359 10331 14399
rect 11171 15279 12131 15319
rect 11171 14399 11211 15279
rect 12091 14399 12131 15279
rect 11171 14359 12131 14399
rect 12971 15279 13931 15319
rect 12971 14399 13011 15279
rect 13891 14399 13931 15279
rect 12971 14359 13931 14399
rect 14771 15279 15731 15319
rect 14771 14399 14811 15279
rect 15691 14399 15731 15279
rect 14771 14359 15731 14399
rect 16571 15279 17531 15319
rect 16571 14399 16611 15279
rect 17491 14399 17531 15279
rect 16571 14359 17531 14399
rect 18371 15279 19331 15319
rect 18371 14399 18411 15279
rect 19291 14399 19331 15279
rect 18371 14359 19331 14399
rect 9371 13479 10331 13519
rect 9371 12599 9411 13479
rect 10291 12599 10331 13479
rect 9371 12559 10331 12599
rect 11171 13479 12131 13519
rect 11171 12599 11211 13479
rect 12091 12599 12131 13479
rect 11171 12559 12131 12599
rect 12971 13479 13931 13519
rect 12971 12599 13011 13479
rect 13891 12599 13931 13479
rect 12971 12559 13931 12599
rect 14771 13479 15731 13519
rect 14771 12599 14811 13479
rect 15691 12599 15731 13479
rect 14771 12559 15731 12599
rect 16571 13479 17531 13519
rect 16571 12599 16611 13479
rect 17491 12599 17531 13479
rect 16571 12559 17531 12599
rect 18371 13479 19331 13519
rect 18371 12599 18411 13479
rect 19291 12599 19331 13479
rect 18371 12559 19331 12599
rect 9371 11679 10331 11719
rect 9371 10799 9411 11679
rect 10291 10799 10331 11679
rect 9371 10759 10331 10799
rect 11171 11679 12131 11719
rect 11171 10799 11211 11679
rect 12091 10799 12131 11679
rect 11171 10759 12131 10799
rect 12971 11679 13931 11719
rect 12971 10799 13011 11679
rect 13891 10799 13931 11679
rect 12971 10759 13931 10799
rect 14771 11679 15731 11719
rect 14771 10799 14811 11679
rect 15691 10799 15731 11679
rect 14771 10759 15731 10799
rect 16571 11679 17531 11719
rect 16571 10799 16611 11679
rect 17491 10799 17531 11679
rect 16571 10759 17531 10799
rect 18371 11679 19331 11719
rect 18371 10799 18411 11679
rect 19291 10799 19331 11679
rect 18371 10759 19331 10799
rect 9371 9879 10331 9919
rect 9371 8999 9411 9879
rect 10291 8999 10331 9879
rect 9371 8959 10331 8999
rect 11171 9879 12131 9919
rect 11171 8999 11211 9879
rect 12091 8999 12131 9879
rect 11171 8959 12131 8999
rect 12971 9879 13931 9919
rect 12971 8999 13011 9879
rect 13891 8999 13931 9879
rect 12971 8959 13931 8999
rect 14771 9879 15731 9919
rect 14771 8999 14811 9879
rect 15691 8999 15731 9879
rect 14771 8959 15731 8999
rect 16571 9879 17531 9919
rect 16571 8999 16611 9879
rect 17491 8999 17531 9879
rect 16571 8959 17531 8999
rect 18371 9879 19331 9919
rect 18371 8999 18411 9879
rect 19291 8999 19331 9879
rect 18371 8959 19331 8999
<< mimcapcontact >>
rect 9411 17999 10291 18879
rect 11211 17999 12091 18879
rect 13011 17999 13891 18879
rect 14811 17999 15691 18879
rect 16611 17999 17491 18879
rect 18411 17999 19291 18879
rect 9411 16199 10291 17079
rect 11211 16199 12091 17079
rect 13011 16199 13891 17079
rect 14811 16199 15691 17079
rect 16611 16199 17491 17079
rect 18411 16199 19291 17079
rect 9411 14399 10291 15279
rect 11211 14399 12091 15279
rect 13011 14399 13891 15279
rect 14811 14399 15691 15279
rect 16611 14399 17491 15279
rect 18411 14399 19291 15279
rect 9411 12599 10291 13479
rect 11211 12599 12091 13479
rect 13011 12599 13891 13479
rect 14811 12599 15691 13479
rect 16611 12599 17491 13479
rect 18411 12599 19291 13479
rect 9411 10799 10291 11679
rect 11211 10799 12091 11679
rect 13011 10799 13891 11679
rect 14811 10799 15691 11679
rect 16611 10799 17491 11679
rect 18411 10799 19291 11679
rect 9411 8999 10291 9879
rect 11211 8999 12091 9879
rect 13011 8999 13891 9879
rect 14811 8999 15691 9879
rect 16611 8999 17491 9879
rect 18411 8999 19291 9879
<< metal4 >>
rect 7288 20620 7354 20621
rect 21190 20620 21256 20621
rect 7272 20556 7289 20620
rect 7353 20556 21191 20620
rect 21255 20556 21256 20620
rect 7288 20555 7354 20556
rect 21190 20555 21256 20556
rect 7580 20222 7646 20223
rect 7580 20220 7581 20222
rect 7272 20158 7581 20220
rect 7645 20220 7646 20222
rect 20866 20220 20932 20221
rect 7645 20158 20867 20220
rect 7272 20156 20867 20158
rect 20931 20156 21255 20220
rect 20866 20155 20932 20156
rect 20576 19820 20642 19821
rect 7272 19819 20577 19820
rect 7272 19756 7872 19819
rect 7871 19755 7872 19756
rect 7936 19756 20577 19819
rect 20641 19756 21255 19820
rect 7936 19755 7937 19756
rect 20576 19755 20642 19756
rect 7871 19754 7937 19755
rect 8181 19421 8247 19422
rect 8181 19420 8182 19421
rect 7272 19357 8182 19420
rect 8246 19420 8247 19421
rect 20268 19420 20334 19421
rect 8246 19357 20269 19420
rect 7272 19356 20269 19357
rect 20333 19356 21255 19420
rect 20268 19355 20334 19356
rect 9410 18879 10292 18880
rect 9410 17999 9411 18879
rect 10291 17999 10292 18879
rect 9410 17998 10292 17999
rect 11210 18879 12092 18880
rect 11210 17999 11211 18879
rect 12091 17999 12092 18879
rect 11210 17998 12092 17999
rect 13010 18879 13892 18880
rect 13010 17999 13011 18879
rect 13891 17999 13892 18879
rect 13010 17998 13892 17999
rect 14810 18879 15692 18880
rect 14810 17999 14811 18879
rect 15691 17999 15692 18879
rect 14810 17998 15692 17999
rect 16610 18879 17492 18880
rect 16610 17999 16611 18879
rect 17491 17999 17492 18879
rect 16610 17998 17492 17999
rect 18410 18879 19292 18880
rect 18410 17999 18411 18879
rect 19291 17999 19292 18879
rect 18410 17998 19292 17999
rect 13066 17415 13132 17416
rect 13066 17351 13067 17415
rect 13131 17351 13132 17415
rect 13066 17350 13132 17351
rect 13067 17080 13131 17350
rect 9410 17079 10292 17080
rect 9410 16199 9411 17079
rect 10291 16199 10292 17079
rect 11210 17079 12092 17080
rect 10593 16552 10659 16553
rect 11210 16552 11211 17079
rect 10593 16488 10594 16552
rect 10658 16488 11211 16552
rect 10593 16487 10659 16488
rect 9410 16198 10292 16199
rect 11210 16199 11211 16488
rect 12091 16199 12092 17079
rect 13010 17079 13892 17080
rect 12700 16272 12766 16273
rect 13010 16272 13011 17079
rect 12700 16208 12701 16272
rect 12765 16208 13011 16272
rect 12700 16207 12766 16208
rect 11210 16198 12092 16199
rect 13010 16199 13011 16208
rect 13891 16199 13892 17079
rect 14810 17079 15692 17080
rect 14480 16440 14546 16441
rect 14810 16440 14811 17079
rect 14480 16376 14481 16440
rect 14545 16376 14811 16440
rect 14480 16375 14546 16376
rect 13010 16198 13892 16199
rect 14810 16199 14811 16376
rect 15691 16199 15692 17079
rect 14810 16198 15692 16199
rect 16610 17079 17492 17080
rect 16610 16199 16611 17079
rect 17491 16554 17492 17079
rect 18410 17079 19292 17080
rect 17774 16554 17840 16555
rect 17491 16490 17775 16554
rect 17839 16490 17840 16554
rect 17491 16199 17492 16490
rect 17774 16489 17840 16490
rect 16610 16198 17492 16199
rect 18410 16199 18411 17079
rect 19291 16199 19292 17079
rect 18410 16198 19292 16199
rect 11615 15970 11679 16198
rect 11615 15906 16176 15970
rect 10873 15829 10939 15830
rect 10873 15765 10874 15829
rect 10938 15828 10939 15829
rect 14480 15828 14546 15829
rect 10938 15765 14481 15828
rect 10873 15764 14481 15765
rect 14545 15764 14546 15828
rect 11391 15280 11455 15764
rect 14480 15763 14546 15764
rect 15154 15587 15220 15588
rect 12313 15523 15155 15587
rect 15219 15523 15221 15587
rect 9410 15279 10292 15280
rect 9410 14399 9411 15279
rect 10291 14399 10292 15279
rect 9410 14398 10292 14399
rect 11210 15279 12092 15280
rect 11210 14399 11211 15279
rect 12091 14399 12092 15279
rect 11210 14398 12092 14399
rect 11836 14143 11900 14398
rect 11835 14142 11901 14143
rect 11835 14078 11836 14142
rect 11900 14078 11901 14142
rect 11835 14077 11901 14078
rect 11834 13812 11900 13813
rect 11834 13748 11835 13812
rect 11899 13748 11900 13812
rect 11834 13747 11900 13748
rect 11835 13480 11899 13747
rect 9410 13479 10292 13480
rect 9410 12599 9411 13479
rect 10291 12599 10292 13479
rect 11210 13479 12092 13480
rect 11210 12708 11211 13479
rect 9410 12598 10292 12599
rect 10707 12644 11211 12708
rect 9410 11679 10292 11680
rect 9410 10799 9411 11679
rect 10291 10799 10292 11679
rect 9410 10798 10292 10799
rect 9410 9879 10292 9880
rect 9410 8999 9411 9879
rect 10291 8999 10292 9879
rect 10707 9586 10771 12644
rect 11210 12599 11211 12644
rect 12091 12599 12092 13479
rect 11210 12598 12092 12599
rect 12001 12001 12065 12598
rect 12000 12000 12066 12001
rect 12000 11936 12001 12000
rect 12065 11936 12066 12000
rect 12000 11935 12066 11936
rect 11210 11679 12092 11680
rect 11210 10799 11211 11679
rect 12091 11518 12092 11679
rect 12313 11518 12377 15523
rect 15154 15522 15220 15523
rect 13010 15279 13892 15280
rect 13010 14399 13011 15279
rect 13891 15222 13892 15279
rect 14810 15279 15692 15280
rect 14176 15222 14242 15223
rect 13891 15158 14177 15222
rect 14241 15158 14242 15222
rect 13891 14399 13892 15158
rect 14176 15157 14242 15158
rect 14376 14521 14442 14522
rect 14810 14521 14811 15279
rect 14376 14457 14377 14521
rect 14441 14457 14811 14521
rect 14376 14456 14442 14457
rect 13010 14398 13892 14399
rect 14810 14399 14811 14457
rect 15691 14399 15692 15279
rect 15946 14639 16012 14640
rect 15946 14575 15947 14639
rect 16011 14575 16012 14639
rect 15946 14574 16012 14575
rect 14810 14398 15692 14399
rect 12478 14142 12544 14143
rect 12478 14078 12479 14142
rect 12543 14078 12544 14142
rect 12478 14077 12544 14078
rect 13419 14091 13483 14398
rect 15581 14122 15645 14398
rect 15580 14121 15646 14122
rect 12091 11454 12377 11518
rect 12479 11472 12543 14077
rect 13419 14027 14983 14091
rect 15580 14057 15581 14121
rect 15645 14057 15646 14121
rect 15580 14056 15646 14057
rect 14919 13480 14983 14027
rect 15578 13810 15644 13811
rect 15578 13746 15579 13810
rect 15643 13746 15644 13810
rect 15578 13745 15644 13746
rect 15579 13480 15643 13745
rect 13010 13479 13892 13480
rect 13010 12599 13011 13479
rect 13891 13282 13892 13479
rect 14810 13479 15692 13480
rect 14376 13282 14442 13283
rect 13891 13218 14377 13282
rect 14441 13218 14442 13282
rect 13891 12599 13892 13218
rect 14376 13217 14442 13218
rect 13010 12598 13892 12599
rect 14810 12599 14811 13479
rect 15691 12599 15692 13479
rect 14810 12598 15692 12599
rect 13401 12300 13465 12598
rect 13400 12299 13466 12300
rect 13400 12235 13401 12299
rect 13465 12235 13466 12299
rect 13400 12234 13466 12235
rect 14964 12181 15030 12182
rect 14154 12117 14965 12181
rect 15029 12117 15030 12181
rect 13010 11679 13892 11680
rect 13010 11472 13011 11679
rect 12091 10799 12092 11454
rect 12479 11408 13011 11472
rect 12493 11008 12559 11009
rect 13010 11008 13011 11408
rect 12491 10944 12494 11008
rect 12558 10944 13011 11008
rect 12493 10943 12559 10944
rect 11210 10798 12092 10799
rect 13010 10799 13011 10944
rect 13891 11471 13892 11679
rect 14154 11471 14218 12117
rect 14964 12116 15030 12117
rect 15014 12001 15078 12004
rect 15013 12000 15079 12001
rect 15013 11936 15014 12000
rect 15078 11936 15079 12000
rect 15013 11935 15079 11936
rect 15014 11680 15078 11935
rect 13891 11407 14218 11471
rect 14810 11679 15692 11680
rect 13891 10799 13892 11407
rect 13010 10798 13892 10799
rect 14810 10799 14811 11679
rect 15691 11503 15692 11679
rect 15947 11503 16011 14574
rect 15691 11439 16011 11503
rect 15691 10799 15692 11439
rect 16112 11275 16176 15906
rect 16777 15588 16841 16198
rect 16776 15587 16842 15588
rect 16776 15523 16777 15587
rect 16841 15523 16842 15587
rect 16776 15522 16842 15523
rect 16610 15279 17492 15280
rect 16276 14639 16342 14640
rect 16610 14639 16611 15279
rect 16276 14575 16277 14639
rect 16341 14575 16611 14639
rect 16276 14574 16342 14575
rect 16610 14399 16611 14575
rect 17491 14399 17492 15279
rect 16610 14398 17492 14399
rect 18410 15279 19292 15280
rect 18410 14399 18411 15279
rect 19291 14399 19292 15279
rect 18410 14398 19292 14399
rect 16610 13479 17492 13480
rect 16610 12599 16611 13479
rect 17491 12599 17492 13479
rect 16610 12598 17492 12599
rect 18410 13479 19292 13480
rect 18410 12599 18411 13479
rect 19291 12599 19292 13479
rect 18410 12598 19292 12599
rect 16807 12182 16871 12598
rect 16806 12181 16872 12182
rect 16806 12117 16807 12181
rect 16871 12117 16872 12181
rect 16806 12116 16872 12117
rect 16610 11679 17492 11680
rect 16610 11275 16611 11679
rect 16112 11211 16611 11275
rect 14810 10798 15692 10799
rect 16610 10799 16611 11211
rect 17491 11152 17492 11679
rect 18410 11679 19292 11680
rect 17770 11152 17836 11153
rect 17491 11088 17771 11152
rect 17835 11088 17837 11152
rect 17491 10799 17492 11088
rect 17770 11087 17836 11088
rect 16610 10798 17492 10799
rect 18410 10799 18411 11679
rect 19291 10799 19292 11679
rect 18410 10798 19292 10799
rect 11231 10442 11295 10798
rect 11230 10441 11296 10442
rect 11230 10377 11231 10441
rect 11295 10377 11296 10441
rect 11230 10376 11296 10377
rect 11210 9879 12092 9880
rect 10706 9585 10772 9586
rect 10706 9521 10707 9585
rect 10771 9521 10772 9585
rect 10706 9520 10772 9521
rect 9410 8998 10292 8999
rect 11210 8999 11211 9879
rect 12091 8999 12092 9879
rect 11210 8998 12092 8999
rect 13010 9879 13892 9880
rect 13010 8999 13011 9879
rect 13891 8999 13892 9879
rect 13010 8998 13892 8999
rect 14810 9879 15692 9880
rect 14810 8999 14811 9879
rect 15691 8999 15692 9879
rect 14810 8998 15692 8999
rect 16610 9879 17492 9880
rect 16610 8999 16611 9879
rect 17491 8999 17492 9879
rect 16610 8998 17492 8999
rect 18410 9879 19292 9880
rect 18410 8999 18411 9879
rect 19291 8999 19292 9879
rect 18410 8998 19292 8999
<< labels >>
flabel metal1 2965 4960 2965 4960 1 FreeSans 800 0 0 0 in
port 2 n
flabel metal1 4751 4964 4751 4964 1 FreeSans 800 0 0 0 ip
port 1 n
flabel metal4 7524 20588 7524 20588 1 FreeSans 800 0 0 0 p2_b
port 6 n
flabel metal4 7520 20183 7520 20183 1 FreeSans 800 0 0 0 p2
port 5 n
flabel metal4 7522 19788 7522 19788 1 FreeSans 800 0 0 0 p1_b
port 4 n
flabel metal4 7522 19380 7522 19380 1 FreeSans 800 0 0 0 p1
port 3 n
flabel metal2 5790 8141 5790 8141 1 FreeSans 800 0 0 0 op
port 7 n
flabel metal2 6403 8150 6403 8150 1 FreeSans 800 0 0 0 on
port 8 n
flabel metal1 22248 1153 22248 1153 1 FreeSans 800 0 0 0 i_bias
port 9 n
flabel metal3 -153 2588 -153 2588 1 FreeSans 800 0 0 0 cm
port 10 n
flabel locali 6730 20089 6730 20089 1 FreeSans 800 0 0 0 VDD
port 16 n power bidirectional
flabel locali 11 93 11 93 1 FreeSans 800 0 0 0 VSS
port 17 n power bidirectional
flabel metal2 22492 5814 22492 5814 1 FreeSans 800 0 0 0 bias_a
port 11 n
flabel metal2 19379 5290 19379 5290 1 FreeSans 800 0 0 0 bias_c
port 13 n
flabel metal2 20397 5292 20397 5292 1 FreeSans 800 0 0 0 bias_b
port 12 n
flabel metal2 708 5110 708 5110 1 FreeSans 800 0 0 0 cmc
port 15 n
flabel metal1 16024 4072 16024 4072 1 FreeSans 800 0 0 0 bias_d
port 14 n
flabel metal1 714 3718 714 3718 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/cmc
flabel metal1 4751 5099 4751 5099 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/ip
flabel metal1 2965 5094 2965 5094 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/in
flabel metal1 14888 2933 14888 2933 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_e
flabel metal1 21565 1108 21565 1108 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/i_bias
flabel metal1 22056 80 22056 80 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/VSS
flabel metal1 21868 6983 21868 6983 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/VDD
flabel metal1 5374 348 5374 348 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_a
flabel metal2 11509 4000 11509 4000 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/on
flabel metal2 8818 4007 8818 4007 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/op
flabel metal2 20392 5317 20392 5317 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_b
flabel space 13687 4065 13687 4065 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_d
flabel metal2 20456 2783 20456 2783 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_c
flabel metal2 20358 5383 20358 5383 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/bias_b
flabel metal3 14892 3288 14892 3288 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/bias_e
flabel metal2 20451 2884 20451 2884 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/bias_c
flabel metal1 21684 1146 21684 1146 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/i_bias
flabel metal1 13352 4057 13352 4057 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/bias_d
flabel metal1 13085 361 13085 361 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/bias_a
flabel locali 21942 86 21942 86 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/VSS
flabel locali 22031 6978 22031 6978 1 FreeSans 800 0 0 0 ota_v2_without_cmfb_0/bias_circuit_0/VDD
flabel metal1 5767 14028 5767 14028 1 FreeSans 400 0 0 0 sc_cmfb_0/op
flabel metal1 6379 14027 6379 14027 1 FreeSans 400 0 0 0 sc_cmfb_0/on
flabel metal1 6839 14030 6839 14030 1 FreeSans 400 0 0 0 sc_cmfb_0/cmc
flabel metal1 21971 13954 21971 13954 1 FreeSans 400 0 0 0 sc_cmfb_0/cm
flabel metal1 22473 13957 22473 13957 1 FreeSans 400 0 0 0 sc_cmfb_0/bias_a
flabel locali 9169 20082 9169 20082 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel locali 9187 19124 9187 19124 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal4 7420 20585 7420 20585 1 FreeSans 400 0 0 0 sc_cmfb_0/p2_b
flabel metal4 7418 20189 7418 20189 1 FreeSans 400 0 0 0 sc_cmfb_0/p2
flabel metal4 7419 19782 7419 19782 1 FreeSans 400 0 0 0 sc_cmfb_0/p1_b
flabel metal4 7418 19392 7418 19392 1 FreeSans 400 0 0 0 sc_cmfb_0/p1
flabel locali 7206 8912 7206 8912 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/VSS
flabel locali 7206 9920 7206 9920 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/VDD
flabel metal1 8428 9320 8428 9320 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/in
flabel metal1 7320 9322 7320 9322 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/out
flabel locali 8306 9008 8306 9008 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/en
flabel locali 8306 9820 8306 9820 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/en_b
flabel locali 20136 8912 20136 8912 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/VSS
flabel locali 20136 9920 20136 9920 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/VDD
flabel metal1 21358 9320 21358 9320 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/in
flabel metal1 20250 9322 20250 9322 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/out
flabel locali 21236 9008 21236 9008 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/en
flabel locali 21236 9820 21236 9820 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/en_b
flabel locali 7206 10712 7206 10712 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/VSS
flabel locali 7206 11720 7206 11720 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/VDD
flabel metal1 8428 11120 8428 11120 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/in
flabel metal1 7320 11122 7320 11122 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/out
flabel locali 8306 10808 8306 10808 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/en
flabel locali 8306 11620 8306 11620 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/en_b
flabel locali 20136 10712 20136 10712 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/VSS
flabel locali 20136 11720 20136 11720 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/VDD
flabel metal1 21358 11120 21358 11120 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/in
flabel metal1 20250 11122 20250 11122 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/out
flabel locali 21236 10808 21236 10808 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/en
flabel locali 21236 11620 21236 11620 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/en_b
flabel locali 7206 12512 7206 12512 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/VSS
flabel locali 7206 13520 7206 13520 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/VDD
flabel metal1 8428 12920 8428 12920 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/in
flabel metal1 7320 12922 7320 12922 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/out
flabel locali 8306 12608 8306 12608 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/en
flabel locali 8306 13420 8306 13420 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/en_b
flabel locali 20136 12512 20136 12512 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/VSS
flabel locali 20136 13520 20136 13520 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/VDD
flabel metal1 21358 12920 21358 12920 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/in
flabel metal1 20250 12922 20250 12922 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/out
flabel locali 21236 12608 21236 12608 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/en
flabel locali 21236 13420 21236 13420 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/en_b
flabel locali 7206 14312 7206 14312 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/VSS
flabel locali 7206 15320 7206 15320 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/VDD
flabel metal1 8428 14720 8428 14720 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/in
flabel metal1 7320 14722 7320 14722 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/out
flabel locali 8306 14408 8306 14408 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/en
flabel locali 8306 15220 8306 15220 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/en_b
flabel locali 20136 14312 20136 14312 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/VSS
flabel locali 20136 15320 20136 15320 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/VDD
flabel metal1 21358 14720 21358 14720 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/in
flabel metal1 20250 14722 20250 14722 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/out
flabel locali 21236 14408 21236 14408 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/en
flabel locali 21236 15220 21236 15220 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/en_b
flabel locali 7206 16112 7206 16112 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/VSS
flabel locali 7206 17120 7206 17120 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/VDD
flabel metal1 8428 16520 8428 16520 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/in
flabel metal1 7320 16522 7320 16522 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/out
flabel locali 8306 16208 8306 16208 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/en
flabel locali 8306 17020 8306 17020 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/en_b
flabel locali 20136 16112 20136 16112 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/VSS
flabel locali 20136 17120 20136 17120 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/VDD
flabel metal1 21358 16520 21358 16520 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/in
flabel metal1 20250 16522 20250 16522 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/out
flabel locali 21236 16208 21236 16208 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/en
flabel locali 21236 17020 21236 17020 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/en_b
flabel locali 7206 17912 7206 17912 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/VSS
flabel locali 7206 18920 7206 18920 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/VDD
flabel metal1 8428 18320 8428 18320 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/in
flabel metal1 7320 18322 7320 18322 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/out
flabel locali 8306 18008 8306 18008 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/en
flabel locali 8306 18820 8306 18820 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/en_b
flabel locali 20136 17912 20136 17912 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/VSS
flabel locali 20136 18920 20136 18920 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/VDD
flabel metal1 21358 18320 21358 18320 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/in
flabel metal1 20250 18322 20250 18322 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/out
flabel locali 21236 18008 21236 18008 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/en
flabel locali 21236 18820 21236 18820 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/en_b
<< end >>
