magic
tech sky130A
magscale 1 2
timestamp 1654583406
<< locali >>
rect 10718 21777 10827 21811
rect 5641 21403 5675 21607
rect 5457 21369 5675 21403
rect 5457 19703 5491 21369
rect 6929 20689 7406 20723
rect 6929 20655 6963 20689
rect 6670 20621 6963 20655
rect 5457 19669 5675 19703
rect 5641 19567 5675 19669
rect 5641 19533 5934 19567
rect 11253 18513 11362 18547
rect 11253 18309 11287 18513
rect 14933 18377 15042 18411
rect 13461 17935 13495 18139
rect 13386 17901 13495 17935
rect 19625 17459 19659 17595
rect 5641 17425 6118 17459
rect 19550 17425 19659 17459
rect 5641 17323 5675 17425
rect 5457 17289 5675 17323
rect 5457 15895 5491 17289
rect 22586 16813 23155 16847
rect 21833 16439 21867 16507
rect 21758 16405 21867 16439
rect 23121 16371 23155 16813
rect 22517 16337 23155 16371
rect 23121 16235 23155 16337
rect 23121 16201 23339 16235
rect 5457 15861 5675 15895
rect 5641 15759 5675 15861
rect 5917 15793 6118 15827
rect 5917 15759 5951 15793
rect 5641 15725 5951 15759
rect 18613 15759 18647 15827
rect 18613 15725 18814 15759
rect 15686 15589 15795 15623
rect 14565 15283 14599 15419
rect 11529 15249 11638 15283
rect 14490 15249 14599 15283
rect 23305 14739 23339 16201
rect 23121 14705 23339 14739
rect 12817 14637 12926 14671
rect 12817 14569 12851 14637
rect 15209 14569 15303 14603
rect 23121 14501 23155 14705
rect 11529 14195 11563 14331
rect 15669 14195 15703 14331
rect 11529 14161 11638 14195
rect 15669 14161 15778 14195
rect 22402 14161 22678 14195
rect 22477 14025 22511 14161
rect 7573 13617 7659 13651
rect 7573 13413 7607 13617
rect 16069 13549 16163 13583
rect 22954 13481 23155 13515
rect 12817 13413 12926 13447
rect 17081 13209 17175 13243
rect 8602 13073 9783 13107
rect 10057 13073 10166 13107
rect 16405 13073 16514 13107
rect 10057 13005 10091 13073
rect 23121 13005 23155 13481
rect 23029 12937 23155 12971
rect 23121 12495 23155 12937
rect 10977 12461 11454 12495
rect 22954 12461 23155 12495
rect 15778 12325 15887 12359
rect 11178 11985 11287 12019
rect 22862 11985 23155 12019
rect 23121 11883 23155 11985
rect 6101 11849 6210 11883
rect 21942 11849 22034 11883
rect 23121 11849 23247 11883
rect 6101 11781 6135 11849
rect 11253 11577 11347 11611
rect 5641 11373 6026 11407
rect 5641 10999 5675 11373
rect 23213 11271 23247 11849
rect 23121 11237 23247 11271
rect 23121 10999 23155 11237
rect 5641 10965 5767 10999
rect 5733 10795 5767 10965
rect 6210 10897 6411 10931
rect 6377 10863 6411 10897
rect 6469 10863 6503 10999
rect 22862 10965 23155 10999
rect 19901 10897 20470 10931
rect 19901 10863 19935 10897
rect 6377 10829 6578 10863
rect 19642 10829 19935 10863
rect 5733 10761 6026 10795
rect 23213 10523 23247 11067
rect 22770 10489 23247 10523
rect 16069 10285 16163 10319
rect 7021 9809 7483 9843
rect 7021 9775 7055 9809
rect 6762 9741 7055 9775
rect 11897 8687 11931 8823
rect 13938 8721 14139 8755
rect 19090 8721 19291 8755
rect 22218 8721 22310 8755
rect 11822 8653 11931 8687
rect 14105 8517 14139 8721
rect 6009 7497 6118 7531
rect 6009 7429 6043 7497
rect 5641 7021 5934 7055
rect 13110 7021 13202 7055
rect 5641 6579 5675 7021
rect 15502 6885 15795 6919
rect 5641 6545 5934 6579
rect 7665 6545 7774 6579
rect 12357 6545 12466 6579
rect 5641 5967 5675 6545
rect 5825 6341 5859 6545
rect 7665 6409 7699 6545
rect 12357 6409 12391 6545
rect 12817 6511 12851 6715
rect 19090 6545 19167 6579
rect 19533 6545 19642 6579
rect 19941 6545 20119 6579
rect 12817 6477 12926 6511
rect 19533 6409 19567 6545
rect 20085 6341 20119 6545
rect 8125 5967 8159 6171
rect 8878 6001 9062 6035
rect 10057 5967 10091 6103
rect 10718 6069 10827 6103
rect 10793 6001 10827 6069
rect 13386 6001 13495 6035
rect 13461 5967 13495 6001
rect 18153 5967 18187 6171
rect 18981 6001 19090 6035
rect 5641 5933 6210 5967
rect 8050 5933 8159 5967
rect 9522 5933 9798 5967
rect 9982 5933 10091 5967
rect 10241 5933 10442 5967
rect 13461 5933 14030 5967
rect 18153 5933 18262 5967
rect 9597 5797 9631 5933
rect 10241 5865 10275 5933
<< metal1 >>
rect 216 24500 12296 24528
rect 5796 21984 23000 22080
rect 9232 21848 10640 21876
rect 9232 21808 9260 21848
rect 7576 21780 7880 21808
rect 9048 21780 9260 21808
rect 10612 21808 10640 21848
rect 10612 21780 10824 21808
rect 11440 21780 11836 21808
rect 5828 21712 7052 21740
rect 7595 21712 7682 21740
rect 9140 21712 10088 21740
rect 5828 21604 5856 21712
rect 5644 21576 5856 21604
rect 7024 21604 7052 21712
rect 10428 21672 10456 21740
rect 10520 21712 11652 21740
rect 11716 21712 13400 21740
rect 15488 21712 16528 21740
rect 19076 21712 21588 21740
rect 9232 21644 9444 21672
rect 10428 21644 11284 21672
rect 16684 21644 16988 21672
rect 20088 21644 20208 21672
rect 7024 21576 7236 21604
rect 9876 21576 9996 21604
rect 12011 21576 12098 21604
rect 16224 21576 16344 21604
rect 20272 21576 20576 21604
rect 5796 21440 23000 21536
rect 13299 21372 13386 21400
rect 16887 21372 16974 21400
rect 17420 21338 18184 21366
rect 17420 21332 17448 21338
rect 9968 21304 10088 21332
rect 11624 21304 12112 21332
rect 13096 21304 14044 21332
rect 14660 21304 15148 21332
rect 15488 21304 16804 21332
rect 7852 21236 8616 21264
rect 8772 21236 8892 21264
rect 13096 21236 13124 21304
rect 14660 21264 14688 21304
rect 14476 21236 14688 21264
rect 16776 21264 16804 21304
rect 17236 21304 17448 21332
rect 18156 21332 18184 21338
rect 18156 21304 18368 21332
rect 17236 21264 17264 21304
rect 18340 21264 18368 21304
rect 16776 21236 17264 21264
rect 17512 21236 18276 21264
rect 18340 21236 19104 21264
rect 19168 21236 19932 21264
rect 7852 21196 7880 21236
rect 6564 21168 7880 21196
rect 8588 21196 8616 21236
rect 8588 21168 9076 21196
rect 9876 21168 12204 21196
rect 13188 21168 13492 21196
rect 14200 21168 14320 21196
rect 15304 21168 15516 21196
rect 15580 21168 16252 21196
rect 17420 21168 17632 21196
rect 15488 21128 15516 21168
rect 16224 21128 16252 21168
rect 15488 21100 15884 21128
rect 16224 21100 17264 21128
rect 17236 21060 17264 21100
rect 7944 21032 8616 21060
rect 8680 21032 9444 21060
rect 10428 21032 10548 21060
rect 11919 21032 12006 21060
rect 12544 21032 12664 21060
rect 14384 21032 14872 21060
rect 15672 21032 15976 21060
rect 17236 21032 17816 21060
rect 18727 21032 18814 21060
rect 5796 20896 23000 20992
rect 7852 20828 8248 20856
rect 11551 20828 11638 20856
rect 11808 20828 14504 20856
rect 17328 20828 17448 20856
rect 10505 20760 10609 20788
rect 11992 20760 13109 20788
rect 16151 20760 16252 20788
rect 18727 20760 18828 20788
rect 20272 20760 20837 20788
rect 7852 20726 8524 20754
rect 7852 20720 7880 20726
rect 7668 20692 7880 20720
rect 8496 20720 8524 20726
rect 13280 20726 13860 20754
rect 13280 20720 13308 20726
rect 8496 20692 8708 20720
rect 9876 20692 9996 20720
rect 12636 20692 13308 20720
rect 13832 20720 13860 20726
rect 13832 20692 15516 20720
rect 15875 20692 15962 20720
rect 20364 20692 20576 20720
rect 7668 20652 7696 20692
rect 12636 20652 12664 20692
rect 5920 20624 7696 20652
rect 7871 20624 7958 20652
rect 8050 20624 8137 20652
rect 8496 20624 8616 20652
rect 9232 20624 9812 20652
rect 10171 20624 10258 20652
rect 12176 20624 12664 20652
rect 12747 20624 12834 20652
rect 14292 20624 14412 20652
rect 18451 20624 18538 20652
rect 12636 20556 12756 20584
rect 6288 20488 6408 20516
rect 8864 20488 9076 20516
rect 10152 20488 10456 20516
rect 11624 20488 11836 20516
rect 12176 20488 12388 20516
rect 14587 20488 14674 20516
rect 18708 20488 19932 20516
rect 21744 20488 21956 20516
rect 5796 20352 23000 20448
rect 7668 20284 9168 20312
rect 13391 20284 13478 20312
rect 18248 20284 18920 20312
rect 19720 20284 19932 20312
rect 8496 20216 8892 20244
rect 15396 20216 15700 20244
rect 15488 20148 15608 20176
rect 21376 20148 22324 20176
rect 6104 20080 6316 20108
rect 6380 20080 6577 20108
rect 9048 20080 9643 20108
rect 9876 20080 10272 20108
rect 11624 20080 12112 20108
rect 12176 20080 12373 20108
rect 14660 20080 14979 20108
rect 15139 20080 15226 20108
rect 15948 20080 16528 20108
rect 17531 20080 17618 20108
rect 18708 20080 19104 20108
rect 19352 20080 21312 20108
rect 21487 20080 21574 20108
rect 15948 20040 15976 20080
rect 15764 20012 15976 20040
rect 16500 20040 16528 20080
rect 16500 20012 17371 20040
rect 13832 19944 14320 19972
rect 15856 19944 16252 19972
rect 21744 19944 21956 19972
rect 5796 19808 23000 19904
rect 10060 19740 10272 19768
rect 20180 19740 20668 19768
rect 21284 19740 21496 19768
rect 7668 19672 8156 19700
rect 10428 19672 11391 19700
rect 14231 19672 14335 19700
rect 15289 19672 15884 19700
rect 17420 19672 17985 19700
rect 7668 19632 7696 19672
rect 5920 19604 6132 19632
rect 7484 19604 7696 19632
rect 8128 19632 8156 19672
rect 8128 19604 8355 19632
rect 8588 19604 8708 19632
rect 11551 19604 11638 19632
rect 19904 19604 21772 19632
rect 14568 19536 15056 19564
rect 17623 19536 17710 19564
rect 21027 19536 21114 19564
rect 21928 19536 23060 19564
rect 21928 19496 21956 19536
rect 16960 19468 17448 19496
rect 16960 19428 16988 19468
rect 6288 19400 6408 19428
rect 7116 19400 7236 19428
rect 13115 19400 13202 19428
rect 15672 19400 16436 19428
rect 16776 19400 16988 19428
rect 17420 19428 17448 19468
rect 19260 19468 20852 19496
rect 19260 19428 19288 19468
rect 17420 19400 19288 19428
rect 20824 19428 20852 19468
rect 21284 19468 21956 19496
rect 21284 19428 21312 19468
rect 20824 19400 21312 19428
rect 23032 19428 23060 19536
rect 23032 19400 26096 19428
rect 5796 19264 23000 19360
rect 8423 19060 8510 19088
rect 12452 19060 12848 19088
rect 14955 19060 15042 19088
rect 16592 19060 17172 19088
rect 18724 19060 18814 19088
rect 20364 19060 21496 19088
rect 16592 19020 16620 19060
rect 6031 18992 6118 19020
rect 6307 18992 6408 19020
rect 8680 18992 8785 19020
rect 11808 18992 12219 19020
rect 14476 18992 14795 19020
rect 16408 18992 16620 19020
rect 17144 19020 17172 19060
rect 17144 18992 17356 19020
rect 7484 18856 7972 18884
rect 8680 18856 8708 18992
rect 13004 18924 13492 18952
rect 13004 18918 13032 18924
rect 11808 18890 13032 18918
rect 11808 18884 11836 18890
rect 9876 18856 10272 18884
rect 10704 18856 11100 18884
rect 11624 18856 11836 18884
rect 13464 18884 13492 18924
rect 17512 18924 18184 18952
rect 18708 18924 19089 18952
rect 19260 18924 20024 18952
rect 17512 18918 17540 18924
rect 16040 18890 17540 18918
rect 16040 18884 16068 18890
rect 13464 18856 13676 18884
rect 15856 18856 16068 18884
rect 18156 18884 18184 18924
rect 19260 18884 19288 18924
rect 18156 18856 18368 18884
rect 18432 18856 19288 18884
rect 19996 18884 20024 18924
rect 20364 18884 20392 19060
rect 21468 18952 21496 19060
rect 21928 18992 22523 19020
rect 22683 18992 22770 19020
rect 21468 18924 22140 18952
rect 19996 18856 20392 18884
rect 21284 18856 21404 18884
rect 5796 18720 23000 18816
rect 6012 18652 6592 18680
rect 7944 18612 7972 18680
rect 8312 18652 8708 18680
rect 13188 18652 14504 18680
rect 14752 18652 17540 18680
rect 22296 18652 22416 18680
rect 7944 18584 8156 18612
rect 8791 18584 8878 18612
rect 8975 18584 9062 18612
rect 11551 18584 11638 18612
rect 14476 18584 14504 18652
rect 16132 18612 16160 18652
rect 15304 18584 15700 18612
rect 15948 18584 16160 18612
rect 18064 18584 18460 18612
rect 18791 18594 19104 18622
rect 8128 18578 8156 18584
rect 8128 18550 8708 18578
rect 8680 18544 8708 18550
rect 7116 18516 7972 18544
rect 8680 18516 8800 18544
rect 11440 18516 11560 18544
rect 6123 18448 6210 18476
rect 6472 18448 6960 18476
rect 7760 18448 8340 18476
rect 8423 18448 8510 18476
rect 9232 18448 10272 18476
rect 6932 18408 6960 18448
rect 9232 18408 9260 18448
rect 6932 18380 7328 18408
rect 8680 18380 9260 18408
rect 10244 18408 10272 18448
rect 10244 18380 10456 18408
rect 11716 18380 11744 18544
rect 13648 18516 14228 18544
rect 14292 18516 14412 18544
rect 14568 18516 15240 18544
rect 15396 18516 15516 18544
rect 15580 18516 15884 18544
rect 16684 18516 18000 18544
rect 18083 18516 18170 18544
rect 18267 18516 18354 18544
rect 18524 18516 18828 18544
rect 19076 18516 19104 18594
rect 20916 18584 21128 18612
rect 22126 18516 22324 18544
rect 15488 18476 15516 18516
rect 14108 18448 15332 18476
rect 15488 18448 16160 18476
rect 17158 18448 17245 18476
rect 17342 18448 17429 18476
rect 21100 18448 21298 18476
rect 12747 18380 12834 18408
rect 13924 18380 14044 18408
rect 14476 18380 14964 18408
rect 15304 18340 15332 18448
rect 21967 18380 22071 18408
rect 16132 18346 17632 18374
rect 16132 18340 16160 18346
rect 6767 18312 6854 18340
rect 7208 18312 8156 18340
rect 8864 18312 8984 18340
rect 11256 18312 11560 18340
rect 11900 18312 12020 18340
rect 14568 18312 14780 18340
rect 15304 18312 15516 18340
rect 15948 18312 16160 18340
rect 17604 18340 17632 18346
rect 17604 18312 17816 18340
rect 19831 18312 19918 18340
rect 5796 18176 23000 18272
rect 6104 18108 6224 18136
rect 6840 18108 7512 18136
rect 7668 18108 8248 18136
rect 8312 18108 9720 18136
rect 10428 18108 10548 18136
rect 11348 18108 11468 18136
rect 11532 18108 13676 18136
rect 14016 18108 15700 18136
rect 18156 18108 18368 18136
rect 7484 18068 7512 18108
rect 7484 18040 7604 18068
rect 7760 17982 7788 18108
rect 8220 18068 8248 18108
rect 8220 18040 8524 18068
rect 9416 18040 9996 18068
rect 12820 18040 12940 18068
rect 9968 17972 9996 18040
rect 12728 17972 13124 18000
rect 14955 17972 15042 18000
rect 7484 17904 7788 17932
rect 8772 17904 8984 17932
rect 9048 17904 9260 17932
rect 9784 17904 10272 17932
rect 12467 17904 12940 17932
rect 13004 17904 14412 17932
rect 15856 17904 16344 17932
rect 16684 17904 16712 18068
rect 16868 18040 16988 18068
rect 22680 17972 22770 18000
rect 16960 17904 17356 17932
rect 18800 17904 18920 17932
rect 19153 17904 19380 17932
rect 13004 17864 13032 17904
rect 17328 17864 17356 17904
rect 19352 17864 19380 17904
rect 19904 17904 21128 17932
rect 19904 17864 19932 17904
rect 7223 17836 7972 17864
rect 11716 17836 13032 17864
rect 13096 17796 13124 17864
rect 13188 17836 13492 17864
rect 14568 17836 14789 17864
rect 16427 17836 16514 17864
rect 16592 17836 16804 17864
rect 6104 17768 6868 17796
rect 8588 17768 8708 17796
rect 12636 17768 13124 17796
rect 13464 17796 13492 17836
rect 17221 17796 17249 17864
rect 17328 17836 17448 17864
rect 17604 17836 18644 17864
rect 19352 17836 19932 17864
rect 22388 17836 22523 17864
rect 17604 17796 17632 17836
rect 13464 17768 13676 17796
rect 17221 17768 17632 17796
rect 18616 17796 18644 17836
rect 18616 17768 19012 17796
rect 20272 17768 20392 17796
rect 21100 17768 21404 17796
rect 5796 17632 23000 17728
rect 6932 17564 7972 17592
rect 7944 17558 7972 17564
rect 8588 17564 8800 17592
rect 8975 17564 9062 17592
rect 10336 17564 12296 17592
rect 12360 17564 12664 17592
rect 16316 17564 16528 17592
rect 17696 17564 18276 17592
rect 18340 17564 19656 17592
rect 8588 17558 8616 17564
rect 7944 17530 8616 17558
rect 7484 17496 7604 17524
rect 6472 17462 7236 17490
rect 6472 17456 6500 17462
rect 5920 17428 6500 17456
rect 7208 17456 7236 17462
rect 10336 17456 10364 17564
rect 10520 17496 10732 17524
rect 7208 17428 7604 17456
rect 7668 17428 7788 17456
rect 7929 17428 8248 17456
rect 9140 17428 9260 17456
rect 9324 17428 9812 17456
rect 10244 17428 10364 17456
rect 10428 17428 10548 17456
rect 10612 17428 11100 17456
rect 6583 17360 6670 17388
rect 6748 17360 7052 17388
rect 7222 17360 7309 17388
rect 7576 17360 7604 17428
rect 10520 17360 10548 17428
rect 11072 17388 11100 17428
rect 11532 17428 11744 17456
rect 11532 17388 11560 17428
rect 11072 17360 11560 17388
rect 12268 17388 12296 17564
rect 18248 17524 18276 17564
rect 13403 17496 13507 17524
rect 15197 17496 15976 17524
rect 18248 17496 18920 17524
rect 19260 17496 19932 17524
rect 21483 17496 21864 17524
rect 22112 17496 22232 17524
rect 18892 17456 18920 17496
rect 12912 17428 13768 17456
rect 14752 17428 14964 17456
rect 17439 17428 17526 17456
rect 17773 17428 18828 17456
rect 18892 17428 19196 17456
rect 19352 17388 19380 17456
rect 21468 17428 21772 17456
rect 12268 17360 12756 17388
rect 18892 17360 19380 17388
rect 18892 17292 18920 17360
rect 18998 17292 19085 17320
rect 22112 17252 22140 17496
rect 22204 17360 22508 17388
rect 9140 17224 9260 17252
rect 10796 17224 10916 17252
rect 20364 17224 22140 17252
rect 22204 17224 22416 17252
rect 5796 17088 23000 17184
rect 7116 17020 7880 17048
rect 7944 17020 8248 17048
rect 10520 17020 10732 17048
rect 7852 16952 7880 17020
rect 10704 16980 10732 17020
rect 11256 17020 11468 17048
rect 13648 17020 14320 17048
rect 16132 17020 16252 17048
rect 18800 17020 19840 17048
rect 11256 16980 11284 17020
rect 19812 17014 19840 17020
rect 20640 17020 20852 17048
rect 21763 17020 21850 17048
rect 22407 17020 22494 17048
rect 20640 17014 20668 17020
rect 19812 16986 20668 17014
rect 8312 16952 8708 16980
rect 8864 16952 9076 16980
rect 10704 16952 11284 16980
rect 13391 16952 13478 16980
rect 21192 16952 28580 16980
rect 21192 16912 21220 16952
rect 7024 16884 7604 16912
rect 7668 16884 8800 16912
rect 9140 16884 9260 16912
rect 12820 16884 13216 16912
rect 14955 16884 15042 16912
rect 20548 16884 21220 16912
rect 21284 16884 21404 16912
rect 21560 16884 21680 16912
rect 22131 16884 22218 16912
rect 7576 16844 7604 16884
rect 20548 16844 20576 16884
rect 6012 16816 6132 16844
rect 6656 16816 7512 16844
rect 7576 16816 7788 16844
rect 7866 16816 7953 16844
rect 8772 16816 8984 16844
rect 9769 16816 10088 16844
rect 11992 16816 12587 16844
rect 12728 16816 12940 16844
rect 13207 16816 13294 16844
rect 14476 16816 14789 16844
rect 16960 16816 17371 16844
rect 17512 16816 18828 16844
rect 19628 16816 20300 16844
rect 20364 16816 20576 16844
rect 20654 16816 20741 16844
rect 22020 16816 22232 16844
rect 22296 16816 22416 16844
rect 6273 16748 6408 16776
rect 7392 16680 7420 16816
rect 8772 16776 8800 16816
rect 22204 16776 22232 16816
rect 7576 16748 8800 16776
rect 12820 16748 13124 16776
rect 7576 16680 7604 16748
rect 13188 16708 13216 16776
rect 18892 16748 19089 16776
rect 20180 16748 20484 16776
rect 22204 16748 22508 16776
rect 7668 16680 7972 16708
rect 8956 16680 9168 16708
rect 10888 16680 11376 16708
rect 12636 16680 13216 16708
rect 20180 16680 20208 16748
rect 21744 16680 22416 16708
rect 5796 16544 23000 16640
rect 8772 16476 8984 16504
rect 20272 16476 21312 16504
rect 21836 16476 22048 16504
rect 22112 16476 22324 16504
rect 22388 16476 22600 16504
rect 8956 16436 8984 16476
rect 8956 16408 9812 16436
rect 10888 16408 11080 16436
rect 9784 16368 9812 16408
rect 22112 16368 22140 16476
rect 22388 16368 22416 16476
rect 7760 16340 7880 16368
rect 7944 16340 8141 16368
rect 9784 16340 10088 16368
rect 10796 16340 11100 16368
rect 11900 16340 12664 16368
rect 13464 16340 13967 16368
rect 14200 16340 14780 16368
rect 17439 16340 17526 16368
rect 17773 16340 18092 16368
rect 21497 16340 22140 16368
rect 22204 16340 22416 16368
rect 9140 16272 9904 16300
rect 11900 16232 11928 16340
rect 11716 16204 11928 16232
rect 12636 16232 12664 16340
rect 22112 16300 22140 16340
rect 17236 16272 17356 16300
rect 19904 16272 20470 16300
rect 22112 16272 22416 16300
rect 12636 16204 12848 16232
rect 15967 16204 16054 16232
rect 16868 16204 17172 16232
rect 20364 16204 20645 16232
rect 11716 16164 11744 16204
rect 9140 16136 9260 16164
rect 10152 16136 10272 16164
rect 10612 16136 11744 16164
rect 11992 16136 12204 16164
rect 18616 16136 18920 16164
rect 21928 16136 22048 16164
rect 5796 16000 23000 16096
rect 6380 15932 6500 15960
rect 10796 15932 12664 15960
rect 12912 15932 13676 15960
rect 14660 15932 15240 15960
rect 16224 15932 16620 15960
rect 17696 15932 17908 15960
rect 11348 15796 11560 15824
rect 14955 15796 15042 15824
rect 11532 15756 11560 15796
rect 15212 15756 15240 15932
rect 17880 15926 17908 15932
rect 18708 15932 18920 15960
rect 21284 15932 21404 15960
rect 18708 15926 18736 15932
rect 17880 15898 18736 15926
rect 15580 15864 16068 15892
rect 15580 15824 15608 15864
rect 15396 15796 15608 15824
rect 16040 15824 16068 15864
rect 16040 15796 16252 15824
rect 17972 15796 18644 15824
rect 22680 15796 22770 15824
rect 6215 15728 6302 15756
rect 7024 15728 7328 15756
rect 8220 15728 8340 15756
rect 9416 15728 9996 15756
rect 11072 15728 11468 15756
rect 11532 15728 11928 15756
rect 11900 15688 11928 15728
rect 12452 15728 12664 15756
rect 12452 15688 12480 15728
rect 9140 15660 9705 15688
rect 11701 15620 11729 15688
rect 11900 15660 12480 15688
rect 13464 15660 14789 15688
rect 15120 15620 15148 15756
rect 15212 15728 15332 15756
rect 15396 15728 15424 15796
rect 15488 15728 15884 15756
rect 16040 15728 17632 15756
rect 17788 15728 17908 15756
rect 17972 15728 18000 15796
rect 18175 15728 18262 15756
rect 19843 15728 19947 15756
rect 20107 15728 20194 15756
rect 20364 15728 21680 15756
rect 17343 15660 17908 15688
rect 18064 15660 18920 15688
rect 19076 15660 19656 15688
rect 11532 15592 11729 15620
rect 12820 15592 13124 15620
rect 15120 15592 15700 15620
rect 15764 15592 16436 15620
rect 17880 15592 17908 15660
rect 19076 15620 19104 15660
rect 19628 15654 19656 15660
rect 20364 15654 20392 15728
rect 21652 15688 21680 15728
rect 21652 15660 22324 15688
rect 22503 15660 23060 15688
rect 19628 15626 20392 15654
rect 18800 15592 19104 15620
rect 22296 15620 22324 15660
rect 22296 15592 22968 15620
rect 5796 15456 23000 15552
rect 23032 15416 23060 15660
rect 6288 15388 6500 15416
rect 6472 15382 6500 15388
rect 7484 15388 7696 15416
rect 11072 15388 13216 15416
rect 14568 15388 15148 15416
rect 7484 15382 7512 15388
rect 6472 15354 7512 15382
rect 15120 15382 15148 15388
rect 17052 15388 17264 15416
rect 18819 15388 18906 15416
rect 22480 15388 23060 15416
rect 15120 15354 15700 15382
rect 15672 15348 15700 15354
rect 17052 15348 17080 15388
rect 7944 15320 8616 15348
rect 10045 15320 10180 15348
rect 11348 15320 11928 15348
rect 12006 15320 12093 15348
rect 15672 15320 17080 15348
rect 7944 15280 7972 15320
rect 6491 15252 6578 15280
rect 7319 15252 7406 15280
rect 7760 15252 7972 15280
rect 8588 15280 8616 15320
rect 8588 15252 8815 15280
rect 8956 15252 9076 15280
rect 9711 15252 9798 15280
rect 11459 15252 11546 15280
rect 11735 15252 11822 15280
rect 12103 15252 12190 15280
rect 13004 15252 13386 15280
rect 14752 15252 14964 15280
rect 15197 15252 15516 15280
rect 17439 15252 17526 15280
rect 17604 15252 17801 15280
rect 21131 15252 21235 15280
rect 22296 15252 22508 15280
rect 6580 15184 6670 15212
rect 7760 15116 7788 15252
rect 17604 15212 17632 15252
rect 16408 15184 17632 15212
rect 21395 15184 21482 15212
rect 21928 15184 22140 15212
rect 10704 15116 13584 15144
rect 10704 15076 10732 15116
rect 13556 15110 13584 15116
rect 14108 15116 14964 15144
rect 14108 15110 14136 15116
rect 13556 15082 14136 15110
rect 14936 15076 14964 15116
rect 16224 15116 16896 15144
rect 16224 15076 16252 15116
rect 7116 15048 7328 15076
rect 10428 15048 10732 15076
rect 10888 15048 11192 15076
rect 14936 15048 16252 15076
rect 16316 15048 16436 15076
rect 19996 15048 20116 15076
rect 5796 14912 23000 15008
rect 7392 14844 7512 14872
rect 7944 14844 8340 14872
rect 10704 14844 12112 14872
rect 7871 14708 7958 14736
rect 10520 14708 10640 14736
rect 6031 14640 6118 14668
rect 7760 14640 8156 14668
rect 8791 14640 8878 14668
rect 5736 14572 6393 14600
rect 8956 14572 9153 14600
rect 5736 14328 5764 14572
rect 10152 14504 10272 14532
rect 10336 14504 10364 14668
rect 10520 14640 10548 14708
rect 10704 14640 10732 14844
rect 12084 14838 12112 14844
rect 13096 14844 13308 14872
rect 13391 14844 13478 14872
rect 13648 14844 14044 14872
rect 16408 14844 17724 14872
rect 17788 14844 18092 14872
rect 13096 14838 13124 14844
rect 12084 14810 13124 14838
rect 12820 14708 13216 14736
rect 10999 14640 11086 14668
rect 13023 14640 13110 14668
rect 13188 14640 13216 14708
rect 13280 14640 13308 14844
rect 15672 14776 16252 14804
rect 14752 14640 15056 14668
rect 10612 14532 10640 14600
rect 10900 14572 11361 14600
rect 11624 14572 13400 14600
rect 14772 14572 15240 14600
rect 15488 14532 15516 14668
rect 15672 14640 15700 14776
rect 17696 14736 17724 14844
rect 17531 14708 17618 14736
rect 17696 14708 18092 14736
rect 20104 14708 20194 14736
rect 18064 14668 18092 14708
rect 15764 14640 15884 14668
rect 17788 14640 18000 14668
rect 18064 14640 18184 14668
rect 18248 14640 18368 14668
rect 20364 14640 21220 14668
rect 22683 14640 22770 14668
rect 15580 14572 16712 14600
rect 17236 14572 17371 14600
rect 17991 14572 18078 14600
rect 19168 14572 19656 14600
rect 19843 14572 19947 14600
rect 16684 14532 16712 14572
rect 19168 14532 19196 14572
rect 10612 14504 10732 14532
rect 12379 14504 12466 14532
rect 15488 14504 15700 14532
rect 16684 14504 18828 14532
rect 18984 14504 19196 14532
rect 19628 14532 19656 14572
rect 20364 14532 20392 14640
rect 19628 14504 20392 14532
rect 21192 14532 21220 14640
rect 21928 14572 22523 14600
rect 21192 14504 22324 14532
rect 5796 14368 23000 14464
rect 23124 14328 23152 14532
rect 5736 14300 6408 14328
rect 7300 14300 7972 14328
rect 10336 14300 10916 14328
rect 10888 14260 10916 14300
rect 11348 14300 11652 14328
rect 11808 14300 12480 14328
rect 12636 14300 15700 14328
rect 16224 14300 16620 14328
rect 16979 14300 17066 14328
rect 17144 14300 17540 14328
rect 20088 14300 20300 14328
rect 11348 14260 11376 14300
rect 10045 14232 10180 14260
rect 10888 14232 11376 14260
rect 11808 14232 11836 14300
rect 16592 14260 16620 14300
rect 17144 14260 17172 14300
rect 20272 14260 20300 14300
rect 21008 14300 21772 14328
rect 22112 14300 23152 14328
rect 21008 14260 21036 14300
rect 16592 14232 17172 14260
rect 18631 14232 19012 14260
rect 20272 14232 21036 14260
rect 22112 14232 22140 14300
rect 22296 14232 22784 14260
rect 22296 14192 22324 14232
rect 6288 14164 6592 14192
rect 9784 14164 9904 14192
rect 11827 14164 11914 14192
rect 12006 14164 12093 14192
rect 13004 14164 16698 14192
rect 18819 14164 18906 14192
rect 21207 14164 21404 14192
rect 21836 14164 22324 14192
rect 22756 14192 22784 14232
rect 22756 14164 22876 14192
rect 6748 14096 7144 14124
rect 8418 14096 9168 14124
rect 21395 14096 21482 14124
rect 7208 14028 7673 14056
rect 11164 14028 12848 14056
rect 14752 14028 15976 14056
rect 22480 14028 22784 14056
rect 7944 13960 8708 13988
rect 12103 13960 12190 13988
rect 21100 13960 22140 13988
rect 5796 13824 23000 13920
rect 8036 13756 8984 13784
rect 15415 13756 15502 13784
rect 17807 13756 17894 13784
rect 21008 13756 21404 13784
rect 21468 13756 22416 13784
rect 7484 13688 7788 13716
rect 16040 13688 16252 13716
rect 20640 13688 21128 13716
rect 7668 13648 7696 13688
rect 16040 13648 16068 13688
rect 21468 13648 21496 13756
rect 21652 13688 22523 13716
rect 7668 13620 8064 13648
rect 8036 13580 8064 13620
rect 8496 13620 8708 13648
rect 12452 13620 13676 13648
rect 15856 13620 16068 13648
rect 17531 13620 17618 13648
rect 17696 13620 18460 13648
rect 8496 13580 8524 13620
rect 6031 13552 6118 13580
rect 8036 13552 8524 13580
rect 11716 13552 13124 13580
rect 13372 13552 13492 13580
rect 13556 13552 13937 13580
rect 14936 13552 15700 13580
rect 15856 13552 15884 13620
rect 17696 13580 17724 13620
rect 16132 13552 17724 13580
rect 17972 13552 18092 13580
rect 18432 13552 18460 13620
rect 21192 13620 21496 13648
rect 21192 13580 21220 13620
rect 20824 13552 21220 13580
rect 17972 13512 18000 13552
rect 6365 13484 6469 13512
rect 6748 13484 7420 13512
rect 12115 13484 12219 13512
rect 12452 13484 13216 13512
rect 13280 13484 13860 13512
rect 6748 13444 6776 13484
rect 6564 13416 6776 13444
rect 7392 13444 7420 13484
rect 13832 13444 13860 13484
rect 14108 13484 14780 13512
rect 15764 13484 16344 13512
rect 17343 13484 17724 13512
rect 17788 13484 18000 13512
rect 18083 13484 18170 13512
rect 18248 13484 18644 13512
rect 20364 13484 20576 13512
rect 14108 13444 14136 13484
rect 7392 13416 7604 13444
rect 10999 13416 11086 13444
rect 12636 13416 12848 13444
rect 13832 13416 14136 13444
rect 14752 13444 14780 13484
rect 16316 13444 16344 13484
rect 14752 13416 15056 13444
rect 16316 13416 16620 13444
rect 17696 13416 17724 13484
rect 20548 13478 20576 13484
rect 21192 13484 21404 13512
rect 21192 13478 21220 13484
rect 20548 13450 21220 13478
rect 5796 13280 23000 13376
rect 6104 13212 6592 13240
rect 6932 13212 7236 13240
rect 11164 13212 11376 13240
rect 9140 13144 9996 13172
rect 10355 13144 10442 13172
rect 9968 13104 9996 13144
rect 10962 13132 11100 13184
rect 11348 13172 11376 13212
rect 12820 13212 14780 13240
rect 12820 13172 12848 13212
rect 11348 13144 11928 13172
rect 11900 13104 11928 13144
rect 12544 13144 12848 13172
rect 12544 13104 12572 13144
rect 7469 13076 8432 13104
rect 9968 13076 10364 13104
rect 10447 13076 10534 13104
rect 10704 13076 10916 13104
rect 11900 13076 12572 13104
rect 8404 13036 8432 13076
rect 6583 13008 6670 13036
rect 6748 12900 6776 13036
rect 6932 13008 7236 13036
rect 8404 13008 10088 13036
rect 10428 12900 10456 13036
rect 10723 13008 10810 13036
rect 13924 13008 13952 13212
rect 14403 13144 14490 13172
rect 15856 13144 16077 13172
rect 16666 13135 16730 13252
rect 17144 13212 17264 13240
rect 17788 13212 18092 13240
rect 19260 13212 20116 13240
rect 21376 13212 21588 13240
rect 21928 13212 22140 13240
rect 19260 13172 19288 13212
rect 16776 13144 19288 13172
rect 20364 13144 21235 13172
rect 22480 13144 22876 13172
rect 14127 13076 14214 13104
rect 14292 13076 14412 13104
rect 14568 13076 14964 13104
rect 16040 13076 16344 13104
rect 16422 13076 16509 13104
rect 16868 13076 17080 13104
rect 17052 13036 17080 13076
rect 17604 13076 17816 13104
rect 18831 13076 18935 13104
rect 19168 13076 21496 13104
rect 21560 13076 22324 13104
rect 22572 13076 22692 13104
rect 22848 13076 22876 13144
rect 17604 13036 17632 13076
rect 14108 13008 14596 13036
rect 17052 13008 17632 13036
rect 12747 12940 12834 12968
rect 14568 12940 14596 13008
rect 21560 12900 21588 13076
rect 22480 13008 23152 13036
rect 21928 12940 23060 12968
rect 6472 12872 6776 12900
rect 9876 12872 10272 12900
rect 10428 12872 11192 12900
rect 12084 12872 12204 12900
rect 14679 12872 14766 12900
rect 14936 12872 15608 12900
rect 20272 12872 21588 12900
rect 22683 12872 22770 12900
rect 5796 12736 23000 12832
rect 8220 12668 8340 12696
rect 9048 12668 10548 12696
rect 10704 12668 10916 12696
rect 11992 12668 13400 12696
rect 13464 12668 14320 12696
rect 14568 12668 15056 12696
rect 16224 12668 18000 12696
rect 19996 12668 20300 12696
rect 21468 12668 21680 12696
rect 6856 12532 6946 12560
rect 9048 12492 9076 12668
rect 11716 12600 12112 12628
rect 15304 12600 15792 12628
rect 17623 12600 17710 12628
rect 5736 12464 6684 12492
rect 5736 12424 5764 12464
rect 4172 12396 5764 12424
rect 6656 12424 6684 12464
rect 7024 12464 7512 12492
rect 7024 12424 7052 12464
rect 7484 12424 7512 12464
rect 7944 12464 9076 12492
rect 9154 12464 9241 12492
rect 9435 12464 9522 12492
rect 10336 12464 11008 12492
rect 11072 12464 11652 12492
rect 11716 12464 11744 12600
rect 15304 12492 15332 12600
rect 15764 12560 15792 12600
rect 15764 12532 16436 12560
rect 7944 12424 7972 12464
rect 6656 12396 7052 12424
rect 7191 12356 7219 12424
rect 7484 12396 7972 12424
rect 9600 12396 9797 12424
rect 9600 12390 9628 12396
rect 9048 12362 9628 12390
rect 9048 12356 9076 12362
rect 11808 12356 11836 12492
rect 12084 12464 12204 12492
rect 12345 12464 12664 12492
rect 13575 12464 13662 12492
rect 15212 12464 15332 12492
rect 15410 12464 15497 12492
rect 15580 12464 15700 12492
rect 17052 12464 17632 12492
rect 17807 12464 17894 12492
rect 17972 12464 18000 12668
rect 18156 12600 18828 12628
rect 20272 12560 20300 12668
rect 22020 12600 22523 12628
rect 20107 12532 20194 12560
rect 20272 12532 21758 12560
rect 18175 12464 18262 12492
rect 13909 12396 14596 12424
rect 15488 12396 15976 12424
rect 16132 12396 16896 12424
rect 17343 12396 18000 12424
rect 18064 12396 18736 12424
rect 19843 12396 19947 12424
rect 16132 12356 16160 12396
rect 7191 12328 7328 12356
rect 8864 12328 9076 12356
rect 11532 12328 11836 12356
rect 15856 12328 16160 12356
rect 16868 12356 16896 12396
rect 16868 12328 17632 12356
rect 17972 12328 18000 12396
rect 5796 12192 23000 12288
rect 11164 12124 11376 12152
rect 11440 12124 11560 12152
rect 18708 12124 18920 12152
rect 21100 12124 21680 12152
rect 9048 12056 10073 12084
rect 15856 12056 16077 12084
rect 17604 12056 17801 12084
rect 6288 11988 6408 12016
rect 7871 11988 7958 12016
rect 8205 11988 8524 12016
rect 9048 11988 9076 12056
rect 21652 12016 21680 12124
rect 22480 12124 22784 12152
rect 22480 12016 22508 12124
rect 9784 11988 9904 12016
rect 11256 11988 11928 12016
rect 12931 11988 13018 12016
rect 16040 11988 17540 12016
rect 21207 11988 21588 12016
rect 21652 11988 21864 12016
rect 22204 11988 22508 12016
rect 22591 11988 22678 12016
rect 16592 11920 17080 11948
rect 21395 11920 21482 11948
rect 22480 11920 22784 11948
rect 17052 11880 17080 11920
rect 13280 11852 13400 11880
rect 16316 11852 16436 11880
rect 16795 11852 16882 11880
rect 17052 11852 17540 11880
rect 5736 11784 6132 11812
rect 6491 11784 6578 11812
rect 8864 11784 9352 11812
rect 14752 11784 14964 11812
rect 16132 11784 16804 11812
rect 17163 11784 17250 11812
rect 20088 11784 22416 11812
rect 5736 11608 5764 11784
rect 5796 11648 23000 11744
rect 5736 11580 6040 11608
rect 8496 11580 8892 11608
rect 11072 11580 11284 11608
rect 12360 11580 12756 11608
rect 14568 11580 15516 11608
rect 15672 11580 15792 11608
rect 19996 11580 20208 11608
rect 12728 11540 12756 11580
rect 12728 11512 12848 11540
rect 20180 11472 20208 11580
rect 21100 11580 22784 11608
rect 21100 11472 21128 11580
rect 6104 11444 6500 11472
rect 7484 11444 8524 11472
rect 19003 11444 19090 11472
rect 20180 11444 21128 11472
rect 21303 11444 21390 11472
rect 6196 11268 6224 11404
rect 6564 11376 6761 11404
rect 8680 11376 9260 11404
rect 10796 11376 10916 11404
rect 12636 11376 12756 11404
rect 12931 11376 13018 11404
rect 13372 11376 13676 11404
rect 14384 11376 15148 11404
rect 15488 11376 15608 11404
rect 17052 11376 17632 11404
rect 6932 11308 7696 11336
rect 10428 11308 10563 11336
rect 12467 11308 13216 11336
rect 13909 11308 14504 11336
rect 14752 11308 15332 11336
rect 6932 11268 6960 11308
rect 5736 11240 6224 11268
rect 6472 11240 6960 11268
rect 7668 11268 7696 11308
rect 15396 11268 15424 11336
rect 16500 11308 17371 11336
rect 19337 11308 19932 11336
rect 21560 11308 21665 11336
rect 21560 11268 21588 11308
rect 7668 11240 7880 11268
rect 9048 11240 9444 11268
rect 15396 11240 16252 11268
rect 20383 11240 20470 11268
rect 21008 11240 21588 11268
rect 5736 11064 5764 11240
rect 5796 11104 23000 11200
rect 5736 11036 7144 11064
rect 7392 11036 7512 11064
rect 14108 11036 14504 11064
rect 17052 11036 17908 11064
rect 17972 11036 18920 11064
rect 19260 11036 19932 11064
rect 21928 11036 23244 11064
rect 6399 10968 6486 10996
rect 10355 10968 10442 10996
rect 12176 10968 12296 10996
rect 13495 10968 13584 10996
rect 17052 10928 17080 11036
rect 17236 10968 17801 10996
rect 17880 10928 17908 11036
rect 21928 10928 21956 11036
rect 22034 10968 22121 10996
rect 22388 10968 22508 10996
rect 6012 10900 6132 10928
rect 8602 10900 8708 10928
rect 9968 10900 10902 10928
rect 13832 10900 17080 10928
rect 17512 10900 17632 10928
rect 17880 10900 18644 10928
rect 6104 10860 6132 10900
rect 18616 10860 18644 10900
rect 19260 10900 20300 10928
rect 21758 10900 21956 10928
rect 19260 10860 19288 10900
rect 22112 10860 22140 10928
rect 22204 10900 22784 10928
rect 6104 10832 6776 10860
rect 8510 10832 8892 10860
rect 9232 10832 10272 10860
rect 13667 10832 13754 10860
rect 18616 10832 19288 10860
rect 20456 10832 20746 10860
rect 22112 10832 22692 10860
rect 7737 10764 7972 10792
rect 9987 10764 10074 10792
rect 11663 10764 11767 10792
rect 14476 10764 14780 10792
rect 20893 10764 21312 10792
rect 10888 10730 11560 10758
rect 10888 10724 10916 10730
rect 8772 10696 8984 10724
rect 10704 10696 10916 10724
rect 11532 10724 11560 10730
rect 11532 10696 12204 10724
rect 12287 10696 12374 10724
rect 21284 10696 21312 10764
rect 22388 10696 22508 10724
rect 5796 10560 23000 10656
rect 8680 10492 9168 10520
rect 8680 10384 8708 10492
rect 9140 10486 9168 10492
rect 9784 10492 10088 10520
rect 13556 10492 14044 10520
rect 9784 10486 9812 10492
rect 9140 10458 9812 10486
rect 8883 10424 8984 10452
rect 9968 10424 10180 10452
rect 8588 10356 8708 10384
rect 10152 10384 10180 10424
rect 11440 10424 11744 10452
rect 13299 10424 13386 10452
rect 11440 10384 11468 10424
rect 10152 10356 11468 10384
rect 13004 10356 13676 10384
rect 13759 10356 13846 10384
rect 17604 10356 17724 10384
rect 18064 10356 18276 10384
rect 18524 10356 18644 10384
rect 6123 10288 6210 10316
rect 14587 10288 14674 10316
rect 14921 10288 15148 10316
rect 15120 10248 15148 10288
rect 15672 10288 16068 10316
rect 16132 10288 16528 10316
rect 17880 10288 18460 10316
rect 18800 10288 19104 10316
rect 21376 10288 21496 10316
rect 21579 10288 21680 10316
rect 15672 10248 15700 10288
rect 6288 10220 6485 10248
rect 15120 10220 15700 10248
rect 17343 10220 17724 10248
rect 18984 10220 19084 10248
rect 6288 10214 6316 10220
rect 5736 10186 6316 10214
rect 5736 9976 5764 10186
rect 18984 10180 19012 10220
rect 7576 10152 7696 10180
rect 16224 10152 16988 10180
rect 18248 10152 19012 10180
rect 19904 10152 20208 10180
rect 5796 10016 23000 10112
rect 5736 9948 6408 9976
rect 9784 9948 10180 9976
rect 10152 9908 10180 9948
rect 11440 9948 11652 9976
rect 12360 9948 12572 9976
rect 15875 9948 15962 9976
rect 16684 9948 17540 9976
rect 19352 9948 19932 9976
rect 21652 9948 22140 9976
rect 11440 9942 11468 9948
rect 10612 9914 11468 9942
rect 10612 9908 10640 9914
rect 19352 9908 19380 9948
rect 10152 9880 10640 9908
rect 12912 9880 13507 9908
rect 16960 9880 17089 9908
rect 18631 9880 19380 9908
rect 19444 9880 20377 9908
rect 20548 9880 21128 9908
rect 20548 9840 20576 9880
rect 6380 9812 7328 9840
rect 7668 9812 7866 9840
rect 10827 9812 10931 9840
rect 12636 9812 13768 9840
rect 17328 9812 18920 9840
rect 20015 9812 20102 9840
rect 20180 9812 20576 9840
rect 21100 9840 21128 9880
rect 21744 9846 22692 9874
rect 21744 9840 21772 9846
rect 21100 9812 21772 9840
rect 22664 9840 22692 9846
rect 22664 9812 22876 9840
rect 20180 9772 20208 9812
rect 7576 9744 7751 9772
rect 11091 9744 11178 9772
rect 14200 9744 15976 9772
rect 19628 9744 19748 9772
rect 19812 9744 20208 9772
rect 21836 9744 22324 9772
rect 22407 9744 22494 9772
rect 22296 9704 22324 9744
rect 7116 9676 7949 9704
rect 14016 9676 14320 9704
rect 18892 9636 18920 9704
rect 22296 9676 22784 9704
rect 19076 9642 20024 9670
rect 19076 9636 19104 9642
rect 8956 9608 9076 9636
rect 14384 9608 14504 9636
rect 18892 9608 19104 9636
rect 19996 9636 20024 9642
rect 19996 9608 21496 9636
rect 5796 9472 23000 9568
rect 6932 9404 7604 9432
rect 9048 9404 9168 9432
rect 10815 9404 10902 9432
rect 19720 9404 20300 9432
rect 20916 9404 21128 9432
rect 21284 9404 21496 9432
rect 22112 9404 22531 9432
rect 19076 9370 19564 9398
rect 19076 9364 19104 9370
rect 8588 9336 8708 9364
rect 16408 9336 16689 9364
rect 18156 9336 19104 9364
rect 19536 9364 19564 9370
rect 19536 9336 19955 9364
rect 18156 9296 18184 9336
rect 7300 9268 9444 9296
rect 10355 9268 10442 9296
rect 10520 9268 10640 9296
rect 16243 9268 16330 9296
rect 17788 9268 18184 9296
rect 20180 9296 20208 9404
rect 20548 9336 20944 9364
rect 20916 9330 20944 9336
rect 21560 9336 22232 9364
rect 21560 9330 21588 9336
rect 20916 9302 21588 9330
rect 20180 9268 20760 9296
rect 22296 9282 22324 9364
rect 22503 9336 22531 9404
rect 6123 9200 6210 9228
rect 9416 9160 9444 9268
rect 9968 9200 10824 9228
rect 12011 9200 12098 9228
rect 13372 9200 14412 9228
rect 14476 9200 14673 9228
rect 16132 9200 16606 9228
rect 18156 9200 19090 9228
rect 22586 9200 23060 9228
rect 9968 9160 9996 9200
rect 6457 9132 6776 9160
rect 8128 9132 8800 9160
rect 9416 9132 9996 9160
rect 10167 9132 10364 9160
rect 8128 9092 8156 9132
rect 7944 9064 8156 9092
rect 8772 9092 8800 9132
rect 10336 9126 10364 9132
rect 11072 9132 11284 9160
rect 12287 9132 12388 9160
rect 11072 9126 11100 9132
rect 10336 9098 11100 9126
rect 8772 9064 8984 9092
rect 13391 9064 13478 9092
rect 15691 9064 15778 9092
rect 18156 9064 18184 9200
rect 18248 9092 18276 9160
rect 18340 9132 18828 9160
rect 18248 9064 20300 9092
rect 22204 9064 22876 9092
rect 5796 8928 23000 9024
rect 10796 8860 11192 8888
rect 11256 8860 11468 8888
rect 12452 8860 13032 8888
rect 14752 8860 15056 8888
rect 18524 8860 18736 8888
rect 7469 8792 7972 8820
rect 9232 8724 10059 8752
rect 11164 8684 11192 8860
rect 18708 8854 18736 8860
rect 19628 8860 20208 8888
rect 22388 8860 22600 8888
rect 19628 8854 19656 8860
rect 18708 8826 19656 8854
rect 22388 8820 22416 8860
rect 11348 8792 11928 8820
rect 16408 8792 16528 8820
rect 22112 8792 22416 8820
rect 19812 8758 20300 8786
rect 19812 8752 19840 8758
rect 14752 8724 15318 8752
rect 17957 8724 18552 8752
rect 19076 8724 19840 8752
rect 20272 8752 20300 8758
rect 22112 8752 22140 8792
rect 23032 8752 23060 9200
rect 20272 8724 20470 8752
rect 21928 8724 22140 8752
rect 22223 8724 22310 8752
rect 22480 8724 23060 8752
rect 22480 8684 22508 8724
rect 7135 8656 7222 8684
rect 11164 8656 12020 8684
rect 17623 8656 17710 8684
rect 19904 8656 20363 8684
rect 22112 8656 22508 8684
rect 8588 8588 8892 8616
rect 10244 8588 10939 8616
rect 12176 8588 12825 8616
rect 14292 8588 15056 8616
rect 14292 8548 14320 8588
rect 9876 8520 10456 8548
rect 14108 8520 14320 8548
rect 15028 8548 15056 8588
rect 15373 8548 15401 8616
rect 20272 8588 20553 8616
rect 21652 8588 21772 8616
rect 21928 8554 22876 8582
rect 21928 8548 21956 8554
rect 15028 8520 15401 8548
rect 21560 8520 21956 8548
rect 22848 8548 22876 8554
rect 22848 8520 23060 8548
rect 5796 8384 23000 8480
rect 9968 8316 10272 8344
rect 13832 8316 14320 8344
rect 21468 8316 22140 8344
rect 8933 8248 9076 8276
rect 13832 8208 13860 8316
rect 23032 8276 23060 8520
rect 14085 8248 14412 8276
rect 15856 8248 15976 8276
rect 20732 8248 21680 8276
rect 22503 8248 23060 8276
rect 15856 8208 15884 8248
rect 8515 8180 8602 8208
rect 8680 8180 8771 8208
rect 12747 8180 12834 8208
rect 13740 8180 13860 8208
rect 15599 8180 15686 8208
rect 15764 8180 15884 8208
rect 21468 8180 21758 8208
rect 22867 8180 22954 8208
rect 8680 8140 8708 8180
rect 7411 8112 7498 8140
rect 7852 8112 8708 8140
rect 15212 8112 15516 8140
rect 15764 8072 15792 8180
rect 16500 8112 18920 8140
rect 20456 8112 20944 8140
rect 21652 8072 21680 8126
rect 7024 8044 7245 8072
rect 15764 8044 16620 8072
rect 17052 8044 17249 8072
rect 19153 8044 19932 8072
rect 20640 8044 21680 8072
rect 15764 8038 15792 8044
rect 12268 8010 13952 8038
rect 12268 8004 12296 8010
rect 6031 7976 6118 8004
rect 7871 7976 7958 8004
rect 12084 7976 12296 8004
rect 13924 8004 13952 8010
rect 15028 8010 15792 8038
rect 15028 8004 15056 8010
rect 16592 8004 16620 8044
rect 20640 8004 20668 8044
rect 13924 7976 15056 8004
rect 15967 7976 16054 8004
rect 16592 7976 17908 8004
rect 18340 7976 18828 8004
rect 20272 7976 20668 8004
rect 21008 7976 21128 8004
rect 5796 7840 23000 7936
rect 6472 7772 7052 7800
rect 7852 7772 8616 7800
rect 12287 7772 12374 7800
rect 18524 7772 19012 7800
rect 19444 7772 19932 7800
rect 22296 7772 22508 7800
rect 10539 7704 10626 7732
rect 14311 7704 14398 7732
rect 16040 7704 16267 7732
rect 17880 7704 18184 7732
rect 18156 7664 18184 7704
rect 7135 7636 7222 7664
rect 7300 7636 7497 7664
rect 10520 7636 10732 7664
rect 12268 7636 12572 7664
rect 16427 7636 16514 7664
rect 17512 7636 17632 7664
rect 17773 7636 18092 7664
rect 18156 7636 18552 7664
rect 18819 7636 20944 7664
rect 21008 7636 21205 7664
rect 10704 7596 10732 7636
rect 18524 7596 18552 7636
rect 6215 7568 6302 7596
rect 10704 7568 10902 7596
rect 11822 7568 12020 7596
rect 12728 7568 12848 7596
rect 12912 7568 13110 7596
rect 18524 7568 20484 7596
rect 10520 7500 11077 7528
rect 12084 7500 12664 7528
rect 12636 7494 12664 7500
rect 13096 7500 13285 7528
rect 19352 7500 19748 7528
rect 19812 7500 19932 7528
rect 13096 7494 13124 7500
rect 12636 7466 13124 7494
rect 19720 7460 19748 7500
rect 5736 7432 6040 7460
rect 10336 7432 10456 7460
rect 15120 7432 15884 7460
rect 18156 7432 18920 7460
rect 19720 7432 20116 7460
rect 5736 7256 5764 7432
rect 5796 7296 23000 7392
rect 5736 7228 6408 7256
rect 6748 7228 6960 7256
rect 7227 7228 7314 7256
rect 12452 7228 12756 7256
rect 16960 7228 17724 7256
rect 17991 7228 18078 7256
rect 18524 7228 18920 7256
rect 20199 7228 20286 7256
rect 17696 7188 17724 7228
rect 12747 7160 12834 7188
rect 17531 7160 17618 7188
rect 17696 7160 18000 7188
rect 18340 7160 19265 7188
rect 6012 7092 6132 7120
rect 6491 7092 6578 7120
rect 7668 7092 7880 7120
rect 8423 7092 8510 7120
rect 13372 7092 13676 7120
rect 15120 7092 15516 7120
rect 17623 7092 17710 7120
rect 6012 7024 6224 7052
rect 6288 7024 7788 7052
rect 8699 7024 8800 7052
rect 10796 7024 11100 7052
rect 11333 7024 11652 7052
rect 12471 7024 12940 7052
rect 13096 7024 13937 7052
rect 15212 7024 15332 7052
rect 16224 7024 16528 7052
rect 17807 7024 17894 7052
rect 6012 6916 6040 7024
rect 17972 6984 18000 7160
rect 18708 7092 19090 7120
rect 20732 7092 21312 7120
rect 18267 7024 18354 7052
rect 18524 7024 18644 7052
rect 18892 7024 19167 7052
rect 12820 6956 13032 6984
rect 16408 6956 16508 6984
rect 17972 6956 18276 6984
rect 18524 6956 18552 7024
rect 16408 6916 16436 6956
rect 18248 6916 18276 6956
rect 5736 6888 6040 6916
rect 9876 6888 9996 6916
rect 12636 6888 13308 6916
rect 13372 6888 14320 6916
rect 14752 6888 15056 6916
rect 15764 6888 16436 6916
rect 17328 6888 18184 6916
rect 18248 6888 18920 6916
rect 20272 6888 20576 6916
rect 5736 6644 5764 6888
rect 5796 6752 23000 6848
rect 6491 6684 6578 6712
rect 7760 6684 8340 6712
rect 9600 6684 9812 6712
rect 11992 6684 12204 6712
rect 12471 6684 12558 6712
rect 12747 6684 12834 6712
rect 14292 6684 14780 6712
rect 15028 6684 15700 6712
rect 16960 6684 17080 6712
rect 17604 6684 17724 6712
rect 19812 6684 20300 6712
rect 8312 6644 8340 6684
rect 9784 6678 9812 6684
rect 9784 6650 11284 6678
rect 11256 6644 11284 6650
rect 5736 6616 7236 6644
rect 8312 6616 8493 6644
rect 11256 6616 12296 6644
rect 12728 6576 12756 6644
rect 13280 6616 13661 6644
rect 18892 6616 19288 6644
rect 19812 6576 19840 6684
rect 6031 6548 6118 6576
rect 6675 6548 6776 6576
rect 7024 6548 7328 6576
rect 7852 6548 7972 6576
rect 8036 6548 8156 6576
rect 8234 6548 8321 6576
rect 10263 6548 10350 6576
rect 10428 6548 10548 6576
rect 10723 6548 10810 6576
rect 10999 6548 11100 6576
rect 12636 6548 12756 6576
rect 13299 6548 13386 6576
rect 17144 6548 17724 6576
rect 19371 6548 19458 6576
rect 19647 6548 19840 6576
rect 6748 6440 6776 6548
rect 13096 6480 13216 6508
rect 14752 6480 15226 6508
rect 16500 6480 16712 6508
rect 17255 6480 17342 6508
rect 17604 6480 17787 6508
rect 20272 6480 22140 6508
rect 16684 6440 16712 6480
rect 6748 6412 7696 6440
rect 7852 6412 8064 6440
rect 12268 6412 12388 6440
rect 15323 6412 15424 6440
rect 16684 6412 17172 6440
rect 12268 6372 12296 6412
rect 17144 6406 17172 6412
rect 17788 6412 17977 6440
rect 19352 6412 19564 6440
rect 19831 6412 19918 6440
rect 17788 6406 17816 6412
rect 17144 6378 17816 6406
rect 20272 6372 20300 6480
rect 5755 6344 5842 6372
rect 6859 6344 6946 6372
rect 10520 6344 12296 6372
rect 18524 6344 19012 6372
rect 19628 6344 20300 6372
rect 22112 6372 22140 6480
rect 22296 6372 22324 6440
rect 22112 6344 22324 6372
rect 5796 6208 23000 6304
rect 6380 6140 6960 6168
rect 6932 6100 6960 6140
rect 7944 6140 8156 6168
rect 8496 6140 8800 6168
rect 11072 6140 11376 6168
rect 11624 6140 11836 6168
rect 12655 6140 12742 6168
rect 12931 6140 13018 6168
rect 15396 6140 15516 6168
rect 18156 6140 18920 6168
rect 19168 6140 19472 6168
rect 19555 6140 19642 6168
rect 7944 6100 7972 6140
rect 20088 6100 20116 6168
rect 6932 6072 7972 6100
rect 9416 6072 10088 6100
rect 11992 6072 12848 6100
rect 14384 6072 14780 6100
rect 19536 6072 20116 6100
rect 8312 6004 8892 6032
rect 10336 5964 10364 6032
rect 10796 6004 11744 6032
rect 11992 5964 12020 6072
rect 12820 6032 12848 6072
rect 12176 6004 12388 6032
rect 12820 6004 13216 6032
rect 14403 6004 14596 6032
rect 6472 5936 6960 5964
rect 7852 5936 7972 5964
rect 9232 5936 9904 5964
rect 10336 5936 10548 5964
rect 10612 5936 10732 5964
rect 11532 5936 12020 5964
rect 12471 5936 12558 5964
rect 12636 5936 12848 5964
rect 14200 5936 14412 5964
rect 14568 5936 14596 6004
rect 14752 5936 14780 6072
rect 18340 6038 18828 6066
rect 18340 6032 18368 6038
rect 9876 5896 9904 5936
rect 10704 5896 10732 5936
rect 12636 5896 12664 5936
rect 6104 5868 6316 5896
rect 8312 5868 9076 5896
rect 9876 5868 10456 5896
rect 10704 5868 11468 5896
rect 8312 5828 8340 5868
rect 7944 5800 8340 5828
rect 9048 5828 9076 5868
rect 11440 5862 11468 5868
rect 12452 5868 12664 5896
rect 14384 5896 14412 5936
rect 15580 5896 15608 6032
rect 17604 5964 17632 6032
rect 17788 6004 18368 6032
rect 18800 6032 18828 6038
rect 18800 6004 19012 6032
rect 15672 5936 17632 5964
rect 18432 5936 18552 5964
rect 19352 5936 19656 5964
rect 19720 5936 19840 5964
rect 14384 5868 15608 5896
rect 12452 5862 12480 5868
rect 11440 5834 12480 5862
rect 9048 5800 9628 5828
rect 17880 5800 18368 5828
rect 5796 5664 23000 5760
<< metal2 >>
rect 216 24474 244 24548
rect 12268 24120 12296 24528
rect 12268 24092 12388 24120
rect 7668 21536 7696 21740
rect 7576 21508 7696 21536
rect 6564 20652 6592 21196
rect 7576 20720 7604 21508
rect 7852 20828 7880 21808
rect 9140 21644 9260 21672
rect 7576 20692 7696 20720
rect 5920 19428 5948 20652
rect 6564 20624 6684 20652
rect 5828 19400 5948 19428
rect 5828 17660 5856 19400
rect 5828 17632 5948 17660
rect 5920 17252 5948 17632
rect 5828 17224 5948 17252
rect 5828 16708 5856 17224
rect 6104 16816 6132 20108
rect 6380 20080 6408 20516
rect 6656 19972 6684 20624
rect 6564 19944 6684 19972
rect 6564 19564 6592 19944
rect 7668 19768 7696 20692
rect 7944 20624 7972 21060
rect 8680 20856 8708 21060
rect 8588 20828 8708 20856
rect 8036 20284 8064 20652
rect 8588 20624 8616 20828
rect 7668 19740 7972 19768
rect 6564 19536 6684 19564
rect 6380 18992 6408 19428
rect 6656 18884 6684 19536
rect 6564 18856 6684 18884
rect 6564 18652 6592 18856
rect 7116 18516 7144 19428
rect 6196 18108 6224 18476
rect 6840 18108 6868 18340
rect 7208 18136 7236 18340
rect 7484 18204 7512 19632
rect 7116 18108 7236 18136
rect 7392 18176 7512 18204
rect 6656 16816 6684 17388
rect 6840 16912 6868 17796
rect 7116 17660 7144 18108
rect 7392 17728 7420 18176
rect 7576 18108 7696 18136
rect 7392 17700 7512 17728
rect 7116 17632 7236 17660
rect 7024 17184 7052 17388
rect 7208 17360 7236 17632
rect 7484 17496 7512 17700
rect 7024 17156 7144 17184
rect 7116 17020 7144 17156
rect 7576 16912 7604 18108
rect 6840 16884 7052 16912
rect 7576 16884 7696 16912
rect 5828 16680 5948 16708
rect 5920 15960 5948 16680
rect 5920 15932 6316 15960
rect 6380 15932 6408 16776
rect 4172 3170 4200 12424
rect 6104 11444 6132 14668
rect 6288 14164 6316 15932
rect 7024 15552 7052 15756
rect 6656 15524 7052 15552
rect 6564 15252 6592 15398
rect 6656 15184 6684 15524
rect 7116 14096 7144 15076
rect 7392 14844 7420 16708
rect 7760 15248 7788 19668
rect 7944 19632 7972 19740
rect 7944 19604 8064 19632
rect 8036 19088 8064 19604
rect 8680 19088 8708 19668
rect 7944 19060 8064 19088
rect 8496 19060 8708 19088
rect 7944 18652 7972 19060
rect 8680 18652 8708 18884
rect 8864 18584 8892 21264
rect 9140 20992 9168 21644
rect 9968 21304 9996 21604
rect 10060 21536 10088 21740
rect 10060 21508 10272 21536
rect 9140 20964 9260 20992
rect 9232 20624 9260 20964
rect 9876 20692 9904 21196
rect 10244 20856 10272 21508
rect 11532 21060 11560 21254
rect 10060 20828 10272 20856
rect 9048 20080 9076 20516
rect 7944 18340 7972 18544
rect 7944 18312 8064 18340
rect 8036 17864 8064 18312
rect 8312 18108 8340 18476
rect 8496 18040 8524 18476
rect 8864 18136 8892 18340
rect 8864 18108 8938 18136
rect 7944 17836 8064 17864
rect 7852 16816 7880 16980
rect 7944 16680 7972 17836
rect 8220 17020 8248 17456
rect 8680 16952 8708 17796
rect 8772 17564 8800 17932
rect 8910 17456 8938 18108
rect 9048 17564 9076 18612
rect 9140 18136 9168 20312
rect 10060 19020 10088 20828
rect 10520 20760 10548 21060
rect 11348 21032 11560 21060
rect 10244 19640 10272 20652
rect 10428 19672 10456 20516
rect 11348 19496 11376 21032
rect 11624 20828 11652 21740
rect 11808 20828 11836 21808
rect 12084 21304 12112 21604
rect 11992 20760 12020 21060
rect 12176 20624 12204 21196
rect 11808 20244 11836 20516
rect 11808 20216 11928 20244
rect 11624 19604 11652 20108
rect 11348 19468 11652 19496
rect 9968 18992 10088 19020
rect 9968 18408 9996 18992
rect 9968 18380 10088 18408
rect 9140 18108 9260 18136
rect 8864 17428 8938 17456
rect 9232 17428 9260 18108
rect 9784 17428 9812 17932
rect 8864 16952 8892 17428
rect 8772 16476 8800 16912
rect 9140 16884 9168 17252
rect 9508 16884 9996 16912
rect 6380 13376 6408 13512
rect 6288 13348 6408 13376
rect 6104 10656 6132 10860
rect 5920 10628 6132 10656
rect 6288 10656 6316 13348
rect 6564 13212 6592 13444
rect 7208 13212 7236 14056
rect 7576 13104 7604 14192
rect 7760 13688 7788 15144
rect 7944 14844 7972 16368
rect 9140 16272 9168 16708
rect 8312 15690 8340 15764
rect 8864 15144 8892 15276
rect 8956 15144 8984 15280
rect 8864 15116 8984 15144
rect 7944 14300 7972 14736
rect 8864 14640 8892 15116
rect 6656 13008 6684 13080
rect 7576 13076 7696 13104
rect 6472 12696 6500 12900
rect 6472 12668 6592 12696
rect 6564 12016 6592 12668
rect 6472 11988 6592 12016
rect 6472 10968 6500 11988
rect 6932 11954 6960 13036
rect 7300 12277 7328 12356
rect 6564 11376 6592 11812
rect 6288 10628 6500 10656
rect 5920 8344 5948 10628
rect 5920 8316 6132 8344
rect 5828 6220 5856 6372
rect 6104 5868 6132 8316
rect 6196 8172 6224 10316
rect 6472 10044 6500 10628
rect 6380 10016 6500 10044
rect 6380 9812 6408 10016
rect 7116 9676 7144 11064
rect 7484 11036 7512 11472
rect 6748 8956 6776 9160
rect 6656 8928 6776 8956
rect 6656 8276 6684 8928
rect 6564 8248 6684 8276
rect 6288 6508 6316 7596
rect 6564 7460 6592 8248
rect 6932 8208 6960 9432
rect 7300 9268 7328 9840
rect 7668 9812 7696 13076
rect 7944 12152 7972 13988
rect 8956 13756 8984 14600
rect 9140 14096 9168 16164
rect 9784 15248 9812 15280
rect 9968 14192 9996 16884
rect 10060 16816 10088 18380
rect 10244 17904 10272 18884
rect 10428 18108 10456 18408
rect 10704 17496 10732 18884
rect 11624 18584 11652 19468
rect 11900 19224 11928 20216
rect 12176 20080 12204 20516
rect 12360 20448 12388 24092
rect 13188 21876 13216 27598
rect 13096 21848 13216 21876
rect 13096 21264 13124 21848
rect 16408 21740 16436 27598
rect 13372 21372 13400 21740
rect 13096 21236 13216 21264
rect 12636 20556 12664 21060
rect 12360 20420 12572 20448
rect 12544 19564 12572 20420
rect 12820 19640 12848 20652
rect 12544 19536 12664 19564
rect 12636 19224 12664 19536
rect 11808 19196 11928 19224
rect 12544 19196 12664 19224
rect 11808 18992 11836 19196
rect 11440 18108 11468 18544
rect 11532 17564 11560 18340
rect 10520 17020 10548 17388
rect 10888 16408 10916 17252
rect 10152 14638 10180 16164
rect 10428 14532 10456 15076
rect 10612 14708 10640 16164
rect 9876 14164 9996 14192
rect 8220 12668 8248 13104
rect 7944 12124 8064 12152
rect 7944 11954 7972 12016
rect 8036 11880 8064 12124
rect 7944 11852 8064 11880
rect 7944 10764 7972 11852
rect 8496 11580 8524 12016
rect 8680 11376 8708 13648
rect 9140 12464 9168 13172
rect 9508 12413 9536 12492
rect 8680 10248 8708 10928
rect 8864 10832 8892 12356
rect 9968 12016 9996 14164
rect 10152 13052 10180 14532
rect 10336 12464 10364 14532
rect 10428 14504 10548 14532
rect 10520 13376 10548 14504
rect 10428 13348 10548 13376
rect 10428 13144 10456 13348
rect 10520 12668 10548 13104
rect 10704 12668 10732 14532
rect 10888 13052 10916 15076
rect 11072 14640 11100 16368
rect 10796 12442 10824 13036
rect 8956 10424 8984 10724
rect 9048 10356 9076 12016
rect 9876 11988 9996 12016
rect 10980 12016 11008 13172
rect 11072 12464 11100 13444
rect 11164 13212 11192 14666
rect 11348 14124 11376 16708
rect 11532 15252 11560 15620
rect 11716 15552 11744 18408
rect 11992 16816 12020 18340
rect 12544 18000 12572 19196
rect 12544 17972 12664 18000
rect 12636 17564 12664 17972
rect 12820 17456 12848 19088
rect 13188 18652 13216 21236
rect 12912 17904 12940 18068
rect 12820 17428 12940 17456
rect 11716 15524 11836 15552
rect 11808 14872 11836 15524
rect 11992 15320 12020 16164
rect 12268 15552 12296 17388
rect 12728 16816 12756 17388
rect 12636 15932 12664 16708
rect 12820 15960 12848 16776
rect 12820 15932 12940 15960
rect 12176 15524 12296 15552
rect 11808 14844 12020 14872
rect 11624 14300 11652 14600
rect 11992 14328 12020 14844
rect 12176 14572 12204 15524
rect 11716 14300 12020 14328
rect 12452 14300 12480 14532
rect 12636 14300 12664 15756
rect 11348 14096 11468 14124
rect 11164 12124 11192 12900
rect 11440 12560 11468 14096
rect 11348 12532 11468 12560
rect 10980 11988 11100 12016
rect 9232 10832 9260 11404
rect 10888 11376 10916 11982
rect 10428 10968 10456 11336
rect 8680 10220 8892 10248
rect 7576 9404 7604 9772
rect 7944 8792 7972 9092
rect 8680 8888 8708 9364
rect 8588 8860 8708 8888
rect 6840 8180 6960 8208
rect 6840 7664 6868 8180
rect 7024 7772 7052 8072
rect 6840 7636 6960 7664
rect 7208 7636 7236 8684
rect 7484 8112 7512 8200
rect 8588 8180 8616 8860
rect 7852 7772 7880 8140
rect 6564 7432 6776 7460
rect 6748 7228 6776 7432
rect 6564 6684 6592 7120
rect 6288 6480 6408 6508
rect 6380 5760 6408 6480
rect 6748 6140 6776 6576
rect 6932 5936 6960 7636
rect 7300 7228 7328 7664
rect 7760 6684 7788 7052
rect 7852 6412 7880 7120
rect 7944 5936 7972 8004
rect 8680 7120 8708 8200
rect 8864 8112 8892 10220
rect 9048 8248 9076 9636
rect 9140 9432 9168 10316
rect 9968 9948 9996 10928
rect 10244 10810 10272 10884
rect 11072 10832 11100 11988
rect 10060 10492 10088 10792
rect 9140 9404 9260 9432
rect 10888 9404 10916 9840
rect 9232 8724 9260 9404
rect 9968 9268 10456 9296
rect 9968 8172 9996 9268
rect 10152 8072 10180 8684
rect 10244 8316 10272 8616
rect 8496 7092 8708 7120
rect 8128 5800 8156 6576
rect 8220 6548 8248 6614
rect 8312 6004 8340 6712
rect 8680 6586 8708 7092
rect 9968 8044 10180 8072
rect 8772 6140 8800 7052
rect 9968 6072 9996 8044
rect 10428 7800 10456 8548
rect 10428 7772 10548 7800
rect 10520 7500 10548 7772
rect 10612 7704 10640 9296
rect 10796 8860 10824 9228
rect 11164 9148 11192 9772
rect 11348 9392 11376 12532
rect 11532 12124 11560 12356
rect 11716 12328 11744 14300
rect 11900 11988 11928 14192
rect 11992 14164 12020 14300
rect 12820 14028 12848 14736
rect 12176 13484 12204 13988
rect 12084 12600 12112 12900
rect 12176 12464 12204 12714
rect 12268 11580 12388 11608
rect 12268 10968 12296 11580
rect 12452 11336 12480 13512
rect 12636 12464 12664 13444
rect 12636 11376 12664 11982
rect 12452 11308 12572 11336
rect 11716 10424 11744 10792
rect 12176 10520 12204 10724
rect 12084 10492 12204 10520
rect 11256 8860 11284 9160
rect 11440 8684 11468 8932
rect 11348 8656 11468 8684
rect 8864 5976 8892 6032
rect 10336 6004 10364 7460
rect 10428 5868 10456 6576
rect 10796 6548 10824 8200
rect 11348 7528 11376 8656
rect 11624 7636 11652 9976
rect 12084 9636 12112 10492
rect 12360 9704 12388 10724
rect 12544 9948 12572 11308
rect 12820 9840 12848 12968
rect 13004 11988 13032 18544
rect 13096 17972 13216 18000
rect 13096 14638 13124 15620
rect 13188 13648 13216 17972
rect 13464 17496 13492 21196
rect 14292 20788 14320 21196
rect 14200 20760 14320 20788
rect 14200 20176 14228 20760
rect 14384 20624 14412 21060
rect 14200 20148 14320 20176
rect 14292 19672 14320 20148
rect 14476 18992 14504 20856
rect 14660 20080 14688 20516
rect 15212 20080 15240 20156
rect 15488 20148 15516 21740
rect 16408 21712 16528 21740
rect 15672 20216 15700 21060
rect 15856 19672 15884 21128
rect 16224 20760 16252 21604
rect 15948 20128 15976 20720
rect 16500 20652 16528 21712
rect 16960 21372 16988 21672
rect 16408 20624 16528 20652
rect 14752 19088 14780 19564
rect 14752 19060 15056 19088
rect 14752 18908 14780 19060
rect 13648 18054 13676 18544
rect 14016 18108 14044 18408
rect 14292 18340 14320 18544
rect 14200 18312 14320 18340
rect 14384 18516 14596 18544
rect 14200 17864 14228 18312
rect 14384 17904 14412 18516
rect 14200 17836 14320 17864
rect 14292 17020 14320 17836
rect 13280 16788 13308 16862
rect 13464 16340 13492 16980
rect 14476 16816 14504 18408
rect 14568 17836 14596 18340
rect 14752 18000 14780 18680
rect 15672 18584 15700 19428
rect 16408 19400 16436 20624
rect 17420 19672 17448 21196
rect 18248 20284 18276 21264
rect 19076 21236 19104 21740
rect 18800 20760 18828 21060
rect 17604 20080 17632 20156
rect 18524 20128 18552 20652
rect 15212 18496 15240 18570
rect 15488 18068 15516 18340
rect 15396 18040 15516 18068
rect 14752 17972 15056 18000
rect 14752 16912 14780 17972
rect 15396 17320 15424 18040
rect 15396 17292 15516 17320
rect 15488 16980 15516 17292
rect 15396 16952 15516 16980
rect 15672 16956 15700 18136
rect 14752 16884 15056 16912
rect 14292 15932 14688 15960
rect 13464 14844 13492 15688
rect 14292 15416 14320 15932
rect 14016 15388 14320 15416
rect 14752 15824 14780 16368
rect 15396 16232 15424 16952
rect 15856 16776 15884 18884
rect 15948 17496 15976 18340
rect 16132 17020 16160 18476
rect 15672 16748 15884 16776
rect 15396 16204 15516 16232
rect 14752 15796 15056 15824
rect 14016 14844 14044 15388
rect 14752 14640 14780 15796
rect 15488 15416 15516 16204
rect 15672 15416 15700 16748
rect 15488 15388 15608 15416
rect 15672 15388 15746 15416
rect 15488 14804 15516 15280
rect 15396 14776 15516 14804
rect 15396 14668 15424 14776
rect 15304 14640 15424 14668
rect 13188 13620 13308 13648
rect 13188 12686 13216 13620
rect 13372 13540 13400 14600
rect 13556 13444 13584 13580
rect 13464 13416 13584 13444
rect 13464 13376 13492 13416
rect 13372 13348 13492 13376
rect 13372 12668 13400 13348
rect 14292 13240 14320 13568
rect 14200 13212 14320 13240
rect 14200 13104 14228 13212
rect 14108 13076 14228 13104
rect 13648 12413 13676 12492
rect 14108 12424 14136 13076
rect 14292 12668 14320 13104
rect 14476 12696 14504 13172
rect 14568 12940 14596 14328
rect 15304 14192 15332 14640
rect 15580 14300 15608 15388
rect 15718 14872 15746 15388
rect 15718 14844 15792 14872
rect 15764 14640 15792 14844
rect 15672 14464 15700 14532
rect 15856 14464 15884 15756
rect 15672 14436 15884 14464
rect 15304 14164 15424 14192
rect 15396 14056 15424 14164
rect 14752 13212 14780 14056
rect 15396 14028 15516 14056
rect 15488 13756 15516 14028
rect 14936 13076 14964 13580
rect 14476 12668 14596 12696
rect 14108 12396 14412 12424
rect 14384 12084 14412 12396
rect 14292 12056 14412 12084
rect 13188 11852 13308 11880
rect 13004 10856 13032 11404
rect 12636 9812 12848 9840
rect 12912 9704 12940 9908
rect 12360 9676 12940 9704
rect 12084 9608 12204 9636
rect 12084 9148 12112 9228
rect 11992 8480 12020 8684
rect 12176 8588 12204 9608
rect 11992 8452 12112 8480
rect 12084 7664 12112 8452
rect 12360 7772 12388 9160
rect 12636 8656 12664 9676
rect 12820 8172 12848 9176
rect 13004 8860 13032 10384
rect 13188 8112 13216 11852
rect 14292 11608 14320 12056
rect 14292 11580 14412 11608
rect 14568 11580 14596 12424
rect 14752 12076 14780 12900
rect 15580 12696 15608 12900
rect 15396 12668 15608 12696
rect 15396 12464 15424 12668
rect 12084 7636 12296 7664
rect 11348 7500 11468 7528
rect 11440 7188 11468 7500
rect 11348 7160 11468 7188
rect 10612 5936 10640 6372
rect 11072 6140 11100 6576
rect 11348 5828 11376 7160
rect 11624 6140 11652 7052
rect 11992 6684 12020 7596
rect 12268 6616 12296 7636
rect 12912 7392 12940 7596
rect 12728 7364 12940 7392
rect 11532 5936 11560 6004
rect 12544 5936 12572 7052
rect 12728 6140 12756 7364
rect 12820 6684 12848 7188
rect 13004 6906 13032 6984
rect 13096 6576 13124 7052
rect 13004 6548 13124 6576
rect 13004 6140 13032 6548
rect 13188 6004 13216 6614
rect 13372 6548 13400 11404
rect 14384 11376 14412 11580
rect 14476 11036 14504 11336
rect 14752 11308 14780 11812
rect 13556 10492 13584 10996
rect 13740 10246 13768 10860
rect 13832 10356 13860 10928
rect 14660 10246 14688 10316
rect 13464 8548 13492 9092
rect 13464 8520 13584 8548
rect 13556 8072 13584 8520
rect 14292 8316 14320 9704
rect 14476 9200 14504 9636
rect 14752 8860 14780 10792
rect 14200 8180 14320 8208
rect 13464 8044 13584 8072
rect 13464 7636 13492 8044
rect 14292 6684 14320 8180
rect 14384 7704 14412 8276
rect 14752 8112 14780 8752
rect 15488 8656 15516 11608
rect 15580 11376 15608 12492
rect 15672 12464 15700 14436
rect 15764 13982 15792 14042
rect 15856 12424 15884 13172
rect 15764 12396 15884 12424
rect 15764 11580 15792 12396
rect 15856 12030 15884 12104
rect 15948 11404 15976 12424
rect 16040 11988 16068 16252
rect 16224 14300 16252 15824
rect 16316 15736 16344 18544
rect 16684 18040 16712 18570
rect 16500 17564 16528 17864
rect 16776 17836 16804 19428
rect 16960 17660 16988 18068
rect 16868 17632 16988 17660
rect 16868 17048 16896 17632
rect 16868 17020 16988 17048
rect 16960 16816 16988 17020
rect 17144 16504 17172 18476
rect 17328 16776 17356 19020
rect 17696 18908 17724 19564
rect 18708 18924 18736 20516
rect 19904 20284 19932 21264
rect 20088 20312 20116 21672
rect 20272 20760 20300 21604
rect 20088 20284 20208 20312
rect 20180 19740 20208 20284
rect 20364 20128 20392 20720
rect 21284 19740 21312 20108
rect 17512 17864 17540 18680
rect 17696 18340 17724 18544
rect 17696 18312 17816 18340
rect 17420 17836 17540 17864
rect 16868 16476 17172 16504
rect 17236 16748 17356 16776
rect 16408 15184 16436 15620
rect 16592 15144 16620 15960
rect 16592 15116 16712 15144
rect 16868 15116 16896 16476
rect 17236 15388 17264 16748
rect 17512 15252 17540 17836
rect 17788 17796 17816 18312
rect 18156 18108 18184 18544
rect 17696 17768 17816 17796
rect 17696 17320 17724 17768
rect 17696 17292 17816 17320
rect 16408 14844 16436 15076
rect 16408 12532 16436 13580
rect 16592 13036 16620 13444
rect 16684 13212 16712 15116
rect 16592 13008 16712 13036
rect 16684 12424 16712 13008
rect 16592 12396 16712 12424
rect 15856 11376 15976 11404
rect 15856 10724 15884 11376
rect 15764 10696 15884 10724
rect 15764 10180 15792 10696
rect 16132 10656 16160 11812
rect 16040 10628 16160 10656
rect 16040 10288 16068 10628
rect 15764 10152 15976 10180
rect 15948 9948 15976 10152
rect 16316 10112 16344 11880
rect 16592 11472 16620 12396
rect 16592 11444 16712 11472
rect 16224 10084 16344 10112
rect 15764 8752 15792 9092
rect 15672 8724 15792 8752
rect 15948 8248 15976 9772
rect 16224 9500 16252 10084
rect 16224 9472 16344 9500
rect 16316 9268 16344 9472
rect 16132 8208 16160 9228
rect 16408 8792 16436 9364
rect 16500 9268 16528 11336
rect 16684 9948 16712 11444
rect 16868 10316 16896 11880
rect 16822 10288 16896 10316
rect 16822 9772 16850 10288
rect 16960 9880 16988 10180
rect 17052 10112 17080 14328
rect 17236 13212 17264 14600
rect 17236 10968 17264 11812
rect 17052 10084 17264 10112
rect 17236 9840 17264 10084
rect 17236 9812 17356 9840
rect 16822 9744 16896 9772
rect 15488 7256 15516 8140
rect 15396 7228 15516 7256
rect 14476 6004 14504 6980
rect 14752 6072 14780 6916
rect 15212 6586 15240 7052
rect 15396 6412 15424 7228
rect 15488 6140 15516 7120
rect 15672 6684 15700 8208
rect 15856 8180 16160 8208
rect 15856 7256 15884 8180
rect 16040 7704 16068 8004
rect 15856 7228 15976 7256
rect 15948 6780 15976 7228
rect 16500 7024 16528 8140
rect 16868 7256 16896 9744
rect 17052 7868 17080 8072
rect 17052 7840 17172 7868
rect 16868 7228 16988 7256
rect 17144 7120 17172 7840
rect 17052 7092 17172 7120
rect 15856 6752 15976 6780
rect 15856 6548 15884 6752
rect 17052 6684 17080 7092
rect 17420 7074 17448 14328
rect 17604 13620 17632 15756
rect 17696 12600 17724 13444
rect 17788 13418 17816 17292
rect 18340 16776 18368 18884
rect 18432 18584 18460 18884
rect 18800 17904 18828 19088
rect 19076 18496 19104 18570
rect 19904 18542 19932 19632
rect 21100 18584 21128 19564
rect 18800 17020 18828 17456
rect 18984 17292 19012 17796
rect 19168 16834 19196 17456
rect 19628 16816 19656 17592
rect 19904 17444 19932 18340
rect 21100 18272 21128 18476
rect 21284 18272 21312 18884
rect 21100 18244 21312 18272
rect 21100 17904 21128 18244
rect 20364 16816 20392 17796
rect 21100 16980 21128 17796
rect 21008 16952 21128 16980
rect 20640 16788 20668 16862
rect 18248 16748 18368 16776
rect 18248 16504 18276 16748
rect 18248 16476 18368 16504
rect 17880 15416 17908 15620
rect 17880 15388 17954 15416
rect 17926 13988 17954 15388
rect 18064 14844 18092 16368
rect 18340 15960 18368 16476
rect 18248 15932 18368 15960
rect 18248 15552 18276 15932
rect 18248 15524 18368 15552
rect 18340 14872 18368 15524
rect 18248 14844 18368 14872
rect 17880 13960 17954 13988
rect 17880 13756 17908 13960
rect 17880 13104 17908 13512
rect 18064 13212 18092 14600
rect 18248 14464 18276 14844
rect 18248 14436 18368 14464
rect 18340 13852 18368 14436
rect 18248 13824 18368 13852
rect 17788 13076 17908 13104
rect 17880 12464 17908 13076
rect 18156 12600 18184 13512
rect 18248 13444 18276 13824
rect 18616 13484 18644 16164
rect 18892 15932 18920 16776
rect 21008 16504 21036 16952
rect 21008 16476 21128 16504
rect 21284 16476 21312 16912
rect 19904 15728 19932 16300
rect 21100 16272 21128 16476
rect 20364 15892 20392 16232
rect 21284 15932 21312 16368
rect 20364 15864 20484 15892
rect 18892 15388 18920 15688
rect 19996 14600 20024 15076
rect 19904 14572 20024 14600
rect 18984 14232 19012 14532
rect 19996 14260 20024 14572
rect 19904 14232 20024 14260
rect 18892 14150 18920 14192
rect 19904 13512 19932 14232
rect 19904 13484 20024 13512
rect 18248 13416 18368 13444
rect 18340 13308 18368 13416
rect 18340 13280 18460 13308
rect 18432 12696 18460 13280
rect 18248 12668 18460 12696
rect 18248 12464 18276 12668
rect 17604 12056 17632 12356
rect 17512 11852 17632 11880
rect 17604 11744 17632 11852
rect 17604 11716 17724 11744
rect 17696 11268 17724 11716
rect 17604 11240 17724 11268
rect 17604 11036 17632 11240
rect 17972 11036 18000 12356
rect 18708 12124 18736 12424
rect 17604 10900 17724 10928
rect 17696 7664 17724 10900
rect 17880 10288 17908 10996
rect 18248 9132 18276 10384
rect 18156 8888 18184 9092
rect 18064 8860 18184 8888
rect 18064 8208 18092 8860
rect 18064 8180 18184 8208
rect 17604 7636 17724 7664
rect 17328 6480 17356 6916
rect 17604 6004 17632 7188
rect 17696 6684 17724 7120
rect 17880 6576 17908 8004
rect 18064 7228 18092 7664
rect 17696 6548 17908 6576
rect 18156 6548 18184 8180
rect 18340 7160 18368 9160
rect 18524 8860 18552 10384
rect 18708 9500 18736 11064
rect 18892 9676 18920 13104
rect 19996 12668 20024 13484
rect 20180 12532 20208 15756
rect 20456 15144 20484 15864
rect 20364 15116 20484 15144
rect 20364 14804 20392 15116
rect 20364 14776 20484 14804
rect 20456 14056 20484 14776
rect 20364 14028 20484 14056
rect 21192 14056 21220 15280
rect 21192 14028 21312 14056
rect 20364 13484 20392 14028
rect 21100 13688 21128 13988
rect 19904 11744 19932 12424
rect 19904 11716 20024 11744
rect 19996 11580 20024 11716
rect 19076 10246 19104 11494
rect 19904 11036 19932 11336
rect 20272 10384 20300 12900
rect 20364 12628 20392 13172
rect 20364 12600 20484 12628
rect 20456 12492 20484 12600
rect 20456 12464 20576 12492
rect 20548 12016 20576 12464
rect 21100 12124 21128 13580
rect 21284 13240 21312 14028
rect 21376 13756 21404 14192
rect 21284 13212 21404 13240
rect 20456 11988 20576 12016
rect 20456 11880 20484 11988
rect 20364 11852 20484 11880
rect 20364 11608 20392 11852
rect 20364 11580 20484 11608
rect 20456 10832 20484 11580
rect 21376 11336 21404 11472
rect 21468 11336 21496 20156
rect 21560 19904 21588 21740
rect 21560 19876 21680 19904
rect 21652 18816 21680 19876
rect 21744 19604 21772 20516
rect 21928 18992 21956 19972
rect 22112 18924 22140 20888
rect 22296 19972 22324 20176
rect 22296 19944 22416 19972
rect 22388 18884 22416 19944
rect 26068 19400 26096 24304
rect 22296 18856 22416 18884
rect 21652 18788 21772 18816
rect 21744 17728 21772 18788
rect 22296 18652 22324 18856
rect 21652 17700 21772 17728
rect 21652 14736 21680 17700
rect 21836 17020 21864 17524
rect 22020 16476 22048 18408
rect 22296 18272 22324 18544
rect 22204 18244 22324 18272
rect 22204 17496 22232 18244
rect 22388 17660 22416 17864
rect 22342 17632 22416 17660
rect 22204 16884 22232 17252
rect 22342 17048 22370 17632
rect 22480 17048 22508 17388
rect 22342 17020 22416 17048
rect 22480 17020 22600 17048
rect 22296 16476 22324 16844
rect 22388 16680 22416 17020
rect 21928 15184 21956 16164
rect 21652 14708 22140 14736
rect 21744 13784 21772 14328
rect 21744 13756 21864 13784
rect 21652 12668 21680 13716
rect 21836 13552 21864 13756
rect 21928 13212 21956 14600
rect 22112 13076 22140 14708
rect 22296 13648 22324 14532
rect 22480 13784 22508 16776
rect 22572 16476 22600 17020
rect 22756 14638 22784 19020
rect 22940 15416 22968 15620
rect 22940 15388 23060 15416
rect 23032 14532 23060 15388
rect 22940 14504 23060 14532
rect 22940 14192 22968 14504
rect 22940 14164 23060 14192
rect 22388 13756 22508 13784
rect 22296 13620 22416 13648
rect 22480 12968 22508 13172
rect 22388 12940 22508 12968
rect 22388 12832 22416 12940
rect 22296 12804 22416 12832
rect 21652 11784 21680 12492
rect 21376 11308 21496 11336
rect 21008 10724 21036 11268
rect 21008 10696 21128 10724
rect 21100 10452 21128 10696
rect 21008 10424 21128 10452
rect 20272 10356 20392 10384
rect 18708 9472 18828 9500
rect 18524 7772 18552 8752
rect 18800 8480 18828 9472
rect 19168 9268 19196 9908
rect 19720 9404 19748 9772
rect 18708 8452 18828 8480
rect 18708 8344 18736 8452
rect 18662 8316 18736 8344
rect 18662 7324 18690 8316
rect 18800 7528 18828 8004
rect 18892 7636 18920 8322
rect 19076 7732 19104 8752
rect 19904 8656 19932 10180
rect 20088 9812 20116 10274
rect 20364 9704 20392 10356
rect 20272 9676 20392 9704
rect 21008 9704 21036 10424
rect 21008 9676 21128 9704
rect 20272 9404 20300 9676
rect 21100 9404 21128 9676
rect 21284 9404 21312 10724
rect 21468 10288 21496 11308
rect 21836 10452 21864 12016
rect 22020 10968 22048 12628
rect 22296 12152 22324 12804
rect 22572 12464 22600 13104
rect 22296 12124 22508 12152
rect 22756 12124 22784 14056
rect 22296 10792 22324 11608
rect 22480 10968 22508 12124
rect 23032 12016 23060 14164
rect 28552 13906 28580 16980
rect 22204 10764 22324 10792
rect 21836 10424 21956 10452
rect 21652 9948 21680 10316
rect 21928 9976 21956 10424
rect 21836 9948 21956 9976
rect 21836 9744 21864 9948
rect 22204 9636 22232 10764
rect 22480 9744 22508 10724
rect 22664 9704 22692 12016
rect 22940 11988 23060 12016
rect 22940 10490 22968 11988
rect 22848 9812 22968 9840
rect 22940 9704 22968 9812
rect 22572 9676 22692 9704
rect 20272 8344 20300 8616
rect 20180 8316 20300 8344
rect 19904 7772 19932 8072
rect 19076 7704 19196 7732
rect 18800 7500 18920 7528
rect 18662 7296 18736 7324
rect 18708 7092 18736 7296
rect 11348 5800 11468 5828
rect 18340 5800 18368 7052
rect 18524 5936 18552 6984
rect 18892 6140 18920 7500
rect 19168 6984 19196 7704
rect 20180 7664 20208 8316
rect 20180 7636 20300 7664
rect 19076 6956 19196 6984
rect 19076 6712 19104 6956
rect 19076 6684 19472 6712
rect 19352 5936 19380 6440
rect 19444 6140 19472 6684
rect 19628 6140 19656 6372
rect 19720 5936 19748 6576
rect 19904 6412 19932 7528
rect 20088 6140 20116 7460
rect 20272 7228 20300 7636
rect 20456 7568 20484 8200
rect 21468 8180 21496 9636
rect 22204 9608 22324 9636
rect 22112 9228 22140 9432
rect 22020 9200 22140 9228
rect 21652 8248 21680 8616
rect 22020 8548 22048 9200
rect 22204 9064 22232 9364
rect 22296 9336 22324 9608
rect 22572 8860 22600 9676
rect 22020 8520 22140 8548
rect 22112 8316 22140 8520
rect 22296 8140 22324 8752
rect 22204 8112 22324 8140
rect 21008 7636 21036 8004
rect 21284 7092 21312 8072
rect 22204 7664 22232 8112
rect 22480 7772 22508 8752
rect 22756 8172 22784 9704
rect 22940 9676 23060 9704
rect 23032 8412 23060 9676
rect 22940 8384 23060 8412
rect 22940 8180 22968 8384
rect 22204 7636 22324 7664
rect 20272 6684 20300 6916
rect 22296 6412 22324 7636
rect 6288 5732 6408 5760
rect 6288 120 6316 5732
rect 11440 3856 11468 5800
rect 11440 3828 11560 3856
rect 11532 3658 11560 3828
<< metal3 >>
rect 0 27676 4860 27736
rect 4800 27614 4860 27676
rect 22648 27676 28796 27736
rect 22648 27614 22708 27676
rect 4800 27554 13232 27614
rect 16392 27554 22708 27614
rect 0 24504 260 24564
rect 26052 24260 28796 24320
rect 0 21454 5780 21514
rect 5720 21270 5780 21454
rect 5720 21210 11576 21270
rect 22096 20844 28796 20904
rect 15196 20112 21512 20172
rect 7744 19624 12864 19684
rect 12804 18892 18844 18952
rect 15196 18526 16728 18586
rect 19060 18526 19948 18586
rect 0 18404 10748 18464
rect 13632 18038 15900 18098
rect 19888 17428 28796 17488
rect 15653 16937 15816 17003
rect 6088 16818 7804 16878
rect 11700 16818 13324 16878
rect 19152 16818 20684 16878
rect 14736 16208 16084 16268
rect 8296 15720 16360 15780
rect 0 15354 6608 15414
rect 7744 15232 12910 15292
rect 10136 14622 11208 14682
rect 13080 14622 13324 14682
rect 21452 14622 22800 14682
rect 17036 14134 20224 14194
rect 15656 14012 15778 14072
rect 28536 13890 28796 13950
rect 13356 13524 14336 13584
rect 15656 13402 17832 13462
rect 6640 13036 10196 13096
rect 10872 13036 11254 13096
rect 12160 12670 13232 12730
rect 9492 12426 13692 12486
rect 0 12304 4768 12364
rect 6778 12304 7344 12364
rect 14736 12060 15900 12120
rect 6088 11938 12910 11998
rect 19060 11450 21512 11510
rect 10228 10840 13876 10900
rect 22924 10474 28796 10534
rect 13356 10230 20132 10290
rect 16944 9864 19212 9924
rect 11056 9376 11392 9436
rect 11056 9314 11116 9376
rect 0 9254 11116 9314
rect 11148 9132 12864 9192
rect 11194 8888 11484 8948
rect 17680 8278 18936 8338
rect 6180 8156 12910 8216
rect 20440 8156 22800 8216
rect 17404 7058 28796 7118
rect 12988 6936 14520 6996
rect 8204 6570 8724 6630
rect 13172 6570 15256 6630
rect 0 6204 5872 6264
rect 8848 5960 11576 6020
rect 11516 3642 28796 3702
rect 0 3154 4216 3214
rect 13264 164 13324 286
rect 0 104 6332 164
rect 13264 104 28796 164
<< metal4 >>
rect 3936 0 4556 27744
rect 4708 12304 4906 12364
rect 5176 0 5796 27744
rect 6640 12304 6838 12364
rect 8000 3852 8620 23892
rect 9240 5092 9860 22652
rect 11194 8888 11254 13096
rect 12850 8156 12910 15292
rect 13264 7850 13324 14682
rect 13126 7790 13324 7850
rect 13126 3702 13186 7790
rect 13600 3852 14220 23892
rect 14840 5092 15460 22652
rect 15748 16634 15808 17000
rect 15748 16574 15946 16634
rect 15886 14438 15946 16574
rect 15748 14378 15946 14438
rect 15748 14012 15808 14378
rect 19200 3852 19820 23892
rect 20440 5092 21060 22652
rect 13126 3642 13324 3702
rect 13264 226 13324 3642
rect 23000 0 23620 27744
rect 24240 0 24860 27744
<< metal5 >>
rect 0 23272 28796 23892
rect 0 22032 28796 22652
rect 4716 12174 6830 12494
rect 0 5092 28796 5712
rect 0 3852 28796 4472
use L1M1_PR  L1M1_PR_0
timestamp 1654583406
transform 1 0 13662 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1
timestamp 1654583406
transform 1 0 13110 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2
timestamp 1654583406
transform 1 0 12834 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3
timestamp 1654583406
transform 1 0 10534 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_4
timestamp 1654583406
transform 1 0 12466 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_5
timestamp 1654583406
transform 1 0 11822 0 1 14246
box -29 -23 29 23
use L1M1_PR  L1M1_PR_6
timestamp 1654583406
transform 1 0 11638 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_7
timestamp 1654583406
transform 1 0 11086 0 1 13430
box -29 -23 29 23
use L1M1_PR  L1M1_PR_8
timestamp 1654583406
transform 1 0 15042 0 1 13430
box -29 -23 29 23
use L1M1_PR  L1M1_PR_9
timestamp 1654583406
transform 1 0 13294 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_10
timestamp 1654583406
transform 1 0 14398 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_11
timestamp 1654583406
transform 1 0 13478 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_12
timestamp 1654583406
transform 1 0 15318 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_13
timestamp 1654583406
transform 1 0 14950 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_14
timestamp 1654583406
transform 1 0 15410 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_15
timestamp 1654583406
transform 1 0 14950 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_16
timestamp 1654583406
transform 1 0 18906 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_17
timestamp 1654583406
transform 1 0 18078 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_18
timestamp 1654583406
transform 1 0 16238 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_19
timestamp 1654583406
transform 1 0 15870 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_20
timestamp 1654583406
transform 1 0 18170 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_21
timestamp 1654583406
transform 1 0 16330 0 1 15062
box -29 -23 29 23
use L1M1_PR  L1M1_PR_22
timestamp 1654583406
transform 1 0 18906 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_23
timestamp 1654583406
transform 1 0 18262 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_24
timestamp 1654583406
transform 1 0 16698 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_25
timestamp 1654583406
transform 1 0 16238 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_26
timestamp 1654583406
transform 1 0 16238 0 1 14790
box -29 -23 29 23
use L1M1_PR  L1M1_PR_27
timestamp 1654583406
transform 1 0 15686 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_28
timestamp 1654583406
transform 1 0 15318 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_29
timestamp 1654583406
transform 1 0 13662 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_30
timestamp 1654583406
transform 1 0 18906 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_31
timestamp 1654583406
transform 1 0 18078 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_32
timestamp 1654583406
transform 1 0 20470 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_33
timestamp 1654583406
transform 1 0 20194 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_34
timestamp 1654583406
transform 1 0 19366 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_35
timestamp 1654583406
transform 1 0 18906 0 1 17306
box -29 -23 29 23
use L1M1_PR  L1M1_PR_36
timestamp 1654583406
transform 1 0 18354 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_37
timestamp 1654583406
transform 1 0 18170 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_38
timestamp 1654583406
transform 1 0 16514 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_39
timestamp 1654583406
transform 1 0 16330 0 1 17578
box -29 -23 29 23
use L1M1_PR  L1M1_PR_40
timestamp 1654583406
transform 1 0 16238 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_41
timestamp 1654583406
transform 1 0 15410 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_42
timestamp 1654583406
transform 1 0 14398 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_43
timestamp 1654583406
transform 1 0 13662 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_44
timestamp 1654583406
transform 1 0 13662 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_45
timestamp 1654583406
transform 1 0 13202 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_46
timestamp 1654583406
transform 1 0 11546 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_47
timestamp 1654583406
transform 1 0 11362 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_48
timestamp 1654583406
transform 1 0 11454 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_49
timestamp 1654583406
transform 1 0 10442 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_50
timestamp 1654583406
transform 1 0 12190 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_51
timestamp 1654583406
transform 1 0 12006 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_52
timestamp 1654583406
transform 1 0 10074 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_53
timestamp 1654583406
transform 1 0 8326 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_54
timestamp 1654583406
transform 1 0 7483 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_55
timestamp 1654583406
transform 1 0 20654 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_56
timestamp 1654583406
transform 1 0 19182 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_57
timestamp 1654583406
transform 1 0 18078 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_58
timestamp 1654583406
transform 1 0 17986 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_59
timestamp 1654583406
transform 1 0 17986 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_60
timestamp 1654583406
transform 1 0 17894 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_61
timestamp 1654583406
transform 1 0 17894 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_62
timestamp 1654583406
transform 1 0 16882 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_63
timestamp 1654583406
transform 1 0 16698 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_64
timestamp 1654583406
transform 1 0 15686 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_65
timestamp 1654583406
transform 1 0 15594 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_66
timestamp 1654583406
transform 1 0 15502 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_67
timestamp 1654583406
transform 1 0 15502 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_68
timestamp 1654583406
transform 1 0 15502 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_69
timestamp 1654583406
transform 1 0 15226 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_70
timestamp 1654583406
transform 1 0 14582 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_71
timestamp 1654583406
transform 1 0 14582 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_72
timestamp 1654583406
transform 1 0 13294 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_73
timestamp 1654583406
transform 1 0 13294 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_74
timestamp 1654583406
transform 1 0 13110 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_75
timestamp 1654583406
transform 1 0 13018 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_76
timestamp 1654583406
transform 1 0 12006 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_77
timestamp 1654583406
transform 1 0 11822 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_78
timestamp 1654583406
transform 1 0 11822 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_79
timestamp 1654583406
transform 1 0 11730 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_80
timestamp 1654583406
transform 1 0 11454 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_81
timestamp 1654583406
transform 1 0 10718 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_82
timestamp 1654583406
transform 1 0 10626 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_83
timestamp 1654583406
transform 1 0 20286 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_84
timestamp 1654583406
transform 1 0 19642 0 1 17578
box -29 -23 29 23
use L1M1_PR  L1M1_PR_85
timestamp 1654583406
transform 1 0 18446 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_86
timestamp 1654583406
transform 1 0 18354 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_87
timestamp 1654583406
transform 1 0 18354 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_88
timestamp 1654583406
transform 1 0 18262 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_89
timestamp 1654583406
transform 1 0 18262 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_90
timestamp 1654583406
transform 1 0 16422 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_91
timestamp 1654583406
transform 1 0 16330 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_92
timestamp 1654583406
transform 1 0 16146 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_93
timestamp 1654583406
transform 1 0 15870 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_94
timestamp 1654583406
transform 1 0 15594 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_95
timestamp 1654583406
transform 1 0 15226 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_96
timestamp 1654583406
transform 1 0 15134 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_97
timestamp 1654583406
transform 1 0 15134 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_98
timestamp 1654583406
transform 1 0 14214 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_99
timestamp 1654583406
transform 1 0 14214 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_100
timestamp 1654583406
transform 1 0 13478 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_101
timestamp 1654583406
transform 1 0 13478 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_102
timestamp 1654583406
transform 1 0 12926 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_103
timestamp 1654583406
transform 1 0 12834 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_104
timestamp 1654583406
transform 1 0 12190 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_105
timestamp 1654583406
transform 1 0 11546 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_106
timestamp 1654583406
transform 1 0 11270 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_107
timestamp 1654583406
transform 1 0 10994 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_108
timestamp 1654583406
transform 1 0 10350 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_109
timestamp 1654583406
transform 1 0 10258 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_110
timestamp 1654583406
transform 1 0 9982 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_111
timestamp 1654583406
transform 1 0 9154 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_112
timestamp 1654583406
transform 1 0 10258 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_113
timestamp 1654583406
transform 1 0 9890 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_114
timestamp 1654583406
transform 1 0 11362 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_115
timestamp 1654583406
transform 1 0 10626 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_116
timestamp 1654583406
transform 1 0 10442 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_117
timestamp 1654583406
transform 1 0 17342 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_118
timestamp 1654583406
transform 1 0 17342 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_119
timestamp 1654583406
transform 1 0 16422 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_120
timestamp 1654583406
transform 1 0 14582 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_121
timestamp 1654583406
transform 1 0 11715 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_122
timestamp 1654583406
transform 1 0 11546 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_123
timestamp 1654583406
transform 1 0 11066 0 1 16431
box -29 -23 29 23
use L1M1_PR  L1M1_PR_124
timestamp 1654583406
transform 1 0 10810 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_125
timestamp 1654583406
transform 1 0 12573 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_126
timestamp 1654583406
transform 1 0 11914 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_127
timestamp 1654583406
transform 1 0 12834 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_128
timestamp 1654583406
transform 1 0 12481 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_129
timestamp 1654583406
transform 1 0 14775 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_130
timestamp 1654583406
transform 1 0 14766 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_131
timestamp 1654583406
transform 1 0 14950 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_132
timestamp 1654583406
transform 1 0 14775 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_133
timestamp 1654583406
transform 1 0 17357 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_134
timestamp 1654583406
transform 1 0 16882 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_135
timestamp 1654583406
transform 1 0 17802 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_136
timestamp 1654583406
transform 1 0 15211 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_137
timestamp 1654583406
transform 1 0 18998 0 1 17306
box -29 -23 29 23
use L1M1_PR  L1M1_PR_138
timestamp 1654583406
transform 1 0 17235 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_139
timestamp 1654583406
transform 1 0 20838 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_140
timestamp 1654583406
transform 1 0 17787 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_141
timestamp 1654583406
transform 1 0 19075 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_142
timestamp 1654583406
transform 1 0 17710 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_143
timestamp 1654583406
transform 1 0 17787 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_144
timestamp 1654583406
transform 1 0 15778 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_145
timestamp 1654583406
transform 1 0 15226 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_146
timestamp 1654583406
transform 1 0 14786 0 1 14577
box -29 -23 29 23
use L1M1_PR  L1M1_PR_147
timestamp 1654583406
transform 1 0 17357 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_148
timestamp 1654583406
transform 1 0 17158 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_149
timestamp 1654583406
transform 1 0 17894 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_150
timestamp 1654583406
transform 1 0 17357 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_151
timestamp 1654583406
transform 1 0 17802 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_152
timestamp 1654583406
transform 1 0 17787 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_153
timestamp 1654583406
transform 1 0 15502 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_154
timestamp 1654583406
transform 1 0 15211 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_155
timestamp 1654583406
transform 1 0 17710 0 1 12614
box -29 -23 29 23
use L1M1_PR  L1M1_PR_156
timestamp 1654583406
transform 1 0 17357 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_157
timestamp 1654583406
transform 1 0 17787 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_158
timestamp 1654583406
transform 1 0 15870 0 1 12342
box -29 -23 29 23
use L1M1_PR  L1M1_PR_159
timestamp 1654583406
transform 1 0 16063 0 1 13167
box -29 -23 29 23
use L1M1_PR  L1M1_PR_160
timestamp 1654583406
transform 1 0 15686 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_161
timestamp 1654583406
transform 1 0 16063 0 1 12079
box -29 -23 29 23
use L1M1_PR  L1M1_PR_162
timestamp 1654583406
transform 1 0 14766 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_163
timestamp 1654583406
transform 1 0 12834 0 1 13430
box -29 -23 29 23
use L1M1_PR  L1M1_PR_164
timestamp 1654583406
transform 1 0 12359 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_165
timestamp 1654583406
transform 1 0 13923 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_166
timestamp 1654583406
transform 1 0 12006 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_167
timestamp 1654583406
transform 1 0 12205 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_168
timestamp 1654583406
transform 1 0 12190 0 1 13974
box -29 -23 29 23
use L1M1_PR  L1M1_PR_169
timestamp 1654583406
transform 1 0 11347 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_170
timestamp 1654583406
transform 1 0 10914 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_171
timestamp 1654583406
transform 1 0 13953 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_172
timestamp 1654583406
transform 1 0 13478 0 1 16966
box -29 -23 29 23
use L1M1_PR  L1M1_PR_173
timestamp 1654583406
transform 1 0 14775 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_174
timestamp 1654583406
transform 1 0 13478 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_175
timestamp 1654583406
transform 1 0 17158 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_176
timestamp 1654583406
transform 1 0 17158 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_177
timestamp 1654583406
transform 1 0 14306 0 1 15130
box -29 -23 29 23
use L1M1_PR  L1M1_PR_178
timestamp 1654583406
transform 1 0 10442 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_179
timestamp 1654583406
transform 1 0 13662 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_180
timestamp 1654583406
transform 1 0 13018 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_181
timestamp 1654583406
transform 1 0 12834 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_182
timestamp 1654583406
transform 1 0 12742 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_183
timestamp 1654583406
transform 1 0 12466 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_184
timestamp 1654583406
transform 1 0 12098 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_185
timestamp 1654583406
transform 1 0 11454 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_186
timestamp 1654583406
transform 1 0 11086 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_187
timestamp 1654583406
transform 1 0 10810 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_188
timestamp 1654583406
transform 1 0 17618 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_189
timestamp 1654583406
transform 1 0 17618 0 1 14722
box -29 -23 29 23
use L1M1_PR  L1M1_PR_190
timestamp 1654583406
transform 1 0 17618 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_191
timestamp 1654583406
transform 1 0 17526 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_192
timestamp 1654583406
transform 1 0 16330 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_193
timestamp 1654583406
transform 1 0 16330 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_194
timestamp 1654583406
transform 1 0 16054 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_195
timestamp 1654583406
transform 1 0 15042 0 1 15810
box -29 -23 29 23
use L1M1_PR  L1M1_PR_196
timestamp 1654583406
transform 1 0 15042 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_197
timestamp 1654583406
transform 1 0 14950 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_198
timestamp 1654583406
transform 1 0 14214 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_199
timestamp 1654583406
transform 1 0 18814 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_200
timestamp 1654583406
transform 1 0 17618 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_201
timestamp 1654583406
transform 1 0 17526 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_202
timestamp 1654583406
transform 1 0 17526 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_203
timestamp 1654583406
transform 1 0 17526 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_204
timestamp 1654583406
transform 1 0 16974 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_205
timestamp 1654583406
transform 1 0 15962 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_206
timestamp 1654583406
transform 1 0 15042 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_207
timestamp 1654583406
transform 1 0 15042 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_208
timestamp 1654583406
transform 1 0 14950 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_209
timestamp 1654583406
transform 1 0 8602 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_210
timestamp 1654583406
transform 1 0 7958 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_211
timestamp 1654583406
transform 1 0 9062 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_212
timestamp 1654583406
transform 1 0 6026 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_213
timestamp 1654583406
transform 1 0 7314 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_214
timestamp 1654583406
transform 1 0 6486 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_215
timestamp 1654583406
transform 1 0 9706 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_216
timestamp 1654583406
transform 1 0 7774 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_217
timestamp 1654583406
transform 1 0 9982 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_218
timestamp 1654583406
transform 1 0 9430 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_219
timestamp 1654583406
transform 1 0 8970 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_220
timestamp 1654583406
transform 1 0 6946 0 1 17578
box -29 -23 29 23
use L1M1_PR  L1M1_PR_221
timestamp 1654583406
transform 1 0 8234 0 1 20842
box -29 -23 29 23
use L1M1_PR  L1M1_PR_222
timestamp 1654583406
transform 1 0 7590 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_223
timestamp 1654583406
transform 1 0 7498 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_224
timestamp 1654583406
transform 1 0 7498 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_225
timestamp 1654583406
transform 1 0 7406 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_226
timestamp 1654583406
transform 1 0 6670 0 1 17374
box -29 -23 29 23
use L1M1_PR  L1M1_PR_227
timestamp 1654583406
transform 1 0 7866 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_228
timestamp 1654583406
transform 1 0 7406 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_229
timestamp 1654583406
transform 1 0 6762 0 1 17374
box -29 -23 29 23
use L1M1_PR  L1M1_PR_230
timestamp 1654583406
transform 1 0 9246 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_231
timestamp 1654583406
transform 1 0 9062 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_232
timestamp 1654583406
transform 1 0 9062 0 1 17578
box -29 -23 29 23
use L1M1_PR  L1M1_PR_233
timestamp 1654583406
transform 1 0 9890 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_234
timestamp 1654583406
transform 1 0 9890 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_235
timestamp 1654583406
transform 1 0 9338 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_236
timestamp 1654583406
transform 1 0 7682 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_237
timestamp 1654583406
transform 1 0 7498 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_238
timestamp 1654583406
transform 1 0 7222 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_239
timestamp 1654583406
transform 1 0 7774 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_240
timestamp 1654583406
transform 1 0 6210 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_241
timestamp 1654583406
transform 1 0 6118 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_242
timestamp 1654583406
transform 1 0 6118 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_243
timestamp 1654583406
transform 1 0 8878 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_244
timestamp 1654583406
transform 1 0 8786 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_245
timestamp 1654583406
transform 1 0 8510 0 1 20230
box -29 -23 29 23
use L1M1_PR  L1M1_PR_246
timestamp 1654583406
transform 1 0 9154 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_247
timestamp 1654583406
transform 1 0 8050 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_248
timestamp 1654583406
transform 1 0 7682 0 1 20298
box -29 -23 29 23
use L1M1_PR  L1M1_PR_249
timestamp 1654583406
transform 1 0 8786 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_250
timestamp 1654583406
transform 1 0 7682 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_251
timestamp 1654583406
transform 1 0 7498 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_252
timestamp 1654583406
transform 1 0 9246 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_253
timestamp 1654583406
transform 1 0 9246 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_254
timestamp 1654583406
transform 1 0 9062 0 1 16966
box -29 -23 29 23
use L1M1_PR  L1M1_PR_255
timestamp 1654583406
transform 1 0 8970 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_256
timestamp 1654583406
transform 1 0 8970 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_257
timestamp 1654583406
transform 1 0 7590 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_258
timestamp 1654583406
transform 1 0 6379 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_259
timestamp 1654583406
transform 1 0 6302 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_260
timestamp 1654583406
transform 1 0 6563 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_261
timestamp 1654583406
transform 1 0 6302 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_262
timestamp 1654583406
transform 1 0 9629 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_263
timestamp 1654583406
transform 1 0 8878 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_264
timestamp 1654583406
transform 1 0 7958 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_265
timestamp 1654583406
transform 1 0 7237 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_266
timestamp 1654583406
transform 1 0 8341 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_267
timestamp 1654583406
transform 1 0 7590 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_268
timestamp 1654583406
transform 1 0 8771 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_269
timestamp 1654583406
transform 1 0 8326 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_270
timestamp 1654583406
transform 1 0 7958 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_271
timestamp 1654583406
transform 1 0 7943 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_272
timestamp 1654583406
transform 1 0 6486 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_273
timestamp 1654583406
transform 1 0 6287 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_274
timestamp 1654583406
transform 1 0 6394 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_275
timestamp 1654583406
transform 1 0 6379 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_276
timestamp 1654583406
transform 1 0 15962 0 1 14042
box -29 -23 29 23
use L1M1_PR  L1M1_PR_277
timestamp 1654583406
transform 1 0 13938 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_278
timestamp 1654583406
transform 1 0 13938 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_279
timestamp 1654583406
transform 1 0 10258 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_280
timestamp 1654583406
transform 1 0 10059 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_281
timestamp 1654583406
transform 1 0 15686 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_282
timestamp 1654583406
transform 1 0 14122 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_283
timestamp 1654583406
transform 1 0 14122 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_284
timestamp 1654583406
transform 1 0 11362 0 1 15810
box -29 -23 29 23
use L1M1_PR  L1M1_PR_285
timestamp 1654583406
transform 1 0 9890 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_286
timestamp 1654583406
transform 1 0 8970 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_287
timestamp 1654583406
transform 1 0 7222 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_288
timestamp 1654583406
transform 1 0 5658 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_289
timestamp 1654583406
transform 1 0 9430 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_290
timestamp 1654583406
transform 1 0 8510 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_291
timestamp 1654583406
transform 1 0 7590 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_292
timestamp 1654583406
transform 1 0 6854 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_293
timestamp 1654583406
transform 1 0 8142 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_294
timestamp 1654583406
transform 1 0 7222 0 1 17374
box -29 -23 29 23
use L1M1_PR  L1M1_PR_295
timestamp 1654583406
transform 1 0 10534 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_296
timestamp 1654583406
transform 1 0 8694 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_297
timestamp 1654583406
transform 1 0 8602 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_298
timestamp 1654583406
transform 1 0 8326 0 1 16966
box -29 -23 29 23
use L1M1_PR  L1M1_PR_299
timestamp 1654583406
transform 1 0 7314 0 1 15062
box -29 -23 29 23
use L1M1_PR  L1M1_PR_300
timestamp 1654583406
transform 1 0 6762 0 1 14110
box -29 -23 29 23
use L1M1_PR  L1M1_PR_301
timestamp 1654583406
transform 1 0 13754 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_302
timestamp 1654583406
transform 1 0 13662 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_303
timestamp 1654583406
transform 1 0 12834 0 1 12954
box -29 -23 29 23
use L1M1_PR  L1M1_PR_304
timestamp 1654583406
transform 1 0 10810 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_305
timestamp 1654583406
transform 1 0 9798 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_306
timestamp 1654583406
transform 1 0 9798 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_307
timestamp 1654583406
transform 1 0 9522 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_308
timestamp 1654583406
transform 1 0 9522 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_309
timestamp 1654583406
transform 1 0 9430 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_310
timestamp 1654583406
transform 1 0 21482 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_311
timestamp 1654583406
transform 1 0 20194 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_312
timestamp 1654583406
transform 1 0 20194 0 1 14722
box -29 -23 29 23
use L1M1_PR  L1M1_PR_313
timestamp 1654583406
transform 1 0 20194 0 1 12546
box -29 -23 29 23
use L1M1_PR  L1M1_PR_314
timestamp 1654583406
transform 1 0 19182 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_315
timestamp 1654583406
transform 1 0 18906 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_316
timestamp 1654583406
transform 1 0 18906 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_317
timestamp 1654583406
transform 1 0 17618 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_318
timestamp 1654583406
transform 1 0 17618 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_319
timestamp 1654583406
transform 1 0 17342 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_320
timestamp 1654583406
transform 1 0 17066 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_321
timestamp 1654583406
transform 1 0 18906 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_322
timestamp 1654583406
transform 1 0 18814 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_323
timestamp 1654583406
transform 1 0 18538 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_324
timestamp 1654583406
transform 1 0 17710 0 1 19550
box -29 -23 29 23
use L1M1_PR  L1M1_PR_325
timestamp 1654583406
transform 1 0 15042 0 1 19550
box -29 -23 29 23
use L1M1_PR  L1M1_PR_326
timestamp 1654583406
transform 1 0 15042 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_327
timestamp 1654583406
transform 1 0 14582 0 1 19550
box -29 -23 29 23
use L1M1_PR  L1M1_PR_328
timestamp 1654583406
transform 1 0 13754 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_329
timestamp 1654583406
transform 1 0 12834 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_330
timestamp 1654583406
transform 1 0 12466 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_331
timestamp 1654583406
transform 1 0 11270 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_332
timestamp 1654583406
transform 1 0 10442 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_333
timestamp 1654583406
transform 1 0 13386 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_334
timestamp 1654583406
transform 1 0 11730 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_335
timestamp 1654583406
transform 1 0 14030 0 1 21318
box -29 -23 29 23
use L1M1_PR  L1M1_PR_336
timestamp 1654583406
transform 1 0 13110 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_337
timestamp 1654583406
transform 1 0 15134 0 1 21318
box -29 -23 29 23
use L1M1_PR  L1M1_PR_338
timestamp 1654583406
transform 1 0 14490 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_339
timestamp 1654583406
transform 1 0 17802 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_340
timestamp 1654583406
transform 1 0 15594 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_341
timestamp 1654583406
transform 1 0 18906 0 1 20298
box -29 -23 29 23
use L1M1_PR  L1M1_PR_342
timestamp 1654583406
transform 1 0 17526 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_343
timestamp 1654583406
transform 1 0 21482 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_344
timestamp 1654583406
transform 1 0 19366 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_345
timestamp 1654583406
transform 1 0 21114 0 1 19550
box -29 -23 29 23
use L1M1_PR  L1M1_PR_346
timestamp 1654583406
transform 1 0 20930 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_347
timestamp 1654583406
transform 1 0 22057 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_348
timestamp 1654583406
transform 1 0 21850 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_349
timestamp 1654583406
transform 1 0 21390 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_350
timestamp 1654583406
transform 1 0 20631 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_351
timestamp 1654583406
transform 1 0 22509 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_352
timestamp 1654583406
transform 1 0 21482 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_353
timestamp 1654583406
transform 1 0 22509 0 1 12614
box -29 -23 29 23
use L1M1_PR  L1M1_PR_354
timestamp 1654583406
transform 1 0 22034 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_355
timestamp 1654583406
transform 1 0 21482 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_356
timestamp 1654583406
transform 1 0 20907 0 1 10778
box -29 -23 29 23
use L1M1_PR  L1M1_PR_357
timestamp 1654583406
transform 1 0 22517 0 1 9350
box -29 -23 29 23
use L1M1_PR  L1M1_PR_358
timestamp 1654583406
transform 1 0 21482 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_359
timestamp 1654583406
transform 1 0 22517 0 1 8262
box -29 -23 29 23
use L1M1_PR  L1M1_PR_360
timestamp 1654583406
transform 1 0 21574 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_361
timestamp 1654583406
transform 1 0 20539 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_362
timestamp 1654583406
transform 1 0 20286 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_363
timestamp 1654583406
transform 1 0 19251 0 1 7174
box -29 -23 29 23
use L1M1_PR  L1M1_PR_364
timestamp 1654583406
transform 1 0 18814 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_365
timestamp 1654583406
transform 1 0 19941 0 1 9350
box -29 -23 29 23
use L1M1_PR  L1M1_PR_366
timestamp 1654583406
transform 1 0 17802 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_367
timestamp 1654583406
transform 1 0 16675 0 1 9350
box -29 -23 29 23
use L1M1_PR  L1M1_PR_368
timestamp 1654583406
transform 1 0 16514 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_369
timestamp 1654583406
transform 1 0 15387 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_370
timestamp 1654583406
transform 1 0 14122 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_371
timestamp 1654583406
transform 1 0 12811 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_372
timestamp 1654583406
transform 1 0 10718 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_373
timestamp 1654583406
transform 1 0 11753 0 1 10778
box -29 -23 29 23
use L1M1_PR  L1M1_PR_374
timestamp 1654583406
transform 1 0 9982 0 1 10438
box -29 -23 29 23
use L1M1_PR  L1M1_PR_375
timestamp 1654583406
transform 1 0 8947 0 1 10438
box -29 -23 29 23
use L1M1_PR  L1M1_PR_376
timestamp 1654583406
transform 1 0 8786 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_377
timestamp 1654583406
transform 1 0 8694 0 1 13974
box -29 -23 29 23
use L1M1_PR  L1M1_PR_378
timestamp 1654583406
transform 1 0 7751 0 1 10778
box -29 -23 29 23
use L1M1_PR  L1M1_PR_379
timestamp 1654583406
transform 1 0 7659 0 1 14042
box -29 -23 29 23
use L1M1_PR  L1M1_PR_380
timestamp 1654583406
transform 1 0 6946 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_381
timestamp 1654583406
transform 1 0 10810 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_382
timestamp 1654583406
transform 1 0 9062 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_383
timestamp 1654583406
transform 1 0 11377 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_384
timestamp 1654583406
transform 1 0 10166 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_385
timestamp 1654583406
transform 1 0 10519 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_386
timestamp 1654583406
transform 1 0 10442 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_387
timestamp 1654583406
transform 1 0 13095 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_388
timestamp 1654583406
transform 1 0 12006 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_389
timestamp 1654583406
transform 1 0 12374 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_390
timestamp 1654583406
transform 1 0 12359 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_391
timestamp 1654583406
transform 1 0 14965 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_392
timestamp 1654583406
transform 1 0 14674 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_393
timestamp 1654583406
transform 1 0 17357 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_394
timestamp 1654583406
transform 1 0 15778 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_395
timestamp 1654583406
transform 1 0 16330 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_396
timestamp 1654583406
transform 1 0 16223 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_397
timestamp 1654583406
transform 1 0 18814 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_398
timestamp 1654583406
transform 1 0 18799 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_399
timestamp 1654583406
transform 1 0 20823 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_400
timestamp 1654583406
transform 1 0 20562 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_401
timestamp 1654583406
transform 1 0 22509 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_402
timestamp 1654583406
transform 1 0 21758 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_403
timestamp 1654583406
transform 1 0 22509 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_404
timestamp 1654583406
transform 1 0 21758 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_405
timestamp 1654583406
transform 1 0 22509 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_406
timestamp 1654583406
transform 1 0 22126 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_407
timestamp 1654583406
transform 1 0 21574 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_408
timestamp 1654583406
transform 1 0 21221 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_409
timestamp 1654583406
transform 1 0 19351 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_410
timestamp 1654583406
transform 1 0 19274 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_411
timestamp 1654583406
transform 1 0 21651 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_412
timestamp 1654583406
transform 1 0 20930 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_413
timestamp 1654583406
transform 1 0 20363 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_414
timestamp 1654583406
transform 1 0 19458 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_415
timestamp 1654583406
transform 1 0 19070 0 1 10225
box -29 -23 29 23
use L1M1_PR  L1M1_PR_416
timestamp 1654583406
transform 1 0 18262 0 1 10166
box -29 -23 29 23
use L1M1_PR  L1M1_PR_417
timestamp 1654583406
transform 1 0 17787 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_418
timestamp 1654583406
transform 1 0 17250 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_419
timestamp 1654583406
transform 1 0 17710 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_420
timestamp 1654583406
transform 1 0 17357 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_421
timestamp 1654583406
transform 1 0 16790 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_422
timestamp 1654583406
transform 1 0 14935 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_423
timestamp 1654583406
transform 1 0 14122 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_424
timestamp 1654583406
transform 1 0 13923 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_425
timestamp 1654583406
transform 1 0 14030 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_426
timestamp 1654583406
transform 1 0 13509 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_427
timestamp 1654583406
transform 1 0 13202 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_428
timestamp 1654583406
transform 1 0 12481 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_429
timestamp 1654583406
transform 1 0 10549 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_430
timestamp 1654583406
transform 1 0 10442 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_431
timestamp 1654583406
transform 1 0 8878 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_432
timestamp 1654583406
transform 1 0 8219 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_433
timestamp 1654583406
transform 1 0 8326 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_434
timestamp 1654583406
transform 1 0 8127 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_435
timestamp 1654583406
transform 1 0 9139 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_436
timestamp 1654583406
transform 1 0 8050 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_437
timestamp 1654583406
transform 1 0 9798 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_438
timestamp 1654583406
transform 1 0 9430 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_439
timestamp 1654583406
transform 1 0 10074 0 1 21318
box -29 -23 29 23
use L1M1_PR  L1M1_PR_440
timestamp 1654583406
transform 1 0 9890 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_441
timestamp 1654583406
transform 1 0 12098 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_442
timestamp 1654583406
transform 1 0 11638 0 1 21318
box -29 -23 29 23
use L1M1_PR  L1M1_PR_443
timestamp 1654583406
transform 1 0 12742 0 1 20570
box -29 -23 29 23
use L1M1_PR  L1M1_PR_444
timestamp 1654583406
transform 1 0 12558 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_445
timestamp 1654583406
transform 1 0 14858 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_446
timestamp 1654583406
transform 1 0 14306 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_447
timestamp 1654583406
transform 1 0 15962 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_448
timestamp 1654583406
transform 1 0 15410 0 1 20230
box -29 -23 29 23
use L1M1_PR  L1M1_PR_449
timestamp 1654583406
transform 1 0 16974 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_450
timestamp 1654583406
transform 1 0 16698 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_451
timestamp 1654583406
transform 1 0 19734 0 1 20298
box -29 -23 29 23
use L1M1_PR  L1M1_PR_452
timestamp 1654583406
transform 1 0 19182 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_453
timestamp 1654583406
transform 1 0 20654 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_454
timestamp 1654583406
transform 1 0 20194 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_455
timestamp 1654583406
transform 1 0 22402 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_456
timestamp 1654583406
transform 1 0 21390 0 1 20162
box -29 -23 29 23
use L1M1_PR  L1M1_PR_457
timestamp 1654583406
transform 1 0 21390 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_458
timestamp 1654583406
transform 1 0 20286 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_459
timestamp 1654583406
transform 1 0 23138 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_460
timestamp 1654583406
transform 1 0 22494 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_461
timestamp 1654583406
transform 1 0 23046 0 1 12954
box -29 -23 29 23
use L1M1_PR  L1M1_PR_462
timestamp 1654583406
transform 1 0 21942 0 1 12954
box -29 -23 29 23
use L1M1_PR  L1M1_PR_463
timestamp 1654583406
transform 1 0 22862 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_464
timestamp 1654583406
transform 1 0 20562 0 1 9350
box -29 -23 29 23
use L1M1_PR  L1M1_PR_465
timestamp 1654583406
transform 1 0 22954 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_466
timestamp 1654583406
transform 1 0 19826 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_467
timestamp 1654583406
transform 1 0 20194 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_468
timestamp 1654583406
transform 1 0 18630 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_469
timestamp 1654583406
transform 1 0 18906 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_470
timestamp 1654583406
transform 1 0 16882 0 1 11866
box -29 -23 29 23
use L1M1_PR  L1M1_PR_471
timestamp 1654583406
transform 1 0 20286 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_472
timestamp 1654583406
transform 1 0 18078 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_473
timestamp 1654583406
transform 1 0 16422 0 1 11866
box -29 -23 29 23
use L1M1_PR  L1M1_PR_474
timestamp 1654583406
transform 1 0 16330 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_475
timestamp 1654583406
transform 1 0 15042 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_476
timestamp 1654583406
transform 1 0 14490 0 1 10778
box -29 -23 29 23
use L1M1_PR  L1M1_PR_477
timestamp 1654583406
transform 1 0 13662 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_478
timestamp 1654583406
transform 1 0 12466 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_479
timestamp 1654583406
transform 1 0 12834 0 1 11526
box -29 -23 29 23
use L1M1_PR  L1M1_PR_480
timestamp 1654583406
transform 1 0 12190 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_481
timestamp 1654583406
transform 1 0 10074 0 1 10778
box -29 -23 29 23
use L1M1_PR  L1M1_PR_482
timestamp 1654583406
transform 1 0 8602 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_483
timestamp 1654583406
transform 1 0 8510 0 1 11458
box -29 -23 29 23
use L1M1_PR  L1M1_PR_484
timestamp 1654583406
transform 1 0 7406 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_485
timestamp 1654583406
transform 1 0 7958 0 1 14722
box -29 -23 29 23
use L1M1_PR  L1M1_PR_486
timestamp 1654583406
transform 1 0 7314 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_487
timestamp 1654583406
transform 1 0 7590 0 1 13430
box -29 -23 29 23
use L1M1_PR  L1M1_PR_488
timestamp 1654583406
transform 1 0 6118 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_489
timestamp 1654583406
transform 1 0 23138 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_490
timestamp 1654583406
transform 1 0 22770 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_491
timestamp 1654583406
transform 1 0 22126 0 1 14246
box -29 -23 29 23
use L1M1_PR  L1M1_PR_492
timestamp 1654583406
transform 1 0 22494 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_493
timestamp 1654583406
transform 1 0 22218 0 1 17374
box -29 -23 29 23
use L1M1_PR  L1M1_PR_494
timestamp 1654583406
transform 1 0 22218 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_495
timestamp 1654583406
transform 1 0 22862 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_496
timestamp 1654583406
transform 1 0 22310 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_497
timestamp 1654583406
transform 1 0 21850 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_498
timestamp 1654583406
transform 1 0 22770 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_499
timestamp 1654583406
transform 1 0 22494 0 1 14042
box -29 -23 29 23
use L1M1_PR  L1M1_PR_500
timestamp 1654583406
transform 1 0 22218 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_501
timestamp 1654583406
transform 1 0 22862 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_502
timestamp 1654583406
transform 1 0 22770 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_503
timestamp 1654583406
transform 1 0 22494 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_504
timestamp 1654583406
transform 1 0 22402 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_505
timestamp 1654583406
transform 1 0 22770 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_506
timestamp 1654583406
transform 1 0 22218 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_507
timestamp 1654583406
transform 1 0 22678 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_508
timestamp 1654583406
transform 1 0 22402 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_509
timestamp 1654583406
transform 1 0 22126 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_510
timestamp 1654583406
transform 1 0 21942 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_511
timestamp 1654583406
transform 1 0 22310 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_512
timestamp 1654583406
transform 1 0 20102 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_513
timestamp 1654583406
transform 1 0 19642 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_514
timestamp 1654583406
transform 1 0 20562 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_515
timestamp 1654583406
transform 1 0 19826 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_516
timestamp 1654583406
transform 1 0 19734 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_517
timestamp 1654583406
transform 1 0 19642 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_518
timestamp 1654583406
transform 1 0 19550 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_519
timestamp 1654583406
transform 1 0 19366 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_520
timestamp 1654583406
transform 1 0 19366 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_521
timestamp 1654583406
transform 1 0 18998 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_522
timestamp 1654583406
transform 1 0 17802 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_523
timestamp 1654583406
transform 1 0 18354 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_524
timestamp 1654583406
transform 1 0 18354 0 1 5814
box -29 -23 29 23
use L1M1_PR  L1M1_PR_525
timestamp 1654583406
transform 1 0 17894 0 1 5814
box -29 -23 29 23
use L1M1_PR  L1M1_PR_526
timestamp 1654583406
transform 1 0 18998 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_527
timestamp 1654583406
transform 1 0 18630 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_528
timestamp 1654583406
transform 1 0 18446 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_529
timestamp 1654583406
transform 1 0 17963 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_530
timestamp 1654583406
transform 1 0 16514 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_531
timestamp 1654583406
transform 1 0 15387 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_532
timestamp 1654583406
transform 1 0 15226 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_533
timestamp 1654583406
transform 1 0 14398 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_534
timestamp 1654583406
transform 1 0 14099 0 1 8262
box -29 -23 29 23
use L1M1_PR  L1M1_PR_535
timestamp 1654583406
transform 1 0 13271 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_536
timestamp 1654583406
transform 1 0 12098 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_537
timestamp 1654583406
transform 1 0 11063 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_538
timestamp 1654583406
transform 1 0 9890 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_539
timestamp 1654583406
transform 1 0 10925 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_540
timestamp 1654583406
transform 1 0 9982 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_541
timestamp 1654583406
transform 1 0 8970 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_542
timestamp 1654583406
transform 1 0 8947 0 1 8262
box -29 -23 29 23
use L1M1_PR  L1M1_PR_543
timestamp 1654583406
transform 1 0 7935 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_544
timestamp 1654583406
transform 1 0 6946 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_545
timestamp 1654583406
transform 1 0 6210 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_546
timestamp 1654583406
transform 1 0 6747 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_547
timestamp 1654583406
transform 1 0 6578 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_548
timestamp 1654583406
transform 1 0 6471 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_549
timestamp 1654583406
transform 1 0 6394 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_550
timestamp 1654583406
transform 1 0 8970 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_551
timestamp 1654583406
transform 1 0 7483 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_552
timestamp 1654583406
transform 1 0 11454 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_553
timestamp 1654583406
transform 1 0 10181 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_554
timestamp 1654583406
transform 1 0 10917 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_555
timestamp 1654583406
transform 1 0 10902 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_556
timestamp 1654583406
transform 1 0 12374 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_557
timestamp 1654583406
transform 1 0 12359 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_558
timestamp 1654583406
transform 1 0 14659 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_559
timestamp 1654583406
transform 1 0 14398 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_560
timestamp 1654583406
transform 1 0 16253 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_561
timestamp 1654583406
transform 1 0 16054 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_562
timestamp 1654583406
transform 1 0 18078 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_563
timestamp 1654583406
transform 1 0 17787 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_564
timestamp 1654583406
transform 1 0 17235 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_565
timestamp 1654583406
transform 1 0 16974 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_566
timestamp 1654583406
transform 1 0 18998 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_567
timestamp 1654583406
transform 1 0 17971 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_568
timestamp 1654583406
transform 1 0 19458 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_569
timestamp 1654583406
transform 1 0 19167 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_570
timestamp 1654583406
transform 1 0 21191 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_571
timestamp 1654583406
transform 1 0 21114 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_572
timestamp 1654583406
transform 1 0 22126 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_573
timestamp 1654583406
transform 1 0 21651 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_574
timestamp 1654583406
transform 1 0 21574 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_575
timestamp 1654583406
transform 1 0 21221 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_576
timestamp 1654583406
transform 1 0 21221 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_577
timestamp 1654583406
transform 1 0 21022 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_578
timestamp 1654583406
transform 1 0 21850 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_579
timestamp 1654583406
transform 1 0 21497 0 1 17519
box -29 -23 29 23
use L1M1_PR  L1M1_PR_580
timestamp 1654583406
transform 1 0 22517 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_581
timestamp 1654583406
transform 1 0 22494 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_582
timestamp 1654583406
transform 1 0 22402 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_583
timestamp 1654583406
transform 1 0 22218 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_584
timestamp 1654583406
transform 1 0 22126 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_585
timestamp 1654583406
transform 1 0 22034 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_586
timestamp 1654583406
transform 1 0 22126 0 1 13974
box -29 -23 29 23
use L1M1_PR  L1M1_PR_587
timestamp 1654583406
transform 1 0 20654 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_588
timestamp 1654583406
transform 1 0 22494 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_589
timestamp 1654583406
transform 1 0 22402 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_590
timestamp 1654583406
transform 1 0 21758 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_591
timestamp 1654583406
transform 1 0 20746 0 1 8262
box -29 -23 29 23
use L1M1_PR  L1M1_PR_592
timestamp 1654583406
transform 1 0 19918 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_593
timestamp 1654583406
transform 1 0 19826 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_594
timestamp 1654583406
transform 1 0 19550 0 1 6086
box -29 -23 29 23
use L1M1_PR  L1M1_PR_595
timestamp 1654583406
transform 1 0 19366 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_596
timestamp 1654583406
transform 1 0 18170 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_597
timestamp 1654583406
transform 1 0 17342 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_598
timestamp 1654583406
transform 1 0 17710 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_599
timestamp 1654583406
transform 1 0 17618 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_600
timestamp 1654583406
transform 1 0 15686 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_601
timestamp 1654583406
transform 1 0 15042 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_602
timestamp 1654583406
transform 1 0 14030 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_603
timestamp 1654583406
transform 1 0 13754 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_604
timestamp 1654583406
transform 1 0 12834 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_605
timestamp 1654583406
transform 1 0 12742 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_606
timestamp 1654583406
transform 1 0 10626 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_607
timestamp 1654583406
transform 1 0 10534 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_608
timestamp 1654583406
transform 1 0 11914 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_609
timestamp 1654583406
transform 1 0 11362 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_610
timestamp 1654583406
transform 1 0 8602 0 1 9350
box -29 -23 29 23
use L1M1_PR  L1M1_PR_611
timestamp 1654583406
transform 1 0 8602 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_612
timestamp 1654583406
transform 1 0 6118 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_613
timestamp 1654583406
transform 1 0 6026 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_614
timestamp 1654583406
transform 1 0 14582 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_615
timestamp 1654583406
transform 1 0 14490 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_616
timestamp 1654583406
transform 1 0 13018 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_617
timestamp 1654583406
transform 1 0 12834 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_618
timestamp 1654583406
transform 1 0 15594 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_619
timestamp 1654583406
transform 1 0 14674 0 1 5882
box -29 -23 29 23
use L1M1_PR  L1M1_PR_620
timestamp 1654583406
transform 1 0 14214 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_621
timestamp 1654583406
transform 1 0 13294 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_622
timestamp 1654583406
transform 1 0 12650 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_623
timestamp 1654583406
transform 1 0 12926 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_624
timestamp 1654583406
transform 1 0 12558 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_625
timestamp 1654583406
transform 1 0 12558 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_626
timestamp 1654583406
transform 1 0 12558 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_627
timestamp 1654583406
transform 1 0 12834 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_628
timestamp 1654583406
transform 1 0 12374 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_629
timestamp 1654583406
transform 1 0 10718 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_630
timestamp 1654583406
transform 1 0 10534 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_631
timestamp 1654583406
transform 1 0 10534 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_632
timestamp 1654583406
transform 1 0 10442 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_633
timestamp 1654583406
transform 1 0 10350 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_634
timestamp 1654583406
transform 1 0 10534 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_635
timestamp 1654583406
transform 1 0 10258 0 1 5882
box -29 -23 29 23
use L1M1_PR  L1M1_PR_636
timestamp 1654583406
transform 1 0 9890 0 1 5882
box -29 -23 29 23
use L1M1_PR  L1M1_PR_637
timestamp 1654583406
transform 1 0 9246 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_638
timestamp 1654583406
transform 1 0 9614 0 1 5814
box -29 -23 29 23
use L1M1_PR  L1M1_PR_639
timestamp 1654583406
transform 1 0 8050 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_640
timestamp 1654583406
transform 1 0 7958 0 1 5814
box -29 -23 29 23
use L1M1_PR  L1M1_PR_641
timestamp 1654583406
transform 1 0 7958 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_642
timestamp 1654583406
transform 1 0 7866 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_643
timestamp 1654583406
transform 1 0 7866 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_644
timestamp 1654583406
transform 1 0 8142 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_645
timestamp 1654583406
transform 1 0 7682 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_646
timestamp 1654583406
transform 1 0 6762 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_647
timestamp 1654583406
transform 1 0 6394 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_648
timestamp 1654583406
transform 1 0 7314 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_649
timestamp 1654583406
transform 1 0 7038 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_650
timestamp 1654583406
transform 1 0 7222 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_651
timestamp 1654583406
transform 1 0 6210 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_652
timestamp 1654583406
transform 1 0 6026 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_653
timestamp 1654583406
transform 1 0 7231 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_654
timestamp 1654583406
transform 1 0 6486 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_655
timestamp 1654583406
transform 1 0 6946 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_656
timestamp 1654583406
transform 1 0 6471 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_657
timestamp 1654583406
transform 1 0 7483 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_658
timestamp 1654583406
transform 1 0 7314 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_659
timestamp 1654583406
transform 1 0 8771 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_660
timestamp 1654583406
transform 1 0 8510 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_661
timestamp 1654583406
transform 1 0 11362 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_662
timestamp 1654583406
transform 1 0 11071 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_663
timestamp 1654583406
transform 1 0 11822 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_664
timestamp 1654583406
transform 1 0 11347 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_665
timestamp 1654583406
transform 1 0 13647 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_666
timestamp 1654583406
transform 1 0 13294 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_667
timestamp 1654583406
transform 1 0 16494 0 1 6961
box -29 -23 29 23
use L1M1_PR  L1M1_PR_668
timestamp 1654583406
transform 1 0 15778 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_669
timestamp 1654583406
transform 1 0 13923 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_670
timestamp 1654583406
transform 1 0 13018 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_671
timestamp 1654583406
transform 1 0 15410 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_672
timestamp 1654583406
transform 1 0 15134 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_673
timestamp 1654583406
transform 1 0 12834 0 1 7174
box -29 -23 29 23
use L1M1_PR  L1M1_PR_674
timestamp 1654583406
transform 1 0 12834 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_675
timestamp 1654583406
transform 1 0 12374 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_676
timestamp 1654583406
transform 1 0 12190 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_677
timestamp 1654583406
transform 1 0 11730 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_678
timestamp 1654583406
transform 1 0 10810 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_679
timestamp 1654583406
transform 1 0 8050 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_680
timestamp 1654583406
transform 1 0 7682 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_681
timestamp 1654583406
transform 1 0 6578 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_682
timestamp 1654583406
transform 1 0 6578 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_683
timestamp 1654583406
transform 1 0 6394 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_684
timestamp 1654583406
transform 1 0 6026 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_685
timestamp 1654583406
transform 1 0 10258 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_686
timestamp 1654583406
transform 1 0 10059 0 1 14246
box -29 -23 29 23
use L1M1_PR  L1M1_PR_687
timestamp 1654583406
transform 1 0 6670 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_688
timestamp 1654583406
transform 1 0 9691 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_689
timestamp 1654583406
transform 1 0 9246 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_690
timestamp 1654583406
transform 1 0 9783 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_691
timestamp 1654583406
transform 1 0 9338 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_692
timestamp 1654583406
transform 1 0 10059 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_693
timestamp 1654583406
transform 1 0 9430 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_694
timestamp 1654583406
transform 1 0 11270 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_695
timestamp 1654583406
transform 1 0 11071 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_696
timestamp 1654583406
transform 1 0 13493 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_697
timestamp 1654583406
transform 1 0 12374 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_698
timestamp 1654583406
transform 1 0 15042 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_699
timestamp 1654583406
transform 1 0 13923 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_700
timestamp 1654583406
transform 1 0 17357 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_701
timestamp 1654583406
transform 1 0 16146 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_702
timestamp 1654583406
transform 1 0 17075 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_703
timestamp 1654583406
transform 1 0 16238 0 1 10166
box -29 -23 29 23
use L1M1_PR  L1M1_PR_704
timestamp 1654583406
transform 1 0 18906 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_705
timestamp 1654583406
transform 1 0 17357 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_706
timestamp 1654583406
transform 1 0 20194 0 1 10166
box -29 -23 29 23
use L1M1_PR  L1M1_PR_707
timestamp 1654583406
transform 1 0 18645 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_708
timestamp 1654583406
transform 1 0 21482 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_709
timestamp 1654583406
transform 1 0 18921 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_710
timestamp 1654583406
transform 1 0 22770 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_711
timestamp 1654583406
transform 1 0 19933 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_712
timestamp 1654583406
transform 1 0 21221 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_713
timestamp 1654583406
transform 1 0 20470 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_714
timestamp 1654583406
transform 1 0 20102 0 1 15062
box -29 -23 29 23
use L1M1_PR  L1M1_PR_715
timestamp 1654583406
transform 1 0 19933 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_716
timestamp 1654583406
transform 1 0 21390 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_717
timestamp 1654583406
transform 1 0 18645 0 1 14246
box -29 -23 29 23
use L1M1_PR  L1M1_PR_718
timestamp 1654583406
transform 1 0 21390 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_719
timestamp 1654583406
transform 1 0 19933 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_720
timestamp 1654583406
transform 1 0 21390 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_721
timestamp 1654583406
transform 1 0 19167 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_722
timestamp 1654583406
transform 1 0 21942 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_723
timestamp 1654583406
transform 1 0 21298 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_724
timestamp 1654583406
transform 1 0 18805 0 1 18608
box -29 -23 29 23
use L1M1_PR  L1M1_PR_725
timestamp 1654583406
transform 1 0 19918 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_726
timestamp 1654583406
transform 1 0 19090 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_727
timestamp 1654583406
transform 1 0 19075 0 1 18938
box -29 -23 29 23
use L1M1_PR  L1M1_PR_728
timestamp 1654583406
transform 1 0 17971 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_729
timestamp 1654583406
transform 1 0 17618 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_730
timestamp 1654583406
transform 1 0 17342 0 1 20842
box -29 -23 29 23
use L1M1_PR  L1M1_PR_731
timestamp 1654583406
transform 1 0 16238 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_732
timestamp 1654583406
transform 1 0 15318 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_733
timestamp 1654583406
transform 1 0 15303 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_734
timestamp 1654583406
transform 1 0 14321 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_735
timestamp 1654583406
transform 1 0 14214 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_736
timestamp 1654583406
transform 1 0 13846 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_737
timestamp 1654583406
transform 1 0 13493 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_738
timestamp 1654583406
transform 1 0 13478 0 1 20298
box -29 -23 29 23
use L1M1_PR  L1M1_PR_739
timestamp 1654583406
transform 1 0 13202 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_740
timestamp 1654583406
transform 1 0 14781 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_741
timestamp 1654583406
transform 1 0 14214 0 1 20842
box -29 -23 29 23
use L1M1_PR  L1M1_PR_742
timestamp 1654583406
transform 1 0 11454 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_743
timestamp 1654583406
transform 1 0 12205 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_744
timestamp 1654583406
transform 1 0 11638 0 1 20842
box -29 -23 29 23
use L1M1_PR  L1M1_PR_745
timestamp 1654583406
transform 1 0 11638 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_746
timestamp 1654583406
transform 1 0 10534 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_747
timestamp 1654583406
transform 1 0 10258 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_748
timestamp 1654583406
transform 1 0 9783 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_749
timestamp 1654583406
transform 1 0 9154 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_750
timestamp 1654583406
transform 1 0 7866 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_751
timestamp 1654583406
transform 1 0 6762 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_752
timestamp 1654583406
transform 1 0 6486 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_753
timestamp 1654583406
transform 1 0 7590 0 1 10166
box -29 -23 29 23
use L1M1_PR  L1M1_PR_754
timestamp 1654583406
transform 1 0 8602 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_755
timestamp 1654583406
transform 1 0 9062 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_756
timestamp 1654583406
transform 1 0 9798 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_757
timestamp 1654583406
transform 1 0 13478 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_758
timestamp 1654583406
transform 1 0 15778 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_759
timestamp 1654583406
transform 1 0 15134 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_760
timestamp 1654583406
transform 1 0 18906 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_761
timestamp 1654583406
transform 1 0 19274 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_762
timestamp 1654583406
transform 1 0 18538 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_763
timestamp 1654583406
transform 1 0 18354 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_764
timestamp 1654583406
transform 1 0 18170 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_765
timestamp 1654583406
transform 1 0 19458 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_766
timestamp 1654583406
transform 1 0 19274 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_767
timestamp 1654583406
transform 1 0 19182 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_768
timestamp 1654583406
transform 1 0 20746 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_769
timestamp 1654583406
transform 1 0 20286 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_770
timestamp 1654583406
transform 1 0 22494 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_771
timestamp 1654583406
transform 1 0 22310 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_772
timestamp 1654583406
transform 1 0 22126 0 1 8670
box -29 -23 29 23
use L1M1_PR  L1M1_PR_773
timestamp 1654583406
transform 1 0 23230 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_774
timestamp 1654583406
transform 1 0 22678 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_775
timestamp 1654583406
transform 1 0 22678 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_776
timestamp 1654583406
transform 1 0 22402 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_777
timestamp 1654583406
transform 1 0 20102 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_778
timestamp 1654583406
transform 1 0 21666 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_779
timestamp 1654583406
transform 1 0 20102 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_780
timestamp 1654583406
transform 1 0 22402 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_781
timestamp 1654583406
transform 1 0 22402 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_782
timestamp 1654583406
transform 1 0 21390 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_783
timestamp 1654583406
transform 1 0 22126 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_784
timestamp 1654583406
transform 1 0 20378 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_785
timestamp 1654583406
transform 1 0 6762 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_786
timestamp 1654583406
transform 1 0 6302 0 1 5882
box -29 -23 29 23
use L1M1_PR  L1M1_PR_787
timestamp 1654583406
transform 1 0 6118 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_788
timestamp 1654583406
transform 1 0 6118 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_789
timestamp 1654583406
transform 1 0 6026 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_790
timestamp 1654583406
transform 1 0 6026 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_791
timestamp 1654583406
transform 1 0 7590 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_792
timestamp 1654583406
transform 1 0 6946 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_793
timestamp 1654583406
transform 1 0 6486 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_794
timestamp 1654583406
transform 1 0 8602 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_795
timestamp 1654583406
transform 1 0 8050 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_796
timestamp 1654583406
transform 1 0 10074 0 1 6086
box -29 -23 29 23
use L1M1_PR  L1M1_PR_797
timestamp 1654583406
transform 1 0 9890 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_798
timestamp 1654583406
transform 1 0 9430 0 1 6086
box -29 -23 29 23
use L1M1_PR  L1M1_PR_799
timestamp 1654583406
transform 1 0 12190 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_800
timestamp 1654583406
transform 1 0 10534 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_801
timestamp 1654583406
transform 1 0 12742 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_802
timestamp 1654583406
transform 1 0 12650 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_803
timestamp 1654583406
transform 1 0 12466 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_804
timestamp 1654583406
transform 1 0 14766 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_805
timestamp 1654583406
transform 1 0 13386 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_806
timestamp 1654583406
transform 1 0 15042 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_807
timestamp 1654583406
transform 1 0 14766 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_808
timestamp 1654583406
transform 1 0 14398 0 1 6086
box -29 -23 29 23
use L1M1_PR  L1M1_PR_809
timestamp 1654583406
transform 1 0 17618 0 1 7174
box -29 -23 29 23
use L1M1_PR  L1M1_PR_810
timestamp 1654583406
transform 1 0 15686 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_811
timestamp 1654583406
transform 1 0 13202 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_812
timestamp 1654583406
transform 1 0 11178 0 1 14042
box -29 -23 29 23
use L1M1_PR  L1M1_PR_813
timestamp 1654583406
transform 1 0 13202 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_814
timestamp 1654583406
transform 1 0 10810 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_815
timestamp 1654583406
transform 1 0 10902 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_816
timestamp 1654583406
transform 1 0 10626 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_817
timestamp 1654583406
transform 1 0 11914 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_818
timestamp 1654583406
transform 1 0 11270 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_819
timestamp 1654583406
transform 1 0 12190 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_820
timestamp 1654583406
transform 1 0 11730 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_821
timestamp 1654583406
transform 1 0 13202 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_822
timestamp 1654583406
transform 1 0 12374 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_823
timestamp 1654583406
transform 1 0 15042 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_824
timestamp 1654583406
transform 1 0 14490 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_825
timestamp 1654583406
transform 1 0 16238 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_826
timestamp 1654583406
transform 1 0 15410 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_827
timestamp 1654583406
transform 1 0 15962 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_828
timestamp 1654583406
transform 1 0 15502 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_829
timestamp 1654583406
transform 1 0 17986 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_830
timestamp 1654583406
transform 1 0 16238 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_831
timestamp 1654583406
transform 1 0 17526 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_832
timestamp 1654583406
transform 1 0 15778 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_833
timestamp 1654583406
transform 1 0 18078 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_834
timestamp 1654583406
transform 1 0 17802 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_835
timestamp 1654583406
transform 1 0 18814 0 1 12614
box -29 -23 29 23
use L1M1_PR  L1M1_PR_836
timestamp 1654583406
transform 1 0 18170 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_837
timestamp 1654583406
transform 1 0 20102 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_838
timestamp 1654583406
transform 1 0 16790 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_839
timestamp 1654583406
transform 1 0 18814 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_840
timestamp 1654583406
transform 1 0 15594 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_841
timestamp 1654583406
transform 1 0 10074 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_842
timestamp 1654583406
transform 1 0 8694 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_843
timestamp 1654583406
transform 1 0 8510 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_844
timestamp 1654583406
transform 1 0 8142 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_845
timestamp 1654583406
transform 1 0 7774 0 1 17996
box -29 -23 29 23
use L1M1_PR  L1M1_PR_846
timestamp 1654583406
transform 1 0 7682 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_847
timestamp 1654583406
transform 1 0 7406 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_848
timestamp 1654583406
transform 1 0 6578 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_849
timestamp 1654583406
transform 1 0 6486 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_850
timestamp 1654583406
transform 1 0 6302 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_851
timestamp 1654583406
transform 1 0 6118 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_852
timestamp 1654583406
transform 1 0 22310 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_853
timestamp 1654583406
transform 1 0 21758 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_854
timestamp 1654583406
transform 1 0 21574 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_855
timestamp 1654583406
transform 1 0 21574 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_856
timestamp 1654583406
transform 1 0 20746 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_857
timestamp 1654583406
transform 1 0 20378 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_858
timestamp 1654583406
transform 1 0 19642 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_859
timestamp 1654583406
transform 1 0 19458 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_860
timestamp 1654583406
transform 1 0 18998 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_861
timestamp 1654583406
transform 1 0 18446 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_862
timestamp 1654583406
transform 1 0 17894 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_863
timestamp 1654583406
transform 1 0 17066 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_864
timestamp 1654583406
transform 1 0 16606 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_865
timestamp 1654583406
transform 1 0 16514 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_866
timestamp 1654583406
transform 1 0 15594 0 1 20162
box -29 -23 29 23
use L1M1_PR  L1M1_PR_867
timestamp 1654583406
transform 1 0 14490 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_868
timestamp 1654583406
transform 1 0 14306 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_869
timestamp 1654583406
transform 1 0 13846 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_870
timestamp 1654583406
transform 1 0 13018 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_871
timestamp 1654583406
transform 1 0 12558 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_872
timestamp 1654583406
transform 1 0 11822 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_873
timestamp 1654583406
transform 1 0 10258 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_874
timestamp 1654583406
transform 1 0 10258 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_875
timestamp 1654583406
transform 1 0 9982 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_876
timestamp 1654583406
transform 1 0 8801 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_877
timestamp 1654583406
transform 1 0 8694 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_878
timestamp 1654583406
transform 1 0 8142 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_879
timestamp 1654583406
transform 1 0 7866 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_880
timestamp 1654583406
transform 1 0 7498 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_881
timestamp 1654583406
transform 1 0 22310 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_882
timestamp 1654583406
transform 1 0 22310 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_883
timestamp 1654583406
transform 1 0 22034 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_884
timestamp 1654583406
transform 1 0 21758 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_885
timestamp 1654583406
transform 1 0 20930 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_886
timestamp 1654583406
transform 1 0 20838 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_887
timestamp 1654583406
transform 1 0 19642 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_888
timestamp 1654583406
transform 1 0 19182 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_889
timestamp 1654583406
transform 1 0 17894 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_890
timestamp 1654583406
transform 1 0 17158 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_891
timestamp 1654583406
transform 1 0 15870 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_892
timestamp 1654583406
transform 1 0 14214 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_893
timestamp 1654583406
transform 1 0 12558 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_894
timestamp 1654583406
transform 1 0 11638 0 1 8670
box -29 -23 29 23
use L1M1_PR  L1M1_PR_895
timestamp 1654583406
transform 1 0 10718 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_896
timestamp 1654583406
transform 1 0 9614 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_897
timestamp 1654583406
transform 1 0 8786 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_898
timestamp 1654583406
transform 1 0 6578 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_899
timestamp 1654583406
transform 1 0 6394 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_900
timestamp 1654583406
transform 1 0 6379 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_901
timestamp 1654583406
transform 1 0 12834 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_902
timestamp 1654583406
transform 1 0 12834 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_903
timestamp 1654583406
transform 1 0 12742 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_904
timestamp 1654583406
transform 1 0 12098 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_905
timestamp 1654583406
transform 1 0 12098 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_906
timestamp 1654583406
transform 1 0 11638 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_907
timestamp 1654583406
transform 1 0 11178 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_908
timestamp 1654583406
transform 1 0 11086 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_909
timestamp 1654583406
transform 1 0 10810 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_910
timestamp 1654583406
transform 1 0 10810 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_911
timestamp 1654583406
transform 1 0 10442 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_912
timestamp 1654583406
transform 1 0 10258 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_913
timestamp 1654583406
transform 1 0 9890 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_914
timestamp 1654583406
transform 1 0 9798 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_915
timestamp 1654583406
transform 1 0 9062 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_916
timestamp 1654583406
transform 1 0 8878 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_917
timestamp 1654583406
transform 1 0 8602 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_918
timestamp 1654583406
transform 1 0 8510 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_919
timestamp 1654583406
transform 1 0 8510 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_920
timestamp 1654583406
transform 1 0 8234 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_921
timestamp 1654583406
transform 1 0 7958 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_922
timestamp 1654583406
transform 1 0 7866 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_923
timestamp 1654583406
transform 1 0 7682 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_924
timestamp 1654583406
transform 1 0 7498 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_925
timestamp 1654583406
transform 1 0 7498 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_926
timestamp 1654583406
transform 1 0 7222 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_927
timestamp 1654583406
transform 1 0 7222 0 1 8670
box -29 -23 29 23
use L1M1_PR  L1M1_PR_928
timestamp 1654583406
transform 1 0 7222 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_929
timestamp 1654583406
transform 1 0 6946 0 1 12546
box -29 -23 29 23
use L1M1_PR  L1M1_PR_930
timestamp 1654583406
transform 1 0 6486 0 1 11458
box -29 -23 29 23
use L1M1_PR  L1M1_PR_931
timestamp 1654583406
transform 1 0 6302 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_932
timestamp 1654583406
transform 1 0 6210 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_933
timestamp 1654583406
transform 1 0 6210 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_934
timestamp 1654583406
transform 1 0 6118 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_935
timestamp 1654583406
transform 1 0 6118 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_936
timestamp 1654583406
transform 1 0 6118 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_937
timestamp 1654583406
transform 1 0 6026 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_938
timestamp 1654583406
transform 1 0 22770 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_939
timestamp 1654583406
transform 1 0 22770 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_940
timestamp 1654583406
transform 1 0 22770 0 1 15810
box -29 -23 29 23
use L1M1_PR  L1M1_PR_941
timestamp 1654583406
transform 1 0 22770 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_942
timestamp 1654583406
transform 1 0 21758 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_943
timestamp 1654583406
transform 1 0 21482 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_944
timestamp 1654583406
transform 1 0 21482 0 1 14110
box -29 -23 29 23
use L1M1_PR  L1M1_PR_945
timestamp 1654583406
transform 1 0 21482 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_946
timestamp 1654583406
transform 1 0 21390 0 1 11458
box -29 -23 29 23
use L1M1_PR  L1M1_PR_947
timestamp 1654583406
transform 1 0 21390 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_948
timestamp 1654583406
transform 1 0 20930 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_949
timestamp 1654583406
transform 1 0 20562 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_950
timestamp 1654583406
transform 1 0 20102 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_951
timestamp 1654583406
transform 1 0 19090 0 1 11458
box -29 -23 29 23
use L1M1_PR  L1M1_PR_952
timestamp 1654583406
transform 1 0 18906 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_953
timestamp 1654583406
transform 1 0 18814 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_954
timestamp 1654583406
transform 1 0 18538 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_955
timestamp 1654583406
transform 1 0 17710 0 1 8670
box -29 -23 29 23
use L1M1_PR  L1M1_PR_956
timestamp 1654583406
transform 1 0 17618 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_957
timestamp 1654583406
transform 1 0 17618 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_958
timestamp 1654583406
transform 1 0 17526 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_959
timestamp 1654583406
transform 1 0 17526 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_960
timestamp 1654583406
transform 1 0 16974 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_961
timestamp 1654583406
transform 1 0 16514 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_962
timestamp 1654583406
transform 1 0 16238 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_963
timestamp 1654583406
transform 1 0 15962 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_964
timestamp 1654583406
transform 1 0 15226 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_965
timestamp 1654583406
transform 1 0 14674 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_966
timestamp 1654583406
transform 1 0 14398 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_967
timestamp 1654583406
transform 1 0 13754 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_968
timestamp 1654583406
transform 1 0 13662 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_969
timestamp 1654583406
transform 1 0 13662 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_970
timestamp 1654583406
transform 1 0 13386 0 1 10438
box -29 -23 29 23
use L1M1_PR  L1M1_PR_971
timestamp 1654583406
transform 1 0 13386 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_972
timestamp 1654583406
transform 1 0 13386 0 1 11866
box -29 -23 29 23
use L1M1_PR  L1M1_PR_973
timestamp 1654583406
transform 1 0 13018 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_974
timestamp 1654583406
transform 1 0 8234 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_975
timestamp 1654583406
transform 1 0 7314 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_976
timestamp 1654583406
transform 1 0 6670 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_977
timestamp 1654583406
transform 1 0 13110 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_978
timestamp 1654583406
transform 1 0 12834 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_979
timestamp 1654583406
transform 1 0 11178 0 1 15062
box -29 -23 29 23
use L1M1_PR  L1M1_PR_980
timestamp 1654583406
transform 1 0 10718 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_981
timestamp 1654583406
transform 1 0 17526 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_982
timestamp 1654583406
transform 1 0 15410 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_983
timestamp 1654583406
transform 1 0 18814 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_984
timestamp 1654583406
transform 1 0 18630 0 1 15810
box -29 -23 29 23
use L1M1_PR  L1M1_PR_985
timestamp 1654583406
transform 1 0 17986 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_986
timestamp 1654583406
transform 1 0 20562 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_987
timestamp 1654583406
transform 1 0 20286 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_988
timestamp 1654583406
transform 1 0 19918 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_989
timestamp 1654583406
transform 1 0 19274 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_990
timestamp 1654583406
transform 1 0 20194 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_991
timestamp 1654583406
transform 1 0 18078 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_992
timestamp 1654583406
transform 1 0 19090 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_993
timestamp 1654583406
transform 1 0 16606 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_994
timestamp 1654583406
transform 1 0 16422 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_995
timestamp 1654583406
transform 1 0 15318 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_996
timestamp 1654583406
transform 1 0 14490 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_997
timestamp 1654583406
transform 1 0 13202 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_998
timestamp 1654583406
transform 1 0 13110 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_999
timestamp 1654583406
transform 1 0 12374 0 1 17578
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1000
timestamp 1654583406
transform 1 0 13662 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1001
timestamp 1654583406
transform 1 0 11638 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1002
timestamp 1654583406
transform 1 0 11086 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1003
timestamp 1654583406
transform 1 0 10534 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1004
timestamp 1654583406
transform 1 0 11914 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1005
timestamp 1654583406
transform 1 0 10902 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1006
timestamp 1654583406
transform 1 0 5842 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1007
timestamp 1654583406
transform 1 0 10534 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1008
timestamp 1654583406
transform 1 0 8970 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1009
timestamp 1654583406
transform 1 0 7205 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1010
timestamp 1654583406
transform 1 0 15318 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1011
timestamp 1654583406
transform 1 0 13202 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1012
timestamp 1654583406
transform 1 0 13110 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1013
timestamp 1654583406
transform 1 0 12006 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1014
timestamp 1654583406
transform 1 0 11546 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1015
timestamp 1654583406
transform 1 0 8694 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1016
timestamp 1654583406
transform 1 0 8479 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1017
timestamp 1654583406
transform 1 0 7498 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1018
timestamp 1654583406
transform 1 0 6762 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1019
timestamp 1654583406
transform 1 0 6302 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1020
timestamp 1654583406
transform 1 0 6578 0 1 15266
box -29 -23 29 23
use M1M2_PR  M1M2_PR_0
timestamp 1654583406
transform 1 0 12926 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1
timestamp 1654583406
transform 1 0 12834 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2
timestamp 1654583406
transform 1 0 10626 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3
timestamp 1654583406
transform 1 0 10626 0 1 14722
box -32 -32 32 32
use M1M2_PR  M1M2_PR_4
timestamp 1654583406
transform 1 0 12466 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_5
timestamp 1654583406
transform 1 0 12466 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_6
timestamp 1654583406
transform 1 0 11086 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_7
timestamp 1654583406
transform 1 0 11086 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_8
timestamp 1654583406
transform 1 0 14306 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_9
timestamp 1654583406
transform 1 0 14306 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_10
timestamp 1654583406
transform 1 0 14766 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_11
timestamp 1654583406
transform 1 0 14766 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_12
timestamp 1654583406
transform 1 0 15594 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_13
timestamp 1654583406
transform 1 0 15410 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_14
timestamp 1654583406
transform 1 0 18722 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_15
timestamp 1654583406
transform 1 0 18722 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_16
timestamp 1654583406
transform 1 0 16422 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_17
timestamp 1654583406
transform 1 0 16422 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_18
timestamp 1654583406
transform 1 0 18630 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_19
timestamp 1654583406
transform 1 0 18630 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_20
timestamp 1654583406
transform 1 0 16698 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_21
timestamp 1654583406
transform 1 0 16606 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_22
timestamp 1654583406
transform 1 0 14674 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_23
timestamp 1654583406
transform 1 0 14030 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_24
timestamp 1654583406
transform 1 0 18906 0 1 15674
box -32 -32 32 32
use M1M2_PR  M1M2_PR_25
timestamp 1654583406
transform 1 0 18906 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_26
timestamp 1654583406
transform 1 0 18170 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_27
timestamp 1654583406
transform 1 0 18170 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_28
timestamp 1654583406
transform 1 0 16514 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_29
timestamp 1654583406
transform 1 0 16514 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_30
timestamp 1654583406
transform 1 0 16146 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_31
timestamp 1654583406
transform 1 0 16146 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_32
timestamp 1654583406
transform 1 0 14306 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_33
timestamp 1654583406
transform 1 0 14306 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_34
timestamp 1654583406
transform 1 0 11454 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_35
timestamp 1654583406
transform 1 0 11454 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_36
timestamp 1654583406
transform 1 0 10534 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_37
timestamp 1654583406
transform 1 0 10534 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_38
timestamp 1654583406
transform 1 0 12006 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_39
timestamp 1654583406
transform 1 0 12006 0 1 15334
box -32 -32 32 32
use M1M2_PR  M1M2_PR_40
timestamp 1654583406
transform 1 0 8234 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_41
timestamp 1654583406
transform 1 0 8234 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_42
timestamp 1654583406
transform 1 0 20654 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_43
timestamp 1654583406
transform 1 0 19182 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_44
timestamp 1654583406
transform 1 0 17894 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_45
timestamp 1654583406
transform 1 0 17894 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_46
timestamp 1654583406
transform 1 0 17802 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_47
timestamp 1654583406
transform 1 0 17802 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_48
timestamp 1654583406
transform 1 0 17802 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_49
timestamp 1654583406
transform 1 0 17802 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_50
timestamp 1654583406
transform 1 0 17710 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_51
timestamp 1654583406
transform 1 0 17710 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_52
timestamp 1654583406
transform 1 0 16698 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_53
timestamp 1654583406
transform 1 0 16698 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_54
timestamp 1654583406
transform 1 0 15870 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_55
timestamp 1654583406
transform 1 0 15686 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_56
timestamp 1654583406
transform 1 0 15686 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_57
timestamp 1654583406
transform 1 0 15594 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_58
timestamp 1654583406
transform 1 0 15594 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_59
timestamp 1654583406
transform 1 0 15226 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_60
timestamp 1654583406
transform 1 0 14950 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_61
timestamp 1654583406
transform 1 0 14950 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_62
timestamp 1654583406
transform 1 0 14582 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_63
timestamp 1654583406
transform 1 0 14398 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_64
timestamp 1654583406
transform 1 0 13294 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_65
timestamp 1654583406
transform 1 0 12006 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_66
timestamp 1654583406
transform 1 0 11822 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_67
timestamp 1654583406
transform 1 0 11822 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_68
timestamp 1654583406
transform 1 0 11730 0 1 18394
box -32 -32 32 32
use M1M2_PR  M1M2_PR_69
timestamp 1654583406
transform 1 0 11730 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_70
timestamp 1654583406
transform 1 0 11730 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_71
timestamp 1654583406
transform 1 0 11730 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_72
timestamp 1654583406
transform 1 0 11730 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_73
timestamp 1654583406
transform 1 0 11546 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_74
timestamp 1654583406
transform 1 0 11546 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_75
timestamp 1654583406
transform 1 0 19642 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_76
timestamp 1654583406
transform 1 0 18354 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_77
timestamp 1654583406
transform 1 0 18354 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_78
timestamp 1654583406
transform 1 0 18354 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_79
timestamp 1654583406
transform 1 0 18262 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_80
timestamp 1654583406
transform 1 0 18262 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_81
timestamp 1654583406
transform 1 0 18262 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_82
timestamp 1654583406
transform 1 0 18262 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_83
timestamp 1654583406
transform 1 0 16422 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_84
timestamp 1654583406
transform 1 0 16422 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_85
timestamp 1654583406
transform 1 0 16422 0 1 12546
box -32 -32 32 32
use M1M2_PR  M1M2_PR_86
timestamp 1654583406
transform 1 0 15870 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_87
timestamp 1654583406
transform 1 0 15870 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_88
timestamp 1654583406
transform 1 0 15870 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_89
timestamp 1654583406
transform 1 0 15778 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_90
timestamp 1654583406
transform 1 0 15686 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_91
timestamp 1654583406
transform 1 0 14398 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_92
timestamp 1654583406
transform 1 0 14214 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_93
timestamp 1654583406
transform 1 0 13662 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_94
timestamp 1654583406
transform 1 0 13662 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_95
timestamp 1654583406
transform 1 0 13386 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_96
timestamp 1654583406
transform 1 0 13386 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_97
timestamp 1654583406
transform 1 0 12742 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_98
timestamp 1654583406
transform 1 0 12742 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_99
timestamp 1654583406
transform 1 0 12282 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_100
timestamp 1654583406
transform 1 0 12190 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_101
timestamp 1654583406
transform 1 0 12190 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_102
timestamp 1654583406
transform 1 0 11638 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_103
timestamp 1654583406
transform 1 0 11638 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_104
timestamp 1654583406
transform 1 0 11546 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_105
timestamp 1654583406
transform 1 0 11546 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_106
timestamp 1654583406
transform 1 0 11546 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_107
timestamp 1654583406
transform 1 0 10350 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_108
timestamp 1654583406
transform 1 0 10350 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_109
timestamp 1654583406
transform 1 0 10350 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_110
timestamp 1654583406
transform 1 0 10350 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_111
timestamp 1654583406
transform 1 0 9154 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_112
timestamp 1654583406
transform 1 0 9154 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_113
timestamp 1654583406
transform 1 0 11178 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_114
timestamp 1654583406
transform 1 0 11178 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_115
timestamp 1654583406
transform 1 0 17342 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_116
timestamp 1654583406
transform 1 0 17342 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_117
timestamp 1654583406
transform 1 0 17250 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_118
timestamp 1654583406
transform 1 0 17250 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_119
timestamp 1654583406
transform 1 0 11546 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_120
timestamp 1654583406
transform 1 0 11546 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_121
timestamp 1654583406
transform 1 0 10902 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_122
timestamp 1654583406
transform 1 0 10902 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_123
timestamp 1654583406
transform 1 0 12006 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_124
timestamp 1654583406
transform 1 0 12006 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_125
timestamp 1654583406
transform 1 0 12926 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_126
timestamp 1654583406
transform 1 0 12926 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_127
timestamp 1654583406
transform 1 0 14582 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_128
timestamp 1654583406
transform 1 0 14582 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_129
timestamp 1654583406
transform 1 0 14490 0 1 18394
box -32 -32 32 32
use M1M2_PR  M1M2_PR_130
timestamp 1654583406
transform 1 0 14490 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_131
timestamp 1654583406
transform 1 0 16974 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_132
timestamp 1654583406
transform 1 0 16974 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_133
timestamp 1654583406
transform 1 0 15962 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_134
timestamp 1654583406
transform 1 0 15962 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_135
timestamp 1654583406
transform 1 0 18998 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_136
timestamp 1654583406
transform 1 0 18998 0 1 17306
box -32 -32 32 32
use M1M2_PR  M1M2_PR_137
timestamp 1654583406
transform 1 0 18814 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_138
timestamp 1654583406
transform 1 0 18814 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_139
timestamp 1654583406
transform 1 0 18906 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_140
timestamp 1654583406
transform 1 0 18906 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_141
timestamp 1654583406
transform 1 0 16422 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_142
timestamp 1654583406
transform 1 0 16422 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_143
timestamp 1654583406
transform 1 0 17250 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_144
timestamp 1654583406
transform 1 0 17250 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_145
timestamp 1654583406
transform 1 0 17894 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_146
timestamp 1654583406
transform 1 0 17894 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_147
timestamp 1654583406
transform 1 0 18078 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_148
timestamp 1654583406
transform 1 0 18078 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_149
timestamp 1654583406
transform 1 0 15502 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_150
timestamp 1654583406
transform 1 0 17710 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_151
timestamp 1654583406
transform 1 0 17710 0 1 12614
box -32 -32 32 32
use M1M2_PR  M1M2_PR_152
timestamp 1654583406
transform 1 0 17618 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_153
timestamp 1654583406
transform 1 0 17618 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_154
timestamp 1654583406
transform 1 0 15870 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_155
timestamp 1654583406
transform 1 0 15778 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_156
timestamp 1654583406
transform 1 0 15870 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_157
timestamp 1654583406
transform 1 0 14766 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_158
timestamp 1654583406
transform 1 0 12650 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_159
timestamp 1654583406
transform 1 0 12650 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_160
timestamp 1654583406
transform 1 0 13570 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_161
timestamp 1654583406
transform 1 0 13386 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_162
timestamp 1654583406
transform 1 0 12190 0 1 13974
box -32 -32 32 32
use M1M2_PR  M1M2_PR_163
timestamp 1654583406
transform 1 0 12190 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_164
timestamp 1654583406
transform 1 0 13478 0 1 16966
box -32 -32 32 32
use M1M2_PR  M1M2_PR_165
timestamp 1654583406
transform 1 0 13478 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_166
timestamp 1654583406
transform 1 0 13478 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_167
timestamp 1654583406
transform 1 0 17158 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_168
timestamp 1654583406
transform 1 0 16882 0 1 16218
box -32 -32 32 32
use M1M2_PR  M1M2_PR_169
timestamp 1654583406
transform 1 0 16882 0 1 15130
box -32 -32 32 32
use M1M2_PR  M1M2_PR_170
timestamp 1654583406
transform 1 0 10442 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_171
timestamp 1654583406
transform 1 0 10442 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_172
timestamp 1654583406
transform 1 0 13294 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_173
timestamp 1654583406
transform 1 0 13202 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_174
timestamp 1654583406
transform 1 0 13110 0 1 17986
box -32 -32 32 32
use M1M2_PR  M1M2_PR_175
timestamp 1654583406
transform 1 0 12190 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_176
timestamp 1654583406
transform 1 0 11086 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_177
timestamp 1654583406
transform 1 0 11086 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_178
timestamp 1654583406
transform 1 0 11086 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_179
timestamp 1654583406
transform 1 0 11086 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_180
timestamp 1654583406
transform 1 0 17618 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_181
timestamp 1654583406
transform 1 0 17618 0 1 14722
box -32 -32 32 32
use M1M2_PR  M1M2_PR_182
timestamp 1654583406
transform 1 0 17618 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_183
timestamp 1654583406
transform 1 0 16054 0 1 16218
box -32 -32 32 32
use M1M2_PR  M1M2_PR_184
timestamp 1654583406
transform 1 0 16054 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_185
timestamp 1654583406
transform 1 0 16054 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_186
timestamp 1654583406
transform 1 0 16054 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_187
timestamp 1654583406
transform 1 0 15042 0 1 15810
box -32 -32 32 32
use M1M2_PR  M1M2_PR_188
timestamp 1654583406
transform 1 0 14766 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_189
timestamp 1654583406
transform 1 0 14766 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_190
timestamp 1654583406
transform 1 0 14766 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_191
timestamp 1654583406
transform 1 0 17526 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_192
timestamp 1654583406
transform 1 0 17526 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_193
timestamp 1654583406
transform 1 0 17526 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_194
timestamp 1654583406
transform 1 0 17526 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_195
timestamp 1654583406
transform 1 0 17526 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_196
timestamp 1654583406
transform 1 0 17434 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_197
timestamp 1654583406
transform 1 0 15042 0 1 17986
box -32 -32 32 32
use M1M2_PR  M1M2_PR_198
timestamp 1654583406
transform 1 0 15042 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_199
timestamp 1654583406
transform 1 0 14766 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_200
timestamp 1654583406
transform 1 0 14766 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_201
timestamp 1654583406
transform 1 0 7958 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_202
timestamp 1654583406
transform 1 0 6578 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_203
timestamp 1654583406
transform 1 0 6578 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_204
timestamp 1654583406
transform 1 0 8326 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_205
timestamp 1654583406
transform 1 0 8326 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_206
timestamp 1654583406
transform 1 0 8786 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_207
timestamp 1654583406
transform 1 0 8786 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_208
timestamp 1654583406
transform 1 0 7866 0 1 21794
box -32 -32 32 32
use M1M2_PR  M1M2_PR_209
timestamp 1654583406
transform 1 0 7866 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_210
timestamp 1654583406
transform 1 0 7406 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_211
timestamp 1654583406
transform 1 0 7406 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_212
timestamp 1654583406
transform 1 0 7406 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_213
timestamp 1654583406
transform 1 0 6670 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_214
timestamp 1654583406
transform 1 0 6670 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_215
timestamp 1654583406
transform 1 0 7866 0 1 16966
box -32 -32 32 32
use M1M2_PR  M1M2_PR_216
timestamp 1654583406
transform 1 0 7866 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_217
timestamp 1654583406
transform 1 0 7130 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_218
timestamp 1654583406
transform 1 0 7038 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_219
timestamp 1654583406
transform 1 0 9062 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_220
timestamp 1654583406
transform 1 0 9062 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_221
timestamp 1654583406
transform 1 0 9062 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_222
timestamp 1654583406
transform 1 0 10258 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_223
timestamp 1654583406
transform 1 0 10258 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_224
timestamp 1654583406
transform 1 0 9798 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_225
timestamp 1654583406
transform 1 0 9798 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_226
timestamp 1654583406
transform 1 0 7958 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_227
timestamp 1654583406
transform 1 0 7130 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_228
timestamp 1654583406
transform 1 0 7130 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_229
timestamp 1654583406
transform 1 0 7038 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_230
timestamp 1654583406
transform 1 0 6854 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_231
timestamp 1654583406
transform 1 0 6210 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_232
timestamp 1654583406
transform 1 0 6210 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_233
timestamp 1654583406
transform 1 0 8878 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_234
timestamp 1654583406
transform 1 0 8878 0 1 20230
box -32 -32 32 32
use M1M2_PR  M1M2_PR_235
timestamp 1654583406
transform 1 0 8878 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_236
timestamp 1654583406
transform 1 0 9246 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_237
timestamp 1654583406
transform 1 0 9154 0 1 20298
box -32 -32 32 32
use M1M2_PR  M1M2_PR_238
timestamp 1654583406
transform 1 0 8050 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_239
timestamp 1654583406
transform 1 0 8050 0 1 20298
box -32 -32 32 32
use M1M2_PR  M1M2_PR_240
timestamp 1654583406
transform 1 0 7682 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_241
timestamp 1654583406
transform 1 0 9154 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_242
timestamp 1654583406
transform 1 0 9154 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_243
timestamp 1654583406
transform 1 0 8878 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_244
timestamp 1654583406
transform 1 0 8878 0 1 16966
box -32 -32 32 32
use M1M2_PR  M1M2_PR_245
timestamp 1654583406
transform 1 0 6394 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_246
timestamp 1654583406
transform 1 0 6394 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_247
timestamp 1654583406
transform 1 0 6394 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_248
timestamp 1654583406
transform 1 0 6394 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_249
timestamp 1654583406
transform 1 0 9062 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_250
timestamp 1654583406
transform 1 0 9062 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_251
timestamp 1654583406
transform 1 0 7498 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_252
timestamp 1654583406
transform 1 0 7498 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_253
timestamp 1654583406
transform 1 0 8694 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_254
timestamp 1654583406
transform 1 0 8694 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_255
timestamp 1654583406
transform 1 0 8234 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_256
timestamp 1654583406
transform 1 0 8234 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_257
timestamp 1654583406
transform 1 0 6394 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_258
timestamp 1654583406
transform 1 0 6394 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_259
timestamp 1654583406
transform 1 0 15778 0 1 14042
box -32 -32 32 32
use M1M2_PR  M1M2_PR_260
timestamp 1654583406
transform 1 0 15686 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_261
timestamp 1654583406
transform 1 0 14766 0 1 14042
box -32 -32 32 32
use M1M2_PR  M1M2_PR_262
timestamp 1654583406
transform 1 0 14766 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_263
timestamp 1654583406
transform 1 0 14030 0 1 18394
box -32 -32 32 32
use M1M2_PR  M1M2_PR_264
timestamp 1654583406
transform 1 0 14030 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_265
timestamp 1654583406
transform 1 0 11178 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_266
timestamp 1654583406
transform 1 0 10166 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_267
timestamp 1654583406
transform 1 0 10166 0 1 15334
box -32 -32 32 32
use M1M2_PR  M1M2_PR_268
timestamp 1654583406
transform 1 0 15594 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_269
timestamp 1654583406
transform 1 0 14582 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_270
timestamp 1654583406
transform 1 0 14582 0 1 12954
box -32 -32 32 32
use M1M2_PR  M1M2_PR_271
timestamp 1654583406
transform 1 0 12650 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_272
timestamp 1654583406
transform 1 0 12650 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_273
timestamp 1654583406
transform 1 0 9154 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_274
timestamp 1654583406
transform 1 0 9154 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_275
timestamp 1654583406
transform 1 0 8694 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_276
timestamp 1654583406
transform 1 0 8602 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_277
timestamp 1654583406
transform 1 0 6854 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_278
timestamp 1654583406
transform 1 0 6854 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_279
timestamp 1654583406
transform 1 0 7222 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_280
timestamp 1654583406
transform 1 0 7222 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_281
timestamp 1654583406
transform 1 0 10442 0 1 18394
box -32 -32 32 32
use M1M2_PR  M1M2_PR_282
timestamp 1654583406
transform 1 0 10442 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_283
timestamp 1654583406
transform 1 0 8694 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_284
timestamp 1654583406
transform 1 0 8694 0 1 16966
box -32 -32 32 32
use M1M2_PR  M1M2_PR_285
timestamp 1654583406
transform 1 0 7130 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_286
timestamp 1654583406
transform 1 0 7130 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_287
timestamp 1654583406
transform 1 0 13662 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_288
timestamp 1654583406
transform 1 0 12834 0 1 12954
box -32 -32 32 32
use M1M2_PR  M1M2_PR_289
timestamp 1654583406
transform 1 0 12650 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_290
timestamp 1654583406
transform 1 0 10810 0 1 13022
box -32 -32 32 32
use M1M2_PR  M1M2_PR_291
timestamp 1654583406
transform 1 0 9982 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_292
timestamp 1654583406
transform 1 0 9890 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_293
timestamp 1654583406
transform 1 0 9890 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_294
timestamp 1654583406
transform 1 0 9522 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_295
timestamp 1654583406
transform 1 0 9522 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_296
timestamp 1654583406
transform 1 0 20194 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_297
timestamp 1654583406
transform 1 0 20194 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_298
timestamp 1654583406
transform 1 0 20194 0 1 12546
box -32 -32 32 32
use M1M2_PR  M1M2_PR_299
timestamp 1654583406
transform 1 0 18906 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_300
timestamp 1654583406
transform 1 0 17342 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_301
timestamp 1654583406
transform 1 0 17066 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_302
timestamp 1654583406
transform 1 0 17066 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_303
timestamp 1654583406
transform 1 0 17066 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_304
timestamp 1654583406
transform 1 0 18814 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_305
timestamp 1654583406
transform 1 0 18814 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_306
timestamp 1654583406
transform 1 0 17710 0 1 19550
box -32 -32 32 32
use M1M2_PR  M1M2_PR_307
timestamp 1654583406
transform 1 0 15042 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_308
timestamp 1654583406
transform 1 0 14766 0 1 19550
box -32 -32 32 32
use M1M2_PR  M1M2_PR_309
timestamp 1654583406
transform 1 0 12926 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_310
timestamp 1654583406
transform 1 0 12834 0 1 18394
box -32 -32 32 32
use M1M2_PR  M1M2_PR_311
timestamp 1654583406
transform 1 0 13386 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_312
timestamp 1654583406
transform 1 0 13386 0 1 21386
box -32 -32 32 32
use M1M2_PR  M1M2_PR_313
timestamp 1654583406
transform 1 0 18262 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_314
timestamp 1654583406
transform 1 0 18262 0 1 20298
box -32 -32 32 32
use M1M2_PR  M1M2_PR_315
timestamp 1654583406
transform 1 0 21298 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_316
timestamp 1654583406
transform 1 0 21298 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_317
timestamp 1654583406
transform 1 0 21114 0 1 19550
box -32 -32 32 32
use M1M2_PR  M1M2_PR_318
timestamp 1654583406
transform 1 0 21114 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_319
timestamp 1654583406
transform 1 0 22034 0 1 18394
box -32 -32 32 32
use M1M2_PR  M1M2_PR_320
timestamp 1654583406
transform 1 0 22034 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_321
timestamp 1654583406
transform 1 0 20378 0 1 16218
box -32 -32 32 32
use M1M2_PR  M1M2_PR_322
timestamp 1654583406
transform 1 0 20378 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_323
timestamp 1654583406
transform 1 0 21666 0 1 13702
box -32 -32 32 32
use M1M2_PR  M1M2_PR_324
timestamp 1654583406
transform 1 0 21666 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_325
timestamp 1654583406
transform 1 0 22034 0 1 12614
box -32 -32 32 32
use M1M2_PR  M1M2_PR_326
timestamp 1654583406
transform 1 0 22034 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_327
timestamp 1654583406
transform 1 0 21298 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_328
timestamp 1654583406
transform 1 0 21298 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_329
timestamp 1654583406
transform 1 0 22126 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_330
timestamp 1654583406
transform 1 0 22126 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_331
timestamp 1654583406
transform 1 0 20286 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_332
timestamp 1654583406
transform 1 0 20286 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_333
timestamp 1654583406
transform 1 0 18354 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_334
timestamp 1654583406
transform 1 0 18354 0 1 7174
box -32 -32 32 32
use M1M2_PR  M1M2_PR_335
timestamp 1654583406
transform 1 0 16422 0 1 9350
box -32 -32 32 32
use M1M2_PR  M1M2_PR_336
timestamp 1654583406
transform 1 0 16422 0 1 8806
box -32 -32 32 32
use M1M2_PR  M1M2_PR_337
timestamp 1654583406
transform 1 0 12190 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_338
timestamp 1654583406
transform 1 0 12190 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_339
timestamp 1654583406
transform 1 0 11730 0 1 10778
box -32 -32 32 32
use M1M2_PR  M1M2_PR_340
timestamp 1654583406
transform 1 0 11730 0 1 10438
box -32 -32 32 32
use M1M2_PR  M1M2_PR_341
timestamp 1654583406
transform 1 0 8970 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_342
timestamp 1654583406
transform 1 0 8970 0 1 10438
box -32 -32 32 32
use M1M2_PR  M1M2_PR_343
timestamp 1654583406
transform 1 0 7958 0 1 13974
box -32 -32 32 32
use M1M2_PR  M1M2_PR_344
timestamp 1654583406
transform 1 0 7958 0 1 10778
box -32 -32 32 32
use M1M2_PR  M1M2_PR_345
timestamp 1654583406
transform 1 0 7222 0 1 14042
box -32 -32 32 32
use M1M2_PR  M1M2_PR_346
timestamp 1654583406
transform 1 0 7222 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_347
timestamp 1654583406
transform 1 0 10442 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_348
timestamp 1654583406
transform 1 0 10442 0 1 19686
box -32 -32 32 32
use M1M2_PR  M1M2_PR_349
timestamp 1654583406
transform 1 0 10534 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_350
timestamp 1654583406
transform 1 0 10534 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_351
timestamp 1654583406
transform 1 0 12006 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_352
timestamp 1654583406
transform 1 0 12006 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_353
timestamp 1654583406
transform 1 0 12190 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_354
timestamp 1654583406
transform 1 0 12190 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_355
timestamp 1654583406
transform 1 0 14674 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_356
timestamp 1654583406
transform 1 0 14674 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_357
timestamp 1654583406
transform 1 0 16238 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_358
timestamp 1654583406
transform 1 0 16238 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_359
timestamp 1654583406
transform 1 0 18814 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_360
timestamp 1654583406
transform 1 0 18814 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_361
timestamp 1654583406
transform 1 0 20286 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_362
timestamp 1654583406
transform 1 0 20286 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_363
timestamp 1654583406
transform 1 0 21942 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_364
timestamp 1654583406
transform 1 0 21942 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_365
timestamp 1654583406
transform 1 0 22402 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_366
timestamp 1654583406
transform 1 0 22402 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_367
timestamp 1654583406
transform 1 0 21942 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_368
timestamp 1654583406
transform 1 0 21942 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_369
timestamp 1654583406
transform 1 0 21390 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_370
timestamp 1654583406
transform 1 0 21206 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_371
timestamp 1654583406
transform 1 0 19918 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_372
timestamp 1654583406
transform 1 0 19918 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_373
timestamp 1654583406
transform 1 0 21114 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_374
timestamp 1654583406
transform 1 0 21022 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_375
timestamp 1654583406
transform 1 0 17250 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_376
timestamp 1654583406
transform 1 0 17250 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_377
timestamp 1654583406
transform 1 0 16146 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_378
timestamp 1654583406
transform 1 0 16054 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_379
timestamp 1654583406
transform 1 0 14490 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_380
timestamp 1654583406
transform 1 0 14490 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_381
timestamp 1654583406
transform 1 0 13570 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_382
timestamp 1654583406
transform 1 0 13570 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_383
timestamp 1654583406
transform 1 0 10442 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_384
timestamp 1654583406
transform 1 0 10442 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_385
timestamp 1654583406
transform 1 0 8510 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_386
timestamp 1654583406
transform 1 0 8510 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_387
timestamp 1654583406
transform 1 0 7958 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_388
timestamp 1654583406
transform 1 0 7958 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_389
timestamp 1654583406
transform 1 0 8970 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_390
timestamp 1654583406
transform 1 0 8970 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_391
timestamp 1654583406
transform 1 0 9246 0 1 21658
box -32 -32 32 32
use M1M2_PR  M1M2_PR_392
timestamp 1654583406
transform 1 0 9246 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_393
timestamp 1654583406
transform 1 0 9982 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_394
timestamp 1654583406
transform 1 0 9982 0 1 21318
box -32 -32 32 32
use M1M2_PR  M1M2_PR_395
timestamp 1654583406
transform 1 0 12098 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_396
timestamp 1654583406
transform 1 0 12098 0 1 21318
box -32 -32 32 32
use M1M2_PR  M1M2_PR_397
timestamp 1654583406
transform 1 0 12650 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_398
timestamp 1654583406
transform 1 0 12650 0 1 20570
box -32 -32 32 32
use M1M2_PR  M1M2_PR_399
timestamp 1654583406
transform 1 0 14398 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_400
timestamp 1654583406
transform 1 0 14398 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_401
timestamp 1654583406
transform 1 0 15686 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_402
timestamp 1654583406
transform 1 0 15686 0 1 20230
box -32 -32 32 32
use M1M2_PR  M1M2_PR_403
timestamp 1654583406
transform 1 0 16974 0 1 21658
box -32 -32 32 32
use M1M2_PR  M1M2_PR_404
timestamp 1654583406
transform 1 0 16974 0 1 21386
box -32 -32 32 32
use M1M2_PR  M1M2_PR_405
timestamp 1654583406
transform 1 0 19918 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_406
timestamp 1654583406
transform 1 0 19918 0 1 20298
box -32 -32 32 32
use M1M2_PR  M1M2_PR_407
timestamp 1654583406
transform 1 0 20194 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_408
timestamp 1654583406
transform 1 0 20102 0 1 21658
box -32 -32 32 32
use M1M2_PR  M1M2_PR_409
timestamp 1654583406
transform 1 0 22310 0 1 20162
box -32 -32 32 32
use M1M2_PR  M1M2_PR_410
timestamp 1654583406
transform 1 0 22310 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_411
timestamp 1654583406
transform 1 0 21298 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_412
timestamp 1654583406
transform 1 0 21298 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_413
timestamp 1654583406
transform 1 0 22218 0 1 9350
box -32 -32 32 32
use M1M2_PR  M1M2_PR_414
timestamp 1654583406
transform 1 0 22218 0 1 9078
box -32 -32 32 32
use M1M2_PR  M1M2_PR_415
timestamp 1654583406
transform 1 0 22954 0 1 8194
box -32 -32 32 32
use M1M2_PR  M1M2_PR_416
timestamp 1654583406
transform 1 0 22862 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_417
timestamp 1654583406
transform 1 0 18538 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_418
timestamp 1654583406
transform 1 0 18538 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_419
timestamp 1654583406
transform 1 0 16974 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_420
timestamp 1654583406
transform 1 0 16882 0 1 11866
box -32 -32 32 32
use M1M2_PR  M1M2_PR_421
timestamp 1654583406
transform 1 0 18262 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_422
timestamp 1654583406
transform 1 0 18262 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_423
timestamp 1654583406
transform 1 0 16330 0 1 11866
box -32 -32 32 32
use M1M2_PR  M1M2_PR_424
timestamp 1654583406
transform 1 0 16330 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_425
timestamp 1654583406
transform 1 0 14766 0 1 10778
box -32 -32 32 32
use M1M2_PR  M1M2_PR_426
timestamp 1654583406
transform 1 0 14766 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_427
timestamp 1654583406
transform 1 0 13018 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_428
timestamp 1654583406
transform 1 0 13018 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_429
timestamp 1654583406
transform 1 0 12374 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_430
timestamp 1654583406
transform 1 0 12282 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_431
timestamp 1654583406
transform 1 0 10074 0 1 10778
box -32 -32 32 32
use M1M2_PR  M1M2_PR_432
timestamp 1654583406
transform 1 0 10074 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_433
timestamp 1654583406
transform 1 0 7498 0 1 11458
box -32 -32 32 32
use M1M2_PR  M1M2_PR_434
timestamp 1654583406
transform 1 0 7498 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_435
timestamp 1654583406
transform 1 0 7958 0 1 14722
box -32 -32 32 32
use M1M2_PR  M1M2_PR_436
timestamp 1654583406
transform 1 0 6578 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_437
timestamp 1654583406
transform 1 0 6578 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_438
timestamp 1654583406
transform 1 0 22586 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_439
timestamp 1654583406
transform 1 0 22494 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_440
timestamp 1654583406
transform 1 0 22494 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_441
timestamp 1654583406
transform 1 0 22770 0 1 14042
box -32 -32 32 32
use M1M2_PR  M1M2_PR_442
timestamp 1654583406
transform 1 0 22770 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_443
timestamp 1654583406
transform 1 0 22770 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_444
timestamp 1654583406
transform 1 0 22494 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_445
timestamp 1654583406
transform 1 0 22494 0 1 11934
box -32 -32 32 32
use M1M2_PR  M1M2_PR_446
timestamp 1654583406
transform 1 0 22494 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_447
timestamp 1654583406
transform 1 0 22678 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_448
timestamp 1654583406
transform 1 0 22678 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_449
timestamp 1654583406
transform 1 0 22586 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_450
timestamp 1654583406
transform 1 0 22310 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_451
timestamp 1654583406
transform 1 0 22310 0 1 6426
box -32 -32 32 32
use M1M2_PR  M1M2_PR_452
timestamp 1654583406
transform 1 0 19642 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_453
timestamp 1654583406
transform 1 0 19642 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_454
timestamp 1654583406
transform 1 0 20286 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_455
timestamp 1654583406
transform 1 0 20286 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_456
timestamp 1654583406
transform 1 0 19734 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_457
timestamp 1654583406
transform 1 0 19734 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_458
timestamp 1654583406
transform 1 0 19366 0 1 6426
box -32 -32 32 32
use M1M2_PR  M1M2_PR_459
timestamp 1654583406
transform 1 0 19366 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_460
timestamp 1654583406
transform 1 0 18354 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_461
timestamp 1654583406
transform 1 0 18354 0 1 5814
box -32 -32 32 32
use M1M2_PR  M1M2_PR_462
timestamp 1654583406
transform 1 0 18538 0 1 6970
box -32 -32 32 32
use M1M2_PR  M1M2_PR_463
timestamp 1654583406
transform 1 0 18538 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_464
timestamp 1654583406
transform 1 0 18538 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_465
timestamp 1654583406
transform 1 0 15502 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_466
timestamp 1654583406
transform 1 0 15410 0 1 6426
box -32 -32 32 32
use M1M2_PR  M1M2_PR_467
timestamp 1654583406
transform 1 0 14398 0 1 8262
box -32 -32 32 32
use M1M2_PR  M1M2_PR_468
timestamp 1654583406
transform 1 0 14398 0 1 7718
box -32 -32 32 32
use M1M2_PR  M1M2_PR_469
timestamp 1654583406
transform 1 0 10534 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_470
timestamp 1654583406
transform 1 0 10442 0 1 8534
box -32 -32 32 32
use M1M2_PR  M1M2_PR_471
timestamp 1654583406
transform 1 0 10258 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_472
timestamp 1654583406
transform 1 0 10258 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_473
timestamp 1654583406
transform 1 0 9062 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_474
timestamp 1654583406
transform 1 0 9062 0 1 8262
box -32 -32 32 32
use M1M2_PR  M1M2_PR_475
timestamp 1654583406
transform 1 0 7130 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_476
timestamp 1654583406
transform 1 0 7130 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_477
timestamp 1654583406
transform 1 0 6578 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_478
timestamp 1654583406
transform 1 0 6578 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_479
timestamp 1654583406
transform 1 0 7958 0 1 8806
box -32 -32 32 32
use M1M2_PR  M1M2_PR_480
timestamp 1654583406
transform 1 0 11270 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_481
timestamp 1654583406
transform 1 0 11270 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_482
timestamp 1654583406
transform 1 0 10902 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_483
timestamp 1654583406
transform 1 0 10902 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_484
timestamp 1654583406
transform 1 0 12374 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_485
timestamp 1654583406
transform 1 0 12374 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_486
timestamp 1654583406
transform 1 0 14490 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_487
timestamp 1654583406
transform 1 0 14490 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_488
timestamp 1654583406
transform 1 0 16054 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_489
timestamp 1654583406
transform 1 0 16054 0 1 7718
box -32 -32 32 32
use M1M2_PR  M1M2_PR_490
timestamp 1654583406
transform 1 0 18078 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_491
timestamp 1654583406
transform 1 0 18078 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_492
timestamp 1654583406
transform 1 0 17066 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_493
timestamp 1654583406
transform 1 0 17066 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_494
timestamp 1654583406
transform 1 0 18538 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_495
timestamp 1654583406
transform 1 0 18538 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_496
timestamp 1654583406
transform 1 0 19918 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_497
timestamp 1654583406
transform 1 0 19918 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_498
timestamp 1654583406
transform 1 0 21022 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_499
timestamp 1654583406
transform 1 0 21022 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_500
timestamp 1654583406
transform 1 0 21666 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_501
timestamp 1654583406
transform 1 0 21666 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_502
timestamp 1654583406
transform 1 0 21390 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_503
timestamp 1654583406
transform 1 0 21390 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_504
timestamp 1654583406
transform 1 0 21850 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_505
timestamp 1654583406
transform 1 0 21850 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_506
timestamp 1654583406
transform 1 0 22218 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_507
timestamp 1654583406
transform 1 0 22218 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_508
timestamp 1654583406
transform 1 0 21942 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_509
timestamp 1654583406
transform 1 0 21942 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_510
timestamp 1654583406
transform 1 0 21114 0 1 13974
box -32 -32 32 32
use M1M2_PR  M1M2_PR_511
timestamp 1654583406
transform 1 0 21114 0 1 13702
box -32 -32 32 32
use M1M2_PR  M1M2_PR_512
timestamp 1654583406
transform 1 0 22494 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_513
timestamp 1654583406
transform 1 0 22494 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_514
timestamp 1654583406
transform 1 0 21666 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_515
timestamp 1654583406
transform 1 0 21666 0 1 8262
box -32 -32 32 32
use M1M2_PR  M1M2_PR_516
timestamp 1654583406
transform 1 0 19918 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_517
timestamp 1654583406
transform 1 0 19918 0 1 6426
box -32 -32 32 32
use M1M2_PR  M1M2_PR_518
timestamp 1654583406
transform 1 0 20102 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_519
timestamp 1654583406
transform 1 0 20102 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_520
timestamp 1654583406
transform 1 0 17342 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_521
timestamp 1654583406
transform 1 0 17342 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_522
timestamp 1654583406
transform 1 0 17710 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_523
timestamp 1654583406
transform 1 0 17710 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_524
timestamp 1654583406
transform 1 0 15686 0 1 8194
box -32 -32 32 32
use M1M2_PR  M1M2_PR_525
timestamp 1654583406
transform 1 0 15686 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_526
timestamp 1654583406
transform 1 0 14306 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_527
timestamp 1654583406
transform 1 0 14306 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_528
timestamp 1654583406
transform 1 0 10626 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_529
timestamp 1654583406
transform 1 0 10626 0 1 7718
box -32 -32 32 32
use M1M2_PR  M1M2_PR_530
timestamp 1654583406
transform 1 0 8694 0 1 9350
box -32 -32 32 32
use M1M2_PR  M1M2_PR_531
timestamp 1654583406
transform 1 0 8602 0 1 8194
box -32 -32 32 32
use M1M2_PR  M1M2_PR_532
timestamp 1654583406
transform 1 0 14490 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_533
timestamp 1654583406
transform 1 0 13018 0 1 6970
box -32 -32 32 32
use M1M2_PR  M1M2_PR_534
timestamp 1654583406
transform 1 0 12558 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_535
timestamp 1654583406
transform 1 0 12558 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_536
timestamp 1654583406
transform 1 0 12558 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_537
timestamp 1654583406
transform 1 0 10626 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_538
timestamp 1654583406
transform 1 0 10626 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_539
timestamp 1654583406
transform 1 0 10350 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_540
timestamp 1654583406
transform 1 0 10350 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_541
timestamp 1654583406
transform 1 0 10350 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_542
timestamp 1654583406
transform 1 0 10442 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_543
timestamp 1654583406
transform 1 0 10442 0 1 5882
box -32 -32 32 32
use M1M2_PR  M1M2_PR_544
timestamp 1654583406
transform 1 0 8142 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_545
timestamp 1654583406
transform 1 0 7958 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_546
timestamp 1654583406
transform 1 0 7958 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_547
timestamp 1654583406
transform 1 0 6762 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_548
timestamp 1654583406
transform 1 0 6762 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_549
timestamp 1654583406
transform 1 0 7038 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_550
timestamp 1654583406
transform 1 0 7038 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_551
timestamp 1654583406
transform 1 0 6762 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_552
timestamp 1654583406
transform 1 0 6762 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_553
timestamp 1654583406
transform 1 0 7314 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_554
timestamp 1654583406
transform 1 0 7314 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_555
timestamp 1654583406
transform 1 0 8786 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_556
timestamp 1654583406
transform 1 0 8786 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_557
timestamp 1654583406
transform 1 0 11086 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_558
timestamp 1654583406
transform 1 0 11086 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_559
timestamp 1654583406
transform 1 0 11638 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_560
timestamp 1654583406
transform 1 0 11638 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_561
timestamp 1654583406
transform 1 0 13110 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_562
timestamp 1654583406
transform 1 0 13018 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_563
timestamp 1654583406
transform 1 0 15502 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_564
timestamp 1654583406
transform 1 0 12834 0 1 7174
box -32 -32 32 32
use M1M2_PR  M1M2_PR_565
timestamp 1654583406
transform 1 0 12834 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_566
timestamp 1654583406
transform 1 0 7866 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_567
timestamp 1654583406
transform 1 0 7866 0 1 6426
box -32 -32 32 32
use M1M2_PR  M1M2_PR_568
timestamp 1654583406
transform 1 0 6578 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_569
timestamp 1654583406
transform 1 0 6578 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_570
timestamp 1654583406
transform 1 0 10166 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_571
timestamp 1654583406
transform 1 0 10166 0 1 14246
box -32 -32 32 32
use M1M2_PR  M1M2_PR_572
timestamp 1654583406
transform 1 0 6670 0 1 13022
box -32 -32 32 32
use M1M2_PR  M1M2_PR_573
timestamp 1654583406
transform 1 0 9154 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_574
timestamp 1654583406
transform 1 0 9154 0 1 15674
box -32 -32 32 32
use M1M2_PR  M1M2_PR_575
timestamp 1654583406
transform 1 0 9154 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_576
timestamp 1654583406
transform 1 0 8878 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_577
timestamp 1654583406
transform 1 0 8878 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_578
timestamp 1654583406
transform 1 0 8878 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_579
timestamp 1654583406
transform 1 0 9062 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_580
timestamp 1654583406
transform 1 0 9062 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_581
timestamp 1654583406
transform 1 0 9062 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_582
timestamp 1654583406
transform 1 0 11086 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_583
timestamp 1654583406
transform 1 0 11086 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_584
timestamp 1654583406
transform 1 0 10994 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_585
timestamp 1654583406
transform 1 0 12926 0 1 9894
box -32 -32 32 32
use M1M2_PR  M1M2_PR_586
timestamp 1654583406
transform 1 0 12650 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_587
timestamp 1654583406
transform 1 0 12374 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_588
timestamp 1654583406
transform 1 0 15502 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_589
timestamp 1654583406
transform 1 0 14582 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_590
timestamp 1654583406
transform 1 0 14582 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_591
timestamp 1654583406
transform 1 0 16514 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_592
timestamp 1654583406
transform 1 0 16514 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_593
timestamp 1654583406
transform 1 0 16514 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_594
timestamp 1654583406
transform 1 0 19182 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_595
timestamp 1654583406
transform 1 0 16974 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_596
timestamp 1654583406
transform 1 0 16974 0 1 9894
box -32 -32 32 32
use M1M2_PR  M1M2_PR_597
timestamp 1654583406
transform 1 0 18722 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_598
timestamp 1654583406
transform 1 0 18722 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_599
timestamp 1654583406
transform 1 0 17986 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_600
timestamp 1654583406
transform 1 0 17986 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_601
timestamp 1654583406
transform 1 0 19918 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_602
timestamp 1654583406
transform 1 0 19918 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_603
timestamp 1654583406
transform 1 0 19918 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_604
timestamp 1654583406
transform 1 0 21482 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_605
timestamp 1654583406
transform 1 0 21482 0 1 8194
box -32 -32 32 32
use M1M2_PR  M1M2_PR_606
timestamp 1654583406
transform 1 0 18906 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_607
timestamp 1654583406
transform 1 0 18906 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_608
timestamp 1654583406
transform 1 0 22310 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_609
timestamp 1654583406
transform 1 0 22310 0 1 9350
box -32 -32 32 32
use M1M2_PR  M1M2_PR_610
timestamp 1654583406
transform 1 0 20010 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_611
timestamp 1654583406
transform 1 0 19918 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_612
timestamp 1654583406
transform 1 0 20470 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_613
timestamp 1654583406
transform 1 0 20470 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_614
timestamp 1654583406
transform 1 0 20378 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_615
timestamp 1654583406
transform 1 0 20010 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_616
timestamp 1654583406
transform 1 0 20010 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_617
timestamp 1654583406
transform 1 0 19918 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_618
timestamp 1654583406
transform 1 0 22402 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_619
timestamp 1654583406
transform 1 0 22310 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_620
timestamp 1654583406
transform 1 0 18998 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_621
timestamp 1654583406
transform 1 0 18998 0 1 14246
box -32 -32 32 32
use M1M2_PR  M1M2_PR_622
timestamp 1654583406
transform 1 0 21114 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_623
timestamp 1654583406
transform 1 0 21114 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_624
timestamp 1654583406
transform 1 0 19918 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_625
timestamp 1654583406
transform 1 0 19918 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_626
timestamp 1654583406
transform 1 0 21298 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_627
timestamp 1654583406
transform 1 0 21114 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_628
timestamp 1654583406
transform 1 0 21114 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_629
timestamp 1654583406
transform 1 0 21758 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_630
timestamp 1654583406
transform 1 0 21758 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_631
timestamp 1654583406
transform 1 0 19918 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_632
timestamp 1654583406
transform 1 0 19090 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_633
timestamp 1654583406
transform 1 0 18722 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_634
timestamp 1654583406
transform 1 0 18722 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_635
timestamp 1654583406
transform 1 0 18722 0 1 18938
box -32 -32 32 32
use M1M2_PR  M1M2_PR_636
timestamp 1654583406
transform 1 0 17434 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_637
timestamp 1654583406
transform 1 0 17434 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_638
timestamp 1654583406
transform 1 0 17434 0 1 19686
box -32 -32 32 32
use M1M2_PR  M1M2_PR_639
timestamp 1654583406
transform 1 0 15870 0 1 21114
box -32 -32 32 32
use M1M2_PR  M1M2_PR_640
timestamp 1654583406
transform 1 0 15870 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_641
timestamp 1654583406
transform 1 0 15870 0 1 19686
box -32 -32 32 32
use M1M2_PR  M1M2_PR_642
timestamp 1654583406
transform 1 0 14306 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_643
timestamp 1654583406
transform 1 0 14306 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_644
timestamp 1654583406
transform 1 0 14306 0 1 19686
box -32 -32 32 32
use M1M2_PR  M1M2_PR_645
timestamp 1654583406
transform 1 0 13478 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_646
timestamp 1654583406
transform 1 0 13478 0 1 20298
box -32 -32 32 32
use M1M2_PR  M1M2_PR_647
timestamp 1654583406
transform 1 0 13478 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_648
timestamp 1654583406
transform 1 0 14490 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_649
timestamp 1654583406
transform 1 0 14490 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_650
timestamp 1654583406
transform 1 0 11822 0 1 21794
box -32 -32 32 32
use M1M2_PR  M1M2_PR_651
timestamp 1654583406
transform 1 0 11822 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_652
timestamp 1654583406
transform 1 0 11822 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_653
timestamp 1654583406
transform 1 0 11822 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_654
timestamp 1654583406
transform 1 0 11638 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_655
timestamp 1654583406
transform 1 0 11638 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_656
timestamp 1654583406
transform 1 0 10074 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_657
timestamp 1654583406
transform 1 0 10074 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_658
timestamp 1654583406
transform 1 0 10074 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_659
timestamp 1654583406
transform 1 0 6486 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_660
timestamp 1654583406
transform 1 0 6486 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_661
timestamp 1654583406
transform 1 0 6486 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_662
timestamp 1654583406
transform 1 0 7682 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_663
timestamp 1654583406
transform 1 0 7682 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_664
timestamp 1654583406
transform 1 0 7590 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_665
timestamp 1654583406
transform 1 0 8878 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_666
timestamp 1654583406
transform 1 0 8878 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_667
timestamp 1654583406
transform 1 0 8694 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_668
timestamp 1654583406
transform 1 0 9246 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_669
timestamp 1654583406
transform 1 0 9154 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_670
timestamp 1654583406
transform 1 0 9154 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_671
timestamp 1654583406
transform 1 0 11638 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_672
timestamp 1654583406
transform 1 0 11638 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_673
timestamp 1654583406
transform 1 0 9982 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_674
timestamp 1654583406
transform 1 0 9982 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_675
timestamp 1654583406
transform 1 0 13478 0 1 9078
box -32 -32 32 32
use M1M2_PR  M1M2_PR_676
timestamp 1654583406
transform 1 0 13478 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_677
timestamp 1654583406
transform 1 0 13478 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_678
timestamp 1654583406
transform 1 0 15778 0 1 9078
box -32 -32 32 32
use M1M2_PR  M1M2_PR_679
timestamp 1654583406
transform 1 0 15686 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_680
timestamp 1654583406
transform 1 0 14766 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_681
timestamp 1654583406
transform 1 0 14766 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_682
timestamp 1654583406
transform 1 0 16146 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_683
timestamp 1654583406
transform 1 0 15870 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_684
timestamp 1654583406
transform 1 0 15870 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_685
timestamp 1654583406
transform 1 0 18170 0 1 9078
box -32 -32 32 32
use M1M2_PR  M1M2_PR_686
timestamp 1654583406
transform 1 0 18170 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_687
timestamp 1654583406
transform 1 0 18170 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_688
timestamp 1654583406
transform 1 0 18906 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_689
timestamp 1654583406
transform 1 0 18906 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_690
timestamp 1654583406
transform 1 0 18906 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_691
timestamp 1654583406
transform 1 0 18906 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_692
timestamp 1654583406
transform 1 0 18814 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_693
timestamp 1654583406
transform 1 0 19458 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_694
timestamp 1654583406
transform 1 0 19458 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_695
timestamp 1654583406
transform 1 0 19090 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_696
timestamp 1654583406
transform 1 0 21298 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_697
timestamp 1654583406
transform 1 0 21298 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_698
timestamp 1654583406
transform 1 0 22494 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_699
timestamp 1654583406
transform 1 0 22494 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_700
timestamp 1654583406
transform 1 0 22586 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_701
timestamp 1654583406
transform 1 0 22586 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_702
timestamp 1654583406
transform 1 0 21666 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_703
timestamp 1654583406
transform 1 0 21666 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_704
timestamp 1654583406
transform 1 0 21850 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_705
timestamp 1654583406
transform 1 0 21758 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_706
timestamp 1654583406
transform 1 0 22310 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_707
timestamp 1654583406
transform 1 0 22310 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_708
timestamp 1654583406
transform 1 0 21298 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_709
timestamp 1654583406
transform 1 0 21298 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_710
timestamp 1654583406
transform 1 0 22310 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_711
timestamp 1654583406
transform 1 0 22218 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_712
timestamp 1654583406
transform 1 0 6118 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_713
timestamp 1654583406
transform 1 0 6118 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_714
timestamp 1654583406
transform 1 0 6118 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_715
timestamp 1654583406
transform 1 0 6118 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_716
timestamp 1654583406
transform 1 0 6118 0 1 5882
box -32 -32 32 32
use M1M2_PR  M1M2_PR_717
timestamp 1654583406
transform 1 0 7590 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_718
timestamp 1654583406
transform 1 0 7590 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_719
timestamp 1654583406
transform 1 0 6946 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_720
timestamp 1654583406
transform 1 0 6946 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_721
timestamp 1654583406
transform 1 0 6946 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_722
timestamp 1654583406
transform 1 0 7866 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_723
timestamp 1654583406
transform 1 0 7866 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_724
timestamp 1654583406
transform 1 0 10166 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_725
timestamp 1654583406
transform 1 0 9982 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_726
timestamp 1654583406
transform 1 0 9982 0 1 6086
box -32 -32 32 32
use M1M2_PR  M1M2_PR_727
timestamp 1654583406
transform 1 0 12006 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_728
timestamp 1654583406
transform 1 0 12006 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_729
timestamp 1654583406
transform 1 0 12926 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_730
timestamp 1654583406
transform 1 0 12742 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_731
timestamp 1654583406
transform 1 0 12742 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_732
timestamp 1654583406
transform 1 0 12742 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_733
timestamp 1654583406
transform 1 0 14306 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_734
timestamp 1654583406
transform 1 0 14306 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_735
timestamp 1654583406
transform 1 0 14214 0 1 8194
box -32 -32 32 32
use M1M2_PR  M1M2_PR_736
timestamp 1654583406
transform 1 0 14766 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_737
timestamp 1654583406
transform 1 0 14766 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_738
timestamp 1654583406
transform 1 0 14766 0 1 6086
box -32 -32 32 32
use M1M2_PR  M1M2_PR_739
timestamp 1654583406
transform 1 0 17618 0 1 7174
box -32 -32 32 32
use M1M2_PR  M1M2_PR_740
timestamp 1654583406
transform 1 0 17618 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_741
timestamp 1654583406
transform 1 0 17618 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_742
timestamp 1654583406
transform 1 0 12834 0 1 14722
box -32 -32 32 32
use M1M2_PR  M1M2_PR_743
timestamp 1654583406
transform 1 0 12834 0 1 14042
box -32 -32 32 32
use M1M2_PR  M1M2_PR_744
timestamp 1654583406
transform 1 0 12650 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_745
timestamp 1654583406
transform 1 0 12650 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_746
timestamp 1654583406
transform 1 0 10718 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_747
timestamp 1654583406
transform 1 0 10718 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_748
timestamp 1654583406
transform 1 0 11914 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_749
timestamp 1654583406
transform 1 0 11914 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_750
timestamp 1654583406
transform 1 0 12098 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_751
timestamp 1654583406
transform 1 0 12098 0 1 12614
box -32 -32 32 32
use M1M2_PR  M1M2_PR_752
timestamp 1654583406
transform 1 0 12558 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_753
timestamp 1654583406
transform 1 0 12466 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_754
timestamp 1654583406
transform 1 0 14582 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_755
timestamp 1654583406
transform 1 0 14490 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_756
timestamp 1654583406
transform 1 0 15962 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_757
timestamp 1654583406
transform 1 0 15962 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_758
timestamp 1654583406
transform 1 0 16698 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_759
timestamp 1654583406
transform 1 0 16606 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_760
timestamp 1654583406
transform 1 0 18078 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_761
timestamp 1654583406
transform 1 0 18078 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_762
timestamp 1654583406
transform 1 0 18170 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_763
timestamp 1654583406
transform 1 0 18170 0 1 12614
box -32 -32 32 32
use M1M2_PR  M1M2_PR_764
timestamp 1654583406
transform 1 0 8786 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_765
timestamp 1654583406
transform 1 0 8786 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_766
timestamp 1654583406
transform 1 0 8510 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_767
timestamp 1654583406
transform 1 0 8510 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_768
timestamp 1654583406
transform 1 0 7682 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_769
timestamp 1654583406
transform 1 0 7682 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_770
timestamp 1654583406
transform 1 0 7590 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_771
timestamp 1654583406
transform 1 0 6302 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_772
timestamp 1654583406
transform 1 0 6302 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_773
timestamp 1654583406
transform 1 0 6302 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_774
timestamp 1654583406
transform 1 0 5934 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_775
timestamp 1654583406
transform 1 0 5934 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_776
timestamp 1654583406
transform 1 0 5934 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_777
timestamp 1654583406
transform 1 0 22126 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_778
timestamp 1654583406
transform 1 0 21666 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_779
timestamp 1654583406
transform 1 0 21574 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_780
timestamp 1654583406
transform 1 0 21574 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_781
timestamp 1654583406
transform 1 0 20286 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_782
timestamp 1654583406
transform 1 0 20286 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_783
timestamp 1654583406
transform 1 0 20286 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_784
timestamp 1654583406
transform 1 0 19734 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_785
timestamp 1654583406
transform 1 0 19734 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_786
timestamp 1654583406
transform 1 0 19090 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_787
timestamp 1654583406
transform 1 0 19090 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_788
timestamp 1654583406
transform 1 0 17894 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_789
timestamp 1654583406
transform 1 0 17894 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_790
timestamp 1654583406
transform 1 0 17618 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_791
timestamp 1654583406
transform 1 0 17526 0 1 11866
box -32 -32 32 32
use M1M2_PR  M1M2_PR_792
timestamp 1654583406
transform 1 0 15502 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_793
timestamp 1654583406
transform 1 0 15502 0 1 21318
box -32 -32 32 32
use M1M2_PR  M1M2_PR_794
timestamp 1654583406
transform 1 0 15502 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_795
timestamp 1654583406
transform 1 0 15502 0 1 20162
box -32 -32 32 32
use M1M2_PR  M1M2_PR_796
timestamp 1654583406
transform 1 0 13846 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_797
timestamp 1654583406
transform 1 0 13846 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_798
timestamp 1654583406
transform 1 0 13018 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_799
timestamp 1654583406
transform 1 0 12190 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_800
timestamp 1654583406
transform 1 0 12190 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_801
timestamp 1654583406
transform 1 0 10258 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_802
timestamp 1654583406
transform 1 0 9890 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_803
timestamp 1654583406
transform 1 0 9890 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_804
timestamp 1654583406
transform 1 0 9246 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_805
timestamp 1654583406
transform 1 0 9246 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_806
timestamp 1654583406
transform 1 0 8694 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_807
timestamp 1654583406
transform 1 0 8694 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_808
timestamp 1654583406
transform 1 0 7774 0 1 15130
box -32 -32 32 32
use M1M2_PR  M1M2_PR_809
timestamp 1654583406
transform 1 0 7774 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_810
timestamp 1654583406
transform 1 0 7774 0 1 13702
box -32 -32 32 32
use M1M2_PR  M1M2_PR_811
timestamp 1654583406
transform 1 0 22770 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_812
timestamp 1654583406
transform 1 0 22494 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_813
timestamp 1654583406
transform 1 0 22494 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_814
timestamp 1654583406
transform 1 0 22402 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_815
timestamp 1654583406
transform 1 0 21850 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_816
timestamp 1654583406
transform 1 0 21850 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_817
timestamp 1654583406
transform 1 0 21114 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_818
timestamp 1654583406
transform 1 0 21114 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_819
timestamp 1654583406
transform 1 0 20470 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_820
timestamp 1654583406
transform 1 0 20470 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_821
timestamp 1654583406
transform 1 0 17894 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_822
timestamp 1654583406
transform 1 0 17894 0 1 7718
box -32 -32 32 32
use M1M2_PR  M1M2_PR_823
timestamp 1654583406
transform 1 0 17894 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_824
timestamp 1654583406
transform 1 0 17710 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_825
timestamp 1654583406
transform 1 0 15962 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_826
timestamp 1654583406
transform 1 0 12282 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_827
timestamp 1654583406
transform 1 0 12282 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_828
timestamp 1654583406
transform 1 0 12098 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_829
timestamp 1654583406
transform 1 0 12006 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_830
timestamp 1654583406
transform 1 0 10810 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_831
timestamp 1654583406
transform 1 0 10810 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_832
timestamp 1654583406
transform 1 0 7314 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_833
timestamp 1654583406
transform 1 0 7314 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_834
timestamp 1654583406
transform 1 0 6394 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_835
timestamp 1654583406
transform 1 0 6394 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_836
timestamp 1654583406
transform 1 0 6302 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_837
timestamp 1654583406
transform 1 0 12834 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_838
timestamp 1654583406
transform 1 0 12834 0 1 8194
box -32 -32 32 32
use M1M2_PR  M1M2_PR_839
timestamp 1654583406
transform 1 0 12650 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_840
timestamp 1654583406
transform 1 0 12098 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_841
timestamp 1654583406
transform 1 0 11638 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_842
timestamp 1654583406
transform 1 0 11638 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_843
timestamp 1654583406
transform 1 0 11178 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_844
timestamp 1654583406
transform 1 0 10902 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_845
timestamp 1654583406
transform 1 0 10810 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_846
timestamp 1654583406
transform 1 0 10810 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_847
timestamp 1654583406
transform 1 0 10442 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_848
timestamp 1654583406
transform 1 0 10258 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_849
timestamp 1654583406
transform 1 0 10258 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_850
timestamp 1654583406
transform 1 0 9798 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_851
timestamp 1654583406
transform 1 0 8970 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_852
timestamp 1654583406
transform 1 0 8878 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_853
timestamp 1654583406
transform 1 0 8694 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_854
timestamp 1654583406
transform 1 0 8510 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_855
timestamp 1654583406
transform 1 0 8510 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_856
timestamp 1654583406
transform 1 0 8234 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_857
timestamp 1654583406
transform 1 0 7958 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_858
timestamp 1654583406
transform 1 0 7774 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_859
timestamp 1654583406
transform 1 0 7774 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_860
timestamp 1654583406
transform 1 0 7774 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_861
timestamp 1654583406
transform 1 0 7498 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_862
timestamp 1654583406
transform 1 0 7222 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_863
timestamp 1654583406
transform 1 0 7222 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_864
timestamp 1654583406
transform 1 0 6946 0 1 13022
box -32 -32 32 32
use M1M2_PR  M1M2_PR_865
timestamp 1654583406
transform 1 0 6210 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_866
timestamp 1654583406
transform 1 0 6210 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_867
timestamp 1654583406
transform 1 0 6118 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_868
timestamp 1654583406
transform 1 0 6118 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_869
timestamp 1654583406
transform 1 0 6118 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_870
timestamp 1654583406
transform 1 0 6118 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_871
timestamp 1654583406
transform 1 0 6118 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_872
timestamp 1654583406
transform 1 0 6118 0 1 11458
box -32 -32 32 32
use M1M2_PR  M1M2_PR_873
timestamp 1654583406
transform 1 0 22770 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_874
timestamp 1654583406
transform 1 0 22770 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_875
timestamp 1654583406
transform 1 0 21482 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_876
timestamp 1654583406
transform 1 0 21482 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_877
timestamp 1654583406
transform 1 0 21482 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_878
timestamp 1654583406
transform 1 0 21482 0 1 11934
box -32 -32 32 32
use M1M2_PR  M1M2_PR_879
timestamp 1654583406
transform 1 0 21482 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_880
timestamp 1654583406
transform 1 0 21390 0 1 11458
box -32 -32 32 32
use M1M2_PR  M1M2_PR_881
timestamp 1654583406
transform 1 0 20378 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_882
timestamp 1654583406
transform 1 0 20102 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_883
timestamp 1654583406
transform 1 0 19090 0 1 11458
box -32 -32 32 32
use M1M2_PR  M1M2_PR_884
timestamp 1654583406
transform 1 0 19090 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_885
timestamp 1654583406
transform 1 0 18906 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_886
timestamp 1654583406
transform 1 0 18906 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_887
timestamp 1654583406
transform 1 0 18538 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_888
timestamp 1654583406
transform 1 0 17710 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_889
timestamp 1654583406
transform 1 0 17710 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_890
timestamp 1654583406
transform 1 0 17618 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_891
timestamp 1654583406
transform 1 0 17618 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_892
timestamp 1654583406
transform 1 0 17618 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_893
timestamp 1654583406
transform 1 0 16514 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_894
timestamp 1654583406
transform 1 0 16514 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_895
timestamp 1654583406
transform 1 0 16514 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_896
timestamp 1654583406
transform 1 0 15962 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_897
timestamp 1654583406
transform 1 0 15226 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_898
timestamp 1654583406
transform 1 0 14674 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_899
timestamp 1654583406
transform 1 0 13754 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_900
timestamp 1654583406
transform 1 0 13386 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_901
timestamp 1654583406
transform 1 0 13386 0 1 10438
box -32 -32 32 32
use M1M2_PR  M1M2_PR_902
timestamp 1654583406
transform 1 0 13386 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_903
timestamp 1654583406
transform 1 0 13386 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_904
timestamp 1654583406
transform 1 0 13294 0 1 11866
box -32 -32 32 32
use M1M2_PR  M1M2_PR_905
timestamp 1654583406
transform 1 0 13202 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_906
timestamp 1654583406
transform 1 0 13202 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_907
timestamp 1654583406
transform 1 0 13018 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_908
timestamp 1654583406
transform 1 0 13018 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_909
timestamp 1654583406
transform 1 0 13018 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_910
timestamp 1654583406
transform 1 0 13018 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_911
timestamp 1654583406
transform 1 0 13018 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_912
timestamp 1654583406
transform 1 0 8326 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_913
timestamp 1654583406
transform 1 0 7038 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_914
timestamp 1654583406
transform 1 0 13110 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_915
timestamp 1654583406
transform 1 0 13110 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_916
timestamp 1654583406
transform 1 0 10902 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_917
timestamp 1654583406
transform 1 0 10902 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_918
timestamp 1654583406
transform 1 0 17434 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_919
timestamp 1654583406
transform 1 0 16238 0 1 15810
box -32 -32 32 32
use M1M2_PR  M1M2_PR_920
timestamp 1654583406
transform 1 0 16238 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_921
timestamp 1654583406
transform 1 0 22954 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_922
timestamp 1654583406
transform 1 0 28566 0 1 16966
box -32 -32 32 32
use M1M2_PR  M1M2_PR_923
timestamp 1654583406
transform 1 0 20378 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_924
timestamp 1654583406
transform 1 0 20378 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_925
timestamp 1654583406
transform 1 0 19918 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_926
timestamp 1654583406
transform 1 0 19918 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_927
timestamp 1654583406
transform 1 0 22126 0 1 18938
box -32 -32 32 32
use M1M2_PR  M1M2_PR_928
timestamp 1654583406
transform 1 0 18446 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_929
timestamp 1654583406
transform 1 0 18446 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_930
timestamp 1654583406
transform 1 0 26082 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_931
timestamp 1654583406
transform 1 0 16790 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_932
timestamp 1654583406
transform 1 0 16790 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_933
timestamp 1654583406
transform 1 0 16422 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_934
timestamp 1654583406
transform 1 0 15686 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_935
timestamp 1654583406
transform 1 0 15686 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_936
timestamp 1654583406
transform 1 0 13202 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_937
timestamp 1654583406
transform 1 0 13202 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_938
timestamp 1654583406
transform 1 0 12650 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_939
timestamp 1654583406
transform 1 0 12650 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_940
timestamp 1654583406
transform 1 0 12282 0 1 24514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_941
timestamp 1654583406
transform 1 0 230 0 1 24514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_942
timestamp 1654583406
transform 1 0 11638 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_943
timestamp 1654583406
transform 1 0 11638 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_944
timestamp 1654583406
transform 1 0 10718 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_945
timestamp 1654583406
transform 1 0 10718 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_946
timestamp 1654583406
transform 1 0 11362 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_947
timestamp 1654583406
transform 1 0 11362 0 1 15334
box -32 -32 32 32
use M1M2_PR  M1M2_PR_948
timestamp 1654583406
transform 1 0 5842 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_949
timestamp 1654583406
transform 1 0 10534 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_950
timestamp 1654583406
transform 1 0 10534 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_951
timestamp 1654583406
transform 1 0 4186 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_952
timestamp 1654583406
transform 1 0 7314 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_953
timestamp 1654583406
transform 1 0 15226 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_954
timestamp 1654583406
transform 1 0 13202 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_955
timestamp 1654583406
transform 1 0 13202 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_956
timestamp 1654583406
transform 1 0 11546 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_957
timestamp 1654583406
transform 1 0 8878 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_958
timestamp 1654583406
transform 1 0 8326 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_959
timestamp 1654583406
transform 1 0 7774 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_960
timestamp 1654583406
transform 1 0 7774 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_961
timestamp 1654583406
transform 1 0 6302 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_962
timestamp 1654583406
transform 1 0 6302 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_963
timestamp 1654583406
transform 1 0 6578 0 1 15266
box -32 -32 32 32
use M1M2_PR_MR  M1M2_PR_MR_0
timestamp 1654583406
transform 1 0 16330 0 1 18530
box -26 -32 26 32
use M1M2_PR_MR  M1M2_PR_MR_1
timestamp 1654583406
transform 1 0 16330 0 1 16354
box -26 -32 26 32
use M1M2_PR_M  M1M2_PR_M_0
timestamp 1654583406
transform 1 0 15686 0 1 14518
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_1
timestamp 1654583406
transform 1 0 19642 0 1 17578
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_2
timestamp 1654583406
transform 1 0 15502 0 1 13770
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_3
timestamp 1654583406
transform 1 0 13478 0 1 15674
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_4
timestamp 1654583406
transform 1 0 13202 0 1 16898
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_5
timestamp 1654583406
transform 1 0 7958 0 1 21046
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_6
timestamp 1654583406
transform 1 0 7958 0 1 16694
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_7
timestamp 1654583406
transform 1 0 7958 0 1 18870
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_8
timestamp 1654583406
transform 1 0 7958 0 1 18666
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_9
timestamp 1654583406
transform 1 0 15502 0 1 18326
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_10
timestamp 1654583406
transform 1 0 12834 0 1 19074
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_11
timestamp 1654583406
transform 1 0 7958 0 1 14314
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_12
timestamp 1654583406
transform 1 0 7958 0 1 9078
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_13
timestamp 1654583406
transform 1 0 8142 0 1 5814
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_14
timestamp 1654583406
transform 1 0 7958 0 1 7990
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_15
timestamp 1654583406
transform 1 0 15502 0 1 6154
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_16
timestamp 1654583406
transform 1 0 15502 0 1 11594
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_17
timestamp 1654583406
transform 1 0 15962 0 1 8262
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_18
timestamp 1654583406
transform 1 0 13386 0 1 7106
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_19
timestamp 1654583406
transform 1 0 8326 0 1 6698
box -32 -26 32 26
use M1M2_PR_R  M1M2_PR_R_0
timestamp 1654583406
transform 1 0 20194 0 1 14722
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_1
timestamp 1654583406
transform 1 0 18814 0 1 19074
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_2
timestamp 1654583406
transform 1 0 6946 0 1 12546
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_3
timestamp 1654583406
transform 1 0 22770 0 1 17986
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_4
timestamp 1654583406
transform 1 0 22770 0 1 15810
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_5
timestamp 1654583406
transform 1 0 6670 0 1 15198
box -32 -32 32 32
use M2M3_PR  M2M3_PR_0
timestamp 1654583406
transform 1 0 20654 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_1
timestamp 1654583406
transform 1 0 19182 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_2
timestamp 1654583406
transform 1 0 17802 0 1 13432
box -33 -37 33 37
use M2M3_PR  M2M3_PR_3
timestamp 1654583406
transform 1 0 16698 0 1 18556
box -33 -37 33 37
use M2M3_PR  M2M3_PR_4
timestamp 1654583406
transform 1 0 15686 0 1 13432
box -33 -37 33 37
use M2M3_PR  M2M3_PR_5
timestamp 1654583406
transform 1 0 15226 0 1 18556
box -33 -37 33 37
use M2M3_PR  M2M3_PR_6
timestamp 1654583406
transform 1 0 13294 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_7
timestamp 1654583406
transform 1 0 11730 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_8
timestamp 1654583406
transform 1 0 15870 0 1 18068
box -33 -37 33 37
use M2M3_PR  M2M3_PR_9
timestamp 1654583406
transform 1 0 14306 0 1 13554
box -33 -37 33 37
use M2M3_PR  M2M3_PR_10
timestamp 1654583406
transform 1 0 13662 0 1 18068
box -33 -37 33 37
use M2M3_PR  M2M3_PR_11
timestamp 1654583406
transform 1 0 13386 0 1 13554
box -33 -37 33 37
use M2M3_PR  M2M3_PR_12
timestamp 1654583406
transform 1 0 15870 0 1 12090
box -33 -37 33 37
use M2M3_PR  M2M3_PR_13
timestamp 1654583406
transform 1 0 14766 0 1 12090
box -33 -37 33 37
use M2M3_PR  M2M3_PR_14
timestamp 1654583406
transform 1 0 13202 0 1 12700
box -33 -37 33 37
use M2M3_PR  M2M3_PR_15
timestamp 1654583406
transform 1 0 12190 0 1 12700
box -33 -37 33 37
use M2M3_PR  M2M3_PR_16
timestamp 1654583406
transform 1 0 16054 0 1 16238
box -33 -37 33 37
use M2M3_PR  M2M3_PR_17
timestamp 1654583406
transform 1 0 14766 0 1 16238
box -33 -37 33 37
use M2M3_PR  M2M3_PR_18
timestamp 1654583406
transform 1 0 15778 0 1 14042
box -33 -37 33 37
use M2M3_PR  M2M3_PR_19
timestamp 1654583406
transform 1 0 15686 0 1 16970
box -33 -37 33 37
use M2M3_PR  M2M3_PR_20
timestamp 1654583406
transform 1 0 11178 0 1 14652
box -33 -37 33 37
use M2M3_PR  M2M3_PR_21
timestamp 1654583406
transform 1 0 10166 0 1 14652
box -33 -37 33 37
use M2M3_PR  M2M3_PR_22
timestamp 1654583406
transform 1 0 13662 0 1 12456
box -33 -37 33 37
use M2M3_PR  M2M3_PR_23
timestamp 1654583406
transform 1 0 12834 0 1 12456
box -33 -37 33 37
use M2M3_PR  M2M3_PR_24
timestamp 1654583406
transform 1 0 10810 0 1 12456
box -33 -37 33 37
use M2M3_PR  M2M3_PR_25
timestamp 1654583406
transform 1 0 9982 0 1 12456
box -33 -37 33 37
use M2M3_PR  M2M3_PR_26
timestamp 1654583406
transform 1 0 9522 0 1 12456
box -33 -37 33 37
use M2M3_PR  M2M3_PR_27
timestamp 1654583406
transform 1 0 20194 0 1 14164
box -33 -37 33 37
use M2M3_PR  M2M3_PR_28
timestamp 1654583406
transform 1 0 18906 0 1 14164
box -33 -37 33 37
use M2M3_PR  M2M3_PR_29
timestamp 1654583406
transform 1 0 17066 0 1 14164
box -33 -37 33 37
use M2M3_PR  M2M3_PR_30
timestamp 1654583406
transform 1 0 18814 0 1 18922
box -33 -37 33 37
use M2M3_PR  M2M3_PR_31
timestamp 1654583406
transform 1 0 17710 0 1 18922
box -33 -37 33 37
use M2M3_PR  M2M3_PR_32
timestamp 1654583406
transform 1 0 14766 0 1 18922
box -33 -37 33 37
use M2M3_PR  M2M3_PR_33
timestamp 1654583406
transform 1 0 12834 0 1 18922
box -33 -37 33 37
use M2M3_PR  M2M3_PR_34
timestamp 1654583406
transform 1 0 14490 0 1 6966
box -33 -37 33 37
use M2M3_PR  M2M3_PR_35
timestamp 1654583406
transform 1 0 13018 0 1 6966
box -33 -37 33 37
use M2M3_PR  M2M3_PR_36
timestamp 1654583406
transform 1 0 10166 0 1 13066
box -33 -37 33 37
use M2M3_PR  M2M3_PR_37
timestamp 1654583406
transform 1 0 6670 0 1 13066
box -33 -37 33 37
use M2M3_PR  M2M3_PR_38
timestamp 1654583406
transform 1 0 19182 0 1 9894
box -33 -37 33 37
use M2M3_PR  M2M3_PR_39
timestamp 1654583406
transform 1 0 16974 0 1 9894
box -33 -37 33 37
use M2M3_PR  M2M3_PR_40
timestamp 1654583406
transform 1 0 19918 0 1 18556
box -33 -37 33 37
use M2M3_PR  M2M3_PR_41
timestamp 1654583406
transform 1 0 19090 0 1 18556
box -33 -37 33 37
use M2M3_PR  M2M3_PR_42
timestamp 1654583406
transform 1 0 13846 0 1 10870
box -33 -37 33 37
use M2M3_PR  M2M3_PR_43
timestamp 1654583406
transform 1 0 13018 0 1 10870
box -33 -37 33 37
use M2M3_PR  M2M3_PR_44
timestamp 1654583406
transform 1 0 10258 0 1 10870
box -33 -37 33 37
use M2M3_PR  M2M3_PR_45
timestamp 1654583406
transform 1 0 22770 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_46
timestamp 1654583406
transform 1 0 20470 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_47
timestamp 1654583406
transform 1 0 12834 0 1 19654
box -33 -37 33 37
use M2M3_PR  M2M3_PR_48
timestamp 1654583406
transform 1 0 12834 0 1 9162
box -33 -37 33 37
use M2M3_PR  M2M3_PR_49
timestamp 1654583406
transform 1 0 12834 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_50
timestamp 1654583406
transform 1 0 12650 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_51
timestamp 1654583406
transform 1 0 12098 0 1 9162
box -33 -37 33 37
use M2M3_PR  M2M3_PR_52
timestamp 1654583406
transform 1 0 11638 0 1 19654
box -33 -37 33 37
use M2M3_PR  M2M3_PR_53
timestamp 1654583406
transform 1 0 11178 0 1 9162
box -33 -37 33 37
use M2M3_PR  M2M3_PR_54
timestamp 1654583406
transform 1 0 10902 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_55
timestamp 1654583406
transform 1 0 10810 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_56
timestamp 1654583406
transform 1 0 10258 0 1 19654
box -33 -37 33 37
use M2M3_PR  M2M3_PR_57
timestamp 1654583406
transform 1 0 9982 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_58
timestamp 1654583406
transform 1 0 9798 0 1 15262
box -33 -37 33 37
use M2M3_PR  M2M3_PR_59
timestamp 1654583406
transform 1 0 8878 0 1 15262
box -33 -37 33 37
use M2M3_PR  M2M3_PR_60
timestamp 1654583406
transform 1 0 8694 0 1 19654
box -33 -37 33 37
use M2M3_PR  M2M3_PR_61
timestamp 1654583406
transform 1 0 8694 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_62
timestamp 1654583406
transform 1 0 8694 0 1 6600
box -33 -37 33 37
use M2M3_PR  M2M3_PR_63
timestamp 1654583406
transform 1 0 8234 0 1 6600
box -33 -37 33 37
use M2M3_PR  M2M3_PR_64
timestamp 1654583406
transform 1 0 7958 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_65
timestamp 1654583406
transform 1 0 7774 0 1 19654
box -33 -37 33 37
use M2M3_PR  M2M3_PR_66
timestamp 1654583406
transform 1 0 7774 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_67
timestamp 1654583406
transform 1 0 7774 0 1 15262
box -33 -37 33 37
use M2M3_PR  M2M3_PR_68
timestamp 1654583406
transform 1 0 7498 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_69
timestamp 1654583406
transform 1 0 7222 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_70
timestamp 1654583406
transform 1 0 6946 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_71
timestamp 1654583406
transform 1 0 6210 0 1 8186
box -33 -37 33 37
use M2M3_PR  M2M3_PR_72
timestamp 1654583406
transform 1 0 6118 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_73
timestamp 1654583406
transform 1 0 6118 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_74
timestamp 1654583406
transform 1 0 22770 0 1 14652
box -33 -37 33 37
use M2M3_PR  M2M3_PR_75
timestamp 1654583406
transform 1 0 21482 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_76
timestamp 1654583406
transform 1 0 21482 0 1 14652
box -33 -37 33 37
use M2M3_PR  M2M3_PR_77
timestamp 1654583406
transform 1 0 21482 0 1 11480
box -33 -37 33 37
use M2M3_PR  M2M3_PR_78
timestamp 1654583406
transform 1 0 20378 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_79
timestamp 1654583406
transform 1 0 20102 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_80
timestamp 1654583406
transform 1 0 19090 0 1 11480
box -33 -37 33 37
use M2M3_PR  M2M3_PR_81
timestamp 1654583406
transform 1 0 19090 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_82
timestamp 1654583406
transform 1 0 18906 0 1 8308
box -33 -37 33 37
use M2M3_PR  M2M3_PR_83
timestamp 1654583406
transform 1 0 18538 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_84
timestamp 1654583406
transform 1 0 17710 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_85
timestamp 1654583406
transform 1 0 17710 0 1 8308
box -33 -37 33 37
use M2M3_PR  M2M3_PR_86
timestamp 1654583406
transform 1 0 17618 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_87
timestamp 1654583406
transform 1 0 15962 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_88
timestamp 1654583406
transform 1 0 15226 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_89
timestamp 1654583406
transform 1 0 14674 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_90
timestamp 1654583406
transform 1 0 13754 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_91
timestamp 1654583406
transform 1 0 13386 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_92
timestamp 1654583406
transform 1 0 16330 0 1 15750
box -33 -37 33 37
use M2M3_PR  M2M3_PR_93
timestamp 1654583406
transform 1 0 13018 0 1 15750
box -33 -37 33 37
use M2M3_PR  M2M3_PR_94
timestamp 1654583406
transform 1 0 8326 0 1 15750
box -33 -37 33 37
use M2M3_PR  M2M3_PR_95
timestamp 1654583406
transform 1 0 13110 0 1 14652
box -33 -37 33 37
use M2M3_PR  M2M3_PR_96
timestamp 1654583406
transform 1 0 11546 0 1 3672
box -33 -37 33 37
use M2M3_PR  M2M3_PR_97
timestamp 1654583406
transform 1 0 11454 0 1 8918
box -33 -37 33 37
use M2M3_PR  M2M3_PR_98
timestamp 1654583406
transform 1 0 10902 0 1 13066
box -33 -37 33 37
use M2M3_PR  M2M3_PR_99
timestamp 1654583406
transform 1 0 17434 0 1 7088
box -33 -37 33 37
use M2M3_PR  M2M3_PR_100
timestamp 1654583406
transform 1 0 22954 0 1 10504
box -33 -37 33 37
use M2M3_PR  M2M3_PR_101
timestamp 1654583406
transform 1 0 28566 0 1 13920
box -33 -37 33 37
use M2M3_PR  M2M3_PR_102
timestamp 1654583406
transform 1 0 19918 0 1 17458
box -33 -37 33 37
use M2M3_PR  M2M3_PR_103
timestamp 1654583406
transform 1 0 22126 0 1 20874
box -33 -37 33 37
use M2M3_PR  M2M3_PR_104
timestamp 1654583406
transform 1 0 26082 0 1 24290
box -33 -37 33 37
use M2M3_PR  M2M3_PR_105
timestamp 1654583406
transform 1 0 16422 0 1 27584
box -33 -37 33 37
use M2M3_PR  M2M3_PR_106
timestamp 1654583406
transform 1 0 13202 0 1 27584
box -33 -37 33 37
use M2M3_PR  M2M3_PR_107
timestamp 1654583406
transform 1 0 230 0 1 24534
box -33 -37 33 37
use M2M3_PR  M2M3_PR_108
timestamp 1654583406
transform 1 0 11546 0 1 21240
box -33 -37 33 37
use M2M3_PR  M2M3_PR_109
timestamp 1654583406
transform 1 0 10718 0 1 18434
box -33 -37 33 37
use M2M3_PR  M2M3_PR_110
timestamp 1654583406
transform 1 0 11362 0 1 9406
box -33 -37 33 37
use M2M3_PR  M2M3_PR_111
timestamp 1654583406
transform 1 0 5842 0 1 6234
box -33 -37 33 37
use M2M3_PR  M2M3_PR_112
timestamp 1654583406
transform 1 0 4186 0 1 3184
box -33 -37 33 37
use M2M3_PR  M2M3_PR_113
timestamp 1654583406
transform 1 0 7314 0 1 12334
box -33 -37 33 37
use M2M3_PR  M2M3_PR_114
timestamp 1654583406
transform 1 0 15226 0 1 6600
box -33 -37 33 37
use M2M3_PR  M2M3_PR_115
timestamp 1654583406
transform 1 0 13202 0 1 6600
box -33 -37 33 37
use M2M3_PR  M2M3_PR_116
timestamp 1654583406
transform 1 0 11546 0 1 5990
box -33 -37 33 37
use M2M3_PR  M2M3_PR_117
timestamp 1654583406
transform 1 0 8878 0 1 5990
box -33 -37 33 37
use M2M3_PR  M2M3_PR_118
timestamp 1654583406
transform 1 0 6302 0 1 134
box -33 -37 33 37
use M2M3_PR  M2M3_PR_119
timestamp 1654583406
transform 1 0 6578 0 1 15384
box -33 -37 33 37
use M3M4_PR  M3M4_PR_0
timestamp 1654583406
transform 1 0 15778 0 1 16970
box -38 -33 38 33
use M3M4_PR  M3M4_PR_1
timestamp 1654583406
transform 1 0 15778 0 1 14042
box -38 -33 38 33
use M3M4_PR  M3M4_PR_2
timestamp 1654583406
transform 1 0 12880 0 1 15262
box -38 -33 38 33
use M3M4_PR  M3M4_PR_3
timestamp 1654583406
transform 1 0 12880 0 1 11968
box -38 -33 38 33
use M3M4_PR  M3M4_PR_4
timestamp 1654583406
transform 1 0 12880 0 1 8186
box -38 -33 38 33
use M3M4_PR  M3M4_PR_5
timestamp 1654583406
transform 1 0 13294 0 1 14652
box -38 -33 38 33
use M3M4_PR  M3M4_PR_6
timestamp 1654583406
transform 1 0 13294 0 1 256
box -38 -33 38 33
use M3M4_PR  M3M4_PR_7
timestamp 1654583406
transform 1 0 11224 0 1 13066
box -38 -33 38 33
use M3M4_PR  M3M4_PR_8
timestamp 1654583406
transform 1 0 11224 0 1 8918
box -38 -33 38 33
use M3M4_PR  M3M4_PR_9
timestamp 1654583406
transform 1 0 6808 0 1 12334
box -38 -33 38 33
use M3M4_PR  M3M4_PR_10
timestamp 1654583406
transform 1 0 4738 0 1 12334
box -38 -33 38 33
use M4M5_PR  M4M5_PR_0
timestamp 1654583406
transform 1 0 6670 0 1 12334
box -142 -142 178 178
use M4M5_PR  M4M5_PR_1
timestamp 1654583406
transform 1 0 4876 0 1 12334
box -142 -142 178 178
use digital_filter_VIA0  digital_filter_VIA0_0
timestamp 1654583406
transform 1 0 20750 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_1
timestamp 1654583406
transform 1 0 15150 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_2
timestamp 1654583406
transform 1 0 9550 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_3
timestamp 1654583406
transform 1 0 20750 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_4
timestamp 1654583406
transform 1 0 15150 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_5
timestamp 1654583406
transform 1 0 9550 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_6
timestamp 1654583406
transform 1 0 23310 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_7
timestamp 1654583406
transform 1 0 23310 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_8
timestamp 1654583406
transform 1 0 5486 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_9
timestamp 1654583406
transform 1 0 5486 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_10
timestamp 1654583406
transform 1 0 19510 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_11
timestamp 1654583406
transform 1 0 13910 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_12
timestamp 1654583406
transform 1 0 8310 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_13
timestamp 1654583406
transform 1 0 19510 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_14
timestamp 1654583406
transform 1 0 13910 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_15
timestamp 1654583406
transform 1 0 8310 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_16
timestamp 1654583406
transform 1 0 24550 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_17
timestamp 1654583406
transform 1 0 24550 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_18
timestamp 1654583406
transform 1 0 4246 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_19
timestamp 1654583406
transform 1 0 4246 0 1 4162
box -310 -310 310 310
use digital_filter_VIA1  digital_filter_VIA1_0
timestamp 1654583406
transform 1 0 20750 0 1 21488
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_1
timestamp 1654583406
transform 1 0 20750 0 1 20400
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_2
timestamp 1654583406
transform 1 0 20750 0 1 19312
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_3
timestamp 1654583406
transform 1 0 20750 0 1 18224
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_4
timestamp 1654583406
transform 1 0 20750 0 1 17136
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_5
timestamp 1654583406
transform 1 0 20750 0 1 16048
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_6
timestamp 1654583406
transform 1 0 20750 0 1 14960
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_7
timestamp 1654583406
transform 1 0 20750 0 1 13872
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_8
timestamp 1654583406
transform 1 0 20750 0 1 12784
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_9
timestamp 1654583406
transform 1 0 20750 0 1 11696
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_10
timestamp 1654583406
transform 1 0 20750 0 1 10608
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_11
timestamp 1654583406
transform 1 0 20750 0 1 9520
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_12
timestamp 1654583406
transform 1 0 20750 0 1 8432
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_13
timestamp 1654583406
transform 1 0 20750 0 1 7344
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_14
timestamp 1654583406
transform 1 0 20750 0 1 6256
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_15
timestamp 1654583406
transform 1 0 15150 0 1 21488
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_16
timestamp 1654583406
transform 1 0 15150 0 1 20400
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_17
timestamp 1654583406
transform 1 0 15150 0 1 19312
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_18
timestamp 1654583406
transform 1 0 15150 0 1 18224
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_19
timestamp 1654583406
transform 1 0 15150 0 1 17136
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_20
timestamp 1654583406
transform 1 0 15150 0 1 16048
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_21
timestamp 1654583406
transform 1 0 15150 0 1 14960
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_22
timestamp 1654583406
transform 1 0 15150 0 1 13872
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_23
timestamp 1654583406
transform 1 0 15150 0 1 12784
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_24
timestamp 1654583406
transform 1 0 15150 0 1 11696
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_25
timestamp 1654583406
transform 1 0 15150 0 1 10608
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_26
timestamp 1654583406
transform 1 0 15150 0 1 9520
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_27
timestamp 1654583406
transform 1 0 15150 0 1 8432
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_28
timestamp 1654583406
transform 1 0 15150 0 1 7344
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_29
timestamp 1654583406
transform 1 0 15150 0 1 6256
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_30
timestamp 1654583406
transform 1 0 9550 0 1 21488
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_31
timestamp 1654583406
transform 1 0 9550 0 1 20400
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_32
timestamp 1654583406
transform 1 0 9550 0 1 19312
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_33
timestamp 1654583406
transform 1 0 9550 0 1 18224
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_34
timestamp 1654583406
transform 1 0 9550 0 1 17136
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_35
timestamp 1654583406
transform 1 0 9550 0 1 16048
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_36
timestamp 1654583406
transform 1 0 9550 0 1 14960
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_37
timestamp 1654583406
transform 1 0 9550 0 1 13872
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_38
timestamp 1654583406
transform 1 0 9550 0 1 12784
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_39
timestamp 1654583406
transform 1 0 9550 0 1 11696
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_40
timestamp 1654583406
transform 1 0 9550 0 1 10608
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_41
timestamp 1654583406
transform 1 0 9550 0 1 9520
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_42
timestamp 1654583406
transform 1 0 9550 0 1 8432
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_43
timestamp 1654583406
transform 1 0 9550 0 1 7344
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_44
timestamp 1654583406
transform 1 0 9550 0 1 6256
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_45
timestamp 1654583406
transform 1 0 19510 0 1 22032
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_46
timestamp 1654583406
transform 1 0 19510 0 1 20944
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_47
timestamp 1654583406
transform 1 0 19510 0 1 19856
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_48
timestamp 1654583406
transform 1 0 19510 0 1 18768
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_49
timestamp 1654583406
transform 1 0 19510 0 1 17680
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_50
timestamp 1654583406
transform 1 0 19510 0 1 16592
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_51
timestamp 1654583406
transform 1 0 19510 0 1 15504
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_52
timestamp 1654583406
transform 1 0 19510 0 1 14416
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_53
timestamp 1654583406
transform 1 0 19510 0 1 13328
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_54
timestamp 1654583406
transform 1 0 19510 0 1 12240
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_55
timestamp 1654583406
transform 1 0 19510 0 1 11152
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_56
timestamp 1654583406
transform 1 0 19510 0 1 10064
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_57
timestamp 1654583406
transform 1 0 19510 0 1 8976
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_58
timestamp 1654583406
transform 1 0 19510 0 1 7888
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_59
timestamp 1654583406
transform 1 0 19510 0 1 6800
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_60
timestamp 1654583406
transform 1 0 19510 0 1 5712
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_61
timestamp 1654583406
transform 1 0 13910 0 1 22032
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_62
timestamp 1654583406
transform 1 0 13910 0 1 20944
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_63
timestamp 1654583406
transform 1 0 13910 0 1 19856
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_64
timestamp 1654583406
transform 1 0 13910 0 1 18768
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_65
timestamp 1654583406
transform 1 0 13910 0 1 17680
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_66
timestamp 1654583406
transform 1 0 13910 0 1 16592
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_67
timestamp 1654583406
transform 1 0 13910 0 1 15504
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_68
timestamp 1654583406
transform 1 0 13910 0 1 14416
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_69
timestamp 1654583406
transform 1 0 13910 0 1 13328
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_70
timestamp 1654583406
transform 1 0 13910 0 1 12240
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_71
timestamp 1654583406
transform 1 0 13910 0 1 11152
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_72
timestamp 1654583406
transform 1 0 13910 0 1 10064
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_73
timestamp 1654583406
transform 1 0 13910 0 1 8976
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_74
timestamp 1654583406
transform 1 0 13910 0 1 7888
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_75
timestamp 1654583406
transform 1 0 13910 0 1 6800
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_76
timestamp 1654583406
transform 1 0 13910 0 1 5712
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_77
timestamp 1654583406
transform 1 0 8310 0 1 22032
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_78
timestamp 1654583406
transform 1 0 8310 0 1 20944
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_79
timestamp 1654583406
transform 1 0 8310 0 1 19856
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_80
timestamp 1654583406
transform 1 0 8310 0 1 18768
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_81
timestamp 1654583406
transform 1 0 8310 0 1 17680
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_82
timestamp 1654583406
transform 1 0 8310 0 1 16592
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_83
timestamp 1654583406
transform 1 0 8310 0 1 15504
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_84
timestamp 1654583406
transform 1 0 8310 0 1 14416
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_85
timestamp 1654583406
transform 1 0 8310 0 1 13328
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_86
timestamp 1654583406
transform 1 0 8310 0 1 12240
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_87
timestamp 1654583406
transform 1 0 8310 0 1 11152
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_88
timestamp 1654583406
transform 1 0 8310 0 1 10064
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_89
timestamp 1654583406
transform 1 0 8310 0 1 8976
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_90
timestamp 1654583406
transform 1 0 8310 0 1 7888
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_91
timestamp 1654583406
transform 1 0 8310 0 1 6800
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_92
timestamp 1654583406
transform 1 0 8310 0 1 5712
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_0
timestamp 1654583406
transform 1 0 20750 0 1 21488
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_1
timestamp 1654583406
transform 1 0 20750 0 1 20400
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_2
timestamp 1654583406
transform 1 0 20750 0 1 19312
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_3
timestamp 1654583406
transform 1 0 20750 0 1 18224
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_4
timestamp 1654583406
transform 1 0 20750 0 1 17136
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_5
timestamp 1654583406
transform 1 0 20750 0 1 16048
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_6
timestamp 1654583406
transform 1 0 20750 0 1 14960
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_7
timestamp 1654583406
transform 1 0 20750 0 1 13872
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_8
timestamp 1654583406
transform 1 0 20750 0 1 12784
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_9
timestamp 1654583406
transform 1 0 20750 0 1 11696
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_10
timestamp 1654583406
transform 1 0 20750 0 1 10608
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_11
timestamp 1654583406
transform 1 0 20750 0 1 9520
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_12
timestamp 1654583406
transform 1 0 20750 0 1 8432
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_13
timestamp 1654583406
transform 1 0 20750 0 1 7344
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_14
timestamp 1654583406
transform 1 0 20750 0 1 6256
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_15
timestamp 1654583406
transform 1 0 15150 0 1 21488
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_16
timestamp 1654583406
transform 1 0 15150 0 1 20400
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_17
timestamp 1654583406
transform 1 0 15150 0 1 19312
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_18
timestamp 1654583406
transform 1 0 15150 0 1 18224
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_19
timestamp 1654583406
transform 1 0 15150 0 1 17136
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_20
timestamp 1654583406
transform 1 0 15150 0 1 16048
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_21
timestamp 1654583406
transform 1 0 15150 0 1 14960
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_22
timestamp 1654583406
transform 1 0 15150 0 1 13872
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_23
timestamp 1654583406
transform 1 0 15150 0 1 12784
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_24
timestamp 1654583406
transform 1 0 15150 0 1 11696
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_25
timestamp 1654583406
transform 1 0 15150 0 1 10608
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_26
timestamp 1654583406
transform 1 0 15150 0 1 9520
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_27
timestamp 1654583406
transform 1 0 15150 0 1 8432
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_28
timestamp 1654583406
transform 1 0 15150 0 1 7344
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_29
timestamp 1654583406
transform 1 0 15150 0 1 6256
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_30
timestamp 1654583406
transform 1 0 9550 0 1 21488
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_31
timestamp 1654583406
transform 1 0 9550 0 1 20400
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_32
timestamp 1654583406
transform 1 0 9550 0 1 19312
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_33
timestamp 1654583406
transform 1 0 9550 0 1 18224
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_34
timestamp 1654583406
transform 1 0 9550 0 1 17136
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_35
timestamp 1654583406
transform 1 0 9550 0 1 16048
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_36
timestamp 1654583406
transform 1 0 9550 0 1 14960
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_37
timestamp 1654583406
transform 1 0 9550 0 1 13872
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_38
timestamp 1654583406
transform 1 0 9550 0 1 12784
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_39
timestamp 1654583406
transform 1 0 9550 0 1 11696
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_40
timestamp 1654583406
transform 1 0 9550 0 1 10608
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_41
timestamp 1654583406
transform 1 0 9550 0 1 9520
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_42
timestamp 1654583406
transform 1 0 9550 0 1 8432
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_43
timestamp 1654583406
transform 1 0 9550 0 1 7344
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_44
timestamp 1654583406
transform 1 0 9550 0 1 6256
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_45
timestamp 1654583406
transform 1 0 19510 0 1 22032
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_46
timestamp 1654583406
transform 1 0 19510 0 1 20944
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_47
timestamp 1654583406
transform 1 0 19510 0 1 19856
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_48
timestamp 1654583406
transform 1 0 19510 0 1 18768
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_49
timestamp 1654583406
transform 1 0 19510 0 1 17680
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_50
timestamp 1654583406
transform 1 0 19510 0 1 16592
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_51
timestamp 1654583406
transform 1 0 19510 0 1 15504
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_52
timestamp 1654583406
transform 1 0 19510 0 1 14416
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_53
timestamp 1654583406
transform 1 0 19510 0 1 13328
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_54
timestamp 1654583406
transform 1 0 19510 0 1 12240
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_55
timestamp 1654583406
transform 1 0 19510 0 1 11152
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_56
timestamp 1654583406
transform 1 0 19510 0 1 10064
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_57
timestamp 1654583406
transform 1 0 19510 0 1 8976
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_58
timestamp 1654583406
transform 1 0 19510 0 1 7888
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_59
timestamp 1654583406
transform 1 0 19510 0 1 6800
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_60
timestamp 1654583406
transform 1 0 19510 0 1 5712
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_61
timestamp 1654583406
transform 1 0 13910 0 1 22032
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_62
timestamp 1654583406
transform 1 0 13910 0 1 20944
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_63
timestamp 1654583406
transform 1 0 13910 0 1 19856
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_64
timestamp 1654583406
transform 1 0 13910 0 1 18768
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_65
timestamp 1654583406
transform 1 0 13910 0 1 17680
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_66
timestamp 1654583406
transform 1 0 13910 0 1 16592
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_67
timestamp 1654583406
transform 1 0 13910 0 1 15504
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_68
timestamp 1654583406
transform 1 0 13910 0 1 14416
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_69
timestamp 1654583406
transform 1 0 13910 0 1 13328
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_70
timestamp 1654583406
transform 1 0 13910 0 1 12240
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_71
timestamp 1654583406
transform 1 0 13910 0 1 11152
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_72
timestamp 1654583406
transform 1 0 13910 0 1 10064
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_73
timestamp 1654583406
transform 1 0 13910 0 1 8976
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_74
timestamp 1654583406
transform 1 0 13910 0 1 7888
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_75
timestamp 1654583406
transform 1 0 13910 0 1 6800
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_76
timestamp 1654583406
transform 1 0 13910 0 1 5712
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_77
timestamp 1654583406
transform 1 0 8310 0 1 22032
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_78
timestamp 1654583406
transform 1 0 8310 0 1 20944
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_79
timestamp 1654583406
transform 1 0 8310 0 1 19856
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_80
timestamp 1654583406
transform 1 0 8310 0 1 18768
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_81
timestamp 1654583406
transform 1 0 8310 0 1 17680
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_82
timestamp 1654583406
transform 1 0 8310 0 1 16592
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_83
timestamp 1654583406
transform 1 0 8310 0 1 15504
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_84
timestamp 1654583406
transform 1 0 8310 0 1 14416
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_85
timestamp 1654583406
transform 1 0 8310 0 1 13328
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_86
timestamp 1654583406
transform 1 0 8310 0 1 12240
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_87
timestamp 1654583406
transform 1 0 8310 0 1 11152
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_88
timestamp 1654583406
transform 1 0 8310 0 1 10064
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_89
timestamp 1654583406
transform 1 0 8310 0 1 8976
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_90
timestamp 1654583406
transform 1 0 8310 0 1 7888
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_91
timestamp 1654583406
transform 1 0 8310 0 1 6800
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_92
timestamp 1654583406
transform 1 0 8310 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_0
timestamp 1654583406
transform 1 0 20750 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_1
timestamp 1654583406
transform 1 0 20750 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_2
timestamp 1654583406
transform 1 0 20750 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_3
timestamp 1654583406
transform 1 0 20750 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_4
timestamp 1654583406
transform 1 0 20750 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_5
timestamp 1654583406
transform 1 0 20750 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_6
timestamp 1654583406
transform 1 0 20750 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_7
timestamp 1654583406
transform 1 0 20750 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_8
timestamp 1654583406
transform 1 0 20750 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_9
timestamp 1654583406
transform 1 0 20750 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_10
timestamp 1654583406
transform 1 0 20750 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_11
timestamp 1654583406
transform 1 0 20750 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_12
timestamp 1654583406
transform 1 0 20750 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_13
timestamp 1654583406
transform 1 0 20750 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_14
timestamp 1654583406
transform 1 0 20750 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_15
timestamp 1654583406
transform 1 0 15150 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_16
timestamp 1654583406
transform 1 0 15150 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_17
timestamp 1654583406
transform 1 0 15150 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_18
timestamp 1654583406
transform 1 0 15150 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_19
timestamp 1654583406
transform 1 0 15150 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_20
timestamp 1654583406
transform 1 0 15150 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_21
timestamp 1654583406
transform 1 0 15150 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_22
timestamp 1654583406
transform 1 0 15150 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_23
timestamp 1654583406
transform 1 0 15150 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_24
timestamp 1654583406
transform 1 0 15150 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_25
timestamp 1654583406
transform 1 0 15150 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_26
timestamp 1654583406
transform 1 0 15150 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_27
timestamp 1654583406
transform 1 0 15150 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_28
timestamp 1654583406
transform 1 0 15150 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_29
timestamp 1654583406
transform 1 0 15150 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_30
timestamp 1654583406
transform 1 0 9550 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_31
timestamp 1654583406
transform 1 0 9550 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_32
timestamp 1654583406
transform 1 0 9550 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_33
timestamp 1654583406
transform 1 0 9550 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_34
timestamp 1654583406
transform 1 0 9550 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_35
timestamp 1654583406
transform 1 0 9550 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_36
timestamp 1654583406
transform 1 0 9550 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_37
timestamp 1654583406
transform 1 0 9550 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_38
timestamp 1654583406
transform 1 0 9550 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_39
timestamp 1654583406
transform 1 0 9550 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_40
timestamp 1654583406
transform 1 0 9550 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_41
timestamp 1654583406
transform 1 0 9550 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_42
timestamp 1654583406
transform 1 0 9550 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_43
timestamp 1654583406
transform 1 0 9550 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_44
timestamp 1654583406
transform 1 0 9550 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_45
timestamp 1654583406
transform 1 0 19510 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_46
timestamp 1654583406
transform 1 0 19510 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_47
timestamp 1654583406
transform 1 0 19510 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_48
timestamp 1654583406
transform 1 0 19510 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_49
timestamp 1654583406
transform 1 0 19510 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_50
timestamp 1654583406
transform 1 0 19510 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_51
timestamp 1654583406
transform 1 0 19510 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_52
timestamp 1654583406
transform 1 0 19510 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_53
timestamp 1654583406
transform 1 0 19510 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_54
timestamp 1654583406
transform 1 0 19510 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_55
timestamp 1654583406
transform 1 0 19510 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_56
timestamp 1654583406
transform 1 0 19510 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_57
timestamp 1654583406
transform 1 0 19510 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_58
timestamp 1654583406
transform 1 0 19510 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_59
timestamp 1654583406
transform 1 0 19510 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_60
timestamp 1654583406
transform 1 0 19510 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_61
timestamp 1654583406
transform 1 0 13910 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_62
timestamp 1654583406
transform 1 0 13910 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_63
timestamp 1654583406
transform 1 0 13910 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_64
timestamp 1654583406
transform 1 0 13910 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_65
timestamp 1654583406
transform 1 0 13910 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_66
timestamp 1654583406
transform 1 0 13910 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_67
timestamp 1654583406
transform 1 0 13910 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_68
timestamp 1654583406
transform 1 0 13910 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_69
timestamp 1654583406
transform 1 0 13910 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_70
timestamp 1654583406
transform 1 0 13910 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_71
timestamp 1654583406
transform 1 0 13910 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_72
timestamp 1654583406
transform 1 0 13910 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_73
timestamp 1654583406
transform 1 0 13910 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_74
timestamp 1654583406
transform 1 0 13910 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_75
timestamp 1654583406
transform 1 0 13910 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_76
timestamp 1654583406
transform 1 0 13910 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_77
timestamp 1654583406
transform 1 0 8310 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_78
timestamp 1654583406
transform 1 0 8310 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_79
timestamp 1654583406
transform 1 0 8310 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_80
timestamp 1654583406
transform 1 0 8310 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_81
timestamp 1654583406
transform 1 0 8310 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_82
timestamp 1654583406
transform 1 0 8310 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_83
timestamp 1654583406
transform 1 0 8310 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_84
timestamp 1654583406
transform 1 0 8310 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_85
timestamp 1654583406
transform 1 0 8310 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_86
timestamp 1654583406
transform 1 0 8310 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_87
timestamp 1654583406
transform 1 0 8310 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_88
timestamp 1654583406
transform 1 0 8310 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_89
timestamp 1654583406
transform 1 0 8310 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_90
timestamp 1654583406
transform 1 0 8310 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_91
timestamp 1654583406
transform 1 0 8310 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_92
timestamp 1654583406
transform 1 0 8310 0 1 5712
box -310 -48 310 48
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_0
timestamp 1654583406
transform 1 0 22080 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_1
timestamp 1654583406
transform -1 0 22448 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_2
timestamp 1654583406
transform -1 0 19964 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_3
timestamp 1654583406
transform -1 0 12880 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_4
timestamp 1654583406
transform -1 0 10764 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_5
timestamp 1654583406
transform -1 0 8096 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_0
timestamp 1654583406
transform -1 0 12236 0 -1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_1
timestamp 1654583406
transform 1 0 10212 0 -1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_2
timestamp 1654583406
transform 1 0 11316 0 -1 18768
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_3
timestamp 1654583406
transform -1 0 13432 0 1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_4
timestamp 1654583406
transform 1 0 14168 0 -1 18768
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_5
timestamp 1654583406
transform -1 0 15640 0 -1 18768
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_6
timestamp 1654583406
transform 1 0 16284 0 1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_7
timestamp 1654583406
transform -1 0 18400 0 -1 18768
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_8
timestamp 1654583406
transform -1 0 19596 0 -1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_9
timestamp 1654583406
transform 1 0 20240 0 1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_10
timestamp 1654583406
transform -1 0 18308 0 1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_11
timestamp 1654583406
transform 1 0 15088 0 1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_12
timestamp 1654583406
transform -1 0 15916 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_13
timestamp 1654583406
transform 1 0 16468 0 -1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_14
timestamp 1654583406
transform -1 0 18492 0 1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_15
timestamp 1654583406
transform -1 0 18400 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_16
timestamp 1654583406
transform -1 0 16100 0 1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_17
timestamp 1654583406
transform -1 0 18308 0 1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_18
timestamp 1654583406
transform 1 0 15180 0 1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_19
timestamp 1654583406
transform 1 0 15088 0 1 11152
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_20
timestamp 1654583406
transform 1 0 14168 0 -1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_21
timestamp 1654583406
transform -1 0 13524 0 1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_22
timestamp 1654583406
transform 1 0 11408 0 1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_23
timestamp 1654583406
transform 1 0 11592 0 -1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_24
timestamp 1654583406
transform 1 0 10304 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_25
timestamp 1654583406
transform 1 0 12880 0 1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_26
timestamp 1654583406
transform 1 0 12880 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0
timestamp 1654583406
transform -1 0 6808 0 -1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_1
timestamp 1654583406
transform 1 0 9844 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_2
timestamp 1654583406
transform 1 0 6072 0 1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_3
timestamp 1654583406
transform -1 0 8372 0 1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_4
timestamp 1654583406
transform -1 0 8740 0 -1 18768
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_5
timestamp 1654583406
transform 1 0 7176 0 -1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_6
timestamp 1654583406
transform 1 0 7544 0 1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_7
timestamp 1654583406
transform 1 0 8464 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_8
timestamp 1654583406
transform -1 0 6716 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_9
timestamp 1654583406
transform 1 0 5888 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_10
timestamp 1654583406
transform 1 0 7636 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_11
timestamp 1654583406
transform 1 0 7912 0 1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_12
timestamp 1654583406
transform 1 0 8464 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_13
timestamp 1654583406
transform 1 0 10028 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_14
timestamp 1654583406
transform 1 0 12788 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_15
timestamp 1654583406
transform 1 0 13616 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_16
timestamp 1654583406
transform -1 0 14536 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_17
timestamp 1654583406
transform 1 0 16376 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_18
timestamp 1654583406
transform -1 0 18124 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_19
timestamp 1654583406
transform 1 0 16836 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_20
timestamp 1654583406
transform -1 0 18676 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_21
timestamp 1654583406
transform -1 0 19872 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_22
timestamp 1654583406
transform 1 0 20516 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_23
timestamp 1654583406
transform -1 0 19688 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_24
timestamp 1654583406
transform -1 0 21988 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_25
timestamp 1654583406
transform -1 0 22540 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_26
timestamp 1654583406
transform 1 0 21344 0 1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_27
timestamp 1654583406
transform 1 0 21344 0 1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_28
timestamp 1654583406
transform 1 0 20148 0 -1 22032
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_29
timestamp 1654583406
transform -1 0 19228 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_30
timestamp 1654583406
transform -1 0 16744 0 -1 22032
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_31
timestamp 1654583406
transform 1 0 15364 0 1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_32
timestamp 1654583406
transform 1 0 14260 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_33
timestamp 1654583406
transform -1 0 12788 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_34
timestamp 1654583406
transform 1 0 11592 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_35
timestamp 1654583406
transform 1 0 10028 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_36
timestamp 1654583406
transform 1 0 9752 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_37
timestamp 1654583406
transform 1 0 6532 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_38
timestamp 1654583406
transform 1 0 6164 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_39
timestamp 1654583406
transform -1 0 6808 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_40
timestamp 1654583406
transform 1 0 8556 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_41
timestamp 1654583406
transform -1 0 11868 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_42
timestamp 1654583406
transform 1 0 10488 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_43
timestamp 1654583406
transform -1 0 12788 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_44
timestamp 1654583406
transform 1 0 13984 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_45
timestamp 1654583406
transform 1 0 15640 0 1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_46
timestamp 1654583406
transform 1 0 17664 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_47
timestamp 1654583406
transform -1 0 17388 0 -1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_48
timestamp 1654583406
transform -1 0 19872 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_49
timestamp 1654583406
transform -1 0 19412 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_50
timestamp 1654583406
transform 1 0 20700 0 1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_51
timestamp 1654583406
transform -1 0 22540 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_52
timestamp 1654583406
transform -1 0 21988 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_53
timestamp 1654583406
transform 1 0 20608 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_54
timestamp 1654583406
transform -1 0 22264 0 1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_55
timestamp 1654583406
transform 1 0 22080 0 -1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_56
timestamp 1654583406
transform 1 0 6072 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_57
timestamp 1654583406
transform 1 0 6532 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_58
timestamp 1654583406
transform -1 0 7728 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_59
timestamp 1654583406
transform -1 0 8924 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_60
timestamp 1654583406
transform -1 0 11776 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_61
timestamp 1654583406
transform -1 0 12236 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_62
timestamp 1654583406
transform 1 0 12880 0 -1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_63
timestamp 1654583406
transform -1 0 13432 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_64
timestamp 1654583406
transform 1 0 15088 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0
timestamp 1654583406
transform 1 0 11316 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_1
timestamp 1654583406
transform 1 0 8924 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_2
timestamp 1654583406
transform -1 0 7452 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_3
timestamp 1654583406
transform -1 0 17940 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_4
timestamp 1654583406
transform 1 0 22632 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_5
timestamp 1654583406
transform 1 0 21620 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_6
timestamp 1654583406
transform 1 0 7176 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_7
timestamp 1654583406
transform -1 0 8096 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_8
timestamp 1654583406
transform -1 0 10580 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_9
timestamp 1654583406
transform -1 0 13432 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0
timestamp 1654583406
transform -1 0 6716 0 -1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_0
timestamp 1654583406
transform 1 0 7176 0 1 15504
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_1
timestamp 1654583406
transform -1 0 13524 0 -1 12240
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0
timestamp 1654583406
transform -1 0 13524 0 1 7888
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1654583406
transform 1 0 11316 0 1 10064
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinvlp_2  sky130_fd_sc_hd__clkinvlp_2_0
timestamp 1654583406
transform -1 0 20792 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0
timestamp 1654583406
transform 1 0 16192 0 1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_1
timestamp 1654583406
transform 1 0 11132 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0
timestamp 1654583406
transform 1 0 22632 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1654583406
transform 1 0 22632 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1654583406
transform 1 0 22632 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_3
timestamp 1654583406
transform 1 0 22632 0 -1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_4
timestamp 1654583406
transform 1 0 22632 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_5
timestamp 1654583406
transform 1 0 22632 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_6
timestamp 1654583406
transform 1 0 22632 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_7
timestamp 1654583406
transform 1 0 22632 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_8
timestamp 1654583406
transform 1 0 22632 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_9
timestamp 1654583406
transform 1 0 22632 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_10
timestamp 1654583406
transform 1 0 22632 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_11
timestamp 1654583406
transform 1 0 22264 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_12
timestamp 1654583406
transform 1 0 21344 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_13
timestamp 1654583406
transform 1 0 21344 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_14
timestamp 1654583406
transform 1 0 20976 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_15
timestamp 1654583406
transform 1 0 20976 0 1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_16
timestamp 1654583406
transform 1 0 20056 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_17
timestamp 1654583406
transform 1 0 19596 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_18
timestamp 1654583406
transform 1 0 19228 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_19
timestamp 1654583406
transform 1 0 18952 0 -1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_20
timestamp 1654583406
transform 1 0 18952 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_21
timestamp 1654583406
transform 1 0 18952 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_22
timestamp 1654583406
transform 1 0 18952 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_23
timestamp 1654583406
transform 1 0 18952 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_24
timestamp 1654583406
transform 1 0 18768 0 1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_25
timestamp 1654583406
transform 1 0 18400 0 1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_26
timestamp 1654583406
transform 1 0 18400 0 1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_27
timestamp 1654583406
transform 1 0 18400 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_28
timestamp 1654583406
transform 1 0 17480 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_29
timestamp 1654583406
transform 1 0 17480 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_30
timestamp 1654583406
transform 1 0 17480 0 -1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_31
timestamp 1654583406
transform 1 0 17480 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_32
timestamp 1654583406
transform 1 0 16744 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_33
timestamp 1654583406
transform 1 0 16376 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_34
timestamp 1654583406
transform 1 0 16376 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_35
timestamp 1654583406
transform 1 0 15824 0 1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_36
timestamp 1654583406
transform 1 0 15824 0 1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_37
timestamp 1654583406
transform 1 0 14904 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_38
timestamp 1654583406
transform 1 0 14904 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_39
timestamp 1654583406
transform 1 0 14536 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_40
timestamp 1654583406
transform 1 0 14536 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_41
timestamp 1654583406
transform 1 0 13800 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_42
timestamp 1654583406
transform 1 0 13800 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_43
timestamp 1654583406
transform 1 0 13616 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_44
timestamp 1654583406
transform 1 0 13248 0 1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_45
timestamp 1654583406
transform 1 0 12328 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_46
timestamp 1654583406
transform 1 0 11960 0 -1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_47
timestamp 1654583406
transform 1 0 11776 0 1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_48
timestamp 1654583406
transform 1 0 11776 0 1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_49
timestamp 1654583406
transform 1 0 11040 0 1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_50
timestamp 1654583406
transform 1 0 11040 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_51
timestamp 1654583406
transform 1 0 11224 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_52
timestamp 1654583406
transform 1 0 11040 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_53
timestamp 1654583406
transform 1 0 11040 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_54
timestamp 1654583406
transform 1 0 10672 0 1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_55
timestamp 1654583406
transform 1 0 10672 0 1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_56
timestamp 1654583406
transform 1 0 10672 0 1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_57
timestamp 1654583406
transform 1 0 10672 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_58
timestamp 1654583406
transform 1 0 10672 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_59
timestamp 1654583406
transform 1 0 9752 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_60
timestamp 1654583406
transform 1 0 9384 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_61
timestamp 1654583406
transform 1 0 9200 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_62
timestamp 1654583406
transform 1 0 9384 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_63
timestamp 1654583406
transform 1 0 8648 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_64
timestamp 1654583406
transform 1 0 8648 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_65
timestamp 1654583406
transform 1 0 8648 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_66
timestamp 1654583406
transform 1 0 8096 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_67
timestamp 1654583406
transform 1 0 8096 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_68
timestamp 1654583406
transform 1 0 7544 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_69
timestamp 1654583406
transform 1 0 6808 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_70
timestamp 1654583406
transform 1 0 6992 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_71
timestamp 1654583406
transform 1 0 5796 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_72
timestamp 1654583406
transform 1 0 5888 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_73
timestamp 1654583406
transform 1 0 5888 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_74
timestamp 1654583406
transform 1 0 5888 0 1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1654583406
transform 1 0 22172 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1654583406
transform 1 0 22080 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1654583406
transform 1 0 21712 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1654583406
transform 1 0 21344 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1654583406
transform 1 0 20884 0 1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1654583406
transform 1 0 20884 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1654583406
transform 1 0 20608 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1654583406
transform 1 0 20332 0 1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1654583406
transform 1 0 20148 0 -1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1654583406
transform 1 0 20148 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_10
timestamp 1654583406
transform 1 0 19504 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_11
timestamp 1654583406
transform 1 0 19228 0 1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_12
timestamp 1654583406
transform 1 0 19044 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_13
timestamp 1654583406
transform 1 0 18860 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_14
timestamp 1654583406
transform 1 0 18308 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_15
timestamp 1654583406
transform 1 0 18124 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_16
timestamp 1654583406
transform 1 0 17756 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_17
timestamp 1654583406
transform 1 0 17020 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_18
timestamp 1654583406
transform 1 0 17020 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_19
timestamp 1654583406
transform 1 0 17020 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_20
timestamp 1654583406
transform 1 0 16560 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_21
timestamp 1654583406
transform 1 0 15732 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_22
timestamp 1654583406
transform 1 0 15640 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_23
timestamp 1654583406
transform 1 0 15272 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_24
timestamp 1654583406
transform 1 0 15088 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_25
timestamp 1654583406
transform 1 0 15272 0 1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_26
timestamp 1654583406
transform 1 0 14904 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_27
timestamp 1654583406
transform 1 0 14904 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_28
timestamp 1654583406
transform 1 0 14444 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_29
timestamp 1654583406
transform 1 0 14444 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_30
timestamp 1654583406
transform 1 0 14444 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_31
timestamp 1654583406
transform 1 0 14444 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_32
timestamp 1654583406
transform 1 0 14168 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_33
timestamp 1654583406
transform 1 0 13800 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_34
timestamp 1654583406
transform 1 0 13064 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_35
timestamp 1654583406
transform 1 0 12696 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_36
timestamp 1654583406
transform 1 0 12328 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_37
timestamp 1654583406
transform 1 0 12328 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_38
timestamp 1654583406
transform 1 0 12052 0 1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_39
timestamp 1654583406
transform 1 0 11868 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_40
timestamp 1654583406
transform 1 0 11040 0 1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_41
timestamp 1654583406
transform 1 0 10580 0 1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_42
timestamp 1654583406
transform 1 0 10396 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_43
timestamp 1654583406
transform 1 0 9660 0 1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_44
timestamp 1654583406
transform 1 0 9844 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_45
timestamp 1654583406
transform 1 0 9844 0 -1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_46
timestamp 1654583406
transform 1 0 9844 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_47
timestamp 1654583406
transform 1 0 9292 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_48
timestamp 1654583406
transform 1 0 9016 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_49
timestamp 1654583406
transform 1 0 8464 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_50
timestamp 1654583406
transform 1 0 8464 0 1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_51
timestamp 1654583406
transform 1 0 8464 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_52
timestamp 1654583406
transform 1 0 8464 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_53
timestamp 1654583406
transform 1 0 8004 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_54
timestamp 1654583406
transform 1 0 8004 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_55
timestamp 1654583406
transform 1 0 8004 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_56
timestamp 1654583406
transform 1 0 7544 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_57
timestamp 1654583406
transform 1 0 6716 0 -1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_58
timestamp 1654583406
transform 1 0 6624 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_59
timestamp 1654583406
transform 1 0 6624 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_60
timestamp 1654583406
transform 1 0 6256 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_61
timestamp 1654583406
transform 1 0 6164 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_62
timestamp 1654583406
transform 1 0 5888 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_63
timestamp 1654583406
transform 1 0 5888 0 -1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_64
timestamp 1654583406
transform 1 0 5888 0 1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1654583406
transform 1 0 21988 0 -1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1654583406
transform 1 0 21528 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1654583406
transform 1 0 21528 0 -1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1654583406
transform 1 0 20700 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1654583406
transform 1 0 20608 0 1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1654583406
transform 1 0 17940 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1654583406
transform 1 0 17940 0 1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1654583406
transform 1 0 16284 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1654583406
transform 1 0 14260 0 -1 16592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1654583406
transform 1 0 14076 0 1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1654583406
transform 1 0 12972 0 1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_11
timestamp 1654583406
transform 1 0 12328 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_12
timestamp 1654583406
transform 1 0 11684 0 -1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_13
timestamp 1654583406
transform 1 0 11684 0 -1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_14
timestamp 1654583406
transform 1 0 11684 0 -1 12240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_15
timestamp 1654583406
transform 1 0 11040 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_16
timestamp 1654583406
transform 1 0 9752 0 -1 7888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_17
timestamp 1654583406
transform 1 0 9752 0 -1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_18
timestamp 1654583406
transform 1 0 9108 0 -1 18768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_19
timestamp 1654583406
transform 1 0 9108 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_20
timestamp 1654583406
transform 1 0 9108 0 -1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_21
timestamp 1654583406
transform 1 0 7820 0 1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_22
timestamp 1654583406
transform 1 0 7820 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_23
timestamp 1654583406
transform 1 0 7268 0 -1 16592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_24
timestamp 1654583406
transform 1 0 7268 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_25
timestamp 1654583406
transform 1 0 6532 0 1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_26
timestamp 1654583406
transform 1 0 6532 0 -1 7888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_27
timestamp 1654583406
transform 1 0 6532 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_28
timestamp 1654583406
transform 1 0 5796 0 -1 14416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_29
timestamp 1654583406
transform 1 0 5796 0 -1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0
timestamp 1654583406
transform 1 0 21988 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1654583406
transform 1 0 21804 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_2
timestamp 1654583406
transform 1 0 21436 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_3
timestamp 1654583406
transform 1 0 20424 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_4
timestamp 1654583406
transform 1 0 20148 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_5
timestamp 1654583406
transform 1 0 20424 0 1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_6
timestamp 1654583406
transform 1 0 20424 0 1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_7
timestamp 1654583406
transform 1 0 20424 0 1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_8
timestamp 1654583406
transform 1 0 20424 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_9
timestamp 1654583406
transform 1 0 20424 0 1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_10
timestamp 1654583406
transform 1 0 20148 0 -1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_11
timestamp 1654583406
transform 1 0 19872 0 1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_12
timestamp 1654583406
transform 1 0 19228 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_13
timestamp 1654583406
transform 1 0 19228 0 -1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_14
timestamp 1654583406
transform 1 0 19228 0 -1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_15
timestamp 1654583406
transform 1 0 19228 0 -1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_16
timestamp 1654583406
transform 1 0 19228 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_17
timestamp 1654583406
transform 1 0 19228 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_18
timestamp 1654583406
transform 1 0 18860 0 1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_19
timestamp 1654583406
transform 1 0 17756 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_20
timestamp 1654583406
transform 1 0 17756 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_21
timestamp 1654583406
transform 1 0 17756 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_22
timestamp 1654583406
transform 1 0 17756 0 1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_23
timestamp 1654583406
transform 1 0 17756 0 1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_24
timestamp 1654583406
transform 1 0 16652 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_25
timestamp 1654583406
transform 1 0 16652 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_26
timestamp 1654583406
transform 1 0 16652 0 -1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_27
timestamp 1654583406
transform 1 0 16652 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_28
timestamp 1654583406
transform 1 0 16652 0 -1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_29
timestamp 1654583406
transform 1 0 16192 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_30
timestamp 1654583406
transform 1 0 16192 0 1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_31
timestamp 1654583406
transform 1 0 16192 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_32
timestamp 1654583406
transform 1 0 15180 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_33
timestamp 1654583406
transform 1 0 15180 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_34
timestamp 1654583406
transform 1 0 15180 0 1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_35
timestamp 1654583406
transform 1 0 15180 0 1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_36
timestamp 1654583406
transform 1 0 14996 0 -1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_37
timestamp 1654583406
transform 1 0 15180 0 -1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_38
timestamp 1654583406
transform 1 0 14076 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_39
timestamp 1654583406
transform 1 0 13616 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_40
timestamp 1654583406
transform 1 0 13616 0 1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_41
timestamp 1654583406
transform 1 0 12420 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_42
timestamp 1654583406
transform 1 0 12604 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_43
timestamp 1654583406
transform 1 0 12604 0 -1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_44
timestamp 1654583406
transform 1 0 11500 0 -1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_45
timestamp 1654583406
transform 1 0 11040 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_46
timestamp 1654583406
transform 1 0 11040 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_47
timestamp 1654583406
transform 1 0 11040 0 1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_48
timestamp 1654583406
transform 1 0 10212 0 1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_49
timestamp 1654583406
transform 1 0 10212 0 1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_50
timestamp 1654583406
transform 1 0 9936 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_51
timestamp 1654583406
transform 1 0 9936 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_52
timestamp 1654583406
transform 1 0 9936 0 1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_53
timestamp 1654583406
transform 1 0 9936 0 1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_54
timestamp 1654583406
transform 1 0 8924 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_55
timestamp 1654583406
transform 1 0 8924 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_56
timestamp 1654583406
transform 1 0 8648 0 1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_57
timestamp 1654583406
transform 1 0 8924 0 -1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_58
timestamp 1654583406
transform 1 0 8924 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_59
timestamp 1654583406
transform 1 0 8924 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_60
timestamp 1654583406
transform 1 0 8924 0 -1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_61
timestamp 1654583406
transform 1 0 7636 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_62
timestamp 1654583406
transform 1 0 7636 0 1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_63
timestamp 1654583406
transform 1 0 7636 0 1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_64
timestamp 1654583406
transform 1 0 7176 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_65
timestamp 1654583406
transform 1 0 6348 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_66
timestamp 1654583406
transform 1 0 6164 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0
timestamp 1654583406
transform 1 0 21620 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1654583406
transform 1 0 21620 0 1 6800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_2
timestamp 1654583406
transform 1 0 21160 0 -1 6800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_3
timestamp 1654583406
transform 1 0 20056 0 1 19856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_4
timestamp 1654583406
transform 1 0 20056 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_5
timestamp 1654583406
transform 1 0 19596 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_6
timestamp 1654583406
transform 1 0 16468 0 1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_7
timestamp 1654583406
transform 1 0 14904 0 -1 11152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_8
timestamp 1654583406
transform 1 0 13340 0 -1 14416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_9
timestamp 1654583406
transform 1 0 8648 0 1 13328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_10
timestamp 1654583406
transform 1 0 7084 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_11
timestamp 1654583406
transform 1 0 5980 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_12
timestamp 1654583406
transform 1 0 5980 0 -1 16592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_13
timestamp 1654583406
transform 1 0 5980 0 -1 8976
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0
timestamp 1654583406
transform -1 0 9108 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_1
timestamp 1654583406
transform 1 0 6072 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_2
timestamp 1654583406
transform 1 0 8188 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_3
timestamp 1654583406
transform 1 0 11408 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_4
timestamp 1654583406
transform 1 0 10764 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_5
timestamp 1654583406
transform -1 0 12880 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_6
timestamp 1654583406
transform -1 0 12788 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_7
timestamp 1654583406
transform -1 0 15088 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_8
timestamp 1654583406
transform -1 0 15088 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_9
timestamp 1654583406
transform -1 0 17664 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_10
timestamp 1654583406
transform 1 0 14904 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_11
timestamp 1654583406
transform 1 0 16928 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_12
timestamp 1654583406
transform 1 0 17480 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_13
timestamp 1654583406
transform 1 0 18768 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_14
timestamp 1654583406
transform 1 0 17480 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_15
timestamp 1654583406
transform -1 0 15088 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_16
timestamp 1654583406
transform -1 0 17664 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_17
timestamp 1654583406
transform -1 0 17664 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_18
timestamp 1654583406
transform 1 0 17480 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_19
timestamp 1654583406
transform 1 0 14904 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_20
timestamp 1654583406
transform -1 0 17664 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_21
timestamp 1654583406
transform 1 0 17480 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_22
timestamp 1654583406
transform -1 0 16376 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_23
timestamp 1654583406
transform -1 0 16376 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_24
timestamp 1654583406
transform 1 0 12052 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_25
timestamp 1654583406
transform 1 0 13616 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_26
timestamp 1654583406
transform -1 0 12512 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_27
timestamp 1654583406
transform 1 0 11040 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_28
timestamp 1654583406
transform -1 0 14260 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_29
timestamp 1654583406
transform -1 0 15088 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_30
timestamp 1654583406
transform 1 0 7176 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_31
timestamp 1654583406
transform 1 0 6900 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_32
timestamp 1654583406
transform 1 0 9752 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_33
timestamp 1654583406
transform 1 0 9384 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_34
timestamp 1654583406
transform 1 0 9476 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_35
timestamp 1654583406
transform 1 0 9752 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_36
timestamp 1654583406
transform 1 0 10764 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_37
timestamp 1654583406
transform -1 0 13800 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_38
timestamp 1654583406
transform 1 0 13616 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_39
timestamp 1654583406
transform -1 0 17664 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_40
timestamp 1654583406
transform -1 0 17388 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_41
timestamp 1654583406
transform -1 0 17664 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_42
timestamp 1654583406
transform -1 0 18952 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_43
timestamp 1654583406
transform -1 0 19228 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_44
timestamp 1654583406
transform -1 0 20240 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_45
timestamp 1654583406
transform -1 0 21528 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_46
timestamp 1654583406
transform -1 0 20240 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_47
timestamp 1654583406
transform -1 0 18952 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_48
timestamp 1654583406
transform -1 0 20240 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_49
timestamp 1654583406
transform 1 0 18860 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_50
timestamp 1654583406
transform 1 0 18492 0 -1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_51
timestamp 1654583406
transform 1 0 18768 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_52
timestamp 1654583406
transform 1 0 17664 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_53
timestamp 1654583406
transform 1 0 14996 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_54
timestamp 1654583406
transform -1 0 14628 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_55
timestamp 1654583406
transform -1 0 13800 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_56
timestamp 1654583406
transform -1 0 15088 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_57
timestamp 1654583406
transform -1 0 12512 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_58
timestamp 1654583406
transform 1 0 9476 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_59
timestamp 1654583406
transform 1 0 9752 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_60
timestamp 1654583406
transform 1 0 6072 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_61
timestamp 1654583406
transform 1 0 5980 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_62
timestamp 1654583406
transform 1 0 7636 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_63
timestamp 1654583406
transform 1 0 8464 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_64
timestamp 1654583406
transform -1 0 8648 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_65
timestamp 1654583406
transform -1 0 7544 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_66
timestamp 1654583406
transform -1 0 9936 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_67
timestamp 1654583406
transform 1 0 6256 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_68
timestamp 1654583406
transform 1 0 6072 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_69
timestamp 1654583406
transform 1 0 8832 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_70
timestamp 1654583406
transform 1 0 7820 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_71
timestamp 1654583406
transform 1 0 7912 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_72
timestamp 1654583406
transform -1 0 10856 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_73
timestamp 1654583406
transform -1 0 12788 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_74
timestamp 1654583406
transform -1 0 13800 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_75
timestamp 1654583406
transform 1 0 13616 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_76
timestamp 1654583406
transform 1 0 14628 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_77
timestamp 1654583406
transform -1 0 17664 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_78
timestamp 1654583406
transform 1 0 17480 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_79
timestamp 1654583406
transform 1 0 18768 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_80
timestamp 1654583406
transform 1 0 20056 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_81
timestamp 1654583406
transform 1 0 21344 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_82
timestamp 1654583406
transform 1 0 19044 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_83
timestamp 1654583406
transform -1 0 21528 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_84
timestamp 1654583406
transform -1 0 22816 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_85
timestamp 1654583406
transform -1 0 22816 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_86
timestamp 1654583406
transform -1 0 22816 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_87
timestamp 1654583406
transform 1 0 20516 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_88
timestamp 1654583406
transform 1 0 18492 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_89
timestamp 1654583406
transform 1 0 15916 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_90
timestamp 1654583406
transform -1 0 17664 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_91
timestamp 1654583406
transform -1 0 15272 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_92
timestamp 1654583406
transform 1 0 12052 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_93
timestamp 1654583406
transform 1 0 12788 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_94
timestamp 1654583406
transform 1 0 10212 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_95
timestamp 1654583406
transform -1 0 11684 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_96
timestamp 1654583406
transform -1 0 22816 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_97
timestamp 1654583406
transform -1 0 21804 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_98
timestamp 1654583406
transform -1 0 21528 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_99
timestamp 1654583406
transform -1 0 21528 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_100
timestamp 1654583406
transform 1 0 21344 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_101
timestamp 1654583406
transform 1 0 20884 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_102
timestamp 1654583406
transform 1 0 18860 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_103
timestamp 1654583406
transform 1 0 17664 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_104
timestamp 1654583406
transform 1 0 16928 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_105
timestamp 1654583406
transform 1 0 17480 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_106
timestamp 1654583406
transform -1 0 16560 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_107
timestamp 1654583406
transform 1 0 14352 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_108
timestamp 1654583406
transform 1 0 12052 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_109
timestamp 1654583406
transform -1 0 11224 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_110
timestamp 1654583406
transform -1 0 10488 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_111
timestamp 1654583406
transform 1 0 7176 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_112
timestamp 1654583406
transform 1 0 6164 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_113
timestamp 1654583406
transform 1 0 6440 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_114
timestamp 1654583406
transform 1 0 13616 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_115
timestamp 1654583406
transform 1 0 16192 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_116
timestamp 1654583406
transform 1 0 13340 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_117
timestamp 1654583406
transform 1 0 11040 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_118
timestamp 1654583406
transform 1 0 10764 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_119
timestamp 1654583406
transform 1 0 8464 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_120
timestamp 1654583406
transform 1 0 7176 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_121
timestamp 1654583406
transform 1 0 6164 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_122
timestamp 1654583406
transform -1 0 7544 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_0
timestamp 1654583406
transform 1 0 20884 0 -1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_1
timestamp 1654583406
transform -1 0 21804 0 -1 16592
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_2
timestamp 1654583406
transform 1 0 21344 0 1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_3
timestamp 1654583406
transform 1 0 21344 0 1 12240
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_4
timestamp 1654583406
transform -1 0 22080 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_5
timestamp 1654583406
transform 1 0 21344 0 1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_6
timestamp 1654583406
transform 1 0 21344 0 1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_7
timestamp 1654583406
transform -1 0 21712 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_8
timestamp 1654583406
transform -1 0 20424 0 1 6800
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_9
timestamp 1654583406
transform 1 0 18768 0 1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_10
timestamp 1654583406
transform -1 0 17848 0 1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_11
timestamp 1654583406
transform -1 0 16560 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_12
timestamp 1654583406
transform -1 0 13984 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_13
timestamp 1654583406
transform 1 0 10580 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_14
timestamp 1654583406
transform -1 0 10120 0 1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_15
timestamp 1654583406
transform -1 0 8924 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_16
timestamp 1654583406
transform -1 0 8832 0 -1 14416
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_17
timestamp 1654583406
transform -1 0 19136 0 -1 6800
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_18
timestamp 1654583406
transform -1 0 16560 0 -1 6800
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_19
timestamp 1654583406
transform -1 0 15272 0 1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_20
timestamp 1654583406
transform -1 0 14444 0 -1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_21
timestamp 1654583406
transform -1 0 12236 0 -1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_22
timestamp 1654583406
transform 1 0 9752 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_23
timestamp 1654583406
transform -1 0 10120 0 1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_24
timestamp 1654583406
transform -1 0 9108 0 -1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0
timestamp 1654583406
transform 1 0 22908 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1654583406
transform 1 0 18768 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1654583406
transform 1 0 18492 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1654583406
transform 1 0 22724 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1654583406
transform 1 0 16192 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1654583406
transform 1 0 10488 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1654583406
transform 1 0 9568 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1654583406
transform 1 0 8188 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1654583406
transform 1 0 5888 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1654583406
transform 1 0 22908 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1654583406
transform 1 0 20056 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1654583406
transform 1 0 5796 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1654583406
transform 1 0 18492 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1654583406
transform 1 0 17664 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1654583406
transform 1 0 7728 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1654583406
transform 1 0 22908 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1654583406
transform 1 0 20056 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1654583406
transform 1 0 19136 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1654583406
transform 1 0 12328 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1654583406
transform 1 0 9752 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1654583406
transform 1 0 15916 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21
timestamp 1654583406
transform 1 0 15088 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_22
timestamp 1654583406
transform 1 0 13340 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_23
timestamp 1654583406
transform 1 0 12512 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_24
timestamp 1654583406
transform 1 0 7544 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_25
timestamp 1654583406
transform 1 0 22908 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_26
timestamp 1654583406
transform 1 0 20056 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_27
timestamp 1654583406
transform 1 0 10396 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_28
timestamp 1654583406
transform 1 0 9752 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_29
timestamp 1654583406
transform 1 0 21160 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_30
timestamp 1654583406
transform 1 0 20332 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_31
timestamp 1654583406
transform 1 0 15916 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_32
timestamp 1654583406
transform 1 0 15088 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_33
timestamp 1654583406
transform 1 0 22908 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_34
timestamp 1654583406
transform 1 0 11776 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_35
timestamp 1654583406
transform 1 0 9752 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_36
timestamp 1654583406
transform 1 0 18492 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_37
timestamp 1654583406
transform 1 0 17664 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_38
timestamp 1654583406
transform 1 0 15916 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_39
timestamp 1654583406
transform 1 0 15088 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_40
timestamp 1654583406
transform 1 0 14904 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_41
timestamp 1654583406
transform 1 0 10304 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_42
timestamp 1654583406
transform 1 0 7176 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_43
timestamp 1654583406
transform 1 0 12880 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_44
timestamp 1654583406
transform 1 0 22908 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_45
timestamp 1654583406
transform 1 0 8832 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_46
timestamp 1654583406
transform 1 0 18768 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_47
timestamp 1654583406
transform 1 0 14352 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_48
timestamp 1654583406
transform 1 0 13524 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_49
timestamp 1654583406
transform 1 0 11592 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_50
timestamp 1654583406
transform 1 0 21160 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_51
timestamp 1654583406
transform 1 0 20516 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_52
timestamp 1654583406
transform 1 0 18492 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_53
timestamp 1654583406
transform 1 0 17664 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_54
timestamp 1654583406
transform 1 0 8924 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_55
timestamp 1654583406
transform 1 0 7912 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_56
timestamp 1654583406
transform 1 0 16928 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_57
timestamp 1654583406
transform 1 0 10120 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_58
timestamp 1654583406
transform 1 0 22908 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_59
timestamp 1654583406
transform 1 0 18952 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_60
timestamp 1654583406
transform 1 0 18492 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_61
timestamp 1654583406
transform 1 0 17848 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_62
timestamp 1654583406
transform 1 0 22908 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_63
timestamp 1654583406
transform 1 0 16560 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_64
timestamp 1654583406
transform 1 0 10120 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_65
timestamp 1654583406
transform 1 0 22908 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_66
timestamp 1654583406
transform 1 0 20056 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_67
timestamp 1654583406
transform 1 0 16560 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_68
timestamp 1654583406
transform 1 0 22724 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_69
timestamp 1654583406
transform 1 0 20792 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_70
timestamp 1654583406
transform 1 0 7728 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_71
timestamp 1654583406
transform 1 0 22908 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_72
timestamp 1654583406
transform 1 0 22908 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_73
timestamp 1654583406
transform 1 0 21344 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_74
timestamp 1654583406
transform 1 0 16928 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_75
timestamp 1654583406
transform 1 0 7176 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_76
timestamp 1654583406
transform 1 0 22448 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_77
timestamp 1654583406
transform 1 0 20056 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_78
timestamp 1654583406
transform 1 0 19872 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_79
timestamp 1654583406
transform 1 0 18584 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_80
timestamp 1654583406
transform 1 0 16192 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_81
timestamp 1654583406
transform 1 0 16008 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_82
timestamp 1654583406
transform 1 0 13432 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_83
timestamp 1654583406
transform 1 0 11040 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_84
timestamp 1654583406
transform 1 0 10856 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_85
timestamp 1654583406
transform 1 0 6992 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_86
timestamp 1654583406
transform 1 0 8280 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_87
timestamp 1654583406
transform 1 0 14720 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_88
timestamp 1654583406
transform 1 0 8372 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_89
timestamp 1654583406
transform 1 0 7176 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_90
timestamp 1654583406
transform 1 0 22908 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_91
timestamp 1654583406
transform 1 0 21160 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_92
timestamp 1654583406
transform 1 0 18584 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_93
timestamp 1654583406
transform 1 0 15272 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_94
timestamp 1654583406
transform 1 0 14904 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_95
timestamp 1654583406
transform 1 0 5796 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_96
timestamp 1654583406
transform 1 0 21160 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_97
timestamp 1654583406
transform 1 0 16008 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_98
timestamp 1654583406
transform 1 0 13432 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_99
timestamp 1654583406
transform 1 0 18400 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_100
timestamp 1654583406
transform 1 0 15640 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_101
timestamp 1654583406
transform 1 0 14904 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_102
timestamp 1654583406
transform 1 0 11224 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_103
timestamp 1654583406
transform 1 0 6992 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_104
timestamp 1654583406
transform 1 0 5796 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_105
timestamp 1654583406
transform 1 0 18768 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_106
timestamp 1654583406
transform 1 0 16192 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_107
timestamp 1654583406
transform 1 0 16008 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_108
timestamp 1654583406
transform 1 0 13432 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_109
timestamp 1654583406
transform 1 0 21804 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_110
timestamp 1654583406
transform 1 0 22264 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_111
timestamp 1654583406
transform 1 0 18584 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_112
timestamp 1654583406
transform 1 0 16008 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_113
timestamp 1654583406
transform 1 0 8832 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_114
timestamp 1654583406
transform 1 0 5888 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_115
timestamp 1654583406
transform 1 0 20056 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_116
timestamp 1654583406
transform 1 0 12696 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_117
timestamp 1654583406
transform 1 0 9752 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_118
timestamp 1654583406
transform 1 0 21160 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_119
timestamp 1654583406
transform 1 0 11040 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_120
timestamp 1654583406
transform 1 0 10856 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_121
timestamp 1654583406
transform 1 0 7084 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_122
timestamp 1654583406
transform 1 0 14720 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_123
timestamp 1654583406
transform 1 0 21160 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_124
timestamp 1654583406
transform 1 0 17664 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_125
timestamp 1654583406
transform 1 0 22908 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_126
timestamp 1654583406
transform 1 0 22448 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_127
timestamp 1654583406
transform 1 0 21528 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_128
timestamp 1654583406
transform 1 0 15640 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_129
timestamp 1654583406
transform 1 0 7544 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_130
timestamp 1654583406
transform 1 0 22908 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_131
timestamp 1654583406
transform 1 0 21988 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_132
timestamp 1654583406
transform 1 0 17296 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_133
timestamp 1654583406
transform 1 0 16376 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_134
timestamp 1654583406
transform 1 0 10028 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_135
timestamp 1654583406
transform 1 0 9568 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_136
timestamp 1654583406
transform 1 0 21160 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_137
timestamp 1654583406
transform 1 0 16008 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_138
timestamp 1654583406
transform 1 0 15088 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_139
timestamp 1654583406
transform 1 0 8832 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_140
timestamp 1654583406
transform 1 0 22908 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_141
timestamp 1654583406
transform 1 0 17296 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_142
timestamp 1654583406
transform 1 0 11224 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_143
timestamp 1654583406
transform 1 0 6992 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_144
timestamp 1654583406
transform 1 0 18584 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_145
timestamp 1654583406
transform 1 0 11224 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_146
timestamp 1654583406
transform 1 0 10856 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_147
timestamp 1654583406
transform 1 0 5888 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_148
timestamp 1654583406
transform 1 0 22908 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_149
timestamp 1654583406
transform 1 0 22448 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_150
timestamp 1654583406
transform 1 0 19872 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_151
timestamp 1654583406
transform 1 0 10488 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_152
timestamp 1654583406
transform 1 0 7176 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_153
timestamp 1654583406
transform 1 0 6992 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_154
timestamp 1654583406
transform 1 0 6440 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_155
timestamp 1654583406
transform 1 0 21160 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_156
timestamp 1654583406
transform 1 0 18124 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_157
timestamp 1654583406
transform 1 0 19872 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_158
timestamp 1654583406
transform 1 0 7360 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_159
timestamp 1654583406
transform 1 0 6992 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_160
timestamp 1654583406
transform 1 0 20424 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_161
timestamp 1654583406
transform 1 0 18584 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_162
timestamp 1654583406
transform 1 0 8464 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_163
timestamp 1654583406
transform 1 0 19872 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_164
timestamp 1654583406
transform 1 0 14720 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_165
timestamp 1654583406
transform 1 0 21160 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_166
timestamp 1654583406
transform 1 0 18768 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_167
timestamp 1654583406
transform 1 0 19872 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_168
timestamp 1654583406
transform 1 0 5980 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_169
timestamp 1654583406
transform 1 0 13432 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_170
timestamp 1654583406
transform 1 0 6440 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_171
timestamp 1654583406
transform 1 0 19504 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_172
timestamp 1654583406
transform 1 0 12328 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_173
timestamp 1654583406
transform 1 0 8096 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_174
timestamp 1654583406
transform 1 0 7636 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_175
timestamp 1654583406
transform 1 0 5796 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_176
timestamp 1654583406
transform 1 0 21160 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_177
timestamp 1654583406
transform 1 0 19872 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_178
timestamp 1654583406
transform 1 0 18952 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_179
timestamp 1654583406
transform 1 0 18124 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_180
timestamp 1654583406
transform 1 0 13432 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_181
timestamp 1654583406
transform 1 0 12880 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_182
timestamp 1654583406
transform 1 0 9568 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_183
timestamp 1654583406
transform 1 0 8924 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_184
timestamp 1654583406
transform 1 0 8280 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_185
timestamp 1654583406
transform 1 0 6072 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0
timestamp 1654583406
transform 1 0 13616 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_1
timestamp 1654583406
transform 1 0 7820 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_2
timestamp 1654583406
transform 1 0 18492 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_3
timestamp 1654583406
transform 1 0 22724 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_4
timestamp 1654583406
transform 1 0 21804 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_5
timestamp 1654583406
transform 1 0 19872 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_6
timestamp 1654583406
transform 1 0 21620 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_7
timestamp 1654583406
transform 1 0 16468 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_8
timestamp 1654583406
transform 1 0 20240 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_9
timestamp 1654583406
transform 1 0 18492 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_10
timestamp 1654583406
transform 1 0 17572 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_11
timestamp 1654583406
transform 1 0 10212 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_12
timestamp 1654583406
transform 1 0 10856 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_13
timestamp 1654583406
transform 1 0 5796 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_14
timestamp 1654583406
transform 1 0 20240 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_15
timestamp 1654583406
transform 1 0 8464 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_16
timestamp 1654583406
transform 1 0 20240 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_17
timestamp 1654583406
transform 1 0 9752 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_18
timestamp 1654583406
transform 1 0 8464 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_19
timestamp 1654583406
transform 1 0 20240 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_20
timestamp 1654583406
transform 1 0 16008 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_21
timestamp 1654583406
transform 1 0 20240 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_22
timestamp 1654583406
transform 1 0 5796 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_23
timestamp 1654583406
transform 1 0 9476 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_24
timestamp 1654583406
transform 1 0 22816 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_25
timestamp 1654583406
transform 1 0 13616 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_26
timestamp 1654583406
transform 1 0 17480 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_27
timestamp 1654583406
transform 1 0 14628 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_28
timestamp 1654583406
transform 1 0 22816 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_29
timestamp 1654583406
transform 1 0 5888 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_30
timestamp 1654583406
transform 1 0 12328 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_31
timestamp 1654583406
transform 1 0 22816 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_32
timestamp 1654583406
transform 1 0 5888 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_33
timestamp 1654583406
transform 1 0 5796 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_34
timestamp 1654583406
transform 1 0 9292 0 1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_35
timestamp 1654583406
transform 1 0 21804 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_36
timestamp 1654583406
transform 1 0 22816 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_37
timestamp 1654583406
transform 1 0 5888 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_38
timestamp 1654583406
transform 1 0 14536 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_39
timestamp 1654583406
transform 1 0 7452 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_40
timestamp 1654583406
transform 1 0 22816 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_41
timestamp 1654583406
transform 1 0 15916 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_42
timestamp 1654583406
transform 1 0 15088 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_43
timestamp 1654583406
transform 1 0 5888 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_44
timestamp 1654583406
transform 1 0 21896 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_45
timestamp 1654583406
transform 1 0 21068 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_46
timestamp 1654583406
transform 1 0 18492 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_47
timestamp 1654583406
transform 1 0 17664 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_48
timestamp 1654583406
transform 1 0 5888 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_49
timestamp 1654583406
transform 1 0 17112 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_50
timestamp 1654583406
transform 1 0 12328 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_51
timestamp 1654583406
transform 1 0 9384 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_52
timestamp 1654583406
transform 1 0 5796 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_53
timestamp 1654583406
transform 1 0 15824 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_54
timestamp 1654583406
transform 1 0 22816 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_55
timestamp 1654583406
transform 1 0 11040 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_56
timestamp 1654583406
transform 1 0 6256 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_57
timestamp 1654583406
transform 1 0 19688 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_58
timestamp 1654583406
transform 1 0 6256 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_59
timestamp 1654583406
transform 1 0 5796 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_60
timestamp 1654583406
transform 1 0 22816 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_61
timestamp 1654583406
transform 1 0 13800 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_62
timestamp 1654583406
transform 1 0 7176 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_63
timestamp 1654583406
transform 1 0 6808 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_64
timestamp 1654583406
transform 1 0 17480 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_65
timestamp 1654583406
transform 1 0 5888 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_66
timestamp 1654583406
transform 1 0 22356 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_67
timestamp 1654583406
transform 1 0 14904 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_68
timestamp 1654583406
transform 1 0 5796 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_69
timestamp 1654583406
transform 1 0 22816 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_70
timestamp 1654583406
transform 1 0 15916 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_71
timestamp 1654583406
transform 1 0 12696 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_72
timestamp 1654583406
transform 1 0 10580 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_73
timestamp 1654583406
transform 1 0 7452 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_74
timestamp 1654583406
transform 1 0 18768 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_75
timestamp 1654583406
transform 1 0 18492 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_76
timestamp 1654583406
transform 1 0 17940 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_77
timestamp 1654583406
transform 1 0 17480 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_78
timestamp 1654583406
transform 1 0 15916 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_79
timestamp 1654583406
transform 1 0 10764 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_80
timestamp 1654583406
transform 1 0 8096 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_81
timestamp 1654583406
transform 1 0 5888 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_0
timestamp 1654583406
transform 1 0 20792 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_1
timestamp 1654583406
transform 1 0 6716 0 -1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_2
timestamp 1654583406
transform 1 0 19596 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_3
timestamp 1654583406
transform 1 0 22632 0 1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_4
timestamp 1654583406
transform 1 0 22632 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_5
timestamp 1654583406
transform 1 0 18308 0 1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_6
timestamp 1654583406
transform 1 0 15732 0 1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_7
timestamp 1654583406
transform 1 0 11224 0 -1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_8
timestamp 1654583406
transform 1 0 12512 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_9
timestamp 1654583406
transform 1 0 11224 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_10
timestamp 1654583406
transform 1 0 12512 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_11
timestamp 1654583406
transform 1 0 11040 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_12
timestamp 1654583406
transform 1 0 5796 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_13
timestamp 1654583406
transform 1 0 20056 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_14
timestamp 1654583406
transform 1 0 11868 0 -1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_15
timestamp 1654583406
transform 1 0 15548 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_16
timestamp 1654583406
transform 1 0 13616 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_17
timestamp 1654583406
transform 1 0 10028 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0
timestamp 1654583406
transform 1 0 10488 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1654583406
transform 1 0 14904 0 -1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1654583406
transform 1 0 8648 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3
timestamp 1654583406
transform 1 0 19136 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_4
timestamp 1654583406
transform 1 0 13984 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_5
timestamp 1654583406
transform 1 0 20056 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_0
timestamp 1654583406
transform 1 0 7268 0 -1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_1
timestamp 1654583406
transform -1 0 9568 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_2
timestamp 1654583406
transform -1 0 6992 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_3
timestamp 1654583406
transform -1 0 8280 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_4
timestamp 1654583406
transform -1 0 10672 0 1 17680
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_5
timestamp 1654583406
transform 1 0 8464 0 1 17680
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_6
timestamp 1654583406
transform 1 0 5980 0 -1 17680
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_7
timestamp 1654583406
transform 1 0 9752 0 -1 22032
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_8
timestamp 1654583406
transform -1 0 12236 0 -1 22032
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_9
timestamp 1654583406
transform 1 0 12420 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_10
timestamp 1654583406
transform -1 0 14996 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_11
timestamp 1654583406
transform -1 0 16100 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_12
timestamp 1654583406
transform 1 0 16836 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_13
timestamp 1654583406
transform -1 0 19872 0 1 19856
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_14
timestamp 1654583406
transform 1 0 20516 0 -1 19856
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_15
timestamp 1654583406
transform 1 0 5980 0 -1 13328
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1654583406
transform -1 0 10028 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1654583406
transform -1 0 10764 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2
timestamp 1654583406
transform 1 0 9108 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_3
timestamp 1654583406
transform 1 0 18216 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_4
timestamp 1654583406
transform 1 0 22356 0 1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_5
timestamp 1654583406
transform 1 0 22632 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_6
timestamp 1654583406
transform -1 0 22540 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_7
timestamp 1654583406
transform -1 0 6164 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_8
timestamp 1654583406
transform -1 0 14812 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_9
timestamp 1654583406
transform -1 0 12696 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_10
timestamp 1654583406
transform -1 0 10028 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0
timestamp 1654583406
transform -1 0 9108 0 -1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_1
timestamp 1654583406
transform -1 0 19504 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_2
timestamp 1654583406
transform -1 0 6532 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  sky130_fd_sc_hd__nand4_1_0
timestamp 1654583406
transform -1 0 7912 0 1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1654583406
transform 1 0 5980 0 1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1654583406
transform 1 0 5980 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1654583406
transform 1 0 22632 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1654583406
transform 1 0 22632 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_4
timestamp 1654583406
transform 1 0 19596 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_5
timestamp 1654583406
transform 1 0 12880 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_6
timestamp 1654583406
transform -1 0 10580 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_7
timestamp 1654583406
transform -1 0 8096 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_0
timestamp 1654583406
transform 1 0 8924 0 1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_0
timestamp 1654583406
transform 1 0 21988 0 -1 16592
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_1
timestamp 1654583406
transform 1 0 21988 0 -1 12240
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_2
timestamp 1654583406
transform 1 0 21712 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_3
timestamp 1654583406
transform -1 0 19596 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_4
timestamp 1654583406
transform 1 0 18124 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_5
timestamp 1654583406
transform 1 0 13984 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_6
timestamp 1654583406
transform 1 0 12328 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_7
timestamp 1654583406
transform 1 0 9016 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_8
timestamp 1654583406
transform 1 0 6532 0 -1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_9
timestamp 1654583406
transform -1 0 6440 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  sky130_fd_sc_hd__o21ai_1_0
timestamp 1654583406
transform 1 0 10120 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_0
timestamp 1654583406
transform -1 0 14536 0 -1 15504
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_1
timestamp 1654583406
transform -1 0 17388 0 -1 16592
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_2
timestamp 1654583406
transform -1 0 17388 0 -1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_3
timestamp 1654583406
transform -1 0 14168 0 -1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_4
timestamp 1654583406
transform 1 0 15732 0 -1 14416
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_5
timestamp 1654583406
transform -1 0 14168 0 -1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1654583406
transform 1 0 22540 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1654583406
transform 1 0 21252 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1654583406
transform 1 0 19964 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1654583406
transform 1 0 18676 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1654583406
transform 1 0 17388 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1654583406
transform 1 0 16100 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1654583406
transform 1 0 14812 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1654583406
transform 1 0 13524 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1654583406
transform 1 0 12236 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1654583406
transform 1 0 10948 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1654583406
transform 1 0 9660 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1654583406
transform 1 0 8372 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1654583406
transform 1 0 7084 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1654583406
transform 1 0 5796 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1654583406
transform 1 0 21252 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1654583406
transform 1 0 18676 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1654583406
transform 1 0 16100 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1654583406
transform 1 0 13524 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1654583406
transform 1 0 10948 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1654583406
transform 1 0 8372 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1654583406
transform 1 0 5796 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1654583406
transform 1 0 22540 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1654583406
transform 1 0 19964 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1654583406
transform 1 0 17388 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1654583406
transform 1 0 14812 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1654583406
transform 1 0 12236 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1654583406
transform 1 0 9660 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1654583406
transform 1 0 7084 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1654583406
transform 1 0 21252 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1654583406
transform 1 0 18676 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1654583406
transform 1 0 16100 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1654583406
transform 1 0 13524 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1654583406
transform 1 0 10948 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1654583406
transform 1 0 8372 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1654583406
transform 1 0 5796 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1654583406
transform 1 0 22540 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1654583406
transform 1 0 19964 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1654583406
transform 1 0 17388 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1654583406
transform 1 0 14812 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1654583406
transform 1 0 12236 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1654583406
transform 1 0 9660 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1654583406
transform 1 0 7084 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1654583406
transform 1 0 21252 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1654583406
transform 1 0 18676 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1654583406
transform 1 0 16100 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1654583406
transform 1 0 13524 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1654583406
transform 1 0 10948 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1654583406
transform 1 0 8372 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1654583406
transform 1 0 5796 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1654583406
transform 1 0 22540 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1654583406
transform 1 0 19964 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1654583406
transform 1 0 17388 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1654583406
transform 1 0 14812 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1654583406
transform 1 0 12236 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1654583406
transform 1 0 9660 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1654583406
transform 1 0 7084 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1654583406
transform 1 0 21252 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1654583406
transform 1 0 18676 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1654583406
transform 1 0 16100 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1654583406
transform 1 0 13524 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1654583406
transform 1 0 10948 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1654583406
transform 1 0 8372 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1654583406
transform 1 0 5796 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1654583406
transform 1 0 22540 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1654583406
transform 1 0 19964 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1654583406
transform 1 0 17388 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1654583406
transform 1 0 14812 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1654583406
transform 1 0 12236 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1654583406
transform 1 0 9660 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1654583406
transform 1 0 7084 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1654583406
transform 1 0 21252 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1654583406
transform 1 0 18676 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1654583406
transform 1 0 16100 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1654583406
transform 1 0 13524 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1654583406
transform 1 0 10948 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1654583406
transform 1 0 8372 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1654583406
transform 1 0 5796 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1654583406
transform 1 0 22540 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1654583406
transform 1 0 19964 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1654583406
transform 1 0 17388 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1654583406
transform 1 0 14812 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1654583406
transform 1 0 12236 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1654583406
transform 1 0 9660 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1654583406
transform 1 0 7084 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1654583406
transform 1 0 21252 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1654583406
transform 1 0 18676 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1654583406
transform 1 0 16100 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1654583406
transform 1 0 13524 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1654583406
transform 1 0 10948 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1654583406
transform 1 0 8372 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1654583406
transform 1 0 5796 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1654583406
transform 1 0 22540 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1654583406
transform 1 0 19964 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1654583406
transform 1 0 17388 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1654583406
transform 1 0 14812 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1654583406
transform 1 0 12236 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1654583406
transform 1 0 9660 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1654583406
transform 1 0 7084 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1654583406
transform 1 0 21252 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1654583406
transform 1 0 18676 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1654583406
transform 1 0 16100 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1654583406
transform 1 0 13524 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1654583406
transform 1 0 10948 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1654583406
transform 1 0 8372 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1654583406
transform 1 0 5796 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1654583406
transform 1 0 22540 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1654583406
transform 1 0 19964 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1654583406
transform 1 0 17388 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1654583406
transform 1 0 14812 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1654583406
transform 1 0 12236 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1654583406
transform 1 0 9660 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1654583406
transform 1 0 7084 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1654583406
transform 1 0 21252 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1654583406
transform 1 0 18676 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1654583406
transform 1 0 16100 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1654583406
transform 1 0 13524 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1654583406
transform 1 0 10948 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1654583406
transform 1 0 8372 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_118
timestamp 1654583406
transform 1 0 5796 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_119
timestamp 1654583406
transform 1 0 22540 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_120
timestamp 1654583406
transform 1 0 19964 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_121
timestamp 1654583406
transform 1 0 17388 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_122
timestamp 1654583406
transform 1 0 14812 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_123
timestamp 1654583406
transform 1 0 12236 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_124
timestamp 1654583406
transform 1 0 9660 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_125
timestamp 1654583406
transform 1 0 7084 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1654583406
transform 1 0 21252 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1654583406
transform 1 0 18676 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1654583406
transform 1 0 16100 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1654583406
transform 1 0 13524 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1654583406
transform 1 0 10948 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1654583406
transform 1 0 8372 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1654583406
transform 1 0 5796 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1654583406
transform 1 0 22540 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1654583406
transform 1 0 19964 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1654583406
transform 1 0 17388 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1654583406
transform 1 0 14812 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1654583406
transform 1 0 12236 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1654583406
transform 1 0 9660 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1654583406
transform 1 0 7084 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1654583406
transform 1 0 21252 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1654583406
transform 1 0 18676 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1654583406
transform 1 0 16100 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1654583406
transform 1 0 13524 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1654583406
transform 1 0 10948 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1654583406
transform 1 0 8372 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1654583406
transform 1 0 5796 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1654583406
transform 1 0 22540 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1654583406
transform 1 0 19964 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1654583406
transform 1 0 17388 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1654583406
transform 1 0 14812 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1654583406
transform 1 0 12236 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1654583406
transform 1 0 9660 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1654583406
transform 1 0 7084 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1654583406
transform 1 0 21252 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1654583406
transform 1 0 18676 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1654583406
transform 1 0 16100 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1654583406
transform 1 0 13524 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1654583406
transform 1 0 10948 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1654583406
transform 1 0 8372 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1654583406
transform 1 0 5796 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1654583406
transform 1 0 22540 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_162
timestamp 1654583406
transform 1 0 19964 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_163
timestamp 1654583406
transform 1 0 17388 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_164
timestamp 1654583406
transform 1 0 14812 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_165
timestamp 1654583406
transform 1 0 12236 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_166
timestamp 1654583406
transform 1 0 9660 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_167
timestamp 1654583406
transform 1 0 7084 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_168
timestamp 1654583406
transform 1 0 21252 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_169
timestamp 1654583406
transform 1 0 18676 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_170
timestamp 1654583406
transform 1 0 16100 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_171
timestamp 1654583406
transform 1 0 13524 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_172
timestamp 1654583406
transform 1 0 10948 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_173
timestamp 1654583406
transform 1 0 8372 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_174
timestamp 1654583406
transform 1 0 5796 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_175
timestamp 1654583406
transform 1 0 22540 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_176
timestamp 1654583406
transform 1 0 19964 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_177
timestamp 1654583406
transform 1 0 17388 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_178
timestamp 1654583406
transform 1 0 14812 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_179
timestamp 1654583406
transform 1 0 12236 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_180
timestamp 1654583406
transform 1 0 9660 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_181
timestamp 1654583406
transform 1 0 7084 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_182
timestamp 1654583406
transform 1 0 21252 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_183
timestamp 1654583406
transform 1 0 18676 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1654583406
transform 1 0 16100 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1654583406
transform 1 0 13524 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1654583406
transform 1 0 10948 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1654583406
transform 1 0 8372 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1654583406
transform 1 0 5796 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1654583406
transform 1 0 22540 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1654583406
transform 1 0 19964 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1654583406
transform 1 0 17388 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1654583406
transform 1 0 14812 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1654583406
transform 1 0 12236 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1654583406
transform 1 0 9660 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1654583406
transform 1 0 7084 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_196
timestamp 1654583406
transform 1 0 21252 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_197
timestamp 1654583406
transform 1 0 18676 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_198
timestamp 1654583406
transform 1 0 16100 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_199
timestamp 1654583406
transform 1 0 13524 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_200
timestamp 1654583406
transform 1 0 10948 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_201
timestamp 1654583406
transform 1 0 8372 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_202
timestamp 1654583406
transform 1 0 5796 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_203
timestamp 1654583406
transform 1 0 22540 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_204
timestamp 1654583406
transform 1 0 19964 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_205
timestamp 1654583406
transform 1 0 17388 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_206
timestamp 1654583406
transform 1 0 14812 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_207
timestamp 1654583406
transform 1 0 12236 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_208
timestamp 1654583406
transform 1 0 9660 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_209
timestamp 1654583406
transform 1 0 7084 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_210
timestamp 1654583406
transform 1 0 22540 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_211
timestamp 1654583406
transform 1 0 21252 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_212
timestamp 1654583406
transform 1 0 19964 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_213
timestamp 1654583406
transform 1 0 18676 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_214
timestamp 1654583406
transform 1 0 17388 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_215
timestamp 1654583406
transform 1 0 16100 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_216
timestamp 1654583406
transform 1 0 14812 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_217
timestamp 1654583406
transform 1 0 13524 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_218
timestamp 1654583406
transform 1 0 12236 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_219
timestamp 1654583406
transform 1 0 10948 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_220
timestamp 1654583406
transform 1 0 9660 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_221
timestamp 1654583406
transform 1 0 8372 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_222
timestamp 1654583406
transform 1 0 7084 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_223
timestamp 1654583406
transform 1 0 5796 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  sky130_fd_sc_hd__xnor2_1_0
timestamp 1654583406
transform 1 0 21896 0 -1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  sky130_fd_sc_hd__xnor2_1_1
timestamp 1654583406
transform -1 0 15916 0 1 5712
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1654583406
transform -1 0 7820 0 -1 22032
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1654583406
transform 1 0 8832 0 -1 22032
box -38 -48 682 592
<< labels >>
rlabel metal3 s 0 15354 160 15414 4 clk
port 1 nsew
rlabel metal3 s 0 104 160 164 4 rst_n
port 2 nsew
rlabel metal3 s 0 12304 160 12364 4 sclk
port 3 nsew
rlabel metal3 s 0 3154 160 3214 4 cs_n
port 4 nsew
rlabel metal3 s 0 6204 160 6264 4 data_in
port 5 nsew
rlabel metal3 s 0 9254 160 9314 4 data_out[11]
port 6 nsew
rlabel metal3 s 0 18404 160 18464 4 data_out[10]
port 7 nsew
rlabel metal3 s 0 21454 160 21514 4 data_out[9]
port 8 nsew
rlabel metal3 s 0 24504 160 24564 4 data_out[8]
port 9 nsew
rlabel metal3 s 0 27676 160 27736 4 data_out[7]
port 10 nsew
rlabel metal3 s 28636 27676 28796 27736 4 data_out[6]
port 11 nsew
rlabel metal3 s 28636 24260 28796 24320 4 data_out[5]
port 12 nsew
rlabel metal3 s 28636 20844 28796 20904 4 data_out[4]
port 13 nsew
rlabel metal3 s 28636 17428 28796 17488 4 data_out[3]
port 14 nsew
rlabel metal3 s 28636 13890 28796 13950 4 data_out[2]
port 15 nsew
rlabel metal3 s 28636 10474 28796 10534 4 data_out[1]
port 16 nsew
rlabel metal3 s 28636 7058 28796 7118 4 data_out[0]
port 17 nsew
rlabel metal3 s 28636 3642 28796 3702 4 new_data
port 18 nsew
rlabel metal3 s 28636 104 28796 164 4 serial_data_out
port 19 nsew
rlabel metal5 s 0 3852 620 4472 4 VSS
port 20 nsew
rlabel metal5 s 0 5092 620 5712 4 VDD
port 21 nsew
<< properties >>
string path 64.630 79.730 68.310 79.730 
<< end >>
