magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< nwell >>
rect -1489 -241 1489 241
<< pmoslvt >>
rect -1395 -140 -1275 140
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
rect 1275 -140 1395 140
<< pdiff >>
rect -1453 119 -1395 140
rect -1453 85 -1441 119
rect -1407 85 -1395 119
rect -1453 51 -1395 85
rect -1453 17 -1441 51
rect -1407 17 -1395 51
rect -1453 -17 -1395 17
rect -1453 -51 -1441 -17
rect -1407 -51 -1395 -17
rect -1453 -85 -1395 -51
rect -1453 -119 -1441 -85
rect -1407 -119 -1395 -85
rect -1453 -140 -1395 -119
rect -1275 119 -1217 140
rect -1275 85 -1263 119
rect -1229 85 -1217 119
rect -1275 51 -1217 85
rect -1275 17 -1263 51
rect -1229 17 -1217 51
rect -1275 -17 -1217 17
rect -1275 -51 -1263 -17
rect -1229 -51 -1217 -17
rect -1275 -85 -1217 -51
rect -1275 -119 -1263 -85
rect -1229 -119 -1217 -85
rect -1275 -140 -1217 -119
rect -1097 119 -1039 140
rect -1097 85 -1085 119
rect -1051 85 -1039 119
rect -1097 51 -1039 85
rect -1097 17 -1085 51
rect -1051 17 -1039 51
rect -1097 -17 -1039 17
rect -1097 -51 -1085 -17
rect -1051 -51 -1039 -17
rect -1097 -85 -1039 -51
rect -1097 -119 -1085 -85
rect -1051 -119 -1039 -85
rect -1097 -140 -1039 -119
rect -919 119 -861 140
rect -919 85 -907 119
rect -873 85 -861 119
rect -919 51 -861 85
rect -919 17 -907 51
rect -873 17 -861 51
rect -919 -17 -861 17
rect -919 -51 -907 -17
rect -873 -51 -861 -17
rect -919 -85 -861 -51
rect -919 -119 -907 -85
rect -873 -119 -861 -85
rect -919 -140 -861 -119
rect -741 119 -683 140
rect -741 85 -729 119
rect -695 85 -683 119
rect -741 51 -683 85
rect -741 17 -729 51
rect -695 17 -683 51
rect -741 -17 -683 17
rect -741 -51 -729 -17
rect -695 -51 -683 -17
rect -741 -85 -683 -51
rect -741 -119 -729 -85
rect -695 -119 -683 -85
rect -741 -140 -683 -119
rect -563 119 -505 140
rect -563 85 -551 119
rect -517 85 -505 119
rect -563 51 -505 85
rect -563 17 -551 51
rect -517 17 -505 51
rect -563 -17 -505 17
rect -563 -51 -551 -17
rect -517 -51 -505 -17
rect -563 -85 -505 -51
rect -563 -119 -551 -85
rect -517 -119 -505 -85
rect -563 -140 -505 -119
rect -385 119 -327 140
rect -385 85 -373 119
rect -339 85 -327 119
rect -385 51 -327 85
rect -385 17 -373 51
rect -339 17 -327 51
rect -385 -17 -327 17
rect -385 -51 -373 -17
rect -339 -51 -327 -17
rect -385 -85 -327 -51
rect -385 -119 -373 -85
rect -339 -119 -327 -85
rect -385 -140 -327 -119
rect -207 119 -149 140
rect -207 85 -195 119
rect -161 85 -149 119
rect -207 51 -149 85
rect -207 17 -195 51
rect -161 17 -149 51
rect -207 -17 -149 17
rect -207 -51 -195 -17
rect -161 -51 -149 -17
rect -207 -85 -149 -51
rect -207 -119 -195 -85
rect -161 -119 -149 -85
rect -207 -140 -149 -119
rect -29 119 29 140
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -140 29 -119
rect 149 119 207 140
rect 149 85 161 119
rect 195 85 207 119
rect 149 51 207 85
rect 149 17 161 51
rect 195 17 207 51
rect 149 -17 207 17
rect 149 -51 161 -17
rect 195 -51 207 -17
rect 149 -85 207 -51
rect 149 -119 161 -85
rect 195 -119 207 -85
rect 149 -140 207 -119
rect 327 119 385 140
rect 327 85 339 119
rect 373 85 385 119
rect 327 51 385 85
rect 327 17 339 51
rect 373 17 385 51
rect 327 -17 385 17
rect 327 -51 339 -17
rect 373 -51 385 -17
rect 327 -85 385 -51
rect 327 -119 339 -85
rect 373 -119 385 -85
rect 327 -140 385 -119
rect 505 119 563 140
rect 505 85 517 119
rect 551 85 563 119
rect 505 51 563 85
rect 505 17 517 51
rect 551 17 563 51
rect 505 -17 563 17
rect 505 -51 517 -17
rect 551 -51 563 -17
rect 505 -85 563 -51
rect 505 -119 517 -85
rect 551 -119 563 -85
rect 505 -140 563 -119
rect 683 119 741 140
rect 683 85 695 119
rect 729 85 741 119
rect 683 51 741 85
rect 683 17 695 51
rect 729 17 741 51
rect 683 -17 741 17
rect 683 -51 695 -17
rect 729 -51 741 -17
rect 683 -85 741 -51
rect 683 -119 695 -85
rect 729 -119 741 -85
rect 683 -140 741 -119
rect 861 119 919 140
rect 861 85 873 119
rect 907 85 919 119
rect 861 51 919 85
rect 861 17 873 51
rect 907 17 919 51
rect 861 -17 919 17
rect 861 -51 873 -17
rect 907 -51 919 -17
rect 861 -85 919 -51
rect 861 -119 873 -85
rect 907 -119 919 -85
rect 861 -140 919 -119
rect 1039 119 1097 140
rect 1039 85 1051 119
rect 1085 85 1097 119
rect 1039 51 1097 85
rect 1039 17 1051 51
rect 1085 17 1097 51
rect 1039 -17 1097 17
rect 1039 -51 1051 -17
rect 1085 -51 1097 -17
rect 1039 -85 1097 -51
rect 1039 -119 1051 -85
rect 1085 -119 1097 -85
rect 1039 -140 1097 -119
rect 1217 119 1275 140
rect 1217 85 1229 119
rect 1263 85 1275 119
rect 1217 51 1275 85
rect 1217 17 1229 51
rect 1263 17 1275 51
rect 1217 -17 1275 17
rect 1217 -51 1229 -17
rect 1263 -51 1275 -17
rect 1217 -85 1275 -51
rect 1217 -119 1229 -85
rect 1263 -119 1275 -85
rect 1217 -140 1275 -119
rect 1395 119 1453 140
rect 1395 85 1407 119
rect 1441 85 1453 119
rect 1395 51 1453 85
rect 1395 17 1407 51
rect 1441 17 1453 51
rect 1395 -17 1453 17
rect 1395 -51 1407 -17
rect 1441 -51 1453 -17
rect 1395 -85 1453 -51
rect 1395 -119 1407 -85
rect 1441 -119 1453 -85
rect 1395 -140 1453 -119
<< pdiffc >>
rect -1441 85 -1407 119
rect -1441 17 -1407 51
rect -1441 -51 -1407 -17
rect -1441 -119 -1407 -85
rect -1263 85 -1229 119
rect -1263 17 -1229 51
rect -1263 -51 -1229 -17
rect -1263 -119 -1229 -85
rect -1085 85 -1051 119
rect -1085 17 -1051 51
rect -1085 -51 -1051 -17
rect -1085 -119 -1051 -85
rect -907 85 -873 119
rect -907 17 -873 51
rect -907 -51 -873 -17
rect -907 -119 -873 -85
rect -729 85 -695 119
rect -729 17 -695 51
rect -729 -51 -695 -17
rect -729 -119 -695 -85
rect -551 85 -517 119
rect -551 17 -517 51
rect -551 -51 -517 -17
rect -551 -119 -517 -85
rect -373 85 -339 119
rect -373 17 -339 51
rect -373 -51 -339 -17
rect -373 -119 -339 -85
rect -195 85 -161 119
rect -195 17 -161 51
rect -195 -51 -161 -17
rect -195 -119 -161 -85
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect 161 85 195 119
rect 161 17 195 51
rect 161 -51 195 -17
rect 161 -119 195 -85
rect 339 85 373 119
rect 339 17 373 51
rect 339 -51 373 -17
rect 339 -119 373 -85
rect 517 85 551 119
rect 517 17 551 51
rect 517 -51 551 -17
rect 517 -119 551 -85
rect 695 85 729 119
rect 695 17 729 51
rect 695 -51 729 -17
rect 695 -119 729 -85
rect 873 85 907 119
rect 873 17 907 51
rect 873 -51 907 -17
rect 873 -119 907 -85
rect 1051 85 1085 119
rect 1051 17 1085 51
rect 1051 -51 1085 -17
rect 1051 -119 1085 -85
rect 1229 85 1263 119
rect 1229 17 1263 51
rect 1229 -51 1263 -17
rect 1229 -119 1263 -85
rect 1407 85 1441 119
rect 1407 17 1441 51
rect 1407 -51 1441 -17
rect 1407 -119 1441 -85
<< poly >>
rect -1373 221 -1297 237
rect -1373 205 -1352 221
rect -1395 187 -1352 205
rect -1318 205 -1297 221
rect -1195 221 -1119 237
rect -1195 205 -1174 221
rect -1318 187 -1275 205
rect -1395 140 -1275 187
rect -1217 187 -1174 205
rect -1140 205 -1119 221
rect -1017 221 -941 237
rect -1017 205 -996 221
rect -1140 187 -1097 205
rect -1217 140 -1097 187
rect -1039 187 -996 205
rect -962 205 -941 221
rect -839 221 -763 237
rect -839 205 -818 221
rect -962 187 -919 205
rect -1039 140 -919 187
rect -861 187 -818 205
rect -784 205 -763 221
rect -661 221 -585 237
rect -661 205 -640 221
rect -784 187 -741 205
rect -861 140 -741 187
rect -683 187 -640 205
rect -606 205 -585 221
rect -483 221 -407 237
rect -483 205 -462 221
rect -606 187 -563 205
rect -683 140 -563 187
rect -505 187 -462 205
rect -428 205 -407 221
rect -305 221 -229 237
rect -305 205 -284 221
rect -428 187 -385 205
rect -505 140 -385 187
rect -327 187 -284 205
rect -250 205 -229 221
rect -127 221 -51 237
rect -127 205 -106 221
rect -250 187 -207 205
rect -327 140 -207 187
rect -149 187 -106 205
rect -72 205 -51 221
rect 51 221 127 237
rect 51 205 72 221
rect -72 187 -29 205
rect -149 140 -29 187
rect 29 187 72 205
rect 106 205 127 221
rect 229 221 305 237
rect 229 205 250 221
rect 106 187 149 205
rect 29 140 149 187
rect 207 187 250 205
rect 284 205 305 221
rect 407 221 483 237
rect 407 205 428 221
rect 284 187 327 205
rect 207 140 327 187
rect 385 187 428 205
rect 462 205 483 221
rect 585 221 661 237
rect 585 205 606 221
rect 462 187 505 205
rect 385 140 505 187
rect 563 187 606 205
rect 640 205 661 221
rect 763 221 839 237
rect 763 205 784 221
rect 640 187 683 205
rect 563 140 683 187
rect 741 187 784 205
rect 818 205 839 221
rect 941 221 1017 237
rect 941 205 962 221
rect 818 187 861 205
rect 741 140 861 187
rect 919 187 962 205
rect 996 205 1017 221
rect 1119 221 1195 237
rect 1119 205 1140 221
rect 996 187 1039 205
rect 919 140 1039 187
rect 1097 187 1140 205
rect 1174 205 1195 221
rect 1297 221 1373 237
rect 1297 205 1318 221
rect 1174 187 1217 205
rect 1097 140 1217 187
rect 1275 187 1318 205
rect 1352 205 1373 221
rect 1352 187 1395 205
rect 1275 140 1395 187
rect -1395 -187 -1275 -140
rect -1395 -205 -1352 -187
rect -1373 -221 -1352 -205
rect -1318 -205 -1275 -187
rect -1217 -187 -1097 -140
rect -1217 -205 -1174 -187
rect -1318 -221 -1297 -205
rect -1373 -237 -1297 -221
rect -1195 -221 -1174 -205
rect -1140 -205 -1097 -187
rect -1039 -187 -919 -140
rect -1039 -205 -996 -187
rect -1140 -221 -1119 -205
rect -1195 -237 -1119 -221
rect -1017 -221 -996 -205
rect -962 -205 -919 -187
rect -861 -187 -741 -140
rect -861 -205 -818 -187
rect -962 -221 -941 -205
rect -1017 -237 -941 -221
rect -839 -221 -818 -205
rect -784 -205 -741 -187
rect -683 -187 -563 -140
rect -683 -205 -640 -187
rect -784 -221 -763 -205
rect -839 -237 -763 -221
rect -661 -221 -640 -205
rect -606 -205 -563 -187
rect -505 -187 -385 -140
rect -505 -205 -462 -187
rect -606 -221 -585 -205
rect -661 -237 -585 -221
rect -483 -221 -462 -205
rect -428 -205 -385 -187
rect -327 -187 -207 -140
rect -327 -205 -284 -187
rect -428 -221 -407 -205
rect -483 -237 -407 -221
rect -305 -221 -284 -205
rect -250 -205 -207 -187
rect -149 -187 -29 -140
rect -149 -205 -106 -187
rect -250 -221 -229 -205
rect -305 -237 -229 -221
rect -127 -221 -106 -205
rect -72 -205 -29 -187
rect 29 -187 149 -140
rect 29 -205 72 -187
rect -72 -221 -51 -205
rect -127 -237 -51 -221
rect 51 -221 72 -205
rect 106 -205 149 -187
rect 207 -187 327 -140
rect 207 -205 250 -187
rect 106 -221 127 -205
rect 51 -237 127 -221
rect 229 -221 250 -205
rect 284 -205 327 -187
rect 385 -187 505 -140
rect 385 -205 428 -187
rect 284 -221 305 -205
rect 229 -237 305 -221
rect 407 -221 428 -205
rect 462 -205 505 -187
rect 563 -187 683 -140
rect 563 -205 606 -187
rect 462 -221 483 -205
rect 407 -237 483 -221
rect 585 -221 606 -205
rect 640 -205 683 -187
rect 741 -187 861 -140
rect 741 -205 784 -187
rect 640 -221 661 -205
rect 585 -237 661 -221
rect 763 -221 784 -205
rect 818 -205 861 -187
rect 919 -187 1039 -140
rect 919 -205 962 -187
rect 818 -221 839 -205
rect 763 -237 839 -221
rect 941 -221 962 -205
rect 996 -205 1039 -187
rect 1097 -187 1217 -140
rect 1097 -205 1140 -187
rect 996 -221 1017 -205
rect 941 -237 1017 -221
rect 1119 -221 1140 -205
rect 1174 -205 1217 -187
rect 1275 -187 1395 -140
rect 1275 -205 1318 -187
rect 1174 -221 1195 -205
rect 1119 -237 1195 -221
rect 1297 -221 1318 -205
rect 1352 -205 1395 -187
rect 1352 -221 1373 -205
rect 1297 -237 1373 -221
<< polycont >>
rect -1352 187 -1318 221
rect -1174 187 -1140 221
rect -996 187 -962 221
rect -818 187 -784 221
rect -640 187 -606 221
rect -462 187 -428 221
rect -284 187 -250 221
rect -106 187 -72 221
rect 72 187 106 221
rect 250 187 284 221
rect 428 187 462 221
rect 606 187 640 221
rect 784 187 818 221
rect 962 187 996 221
rect 1140 187 1174 221
rect 1318 187 1352 221
rect -1352 -221 -1318 -187
rect -1174 -221 -1140 -187
rect -996 -221 -962 -187
rect -818 -221 -784 -187
rect -640 -221 -606 -187
rect -462 -221 -428 -187
rect -284 -221 -250 -187
rect -106 -221 -72 -187
rect 72 -221 106 -187
rect 250 -221 284 -187
rect 428 -221 462 -187
rect 606 -221 640 -187
rect 784 -221 818 -187
rect 962 -221 996 -187
rect 1140 -221 1174 -187
rect 1318 -221 1352 -187
<< locali >>
rect -1373 187 -1352 221
rect -1318 187 -1297 221
rect -1195 187 -1174 221
rect -1140 187 -1119 221
rect -1017 187 -996 221
rect -962 187 -941 221
rect -839 187 -818 221
rect -784 187 -763 221
rect -661 187 -640 221
rect -606 187 -585 221
rect -483 187 -462 221
rect -428 187 -407 221
rect -305 187 -284 221
rect -250 187 -229 221
rect -127 187 -106 221
rect -72 187 -51 221
rect 51 187 72 221
rect 106 187 127 221
rect 229 187 250 221
rect 284 187 305 221
rect 407 187 428 221
rect 462 187 483 221
rect 585 187 606 221
rect 640 187 661 221
rect 763 187 784 221
rect 818 187 839 221
rect 941 187 962 221
rect 996 187 1017 221
rect 1119 187 1140 221
rect 1174 187 1195 221
rect 1297 187 1318 221
rect 1352 187 1373 221
rect -1441 125 -1407 144
rect -1441 53 -1407 85
rect -1441 -17 -1407 17
rect -1441 -85 -1407 -53
rect -1441 -144 -1407 -125
rect -1263 125 -1229 144
rect -1263 53 -1229 85
rect -1263 -17 -1229 17
rect -1263 -85 -1229 -53
rect -1263 -144 -1229 -125
rect -1085 125 -1051 144
rect -1085 53 -1051 85
rect -1085 -17 -1051 17
rect -1085 -85 -1051 -53
rect -1085 -144 -1051 -125
rect -907 125 -873 144
rect -907 53 -873 85
rect -907 -17 -873 17
rect -907 -85 -873 -53
rect -907 -144 -873 -125
rect -729 125 -695 144
rect -729 53 -695 85
rect -729 -17 -695 17
rect -729 -85 -695 -53
rect -729 -144 -695 -125
rect -551 125 -517 144
rect -551 53 -517 85
rect -551 -17 -517 17
rect -551 -85 -517 -53
rect -551 -144 -517 -125
rect -373 125 -339 144
rect -373 53 -339 85
rect -373 -17 -339 17
rect -373 -85 -339 -53
rect -373 -144 -339 -125
rect -195 125 -161 144
rect -195 53 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -53
rect -195 -144 -161 -125
rect -17 125 17 144
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -144 17 -125
rect 161 125 195 144
rect 161 53 195 85
rect 161 -17 195 17
rect 161 -85 195 -53
rect 161 -144 195 -125
rect 339 125 373 144
rect 339 53 373 85
rect 339 -17 373 17
rect 339 -85 373 -53
rect 339 -144 373 -125
rect 517 125 551 144
rect 517 53 551 85
rect 517 -17 551 17
rect 517 -85 551 -53
rect 517 -144 551 -125
rect 695 125 729 144
rect 695 53 729 85
rect 695 -17 729 17
rect 695 -85 729 -53
rect 695 -144 729 -125
rect 873 125 907 144
rect 873 53 907 85
rect 873 -17 907 17
rect 873 -85 907 -53
rect 873 -144 907 -125
rect 1051 125 1085 144
rect 1051 53 1085 85
rect 1051 -17 1085 17
rect 1051 -85 1085 -53
rect 1051 -144 1085 -125
rect 1229 125 1263 144
rect 1229 53 1263 85
rect 1229 -17 1263 17
rect 1229 -85 1263 -53
rect 1229 -144 1263 -125
rect 1407 125 1441 144
rect 1407 53 1441 85
rect 1407 -17 1441 17
rect 1407 -85 1441 -53
rect 1407 -144 1441 -125
rect -1373 -221 -1352 -187
rect -1318 -221 -1297 -187
rect -1195 -221 -1174 -187
rect -1140 -221 -1119 -187
rect -1017 -221 -996 -187
rect -962 -221 -941 -187
rect -839 -221 -818 -187
rect -784 -221 -763 -187
rect -661 -221 -640 -187
rect -606 -221 -585 -187
rect -483 -221 -462 -187
rect -428 -221 -407 -187
rect -305 -221 -284 -187
rect -250 -221 -229 -187
rect -127 -221 -106 -187
rect -72 -221 -51 -187
rect 51 -221 72 -187
rect 106 -221 127 -187
rect 229 -221 250 -187
rect 284 -221 305 -187
rect 407 -221 428 -187
rect 462 -221 483 -187
rect 585 -221 606 -187
rect 640 -221 661 -187
rect 763 -221 784 -187
rect 818 -221 839 -187
rect 941 -221 962 -187
rect 996 -221 1017 -187
rect 1119 -221 1140 -187
rect 1174 -221 1195 -187
rect 1297 -221 1318 -187
rect 1352 -221 1373 -187
<< viali >>
rect -1352 187 -1318 221
rect -1174 187 -1140 221
rect -996 187 -962 221
rect -818 187 -784 221
rect -640 187 -606 221
rect -462 187 -428 221
rect -284 187 -250 221
rect -106 187 -72 221
rect 72 187 106 221
rect 250 187 284 221
rect 428 187 462 221
rect 606 187 640 221
rect 784 187 818 221
rect 962 187 996 221
rect 1140 187 1174 221
rect 1318 187 1352 221
rect -1441 119 -1407 125
rect -1441 91 -1407 119
rect -1441 51 -1407 53
rect -1441 19 -1407 51
rect -1441 -51 -1407 -19
rect -1441 -53 -1407 -51
rect -1441 -119 -1407 -91
rect -1441 -125 -1407 -119
rect -1263 119 -1229 125
rect -1263 91 -1229 119
rect -1263 51 -1229 53
rect -1263 19 -1229 51
rect -1263 -51 -1229 -19
rect -1263 -53 -1229 -51
rect -1263 -119 -1229 -91
rect -1263 -125 -1229 -119
rect -1085 119 -1051 125
rect -1085 91 -1051 119
rect -1085 51 -1051 53
rect -1085 19 -1051 51
rect -1085 -51 -1051 -19
rect -1085 -53 -1051 -51
rect -1085 -119 -1051 -91
rect -1085 -125 -1051 -119
rect -907 119 -873 125
rect -907 91 -873 119
rect -907 51 -873 53
rect -907 19 -873 51
rect -907 -51 -873 -19
rect -907 -53 -873 -51
rect -907 -119 -873 -91
rect -907 -125 -873 -119
rect -729 119 -695 125
rect -729 91 -695 119
rect -729 51 -695 53
rect -729 19 -695 51
rect -729 -51 -695 -19
rect -729 -53 -695 -51
rect -729 -119 -695 -91
rect -729 -125 -695 -119
rect -551 119 -517 125
rect -551 91 -517 119
rect -551 51 -517 53
rect -551 19 -517 51
rect -551 -51 -517 -19
rect -551 -53 -517 -51
rect -551 -119 -517 -91
rect -551 -125 -517 -119
rect -373 119 -339 125
rect -373 91 -339 119
rect -373 51 -339 53
rect -373 19 -339 51
rect -373 -51 -339 -19
rect -373 -53 -339 -51
rect -373 -119 -339 -91
rect -373 -125 -339 -119
rect -195 119 -161 125
rect -195 91 -161 119
rect -195 51 -161 53
rect -195 19 -161 51
rect -195 -51 -161 -19
rect -195 -53 -161 -51
rect -195 -119 -161 -91
rect -195 -125 -161 -119
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect 161 119 195 125
rect 161 91 195 119
rect 161 51 195 53
rect 161 19 195 51
rect 161 -51 195 -19
rect 161 -53 195 -51
rect 161 -119 195 -91
rect 161 -125 195 -119
rect 339 119 373 125
rect 339 91 373 119
rect 339 51 373 53
rect 339 19 373 51
rect 339 -51 373 -19
rect 339 -53 373 -51
rect 339 -119 373 -91
rect 339 -125 373 -119
rect 517 119 551 125
rect 517 91 551 119
rect 517 51 551 53
rect 517 19 551 51
rect 517 -51 551 -19
rect 517 -53 551 -51
rect 517 -119 551 -91
rect 517 -125 551 -119
rect 695 119 729 125
rect 695 91 729 119
rect 695 51 729 53
rect 695 19 729 51
rect 695 -51 729 -19
rect 695 -53 729 -51
rect 695 -119 729 -91
rect 695 -125 729 -119
rect 873 119 907 125
rect 873 91 907 119
rect 873 51 907 53
rect 873 19 907 51
rect 873 -51 907 -19
rect 873 -53 907 -51
rect 873 -119 907 -91
rect 873 -125 907 -119
rect 1051 119 1085 125
rect 1051 91 1085 119
rect 1051 51 1085 53
rect 1051 19 1085 51
rect 1051 -51 1085 -19
rect 1051 -53 1085 -51
rect 1051 -119 1085 -91
rect 1051 -125 1085 -119
rect 1229 119 1263 125
rect 1229 91 1263 119
rect 1229 51 1263 53
rect 1229 19 1263 51
rect 1229 -51 1263 -19
rect 1229 -53 1263 -51
rect 1229 -119 1263 -91
rect 1229 -125 1263 -119
rect 1407 119 1441 125
rect 1407 91 1441 119
rect 1407 51 1441 53
rect 1407 19 1441 51
rect 1407 -51 1441 -19
rect 1407 -53 1441 -51
rect 1407 -119 1441 -91
rect 1407 -125 1441 -119
rect -1352 -221 -1318 -187
rect -1174 -221 -1140 -187
rect -996 -221 -962 -187
rect -818 -221 -784 -187
rect -640 -221 -606 -187
rect -462 -221 -428 -187
rect -284 -221 -250 -187
rect -106 -221 -72 -187
rect 72 -221 106 -187
rect 250 -221 284 -187
rect 428 -221 462 -187
rect 606 -221 640 -187
rect 784 -221 818 -187
rect 962 -221 996 -187
rect 1140 -221 1174 -187
rect 1318 -221 1352 -187
<< metal1 >>
rect -1373 221 -1297 237
rect -1373 187 -1352 221
rect -1318 187 -1297 221
rect -1373 181 -1297 187
rect -1195 221 -1119 237
rect -1195 187 -1174 221
rect -1140 187 -1119 221
rect -1195 181 -1119 187
rect -1017 221 -941 237
rect -1017 187 -996 221
rect -962 187 -941 221
rect -1017 181 -941 187
rect -839 221 -763 237
rect -839 187 -818 221
rect -784 187 -763 221
rect -839 181 -763 187
rect -661 221 -585 237
rect -661 187 -640 221
rect -606 187 -585 221
rect -661 181 -585 187
rect -483 221 -407 237
rect -483 187 -462 221
rect -428 187 -407 221
rect -483 181 -407 187
rect -305 221 -229 237
rect -305 187 -284 221
rect -250 187 -229 221
rect -305 181 -229 187
rect -127 221 -51 237
rect -127 187 -106 221
rect -72 187 -51 221
rect -127 181 -51 187
rect 51 221 127 237
rect 51 187 72 221
rect 106 187 127 221
rect 51 181 127 187
rect 229 221 305 237
rect 229 187 250 221
rect 284 187 305 221
rect 229 181 305 187
rect 407 221 483 237
rect 407 187 428 221
rect 462 187 483 221
rect 407 181 483 187
rect 585 221 661 237
rect 585 187 606 221
rect 640 187 661 221
rect 585 181 661 187
rect 763 221 839 237
rect 763 187 784 221
rect 818 187 839 221
rect 763 181 839 187
rect 941 221 1017 237
rect 941 187 962 221
rect 996 187 1017 221
rect 941 181 1017 187
rect 1119 221 1195 237
rect 1119 187 1140 221
rect 1174 187 1195 221
rect 1119 181 1195 187
rect 1297 221 1373 237
rect 1297 187 1318 221
rect 1352 187 1373 221
rect 1297 181 1373 187
rect -1447 125 -1401 140
rect -1447 91 -1441 125
rect -1407 91 -1401 125
rect -1447 53 -1401 91
rect -1447 19 -1441 53
rect -1407 19 -1401 53
rect -1447 -19 -1401 19
rect -1447 -53 -1441 -19
rect -1407 -53 -1401 -19
rect -1447 -91 -1401 -53
rect -1447 -125 -1441 -91
rect -1407 -125 -1401 -91
rect -1447 -140 -1401 -125
rect -1269 125 -1223 140
rect -1269 91 -1263 125
rect -1229 91 -1223 125
rect -1269 53 -1223 91
rect -1269 19 -1263 53
rect -1229 19 -1223 53
rect -1269 -19 -1223 19
rect -1269 -53 -1263 -19
rect -1229 -53 -1223 -19
rect -1269 -91 -1223 -53
rect -1269 -125 -1263 -91
rect -1229 -125 -1223 -91
rect -1269 -140 -1223 -125
rect -1091 125 -1045 140
rect -1091 91 -1085 125
rect -1051 91 -1045 125
rect -1091 53 -1045 91
rect -1091 19 -1085 53
rect -1051 19 -1045 53
rect -1091 -19 -1045 19
rect -1091 -53 -1085 -19
rect -1051 -53 -1045 -19
rect -1091 -91 -1045 -53
rect -1091 -125 -1085 -91
rect -1051 -125 -1045 -91
rect -1091 -140 -1045 -125
rect -913 125 -867 140
rect -913 91 -907 125
rect -873 91 -867 125
rect -913 53 -867 91
rect -913 19 -907 53
rect -873 19 -867 53
rect -913 -19 -867 19
rect -913 -53 -907 -19
rect -873 -53 -867 -19
rect -913 -91 -867 -53
rect -913 -125 -907 -91
rect -873 -125 -867 -91
rect -913 -140 -867 -125
rect -735 125 -689 140
rect -735 91 -729 125
rect -695 91 -689 125
rect -735 53 -689 91
rect -735 19 -729 53
rect -695 19 -689 53
rect -735 -19 -689 19
rect -735 -53 -729 -19
rect -695 -53 -689 -19
rect -735 -91 -689 -53
rect -735 -125 -729 -91
rect -695 -125 -689 -91
rect -735 -140 -689 -125
rect -557 125 -511 140
rect -557 91 -551 125
rect -517 91 -511 125
rect -557 53 -511 91
rect -557 19 -551 53
rect -517 19 -511 53
rect -557 -19 -511 19
rect -557 -53 -551 -19
rect -517 -53 -511 -19
rect -557 -91 -511 -53
rect -557 -125 -551 -91
rect -517 -125 -511 -91
rect -557 -140 -511 -125
rect -379 125 -333 140
rect -379 91 -373 125
rect -339 91 -333 125
rect -379 53 -333 91
rect -379 19 -373 53
rect -339 19 -333 53
rect -379 -19 -333 19
rect -379 -53 -373 -19
rect -339 -53 -333 -19
rect -379 -91 -333 -53
rect -379 -125 -373 -91
rect -339 -125 -333 -91
rect -379 -140 -333 -125
rect -201 125 -155 140
rect -201 91 -195 125
rect -161 91 -155 125
rect -201 53 -155 91
rect -201 19 -195 53
rect -161 19 -155 53
rect -201 -19 -155 19
rect -201 -53 -195 -19
rect -161 -53 -155 -19
rect -201 -91 -155 -53
rect -201 -125 -195 -91
rect -161 -125 -155 -91
rect -201 -140 -155 -125
rect -23 125 23 140
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -140 23 -125
rect 155 125 201 140
rect 155 91 161 125
rect 195 91 201 125
rect 155 53 201 91
rect 155 19 161 53
rect 195 19 201 53
rect 155 -19 201 19
rect 155 -53 161 -19
rect 195 -53 201 -19
rect 155 -91 201 -53
rect 155 -125 161 -91
rect 195 -125 201 -91
rect 155 -140 201 -125
rect 333 125 379 140
rect 333 91 339 125
rect 373 91 379 125
rect 333 53 379 91
rect 333 19 339 53
rect 373 19 379 53
rect 333 -19 379 19
rect 333 -53 339 -19
rect 373 -53 379 -19
rect 333 -91 379 -53
rect 333 -125 339 -91
rect 373 -125 379 -91
rect 333 -140 379 -125
rect 511 125 557 140
rect 511 91 517 125
rect 551 91 557 125
rect 511 53 557 91
rect 511 19 517 53
rect 551 19 557 53
rect 511 -19 557 19
rect 511 -53 517 -19
rect 551 -53 557 -19
rect 511 -91 557 -53
rect 511 -125 517 -91
rect 551 -125 557 -91
rect 511 -140 557 -125
rect 689 125 735 140
rect 689 91 695 125
rect 729 91 735 125
rect 689 53 735 91
rect 689 19 695 53
rect 729 19 735 53
rect 689 -19 735 19
rect 689 -53 695 -19
rect 729 -53 735 -19
rect 689 -91 735 -53
rect 689 -125 695 -91
rect 729 -125 735 -91
rect 689 -140 735 -125
rect 867 125 913 140
rect 867 91 873 125
rect 907 91 913 125
rect 867 53 913 91
rect 867 19 873 53
rect 907 19 913 53
rect 867 -19 913 19
rect 867 -53 873 -19
rect 907 -53 913 -19
rect 867 -91 913 -53
rect 867 -125 873 -91
rect 907 -125 913 -91
rect 867 -140 913 -125
rect 1045 125 1091 140
rect 1045 91 1051 125
rect 1085 91 1091 125
rect 1045 53 1091 91
rect 1045 19 1051 53
rect 1085 19 1091 53
rect 1045 -19 1091 19
rect 1045 -53 1051 -19
rect 1085 -53 1091 -19
rect 1045 -91 1091 -53
rect 1045 -125 1051 -91
rect 1085 -125 1091 -91
rect 1045 -140 1091 -125
rect 1223 125 1269 140
rect 1223 91 1229 125
rect 1263 91 1269 125
rect 1223 53 1269 91
rect 1223 19 1229 53
rect 1263 19 1269 53
rect 1223 -19 1269 19
rect 1223 -53 1229 -19
rect 1263 -53 1269 -19
rect 1223 -91 1269 -53
rect 1223 -125 1229 -91
rect 1263 -125 1269 -91
rect 1223 -140 1269 -125
rect 1401 125 1447 140
rect 1401 91 1407 125
rect 1441 91 1447 125
rect 1401 53 1447 91
rect 1401 19 1407 53
rect 1441 19 1447 53
rect 1401 -19 1447 19
rect 1401 -53 1407 -19
rect 1441 -53 1447 -19
rect 1401 -91 1447 -53
rect 1401 -125 1407 -91
rect 1441 -125 1447 -91
rect 1401 -140 1447 -125
rect -1373 -187 -1297 -181
rect -1373 -221 -1352 -187
rect -1318 -221 -1297 -187
rect -1373 -237 -1297 -221
rect -1195 -187 -1119 -181
rect -1195 -221 -1174 -187
rect -1140 -221 -1119 -187
rect -1195 -237 -1119 -221
rect -1017 -187 -941 -181
rect -1017 -221 -996 -187
rect -962 -221 -941 -187
rect -1017 -237 -941 -221
rect -839 -187 -763 -181
rect -839 -221 -818 -187
rect -784 -221 -763 -187
rect -839 -237 -763 -221
rect -661 -187 -585 -181
rect -661 -221 -640 -187
rect -606 -221 -585 -187
rect -661 -237 -585 -221
rect -483 -187 -407 -181
rect -483 -221 -462 -187
rect -428 -221 -407 -187
rect -483 -237 -407 -221
rect -305 -187 -229 -181
rect -305 -221 -284 -187
rect -250 -221 -229 -187
rect -305 -237 -229 -221
rect -127 -187 -51 -181
rect -127 -221 -106 -187
rect -72 -221 -51 -187
rect -127 -237 -51 -221
rect 51 -187 127 -181
rect 51 -221 72 -187
rect 106 -221 127 -187
rect 51 -237 127 -221
rect 229 -187 305 -181
rect 229 -221 250 -187
rect 284 -221 305 -187
rect 229 -237 305 -221
rect 407 -187 483 -181
rect 407 -221 428 -187
rect 462 -221 483 -187
rect 407 -237 483 -221
rect 585 -187 661 -181
rect 585 -221 606 -187
rect 640 -221 661 -187
rect 585 -237 661 -221
rect 763 -187 839 -181
rect 763 -221 784 -187
rect 818 -221 839 -187
rect 763 -237 839 -221
rect 941 -187 1017 -181
rect 941 -221 962 -187
rect 996 -221 1017 -187
rect 941 -237 1017 -221
rect 1119 -187 1195 -181
rect 1119 -221 1140 -187
rect 1174 -221 1195 -187
rect 1119 -237 1195 -221
rect 1297 -187 1373 -181
rect 1297 -221 1318 -187
rect 1352 -221 1373 -187
rect 1297 -237 1373 -221
<< end >>
