magic
tech sky130A
magscale 1 2
timestamp 1652424873
<< error_p >>
rect -29 1451 29 1457
rect -29 1417 -17 1451
rect -29 1411 29 1417
rect -29 -1417 29 -1411
rect -29 -1451 -17 -1417
rect -29 -1457 29 -1451
<< nwell >>
rect -211 -1589 211 1589
<< pmos >>
rect -15 -1370 15 1370
<< pdiff >>
rect -73 1358 -15 1370
rect -73 -1358 -61 1358
rect -27 -1358 -15 1358
rect -73 -1370 -15 -1358
rect 15 1358 73 1370
rect 15 -1358 27 1358
rect 61 -1358 73 1358
rect 15 -1370 73 -1358
<< pdiffc >>
rect -61 -1358 -27 1358
rect 27 -1358 61 1358
<< nsubdiff >>
rect -175 1519 -79 1553
rect 79 1519 175 1553
rect -175 1457 -141 1519
rect 141 1457 175 1519
rect -175 -1519 -141 -1457
rect 141 -1519 175 -1457
rect -175 -1553 -79 -1519
rect 79 -1553 175 -1519
<< nsubdiffcont >>
rect -79 1519 79 1553
rect -175 -1457 -141 1457
rect 141 -1457 175 1457
rect -79 -1553 79 -1519
<< poly >>
rect -33 1451 33 1467
rect -33 1417 -17 1451
rect 17 1417 33 1451
rect -33 1401 33 1417
rect -15 1370 15 1401
rect -15 -1401 15 -1370
rect -33 -1417 33 -1401
rect -33 -1451 -17 -1417
rect 17 -1451 33 -1417
rect -33 -1467 33 -1451
<< polycont >>
rect -17 1417 17 1451
rect -17 -1451 17 -1417
<< locali >>
rect -175 1519 -79 1553
rect 79 1519 175 1553
rect -175 1457 -141 1519
rect 141 1457 175 1519
rect -33 1417 -17 1451
rect 17 1417 33 1451
rect -61 1358 -27 1374
rect -61 -1374 -27 -1358
rect 27 1358 61 1374
rect 27 -1374 61 -1358
rect -33 -1451 -17 -1417
rect 17 -1451 33 -1417
rect -175 -1519 -141 -1457
rect 141 -1519 175 -1457
rect -175 -1553 -79 -1519
rect 79 -1553 175 -1519
<< viali >>
rect -17 1417 17 1451
rect -61 -1358 -27 1358
rect 27 -1358 61 1358
rect -17 -1451 17 -1417
<< metal1 >>
rect -29 1451 29 1457
rect -29 1417 -17 1451
rect 17 1417 29 1451
rect -29 1411 29 1417
rect -67 1358 -21 1370
rect -67 -1358 -61 1358
rect -27 -1358 -21 1358
rect -67 -1370 -21 -1358
rect 21 1358 67 1370
rect 21 -1358 27 1358
rect 61 -1358 67 1358
rect 21 -1370 67 -1358
rect -29 -1417 29 -1411
rect -29 -1451 -17 -1417
rect 17 -1451 29 -1417
rect -29 -1457 29 -1451
<< properties >>
string FIXED_BBOX -158 -1536 158 1536
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 13.7 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
