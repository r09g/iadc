magic
tech sky130A
magscale 1 2
timestamp 1654408082
<< pwell >>
rect 610 59884 768 60125
rect 344 56750 640 56804
rect 344 56508 668 56750
rect 338 53104 671 53400
rect -27087 49194 -25523 49341
rect 39849 44543 45825 44690
rect 39849 43393 45825 43540
rect 39849 40868 45825 41000
rect 39849 40853 41395 40868
rect 41833 40853 45825 40868
rect 39849 39583 45825 39730
rect 5643 24033 5707 24097
rect 5284 9365 5337 9418
<< viali >>
rect 11189 73428 11223 76698
rect 377 53140 477 60758
rect -5624 50925 -155 51018
rect -26047 49413 -26013 49447
rect -26399 49359 -26176 49404
rect -26047 49327 -26013 49361
rect -4 47771 89 50741
rect 377 44350 477 45818
rect 39984 44783 40018 44817
rect 40603 44782 40637 44816
rect 41005 44776 41039 44810
rect 41161 44782 41195 44816
rect 40128 44702 40162 44736
rect 40905 44717 40939 44751
rect 41808 44596 41842 44936
rect 42537 44713 42936 44747
rect 43003 44648 43038 44818
rect 43281 44802 43315 44836
rect 43453 44802 43487 44836
rect 43625 44802 43659 44836
rect 43797 44802 43831 44836
rect 43969 44802 44003 44836
rect 44174 44802 44208 44836
rect 44351 44802 44385 44836
rect 44523 44802 44557 44836
rect 44695 44802 44729 44836
rect 44867 44802 44901 44836
rect 45039 44802 45073 44836
rect 45211 44802 45245 44836
rect 43253 44716 43408 44750
rect 39984 43633 40018 43667
rect 40603 43632 40637 43666
rect 41005 43626 41039 43660
rect 41161 43632 41195 43666
rect 40128 43552 40162 43586
rect 40905 43567 40939 43601
rect 41808 43446 41842 43786
rect 42537 43563 42936 43597
rect 43003 43498 43038 43668
rect 43281 43652 43315 43686
rect 43453 43652 43487 43686
rect 43625 43652 43659 43686
rect 43797 43652 43831 43686
rect 43969 43652 44003 43686
rect 44174 43652 44208 43686
rect 44351 43652 44385 43686
rect 44523 43652 44557 43686
rect 44695 43652 44729 43686
rect 44867 43652 44901 43686
rect 45039 43652 45073 43686
rect 45211 43652 45245 43686
rect 43253 43566 43408 43600
rect 377 40051 477 41343
rect 39984 41093 40018 41127
rect 40603 41092 40637 41126
rect 41005 41086 41039 41120
rect 41161 41092 41195 41126
rect 40128 41012 40162 41046
rect 40905 41027 40939 41061
rect 41808 40906 41842 41246
rect 42537 41023 42936 41057
rect 43003 40958 43038 41128
rect 43281 41112 43315 41146
rect 43453 41112 43487 41146
rect 43625 41112 43659 41146
rect 43797 41112 43831 41146
rect 43969 41112 44003 41146
rect 44174 41112 44208 41146
rect 44351 41112 44385 41146
rect 44523 41112 44557 41146
rect 44695 41112 44729 41146
rect 44867 41112 44901 41146
rect 45039 41112 45073 41146
rect 45211 41112 45245 41146
rect 43253 41026 43408 41060
rect 39984 39823 40018 39857
rect 40603 39822 40637 39856
rect 41005 39816 41039 39850
rect 41161 39822 41195 39856
rect -5637 39710 -168 39803
rect 40128 39742 40162 39776
rect 40905 39757 40939 39791
rect 41808 39636 41842 39976
rect 42537 39753 42936 39787
rect 43003 39688 43038 39858
rect 43281 39842 43315 39876
rect 43453 39842 43487 39876
rect 43625 39842 43659 39876
rect 43797 39842 43831 39876
rect 43969 39842 44003 39876
rect 44174 39842 44208 39876
rect 44351 39842 44385 39876
rect 44523 39842 44557 39876
rect 44695 39842 44729 39876
rect 44867 39842 44901 39876
rect 45039 39842 45073 39876
rect 45211 39842 45245 39876
rect 43253 39756 43408 39790
rect -31795 38846 -31761 39132
rect -31795 38202 -31761 38576
rect 59 10666 152 16135
rect 11274 14432 11367 16122
rect 11274 12989 11367 13953
rect 11274 11323 11367 12105
rect 6553 10409 11090 10502
rect 400 10021 1790 10121
rect 5748 10021 11698 10121
rect 13915 10021 21107 10121
rect 59 5602 159 9792
rect 59 374 159 2748
rect 21283 493 21383 9911
<< metal1 >>
rect -15420 77904 -15410 78140
rect -15174 77904 -15164 78140
rect -16859 73398 -16849 76723
rect -16748 73398 -16738 76723
rect -15353 75255 -15225 77904
rect 12596 77875 12606 78111
rect 12842 77875 12852 78111
rect 24646 77876 24656 78112
rect 24892 77876 24902 78112
rect 11177 76732 11367 76806
rect -15353 71958 -15225 74801
rect -13858 73404 -13848 76729
rect -13747 73404 -13737 76729
rect 11133 73392 11143 76732
rect 11271 73392 11367 76732
rect 11177 73320 11367 73392
rect 12660 73019 12778 77875
rect 14134 73405 14144 76745
rect 14272 73405 14282 76745
rect -16674 71738 -16664 71802
rect -16600 71738 -16590 71802
rect -15496 71734 -15486 71798
rect -15422 71734 -15412 71798
rect -15279 71741 -15269 71805
rect -15205 71741 -15195 71805
rect -14145 71738 -14135 71802
rect -14071 71738 -14061 71802
rect -16564 70234 -16554 70298
rect -16490 70234 -16480 70298
rect -15450 70220 -15440 70284
rect -15376 70220 -15366 70284
rect -15237 70221 -15227 70285
rect -15163 70221 -15153 70285
rect -14073 70221 -14063 70285
rect -13999 70221 -13989 70285
rect -15973 68105 -15963 68261
rect -15890 68105 -15880 68261
rect -15432 68166 -15422 68515
rect -15358 68166 -15348 68515
rect -14889 68108 -14879 68264
rect -14806 68108 -14796 68264
rect -16587 67549 -16577 67613
rect -16513 67549 -16503 67613
rect -15432 67543 -15422 67607
rect -15358 67543 -15348 67607
rect -14314 67554 -14304 67618
rect -14240 67554 -14230 67618
rect -16123 52998 -15995 66326
rect -14782 53600 -14654 66338
rect -9894 63338 -9884 63402
rect -9442 63338 -9432 63402
rect -9237 63338 -8980 63402
rect -8083 63340 -8073 63404
rect -7631 63340 -7621 63404
rect -9136 62888 -9072 63338
rect -7427 63332 -7188 63396
rect -6288 63336 -6278 63400
rect -5836 63336 -5826 63400
rect -5623 63337 -5392 63401
rect -7341 62888 -7277 63332
rect -6949 62966 -6939 63206
rect -6699 62966 -6689 63206
rect -6857 62888 -6793 62966
rect -5541 62888 -5477 63337
rect -4489 63334 -4479 63398
rect -4037 63334 -4027 63398
rect -3832 63335 -3572 63399
rect -2698 63338 -2688 63402
rect -2246 63338 -2236 63402
rect -2029 63339 -1794 63403
rect -3738 62888 -3674 63335
rect -1934 62888 -1870 63339
rect -896 63334 -886 63398
rect -444 63334 -434 63398
rect -221 63338 -2 63402
rect -138 63141 -74 63338
rect 747 63141 757 63232
rect -138 63077 757 63141
rect -138 62888 -74 63077
rect 747 62992 757 63077
rect 1287 62992 1297 63232
rect -9136 62824 -74 62888
rect -6867 54596 -6803 54597
rect -8567 54531 -8557 54595
rect -8493 54531 -8483 54595
rect -6876 54532 -6866 54596
rect -6802 54532 -6792 54596
rect -9714 54339 -9704 54403
rect -9462 54339 -9452 54403
rect -8557 54401 -8493 54531
rect -6867 54403 -6803 54532
rect -5171 54531 -5161 54595
rect -5097 54531 -5087 54595
rect -3375 54531 -3365 54595
rect -3301 54531 -3291 54595
rect -1546 54531 -1536 54595
rect -1472 54531 -1462 54595
rect -9230 54337 -8491 54401
rect -7919 54338 -7909 54402
rect -7667 54338 -7657 54402
rect -7435 54339 -6803 54403
rect -6119 54340 -6109 54404
rect -5867 54340 -5857 54404
rect -5161 54403 -5097 54531
rect -5632 54339 -5097 54403
rect -4321 54339 -4311 54403
rect -4069 54339 -4059 54403
rect -3365 54401 -3301 54531
rect -3832 54339 -3301 54401
rect -2523 54340 -2513 54404
rect -2271 54340 -2261 54404
rect -1536 54402 -1472 54531
rect -2027 54338 -1472 54402
rect -720 54339 -710 54403
rect -468 54339 -458 54403
rect -225 54340 176 54404
rect 240 54340 250 54404
rect -14793 53536 -14783 53600
rect -14655 53536 -14645 53600
rect -7560 53536 -7550 53600
rect -7486 53536 -7476 53600
rect -6999 53536 -6989 53600
rect -6861 53536 -6851 53600
rect -14782 53520 -14654 53536
rect 337 53121 347 60827
rect 519 53121 529 60827
rect 5400 58752 5410 58930
rect 5588 58752 5598 58930
rect 2037 57297 2047 57475
rect 2225 57297 2235 57475
rect 4037 57297 4047 57475
rect 4225 57297 4235 57475
rect 5400 55752 5410 55930
rect 5588 55752 5598 55930
rect 3997 53001 4007 53179
rect 4185 53001 4195 53179
rect -16123 52992 -9120 52998
rect -16123 52928 -9398 52992
rect -9270 52928 -9120 52992
rect -16123 52923 -9120 52928
rect 7715 51858 7725 52036
rect 7903 51858 7913 52036
rect -8864 51014 -8854 51249
rect -8770 51014 -8760 51249
rect -9408 50873 -9398 50937
rect -9270 50873 -8690 50937
rect -7544 50871 -6989 50935
rect -6861 50871 -6851 50935
rect -5698 50883 -5688 51066
rect -3888 51024 -3878 51066
rect -3372 51024 -3362 51074
rect -3888 51018 -3362 51024
rect -2536 51024 -2526 51074
rect -1665 51024 -1655 51064
rect -2536 51018 -1655 51024
rect -765 51024 -755 51064
rect -765 51018 -143 51024
rect -155 50925 -143 51018
rect -3888 50919 -3362 50925
rect -3888 50883 -3878 50919
rect -3372 50896 -3362 50919
rect -2536 50919 -1655 50925
rect -2536 50896 -2526 50919
rect -1665 50886 -1655 50919
rect -765 50919 -143 50925
rect -765 50886 -755 50919
rect -8884 50378 -8874 50791
rect -8780 50378 -8770 50791
rect -27080 49656 -27070 49720
rect -26726 49656 -26716 49720
rect -26059 49447 -26001 49468
rect -26059 49424 -26047 49447
rect -26013 49424 -26001 49447
rect -26418 49349 -26408 49413
rect -26157 49349 -26147 49413
rect -26070 49360 -26060 49424
rect -25996 49360 -25986 49424
rect -26059 49327 -26047 49360
rect -26013 49327 -26001 49360
rect -26059 49295 -26001 49327
rect -25994 49114 -25984 49178
rect -25640 49114 -25630 49178
rect -5942 47776 -5932 50720
rect -5748 47776 -5738 50720
rect -88 47752 -78 50774
rect 121 47752 131 50774
rect 10167 47617 10177 60836
rect 10551 47617 10561 60836
rect -27097 42779 -27087 43313
rect -26990 42779 -26980 43313
rect -13479 42997 -13469 43061
rect -13405 42997 -13395 43061
rect -27092 41002 -27082 42169
rect -26995 41002 -26985 42169
rect -27087 39476 -27077 40643
rect -26990 39476 -26980 40643
rect -31822 39007 -31812 39166
rect -31831 38973 -31812 39007
rect -31822 38827 -31812 38973
rect -31748 39007 -31738 39166
rect -31146 39126 -31082 39141
rect -31549 39092 -31082 39126
rect -31748 38973 -31710 39007
rect -31748 38827 -31738 38973
rect -31146 38886 -31082 39092
rect -31553 38852 -31082 38886
rect -31821 38407 -31811 38613
rect -31831 38373 -31811 38407
rect -31821 38141 -31811 38373
rect -31747 38407 -31737 38613
rect -31146 38570 -31082 38852
rect -31553 38536 -31082 38570
rect -31747 38373 -31703 38407
rect -31747 38141 -31737 38373
rect -31146 38256 -31082 38536
rect -29624 38349 -29614 38413
rect -29150 38349 -29140 38413
rect -31159 38242 -31030 38256
rect -31553 38208 -31030 38242
rect -31159 38192 -31030 38208
rect -30901 38192 -29704 38256
rect -27092 38232 -27082 39120
rect -26998 38232 -26988 39120
rect -35528 37332 -35518 37568
rect -35282 37475 -35272 37568
rect -35282 37411 -30199 37475
rect -30070 37411 -29696 37475
rect -35282 37332 -35272 37411
rect -29662 37259 -29652 37323
rect -29143 37259 -29133 37323
rect -27089 36465 -27079 37353
rect -26995 36465 -26985 37353
rect -27087 34985 -27077 36160
rect -26996 34985 -26986 36160
rect -18893 36124 -18883 39537
rect -18807 36124 -18797 39537
rect -27089 33498 -27079 34691
rect -27000 33498 -26990 34691
rect -27094 32365 -27084 32899
rect -27005 32365 -26995 32899
rect -13469 29329 -13405 42997
rect -12703 42334 -12693 42398
rect -12629 42334 -12619 42398
rect -12693 29752 -12629 42334
rect -5934 39819 -5924 46274
rect -5722 39819 -5712 46274
rect 93 45365 157 45366
rect -569 45313 157 45365
rect -4111 45129 -4101 45307
rect -3923 45129 -3913 45307
rect -1492 44281 -1482 44459
rect -1304 44281 -1294 44459
rect -6989 39805 -6861 39806
rect -9408 39741 -9398 39805
rect -9270 39741 -9260 39805
rect -6999 39741 -6989 39805
rect -6861 39741 -6851 39805
rect -9398 34676 -9270 39741
rect -9398 34612 -9369 34676
rect -9305 34612 -9270 34676
rect -9398 30305 -9270 34612
rect -6989 33179 -6861 39741
rect -5694 39666 -5684 39846
rect -148 39666 -138 39846
rect 93 38566 157 45313
rect 334 44318 344 45844
rect 558 44318 568 45844
rect 2122 44330 2132 44508
rect 2310 44330 2320 44508
rect 4122 44330 4132 44508
rect 4310 44330 4320 44508
rect 6122 44330 6132 44508
rect 6310 44330 6320 44508
rect 8122 44330 8132 44508
rect 8310 44330 8320 44508
rect 342 39855 352 41383
rect 512 39855 522 41383
rect 7082 41306 7200 43012
rect 2503 38642 2513 38881
rect 2595 38642 2605 38881
rect 5361 38568 5425 40438
rect 83 38502 93 38566
rect 157 38502 167 38566
rect 1220 38502 1230 38566
rect 1294 38502 1304 38566
rect 2439 38504 2626 38568
rect 2690 38504 2700 38568
rect 5351 38504 5361 38568
rect 5425 38504 5435 38568
rect 93 37651 157 38502
rect 2505 37996 2515 38420
rect 2614 37996 2624 38420
rect 5361 38155 5425 38504
rect 5351 38091 5361 38155
rect 5425 38091 5435 38155
rect 83 37587 93 37651
rect 157 37587 167 37651
rect 3417 37587 3427 37651
rect 3491 37587 3501 37651
rect 93 36816 157 37587
rect 2158 36898 2168 37149
rect 2232 36898 2242 37149
rect 2634 37143 2644 37207
rect 2708 37143 2718 37207
rect 2644 36816 2708 37143
rect 83 36752 93 36816
rect 157 36752 167 36816
rect 873 36752 883 36816
rect 947 36752 957 36816
rect 2240 36752 2708 36816
rect 93 36750 157 36752
rect 2159 36250 2169 36668
rect 2233 36250 2243 36668
rect 2928 36030 2938 36088
rect 3343 36030 3353 36088
rect 3427 35950 3491 37587
rect 6701 37207 6765 40449
rect 7082 39210 7318 41306
rect 10170 39867 10180 46128
rect 10551 39867 10561 46128
rect 12542 39210 12778 73019
rect 24656 66701 24892 77876
rect 24750 65741 24796 66701
rect 17420 64169 17430 64743
rect 17496 64169 17506 64743
rect 23948 64169 23958 64743
rect 24024 64169 24034 64743
rect 31564 64169 31574 64743
rect 31640 64169 31650 64743
rect 17965 62166 17975 62740
rect 18041 62166 18051 62740
rect 19053 62166 19063 62740
rect 19129 62166 19139 62740
rect 21229 62166 21239 62740
rect 21305 62166 21315 62740
rect 22317 62166 22327 62740
rect 22393 62166 22403 62740
rect 23405 62166 23415 62740
rect 23481 62166 23491 62740
rect 24493 62166 24503 62740
rect 24569 62166 24579 62740
rect 25581 62166 25591 62740
rect 25657 62166 25667 62740
rect 26669 62166 26679 62740
rect 26745 62166 26755 62740
rect 28845 62166 28855 62740
rect 28921 62166 28931 62740
rect 29933 62166 29943 62740
rect 30009 62166 30019 62740
rect 31021 62166 31031 62740
rect 31097 62166 31107 62740
rect 17420 60169 17430 60743
rect 17496 60169 17506 60743
rect 18508 60169 18518 60743
rect 18584 60169 18594 60743
rect 19596 60169 19606 60743
rect 19672 60169 19682 60743
rect 20684 60169 20694 60743
rect 20760 60169 20770 60743
rect 21772 60169 21782 60743
rect 21848 60169 21858 60743
rect 22860 60169 22870 60743
rect 22936 60169 22946 60743
rect 23948 60169 23958 60743
rect 24024 60169 24034 60743
rect 25036 60169 25046 60743
rect 25112 60169 25122 60743
rect 26124 60169 26134 60743
rect 26200 60169 26210 60743
rect 27212 60169 27222 60743
rect 27288 60169 27298 60743
rect 28300 60169 28310 60743
rect 28376 60169 28386 60743
rect 29388 60169 29398 60743
rect 29464 60169 29474 60743
rect 30476 60169 30486 60743
rect 30552 60169 30562 60743
rect 31564 60169 31574 60743
rect 31640 60169 31650 60743
rect 17965 58166 17975 58740
rect 18041 58166 18051 58740
rect 19053 58166 19063 58740
rect 19129 58166 19139 58740
rect 20141 58166 20151 58740
rect 20217 58166 20227 58740
rect 21229 58166 21239 58740
rect 21305 58166 21315 58740
rect 22317 58166 22327 58740
rect 22393 58166 22403 58740
rect 23405 58166 23415 58740
rect 23481 58166 23491 58740
rect 24493 58166 24503 58740
rect 24569 58166 24579 58740
rect 25581 58166 25591 58740
rect 25657 58166 25667 58740
rect 26669 58166 26679 58740
rect 26745 58166 26755 58740
rect 27757 58166 27767 58740
rect 27833 58166 27843 58740
rect 28845 58166 28855 58740
rect 28921 58166 28931 58740
rect 29933 58166 29943 58740
rect 30009 58166 30019 58740
rect 31021 58166 31031 58740
rect 31097 58166 31107 58740
rect 17420 56169 17430 56743
rect 17496 56169 17506 56743
rect 18508 56169 18518 56743
rect 18584 56169 18594 56743
rect 19596 56169 19606 56743
rect 19672 56169 19682 56743
rect 20684 56169 20694 56743
rect 20760 56169 20770 56743
rect 21772 56169 21782 56743
rect 21848 56169 21858 56743
rect 22860 56169 22870 56743
rect 22936 56169 22946 56743
rect 23948 56169 23958 56743
rect 24024 56169 24034 56743
rect 25036 56169 25046 56743
rect 25112 56169 25122 56743
rect 26124 56169 26134 56743
rect 26200 56169 26210 56743
rect 27212 56169 27222 56743
rect 27288 56169 27298 56743
rect 28300 56169 28310 56743
rect 28376 56169 28386 56743
rect 29388 56169 29398 56743
rect 29464 56169 29474 56743
rect 30476 56169 30486 56743
rect 30552 56169 30562 56743
rect 31564 56169 31574 56743
rect 31640 56169 31650 56743
rect 17965 54166 17975 54740
rect 18041 54166 18051 54740
rect 19053 54166 19063 54740
rect 19129 54166 19139 54740
rect 20141 54166 20151 54740
rect 20217 54166 20227 54740
rect 21229 54166 21239 54740
rect 21305 54166 21315 54740
rect 22317 54166 22327 54740
rect 22393 54166 22403 54740
rect 23405 54166 23415 54740
rect 23481 54166 23491 54740
rect 24493 54166 24503 54740
rect 24569 54166 24579 54740
rect 25581 54166 25591 54740
rect 25657 54166 25667 54740
rect 26669 54166 26679 54740
rect 26745 54166 26755 54740
rect 27757 54166 27767 54740
rect 27833 54166 27843 54740
rect 28845 54166 28855 54740
rect 28921 54166 28931 54740
rect 29933 54166 29943 54740
rect 30009 54166 30019 54740
rect 31021 54166 31031 54740
rect 31097 54166 31107 54740
rect 17420 52169 17430 52743
rect 17496 52169 17506 52743
rect 18508 52169 18518 52743
rect 18584 52169 18594 52743
rect 19596 52169 19606 52743
rect 19672 52169 19682 52743
rect 20684 52169 20694 52743
rect 20760 52169 20770 52743
rect 21772 52169 21782 52743
rect 21848 52169 21858 52743
rect 22860 52169 22870 52743
rect 22936 52169 22946 52743
rect 23948 52169 23958 52743
rect 24024 52169 24034 52743
rect 25036 52169 25046 52743
rect 25112 52169 25122 52743
rect 26124 52169 26134 52743
rect 26200 52169 26210 52743
rect 27212 52169 27222 52743
rect 27288 52169 27298 52743
rect 28300 52169 28310 52743
rect 28376 52169 28386 52743
rect 29388 52169 29398 52743
rect 29464 52169 29474 52743
rect 30476 52169 30486 52743
rect 30552 52169 30562 52743
rect 31564 52169 31574 52743
rect 31640 52169 31650 52743
rect 17965 50166 17975 50740
rect 18041 50166 18051 50740
rect 20141 50166 20151 50740
rect 20217 50166 20227 50740
rect 21229 50166 21239 50740
rect 21305 50166 21315 50740
rect 23405 50166 23415 50740
rect 23481 50166 23491 50740
rect 24493 50166 24503 50740
rect 24569 50166 24579 50740
rect 25581 50166 25591 50740
rect 25657 50166 25667 50740
rect 27757 50166 27767 50740
rect 27833 50166 27843 50740
rect 28845 50166 28855 50740
rect 28921 50166 28931 50740
rect 31021 50166 31031 50740
rect 31097 50166 31107 50740
rect 17420 48169 17430 48743
rect 17496 48169 17506 48743
rect 18508 48169 18518 48743
rect 18584 48169 18594 48743
rect 19596 48169 19606 48743
rect 19672 48169 19682 48743
rect 20684 48169 20694 48743
rect 20760 48169 20770 48743
rect 21772 48169 21782 48743
rect 21848 48169 21858 48743
rect 22860 48169 22870 48743
rect 22936 48169 22946 48743
rect 23948 48169 23958 48743
rect 24024 48169 24034 48743
rect 29388 48169 29398 48743
rect 29464 48169 29474 48743
rect 30476 48169 30486 48743
rect 30552 48169 30562 48743
rect 31564 48169 31574 48743
rect 31640 48169 31650 48743
rect 17965 46166 17975 46740
rect 18041 46166 18051 46740
rect 19053 46166 19063 46740
rect 19129 46166 19139 46740
rect 20141 46166 20151 46740
rect 20217 46166 20227 46740
rect 21229 46166 21239 46740
rect 21305 46166 21315 46740
rect 22317 46166 22327 46740
rect 22393 46166 22403 46740
rect 24493 46166 24503 46740
rect 24569 46166 24579 46740
rect 25581 46166 25591 46740
rect 25657 46166 25667 46740
rect 26669 46166 26679 46740
rect 26745 46166 26755 46740
rect 27757 46166 27767 46740
rect 27833 46166 27843 46740
rect 28845 46166 28855 46740
rect 28921 46166 28931 46740
rect 29933 46166 29943 46740
rect 30009 46166 30019 46740
rect 31021 46166 31031 46740
rect 31097 46166 31107 46740
rect 18235 45684 18245 45748
rect 18309 45684 18319 45748
rect 18781 45684 18791 45748
rect 18855 45684 18865 45748
rect 19327 45675 19337 45739
rect 19401 45675 19411 45739
rect 19872 45674 19882 45738
rect 19946 45674 19956 45738
rect 21507 45684 21517 45748
rect 21581 45684 21591 45748
rect 22041 45671 22051 45735
rect 22115 45671 22125 45735
rect 22588 45677 22598 45741
rect 22662 45677 22672 45741
rect 23133 45677 23143 45741
rect 23207 45677 23217 45741
rect 25853 45674 25863 45738
rect 25927 45674 25937 45738
rect 26396 45678 26406 45742
rect 26470 45678 26480 45742
rect 26938 45672 26948 45736
rect 27012 45672 27022 45736
rect 27495 45663 27505 45727
rect 27569 45663 27579 45727
rect 29119 45674 29129 45738
rect 29193 45674 29203 45738
rect 29663 45667 29673 45731
rect 29737 45667 29747 45731
rect 30213 45671 30223 45735
rect 30287 45671 30297 45735
rect 30746 45671 30756 45735
rect 30820 45671 30830 45735
rect 44744 45007 44754 45074
rect 45306 45007 45316 45074
rect 41802 44936 41848 44948
rect 39547 44827 39557 44891
rect 39621 44861 39631 44891
rect 39621 44827 40018 44861
rect 39972 44823 40018 44827
rect 39972 44817 40030 44823
rect 39972 44783 39984 44817
rect 40018 44783 40030 44817
rect 39972 44777 40030 44783
rect 40585 44778 40595 44830
rect 40647 44778 40657 44830
rect 40591 44776 40649 44778
rect 40985 44767 40995 44819
rect 41047 44767 41057 44819
rect 41142 44771 41152 44823
rect 41204 44771 41214 44823
rect 40116 44736 40174 44742
rect 40116 44702 40128 44736
rect 40162 44702 40174 44736
rect 40884 44710 40894 44762
rect 40946 44710 40956 44762
rect 40116 44701 40174 44702
rect 39547 44637 39557 44701
rect 39621 44696 40174 44701
rect 39621 44667 40162 44696
rect 39621 44637 39631 44667
rect 41802 44596 41808 44936
rect 41842 44753 41848 44936
rect 46284 44853 46294 44939
rect 43269 44836 43327 44842
rect 43441 44836 43499 44842
rect 43613 44836 43671 44842
rect 43785 44836 43843 44842
rect 43957 44836 44015 44842
rect 44162 44836 44220 44842
rect 44339 44836 44397 44842
rect 44511 44836 44569 44842
rect 44683 44836 44741 44842
rect 44855 44836 44913 44842
rect 45027 44836 45085 44842
rect 45199 44836 45257 44842
rect 45864 44836 46294 44853
rect 42997 44818 43044 44830
rect 41842 44747 42948 44753
rect 41842 44713 42537 44747
rect 42936 44713 42948 44747
rect 41842 44708 42948 44713
rect 41842 44596 41848 44708
rect 42525 44707 42948 44708
rect 42997 44648 43003 44818
rect 43038 44756 43044 44818
rect 43269 44802 43281 44836
rect 43315 44802 43453 44836
rect 43487 44802 43625 44836
rect 43659 44802 43797 44836
rect 43831 44802 43969 44836
rect 44003 44802 44174 44836
rect 44208 44802 44351 44836
rect 44385 44802 44523 44836
rect 44557 44802 44695 44836
rect 44729 44802 44867 44836
rect 44901 44802 45039 44836
rect 45073 44802 45211 44836
rect 45245 44802 46294 44836
rect 43269 44796 43327 44802
rect 43441 44796 43499 44802
rect 43613 44796 43671 44802
rect 43785 44796 43843 44802
rect 43957 44796 44015 44802
rect 44162 44796 44220 44802
rect 44339 44796 44397 44802
rect 44511 44796 44569 44802
rect 44683 44796 44741 44802
rect 44855 44796 44913 44802
rect 45027 44796 45085 44802
rect 45199 44796 45257 44802
rect 45864 44789 46294 44802
rect 43038 44750 43507 44756
rect 43038 44716 43253 44750
rect 43408 44716 43507 44750
rect 43038 44710 43507 44716
rect 43038 44648 43044 44710
rect 46284 44703 46294 44789
rect 46530 44703 46540 44939
rect 42997 44636 43044 44648
rect 41802 44584 41848 44596
rect 41506 44462 41516 44527
rect 41874 44462 41884 44527
rect 44756 43854 44766 43925
rect 45293 43854 45303 43925
rect 41802 43786 41848 43798
rect 39547 43677 39557 43741
rect 39621 43711 39631 43741
rect 39621 43677 40018 43711
rect 39972 43673 40018 43677
rect 39972 43667 40030 43673
rect 39972 43633 39984 43667
rect 40018 43633 40030 43667
rect 39972 43627 40030 43633
rect 40585 43628 40595 43680
rect 40647 43628 40657 43680
rect 40591 43626 40649 43628
rect 40985 43617 40995 43669
rect 41047 43617 41057 43669
rect 41142 43621 41152 43673
rect 41204 43621 41214 43673
rect 40116 43586 40174 43592
rect 40116 43552 40128 43586
rect 40162 43552 40174 43586
rect 40884 43560 40894 43612
rect 40946 43560 40956 43612
rect 40116 43551 40174 43552
rect 39547 43487 39557 43551
rect 39621 43546 40174 43551
rect 39621 43517 40162 43546
rect 39621 43487 39631 43517
rect 41802 43446 41808 43786
rect 41842 43603 41848 43786
rect 46272 43703 46282 43788
rect 43269 43686 43327 43692
rect 43441 43686 43499 43692
rect 43613 43686 43671 43692
rect 43785 43686 43843 43692
rect 43957 43686 44015 43692
rect 44162 43686 44220 43692
rect 44339 43686 44397 43692
rect 44511 43686 44569 43692
rect 44683 43686 44741 43692
rect 44855 43686 44913 43692
rect 45027 43686 45085 43692
rect 45199 43686 45257 43692
rect 45864 43686 46282 43703
rect 42997 43668 43044 43680
rect 41842 43597 42948 43603
rect 41842 43563 42537 43597
rect 42936 43563 42948 43597
rect 41842 43558 42948 43563
rect 41842 43446 41848 43558
rect 42525 43557 42948 43558
rect 42997 43498 43003 43668
rect 43038 43606 43044 43668
rect 43269 43652 43281 43686
rect 43315 43652 43453 43686
rect 43487 43652 43625 43686
rect 43659 43652 43797 43686
rect 43831 43652 43969 43686
rect 44003 43652 44174 43686
rect 44208 43652 44351 43686
rect 44385 43652 44523 43686
rect 44557 43652 44695 43686
rect 44729 43652 44867 43686
rect 44901 43652 45039 43686
rect 45073 43652 45211 43686
rect 45245 43652 46282 43686
rect 43269 43646 43327 43652
rect 43441 43646 43499 43652
rect 43613 43646 43671 43652
rect 43785 43646 43843 43652
rect 43957 43646 44015 43652
rect 44162 43646 44220 43652
rect 44339 43646 44397 43652
rect 44511 43646 44569 43652
rect 44683 43646 44741 43652
rect 44855 43646 44913 43652
rect 45027 43646 45085 43652
rect 45199 43646 45257 43652
rect 45864 43639 46282 43652
rect 43038 43600 43507 43606
rect 43038 43566 43253 43600
rect 43408 43566 43507 43600
rect 43038 43560 43507 43566
rect 43038 43498 43044 43560
rect 46272 43552 46282 43639
rect 46518 43552 46528 43788
rect 42997 43486 43044 43498
rect 41802 43434 41848 43446
rect 41504 43312 41514 43377
rect 41872 43312 41882 43377
rect 44746 41312 44756 41383
rect 45283 41312 45293 41383
rect 41802 41246 41848 41258
rect 39547 41137 39557 41201
rect 39621 41171 39631 41201
rect 39621 41137 40018 41171
rect 39972 41133 40018 41137
rect 39972 41127 40030 41133
rect 39972 41093 39984 41127
rect 40018 41093 40030 41127
rect 39972 41087 40030 41093
rect 40585 41088 40595 41140
rect 40647 41088 40657 41140
rect 40591 41086 40649 41088
rect 40985 41077 40995 41129
rect 41047 41077 41057 41129
rect 41142 41081 41152 41133
rect 41204 41081 41214 41133
rect 40116 41046 40174 41052
rect 40116 41012 40128 41046
rect 40162 41012 40174 41046
rect 40884 41020 40894 41072
rect 40946 41020 40956 41072
rect 40116 41011 40174 41012
rect 39547 40947 39557 41011
rect 39621 41006 40174 41011
rect 39621 40977 40162 41006
rect 39621 40947 39631 40977
rect 41802 40906 41808 41246
rect 41842 41063 41848 41246
rect 46130 41162 46140 41256
rect 43269 41146 43327 41152
rect 43441 41146 43499 41152
rect 43613 41146 43671 41152
rect 43785 41146 43843 41152
rect 43957 41146 44015 41152
rect 44162 41146 44220 41152
rect 44339 41146 44397 41152
rect 44511 41146 44569 41152
rect 44683 41146 44741 41152
rect 44855 41146 44913 41152
rect 45027 41146 45085 41152
rect 45199 41146 45257 41152
rect 45864 41146 46140 41162
rect 42997 41128 43044 41140
rect 41842 41057 42948 41063
rect 41842 41023 42537 41057
rect 42936 41023 42948 41057
rect 41842 41018 42948 41023
rect 41842 40906 41848 41018
rect 42525 41017 42948 41018
rect 42997 40958 43003 41128
rect 43038 41066 43044 41128
rect 43269 41112 43281 41146
rect 43315 41112 43453 41146
rect 43487 41112 43625 41146
rect 43659 41112 43797 41146
rect 43831 41112 43969 41146
rect 44003 41112 44174 41146
rect 44208 41112 44351 41146
rect 44385 41112 44523 41146
rect 44557 41112 44695 41146
rect 44729 41112 44867 41146
rect 44901 41112 45039 41146
rect 45073 41112 45211 41146
rect 45245 41112 46140 41146
rect 43269 41106 43327 41112
rect 43441 41106 43499 41112
rect 43613 41106 43671 41112
rect 43785 41106 43843 41112
rect 43957 41106 44015 41112
rect 44162 41106 44220 41112
rect 44339 41106 44397 41112
rect 44511 41106 44569 41112
rect 44683 41106 44741 41112
rect 44855 41106 44913 41112
rect 45027 41106 45085 41112
rect 45199 41106 45257 41112
rect 45864 41098 46140 41112
rect 43038 41060 43507 41066
rect 43038 41026 43253 41060
rect 43408 41026 43507 41060
rect 43038 41020 43507 41026
rect 46130 41020 46140 41098
rect 46376 41020 46386 41256
rect 43038 40958 43044 41020
rect 42997 40946 43044 40958
rect 41802 40894 41848 40906
rect 41422 40771 41432 40836
rect 41790 40771 41800 40836
rect 44746 40042 44756 40113
rect 45283 40042 45293 40113
rect 41802 39976 41848 39988
rect 39547 39867 39557 39931
rect 39621 39901 39631 39931
rect 39621 39867 40018 39901
rect 39972 39863 40018 39867
rect 39972 39857 40030 39863
rect 39972 39823 39984 39857
rect 40018 39823 40030 39857
rect 39972 39817 40030 39823
rect 40585 39818 40595 39870
rect 40647 39818 40657 39870
rect 40591 39816 40649 39818
rect 40985 39807 40995 39859
rect 41047 39807 41057 39859
rect 41142 39811 41152 39863
rect 41204 39811 41214 39863
rect 40116 39776 40174 39782
rect 40116 39742 40128 39776
rect 40162 39742 40174 39776
rect 40884 39750 40894 39802
rect 40946 39750 40956 39802
rect 40116 39741 40174 39742
rect 39547 39677 39557 39741
rect 39621 39736 40174 39741
rect 39621 39707 40162 39736
rect 39621 39677 39631 39707
rect 41802 39636 41808 39976
rect 41842 39793 41848 39976
rect 46101 39892 46111 39966
rect 43269 39876 43327 39882
rect 43441 39876 43499 39882
rect 43613 39876 43671 39882
rect 43785 39876 43843 39882
rect 43957 39876 44015 39882
rect 44162 39876 44220 39882
rect 44339 39876 44397 39882
rect 44511 39876 44569 39882
rect 44683 39876 44741 39882
rect 44855 39876 44913 39882
rect 45027 39876 45085 39882
rect 45199 39876 45257 39882
rect 45864 39876 46111 39892
rect 42997 39858 43044 39870
rect 41842 39787 42948 39793
rect 41842 39753 42537 39787
rect 42936 39753 42948 39787
rect 41842 39748 42948 39753
rect 41842 39636 41848 39748
rect 42525 39747 42948 39748
rect 42997 39688 43003 39858
rect 43038 39796 43044 39858
rect 43269 39842 43281 39876
rect 43315 39842 43453 39876
rect 43487 39842 43625 39876
rect 43659 39842 43797 39876
rect 43831 39842 43969 39876
rect 44003 39842 44174 39876
rect 44208 39842 44351 39876
rect 44385 39842 44523 39876
rect 44557 39842 44695 39876
rect 44729 39842 44867 39876
rect 44901 39842 45039 39876
rect 45073 39842 45211 39876
rect 45245 39842 46111 39876
rect 43269 39836 43327 39842
rect 43441 39836 43499 39842
rect 43613 39836 43671 39842
rect 43785 39836 43843 39842
rect 43957 39836 44015 39842
rect 44162 39836 44220 39842
rect 44339 39836 44397 39842
rect 44511 39836 44569 39842
rect 44683 39836 44741 39842
rect 44855 39836 44913 39842
rect 45027 39836 45085 39842
rect 45199 39836 45257 39842
rect 45864 39828 46111 39842
rect 43038 39790 43507 39796
rect 43038 39756 43253 39790
rect 43408 39756 43507 39790
rect 43038 39750 43507 39756
rect 43038 39688 43044 39750
rect 46101 39730 46111 39828
rect 46347 39730 46357 39966
rect 42997 39676 43044 39688
rect 41802 39624 41848 39636
rect 41420 39502 41430 39567
rect 41788 39502 41798 39567
rect 7072 38974 7082 39210
rect 7318 38974 7328 39210
rect 12532 38974 12542 39210
rect 12778 38974 12788 39210
rect 12660 38964 12778 38974
rect 7236 38155 7300 38168
rect 7226 38091 7236 38155
rect 7300 38091 7310 38155
rect 5419 37143 5429 37207
rect 5493 37143 5503 37207
rect 6691 37143 6701 37207
rect 6765 37143 6775 37207
rect 3572 36030 3582 36094
rect 3811 36030 3821 36094
rect 5045 36018 5055 36104
rect 5351 36018 5361 36104
rect 5429 35945 5493 37143
rect 7236 36107 7300 38091
rect 9418 37587 9428 37651
rect 9492 37587 9502 37651
rect 5564 36027 5574 36097
rect 5801 36027 5811 36097
rect 6926 36020 6936 36089
rect 7157 36020 7167 36089
rect 7373 36028 7383 36094
rect 7681 36028 7691 36094
rect 8911 36028 8921 36093
rect 9348 36028 9358 36093
rect 9428 35940 9492 37587
rect 9565 36023 9575 36091
rect 9802 36023 9812 36091
rect 5420 34956 5430 35020
rect 5494 34956 5504 35020
rect 7232 34954 7242 35018
rect 7306 34954 7316 35018
rect 3866 34780 4878 34844
rect 7854 34781 8873 34845
rect 3745 33850 3797 34654
rect 3735 33798 3745 33850
rect 3797 33798 3807 33850
rect -6989 33115 -6948 33179
rect -6884 33115 -6861 33179
rect -6989 31811 -6861 33115
rect -6999 31747 -6989 31811
rect -6861 31747 -6851 31811
rect -6989 31712 -6861 31747
rect 4354 30432 4418 34780
rect 5420 34361 5430 34425
rect 5494 34361 5504 34425
rect 7232 34361 7242 34425
rect 7306 34361 7316 34425
rect 5430 33561 5494 34361
rect 7242 34328 7306 34361
rect 7242 34264 7492 34328
rect 7428 33569 7492 34264
rect 5420 33497 5430 33561
rect 5494 33497 5504 33561
rect 7418 33505 7428 33569
rect 7492 33505 7502 33569
rect 5430 33480 5494 33497
rect 8328 30437 8392 34781
rect 9745 33850 9797 34662
rect 9735 33798 9745 33850
rect 9797 33798 9807 33850
rect 9745 33795 9797 33798
rect 4344 30368 4354 30432
rect 4418 30368 4428 30432
rect 8318 30373 8328 30437
rect 8392 30373 8402 30437
rect -9407 30241 -9397 30305
rect -9269 30241 -9259 30305
rect -9398 30201 -9270 30241
rect -12703 29688 -12693 29752
rect -12629 29688 -12619 29752
rect -30209 29159 -30199 29288
rect -30070 29159 -18523 29288
rect -18394 29159 -18384 29288
rect -13479 29265 -13469 29329
rect -13405 29265 -13395 29329
rect 1941 28744 1951 28808
rect 2079 28744 2089 28808
rect 7950 28782 7960 28846
rect 8024 28782 8034 28846
rect 1951 28644 2079 28744
rect -11888 28608 2079 28644
rect -11888 28544 -6086 28608
rect -5958 28544 2079 28608
rect -11888 28516 2079 28544
rect 3368 28595 3496 28627
rect 3368 28531 3399 28595
rect 3463 28531 3496 28595
rect -31040 27801 -31030 27930
rect -30901 27801 -19383 27930
rect -19254 27801 -19244 27930
rect -15722 27645 -15712 28098
rect -15613 27645 -15603 28098
rect -13993 28014 -13983 28066
rect -13931 28014 -13694 28066
rect -12399 27670 -12389 28076
rect -12316 27670 -12306 28076
rect -18326 27575 -18262 27600
rect -18336 27511 -18326 27575
rect -18262 27511 -18252 27575
rect -17645 27516 -17635 27644
rect -17507 27568 -17497 27644
rect -11888 27634 -11760 28516
rect -12206 27579 -11760 27634
rect -17507 27516 -17334 27568
rect -14916 27519 -14906 27571
rect -14854 27519 -13619 27571
rect -12491 27515 -11760 27579
rect -18326 27098 -18262 27511
rect -12206 27506 -11760 27515
rect -14414 27207 -14404 27259
rect -14352 27207 -13728 27259
rect -12404 27198 -12394 27427
rect -12297 27198 -12287 27427
rect -18336 27034 -18326 27098
rect -18262 27034 -18252 27098
rect -15239 27082 -14906 27083
rect -18891 26696 -18881 26760
rect -18817 26696 -18807 26760
rect -38200 26514 -38190 26611
rect -34856 26514 -34846 26611
rect -18881 25977 -18817 26696
rect -18892 25913 -18882 25977
rect -18818 25913 -18808 25977
rect -25459 25175 -25449 25482
rect -25369 25175 -25359 25482
rect -40603 24935 -40593 25171
rect -40357 25112 -40347 25171
rect -40357 24984 -32991 25112
rect -32863 24984 -26683 25112
rect -25335 24984 -24122 25112
rect -40357 24935 -40347 24984
rect -25462 24714 -25452 24945
rect -25365 24714 -25355 24945
rect -38192 23503 -38182 23605
rect -34852 23503 -34842 23605
rect -24250 21702 -24122 24984
rect -18881 24456 -18817 25913
rect -18891 24392 -18881 24456
rect -18817 24392 -18807 24456
rect -18326 24117 -18262 27034
rect -15242 27031 -14906 27082
rect -14854 27031 -14844 27083
rect -17266 26696 -17256 26760
rect -17192 26696 -17182 26760
rect -11912 26524 -10016 26588
rect -9888 26524 -9878 26588
rect -17645 26287 -17635 26415
rect -17507 26363 -17334 26415
rect -13993 26414 -13983 26466
rect -13931 26414 -13722 26466
rect -17507 26287 -17497 26363
rect -15735 26044 -15725 26281
rect -15636 26044 -15626 26281
rect -12406 26057 -12396 26486
rect -12301 26057 -12291 26486
rect -11912 25978 -11848 26524
rect -14916 25915 -14906 25967
rect -14854 25915 -13624 25967
rect -12478 25914 -11848 25978
rect -14414 25607 -14404 25659
rect -14352 25607 -13741 25659
rect -12394 25604 -12384 25823
rect -12321 25604 -12311 25823
rect 1952 25820 2080 25825
rect 1942 25756 1952 25820
rect 2080 25756 2090 25820
rect 1952 25448 2080 25756
rect -15737 25018 -15727 25447
rect -15632 25018 -15622 25447
rect -11886 25414 2080 25448
rect -11886 25350 -3501 25414
rect -3373 25350 2080 25414
rect -11886 25320 2080 25350
rect -17645 24874 -17635 25002
rect -17507 24926 -17497 25002
rect -17507 24874 -17339 24926
rect -13993 24814 -13983 24866
rect -13931 24814 -13749 24866
rect -12403 24458 -12393 24712
rect -12328 24458 -12318 24712
rect -15202 24389 -14908 24441
rect -14856 24389 -14850 24441
rect -11886 24408 -11758 25320
rect -14908 24369 -14850 24389
rect -12198 24376 -11758 24408
rect -14908 24317 -13620 24369
rect -12469 24312 -11758 24376
rect -12198 24280 -11758 24312
rect -18336 24053 -18326 24117
rect -18262 24053 -18252 24117
rect -17265 24053 -17255 24117
rect -17191 24053 -17181 24117
rect -14414 24007 -14404 24059
rect -14352 24007 -13733 24059
rect -12408 24003 -12398 24239
rect -12316 24003 -12306 24239
rect 3368 24101 3496 28531
rect 7960 25820 8024 28782
rect 9366 28592 9494 28632
rect 9366 28528 9399 28592
rect 9463 28528 9494 28592
rect 7950 25756 7960 25820
rect 8024 25756 8034 25820
rect 5705 24186 5715 24594
rect 5783 24186 5793 24594
rect 9366 24101 9494 28528
rect 3368 24037 3399 24101
rect 3463 24037 3496 24101
rect -17645 23645 -17635 23773
rect -17507 23721 -17338 23773
rect -17507 23645 -17497 23721
rect -15735 23405 -15725 23637
rect -15658 23405 -15648 23637
rect 3368 23415 3496 24037
rect 5633 24033 5643 24097
rect 5707 24033 5717 24097
rect 7007 24037 7017 24101
rect 7081 24037 7091 24101
rect 9366 24037 9399 24101
rect 9463 24037 9494 24101
rect 42846 24065 42856 24174
rect 46190 24065 46200 24174
rect 5724 23395 5788 23661
rect 9366 23423 9494 24037
rect 35142 23802 35152 23866
rect 35216 23802 35226 23866
rect 37809 23492 37819 23611
rect 37892 23492 37902 23611
rect 39336 23493 39346 23714
rect 39420 23493 39430 23714
rect 2550 23328 2850 23392
rect 3860 23356 9002 23395
rect 3860 23331 8787 23356
rect -13993 23214 -13983 23266
rect -13931 23214 -13709 23266
rect -12399 22857 -12389 23277
rect -12319 22857 -12309 23277
rect 2550 23063 2614 23328
rect 8777 23246 8787 23331
rect 8943 23331 9002 23356
rect 8943 23246 8953 23331
rect 10068 23326 10266 23390
rect 10202 23063 10266 23326
rect 13272 23295 33935 23423
rect 39446 23303 39682 23431
rect 2540 22999 2550 23063
rect 2614 22999 2624 23063
rect 10192 22999 10202 23063
rect 10266 22999 10276 23063
rect -12465 22773 -11601 22776
rect -14918 22719 -14908 22771
rect -14856 22719 -13614 22771
rect -12460 22712 -11601 22773
rect -11473 22712 -11463 22776
rect -14414 22407 -14404 22459
rect -14352 22407 -13740 22459
rect -12401 22399 -12391 22624
rect -12323 22399 -12313 22624
rect 3395 22101 3459 22106
rect -24250 21671 -5931 21702
rect -24250 21607 -6086 21671
rect -5958 21607 -5931 21671
rect -24250 21574 -5931 21607
rect -24284 20809 -3339 20842
rect -24284 20745 -3501 20809
rect -3373 20745 -3339 20809
rect -24284 20714 -3339 20745
rect -38178 18987 -38168 19065
rect -34861 18987 -34851 19065
rect -40606 17394 -40596 17630
rect -40360 17582 -40350 17630
rect -25462 17627 -25452 17922
rect -25387 17627 -25377 17922
rect -40360 17454 -31130 17582
rect -31002 17454 -26675 17582
rect -24284 17579 -24156 20714
rect -454 19981 -444 20109
rect -380 19981 -370 20109
rect -444 18993 -380 19981
rect 1674 19282 1684 19410
rect 1748 19282 1812 19410
rect -40360 17394 -40350 17454
rect -25357 17451 -24156 17579
rect -821 17525 -757 17735
rect 223 17708 233 17772
rect 297 17708 307 17772
rect -831 17461 -821 17525
rect -757 17461 -747 17525
rect -25460 17169 -25450 17404
rect -25378 17169 -25368 17404
rect -445 17221 -381 17690
rect 1684 17221 1812 19282
rect 3361 19346 3489 22101
rect 4387 21985 4397 22037
rect 4449 21985 4459 22037
rect 8218 21985 8228 22037
rect 8280 21985 8290 22037
rect 4397 20945 4449 21985
rect 8228 20945 8280 21985
rect 4387 20893 4397 20945
rect 4449 20893 4459 20945
rect 8218 20893 8228 20945
rect 8280 20893 8290 20945
rect 8228 20883 8280 20893
rect 9363 20109 9491 22105
rect 5384 19981 5394 20109
rect 5458 19981 5468 20109
rect 9363 19981 9394 20109
rect 9458 19981 9491 20109
rect 3361 19282 3395 19346
rect 3459 19282 3489 19346
rect 3051 19042 3061 19106
rect 3125 19042 3135 19106
rect 3361 19072 3489 19282
rect 3883 18987 4359 19051
rect 4847 19027 4857 19173
rect 5194 19027 5204 19173
rect 5394 19098 5458 19981
rect 7384 19282 7394 19410
rect 7458 19282 7468 19410
rect 5882 18991 6291 19055
rect 7075 19042 7085 19106
rect 7149 19042 7159 19106
rect 7394 19103 7458 19282
rect -455 17093 -445 17221
rect -381 17093 -371 17221
rect 1674 17093 1684 17221
rect 1748 17093 1812 17221
rect 3393 16866 3457 17769
rect 4295 17289 4359 18987
rect 4285 17225 4295 17289
rect 4359 17225 4369 17289
rect 5393 16866 5457 17768
rect 6227 17289 6291 18991
rect 7877 18989 8344 19053
rect 8971 19042 8981 19106
rect 9045 19042 9055 19106
rect 9363 19074 9491 19981
rect 13272 19716 13347 23295
rect 37809 22946 37819 23194
rect 37905 22946 37915 23194
rect 39325 22952 39335 23200
rect 39421 22952 39431 23200
rect 35090 22610 35100 22790
rect 35280 22610 35290 22790
rect 35750 22668 35760 22730
rect 36021 22668 36031 22730
rect 39554 22677 39682 23303
rect 47546 22677 47556 22734
rect 39554 22549 47556 22677
rect 37816 22151 37826 22280
rect 37896 22151 37906 22280
rect 39336 22167 39346 22388
rect 39420 22167 39430 22388
rect 13877 21996 13887 22124
rect 13951 21996 33915 22124
rect 39556 22107 39684 22549
rect 47546 22498 47556 22549
rect 47792 22498 47802 22734
rect 39464 21979 39684 22107
rect 37804 21621 37814 21823
rect 37899 21621 37909 21823
rect 39331 21586 39341 21834
rect 39427 21586 39437 21834
rect 35142 21521 35152 21585
rect 35216 21521 35226 21585
rect 42844 21069 42854 21178
rect 46188 21069 46198 21178
rect 14678 20963 14688 21027
rect 14752 20963 14762 21027
rect 14688 20497 14752 20963
rect 23660 20152 23670 20216
rect 23734 20152 23744 20216
rect 14686 19278 14750 19343
rect 23679 19318 23689 19382
rect 23753 19318 23763 19382
rect 14676 19214 14686 19278
rect 14750 19214 14760 19278
rect 9877 18994 10232 19058
rect 10296 18994 10306 19058
rect 8280 18718 8344 18989
rect 8270 18654 8280 18718
rect 8344 18654 8354 18718
rect 13564 18624 13574 18688
rect 13638 18624 14728 18688
rect 23648 18364 23658 18428
rect 23722 18364 23732 18428
rect 13877 17983 13887 18047
rect 13951 17983 13961 18047
rect 7393 17359 7457 17775
rect 9396 17359 9460 17774
rect 14679 17485 14689 17549
rect 14753 17485 14763 17549
rect 23679 17488 23689 17552
rect 23753 17488 23763 17552
rect 6217 17225 6227 17289
rect 6291 17225 6301 17289
rect 7383 17231 7393 17359
rect 7457 17231 7467 17359
rect 9386 17231 9396 17359
rect 9460 17231 9470 17359
rect 13875 17231 13885 17359
rect 13949 17231 13959 17359
rect 14680 17019 14690 17083
rect 14754 17019 14764 17083
rect 14690 16894 14754 17019
rect 3383 16738 3393 16866
rect 3457 16738 3467 16866
rect 5383 16738 5393 16866
rect 5457 16738 5467 16866
rect 13267 16738 13277 16866
rect 13341 16738 13351 16866
rect 23062 16656 23727 16720
rect -3926 16288 -3862 16297
rect -3936 16224 -3926 16288
rect -3862 16224 -3852 16288
rect 241 16238 251 16446
rect 11139 16238 11149 16446
rect -38184 15987 -38174 16075
rect -34852 15987 -34842 16075
rect -5787 15708 -3049 15709
rect -5796 15644 -5786 15708
rect -5722 15645 -3049 15708
rect -5722 15644 -5712 15645
rect -3113 15543 -3049 15645
rect -3927 15083 -3914 15135
rect -3862 15083 -2971 15135
rect -1824 15084 -678 15136
rect -626 15084 -616 15136
rect -3154 14719 -3144 14998
rect -3061 14719 -3051 14998
rect -25527 14157 -25517 14446
rect -25444 14157 -25434 14446
rect -4912 14236 -4902 14446
rect -4832 14236 -4822 14446
rect -33001 13974 -32991 14102
rect -32863 13974 -26755 14102
rect -25361 14073 -18140 14105
rect -13074 14077 -13064 14141
rect -13000 14077 -6544 14141
rect -6480 14077 -6287 14141
rect -4816 14087 -3914 14139
rect -3862 14087 -3852 14139
rect -25592 14009 -18223 14073
rect -18159 14009 -18140 14073
rect -25361 13977 -18140 14009
rect -25528 13690 -25518 13925
rect -25446 13690 -25436 13925
rect -4927 13706 -4917 13998
rect -4833 13706 -4823 13998
rect -6554 12828 -6544 12892
rect -6480 12828 -5851 12892
rect -5787 12828 -5777 12892
rect -1818 12726 -1808 13133
rect -1725 12726 -1715 13133
rect -3914 12635 -3027 12636
rect -3924 12583 -3914 12635
rect -3862 12583 -3027 12635
rect -1725 12585 -279 12637
rect -227 12585 -217 12637
rect -1785 12345 -1498 12409
rect -1434 12345 -1424 12409
rect -5861 12155 -5851 12219
rect -5787 12155 -5777 12219
rect -1798 11529 -1703 11530
rect -1798 11140 -1759 11529
rect -1693 11140 -1683 11529
rect -1798 11139 -1703 11140
rect -3425 10982 -3415 11034
rect -3363 10982 -3032 11034
rect -1724 10983 -279 11035
rect -227 10983 -217 11035
rect -5855 10891 -5845 10943
rect -5793 10891 -5783 10943
rect -6172 10758 -6162 10833
rect -5937 10758 -5927 10833
rect -5717 10751 -5707 10838
rect -5401 10751 -5391 10838
rect -1803 10719 -1498 10783
rect -1434 10719 -1424 10783
rect 18 10640 28 16189
rect 187 10640 197 16189
rect 5468 14421 5478 14599
rect 5656 14421 5666 14599
rect 11229 14426 11239 16184
rect 11399 14426 11409 16184
rect 14675 15689 14685 15753
rect 14749 15689 14759 15753
rect 23062 15496 23126 16656
rect 23676 15724 23686 15788
rect 23750 15724 23760 15788
rect 20918 15432 20928 15496
rect 20992 15432 23763 15496
rect 14680 15164 14690 15228
rect 14754 15164 14764 15228
rect 14690 15130 14754 15164
rect 23699 15092 23763 15432
rect 11268 14420 11373 14426
rect 11268 13954 11373 13965
rect 11247 12990 11257 13954
rect 11384 12990 11394 13954
rect 14675 13901 14685 13965
rect 14749 13901 14759 13965
rect 23676 13933 23686 13997
rect 23750 13933 23760 13997
rect 14680 13464 14690 13528
rect 14754 13464 14764 13528
rect 14690 13327 14754 13464
rect 11268 12989 11274 12990
rect 11367 12989 11373 12990
rect 11268 12977 11373 12989
rect 23675 12942 23685 13006
rect 23749 12942 23759 13006
rect 4620 11802 4630 11980
rect 4808 11802 4818 11980
rect 11233 11316 11243 12129
rect 11398 11316 11408 12129
rect 14692 12116 14702 12180
rect 14766 12116 14776 12180
rect 23681 12126 23691 12190
rect 23755 12126 23765 12190
rect 14682 11612 14692 11676
rect 14756 11612 14766 11676
rect 14692 11520 14756 11612
rect 23679 11455 23689 11519
rect 23753 11455 23763 11519
rect 11268 11311 11373 11316
rect 5662 10402 5714 11030
rect -5855 10349 -5845 10402
rect -5792 10350 -678 10402
rect -626 10350 5714 10402
rect 6484 10502 11218 10536
rect 6484 10409 6553 10502
rect 11090 10409 11218 10502
rect 6484 10357 11218 10409
rect -5792 10349 5714 10350
rect 14681 10319 14691 10383
rect 14755 10319 14765 10383
rect 23681 10316 23691 10380
rect 23755 10316 23765 10380
rect 362 10003 372 10144
rect 1812 10003 1822 10144
rect 5717 9990 5727 10135
rect 11722 9990 11732 10135
rect 13866 9993 13876 10150
rect 21118 9993 21128 10150
rect -6177 9513 -6167 9592
rect -5929 9513 -5919 9592
rect -5718 9509 -5708 9595
rect -5399 9509 -5389 9595
rect -1769 9532 -1759 9930
rect -1695 9532 -1685 9930
rect 3748 9911 5265 9945
rect -5855 9400 -5845 9452
rect -5793 9400 -5783 9452
rect -3924 9385 -3914 9437
rect -3862 9385 -3040 9437
rect -1726 9383 -1149 9435
rect -1097 9383 -1087 9435
rect -1779 9061 -1498 9125
rect -1434 9061 -1424 9125
rect -5863 8110 -5853 8174
rect -5789 8110 -5779 8174
rect -1768 7930 -1758 8330
rect -1690 7930 -1680 8330
rect -3425 7783 -3415 7835
rect -3363 7783 -3029 7835
rect -1726 7783 -1149 7835
rect -1097 7783 -1087 7835
rect -6572 7591 -5853 7595
rect -6575 7527 -6565 7591
rect -6501 7531 -5853 7591
rect -5789 7531 -5779 7595
rect -6501 7527 -6491 7531
rect -1796 7522 -1498 7586
rect -1434 7522 -1424 7586
rect -7224 7003 -7214 7243
rect -6751 7175 -6741 7243
rect -1508 7175 -1498 7258
rect -6751 7066 -1498 7175
rect -6751 7003 -6741 7066
rect -1508 6974 -1498 7066
rect -1434 6974 -1424 7258
rect -25531 6408 -25521 6669
rect -25446 6408 -25436 6669
rect -4927 6392 -4917 6695
rect -4836 6392 -4826 6695
rect -3114 6387 -1498 6451
rect -1434 6387 -1424 6451
rect -31140 6209 -31130 6337
rect -31002 6209 -26744 6337
rect -25374 6303 -18149 6336
rect -25603 6239 -18251 6303
rect -18187 6239 -18149 6303
rect -13085 6249 -13075 6313
rect -13011 6249 -6565 6313
rect -6501 6249 -6261 6313
rect -4806 6258 -3415 6310
rect -3363 6258 -3353 6310
rect -25374 6208 -18149 6239
rect -25532 5929 -25522 6174
rect -25447 5929 -25437 6174
rect -4917 5950 -4907 6163
rect -4841 5950 -4831 6163
rect -3114 6161 -3050 6387
rect -3425 5671 -3415 5723
rect -3363 5671 -2970 5723
rect -1832 5671 -678 5723
rect -626 5671 -616 5723
rect -3203 5296 -3193 5577
rect -3110 5296 -3069 5577
rect 19 5570 29 9830
rect 212 5570 222 9830
rect 5231 9418 5265 9911
rect 21277 9911 21389 9923
rect 5213 9365 5223 9418
rect 5276 9365 5286 9418
rect 4669 8188 4679 8366
rect 4857 8188 4867 8366
rect 17636 8273 17646 8451
rect 17824 8273 17834 8451
rect 21277 7514 21283 9911
rect 21383 7514 21389 9911
rect 24534 9360 24544 9424
rect 24608 9360 24618 9424
rect 23198 7792 23208 7845
rect 23261 7792 23271 7845
rect 4669 6188 4679 6366
rect 4857 6188 4867 6366
rect 13340 6313 13350 6491
rect 13528 6313 13538 6491
rect 17636 6273 17646 6451
rect 17824 6273 17834 6451
rect -1149 5129 899 5130
rect -1159 5077 -1149 5129
rect -1097 5077 899 5129
rect -3437 4983 -3427 5047
rect -3363 4983 -3353 5047
rect -3427 4973 -3363 4983
rect 16091 4910 16101 5088
rect 16279 4910 16289 5088
rect 19091 4910 19101 5088
rect 19279 4910 19289 5088
rect 21240 4540 21250 7514
rect 21417 4540 21427 7514
rect 23208 4916 23261 7792
rect 24544 6312 24608 9360
rect 35014 8219 35024 8283
rect 35088 8219 35098 8283
rect 38565 7892 38575 8038
rect 38645 7892 38655 8038
rect 40090 7933 40100 8121
rect 40181 7933 40191 8121
rect 36291 7814 36301 7881
rect 36532 7814 36542 7881
rect 33736 7587 33746 7651
rect 33810 7587 33820 7651
rect 38558 7375 38568 7563
rect 38649 7375 38659 7563
rect 40077 7388 40087 7576
rect 40168 7388 40178 7576
rect 36352 7275 36362 7337
rect 36531 7275 36541 7337
rect 35018 7159 35028 7223
rect 35092 7159 35102 7223
rect 42592 7143 42602 7232
rect 45923 7143 45933 7232
rect 35017 6890 35027 6954
rect 35091 6890 35101 6954
rect 36342 6721 36352 6795
rect 36437 6721 36447 6795
rect 38561 6582 38571 6707
rect 38649 6582 38659 6707
rect 40082 6597 40092 6785
rect 40173 6597 40183 6785
rect 24534 6248 24544 6312
rect 24608 6248 24618 6312
rect 33724 6248 33734 6312
rect 33798 6248 33808 6312
rect 35757 6169 36971 6265
rect 37067 6169 37077 6265
rect 38553 6044 38563 6232
rect 38644 6044 38654 6232
rect 40082 6041 40092 6229
rect 40173 6041 40183 6229
rect 35017 5821 35027 5885
rect 35091 5821 35101 5885
rect 47463 5744 47473 5800
rect 35960 5644 35970 5707
rect 36149 5644 36159 5707
rect 40356 5616 47473 5744
rect 47463 5564 47473 5616
rect 47709 5564 47719 5800
rect 35014 5498 35024 5562
rect 35088 5498 35098 5562
rect 38564 5187 38574 5322
rect 38648 5187 38658 5322
rect 40099 5217 40109 5405
rect 40190 5217 40200 5405
rect 36504 5092 36514 5162
rect 36734 5092 36744 5162
rect 23198 4863 23208 4916
rect 23261 4863 23271 4916
rect 33732 4863 33742 4916
rect 33795 4863 33805 4916
rect 38552 4691 38562 4879
rect 38643 4691 38653 4879
rect 40082 4669 40092 4857
rect 40173 4669 40183 4857
rect 36354 4555 36364 4613
rect 36509 4555 36519 4613
rect 4669 4188 4679 4366
rect 4857 4188 4867 4366
rect -253 3789 867 3790
rect -289 3737 -279 3789
rect -227 3737 867 3789
rect -2121 3298 3361 3416
rect -2121 3180 1661 3298
rect -2121 -6585 -1885 3180
rect 18 359 28 2773
rect 190 359 200 2773
rect 12197 2595 12207 2773
rect 12385 2595 12395 2773
rect 4669 2188 4679 2366
rect 4857 2188 4867 2366
rect 21277 2139 21283 4540
rect 21383 2139 21389 4540
rect 35025 4428 35035 4492
rect 35099 4428 35109 4492
rect 23422 2354 23432 2407
rect 23485 2354 23495 2407
rect 21233 1288 21243 2139
rect 21419 1288 21429 2139
rect 21277 493 21283 1288
rect 21383 493 21389 1288
rect 22579 1044 22589 1097
rect 22642 1044 22652 1097
rect 21277 481 21389 493
rect 312 67 322 232
rect 21107 67 21117 232
rect 22589 -2017 22642 1044
rect 23432 -640 23485 2354
rect 26001 716 26076 4397
rect 35014 4123 35024 4187
rect 35088 4123 35098 4187
rect 42589 4144 42599 4233
rect 45959 4144 45969 4233
rect 36299 3993 36972 4089
rect 37068 3993 37078 4089
rect 38562 3781 38572 3934
rect 38651 3781 38661 3934
rect 40089 3838 40099 4026
rect 40180 3838 40190 4026
rect 36349 3459 36359 3531
rect 36486 3459 36496 3531
rect 38555 3291 38565 3479
rect 38646 3291 38656 3479
rect 40079 3285 40089 3473
rect 40170 3285 40180 3473
rect 35021 3058 35031 3122
rect 35095 3058 35105 3122
rect 35014 1279 35024 1343
rect 35088 1279 35098 1343
rect 38565 952 38575 1098
rect 38645 952 38655 1098
rect 40090 993 40100 1181
rect 40181 993 40191 1181
rect 36291 874 36301 941
rect 36532 874 36542 941
rect 25991 641 26001 716
rect 26076 641 26086 716
rect 33720 641 33730 716
rect 33805 711 33815 716
rect 33810 647 33820 711
rect 33805 641 33815 647
rect 38558 435 38568 623
rect 38649 435 38659 623
rect 40077 448 40087 636
rect 40168 448 40178 636
rect 36352 335 36362 397
rect 36531 335 36541 397
rect 35018 219 35028 283
rect 35092 219 35102 283
rect 42589 199 42599 309
rect 45930 199 45940 309
rect 35017 -50 35027 14
rect 35091 -50 35101 14
rect 36342 -219 36352 -145
rect 36437 -219 36447 -145
rect 38561 -358 38571 -233
rect 38649 -358 38659 -233
rect 40082 -343 40092 -155
rect 40173 -343 40183 -155
rect 23422 -693 23432 -640
rect 23485 -693 23495 -640
rect 33724 -692 33734 -628
rect 33798 -692 33808 -628
rect 33731 -693 33741 -692
rect 33794 -693 33804 -692
rect 35757 -771 36971 -675
rect 37067 -771 37077 -675
rect 38553 -896 38563 -708
rect 38644 -896 38654 -708
rect 40082 -899 40092 -711
rect 40173 -899 40183 -711
rect 35017 -1119 35027 -1055
rect 35091 -1119 35101 -1055
rect 47479 -1196 47489 -1140
rect 35960 -1296 35970 -1233
rect 36149 -1296 36159 -1233
rect 40356 -1324 47489 -1196
rect 47479 -1376 47489 -1324
rect 47725 -1376 47735 -1140
rect 35014 -1442 35024 -1378
rect 35088 -1442 35098 -1378
rect 38564 -1753 38574 -1618
rect 38648 -1753 38658 -1618
rect 40099 -1723 40109 -1535
rect 40190 -1723 40200 -1535
rect 36504 -1848 36514 -1778
rect 36734 -1848 36744 -1778
rect 22579 -2070 22589 -2017
rect 22643 -2070 22653 -2017
rect 33747 -2024 33757 -2017
rect 22589 -2073 22642 -2070
rect 33732 -2077 33742 -2024
rect 33810 -2070 33820 -2017
rect 33795 -2077 33805 -2070
rect 38552 -2249 38562 -2061
rect 38643 -2249 38653 -2061
rect 40082 -2271 40092 -2083
rect 40173 -2271 40183 -2083
rect 36354 -2385 36364 -2327
rect 36509 -2385 36519 -2327
rect 35025 -2512 35035 -2448
rect 35099 -2512 35109 -2448
rect 35014 -2817 35024 -2753
rect 35088 -2817 35098 -2753
rect 42577 -2796 42587 -2708
rect 45933 -2796 45943 -2708
rect 36299 -2947 36972 -2851
rect 37068 -2947 37078 -2851
rect 38562 -3159 38572 -3006
rect 38651 -3159 38661 -3006
rect 40089 -3102 40099 -2914
rect 40180 -3102 40190 -2914
rect 36349 -3481 36359 -3409
rect 36486 -3481 36496 -3409
rect 38555 -3649 38565 -3461
rect 38646 -3649 38656 -3461
rect 40079 -3655 40089 -3467
rect 40170 -3655 40180 -3467
rect 35021 -3882 35031 -3818
rect 35095 -3882 35105 -3818
rect -2121 -6799 -1993 -6585
rect -3605 -10130 -3595 -6822
rect -3503 -10130 -3493 -6822
rect -2121 -10365 -2003 -6799
rect -610 -10140 -600 -6825
rect -486 -10140 -476 -6825
rect -2179 -12082 -1943 -10365
rect -2189 -12318 -2179 -12082
rect -1943 -12318 -1933 -12082
<< via1 >>
rect -15410 77904 -15174 78140
rect -16849 73398 -16748 76723
rect 12606 77875 12842 78111
rect 24656 77876 24892 78112
rect -13848 73404 -13747 76729
rect 11143 76698 11271 76732
rect 11143 73428 11189 76698
rect 11189 73428 11223 76698
rect 11223 73428 11271 76698
rect 11143 73392 11271 73428
rect 14144 73405 14272 76745
rect -16664 71738 -16600 71802
rect -15486 71734 -15422 71798
rect -15269 71741 -15205 71805
rect -14135 71738 -14071 71802
rect -16554 70234 -16490 70298
rect -15440 70220 -15376 70284
rect -15227 70221 -15163 70285
rect -14063 70221 -13999 70285
rect -15963 68105 -15890 68261
rect -15422 68166 -15358 68515
rect -14879 68108 -14806 68264
rect -16577 67549 -16513 67613
rect -15422 67543 -15358 67607
rect -14304 67554 -14240 67618
rect -9884 63338 -9442 63402
rect -8073 63340 -7631 63404
rect -6278 63336 -5836 63400
rect -6939 62966 -6699 63206
rect -4479 63334 -4037 63398
rect -2688 63338 -2246 63402
rect -886 63334 -444 63398
rect 757 62992 1287 63232
rect -8557 54531 -8493 54595
rect -6866 54532 -6802 54596
rect -9704 54339 -9462 54403
rect -5161 54531 -5097 54595
rect -3365 54531 -3301 54595
rect -1536 54531 -1472 54595
rect -7909 54338 -7667 54402
rect -6109 54340 -5867 54404
rect -4311 54339 -4069 54403
rect -2513 54340 -2271 54404
rect -710 54339 -468 54403
rect 176 54340 240 54404
rect -14783 53536 -14655 53600
rect -7550 53536 -7486 53600
rect -6989 53536 -6861 53600
rect 347 60758 519 60827
rect 347 53140 377 60758
rect 377 53140 477 60758
rect 477 53140 519 60758
rect 347 53121 519 53140
rect 5410 58752 5588 58930
rect 2047 57297 2225 57475
rect 4047 57297 4225 57475
rect 5410 55752 5588 55930
rect 4007 53001 4185 53179
rect -9398 52928 -9270 52992
rect 7725 51858 7903 52036
rect -8854 51014 -8770 51249
rect -9398 50873 -9270 50937
rect -6989 50871 -6861 50935
rect -5688 51018 -3888 51066
rect -3362 51018 -2536 51074
rect -1655 51018 -765 51064
rect -5688 50925 -5624 51018
rect -5624 50925 -3888 51018
rect -3362 50925 -2536 51018
rect -1655 50925 -765 51018
rect -5688 50883 -3888 50925
rect -3362 50896 -2536 50925
rect -1655 50886 -765 50925
rect -8874 50378 -8780 50791
rect -27070 49656 -26726 49720
rect -26408 49404 -26157 49413
rect -26408 49359 -26399 49404
rect -26399 49359 -26176 49404
rect -26176 49359 -26157 49404
rect -26408 49349 -26157 49359
rect -26060 49413 -26047 49424
rect -26047 49413 -26013 49424
rect -26013 49413 -25996 49424
rect -26060 49361 -25996 49413
rect -26060 49360 -26047 49361
rect -26047 49360 -26013 49361
rect -26013 49360 -25996 49361
rect -25984 49114 -25640 49178
rect -5932 47776 -5748 50720
rect -78 50741 121 50774
rect -78 47771 -4 50741
rect -4 47771 89 50741
rect 89 47771 121 50741
rect -78 47752 121 47771
rect 10177 47617 10551 60836
rect -27087 42779 -26990 43313
rect -13469 42997 -13405 43061
rect -27082 41002 -26995 42169
rect -27077 39476 -26990 40643
rect -31812 39132 -31748 39166
rect -31812 38846 -31795 39132
rect -31795 38846 -31761 39132
rect -31761 38846 -31748 39132
rect -31812 38827 -31748 38846
rect -31811 38576 -31747 38613
rect -31811 38202 -31795 38576
rect -31795 38202 -31761 38576
rect -31761 38202 -31747 38576
rect -31811 38141 -31747 38202
rect -29614 38349 -29150 38413
rect -31030 38192 -30901 38256
rect -27082 38232 -26998 39120
rect -35518 37332 -35282 37568
rect -30199 37411 -30070 37475
rect -29652 37259 -29143 37323
rect -27079 36465 -26995 37353
rect -27077 34985 -26996 36160
rect -18883 36124 -18807 39537
rect -27079 33498 -27000 34691
rect -27084 32365 -27005 32899
rect -12693 42334 -12629 42398
rect -5924 39819 -5722 46274
rect -4101 45129 -3923 45307
rect -1482 44281 -1304 44459
rect -9398 39741 -9270 39805
rect -6989 39741 -6861 39805
rect -9369 34612 -9305 34676
rect -5684 39803 -148 39846
rect -5684 39710 -5637 39803
rect -5637 39710 -168 39803
rect -168 39710 -148 39803
rect -5684 39666 -148 39710
rect 344 45818 558 45844
rect 344 44350 377 45818
rect 377 44350 477 45818
rect 477 44350 558 45818
rect 344 44318 558 44350
rect 2132 44330 2310 44508
rect 4132 44330 4310 44508
rect 6132 44330 6310 44508
rect 8132 44330 8310 44508
rect 352 41343 512 41383
rect 352 40051 377 41343
rect 377 40051 477 41343
rect 477 40051 512 41343
rect 352 39855 512 40051
rect 2513 38642 2595 38881
rect 93 38502 157 38566
rect 1230 38502 1294 38566
rect 2626 38504 2690 38568
rect 5361 38504 5425 38568
rect 2515 37996 2614 38420
rect 5361 38091 5425 38155
rect 93 37587 157 37651
rect 3427 37587 3491 37651
rect 2168 36898 2232 37149
rect 2644 37143 2708 37207
rect 93 36752 157 36816
rect 883 36752 947 36816
rect 2169 36250 2233 36668
rect 2938 36030 3343 36088
rect 10180 39867 10551 46128
rect 17430 64169 17496 64743
rect 23958 64169 24024 64743
rect 31574 64169 31640 64743
rect 17975 62166 18041 62740
rect 19063 62166 19129 62740
rect 21239 62166 21305 62740
rect 22327 62166 22393 62740
rect 23415 62166 23481 62740
rect 24503 62166 24569 62740
rect 25591 62166 25657 62740
rect 26679 62166 26745 62740
rect 28855 62166 28921 62740
rect 29943 62166 30009 62740
rect 31031 62166 31097 62740
rect 17430 60169 17496 60743
rect 18518 60169 18584 60743
rect 19606 60169 19672 60743
rect 20694 60169 20760 60743
rect 21782 60169 21848 60743
rect 22870 60169 22936 60743
rect 23958 60169 24024 60743
rect 25046 60169 25112 60743
rect 26134 60169 26200 60743
rect 27222 60169 27288 60743
rect 28310 60169 28376 60743
rect 29398 60169 29464 60743
rect 30486 60169 30552 60743
rect 31574 60169 31640 60743
rect 17975 58166 18041 58740
rect 19063 58166 19129 58740
rect 20151 58166 20217 58740
rect 21239 58166 21305 58740
rect 22327 58166 22393 58740
rect 23415 58166 23481 58740
rect 24503 58166 24569 58740
rect 25591 58166 25657 58740
rect 26679 58166 26745 58740
rect 27767 58166 27833 58740
rect 28855 58166 28921 58740
rect 29943 58166 30009 58740
rect 31031 58166 31097 58740
rect 17430 56169 17496 56743
rect 18518 56169 18584 56743
rect 19606 56169 19672 56743
rect 20694 56169 20760 56743
rect 21782 56169 21848 56743
rect 22870 56169 22936 56743
rect 23958 56169 24024 56743
rect 25046 56169 25112 56743
rect 26134 56169 26200 56743
rect 27222 56169 27288 56743
rect 28310 56169 28376 56743
rect 29398 56169 29464 56743
rect 30486 56169 30552 56743
rect 31574 56169 31640 56743
rect 17975 54166 18041 54740
rect 19063 54166 19129 54740
rect 20151 54166 20217 54740
rect 21239 54166 21305 54740
rect 22327 54166 22393 54740
rect 23415 54166 23481 54740
rect 24503 54166 24569 54740
rect 25591 54166 25657 54740
rect 26679 54166 26745 54740
rect 27767 54166 27833 54740
rect 28855 54166 28921 54740
rect 29943 54166 30009 54740
rect 31031 54166 31097 54740
rect 17430 52169 17496 52743
rect 18518 52169 18584 52743
rect 19606 52169 19672 52743
rect 20694 52169 20760 52743
rect 21782 52169 21848 52743
rect 22870 52169 22936 52743
rect 23958 52169 24024 52743
rect 25046 52169 25112 52743
rect 26134 52169 26200 52743
rect 27222 52169 27288 52743
rect 28310 52169 28376 52743
rect 29398 52169 29464 52743
rect 30486 52169 30552 52743
rect 31574 52169 31640 52743
rect 17975 50166 18041 50740
rect 20151 50166 20217 50740
rect 21239 50166 21305 50740
rect 23415 50166 23481 50740
rect 24503 50166 24569 50740
rect 25591 50166 25657 50740
rect 27767 50166 27833 50740
rect 28855 50166 28921 50740
rect 31031 50166 31097 50740
rect 17430 48169 17496 48743
rect 18518 48169 18584 48743
rect 19606 48169 19672 48743
rect 20694 48169 20760 48743
rect 21782 48169 21848 48743
rect 22870 48169 22936 48743
rect 23958 48169 24024 48743
rect 29398 48169 29464 48743
rect 30486 48169 30552 48743
rect 31574 48169 31640 48743
rect 17975 46166 18041 46740
rect 19063 46166 19129 46740
rect 20151 46166 20217 46740
rect 21239 46166 21305 46740
rect 22327 46166 22393 46740
rect 24503 46166 24569 46740
rect 25591 46166 25657 46740
rect 26679 46166 26745 46740
rect 27767 46166 27833 46740
rect 28855 46166 28921 46740
rect 29943 46166 30009 46740
rect 31031 46166 31097 46740
rect 18245 45684 18309 45748
rect 18791 45684 18855 45748
rect 19337 45675 19401 45739
rect 19882 45674 19946 45738
rect 21517 45684 21581 45748
rect 22051 45671 22115 45735
rect 22598 45677 22662 45741
rect 23143 45677 23207 45741
rect 25863 45674 25927 45738
rect 26406 45678 26470 45742
rect 26948 45672 27012 45736
rect 27505 45663 27569 45727
rect 29129 45674 29193 45738
rect 29673 45667 29737 45731
rect 30223 45671 30287 45735
rect 30756 45671 30820 45735
rect 44754 45007 45306 45074
rect 39557 44827 39621 44891
rect 40595 44816 40647 44830
rect 40595 44782 40603 44816
rect 40603 44782 40637 44816
rect 40637 44782 40647 44816
rect 40595 44778 40647 44782
rect 40995 44810 41047 44819
rect 40995 44776 41005 44810
rect 41005 44776 41039 44810
rect 41039 44776 41047 44810
rect 40995 44767 41047 44776
rect 41152 44816 41204 44823
rect 41152 44782 41161 44816
rect 41161 44782 41195 44816
rect 41195 44782 41204 44816
rect 41152 44771 41204 44782
rect 40894 44751 40946 44762
rect 40894 44717 40905 44751
rect 40905 44717 40939 44751
rect 40939 44717 40946 44751
rect 40894 44710 40946 44717
rect 39557 44637 39621 44701
rect 46294 44703 46530 44939
rect 41516 44462 41874 44527
rect 44766 43854 45293 43925
rect 39557 43677 39621 43741
rect 40595 43666 40647 43680
rect 40595 43632 40603 43666
rect 40603 43632 40637 43666
rect 40637 43632 40647 43666
rect 40595 43628 40647 43632
rect 40995 43660 41047 43669
rect 40995 43626 41005 43660
rect 41005 43626 41039 43660
rect 41039 43626 41047 43660
rect 40995 43617 41047 43626
rect 41152 43666 41204 43673
rect 41152 43632 41161 43666
rect 41161 43632 41195 43666
rect 41195 43632 41204 43666
rect 41152 43621 41204 43632
rect 40894 43601 40946 43612
rect 40894 43567 40905 43601
rect 40905 43567 40939 43601
rect 40939 43567 40946 43601
rect 40894 43560 40946 43567
rect 39557 43487 39621 43551
rect 46282 43552 46518 43788
rect 41514 43312 41872 43377
rect 44756 41312 45283 41383
rect 39557 41137 39621 41201
rect 40595 41126 40647 41140
rect 40595 41092 40603 41126
rect 40603 41092 40637 41126
rect 40637 41092 40647 41126
rect 40595 41088 40647 41092
rect 40995 41120 41047 41129
rect 40995 41086 41005 41120
rect 41005 41086 41039 41120
rect 41039 41086 41047 41120
rect 40995 41077 41047 41086
rect 41152 41126 41204 41133
rect 41152 41092 41161 41126
rect 41161 41092 41195 41126
rect 41195 41092 41204 41126
rect 41152 41081 41204 41092
rect 40894 41061 40946 41072
rect 40894 41027 40905 41061
rect 40905 41027 40939 41061
rect 40939 41027 40946 41061
rect 40894 41020 40946 41027
rect 39557 40947 39621 41011
rect 46140 41020 46376 41256
rect 41432 40771 41790 40836
rect 44756 40042 45283 40113
rect 39557 39867 39621 39931
rect 40595 39856 40647 39870
rect 40595 39822 40603 39856
rect 40603 39822 40637 39856
rect 40637 39822 40647 39856
rect 40595 39818 40647 39822
rect 40995 39850 41047 39859
rect 40995 39816 41005 39850
rect 41005 39816 41039 39850
rect 41039 39816 41047 39850
rect 40995 39807 41047 39816
rect 41152 39856 41204 39863
rect 41152 39822 41161 39856
rect 41161 39822 41195 39856
rect 41195 39822 41204 39856
rect 41152 39811 41204 39822
rect 40894 39791 40946 39802
rect 40894 39757 40905 39791
rect 40905 39757 40939 39791
rect 40939 39757 40946 39791
rect 40894 39750 40946 39757
rect 39557 39677 39621 39741
rect 46111 39730 46347 39966
rect 41430 39502 41788 39567
rect 7082 38974 7318 39210
rect 12542 38974 12778 39210
rect 7236 38091 7300 38155
rect 5429 37143 5493 37207
rect 6701 37143 6765 37207
rect 3582 36030 3811 36094
rect 5055 36018 5351 36104
rect 9428 37587 9492 37651
rect 5574 36027 5801 36097
rect 6936 36020 7157 36089
rect 7383 36028 7681 36094
rect 8921 36028 9348 36093
rect 9575 36023 9802 36091
rect 5430 34956 5494 35020
rect 7242 34954 7306 35018
rect 3745 33798 3797 33850
rect -6948 33115 -6884 33179
rect -6989 31747 -6861 31811
rect 5430 34361 5494 34425
rect 7242 34361 7306 34425
rect 5430 33497 5494 33561
rect 7428 33505 7492 33569
rect 9745 33798 9797 33850
rect 4354 30368 4418 30432
rect 8328 30373 8392 30437
rect -9397 30241 -9269 30305
rect -12693 29688 -12629 29752
rect -30199 29159 -30070 29288
rect -18523 29159 -18394 29288
rect -13469 29265 -13405 29329
rect 1951 28744 2079 28808
rect 7960 28782 8024 28846
rect -6086 28544 -5958 28608
rect 3399 28531 3463 28595
rect -31030 27801 -30901 27930
rect -19383 27801 -19254 27930
rect -15712 27645 -15613 28098
rect -13983 28014 -13931 28066
rect -12389 27670 -12316 28076
rect -18326 27511 -18262 27575
rect -17635 27516 -17507 27644
rect -14906 27519 -14854 27571
rect -14404 27207 -14352 27259
rect -12394 27198 -12297 27427
rect -18326 27034 -18262 27098
rect -18881 26696 -18817 26760
rect -38190 26514 -34856 26611
rect -18882 25913 -18818 25977
rect -25449 25175 -25369 25482
rect -40593 24935 -40357 25171
rect -32991 24984 -32863 25112
rect -25452 24714 -25365 24945
rect -38182 23503 -34852 23605
rect -18881 24392 -18817 24456
rect -14906 27031 -14854 27083
rect -17256 26696 -17192 26760
rect -10016 26524 -9888 26588
rect -17635 26287 -17507 26415
rect -13983 26414 -13931 26466
rect -15725 26044 -15636 26281
rect -12396 26057 -12301 26486
rect -14906 25915 -14854 25967
rect -14404 25607 -14352 25659
rect -12384 25604 -12321 25823
rect 1952 25756 2080 25820
rect -15727 25018 -15632 25447
rect -3501 25350 -3373 25414
rect -17635 24874 -17507 25002
rect -13983 24814 -13931 24866
rect -12393 24458 -12328 24712
rect -14908 24389 -14856 24441
rect -18326 24053 -18262 24117
rect -17255 24053 -17191 24117
rect -14404 24007 -14352 24059
rect -12398 24003 -12316 24239
rect 9399 28528 9463 28592
rect 7960 25756 8024 25820
rect 5715 24186 5783 24594
rect 3399 24037 3463 24101
rect -17635 23645 -17507 23773
rect -15725 23405 -15658 23637
rect 5643 24033 5707 24097
rect 7017 24037 7081 24101
rect 9399 24037 9463 24101
rect 42856 24065 46190 24174
rect 35152 23802 35216 23866
rect 37819 23492 37892 23611
rect 39346 23493 39420 23714
rect -13983 23214 -13931 23266
rect -12389 22857 -12319 23277
rect 8787 23246 8943 23356
rect 2550 22999 2614 23063
rect 10202 22999 10266 23063
rect -14908 22719 -14856 22771
rect -11601 22712 -11473 22776
rect -14404 22407 -14352 22459
rect -12391 22399 -12323 22624
rect -6086 21607 -5958 21671
rect -3501 20745 -3373 20809
rect -38168 18987 -34861 19065
rect -40596 17394 -40360 17630
rect -25452 17627 -25387 17922
rect -31130 17454 -31002 17582
rect -444 19981 -380 20109
rect 1684 19282 1748 19410
rect 233 17708 297 17772
rect -821 17461 -757 17525
rect -25450 17169 -25378 17404
rect 4397 21985 4449 22037
rect 8228 21985 8280 22037
rect 4397 20893 4449 20945
rect 8228 20893 8280 20945
rect 5394 19981 5458 20109
rect 9394 19981 9458 20109
rect 3395 19282 3459 19346
rect 3061 19042 3125 19106
rect 4857 19027 5194 19173
rect 7394 19282 7458 19410
rect 7085 19042 7149 19106
rect -445 17093 -381 17221
rect 1684 17093 1748 17221
rect 4295 17225 4359 17289
rect 8981 19042 9045 19106
rect 37819 22946 37905 23194
rect 39335 22952 39421 23200
rect 35100 22610 35280 22790
rect 35760 22668 36021 22730
rect 37826 22151 37896 22280
rect 39346 22167 39420 22388
rect 13887 21996 13951 22124
rect 47556 22498 47792 22734
rect 37814 21621 37899 21823
rect 39341 21586 39427 21834
rect 35152 21521 35216 21585
rect 42854 21069 46188 21178
rect 14688 20963 14752 21027
rect 23670 20152 23734 20216
rect 23689 19318 23753 19382
rect 14686 19214 14750 19278
rect 10232 18994 10296 19058
rect 8280 18654 8344 18718
rect 13574 18624 13638 18688
rect 23658 18364 23722 18428
rect 13887 17983 13951 18047
rect 14689 17485 14753 17549
rect 23689 17488 23753 17552
rect 6227 17225 6291 17289
rect 7393 17231 7457 17359
rect 9396 17231 9460 17359
rect 13885 17231 13949 17359
rect 14690 17019 14754 17083
rect 3393 16738 3457 16866
rect 5393 16738 5457 16866
rect 13277 16738 13341 16866
rect -3926 16224 -3862 16288
rect 251 16238 11139 16446
rect -38174 15987 -34852 16075
rect -5786 15644 -5722 15708
rect -3914 15083 -3862 15135
rect -678 15084 -626 15136
rect -3144 14719 -3061 14998
rect -25517 14157 -25444 14446
rect -4902 14236 -4832 14446
rect -32991 13974 -32863 14102
rect -13064 14077 -13000 14141
rect -6544 14077 -6480 14141
rect -3914 14087 -3862 14139
rect -18223 14009 -18159 14073
rect -25518 13690 -25446 13925
rect -4917 13706 -4833 13998
rect -6544 12828 -6480 12892
rect -5851 12828 -5787 12892
rect -1808 12726 -1725 13133
rect -3914 12583 -3862 12635
rect -279 12585 -227 12637
rect -1498 12345 -1434 12409
rect -5851 12155 -5787 12219
rect -1759 11140 -1693 11529
rect -3415 10982 -3363 11034
rect -279 10983 -227 11035
rect -5845 10891 -5793 10943
rect -6162 10758 -5937 10833
rect -5707 10751 -5401 10838
rect -1498 10719 -1434 10783
rect 28 16135 187 16189
rect 28 10666 59 16135
rect 59 10666 152 16135
rect 152 10666 187 16135
rect 28 10640 187 10666
rect 5478 14421 5656 14599
rect 11239 16122 11399 16184
rect 11239 14432 11274 16122
rect 11274 14432 11367 16122
rect 11367 14432 11399 16122
rect 11239 14426 11399 14432
rect 14685 15689 14749 15753
rect 23686 15724 23750 15788
rect 20928 15432 20992 15496
rect 14690 15164 14754 15228
rect 11257 13953 11384 13954
rect 11257 12990 11274 13953
rect 11274 12990 11367 13953
rect 11367 12990 11384 13953
rect 14685 13901 14749 13965
rect 23686 13933 23750 13997
rect 14690 13464 14754 13528
rect 23685 12942 23749 13006
rect 4630 11802 4808 11980
rect 11243 12105 11398 12129
rect 11243 11323 11274 12105
rect 11274 11323 11367 12105
rect 11367 11323 11398 12105
rect 11243 11316 11398 11323
rect 14702 12116 14766 12180
rect 23691 12126 23755 12190
rect 14692 11612 14756 11676
rect 23689 11455 23753 11519
rect -5845 10349 -5792 10402
rect -678 10350 -626 10402
rect 14691 10319 14755 10383
rect 23691 10316 23755 10380
rect 372 10121 1812 10144
rect 372 10021 400 10121
rect 400 10021 1790 10121
rect 1790 10021 1812 10121
rect 372 10003 1812 10021
rect 5727 10121 11722 10135
rect 5727 10021 5748 10121
rect 5748 10021 11698 10121
rect 11698 10021 11722 10121
rect 5727 9990 11722 10021
rect 13876 10121 21118 10150
rect 13876 10021 13915 10121
rect 13915 10021 21107 10121
rect 21107 10021 21118 10121
rect 13876 9993 21118 10021
rect -6167 9513 -5929 9592
rect -5708 9509 -5399 9595
rect -1759 9532 -1695 9930
rect -5845 9400 -5793 9452
rect -3914 9385 -3862 9437
rect -1149 9383 -1097 9435
rect -1498 9061 -1434 9125
rect -5853 8110 -5789 8174
rect -1758 7930 -1690 8330
rect -3415 7783 -3363 7835
rect -1149 7783 -1097 7835
rect -6565 7527 -6501 7591
rect -5853 7531 -5789 7595
rect -1498 7522 -1434 7586
rect -7214 7003 -6751 7243
rect -1498 6974 -1434 7258
rect -25521 6408 -25446 6669
rect -4917 6392 -4836 6695
rect -1498 6387 -1434 6451
rect -31130 6209 -31002 6337
rect -18251 6239 -18187 6303
rect -13075 6249 -13011 6313
rect -6565 6249 -6501 6313
rect -3415 6258 -3363 6310
rect -25522 5929 -25447 6174
rect -4907 5950 -4841 6163
rect -3415 5671 -3363 5723
rect -678 5671 -626 5723
rect -3193 5296 -3110 5577
rect 29 9792 212 9830
rect 29 5602 59 9792
rect 59 5602 159 9792
rect 159 5602 212 9792
rect 29 5570 212 5602
rect 5223 9365 5276 9418
rect 4679 8188 4857 8366
rect 17646 8273 17824 8451
rect 24544 9360 24608 9424
rect 23208 7792 23261 7845
rect 4679 6188 4857 6366
rect 13350 6313 13528 6491
rect 17646 6273 17824 6451
rect -1149 5077 -1097 5129
rect -3427 4983 -3363 5047
rect 16101 4910 16279 5088
rect 19101 4910 19279 5088
rect 21250 4540 21283 7514
rect 21283 4540 21383 7514
rect 21383 4540 21417 7514
rect 35024 8219 35088 8283
rect 38575 7892 38645 8038
rect 40100 7933 40181 8121
rect 36301 7814 36532 7881
rect 33746 7587 33810 7651
rect 38568 7375 38649 7563
rect 40087 7388 40168 7576
rect 36362 7275 36531 7337
rect 35028 7159 35092 7223
rect 42602 7143 45923 7232
rect 35027 6890 35091 6954
rect 36352 6721 36437 6795
rect 38571 6582 38649 6707
rect 40092 6597 40173 6785
rect 24544 6248 24608 6312
rect 33734 6248 33798 6312
rect 36971 6169 37067 6265
rect 38563 6044 38644 6232
rect 40092 6041 40173 6229
rect 35027 5821 35091 5885
rect 35970 5644 36149 5707
rect 47473 5564 47709 5800
rect 35024 5498 35088 5562
rect 38574 5187 38648 5322
rect 40109 5217 40190 5405
rect 36514 5092 36734 5162
rect 23208 4863 23261 4916
rect 33742 4863 33795 4916
rect 38562 4691 38643 4879
rect 40092 4669 40173 4857
rect 36364 4555 36509 4613
rect 4679 4188 4857 4366
rect -279 3737 -227 3789
rect 28 2748 190 2773
rect 28 374 59 2748
rect 59 374 159 2748
rect 159 374 190 2748
rect 28 359 190 374
rect 12207 2595 12385 2773
rect 4679 2188 4857 2366
rect 35035 4428 35099 4492
rect 23432 2354 23485 2407
rect 21243 1288 21283 2139
rect 21283 1288 21383 2139
rect 21383 1288 21419 2139
rect 22589 1044 22642 1097
rect 322 67 21107 232
rect 35024 4123 35088 4187
rect 42599 4144 45959 4233
rect 36972 3993 37068 4089
rect 38572 3781 38651 3934
rect 40099 3838 40180 4026
rect 36359 3459 36486 3531
rect 38565 3291 38646 3479
rect 40089 3285 40170 3473
rect 35031 3058 35095 3122
rect 35024 1279 35088 1343
rect 38575 952 38645 1098
rect 40100 993 40181 1181
rect 36301 874 36532 941
rect 26001 641 26076 716
rect 33730 711 33805 716
rect 33730 647 33810 711
rect 33730 641 33805 647
rect 38568 435 38649 623
rect 40087 448 40168 636
rect 36362 335 36531 397
rect 35028 219 35092 283
rect 42599 199 45930 309
rect 35027 -50 35091 14
rect 36352 -219 36437 -145
rect 38571 -358 38649 -233
rect 40092 -343 40173 -155
rect 23432 -693 23485 -640
rect 33734 -692 33798 -628
rect 33741 -693 33794 -692
rect 36971 -771 37067 -675
rect 38563 -896 38644 -708
rect 40092 -899 40173 -711
rect 35027 -1119 35091 -1055
rect 35970 -1296 36149 -1233
rect 47489 -1376 47725 -1140
rect 35024 -1442 35088 -1378
rect 38574 -1753 38648 -1618
rect 40109 -1723 40190 -1535
rect 36514 -1848 36734 -1778
rect 22589 -2070 22643 -2017
rect 33757 -2024 33810 -2017
rect 33742 -2070 33810 -2024
rect 33742 -2077 33795 -2070
rect 38562 -2249 38643 -2061
rect 40092 -2271 40173 -2083
rect 36364 -2385 36509 -2327
rect 35035 -2512 35099 -2448
rect 35024 -2817 35088 -2753
rect 42587 -2796 45933 -2708
rect 36972 -2947 37068 -2851
rect 38572 -3159 38651 -3006
rect 40099 -3102 40180 -2914
rect 36359 -3481 36486 -3409
rect 38565 -3649 38646 -3461
rect 40089 -3655 40170 -3467
rect 35031 -3882 35095 -3818
rect -3595 -10130 -3503 -6822
rect -600 -10140 -486 -6825
rect -2179 -12318 -1943 -12082
<< metal2 >>
rect -15410 78140 -15174 78150
rect -15410 77894 -15174 77904
rect 12606 78111 12842 78121
rect 12606 77865 12842 77875
rect 24656 78112 24892 78122
rect 24656 77866 24892 77876
rect 14144 76745 14272 76755
rect -16849 76723 -16748 76733
rect -16849 73388 -16748 73398
rect -13848 76729 -13747 76739
rect -13848 73394 -13747 73404
rect 11143 76732 11271 76742
rect 14144 73395 14272 73405
rect 11143 73382 11271 73392
rect -16664 71802 -16600 71812
rect -16664 71728 -16600 71738
rect -15486 71798 -15422 71808
rect -15486 71724 -15422 71734
rect -15269 71805 -15205 71815
rect -15269 71731 -15205 71741
rect -14135 71802 -14071 71812
rect -14135 71728 -14071 71738
rect -16554 70298 -16490 70308
rect -16554 70224 -16490 70234
rect -15440 70284 -15376 70294
rect -15440 70210 -15376 70220
rect -15227 70285 -15163 70295
rect -15227 70211 -15163 70221
rect -14063 70285 -13999 70295
rect -14063 70211 -13999 70221
rect -16708 68703 -16644 68713
rect -16708 68629 -16644 68639
rect -16699 68335 -16647 68629
rect -15422 68515 -15358 68525
rect -15963 68261 -15890 68271
rect -15422 68156 -15358 68166
rect -14879 68264 -14806 68274
rect -15963 68095 -15890 68105
rect -14879 68098 -14806 68108
rect -14192 68083 -14140 68387
rect -14199 68073 -14135 68083
rect -14199 67999 -14135 68009
rect -14192 67996 -14140 67999
rect -16577 67613 -16513 67623
rect -14304 67618 -14240 67628
rect -16577 67539 -16513 67549
rect -15422 67607 -15358 67617
rect -14304 67544 -14240 67554
rect -15422 67533 -15358 67543
rect 17430 64743 17496 64753
rect 17430 64159 17496 64169
rect 23958 64743 24024 64753
rect 23958 64159 24024 64169
rect 31574 64743 31640 64753
rect 31574 64159 31640 64169
rect -9884 63402 -9442 63412
rect -9884 63328 -9442 63338
rect -8073 63404 -7631 63414
rect -8073 63330 -7631 63340
rect -6278 63400 -5836 63410
rect -6278 63326 -5836 63336
rect -4479 63398 -4037 63408
rect -4479 63324 -4037 63334
rect -2688 63402 -2246 63412
rect -2688 63328 -2246 63338
rect -886 63398 -444 63408
rect -886 63324 -444 63334
rect 757 63232 1287 63242
rect -6939 63206 -6699 63216
rect 757 62982 1287 62992
rect -6939 62956 -6699 62966
rect 17975 62740 18041 62750
rect 17975 62156 18041 62166
rect 19063 62740 19129 62750
rect 19063 62156 19129 62166
rect 21239 62740 21305 62750
rect 21239 62156 21305 62166
rect 22327 62740 22393 62750
rect 22327 62156 22393 62166
rect 23415 62740 23481 62750
rect 23415 62156 23481 62166
rect 24503 62740 24569 62750
rect 24503 62156 24569 62166
rect 25591 62740 25657 62750
rect 25591 62156 25657 62166
rect 26679 62740 26745 62750
rect 26679 62156 26745 62166
rect 28855 62740 28921 62750
rect 28855 62156 28921 62166
rect 29943 62740 30009 62750
rect 29943 62156 30009 62166
rect 31031 62740 31097 62750
rect 31031 62156 31097 62166
rect 347 60827 519 60837
rect -8557 54595 -8493 54605
rect -8557 54521 -8493 54531
rect -6866 54596 -6802 54606
rect -6866 54522 -6802 54532
rect -5161 54595 -5097 54605
rect -5161 54521 -5097 54531
rect -3365 54595 -3301 54605
rect -3365 54521 -3301 54531
rect -1536 54595 -1472 54605
rect -1536 54521 -1472 54531
rect -9704 54403 -9462 54413
rect -9704 54329 -9462 54339
rect -7909 54402 -7667 54412
rect -7909 54328 -7667 54338
rect -6109 54404 -5867 54414
rect -6109 54330 -5867 54340
rect -4311 54403 -4069 54413
rect -4311 54329 -4069 54339
rect -2513 54404 -2271 54414
rect -2513 54330 -2271 54340
rect -710 54403 -468 54413
rect -710 54329 -468 54339
rect 176 54404 240 54414
rect 176 54330 240 54340
rect -14783 53600 -14655 53610
rect -7550 53600 -7486 53610
rect -14655 53536 -7550 53600
rect -14783 53526 -14655 53536
rect -7550 53526 -7486 53536
rect -6989 53600 -6861 53610
rect -9398 52992 -9270 53002
rect -9398 50937 -9270 52928
rect -8854 51249 -8770 51259
rect -7722 51247 -7658 51257
rect -7722 51173 -7658 51183
rect -8854 51004 -8770 51014
rect -27070 49720 -26726 49730
rect -27070 49646 -26726 49656
rect -26060 49424 -25996 49434
rect -26408 49413 -26157 49423
rect -26060 49350 -25996 49360
rect -26408 49339 -26157 49349
rect -25984 49178 -25640 49188
rect -25984 49104 -25640 49114
rect -27087 43313 -26990 43323
rect -13469 43061 -13405 43071
rect -13469 42987 -13405 42997
rect -27087 42769 -26990 42779
rect -12693 42398 -12629 42408
rect -12693 42324 -12629 42334
rect -27082 42169 -26995 42179
rect -21475 42163 -21411 42173
rect -21475 42089 -21411 42099
rect -27082 40992 -26995 41002
rect -27077 40643 -26990 40653
rect -9398 39805 -9270 50873
rect -6989 50935 -6861 53536
rect 10177 60836 10551 60846
rect 5410 58930 5588 58940
rect 5410 58742 5588 58752
rect 2047 57475 2225 57485
rect 2047 57287 2225 57297
rect 4047 57475 4225 57485
rect 4047 57287 4225 57297
rect 5410 55930 5588 55940
rect 5410 55742 5588 55752
rect 347 53111 519 53121
rect 4007 53179 4185 53189
rect 4007 52991 4185 53001
rect 7725 52036 7903 52046
rect 7725 51848 7903 51858
rect -5688 51066 -3888 51076
rect -3362 51074 -2536 51084
rect -3362 50886 -2536 50896
rect -1655 51064 -765 51074
rect -5688 50873 -3888 50883
rect -1655 50876 -765 50886
rect -8874 50791 -8780 50801
rect -8874 50368 -8780 50378
rect -8480 50441 -8416 50451
rect -8480 50367 -8416 50377
rect -9398 39728 -9270 39741
rect -6989 39805 -6861 50871
rect -78 50774 121 50784
rect -5932 50720 -5748 50730
rect -5932 47766 -5748 47776
rect -78 47742 121 47752
rect 17430 60743 17496 60753
rect 17430 60159 17496 60169
rect 18518 60743 18584 60753
rect 18518 60159 18584 60169
rect 19606 60743 19672 60753
rect 19606 60159 19672 60169
rect 20694 60743 20760 60753
rect 20694 60159 20760 60169
rect 21782 60743 21848 60753
rect 21782 60159 21848 60169
rect 22870 60743 22936 60753
rect 22870 60159 22936 60169
rect 23958 60743 24024 60753
rect 23958 60159 24024 60169
rect 25046 60743 25112 60753
rect 25046 60159 25112 60169
rect 26134 60743 26200 60753
rect 26134 60159 26200 60169
rect 27222 60743 27288 60753
rect 27222 60159 27288 60169
rect 28310 60743 28376 60753
rect 28310 60159 28376 60169
rect 29398 60743 29464 60753
rect 29398 60159 29464 60169
rect 30486 60743 30552 60753
rect 30486 60159 30552 60169
rect 31574 60743 31640 60753
rect 31574 60159 31640 60169
rect 17975 58740 18041 58750
rect 17975 58156 18041 58166
rect 19063 58740 19129 58750
rect 19063 58156 19129 58166
rect 20151 58740 20217 58750
rect 20151 58156 20217 58166
rect 21239 58740 21305 58750
rect 21239 58156 21305 58166
rect 22327 58740 22393 58750
rect 22327 58156 22393 58166
rect 23415 58740 23481 58750
rect 23415 58156 23481 58166
rect 24503 58740 24569 58750
rect 24503 58156 24569 58166
rect 25591 58740 25657 58750
rect 25591 58156 25657 58166
rect 26679 58740 26745 58750
rect 26679 58156 26745 58166
rect 27767 58740 27833 58750
rect 27767 58156 27833 58166
rect 28855 58740 28921 58750
rect 28855 58156 28921 58166
rect 29943 58740 30009 58750
rect 29943 58156 30009 58166
rect 31031 58740 31097 58750
rect 31031 58156 31097 58166
rect 17430 56743 17496 56753
rect 17430 56159 17496 56169
rect 18518 56743 18584 56753
rect 18518 56159 18584 56169
rect 19606 56743 19672 56753
rect 19606 56159 19672 56169
rect 20694 56743 20760 56753
rect 20694 56159 20760 56169
rect 21782 56743 21848 56753
rect 21782 56159 21848 56169
rect 22870 56743 22936 56753
rect 22870 56159 22936 56169
rect 23958 56743 24024 56753
rect 23958 56159 24024 56169
rect 25046 56743 25112 56753
rect 25046 56159 25112 56169
rect 26134 56743 26200 56753
rect 26134 56159 26200 56169
rect 27222 56743 27288 56753
rect 27222 56159 27288 56169
rect 28310 56743 28376 56753
rect 28310 56159 28376 56169
rect 29398 56743 29464 56753
rect 29398 56159 29464 56169
rect 30486 56743 30552 56753
rect 30486 56159 30552 56169
rect 31574 56743 31640 56753
rect 31574 56159 31640 56169
rect 17975 54740 18041 54750
rect 17975 54156 18041 54166
rect 19063 54740 19129 54750
rect 19063 54156 19129 54166
rect 20151 54740 20217 54750
rect 20151 54156 20217 54166
rect 21239 54740 21305 54750
rect 21239 54156 21305 54166
rect 22327 54740 22393 54750
rect 22327 54156 22393 54166
rect 23415 54740 23481 54750
rect 23415 54156 23481 54166
rect 24503 54740 24569 54750
rect 24503 54156 24569 54166
rect 25591 54740 25657 54750
rect 25591 54156 25657 54166
rect 26679 54740 26745 54750
rect 26679 54156 26745 54166
rect 27767 54740 27833 54750
rect 27767 54156 27833 54166
rect 28855 54740 28921 54750
rect 28855 54156 28921 54166
rect 29943 54740 30009 54750
rect 29943 54156 30009 54166
rect 31031 54740 31097 54750
rect 31031 54156 31097 54166
rect 17430 52743 17496 52753
rect 17430 52159 17496 52169
rect 18518 52743 18584 52753
rect 18518 52159 18584 52169
rect 19606 52743 19672 52753
rect 19606 52159 19672 52169
rect 20694 52743 20760 52753
rect 20694 52159 20760 52169
rect 21782 52743 21848 52753
rect 21782 52159 21848 52169
rect 22870 52743 22936 52753
rect 22870 52159 22936 52169
rect 23958 52743 24024 52753
rect 23958 52159 24024 52169
rect 25046 52743 25112 52753
rect 25046 52159 25112 52169
rect 26134 52743 26200 52753
rect 26134 52159 26200 52169
rect 27222 52743 27288 52753
rect 27222 52159 27288 52169
rect 28310 52743 28376 52753
rect 28310 52159 28376 52169
rect 29398 52743 29464 52753
rect 29398 52159 29464 52169
rect 30486 52743 30552 52753
rect 30486 52159 30552 52169
rect 31574 52743 31640 52753
rect 31574 52159 31640 52169
rect 17975 50740 18041 50750
rect 17975 50156 18041 50166
rect 20151 50740 20217 50750
rect 20151 50156 20217 50166
rect 21239 50740 21305 50750
rect 21239 50156 21305 50166
rect 23415 50740 23481 50750
rect 23415 50156 23481 50166
rect 24503 50740 24569 50750
rect 24503 50156 24569 50166
rect 25591 50740 25657 50750
rect 25591 50156 25657 50166
rect 27767 50740 27833 50750
rect 27767 50156 27833 50166
rect 28855 50740 28921 50750
rect 28855 50156 28921 50166
rect 31031 50740 31097 50750
rect 31031 50156 31097 50166
rect 17430 48743 17496 48753
rect 17430 48159 17496 48169
rect 18518 48743 18584 48753
rect 18518 48159 18584 48169
rect 19606 48743 19672 48753
rect 19606 48159 19672 48169
rect 20694 48743 20760 48753
rect 20694 48159 20760 48169
rect 21782 48743 21848 48753
rect 21782 48159 21848 48169
rect 22870 48743 22936 48753
rect 22870 48159 22936 48169
rect 23958 48743 24024 48753
rect 23958 48159 24024 48169
rect 29398 48743 29464 48753
rect 29398 48159 29464 48169
rect 30486 48743 30552 48753
rect 30486 48159 30552 48169
rect 31574 48743 31640 48753
rect 31574 48159 31640 48169
rect 10177 47607 10551 47617
rect 17975 46740 18041 46750
rect -5924 46274 -5722 46284
rect 17975 46156 18041 46166
rect 19063 46740 19129 46750
rect 19063 46156 19129 46166
rect 20151 46740 20217 46750
rect 20151 46156 20217 46166
rect 21239 46740 21305 46750
rect 21239 46156 21305 46166
rect 22327 46740 22393 46750
rect 22327 46156 22393 46166
rect 24503 46740 24569 46750
rect 24503 46156 24569 46166
rect 25591 46740 25657 46750
rect 25591 46156 25657 46166
rect 26679 46740 26745 46750
rect 26679 46156 26745 46166
rect 27767 46740 27833 46750
rect 27767 46156 27833 46166
rect 28855 46740 28921 46750
rect 28855 46156 28921 46166
rect 29943 46740 30009 46750
rect 29943 46156 30009 46166
rect 31031 46740 31097 46750
rect 40589 46375 40653 46385
rect 40589 46301 40653 46311
rect 31031 46156 31097 46166
rect 10180 46128 10551 46138
rect 344 45844 558 45854
rect -4101 45307 -3923 45317
rect -4101 45119 -3923 45129
rect -1482 44459 -1304 44469
rect 2132 44508 2310 44518
rect 2132 44320 2310 44330
rect 4132 44508 4310 44518
rect 4132 44320 4310 44330
rect 6132 44508 6310 44518
rect 6132 44320 6310 44330
rect 8132 44508 8310 44518
rect 8132 44320 8310 44330
rect 344 44308 558 44318
rect -1482 44271 -1304 44281
rect 352 41383 512 41393
rect -5924 39809 -5722 39819
rect -5684 39846 -148 39856
rect -6989 39731 -6861 39741
rect 18245 45748 18309 45758
rect 18245 45674 18309 45684
rect 18791 45748 18855 45758
rect 18791 45674 18855 45684
rect 19337 45739 19401 45749
rect 21517 45748 21581 45758
rect 19337 45665 19401 45675
rect 19882 45738 19946 45748
rect 21517 45674 21581 45684
rect 22051 45735 22115 45745
rect 19882 45664 19946 45674
rect 22051 45661 22115 45671
rect 22598 45741 22662 45751
rect 22598 45667 22662 45677
rect 23143 45741 23207 45751
rect 23143 45667 23207 45677
rect 25863 45738 25927 45748
rect 25863 45664 25927 45674
rect 26406 45742 26470 45752
rect 26406 45668 26470 45678
rect 26948 45736 27012 45746
rect 29129 45738 29193 45748
rect 26948 45662 27012 45672
rect 27505 45727 27569 45737
rect 29129 45664 29193 45674
rect 29673 45731 29737 45741
rect 27505 45653 27569 45663
rect 29673 45657 29737 45667
rect 30223 45735 30287 45745
rect 30223 45661 30287 45671
rect 30756 45735 30820 45745
rect 30756 45661 30820 45671
rect 39557 44891 39621 44901
rect 39557 44817 39621 44827
rect 40595 44830 40647 46301
rect 41146 45819 41210 45829
rect 41146 45745 41210 45755
rect 40988 44991 41052 45001
rect 40988 44917 41052 44927
rect 39557 44701 39621 44711
rect 39557 44627 39621 44637
rect 39557 43741 39621 43751
rect 39557 43667 39621 43677
rect 40595 43680 40647 44778
rect 40995 44819 41047 44917
rect 40894 44762 40946 44772
rect 40995 44757 41047 44767
rect 41152 44823 41204 45745
rect 44754 45074 45306 45084
rect 44754 44997 45306 45007
rect 40894 44617 40946 44710
rect 40888 44607 40952 44617
rect 40888 44533 40952 44543
rect 40988 43841 41052 43851
rect 40988 43767 41052 43777
rect 40595 43618 40647 43628
rect 40995 43669 41047 43767
rect 40894 43612 40946 43622
rect 39557 43551 39621 43561
rect 39557 43477 39621 43487
rect 40995 43607 41047 43617
rect 41152 43673 41204 44771
rect 46294 44939 46530 44949
rect 46294 44693 46530 44703
rect 41516 44527 41874 44537
rect 41516 44452 41874 44462
rect 44766 43925 45293 43935
rect 44766 43844 45293 43854
rect 41152 43611 41204 43621
rect 46282 43788 46518 43798
rect 40894 43467 40946 43560
rect 46282 43542 46518 43552
rect 40888 43457 40952 43467
rect 40888 43383 40952 43393
rect 41514 43377 41872 43387
rect 41514 43302 41872 43312
rect 40589 42685 40653 42695
rect 40589 42611 40653 42621
rect 39557 41201 39621 41211
rect 39557 41127 39621 41137
rect 40595 41140 40647 42611
rect 41146 42129 41210 42139
rect 41146 42055 41210 42065
rect 40988 41301 41052 41311
rect 40988 41227 41052 41237
rect 39557 41011 39621 41021
rect 39557 40937 39621 40947
rect 10180 39857 10551 39867
rect 39557 39931 39621 39941
rect 39557 39857 39621 39867
rect 40595 39870 40647 41088
rect 40995 41129 41047 41227
rect 40894 41072 40946 41082
rect 40995 41067 41047 41077
rect 41152 41133 41204 42055
rect 44756 41383 45283 41393
rect 44756 41302 45283 41312
rect 40894 40927 40946 41020
rect 40888 40917 40952 40927
rect 40888 40843 40952 40853
rect 40988 40031 41052 40041
rect 40988 39957 41052 39967
rect 352 39845 512 39855
rect 40595 39808 40647 39818
rect 40995 39859 41047 39957
rect 40894 39802 40946 39812
rect 39557 39741 39621 39751
rect 39557 39667 39621 39677
rect 40995 39797 41047 39807
rect 41152 39863 41204 41081
rect 46140 41256 46376 41266
rect 46140 41010 46376 41020
rect 41432 40836 41790 40846
rect 41432 40761 41790 40771
rect 44756 40113 45283 40123
rect 44756 40032 45283 40042
rect 41152 39801 41204 39811
rect 46111 39966 46347 39976
rect -5684 39656 -148 39666
rect 40894 39657 40946 39750
rect 46111 39720 46347 39730
rect 40888 39647 40952 39657
rect 40888 39573 40952 39583
rect 41430 39567 41788 39577
rect -27077 39466 -26990 39476
rect -18883 39537 -18807 39547
rect -31812 39166 -31748 39176
rect -31812 38817 -31748 38827
rect -27082 39120 -26998 39130
rect -31811 38613 -31747 38623
rect -29614 38413 -29150 38423
rect -29614 38339 -29150 38349
rect -31030 38256 -30901 38266
rect -31047 38192 -31030 38256
rect -30901 38192 -30885 38256
rect -27082 38222 -26998 38232
rect -31811 38131 -31747 38141
rect -35518 37568 -35282 37578
rect -35518 37322 -35282 37332
rect -31030 27930 -30901 38192
rect -30199 37475 -30070 37496
rect -30217 37411 -30199 37475
rect -30070 37411 -30055 37475
rect -30199 29288 -30070 37411
rect -27079 37353 -26995 37363
rect -29652 37323 -29143 37333
rect -29652 37249 -29143 37259
rect -27079 36455 -26995 36465
rect -27077 36160 -26996 36170
rect 41430 39492 41788 39502
rect 7082 39210 7318 39220
rect 12542 39210 12778 39220
rect 7318 38974 12542 39210
rect 7082 38964 7318 38974
rect 12542 38964 12778 38974
rect 1473 38878 1537 38888
rect 1473 38804 1537 38814
rect 2513 38881 2595 38891
rect 2513 38632 2595 38642
rect 93 38566 157 38576
rect 1230 38566 1294 38576
rect 87 38502 93 38566
rect 157 38502 1230 38566
rect 93 38492 157 38502
rect 1230 38492 1294 38502
rect 2626 38568 2690 38578
rect 5361 38568 5425 38578
rect 2690 38504 5361 38568
rect 2626 38494 2690 38504
rect 5361 38494 5425 38504
rect 2515 38420 2614 38430
rect 1996 38069 2060 38079
rect 1996 37995 2060 38005
rect 5361 38155 5425 38165
rect 7236 38155 7300 38165
rect 5425 38091 7236 38155
rect 5361 38081 5425 38091
rect 7236 38081 7300 38091
rect 2515 37986 2614 37996
rect 93 37651 157 37661
rect 3427 37651 3491 37661
rect 9428 37651 9492 37661
rect 157 37587 3427 37651
rect 3491 37587 9428 37651
rect 93 37577 157 37587
rect 3427 37577 3491 37587
rect 9428 37577 9492 37587
rect 2644 37207 2708 37217
rect 5429 37207 5493 37217
rect 6701 37207 6765 37217
rect 2168 37149 2232 37159
rect 1473 37129 1537 37139
rect 1473 37055 1537 37065
rect 2708 37143 5429 37207
rect 5493 37143 6701 37207
rect 2644 37133 2708 37143
rect 5429 37133 5493 37143
rect 6701 37133 6765 37143
rect 2168 36888 2232 36898
rect 93 36816 157 36826
rect 883 36816 947 36826
rect 90 36752 93 36816
rect 157 36752 883 36816
rect 93 36742 157 36752
rect 883 36742 947 36752
rect 2169 36668 2233 36678
rect 1996 36319 2060 36329
rect 1996 36245 2060 36255
rect 6345 36597 6409 36607
rect 2169 36240 2233 36250
rect 4938 36539 6345 36591
rect -18883 36114 -18807 36124
rect 2938 36088 3343 36098
rect 2938 36020 3343 36030
rect 3582 36094 3811 36104
rect 3582 36020 3811 36030
rect 4938 35863 4990 36539
rect 6409 36539 7804 36591
rect 6345 36523 6409 36533
rect 6345 36253 6409 36263
rect 5990 36195 6345 36247
rect 5055 36104 5351 36114
rect 5055 36008 5351 36018
rect 5574 36097 5801 36107
rect 5574 36017 5801 36027
rect 5990 35969 6042 36195
rect 6409 36195 6740 36247
rect 6345 36179 6409 36189
rect 5747 35917 6042 35969
rect 6688 35969 6740 36195
rect 6936 36089 7157 36099
rect 6936 36010 7157 36020
rect 7383 36094 7681 36104
rect 7383 36018 7681 36028
rect 6688 35917 6989 35969
rect 7752 35941 7804 36539
rect 8921 36093 9348 36103
rect 8921 36018 9348 36028
rect 9575 36091 9802 36101
rect 9575 36013 9802 36023
rect -27077 34975 -26996 34985
rect 5430 35020 5494 35030
rect -27079 34691 -27000 34701
rect -9369 34676 -9305 34686
rect -9369 34602 -9305 34612
rect 2938 34183 2990 34704
rect 5430 34425 5494 34956
rect 5430 34351 5494 34361
rect 7242 35018 7306 35028
rect 7242 34425 7306 34954
rect 7242 34351 7306 34361
rect 5932 34195 5996 34205
rect 2938 34131 5932 34183
rect 8938 34183 8990 34790
rect 5996 34131 8990 34183
rect 5932 34121 5996 34131
rect 3745 33850 3797 33860
rect 6738 33850 6802 33860
rect 9745 33850 9797 33860
rect 3797 33798 6738 33850
rect 3745 33788 3797 33798
rect 6802 33798 9745 33850
rect 9797 33798 9798 33850
rect 9745 33788 9797 33798
rect 6738 33776 6802 33786
rect 5430 33561 5494 33574
rect -27079 33488 -27000 33498
rect -21518 33551 -21454 33561
rect -21518 33477 -21454 33487
rect -6948 33179 -6884 33189
rect -6948 33105 -6884 33115
rect -27084 32899 -27005 32909
rect -27084 32355 -27005 32365
rect 5317 32345 5381 32355
rect 5430 32345 5494 33497
rect 7428 33569 7492 33579
rect 7428 32362 7492 33505
rect 5381 32281 5494 32345
rect 7364 32352 7492 32362
rect 7428 32288 7492 32352
rect 5317 32271 5381 32281
rect 7364 32278 7428 32288
rect -6989 31811 8057 31840
rect -6861 31747 7965 31811
rect 8029 31747 8057 31811
rect -6989 31712 8057 31747
rect 4354 30432 4418 30442
rect 4354 30358 4418 30368
rect 8328 30437 8392 30447
rect 8328 30363 8392 30373
rect -9347 30315 2453 30338
rect -9397 30305 2453 30315
rect 3326 30305 3390 30315
rect -9269 30241 3326 30305
rect -9397 30231 2453 30241
rect 3326 30231 3390 30241
rect -9347 30210 2453 30231
rect -12693 29752 -12629 29762
rect -12693 29678 -12629 29688
rect 1913 29752 1977 29762
rect 16721 29752 16785 29762
rect 1977 29688 16721 29752
rect 1913 29678 1977 29688
rect 16721 29678 16785 29688
rect -13469 29329 -13405 29339
rect -30199 29149 -30070 29159
rect -18523 29288 -18394 29298
rect -13469 29255 -13405 29265
rect 1913 29329 1977 29339
rect 17412 29329 17476 29339
rect 1977 29265 17412 29329
rect 1913 29255 1977 29265
rect 17412 29255 17476 29265
rect -31030 27791 -30901 27801
rect -19383 27930 -19254 27940
rect -38190 26611 -34856 26621
rect -38190 26504 -34856 26514
rect -19383 26015 -19254 27801
rect -18523 27609 -18394 29159
rect 7960 28846 8024 28856
rect 1951 28808 2079 28818
rect 4701 28808 4765 28818
rect 2079 28744 4701 28808
rect 7960 28772 8024 28782
rect 1951 28734 2079 28744
rect 4701 28734 4765 28744
rect -6086 28608 -5958 28633
rect -15712 28098 -15613 28108
rect -17635 27644 -17507 27654
rect -18523 27575 -18246 27609
rect -18523 27511 -18326 27575
rect -18262 27511 -18246 27575
rect -18523 27480 -18246 27511
rect -12389 28076 -12316 28086
rect -15712 27635 -15613 27645
rect -13983 28066 -13931 28076
rect -17635 27506 -17507 27516
rect -14906 27571 -14854 27581
rect -18326 27098 -18262 27108
rect -18262 27034 -17257 27098
rect -14906 27083 -14854 27519
rect -18326 27024 -18262 27034
rect -18881 26760 -18817 26770
rect -17256 26760 -17192 26770
rect -18817 26696 -17256 26760
rect -18881 26686 -18817 26696
rect -17256 26686 -17192 26696
rect -17635 26415 -17507 26425
rect -17635 26277 -17507 26287
rect -15725 26281 -15636 26291
rect -15725 26034 -15636 26044
rect -19383 25977 -18816 26015
rect -19383 25913 -18882 25977
rect -18818 25913 -18816 25977
rect -19383 25886 -18816 25913
rect -14906 25967 -14854 27031
rect -14906 25905 -14854 25915
rect -14404 27259 -14352 27269
rect -14404 25659 -14352 27207
rect -13983 26466 -13931 28014
rect -12389 27660 -12316 27670
rect -12394 27427 -12297 27437
rect -12394 27188 -12297 27198
rect -10016 26588 -9888 26598
rect -13983 25674 -13931 26414
rect -12396 26486 -12301 26496
rect -12396 26047 -12301 26057
rect -12384 25823 -12321 25833
rect -25551 25527 -24848 25579
rect -25449 25482 -25369 25492
rect -40593 25171 -40357 25181
rect -25449 25165 -25369 25175
rect -40593 24925 -40357 24935
rect -32991 25112 -32863 25122
rect -38182 23605 -34852 23615
rect -38182 23493 -34852 23503
rect -38168 19065 -34861 19075
rect -38168 18977 -34861 18987
rect -40596 17630 -40360 17640
rect -40596 17384 -40360 17394
rect -38174 16075 -34852 16085
rect -38174 15977 -34852 15987
rect -32991 14102 -32863 24984
rect -25452 24945 -25365 24955
rect -27178 24719 -26676 24771
rect -27178 21000 -27126 24719
rect -25452 24704 -25365 24714
rect -27939 20948 -27126 21000
rect -32991 13964 -32863 13974
rect -31130 17582 -31002 17592
rect -31130 6337 -31002 17454
rect -27939 15451 -27887 20948
rect -27178 17229 -27126 20948
rect -24900 21808 -24848 25527
rect -15727 25447 -15632 25457
rect -17635 25002 -17507 25012
rect -15727 25008 -15632 25018
rect -14404 24882 -14352 25607
rect -13989 25664 -13925 25674
rect -13989 25590 -13925 25600
rect -12384 25594 -12321 25604
rect -17635 24864 -17507 24874
rect -14410 24872 -14346 24882
rect -14410 24798 -14346 24808
rect -13983 24866 -13931 25590
rect -18881 24456 -18817 24466
rect -18885 24392 -18881 24456
rect -18817 24392 -17231 24456
rect -14908 24441 -14856 24451
rect -18881 24382 -18817 24392
rect -18326 24117 -18262 24127
rect -17255 24117 -17191 24127
rect -18334 24053 -18326 24117
rect -18262 24053 -17255 24117
rect -18326 24043 -18262 24053
rect -17255 24043 -17191 24053
rect -17635 23773 -17507 23783
rect -17635 23635 -17507 23645
rect -15725 23637 -15658 23647
rect -15725 23395 -15658 23405
rect -14908 22771 -14856 24389
rect -14908 22713 -14856 22719
rect -14404 24059 -14352 24798
rect -14404 22459 -14352 24007
rect -13983 23266 -13931 24814
rect -12393 24712 -12328 24722
rect -12393 24448 -12328 24458
rect -12398 24239 -12316 24249
rect -12398 23993 -12316 24003
rect -13983 23203 -13931 23214
rect -12389 23277 -12319 23287
rect -12389 22847 -12319 22857
rect -11601 22776 -11473 22786
rect -14404 22397 -14352 22407
rect -12391 22624 -12323 22634
rect -12391 22389 -12323 22399
rect -11601 21851 -11473 22712
rect -24900 21756 -24087 21808
rect -24900 18038 -24848 21756
rect -25557 17986 -24848 18038
rect -25452 17922 -25387 17932
rect -25452 17617 -25387 17627
rect -25450 17404 -25378 17414
rect -27178 17177 -26752 17229
rect -25450 17159 -25378 17169
rect -24139 16259 -24087 21756
rect -24191 16249 -24087 16259
rect -24191 16185 -24170 16249
rect -24106 16185 -24087 16249
rect -24191 16175 -24087 16185
rect -27939 15441 -27835 15451
rect -27939 15377 -27920 15441
rect -27856 15377 -27835 15441
rect -27939 15367 -27835 15377
rect -27939 9871 -27887 15367
rect -25572 14514 -24916 14562
rect -25575 14513 -24916 14514
rect -25572 14510 -24916 14513
rect -25517 14446 -25444 14456
rect -25517 14147 -25444 14157
rect -25518 13925 -25446 13935
rect -27246 13723 -26815 13755
rect -27246 13714 -26812 13723
rect -27246 13703 -26815 13714
rect -27246 9871 -27194 13703
rect -25518 13680 -25446 13690
rect -27939 9819 -27194 9871
rect -31130 6199 -31002 6209
rect -27246 5987 -27194 9819
rect -24968 10677 -24916 14510
rect -24139 10677 -24087 16175
rect -13972 21723 -11473 21851
rect -18223 14073 -18159 14083
rect -18223 13999 -18159 14009
rect -24968 10625 -24087 10677
rect -24968 6793 -24916 10625
rect -13972 10181 -13844 21723
rect -10016 21076 -9888 26524
rect -6086 21671 -5958 28544
rect 3399 28595 3463 28605
rect 4328 28595 4392 28605
rect 3463 28531 4328 28595
rect 4392 28531 4398 28595
rect 8338 28592 8402 28602
rect 9399 28592 9463 28602
rect 3399 28521 3463 28531
rect 4328 28521 4392 28531
rect 8402 28528 9399 28592
rect 9463 28528 9473 28592
rect 8338 28518 8402 28528
rect 9399 28518 9463 28528
rect -5279 27532 -5215 27542
rect -5215 27468 19935 27532
rect -5279 27458 -5215 27468
rect -3918 26855 -3854 26865
rect -3854 26791 17577 26855
rect -3918 26781 -3854 26791
rect 1952 25820 2080 25830
rect 7960 25820 8024 25830
rect 2080 25756 7960 25820
rect 1952 25746 2080 25756
rect 7960 25746 8024 25756
rect -6086 21597 -5958 21607
rect -3501 25414 -3373 25433
rect -12387 20948 -9888 21076
rect -12387 17968 -12259 20948
rect -3501 20809 -3373 25350
rect 17513 24802 17577 26791
rect 19871 26009 19935 27468
rect 19871 25935 19935 25945
rect 19873 25598 19937 25608
rect 19873 24802 19937 25534
rect 17513 24738 19937 24802
rect 5715 24594 5783 24604
rect 7068 24592 7132 24602
rect 7068 24518 7132 24528
rect 5715 24176 5783 24186
rect 42856 24174 46190 24184
rect 3399 24101 3463 24109
rect 5643 24097 5707 24107
rect 3463 24037 5643 24097
rect 3399 24033 5643 24037
rect 3399 24027 3463 24033
rect 5643 24023 5707 24033
rect 7017 24101 7081 24111
rect 9399 24101 9463 24111
rect 7081 24037 9399 24101
rect 9463 24037 9467 24101
rect 42856 24055 46190 24065
rect 7017 24027 7081 24037
rect 9399 24027 9463 24037
rect 36066 24018 36130 24028
rect 35939 23960 36066 24012
rect 36066 23944 36130 23954
rect 35152 23866 35216 23876
rect 35152 23792 35216 23802
rect 7091 23652 7155 23782
rect 39346 23714 39420 23724
rect 7091 23578 7155 23588
rect 37819 23611 37892 23621
rect 37819 23482 37892 23492
rect 39346 23483 39420 23493
rect 8787 23356 8943 23366
rect 8787 23236 8943 23246
rect 37819 23194 37905 23204
rect 2550 23063 2614 23073
rect 2550 22989 2614 22999
rect 10202 23063 10266 23073
rect 10202 22989 10266 22999
rect 37819 22936 37905 22946
rect 39335 23200 39421 23210
rect 39335 22942 39421 22952
rect 35100 22790 35280 22800
rect 35760 22730 36021 22740
rect 35760 22658 36021 22668
rect 47556 22734 47792 22744
rect 35100 22600 35280 22610
rect 47556 22488 47792 22498
rect 39346 22388 39420 22398
rect 37826 22280 37896 22290
rect 39346 22157 39420 22167
rect 37826 22141 37896 22151
rect 13887 22124 13951 22134
rect 4397 22037 4449 22047
rect -3501 20735 -3373 20745
rect -971 21625 -907 21635
rect -971 20715 -907 21561
rect 2910 21612 2962 22014
rect 3779 21985 4397 22037
rect 4397 21975 4449 21985
rect 8228 22037 8280 22047
rect 8280 21985 9098 22037
rect 8228 21975 8280 21985
rect 6312 21635 6364 21664
rect 6307 21625 6371 21635
rect 2910 21561 6307 21612
rect 9905 21612 9957 22096
rect 6371 21561 9957 21612
rect 2910 21560 9957 21561
rect 6307 21551 6371 21560
rect 6312 20967 6364 20997
rect 6310 20957 6374 20967
rect 4397 20945 4449 20955
rect 4387 20893 4397 20945
rect 4449 20893 6310 20945
rect 8228 20945 8280 20955
rect 6374 20893 8228 20945
rect 8280 20893 8290 20945
rect 4397 20883 4449 20893
rect 6310 20883 6374 20893
rect 8228 20883 8280 20893
rect -971 20641 -907 20651
rect -444 20109 -380 20119
rect 5394 20109 5458 20119
rect 9394 20109 9458 20119
rect -12387 17904 -12355 17968
rect -12291 17904 -12259 17968
rect -10970 19981 -444 20109
rect -380 19981 5394 20109
rect 5458 19981 9394 20109
rect 9458 19981 9474 20109
rect -12355 17894 -12291 17904
rect -13064 14141 -13000 14151
rect -13064 14067 -13000 14077
rect -13972 10117 -13941 10181
rect -13877 10117 -13844 10181
rect -10970 10223 -10842 19981
rect -444 19971 -380 19981
rect 5394 19971 5458 19981
rect 9394 19971 9458 19981
rect 51 19513 115 19523
rect -756 19212 -692 19222
rect -756 19049 -692 19148
rect 51 19051 115 19449
rect 1684 19410 1748 19420
rect 7394 19410 7458 19420
rect 1748 19346 7394 19410
rect 1748 19282 3395 19346
rect 3459 19282 7394 19346
rect 7458 19282 7468 19410
rect 1684 19272 1748 19282
rect 3395 19272 3459 19282
rect 7394 19272 7458 19282
rect 4857 19173 5194 19183
rect 3061 19106 3125 19116
rect 3061 19032 3125 19042
rect 7085 19106 7149 19116
rect 7085 19032 7149 19042
rect 8981 19106 9045 19116
rect 8981 19032 9045 19042
rect 10232 19058 10296 19068
rect 4857 19017 5194 19027
rect 10232 18984 10296 18994
rect 5707 18910 5771 18920
rect 5707 18836 5771 18846
rect 7706 18910 7770 18920
rect 7706 18836 7770 18846
rect 8280 18718 8344 18728
rect 4899 18651 4963 18661
rect 4899 18577 4963 18587
rect 6897 18651 6961 18661
rect 8280 18644 8344 18654
rect 13574 18688 13638 18698
rect 13574 18614 13638 18624
rect 6897 18577 6961 18587
rect 3707 18312 3771 18322
rect 3707 18238 3771 18248
rect 9706 18312 9770 18322
rect 9706 18238 9770 18248
rect 13887 18047 13951 21996
rect 39341 21834 39427 21844
rect 37814 21823 37899 21833
rect 37814 21611 37899 21621
rect 35152 21585 35216 21595
rect 39341 21576 39427 21586
rect 35152 21511 35216 21521
rect 35477 21379 35541 21389
rect 35475 21321 35477 21373
rect 35939 21373 35991 21544
rect 35541 21321 35991 21373
rect 35477 21305 35541 21315
rect 42854 21178 46188 21188
rect 42854 21059 46188 21069
rect 14688 21027 14752 21037
rect 14688 20953 14752 20963
rect 23670 20216 23734 20226
rect 22767 20152 23670 20216
rect 14686 19278 14750 19288
rect 14686 19204 14750 19214
rect 20971 19062 21035 19072
rect 22767 19062 22831 20152
rect 23670 20142 23734 20152
rect 23689 19382 23753 19392
rect 23689 19308 23753 19318
rect 21035 18998 22831 19062
rect 20971 18988 21035 18998
rect 22767 18428 22831 18998
rect 23658 18428 23722 18438
rect 22767 18364 23658 18428
rect 23658 18354 23722 18364
rect 2898 18031 2962 18041
rect 2898 17957 2962 17967
rect 8899 18031 8963 18041
rect 13887 17973 13951 17983
rect 8899 17957 8963 17967
rect 233 17772 297 17782
rect 233 17698 297 17708
rect 14689 17549 14753 17559
rect -821 17525 -757 17535
rect 14689 17475 14753 17485
rect 23689 17552 23753 17562
rect 23689 17478 23753 17488
rect -821 17451 -757 17461
rect 7393 17359 7457 17369
rect 9396 17359 9460 17369
rect 13885 17359 13949 17369
rect 4295 17289 4359 17299
rect -445 17221 -381 17231
rect 1684 17221 1748 17231
rect -10479 17157 -445 17221
rect -10479 17093 -10416 17157
rect -10352 17093 -445 17157
rect -381 17093 1684 17221
rect 4295 17215 4359 17225
rect 6227 17289 6291 17299
rect 6227 17215 6291 17225
rect 7457 17231 9396 17359
rect 9460 17231 13885 17359
rect 13949 17231 13962 17359
rect 7393 17221 7457 17231
rect 9396 17221 9460 17231
rect 13885 17221 13949 17231
rect -10479 17092 1748 17093
rect -10416 17083 -10352 17092
rect -445 17083 -381 17092
rect 1684 17083 1748 17092
rect 13603 17083 13667 17093
rect 14690 17083 14754 17093
rect 13667 17019 14690 17083
rect 13603 17009 13667 17019
rect 14690 17009 14754 17019
rect 3393 16866 3457 16876
rect 5393 16866 5457 16876
rect 13277 16866 13341 16876
rect 3457 16738 5393 16866
rect 5457 16738 13277 16866
rect 13341 16738 13351 16866
rect 3393 16728 3457 16738
rect 5393 16728 5457 16738
rect 13277 16728 13341 16738
rect 251 16446 11139 16456
rect -10415 16288 -10351 16298
rect -3926 16288 -3862 16298
rect -10351 16224 -3926 16288
rect 251 16228 11139 16238
rect -10415 16214 -10351 16224
rect -3926 16214 -3862 16224
rect -5786 15708 -5722 15718
rect -5786 15634 -5722 15644
rect -3914 15135 -3862 16214
rect 28 16189 187 16199
rect -3008 15454 -2944 15464
rect -3008 15380 -2944 15390
rect -5026 14663 -4390 14715
rect -5026 14411 -4974 14663
rect -4902 14446 -4832 14456
rect -4902 14226 -4832 14236
rect -6544 14141 -6480 14151
rect -6544 12892 -6480 14077
rect -4917 13998 -4833 14008
rect -4917 13696 -4833 13706
rect -5006 13597 -4731 13649
rect -6544 12818 -6480 12828
rect -5851 12892 -5787 12902
rect -5851 12219 -5787 12828
rect -5851 12145 -5787 12155
rect -5845 10943 -5793 10953
rect -6411 10890 -6103 10942
rect -6411 10701 -6359 10890
rect -6162 10833 -5937 10843
rect -6162 10748 -5937 10758
rect -6411 10649 -6104 10701
rect -10906 10159 -10842 10223
rect -10970 10139 -10842 10159
rect -6156 10214 -6104 10649
rect -5845 10412 -5793 10891
rect -5707 10838 -5401 10848
rect -5707 10741 -5401 10751
rect -5845 10402 -5792 10412
rect -5845 10339 -5792 10349
rect -6156 10204 -6092 10214
rect -13972 10113 -13844 10117
rect -6156 10130 -6092 10140
rect -13941 10107 -13877 10113
rect -6156 9717 -6104 10130
rect -6383 9665 -6104 9717
rect -6383 9453 -6331 9665
rect -6167 9592 -5929 9602
rect -6167 9503 -5929 9513
rect -6383 9401 -6110 9453
rect -5845 9452 -5793 10339
rect -5348 10214 -5296 10935
rect -4783 10243 -4731 13597
rect -4442 10243 -4390 14663
rect -3914 14139 -3862 15083
rect -678 15136 -626 15146
rect -3144 14998 -3061 15008
rect -3144 14709 -3061 14719
rect -3023 14644 -2959 14654
rect -3023 14570 -2959 14580
rect -3914 12635 -3862 14087
rect -2598 13137 -2534 13147
rect -2598 13063 -2534 13073
rect -1808 13133 -1725 13143
rect -1808 12716 -1725 12726
rect -5361 10204 -5296 10214
rect -5363 10146 -5361 10198
rect -5297 10140 -5296 10204
rect -4789 10233 -4725 10243
rect -4789 10159 -4725 10169
rect -4448 10233 -4384 10243
rect -4448 10159 -4384 10169
rect -5361 10130 -5296 10140
rect -5708 9595 -5399 9605
rect -5708 9499 -5399 9509
rect -5348 9406 -5296 10130
rect -5845 9390 -5793 9400
rect -5853 8174 -5789 8184
rect -6565 7591 -6501 7601
rect -7214 7243 -6751 7253
rect -7214 6993 -6751 7003
rect -25628 6741 -24916 6793
rect -25521 6669 -25446 6679
rect -25521 6398 -25446 6408
rect -13075 6313 -13011 6323
rect -18251 6303 -18187 6313
rect -13075 6239 -13011 6249
rect -6565 6313 -6501 7527
rect -5853 7595 -5789 8110
rect -5853 7521 -5789 7531
rect -4783 6803 -4731 10159
rect -5036 6751 -4731 6803
rect -4917 6695 -4836 6705
rect -4917 6382 -4836 6392
rect -6565 6239 -6501 6249
rect -18251 6229 -18187 6239
rect -25522 6174 -25447 6184
rect -27246 5936 -26782 5987
rect -27165 5935 -26782 5936
rect -4907 6163 -4841 6173
rect -25522 5919 -25447 5929
rect -5029 5826 -4977 5994
rect -4907 5940 -4841 5950
rect -4442 5826 -4390 10159
rect -3914 9437 -3862 12583
rect -1498 12409 -1434 12419
rect -2885 12328 -2821 12338
rect -1498 12335 -1434 12345
rect -2885 12254 -2821 12264
rect -1926 11535 -1862 11545
rect -1926 11461 -1862 11471
rect -1759 11529 -1693 11539
rect -1759 11130 -1693 11140
rect -3914 9375 -3862 9385
rect -3415 11034 -3363 11044
rect -5029 5774 -4390 5826
rect -3415 7835 -3363 10982
rect -1498 10783 -1434 10793
rect -2212 10729 -2148 10739
rect -1498 10709 -1434 10719
rect -2212 10655 -2148 10665
rect -678 10402 -626 15084
rect -1926 9937 -1862 9947
rect -1926 9863 -1862 9873
rect -1759 9930 -1695 9940
rect -1759 9522 -1695 9532
rect -1149 9435 -1097 9451
rect -2212 9129 -2148 9139
rect -2212 9055 -2148 9065
rect -1498 9125 -1434 9135
rect -1498 9051 -1434 9061
rect -2598 8335 -2534 8345
rect -2598 8261 -2534 8271
rect -1758 8330 -1690 8340
rect -1758 7920 -1690 7930
rect -3415 6310 -3363 7783
rect -1149 7835 -1097 9383
rect -1498 7586 -1434 7596
rect -2885 7527 -2821 7537
rect -1498 7512 -1434 7522
rect -2885 7453 -2821 7463
rect -1498 7258 -1434 7268
rect -1498 6964 -1434 6974
rect -1498 6451 -1434 6461
rect -1498 6377 -1434 6387
rect -3415 5723 -3363 6258
rect -3050 6042 -2986 6052
rect -3050 5968 -2986 5978
rect -3415 5057 -3363 5671
rect -3193 5577 -3110 5587
rect -3193 5286 -3110 5296
rect -3028 5233 -2964 5243
rect -3028 5159 -2964 5169
rect -1149 5129 -1097 7783
rect -678 5723 -626 10350
rect -678 5661 -626 5671
rect -279 12637 -227 12647
rect -279 11035 -227 12585
rect -1149 5067 -1097 5077
rect -10766 5047 -10702 5057
rect -3427 5047 -3363 5057
rect -10702 4983 -3427 5047
rect -10766 4973 -10702 4983
rect -3427 4973 -3363 4983
rect -279 3789 -227 10983
rect 11239 16184 11399 16194
rect 5478 14599 5656 14609
rect 5478 14411 5656 14421
rect 23686 15788 23750 15798
rect 14685 15753 14749 15763
rect 23686 15714 23750 15724
rect 14685 15679 14749 15689
rect 20928 15496 20992 15506
rect 20928 15422 20992 15432
rect 14690 15228 14754 15238
rect 14690 15154 14754 15164
rect 11239 14416 11399 14426
rect 23686 13997 23750 14007
rect 14685 13965 14749 13975
rect 11257 13954 11384 13964
rect 23686 13923 23750 13933
rect 14685 13891 14749 13901
rect 13636 13528 13700 13538
rect 14690 13528 14754 13538
rect 13700 13464 14690 13528
rect 13636 13454 13700 13464
rect 14690 13454 14754 13464
rect 23685 13006 23749 13016
rect 11257 12980 11384 12990
rect 23094 12942 23685 13006
rect 14702 12180 14766 12190
rect 11243 12129 11398 12139
rect 4630 11980 4808 11990
rect 4630 11792 4808 11802
rect 14702 12106 14766 12116
rect 20985 11906 21049 11916
rect 23094 11906 23158 12942
rect 23685 12932 23749 12942
rect 23691 12190 23755 12200
rect 23691 12116 23755 12126
rect 20968 11842 20985 11906
rect 21049 11842 23753 11906
rect 20985 11832 21049 11842
rect 13699 11676 13763 11686
rect 14692 11676 14756 11686
rect 13763 11612 14692 11676
rect 13699 11602 13763 11612
rect 14692 11602 14756 11612
rect 23689 11519 23753 11842
rect 23689 11445 23753 11455
rect 11243 11306 11398 11316
rect 28 10630 187 10640
rect 6483 10537 11218 10547
rect 6483 10346 11218 10356
rect 14691 10383 14755 10393
rect 14691 10309 14755 10319
rect 23691 10380 23755 10390
rect 23691 10306 23755 10316
rect 372 10144 1812 10154
rect 13876 10150 21118 10160
rect 372 9993 1812 10003
rect 5727 10135 11722 10145
rect 5727 9980 11722 9990
rect 13876 9983 21118 9993
rect 29 9830 212 9840
rect 5223 9418 5276 9428
rect 24544 9424 24608 9434
rect 5276 9365 24544 9418
rect 5223 9355 5276 9365
rect 24544 9350 24608 9360
rect 36066 9154 36130 9164
rect 17646 8451 17824 8461
rect 4679 8366 4857 8376
rect 17646 8263 17824 8273
rect 4679 8178 4857 8188
rect 23208 7845 23261 7855
rect 17672 7792 23208 7845
rect 17672 7717 17725 7792
rect 23208 7782 23261 7792
rect 12920 7664 17725 7717
rect 25495 7651 25559 9116
rect 35842 9096 36066 9150
rect 35489 8531 35553 8541
rect 35489 8457 35553 8467
rect 35842 8400 35896 9096
rect 36066 9080 36130 9090
rect 36631 8469 36695 8479
rect 35982 8413 36631 8465
rect 36631 8395 36695 8405
rect 35024 8283 35088 8293
rect 35024 8209 35088 8219
rect 40100 8121 40181 8131
rect 38575 8038 38645 8048
rect 40100 7923 40181 7933
rect 36301 7881 36532 7891
rect 38575 7882 38645 7892
rect 36301 7804 36532 7814
rect 33746 7651 33810 7661
rect 25495 7587 33746 7651
rect 33746 7577 33810 7587
rect 40087 7576 40168 7586
rect 38568 7563 38649 7573
rect 21250 7514 21417 7524
rect 13350 6491 13528 6501
rect 4679 6366 4857 6376
rect 13350 6303 13528 6313
rect 17646 6451 17824 6461
rect 17646 6263 17824 6273
rect 4679 6178 4857 6188
rect 29 5560 212 5570
rect 16101 5088 16279 5098
rect 16101 4900 16279 4910
rect 19101 5088 19279 5098
rect 19101 4900 19279 4910
rect 40087 7378 40168 7388
rect 38568 7365 38649 7375
rect 36362 7337 36531 7347
rect 36362 7265 36531 7275
rect 35028 7223 35092 7233
rect 35028 7149 35092 7159
rect 42602 7232 45923 7242
rect 42602 7133 45923 7143
rect 35027 6954 35091 6964
rect 35027 6880 35091 6890
rect 36352 6795 36437 6805
rect 36352 6711 36437 6721
rect 40092 6785 40173 6795
rect 38571 6707 38649 6717
rect 40092 6587 40173 6597
rect 38571 6572 38649 6582
rect 24544 6312 24608 6322
rect 33734 6312 33798 6322
rect 24608 6248 33734 6312
rect 24544 6238 24608 6248
rect 33734 6238 33798 6248
rect 36971 6265 37067 6275
rect 36971 6159 37067 6169
rect 38563 6232 38644 6242
rect 38563 6034 38644 6044
rect 40092 6229 40173 6239
rect 40092 6031 40173 6041
rect 35027 5885 35091 5895
rect 35027 5811 35091 5821
rect 47473 5800 47709 5810
rect 35970 5707 36149 5717
rect 35970 5634 36149 5644
rect 35024 5562 35088 5572
rect 47473 5554 47709 5564
rect 35024 5488 35088 5498
rect 40109 5405 40190 5415
rect 38574 5322 38648 5332
rect 40109 5207 40190 5217
rect 38574 5177 38648 5187
rect 36514 5162 36734 5172
rect 36514 5082 36734 5092
rect 23208 4916 23261 4926
rect 33742 4916 33795 4926
rect 23261 4863 33742 4916
rect 23208 4853 23261 4863
rect 33742 4853 33795 4863
rect 38562 4879 38643 4889
rect 38562 4681 38643 4691
rect 40092 4857 40173 4867
rect 40092 4659 40173 4669
rect 36364 4613 36509 4623
rect 36364 4545 36509 4555
rect 21250 4530 21417 4540
rect 35035 4492 35099 4502
rect 35035 4418 35099 4428
rect 4679 4366 4857 4376
rect 42599 4233 45959 4243
rect 4679 4178 4857 4188
rect 35024 4187 35088 4197
rect 42599 4134 45959 4144
rect 35024 4113 35088 4123
rect 36972 4089 37068 4099
rect 36972 3983 37068 3993
rect 40099 4026 40180 4036
rect 38572 3934 38651 3944
rect 40099 3828 40180 3838
rect 38572 3771 38651 3781
rect -279 3727 -227 3737
rect 36359 3531 36486 3541
rect 36359 3449 36486 3459
rect 38565 3479 38646 3489
rect 38565 3281 38646 3291
rect 40089 3473 40170 3483
rect 40089 3275 40170 3285
rect 35031 3122 35095 3132
rect 35031 3048 35095 3058
rect 28 2773 190 2783
rect 12207 2773 12385 2783
rect 3670 2688 5404 2741
rect 5351 2407 5404 2688
rect 12207 2585 12385 2595
rect 23432 2407 23485 2417
rect 4679 2366 4857 2376
rect 5351 2354 23432 2407
rect 23432 2344 23485 2354
rect 36066 2214 36130 2224
rect 4679 2178 4857 2188
rect 35842 2156 36066 2210
rect 21243 2139 21419 2149
rect 35489 1591 35553 1601
rect 35489 1517 35553 1527
rect 35842 1460 35896 2156
rect 36066 2140 36130 2150
rect 36631 1529 36695 1539
rect 35982 1473 36631 1525
rect 36631 1455 36695 1465
rect 21243 1278 21419 1288
rect 35024 1343 35088 1353
rect 35024 1269 35088 1279
rect 40100 1181 40181 1191
rect 22589 1097 22642 1107
rect 18808 1044 22589 1097
rect 22589 1034 22642 1044
rect 38575 1098 38645 1108
rect 40100 983 40181 993
rect 36301 941 36532 951
rect 38575 942 38645 952
rect 36301 864 36532 874
rect 26001 716 26076 726
rect 33730 721 33805 726
rect 33730 716 33810 721
rect 26076 641 33730 716
rect 33805 711 33810 716
rect 33805 641 33810 647
rect 26001 631 26076 641
rect 33730 637 33810 641
rect 33730 631 33805 637
rect 40087 636 40168 646
rect 38568 623 38649 633
rect 40087 438 40168 448
rect 38568 425 38649 435
rect 28 349 190 359
rect 36362 397 36531 407
rect 36362 325 36531 335
rect 42599 309 45930 319
rect 35028 283 35092 293
rect 322 232 21107 242
rect 35028 209 35092 219
rect 42599 189 45930 199
rect 322 57 21107 67
rect 35027 14 35091 24
rect 35027 -60 35091 -50
rect 36352 -145 36437 -135
rect 36352 -229 36437 -219
rect 40092 -155 40173 -145
rect 38571 -233 38649 -223
rect 40092 -353 40173 -343
rect 38571 -368 38649 -358
rect 33734 -628 33798 -618
rect 23417 -640 33734 -628
rect 23417 -693 23432 -640
rect 23485 -692 33734 -640
rect 23485 -693 33741 -692
rect 33794 -693 33798 -692
rect 23432 -703 23485 -693
rect 33734 -702 33798 -693
rect 36971 -675 37067 -665
rect 33741 -703 33794 -702
rect 36971 -781 37067 -771
rect 38563 -708 38644 -698
rect 38563 -906 38644 -896
rect 40092 -711 40173 -701
rect 40092 -909 40173 -899
rect 35027 -1055 35091 -1045
rect 35027 -1129 35091 -1119
rect 47489 -1140 47725 -1130
rect 35970 -1233 36149 -1223
rect 35970 -1306 36149 -1296
rect 35024 -1378 35088 -1368
rect 47489 -1386 47725 -1376
rect 35024 -1452 35088 -1442
rect 40109 -1535 40190 -1525
rect 38574 -1618 38648 -1608
rect 40109 -1733 40190 -1723
rect 38574 -1763 38648 -1753
rect 36514 -1778 36734 -1768
rect 36514 -1858 36734 -1848
rect 22589 -2017 22643 -2007
rect 33757 -2014 33810 -2007
rect 33742 -2017 33810 -2014
rect 22587 -2070 22589 -2017
rect 22643 -2024 33757 -2017
rect 22643 -2070 33742 -2024
rect 22587 -2077 33742 -2070
rect 33795 -2077 33810 -2070
rect 22589 -2080 22643 -2077
rect 33742 -2080 33810 -2077
rect 38562 -2061 38643 -2051
rect 33742 -2087 33795 -2080
rect 38562 -2259 38643 -2249
rect 40092 -2083 40173 -2073
rect 40092 -2281 40173 -2271
rect 36364 -2327 36509 -2317
rect 36364 -2395 36509 -2385
rect 35035 -2448 35099 -2438
rect 35035 -2522 35099 -2512
rect 42587 -2708 45933 -2698
rect 35024 -2753 35088 -2743
rect 42587 -2806 45933 -2796
rect 35024 -2827 35088 -2817
rect 36972 -2851 37068 -2841
rect 36972 -2957 37068 -2947
rect 40099 -2914 40180 -2904
rect 38572 -3006 38651 -2996
rect 40099 -3112 40180 -3102
rect 38572 -3169 38651 -3159
rect 36359 -3409 36486 -3399
rect 36359 -3491 36486 -3481
rect 38565 -3461 38646 -3451
rect 38565 -3659 38646 -3649
rect 40089 -3467 40170 -3457
rect 40089 -3665 40170 -3655
rect 35031 -3818 35095 -3808
rect 35031 -3892 35095 -3882
rect -3595 -6822 -3503 -6812
rect -3595 -10140 -3503 -10130
rect -600 -6825 -486 -6815
rect -600 -10150 -486 -10140
rect -2179 -12082 -1943 -12072
rect -2179 -12328 -1943 -12318
<< via2 >>
rect -15410 77904 -15174 78140
rect 12606 77875 12842 78111
rect 24656 77876 24892 78112
rect -16849 73398 -16748 76723
rect -13848 73404 -13747 76729
rect 11143 73392 11271 76732
rect 14144 73405 14272 76745
rect -16664 71738 -16600 71802
rect -15486 71734 -15422 71798
rect -15269 71741 -15205 71805
rect -14135 71738 -14071 71802
rect -16554 70234 -16490 70298
rect -15440 70220 -15376 70284
rect -15227 70221 -15163 70285
rect -14063 70221 -13999 70285
rect -16708 68639 -16644 68703
rect -15963 68105 -15890 68261
rect -15422 68166 -15358 68515
rect -14879 68108 -14806 68264
rect -14199 68009 -14135 68073
rect -16577 67549 -16513 67613
rect -15422 67543 -15358 67607
rect -14304 67554 -14240 67618
rect 17430 64169 17496 64743
rect 23958 64169 24024 64743
rect 31574 64169 31640 64743
rect -9884 63338 -9442 63402
rect -8073 63340 -7631 63404
rect -6278 63336 -5836 63400
rect -4479 63334 -4037 63398
rect -2688 63338 -2246 63402
rect -886 63334 -444 63398
rect -6939 62966 -6699 63206
rect 757 62992 1287 63232
rect 17975 62166 18041 62740
rect 19063 62166 19129 62740
rect 21239 62166 21305 62740
rect 22327 62166 22393 62740
rect 23415 62166 23481 62740
rect 24503 62166 24569 62740
rect 25591 62166 25657 62740
rect 26679 62166 26745 62740
rect 28855 62166 28921 62740
rect 29943 62166 30009 62740
rect 31031 62166 31097 62740
rect -8557 54531 -8493 54595
rect -6866 54532 -6802 54596
rect -5161 54531 -5097 54595
rect -3365 54531 -3301 54595
rect -1536 54531 -1472 54595
rect -9704 54339 -9462 54403
rect -7909 54338 -7667 54402
rect -6109 54340 -5867 54404
rect -4311 54339 -4069 54403
rect -2513 54340 -2271 54404
rect -710 54339 -468 54403
rect 176 54340 240 54404
rect -8854 51014 -8770 51249
rect -7722 51183 -7658 51247
rect -27070 49656 -26726 49720
rect -26408 49349 -26157 49413
rect -26060 49360 -25996 49424
rect -25984 49114 -25640 49178
rect -27087 42779 -26990 43313
rect -13469 42997 -13405 43061
rect -12693 42334 -12629 42398
rect -27082 41002 -26995 42169
rect -21475 42099 -21411 42163
rect -27077 39476 -26990 40643
rect 347 53121 519 60827
rect 5410 58752 5588 58930
rect 2047 57297 2225 57475
rect 4047 57297 4225 57475
rect 5410 55752 5588 55930
rect 4007 53001 4185 53179
rect 7725 51858 7903 52036
rect -5688 50883 -3888 51066
rect -3362 50896 -2536 51074
rect -1655 50886 -765 51064
rect -8874 50378 -8780 50791
rect -8480 50377 -8416 50441
rect -5932 47776 -5748 50720
rect -78 47752 121 50774
rect 10177 47617 10551 60836
rect 17430 60169 17496 60743
rect 18518 60169 18584 60743
rect 19606 60169 19672 60743
rect 20694 60169 20760 60743
rect 21782 60169 21848 60743
rect 22870 60169 22936 60743
rect 23958 60169 24024 60743
rect 25046 60169 25112 60743
rect 26134 60169 26200 60743
rect 27222 60169 27288 60743
rect 28310 60169 28376 60743
rect 29398 60169 29464 60743
rect 30486 60169 30552 60743
rect 31574 60169 31640 60743
rect 17975 58166 18041 58740
rect 19063 58166 19129 58740
rect 20151 58166 20217 58740
rect 21239 58166 21305 58740
rect 22327 58166 22393 58740
rect 23415 58166 23481 58740
rect 24503 58166 24569 58740
rect 25591 58166 25657 58740
rect 26679 58166 26745 58740
rect 27767 58166 27833 58740
rect 28855 58166 28921 58740
rect 29943 58166 30009 58740
rect 31031 58166 31097 58740
rect 17430 56169 17496 56743
rect 18518 56169 18584 56743
rect 19606 56169 19672 56743
rect 20694 56169 20760 56743
rect 21782 56169 21848 56743
rect 22870 56169 22936 56743
rect 23958 56169 24024 56743
rect 25046 56169 25112 56743
rect 26134 56169 26200 56743
rect 27222 56169 27288 56743
rect 28310 56169 28376 56743
rect 29398 56169 29464 56743
rect 30486 56169 30552 56743
rect 31574 56169 31640 56743
rect 17975 54166 18041 54740
rect 19063 54166 19129 54740
rect 20151 54166 20217 54740
rect 21239 54166 21305 54740
rect 22327 54166 22393 54740
rect 23415 54166 23481 54740
rect 24503 54166 24569 54740
rect 25591 54166 25657 54740
rect 26679 54166 26745 54740
rect 27767 54166 27833 54740
rect 28855 54166 28921 54740
rect 29943 54166 30009 54740
rect 31031 54166 31097 54740
rect 17430 52169 17496 52743
rect 18518 52169 18584 52743
rect 19606 52169 19672 52743
rect 20694 52169 20760 52743
rect 21782 52169 21848 52743
rect 22870 52169 22936 52743
rect 23958 52169 24024 52743
rect 25046 52169 25112 52743
rect 26134 52169 26200 52743
rect 27222 52169 27288 52743
rect 28310 52169 28376 52743
rect 29398 52169 29464 52743
rect 30486 52169 30552 52743
rect 31574 52169 31640 52743
rect 17975 50166 18041 50740
rect 20151 50166 20217 50740
rect 21239 50166 21305 50740
rect 23415 50166 23481 50740
rect 24503 50166 24569 50740
rect 25591 50166 25657 50740
rect 27767 50166 27833 50740
rect 28855 50166 28921 50740
rect 31031 50166 31097 50740
rect 17430 48169 17496 48743
rect 18518 48169 18584 48743
rect 19606 48169 19672 48743
rect 20694 48169 20760 48743
rect 21782 48169 21848 48743
rect 22870 48169 22936 48743
rect 23958 48169 24024 48743
rect 29398 48169 29464 48743
rect 30486 48169 30552 48743
rect 31574 48169 31640 48743
rect -5924 39819 -5722 46274
rect 17975 46166 18041 46740
rect 19063 46166 19129 46740
rect 20151 46166 20217 46740
rect 21239 46166 21305 46740
rect 22327 46166 22393 46740
rect 24503 46166 24569 46740
rect 25591 46166 25657 46740
rect 26679 46166 26745 46740
rect 27767 46166 27833 46740
rect 28855 46166 28921 46740
rect 29943 46166 30009 46740
rect 31031 46166 31097 46740
rect 40589 46311 40653 46375
rect -4101 45129 -3923 45307
rect -1482 44281 -1304 44459
rect 344 44318 558 45844
rect 2132 44330 2310 44508
rect 4132 44330 4310 44508
rect 6132 44330 6310 44508
rect 8132 44330 8310 44508
rect -5684 39666 -148 39846
rect 352 39855 512 41383
rect 10180 39867 10551 46128
rect 18245 45684 18309 45748
rect 18791 45684 18855 45748
rect 19337 45675 19401 45739
rect 19882 45674 19946 45738
rect 21517 45684 21581 45748
rect 22051 45671 22115 45735
rect 22598 45677 22662 45741
rect 23143 45677 23207 45741
rect 25863 45674 25927 45738
rect 26406 45678 26470 45742
rect 26948 45672 27012 45736
rect 27505 45663 27569 45727
rect 29129 45674 29193 45738
rect 29673 45667 29737 45731
rect 30223 45671 30287 45735
rect 30756 45671 30820 45735
rect 39557 44827 39621 44891
rect 41146 45755 41210 45819
rect 40988 44927 41052 44991
rect 39557 44637 39621 44701
rect 39557 43677 39621 43741
rect 44754 45007 45306 45074
rect 40888 44543 40952 44607
rect 40988 43777 41052 43841
rect 39557 43487 39621 43551
rect 46294 44703 46530 44939
rect 41516 44462 41874 44527
rect 44766 43854 45293 43925
rect 46282 43552 46518 43788
rect 40888 43393 40952 43457
rect 41514 43312 41872 43377
rect 40589 42621 40653 42685
rect 39557 41137 39621 41201
rect 41146 42065 41210 42129
rect 40988 41237 41052 41301
rect 39557 40947 39621 41011
rect 39557 39867 39621 39931
rect 44756 41312 45283 41383
rect 40888 40853 40952 40917
rect 40988 39967 41052 40031
rect 39557 39677 39621 39741
rect 46140 41020 46376 41256
rect 41432 40771 41790 40836
rect 44756 40042 45283 40113
rect 46111 39730 46347 39966
rect 40888 39583 40952 39647
rect -31812 38827 -31748 39166
rect -31811 38141 -31747 38613
rect -29614 38349 -29150 38413
rect -27082 38232 -26998 39120
rect -35518 37332 -35282 37568
rect -29652 37259 -29143 37323
rect -27079 36465 -26995 37353
rect -27077 34985 -26996 36160
rect -18883 36124 -18807 39537
rect 41430 39502 41788 39567
rect 1473 38814 1537 38878
rect 2513 38642 2595 38881
rect 1996 38005 2060 38069
rect 2515 37996 2614 38420
rect 1473 37065 1537 37129
rect 2168 36898 2232 37149
rect 1996 36255 2060 36319
rect 2169 36250 2233 36668
rect 2938 36030 3343 36088
rect 3582 36030 3811 36094
rect 6345 36533 6409 36597
rect 5055 36018 5351 36104
rect 5574 36027 5801 36097
rect 6345 36189 6409 36253
rect 6936 36020 7157 36089
rect 7383 36028 7681 36094
rect 8921 36028 9348 36093
rect 9575 36023 9802 36091
rect -27079 33498 -27000 34691
rect -9369 34612 -9305 34676
rect 5932 34131 5996 34195
rect 6738 33786 6802 33850
rect -21518 33487 -21454 33551
rect -6948 33115 -6884 33179
rect -27084 32365 -27005 32899
rect 5317 32281 5381 32345
rect 7364 32288 7428 32352
rect 7965 31747 8029 31811
rect 4354 30368 4418 30432
rect 8328 30373 8392 30437
rect 3326 30241 3390 30305
rect -12693 29688 -12629 29752
rect 1913 29688 1977 29752
rect 16721 29688 16785 29752
rect -13469 29265 -13405 29329
rect 1913 29265 1977 29329
rect 17412 29265 17476 29329
rect -38190 26514 -34856 26611
rect 4701 28744 4765 28808
rect 7960 28782 8024 28846
rect -17635 27516 -17507 27644
rect -15712 27645 -15613 28098
rect -17635 26287 -17507 26415
rect -15725 26044 -15636 26281
rect -12389 27670 -12316 28076
rect -12394 27198 -12297 27427
rect -12396 26057 -12301 26486
rect -40593 24935 -40357 25171
rect -25449 25175 -25369 25482
rect -38182 23503 -34852 23605
rect -38168 18987 -34861 19065
rect -40596 17394 -40360 17630
rect -38174 15987 -34852 16075
rect -25452 24714 -25365 24945
rect -15727 25018 -15632 25447
rect -17635 24874 -17507 25002
rect -13989 25600 -13925 25664
rect -12384 25604 -12321 25823
rect -14410 24808 -14346 24872
rect -17635 23645 -17507 23773
rect -15725 23405 -15658 23637
rect -12393 24458 -12328 24712
rect -12398 24003 -12316 24239
rect -12389 22857 -12319 23277
rect -12391 22399 -12323 22624
rect -25452 17627 -25387 17922
rect -25450 17169 -25378 17404
rect -24170 16185 -24106 16249
rect -27920 15377 -27856 15441
rect -25517 14157 -25444 14446
rect -25518 13690 -25446 13925
rect -18223 14009 -18159 14073
rect 4328 28531 4392 28595
rect 8338 28528 8402 28592
rect -5279 27468 -5215 27532
rect -3918 26791 -3854 26855
rect 19871 25945 19935 26009
rect 19873 25534 19937 25598
rect 5715 24186 5783 24594
rect 7068 24528 7132 24592
rect 42856 24065 46190 24174
rect 36066 23954 36130 24018
rect 35152 23802 35216 23866
rect 7091 23588 7155 23652
rect 37819 23492 37892 23611
rect 39346 23493 39420 23714
rect 8787 23246 8943 23356
rect 2550 22999 2614 23063
rect 10202 22999 10266 23063
rect 37819 22946 37905 23194
rect 39335 22952 39421 23200
rect 35100 22610 35280 22790
rect 35760 22668 36021 22730
rect 47556 22498 47792 22734
rect 37826 22151 37896 22280
rect 39346 22167 39420 22388
rect -971 21561 -907 21625
rect 6307 21561 6371 21625
rect 6310 20893 6374 20957
rect -971 20651 -907 20715
rect -12355 17904 -12291 17968
rect -13064 14077 -13000 14141
rect -13941 10117 -13877 10181
rect 51 19449 115 19513
rect -756 19148 -692 19212
rect 3061 19042 3125 19106
rect 4857 19027 5194 19173
rect 7085 19042 7149 19106
rect 8981 19042 9045 19106
rect 10232 18994 10296 19058
rect 5707 18846 5771 18910
rect 7706 18846 7770 18910
rect 4899 18587 4963 18651
rect 6897 18587 6961 18651
rect 8280 18654 8344 18718
rect 13574 18624 13638 18688
rect 3707 18248 3771 18312
rect 9706 18248 9770 18312
rect 37814 21621 37899 21823
rect 35152 21521 35216 21585
rect 39341 21586 39427 21834
rect 35477 21315 35541 21379
rect 42854 21069 46188 21178
rect 14688 20963 14752 21027
rect 14686 19214 14750 19278
rect 23689 19318 23753 19382
rect 20971 18998 21035 19062
rect 2898 17967 2962 18031
rect 8899 17967 8963 18031
rect 233 17708 297 17772
rect -821 17461 -757 17525
rect 14689 17485 14753 17549
rect 23689 17488 23753 17552
rect -10416 17093 -10352 17157
rect 4295 17225 4359 17289
rect 6227 17225 6291 17289
rect 13603 17019 13667 17083
rect -10415 16224 -10351 16288
rect 251 16238 11139 16446
rect -5786 15644 -5722 15708
rect -3008 15390 -2944 15454
rect -4902 14236 -4832 14446
rect -4917 13706 -4833 13998
rect -6162 10758 -5937 10833
rect -10970 10159 -10906 10223
rect -5707 10751 -5401 10838
rect -6156 10140 -6092 10204
rect -6167 9513 -5929 9592
rect -3144 14719 -3061 14998
rect -3023 14580 -2959 14644
rect -2598 13073 -2534 13137
rect -1808 12726 -1725 13133
rect -5361 10140 -5297 10204
rect -4789 10169 -4725 10233
rect -4448 10169 -4384 10233
rect -5708 9509 -5399 9595
rect -7214 7003 -6751 7243
rect -25521 6408 -25446 6669
rect -18251 6239 -18187 6303
rect -13075 6249 -13011 6313
rect -4917 6392 -4836 6695
rect -25522 5929 -25447 6174
rect -4907 5950 -4841 6163
rect -1498 12345 -1434 12409
rect -2885 12264 -2821 12328
rect -1926 11471 -1862 11535
rect -1759 11140 -1693 11529
rect -2212 10665 -2148 10729
rect -1498 10719 -1434 10783
rect -1926 9873 -1862 9937
rect -1759 9532 -1695 9930
rect -2212 9065 -2148 9129
rect -1498 9061 -1434 9125
rect -2598 8271 -2534 8335
rect -1758 7930 -1690 8330
rect -2885 7463 -2821 7527
rect -1498 7522 -1434 7586
rect -1498 6974 -1434 7258
rect -1498 6387 -1434 6451
rect -3050 5978 -2986 6042
rect -3193 5296 -3110 5577
rect -3028 5169 -2964 5233
rect -10766 4983 -10702 5047
rect 28 10640 187 16189
rect 5478 14421 5656 14599
rect 11239 14426 11399 16184
rect 14685 15689 14749 15753
rect 23686 15724 23750 15788
rect 20928 15432 20992 15496
rect 14690 15164 14754 15228
rect 11257 12990 11384 13954
rect 14685 13901 14749 13965
rect 23686 13933 23750 13997
rect 13636 13464 13700 13528
rect 4630 11802 4808 11980
rect 11243 11316 11398 12129
rect 14702 12116 14766 12180
rect 23691 12126 23755 12190
rect 20985 11842 21049 11906
rect 13699 11612 13763 11676
rect 6483 10356 11218 10537
rect 14691 10319 14755 10383
rect 23691 10316 23755 10380
rect 372 10003 1812 10144
rect 5727 9990 11722 10135
rect 13876 9993 21118 10150
rect 29 5570 212 9830
rect 4679 8188 4857 8366
rect 17646 8273 17824 8451
rect 35489 8467 35553 8531
rect 36066 9090 36130 9154
rect 36631 8405 36695 8469
rect 35024 8219 35088 8283
rect 38575 7892 38645 8038
rect 40100 7933 40181 8121
rect 36301 7814 36532 7881
rect 4679 6188 4857 6366
rect 13350 6313 13528 6491
rect 17646 6273 17824 6451
rect 16101 4910 16279 5088
rect 19101 4910 19279 5088
rect 21250 4540 21417 7514
rect 38568 7375 38649 7563
rect 40087 7388 40168 7576
rect 36362 7275 36531 7337
rect 35028 7159 35092 7223
rect 42602 7143 45923 7232
rect 35027 6890 35091 6954
rect 36352 6721 36437 6795
rect 38571 6582 38649 6707
rect 40092 6597 40173 6785
rect 36971 6169 37067 6265
rect 38563 6044 38644 6232
rect 40092 6041 40173 6229
rect 35027 5821 35091 5885
rect 35970 5644 36149 5707
rect 35024 5498 35088 5562
rect 47473 5564 47709 5800
rect 38574 5187 38648 5322
rect 40109 5217 40190 5405
rect 36514 5092 36734 5162
rect 38562 4691 38643 4879
rect 40092 4669 40173 4857
rect 36364 4555 36509 4613
rect 35035 4428 35099 4492
rect 4679 4188 4857 4366
rect 35024 4123 35088 4187
rect 42599 4144 45959 4233
rect 36972 3993 37068 4089
rect 38572 3781 38651 3934
rect 40099 3838 40180 4026
rect 36359 3459 36486 3531
rect 38565 3291 38646 3479
rect 40089 3285 40170 3473
rect 35031 3058 35095 3122
rect 28 359 190 2773
rect 12207 2595 12385 2773
rect 4679 2188 4857 2366
rect 21243 1288 21419 2139
rect 35489 1527 35553 1591
rect 36066 2150 36130 2214
rect 36631 1465 36695 1529
rect 35024 1279 35088 1343
rect 38575 952 38645 1098
rect 40100 993 40181 1181
rect 36301 874 36532 941
rect 38568 435 38649 623
rect 40087 448 40168 636
rect 36362 335 36531 397
rect 322 67 21107 232
rect 35028 219 35092 283
rect 42599 199 45930 309
rect 35027 -50 35091 14
rect 36352 -219 36437 -145
rect 38571 -358 38649 -233
rect 40092 -343 40173 -155
rect 36971 -771 37067 -675
rect 38563 -896 38644 -708
rect 40092 -899 40173 -711
rect 35027 -1119 35091 -1055
rect 35970 -1296 36149 -1233
rect 35024 -1442 35088 -1378
rect 47489 -1376 47725 -1140
rect 38574 -1753 38648 -1618
rect 40109 -1723 40190 -1535
rect 36514 -1848 36734 -1778
rect 38562 -2249 38643 -2061
rect 40092 -2271 40173 -2083
rect 36364 -2385 36509 -2327
rect 35035 -2512 35099 -2448
rect 35024 -2817 35088 -2753
rect 42587 -2796 45933 -2708
rect 36972 -2947 37068 -2851
rect 38572 -3159 38651 -3006
rect 40099 -3102 40180 -2914
rect 36359 -3481 36486 -3409
rect 38565 -3649 38646 -3461
rect 40089 -3655 40170 -3467
rect 35031 -3882 35095 -3818
rect -3595 -10130 -3503 -6822
rect -600 -10140 -486 -6825
rect -2179 -12318 -1943 -12082
<< metal3 >>
rect -17013 85607 -16777 90441
rect -17013 85371 -15174 85607
rect -15410 78145 -15174 85371
rect 10990 85579 11226 90441
rect 22915 85752 23151 90441
rect 10990 85343 12843 85579
rect 22915 85516 24892 85752
rect -15420 78140 -15164 78145
rect -15420 77904 -15410 78140
rect -15174 77904 -15164 78140
rect 12607 78116 12843 85343
rect 24656 78117 24892 85516
rect -15420 77899 -15164 77904
rect 12596 78111 12852 78116
rect 12596 77875 12606 78111
rect 12842 77875 12852 78111
rect 12596 77870 12852 77875
rect 24646 78112 24902 78117
rect 24646 77876 24656 78112
rect 24892 77876 24902 78112
rect 24646 77871 24902 77876
rect 14134 76745 14282 76750
rect -13858 76729 -13737 76734
rect -16859 76723 -16738 76728
rect -16859 73398 -16849 76723
rect -16748 73398 -16738 76723
rect -13858 73404 -13848 76729
rect -13747 73404 -13737 76729
rect -13858 73399 -13737 73404
rect 11133 76732 11281 76737
rect -16859 73393 -16738 73398
rect 11133 73392 11143 76732
rect 11271 73392 11281 76732
rect 14134 73405 14144 76745
rect 14272 73405 14282 76745
rect 14134 73400 14282 73405
rect 57721 75975 62907 76211
rect 11133 73387 11281 73392
rect -16697 71802 -16560 71832
rect -16697 71738 -16664 71802
rect -16600 71738 -16560 71802
rect -16697 71706 -16560 71738
rect -15509 71798 -15392 71820
rect -15509 71734 -15486 71798
rect -15422 71734 -15392 71798
rect -15509 71709 -15392 71734
rect -15292 71805 -15176 71835
rect -15292 71741 -15269 71805
rect -15205 71741 -15176 71805
rect -15292 71714 -15176 71741
rect -14161 71802 -14041 71826
rect -14161 71738 -14135 71802
rect -14071 71738 -14041 71802
rect -14161 71709 -14041 71738
rect -16577 70298 -16469 70319
rect -16577 70234 -16554 70298
rect -16490 70234 -16469 70298
rect -16577 70206 -16469 70234
rect -15464 70284 -15355 70304
rect -15464 70220 -15440 70284
rect -15376 70220 -15355 70284
rect -15464 70197 -15355 70220
rect -15249 70285 -15140 70310
rect -15249 70221 -15227 70285
rect -15163 70221 -15140 70285
rect -15249 70197 -15140 70221
rect -14091 70285 -13954 70311
rect -14091 70221 -14063 70285
rect -13999 70221 -13954 70285
rect -14091 70197 -13954 70221
rect 57721 69420 57957 75975
rect 36555 69334 57957 69420
rect 36555 69270 36631 69334
rect 36695 69270 57957 69334
rect 36555 69184 57957 69270
rect -13963 68742 62907 68813
rect -16718 68703 -16634 68708
rect -13963 68703 36065 68742
rect -16718 68639 -16708 68703
rect -16644 68676 36065 68703
rect 36131 68676 62907 68742
rect -16644 68639 62907 68676
rect -16718 68634 -16634 68639
rect -13963 68577 62907 68639
rect -15432 68515 -15348 68520
rect -15973 68261 -15880 68266
rect -15973 68105 -15963 68261
rect -15890 68105 -15880 68261
rect -15432 68166 -15422 68515
rect -15358 68166 -15348 68515
rect -15432 68161 -15348 68166
rect -14889 68264 -14796 68269
rect -15973 68100 -15880 68105
rect -14889 68108 -14879 68264
rect -14806 68108 -14796 68264
rect -14889 68103 -14796 68108
rect -13966 68082 58032 68169
rect -14209 68073 -14125 68078
rect -13966 68073 35476 68082
rect -14209 68009 -14199 68073
rect -14135 68016 35476 68073
rect 35542 68016 58032 68082
rect -14135 68009 58032 68016
rect -14209 68004 -14125 68009
rect -13966 67933 58032 68009
rect -16605 67613 -16482 67643
rect -16605 67549 -16577 67613
rect -16513 67549 -16482 67613
rect -16605 67518 -16482 67549
rect -15449 67607 -15330 67633
rect -15449 67543 -15422 67607
rect -15358 67543 -15330 67607
rect -15449 67513 -15330 67543
rect -14328 67618 -14211 67641
rect -14328 67554 -14304 67618
rect -14240 67554 -14211 67618
rect -14328 67526 -14211 67554
rect -13106 66705 -13096 66769
rect -13032 66705 -8073 66769
rect -8009 66705 -7999 66769
rect -12325 66382 -12315 66446
rect -12251 66382 -7266 66446
rect -7202 66382 -7192 66446
rect -11313 65949 -11305 66013
rect -11241 65949 -2673 66013
rect -2609 65949 -2599 66013
rect -10544 65696 -10536 65760
rect -10472 65696 -1866 65760
rect -1802 65696 -1792 65760
rect -8083 65265 -8073 65329
rect -8009 65265 -7999 65329
rect -2683 65265 -2673 65329
rect -2609 65265 -2599 65329
rect -7276 65012 -7266 65076
rect -7202 65012 -7192 65076
rect -1876 65012 -1866 65076
rect -1802 65012 -1792 65076
rect 17420 64743 17506 64748
rect 17420 64169 17430 64743
rect 17496 64169 17506 64743
rect 17420 64164 17506 64169
rect 23948 64743 24034 64748
rect 23948 64169 23958 64743
rect 24024 64169 24034 64743
rect 23948 64164 24034 64169
rect 31564 64743 31650 64748
rect 31564 64169 31574 64743
rect 31640 64169 31650 64743
rect 31564 64164 31650 64169
rect -11081 63205 -11071 63557
rect -10737 63402 -10727 63557
rect -9894 63402 -9432 63407
rect -10737 63338 -10187 63402
rect -10123 63338 -10113 63402
rect -9894 63338 -9884 63402
rect -9442 63338 -9432 63402
rect -10737 63205 -10727 63338
rect -9894 63333 -9432 63338
rect -8083 63404 -7621 63409
rect -8083 63340 -8073 63404
rect -7631 63340 -7621 63404
rect -8083 63335 -7621 63340
rect -6288 63400 -5826 63405
rect -6288 63336 -6278 63400
rect -5836 63336 -5826 63400
rect -6288 63331 -5826 63336
rect -4489 63398 -4027 63403
rect -4489 63334 -4479 63398
rect -4037 63334 -4027 63398
rect -4489 63329 -4027 63334
rect -2698 63402 -2236 63407
rect -2698 63338 -2688 63402
rect -2246 63338 -2236 63402
rect -2698 63333 -2236 63338
rect -896 63398 -434 63403
rect -896 63334 -886 63398
rect -444 63334 -434 63398
rect -896 63329 -434 63334
rect 747 63232 1297 63237
rect -6949 63206 -6689 63211
rect -6949 62966 -6939 63206
rect -6699 62966 -6689 63206
rect 747 62992 757 63232
rect 1287 62992 1297 63232
rect 747 62987 1297 62992
rect -6949 62961 -6689 62966
rect 17965 62740 18051 62745
rect 17965 62166 17975 62740
rect 18041 62166 18051 62740
rect 17965 62161 18051 62166
rect 19053 62740 19139 62745
rect 19053 62166 19063 62740
rect 19129 62166 19139 62740
rect 19053 62161 19139 62166
rect 21229 62740 21315 62745
rect 21229 62166 21239 62740
rect 21305 62166 21315 62740
rect 21229 62161 21315 62166
rect 22317 62740 22403 62745
rect 22317 62166 22327 62740
rect 22393 62166 22403 62740
rect 22317 62161 22403 62166
rect 23405 62740 23491 62745
rect 23405 62166 23415 62740
rect 23481 62166 23491 62740
rect 23405 62161 23491 62166
rect 24493 62740 24579 62745
rect 24493 62166 24503 62740
rect 24569 62166 24579 62740
rect 24493 62161 24579 62166
rect 25581 62740 25667 62745
rect 25581 62166 25591 62740
rect 25657 62166 25667 62740
rect 25581 62161 25667 62166
rect 26669 62740 26755 62745
rect 26669 62166 26679 62740
rect 26745 62166 26755 62740
rect 26669 62161 26755 62166
rect 28845 62740 28931 62745
rect 28845 62166 28855 62740
rect 28921 62166 28931 62740
rect 28845 62161 28931 62166
rect 29933 62740 30019 62745
rect 29933 62166 29943 62740
rect 30009 62166 30019 62740
rect 29933 62161 30019 62166
rect 31021 62740 31107 62745
rect 31021 62166 31031 62740
rect 31097 62166 31107 62740
rect 31021 62161 31107 62166
rect 57796 61375 58032 67933
rect 57796 61139 62907 61375
rect 10167 60836 10561 60841
rect 337 60827 529 60832
rect -8583 54595 -8471 54619
rect -8583 54531 -8557 54595
rect -8493 54531 -8471 54595
rect -8583 54507 -8471 54531
rect -6889 54596 -6772 54625
rect -6889 54532 -6866 54596
rect -6802 54532 -6772 54596
rect -6889 54508 -6772 54532
rect -5179 54595 -5082 54614
rect -5179 54531 -5161 54595
rect -5097 54531 -5082 54595
rect -5179 54511 -5082 54531
rect -3385 54595 -3280 54622
rect -3385 54531 -3365 54595
rect -3301 54531 -3280 54595
rect -3385 54512 -3280 54531
rect -1556 54595 -1453 54615
rect -1556 54531 -1536 54595
rect -1472 54531 -1453 54595
rect -1556 54511 -1453 54531
rect -9714 54403 -9452 54408
rect -9714 54339 -9704 54403
rect -9462 54339 -9452 54403
rect -9714 54334 -9452 54339
rect -7919 54402 -7657 54407
rect -7919 54338 -7909 54402
rect -7667 54338 -7657 54402
rect -7919 54333 -7657 54338
rect -6119 54404 -5857 54409
rect -6119 54340 -6109 54404
rect -5867 54340 -5857 54404
rect -6119 54335 -5857 54340
rect -4321 54403 -4059 54408
rect -4321 54339 -4311 54403
rect -4069 54339 -4059 54403
rect -4321 54334 -4059 54339
rect -2523 54404 -2261 54409
rect -2523 54340 -2513 54404
rect -2271 54340 -2261 54404
rect -2523 54335 -2261 54340
rect -720 54403 -458 54408
rect -720 54339 -710 54403
rect -468 54339 -458 54403
rect -720 54334 -458 54339
rect 156 54404 258 54424
rect 156 54340 176 54404
rect 240 54340 258 54404
rect 156 54319 258 54340
rect -7275 54019 -7265 54083
rect -7201 54019 -7191 54083
rect -1875 54019 -1865 54083
rect -1801 54019 -1791 54083
rect -8083 53766 -8073 53830
rect -8009 53766 -7999 53830
rect -2683 53766 -2673 53830
rect -2609 53766 -2599 53830
rect -10546 53338 -10536 53402
rect -10472 53338 -1865 53402
rect -1801 53338 -1791 53402
rect -11315 53082 -11305 53146
rect -11241 53082 -2673 53146
rect -2609 53082 -2599 53146
rect 337 53121 347 60827
rect 519 53121 529 60827
rect 5400 58930 5598 58935
rect 5400 58752 5410 58930
rect 5588 58752 5598 58930
rect 5400 58747 5598 58752
rect 2037 57475 2235 57480
rect 2037 57297 2047 57475
rect 2225 57297 2235 57475
rect 2037 57292 2235 57297
rect 4037 57475 4235 57480
rect 4037 57297 4047 57475
rect 4225 57297 4235 57475
rect 4037 57292 4235 57297
rect 5400 55930 5598 55935
rect 5400 55752 5410 55930
rect 5588 55752 5598 55930
rect 5400 55747 5598 55752
rect 337 53116 529 53121
rect 3997 53179 4195 53184
rect 3997 53001 4007 53179
rect 4185 53001 4195 53179
rect 3997 52996 4195 53001
rect -12325 52649 -12315 52713
rect -12251 52649 -7265 52713
rect -7201 52649 -7191 52713
rect -13106 52326 -13096 52390
rect -13032 52326 -8073 52390
rect -8009 52326 -7999 52390
rect 7715 52036 7913 52041
rect 7715 51858 7725 52036
rect 7903 51858 7913 52036
rect 7715 51853 7913 51858
rect -8864 51249 -8760 51254
rect -8864 51014 -8854 51249
rect -8770 51014 -8760 51249
rect -7742 51247 -7634 51272
rect -7742 51183 -7722 51247
rect -7658 51183 -7634 51247
rect -7742 51162 -7634 51183
rect -3372 51074 -2526 51079
rect -8864 51009 -8760 51014
rect -5698 51066 -3878 51071
rect -5698 50883 -5688 51066
rect -3888 50883 -3878 51066
rect -3372 50896 -3362 51074
rect -2536 50896 -2526 51074
rect -3372 50891 -2526 50896
rect -1665 51064 -755 51069
rect -5698 50878 -3878 50883
rect -1665 50886 -1655 51064
rect -765 50886 -755 51064
rect -1665 50881 -755 50886
rect -8884 50791 -8770 50796
rect -8884 50617 -8874 50791
rect -19102 50512 -8874 50617
rect -8884 50378 -8874 50512
rect -8780 50378 -8770 50791
rect -88 50774 131 50779
rect -5942 50720 -5738 50725
rect -8884 50373 -8770 50378
rect -8497 50441 -8398 50461
rect -8497 50377 -8480 50441
rect -8416 50377 -8398 50441
rect -8497 50357 -8398 50377
rect -57094 50072 -28000 50155
rect -57094 50008 -8480 50072
rect -8416 50008 -8406 50072
rect -57094 49919 -28000 50008
rect -27080 49720 -26716 49725
rect -27080 49656 -27070 49720
rect -26726 49656 -26716 49720
rect -27080 49651 -26716 49656
rect -26472 49418 -26408 50008
rect -26070 49424 -25986 49429
rect -26472 49413 -26147 49418
rect -26472 49349 -26408 49413
rect -26157 49349 -26147 49413
rect -26070 49360 -26060 49424
rect -25996 49360 -7722 49424
rect -7658 49360 -7648 49424
rect -26070 49355 -25986 49360
rect -26418 49344 -26147 49349
rect -25994 49178 -25630 49183
rect -25994 49114 -25984 49178
rect -25640 49114 -25630 49178
rect -25994 49109 -25630 49114
rect -5942 47776 -5932 50720
rect -5748 47776 -5738 50720
rect -5942 47771 -5738 47776
rect -88 47752 -78 50774
rect 121 47752 131 50774
rect -88 47747 131 47752
rect 10167 47617 10177 60836
rect 10551 47617 10561 60836
rect 17420 60743 17506 60748
rect 17420 60169 17430 60743
rect 17496 60169 17506 60743
rect 17420 60164 17506 60169
rect 18508 60743 18594 60748
rect 18508 60169 18518 60743
rect 18584 60169 18594 60743
rect 18508 60164 18594 60169
rect 19596 60743 19682 60748
rect 19596 60169 19606 60743
rect 19672 60169 19682 60743
rect 19596 60164 19682 60169
rect 20684 60743 20770 60748
rect 20684 60169 20694 60743
rect 20760 60169 20770 60743
rect 20684 60164 20770 60169
rect 21772 60743 21858 60748
rect 21772 60169 21782 60743
rect 21848 60169 21858 60743
rect 21772 60164 21858 60169
rect 22860 60743 22946 60748
rect 22860 60169 22870 60743
rect 22936 60169 22946 60743
rect 22860 60164 22946 60169
rect 23948 60743 24034 60748
rect 23948 60169 23958 60743
rect 24024 60169 24034 60743
rect 23948 60164 24034 60169
rect 25036 60743 25122 60748
rect 25036 60169 25046 60743
rect 25112 60169 25122 60743
rect 25036 60164 25122 60169
rect 26124 60743 26210 60748
rect 26124 60169 26134 60743
rect 26200 60169 26210 60743
rect 26124 60164 26210 60169
rect 27212 60743 27298 60748
rect 27212 60169 27222 60743
rect 27288 60169 27298 60743
rect 27212 60164 27298 60169
rect 28300 60743 28386 60748
rect 28300 60169 28310 60743
rect 28376 60169 28386 60743
rect 28300 60164 28386 60169
rect 29388 60743 29474 60748
rect 29388 60169 29398 60743
rect 29464 60169 29474 60743
rect 29388 60164 29474 60169
rect 30476 60743 30562 60748
rect 30476 60169 30486 60743
rect 30552 60169 30562 60743
rect 30476 60164 30562 60169
rect 31564 60743 31650 60748
rect 31564 60169 31574 60743
rect 31640 60169 31650 60743
rect 31564 60164 31650 60169
rect 17965 58740 18051 58745
rect 17965 58166 17975 58740
rect 18041 58166 18051 58740
rect 17965 58161 18051 58166
rect 19053 58740 19139 58745
rect 19053 58166 19063 58740
rect 19129 58166 19139 58740
rect 19053 58161 19139 58166
rect 20141 58740 20227 58745
rect 20141 58166 20151 58740
rect 20217 58166 20227 58740
rect 20141 58161 20227 58166
rect 21229 58740 21315 58745
rect 21229 58166 21239 58740
rect 21305 58166 21315 58740
rect 21229 58161 21315 58166
rect 22317 58740 22403 58745
rect 22317 58166 22327 58740
rect 22393 58166 22403 58740
rect 22317 58161 22403 58166
rect 23405 58740 23491 58745
rect 23405 58166 23415 58740
rect 23481 58166 23491 58740
rect 23405 58161 23491 58166
rect 24493 58740 24579 58745
rect 24493 58166 24503 58740
rect 24569 58166 24579 58740
rect 24493 58161 24579 58166
rect 25581 58740 25667 58745
rect 25581 58166 25591 58740
rect 25657 58166 25667 58740
rect 25581 58161 25667 58166
rect 26669 58740 26755 58745
rect 26669 58166 26679 58740
rect 26745 58166 26755 58740
rect 26669 58161 26755 58166
rect 27757 58740 27843 58745
rect 27757 58166 27767 58740
rect 27833 58166 27843 58740
rect 27757 58161 27843 58166
rect 28845 58740 28931 58745
rect 28845 58166 28855 58740
rect 28921 58166 28931 58740
rect 28845 58161 28931 58166
rect 29933 58740 30019 58745
rect 29933 58166 29943 58740
rect 30009 58166 30019 58740
rect 29933 58161 30019 58166
rect 31021 58740 31107 58745
rect 31021 58166 31031 58740
rect 31097 58166 31107 58740
rect 31021 58161 31107 58166
rect 17420 56743 17506 56748
rect 17420 56169 17430 56743
rect 17496 56169 17506 56743
rect 17420 56164 17506 56169
rect 18508 56743 18594 56748
rect 18508 56169 18518 56743
rect 18584 56169 18594 56743
rect 18508 56164 18594 56169
rect 19596 56743 19682 56748
rect 19596 56169 19606 56743
rect 19672 56169 19682 56743
rect 19596 56164 19682 56169
rect 20684 56743 20770 56748
rect 20684 56169 20694 56743
rect 20760 56169 20770 56743
rect 20684 56164 20770 56169
rect 21772 56743 21858 56748
rect 21772 56169 21782 56743
rect 21848 56169 21858 56743
rect 21772 56164 21858 56169
rect 22860 56743 22946 56748
rect 22860 56169 22870 56743
rect 22936 56169 22946 56743
rect 22860 56164 22946 56169
rect 23948 56743 24034 56748
rect 23948 56169 23958 56743
rect 24024 56169 24034 56743
rect 23948 56164 24034 56169
rect 25036 56743 25122 56748
rect 25036 56169 25046 56743
rect 25112 56169 25122 56743
rect 25036 56164 25122 56169
rect 26124 56743 26210 56748
rect 26124 56169 26134 56743
rect 26200 56169 26210 56743
rect 26124 56164 26210 56169
rect 27212 56743 27298 56748
rect 27212 56169 27222 56743
rect 27288 56169 27298 56743
rect 27212 56164 27298 56169
rect 28300 56743 28386 56748
rect 28300 56169 28310 56743
rect 28376 56169 28386 56743
rect 28300 56164 28386 56169
rect 29388 56743 29474 56748
rect 29388 56169 29398 56743
rect 29464 56169 29474 56743
rect 29388 56164 29474 56169
rect 30476 56743 30562 56748
rect 30476 56169 30486 56743
rect 30552 56169 30562 56743
rect 30476 56164 30562 56169
rect 31564 56743 31650 56748
rect 31564 56169 31574 56743
rect 31640 56169 31650 56743
rect 31564 56164 31650 56169
rect 52756 55101 62907 55337
rect 17965 54740 18051 54745
rect 17965 54166 17975 54740
rect 18041 54166 18051 54740
rect 17965 54161 18051 54166
rect 19053 54740 19139 54745
rect 19053 54166 19063 54740
rect 19129 54166 19139 54740
rect 19053 54161 19139 54166
rect 20141 54740 20227 54745
rect 20141 54166 20151 54740
rect 20217 54166 20227 54740
rect 20141 54161 20227 54166
rect 21229 54740 21315 54745
rect 21229 54166 21239 54740
rect 21305 54166 21315 54740
rect 21229 54161 21315 54166
rect 22317 54740 22403 54745
rect 22317 54166 22327 54740
rect 22393 54166 22403 54740
rect 22317 54161 22403 54166
rect 23405 54740 23491 54745
rect 23405 54166 23415 54740
rect 23481 54166 23491 54740
rect 23405 54161 23491 54166
rect 24493 54740 24579 54745
rect 24493 54166 24503 54740
rect 24569 54166 24579 54740
rect 24493 54161 24579 54166
rect 25581 54740 25667 54745
rect 25581 54166 25591 54740
rect 25657 54166 25667 54740
rect 25581 54161 25667 54166
rect 26669 54740 26755 54745
rect 26669 54166 26679 54740
rect 26745 54166 26755 54740
rect 26669 54161 26755 54166
rect 27757 54740 27843 54745
rect 27757 54166 27767 54740
rect 27833 54166 27843 54740
rect 27757 54161 27843 54166
rect 28845 54740 28931 54745
rect 28845 54166 28855 54740
rect 28921 54166 28931 54740
rect 28845 54161 28931 54166
rect 29933 54740 30019 54745
rect 29933 54166 29943 54740
rect 30009 54166 30019 54740
rect 29933 54161 30019 54166
rect 31021 54740 31107 54745
rect 31021 54166 31031 54740
rect 31097 54166 31107 54740
rect 31021 54161 31107 54166
rect 17420 52743 17506 52748
rect 17420 52169 17430 52743
rect 17496 52169 17506 52743
rect 17420 52164 17506 52169
rect 18508 52743 18594 52748
rect 18508 52169 18518 52743
rect 18584 52169 18594 52743
rect 18508 52164 18594 52169
rect 19596 52743 19682 52748
rect 19596 52169 19606 52743
rect 19672 52169 19682 52743
rect 19596 52164 19682 52169
rect 20684 52743 20770 52748
rect 20684 52169 20694 52743
rect 20760 52169 20770 52743
rect 20684 52164 20770 52169
rect 21772 52743 21858 52748
rect 21772 52169 21782 52743
rect 21848 52169 21858 52743
rect 21772 52164 21858 52169
rect 22860 52743 22946 52748
rect 22860 52169 22870 52743
rect 22936 52169 22946 52743
rect 22860 52164 22946 52169
rect 23948 52743 24034 52748
rect 23948 52169 23958 52743
rect 24024 52169 24034 52743
rect 23948 52164 24034 52169
rect 25036 52743 25122 52748
rect 25036 52169 25046 52743
rect 25112 52169 25122 52743
rect 25036 52164 25122 52169
rect 26124 52743 26210 52748
rect 26124 52169 26134 52743
rect 26200 52169 26210 52743
rect 26124 52164 26210 52169
rect 27212 52743 27298 52748
rect 27212 52169 27222 52743
rect 27288 52169 27298 52743
rect 27212 52164 27298 52169
rect 28300 52743 28386 52748
rect 28300 52169 28310 52743
rect 28376 52169 28386 52743
rect 28300 52164 28386 52169
rect 29388 52743 29474 52748
rect 29388 52169 29398 52743
rect 29464 52169 29474 52743
rect 29388 52164 29474 52169
rect 30476 52743 30562 52748
rect 30476 52169 30486 52743
rect 30552 52169 30562 52743
rect 30476 52164 30562 52169
rect 31564 52743 31650 52748
rect 31564 52169 31574 52743
rect 31640 52169 31650 52743
rect 31564 52164 31650 52169
rect 17965 50740 18051 50745
rect 17965 50166 17975 50740
rect 18041 50166 18051 50740
rect 17965 50161 18051 50166
rect 20141 50740 20227 50745
rect 20141 50166 20151 50740
rect 20217 50166 20227 50740
rect 20141 50161 20227 50166
rect 21229 50740 21315 50745
rect 21229 50166 21239 50740
rect 21305 50166 21315 50740
rect 21229 50161 21315 50166
rect 23405 50740 23491 50745
rect 23405 50166 23415 50740
rect 23481 50166 23491 50740
rect 23405 50161 23491 50166
rect 24493 50740 24579 50745
rect 24493 50166 24503 50740
rect 24569 50166 24579 50740
rect 24493 50161 24579 50166
rect 25581 50740 25667 50745
rect 25581 50166 25591 50740
rect 25657 50166 25667 50740
rect 25581 50161 25667 50166
rect 27757 50740 27843 50745
rect 27757 50166 27767 50740
rect 27833 50166 27843 50740
rect 27757 50161 27843 50166
rect 28845 50740 28931 50745
rect 28845 50166 28855 50740
rect 28921 50166 28931 50740
rect 28845 50161 28931 50166
rect 31021 50740 31107 50745
rect 31021 50166 31031 50740
rect 31097 50166 31107 50740
rect 31021 50161 31107 50166
rect 17420 48743 17506 48748
rect 17420 48169 17430 48743
rect 17496 48169 17506 48743
rect 17420 48164 17506 48169
rect 18508 48743 18594 48748
rect 18508 48169 18518 48743
rect 18584 48169 18594 48743
rect 18508 48164 18594 48169
rect 19596 48743 19682 48748
rect 19596 48169 19606 48743
rect 19672 48169 19682 48743
rect 19596 48164 19682 48169
rect 20684 48743 20770 48748
rect 20684 48169 20694 48743
rect 20760 48169 20770 48743
rect 20684 48164 20770 48169
rect 21772 48743 21858 48748
rect 21772 48169 21782 48743
rect 21848 48169 21858 48743
rect 21772 48164 21858 48169
rect 22860 48743 22946 48748
rect 22860 48169 22870 48743
rect 22936 48169 22946 48743
rect 22860 48164 22946 48169
rect 23948 48743 24034 48748
rect 23948 48169 23958 48743
rect 24024 48169 24034 48743
rect 23948 48164 24034 48169
rect 29388 48743 29474 48748
rect 29388 48169 29398 48743
rect 29464 48169 29474 48743
rect 29388 48164 29474 48169
rect 30476 48743 30562 48748
rect 30476 48169 30486 48743
rect 30552 48169 30562 48743
rect 30476 48164 30562 48169
rect 31564 48743 31650 48748
rect 31564 48169 31574 48743
rect 31640 48169 31650 48743
rect 31564 48164 31650 48169
rect 10167 47612 10561 47617
rect -23498 47192 -11361 47256
rect -11297 47192 -6411 47256
rect -6347 47192 -6337 47256
rect -27097 43313 -26980 43318
rect -27097 42779 -27087 43313
rect -26990 42779 -26980 43313
rect -27097 42774 -26980 42779
rect -27092 42169 -26985 42174
rect -27092 41002 -27082 42169
rect -26995 41002 -26985 42169
rect -27092 40997 -26985 41002
rect -27087 40643 -26980 40648
rect -27087 39476 -27077 40643
rect -26990 39476 -26980 40643
rect -27087 39471 -26980 39476
rect -31822 39166 -31738 39171
rect -31822 38827 -31812 39166
rect -31748 38827 -31738 39166
rect -31822 38822 -31738 38827
rect -27092 39120 -26988 39125
rect -31821 38613 -31737 38618
rect -31821 38141 -31811 38613
rect -31747 38141 -31737 38613
rect -29624 38413 -29140 38418
rect -29624 38349 -29614 38413
rect -29150 38349 -29140 38413
rect -29624 38344 -29140 38349
rect -27092 38232 -27082 39120
rect -26998 38232 -26988 39120
rect -27092 38227 -26988 38232
rect -31821 38136 -31737 38141
rect -23498 37802 -23434 47192
rect 17965 46740 18051 46745
rect -10497 46569 -10487 46633
rect -10423 46569 -6411 46633
rect -6347 46569 -6335 46633
rect -5934 46274 -5712 46279
rect -13479 43061 -13395 43066
rect -13479 42997 -13469 43061
rect -13405 42997 -9208 43061
rect -9144 42997 -9134 43061
rect -13479 42992 -13395 42997
rect -12703 42398 -12619 42403
rect -12703 42334 -12693 42398
rect -12629 42334 -10069 42398
rect -10005 42334 -9995 42398
rect -12703 42329 -12619 42334
rect -21501 42163 -21386 42190
rect -21501 42099 -21475 42163
rect -21411 42099 -21386 42163
rect -21501 42074 -21386 42099
rect -5934 39917 -5924 46274
rect -5967 39819 -5924 39917
rect -5722 39917 -5712 46274
rect 17965 46166 17975 46740
rect 18041 46166 18051 46740
rect 17965 46161 18051 46166
rect 19053 46740 19139 46745
rect 19053 46166 19063 46740
rect 19129 46166 19139 46740
rect 19053 46161 19139 46166
rect 20141 46740 20227 46745
rect 20141 46166 20151 46740
rect 20217 46166 20227 46740
rect 20141 46161 20227 46166
rect 21229 46740 21315 46745
rect 21229 46166 21239 46740
rect 21305 46166 21315 46740
rect 21229 46161 21315 46166
rect 22317 46740 22403 46745
rect 22317 46166 22327 46740
rect 22393 46166 22403 46740
rect 22317 46161 22403 46166
rect 24493 46740 24579 46745
rect 24493 46166 24503 46740
rect 24569 46166 24579 46740
rect 24493 46161 24579 46166
rect 25581 46740 25667 46745
rect 25581 46166 25591 46740
rect 25657 46166 25667 46740
rect 25581 46161 25667 46166
rect 26669 46740 26755 46745
rect 26669 46166 26679 46740
rect 26745 46166 26755 46740
rect 26669 46161 26755 46166
rect 27757 46740 27843 46745
rect 27757 46166 27767 46740
rect 27833 46166 27843 46740
rect 27757 46161 27843 46166
rect 28845 46740 28931 46745
rect 28845 46166 28855 46740
rect 28921 46166 28931 46740
rect 28845 46161 28931 46166
rect 29933 46740 30019 46745
rect 29933 46166 29943 46740
rect 30009 46166 30019 46740
rect 29933 46161 30019 46166
rect 31021 46740 31107 46745
rect 31021 46166 31031 46740
rect 31097 46166 31107 46740
rect 52756 46464 52992 55101
rect 40579 46375 40663 46380
rect 47769 46375 52992 46464
rect 40579 46311 40589 46375
rect 40653 46311 52992 46375
rect 40579 46306 40663 46311
rect 47769 46228 52992 46311
rect 55186 50886 62907 51122
rect 31021 46161 31107 46166
rect 10170 46128 10561 46133
rect 334 45844 568 45849
rect -4111 45307 -3913 45312
rect -4111 45129 -4101 45307
rect -3923 45129 -3913 45307
rect -4111 45124 -3913 45129
rect -1492 44459 -1294 44464
rect -1492 44281 -1482 44459
rect -1304 44281 -1294 44459
rect 334 44318 344 45844
rect 558 44318 568 45844
rect 2122 44508 2320 44513
rect 2122 44330 2132 44508
rect 2310 44330 2320 44508
rect 2122 44325 2320 44330
rect 4122 44508 4320 44513
rect 4122 44330 4132 44508
rect 4310 44330 4320 44508
rect 4122 44325 4320 44330
rect 6122 44508 6320 44513
rect 6122 44330 6132 44508
rect 6310 44330 6320 44508
rect 6122 44325 6320 44330
rect 8122 44508 8320 44513
rect 8122 44330 8132 44508
rect 8310 44330 8320 44508
rect 8122 44325 8320 44330
rect 334 44313 568 44318
rect -1492 44276 -1294 44281
rect 342 41383 522 41388
rect -5722 39851 -5651 39917
rect 342 39855 352 41383
rect 512 39855 522 41383
rect 10170 39867 10180 46128
rect 10551 39867 10561 46128
rect 55186 45902 55422 50886
rect 41136 45819 41220 45824
rect 47769 45819 55422 45902
rect 18221 45748 18339 45774
rect 18221 45684 18245 45748
rect 18309 45684 18339 45748
rect 18221 45659 18339 45684
rect 18766 45748 18884 45773
rect 18766 45684 18791 45748
rect 18855 45684 18884 45748
rect 18766 45658 18884 45684
rect 19308 45739 19426 45769
rect 19308 45675 19337 45739
rect 19401 45675 19426 45739
rect 19308 45654 19426 45675
rect 19856 45738 19974 45767
rect 19856 45674 19882 45738
rect 19946 45674 19974 45738
rect 19856 45652 19974 45674
rect 21487 45748 21605 45772
rect 21487 45684 21517 45748
rect 21581 45684 21605 45748
rect 21487 45657 21605 45684
rect 22023 45735 22141 45761
rect 22023 45671 22051 45735
rect 22115 45671 22141 45735
rect 22023 45646 22141 45671
rect 22573 45741 22691 45770
rect 22573 45677 22598 45741
rect 22662 45677 22691 45741
rect 22573 45655 22691 45677
rect 23116 45741 23234 45766
rect 23116 45677 23143 45741
rect 23207 45677 23234 45741
rect 23116 45651 23234 45677
rect 25837 45738 25955 45766
rect 25837 45674 25863 45738
rect 25927 45674 25955 45738
rect 25837 45651 25955 45674
rect 26381 45742 26499 45766
rect 26381 45678 26406 45742
rect 26470 45678 26499 45742
rect 26381 45651 26499 45678
rect 26920 45736 27038 45764
rect 26920 45672 26948 45736
rect 27012 45672 27038 45736
rect 26920 45649 27038 45672
rect 27479 45727 27597 45753
rect 27479 45663 27505 45727
rect 27569 45663 27597 45727
rect 27479 45638 27597 45663
rect 29103 45738 29221 45765
rect 29103 45674 29129 45738
rect 29193 45674 29221 45738
rect 29103 45650 29221 45674
rect 29645 45731 29763 45756
rect 29645 45667 29673 45731
rect 29737 45667 29763 45731
rect 29645 45641 29763 45667
rect 30198 45735 30316 45760
rect 30198 45671 30223 45735
rect 30287 45671 30316 45735
rect 30198 45645 30316 45671
rect 30728 45735 30846 45762
rect 41136 45755 41146 45819
rect 41210 45755 55422 45819
rect 41136 45750 41220 45755
rect 30728 45671 30756 45735
rect 30820 45671 30846 45735
rect 30728 45647 30846 45671
rect 47769 45666 55422 45755
rect 57721 47147 62907 47383
rect 44744 45074 45316 45079
rect 18762 45008 18791 45072
rect 18855 45008 39775 45072
rect 39711 44991 39775 45008
rect 44744 45007 44754 45074
rect 45306 45007 45316 45074
rect 44744 45002 45316 45007
rect 40978 44991 41062 44996
rect 39711 44927 40988 44991
rect 41052 44927 41062 44991
rect 40978 44922 41062 44927
rect 46284 44939 46540 44944
rect 57721 44939 57957 47147
rect 39547 44891 39631 44896
rect 25844 44827 25863 44891
rect 25927 44827 39557 44891
rect 39621 44827 39631 44891
rect 39547 44822 39631 44827
rect 39547 44701 39631 44706
rect 18231 44637 18245 44701
rect 18309 44637 39557 44701
rect 39621 44637 39631 44701
rect 46284 44703 46294 44939
rect 46530 44703 57957 44939
rect 46284 44698 46540 44703
rect 39547 44632 39631 44637
rect 40878 44607 40962 44612
rect 39711 44543 40888 44607
rect 40952 44543 40962 44607
rect 39711 44526 39775 44543
rect 40878 44538 40962 44543
rect 26392 44462 26406 44526
rect 26470 44462 39775 44526
rect 41506 44527 41884 44532
rect 41506 44462 41516 44527
rect 41874 44462 41884 44527
rect 41506 44457 41884 44462
rect 44756 43925 45303 43930
rect 22582 43858 22598 43922
rect 22662 43858 39775 43922
rect 39711 43841 39775 43858
rect 44756 43854 44766 43925
rect 45293 43854 45303 43925
rect 44756 43849 45303 43854
rect 40978 43841 41062 43846
rect 39711 43777 40988 43841
rect 41052 43777 41062 43841
rect 40978 43772 41062 43777
rect 46272 43788 46528 43793
rect 39547 43741 39631 43746
rect 30746 43677 30756 43741
rect 30820 43677 39557 43741
rect 39621 43677 39631 43741
rect 39547 43672 39631 43677
rect 39547 43551 39631 43556
rect 23126 43487 23143 43551
rect 23207 43487 39557 43551
rect 39621 43487 39631 43551
rect 46272 43552 46282 43788
rect 46518 43552 62907 43788
rect 46272 43547 46528 43552
rect 39547 43482 39631 43487
rect 40878 43457 40962 43462
rect 39711 43393 40888 43457
rect 40952 43393 40962 43457
rect 39711 43376 39775 43393
rect 40878 43388 40962 43393
rect 30214 43375 39775 43376
rect 30212 43311 30222 43375
rect 30286 43312 39775 43375
rect 41504 43377 41882 43382
rect 41504 43312 41514 43377
rect 41872 43312 41882 43377
rect 30286 43311 30296 43312
rect 41504 43307 41882 43312
rect 40579 42685 40663 42690
rect 47760 42685 57965 42777
rect 40579 42621 40589 42685
rect 40653 42621 57965 42685
rect 40579 42616 40663 42621
rect 47760 42541 57965 42621
rect 41136 42129 41220 42134
rect 47751 42129 55382 42223
rect 41136 42065 41146 42129
rect 41210 42065 55382 42129
rect 41136 42060 41220 42065
rect 47751 41987 55382 42065
rect 44746 41383 45293 41388
rect 19872 41318 19882 41382
rect 19946 41318 39775 41382
rect 39711 41301 39775 41318
rect 44746 41312 44756 41383
rect 45283 41312 45293 41383
rect 44746 41307 45293 41312
rect 40978 41301 41062 41306
rect 39711 41237 40988 41301
rect 41052 41237 41062 41301
rect 40978 41232 41062 41237
rect 46130 41256 46386 41261
rect 39547 41201 39631 41206
rect 26938 41137 26948 41201
rect 27012 41137 39557 41201
rect 39621 41137 39631 41201
rect 39547 41132 39631 41137
rect 46130 41020 46140 41256
rect 46376 41020 53037 41256
rect 39547 41011 39631 41016
rect 46130 41015 46386 41020
rect 19305 40947 19337 41011
rect 19401 40947 39557 41011
rect 39621 40947 39631 41011
rect 39547 40942 39631 40947
rect 40878 40917 40962 40922
rect 39711 40853 40888 40917
rect 40952 40853 40962 40917
rect 39711 40836 39775 40853
rect 40878 40848 40962 40853
rect 27490 40772 27505 40836
rect 27569 40772 39775 40836
rect 41422 40836 41800 40841
rect 41422 40771 41432 40836
rect 41790 40771 41800 40836
rect 41422 40766 41800 40771
rect 44746 40113 45293 40118
rect 21507 40048 21517 40112
rect 21581 40048 39775 40112
rect 39711 40031 39775 40048
rect 44746 40042 44756 40113
rect 45283 40042 45293 40113
rect 44746 40037 45293 40042
rect 40978 40031 41062 40036
rect 39711 39967 40988 40031
rect 41052 39967 41062 40031
rect 40978 39962 41062 39967
rect 46101 39966 46357 39971
rect 39547 39931 39631 39936
rect 29663 39867 29673 39931
rect 29737 39867 39557 39931
rect 39621 39867 39631 39931
rect 10170 39862 10561 39867
rect 39547 39862 39631 39867
rect -5722 39846 -138 39851
rect 342 39850 522 39855
rect -5722 39819 -5684 39846
rect -5967 39666 -5684 39819
rect -148 39666 -138 39846
rect 39547 39741 39631 39746
rect 22041 39677 22051 39741
rect 22115 39677 39557 39741
rect 39621 39677 39631 39741
rect 46101 39730 46111 39966
rect 46347 39730 50842 39966
rect 46101 39725 46357 39730
rect 39547 39672 39631 39677
rect -5967 39661 -138 39666
rect -5967 39650 -5651 39661
rect 40878 39647 40962 39652
rect 39711 39583 40888 39647
rect 40952 39583 40962 39647
rect 39711 39566 39775 39583
rect 40878 39578 40962 39583
rect -18893 39537 -18797 39542
rect -35528 37569 -35272 37573
rect -57094 37568 -35272 37569
rect -57094 37333 -35518 37568
rect -35528 37332 -35518 37333
rect -35282 37332 -35272 37568
rect -35528 37327 -35272 37332
rect -27089 37353 -26985 37358
rect -29662 37323 -29133 37328
rect -29662 37259 -29652 37323
rect -29143 37259 -29133 37323
rect -29662 37254 -29133 37259
rect -27089 36465 -27079 37353
rect -26995 36465 -26985 37353
rect -27089 36460 -26985 36465
rect -27087 36160 -26986 36165
rect -27087 34985 -27077 36160
rect -26996 34985 -26986 36160
rect -18893 36124 -18883 39537
rect -18807 36124 -18797 39537
rect 29119 39502 29129 39566
rect 29193 39502 39775 39566
rect 41420 39567 41798 39572
rect 41420 39502 41430 39567
rect 41788 39502 41798 39567
rect 41420 39497 41798 39502
rect 1473 38883 1537 38887
rect 1463 38878 1547 38883
rect 1463 38814 1473 38878
rect 1537 38814 1547 38878
rect 1463 38809 1547 38814
rect 2503 38881 2605 38886
rect -11723 38726 -11713 38790
rect -11649 38726 -4713 38790
rect -4649 38726 -4639 38790
rect -16012 37597 -15860 38546
rect -10912 38383 -10905 38447
rect -10841 38383 -4123 38447
rect -4059 38383 -4049 38447
rect 1473 37899 1537 38809
rect 2503 38642 2513 38881
rect 2595 38642 2605 38881
rect 2503 38637 2605 38642
rect 2505 38420 2624 38425
rect 1996 38074 2060 38083
rect 1986 38069 2070 38074
rect 1986 38005 1996 38069
rect 2060 38005 2070 38069
rect 1986 38000 2070 38005
rect -7732 37835 -7722 37899
rect -7658 37835 -2398 37899
rect -2334 37835 -760 37899
rect -696 37835 -686 37899
rect 1463 37835 1473 37899
rect 1537 37835 1547 37899
rect -8490 37307 -8480 37371
rect -8416 37307 -2815 37371
rect -2751 37370 -729 37371
rect -2751 37307 -760 37370
rect -770 37306 -760 37307
rect -696 37306 -686 37370
rect 1473 37134 1537 37835
rect 1996 37370 2060 38000
rect 2505 37996 2515 38420
rect 2614 37996 2624 38420
rect 13821 38372 13831 38436
rect 13895 38372 18245 38436
rect 18309 38372 18319 38436
rect 25853 38354 25863 38418
rect 25927 38354 32414 38418
rect 32478 38354 32488 38418
rect 2505 37991 2624 37996
rect 14576 37797 14586 37861
rect 14650 37797 18791 37861
rect 18855 37797 18865 37861
rect 26396 37774 26406 37838
rect 26470 37774 31824 37838
rect 31888 37774 31898 37838
rect 1986 37306 1996 37370
rect 2060 37306 2070 37370
rect 1463 37129 1547 37134
rect 1463 37065 1473 37129
rect 1537 37065 1547 37129
rect 1463 37060 1547 37065
rect 1996 36324 2060 37306
rect 15220 37246 15230 37310
rect 15294 37246 19337 37310
rect 19401 37246 19411 37310
rect 30746 37165 30756 37229
rect 30820 37165 31231 37229
rect 31295 37165 31305 37229
rect 2158 37149 2242 37154
rect 2158 36898 2168 37149
rect 2232 36898 2242 37149
rect 2158 36893 2242 36898
rect 2159 36668 2243 36673
rect 1986 36319 2070 36324
rect 1986 36255 1996 36319
rect 2060 36255 2070 36319
rect 1986 36250 2070 36255
rect 2159 36250 2169 36668
rect 2233 36250 2243 36668
rect 15980 36664 15990 36728
rect 16054 36664 19882 36728
rect 19946 36664 19956 36728
rect 6335 36597 6419 36602
rect 2159 36245 2243 36250
rect 2461 36533 6345 36597
rect 6409 36533 6419 36597
rect -18893 36119 -18797 36124
rect 2461 35941 2525 36533
rect 6335 36528 6419 36533
rect 30212 36529 30222 36593
rect 30286 36529 30584 36593
rect 30648 36529 30658 36593
rect 6345 36523 6409 36528
rect 6345 36258 6409 36264
rect 6335 36253 6419 36258
rect 6335 36189 6345 36253
rect 6409 36189 6419 36253
rect 6335 36184 6419 36189
rect 3122 36093 3241 36135
rect 5045 36104 5361 36109
rect 3572 36094 3821 36099
rect 2928 36088 3353 36093
rect 2928 36030 2938 36088
rect 3343 36030 3353 36088
rect 2928 36025 3353 36030
rect 3572 36030 3582 36094
rect 3811 36030 3821 36094
rect 3572 36025 3821 36030
rect -9218 35877 -9208 35941
rect -9144 35877 2525 35941
rect 3122 35672 3241 36025
rect 5045 36018 5055 36104
rect 5351 36018 5361 36104
rect 5564 36097 5811 36102
rect 5564 36027 5574 36097
rect 5801 36027 5811 36097
rect 5564 36022 5811 36027
rect 5045 36013 5361 36018
rect 3111 35553 3121 35672
rect 3240 35553 3250 35672
rect 6345 35351 6409 36184
rect 7503 36099 7622 36121
rect 7373 36094 7691 36099
rect 6926 36089 7167 36094
rect 6926 36020 6936 36089
rect 7157 36020 7167 36089
rect 7373 36028 7383 36094
rect 7681 36028 7691 36094
rect 7373 36023 7691 36028
rect 8911 36093 9358 36098
rect 8911 36028 8921 36093
rect 9348 36028 9358 36093
rect 8911 36023 9358 36028
rect 9565 36091 9812 36096
rect 9565 36023 9575 36091
rect 9802 36023 9812 36091
rect 6926 36015 7167 36020
rect 7503 35641 7622 36023
rect 9070 35650 9189 36023
rect 9565 36018 9812 36023
rect 16711 35986 16721 36050
rect 16785 35986 21517 36050
rect 21581 35986 21591 36050
rect 29663 35906 29673 35970
rect 29737 35906 29990 35970
rect 30054 35906 30064 35970
rect 7493 35522 7503 35641
rect 7622 35522 7632 35641
rect 9060 35531 9070 35650
rect 9189 35531 9199 35650
rect -10079 35287 -10069 35351
rect -10005 35287 6409 35351
rect 17402 35279 17412 35343
rect 17476 35279 22051 35343
rect 22115 35279 22125 35343
rect 29119 35194 29129 35258
rect 29193 35194 29407 35258
rect 29471 35194 29481 35258
rect -27087 34980 -26986 34985
rect -27089 34691 -26990 34696
rect -27089 33498 -27079 34691
rect -27000 33498 -26990 34691
rect -9379 34676 -9295 34681
rect -13405 34612 -13395 34676
rect -13331 34612 -9369 34676
rect -9305 34612 -9295 34676
rect -9379 34607 -9295 34612
rect 18242 34519 18252 34583
rect 18316 34519 22598 34583
rect 22662 34519 22672 34583
rect 26938 34458 26948 34522
rect 27012 34458 28828 34522
rect 28892 34458 28902 34522
rect 5922 34195 6006 34200
rect -4723 34131 -4713 34195
rect -4649 34131 5932 34195
rect 5996 34131 6006 34195
rect 5922 34126 6006 34131
rect 6728 33850 6812 33855
rect -4133 33786 -4123 33850
rect -4059 33786 6738 33850
rect 6802 33786 6812 33850
rect 6728 33781 6812 33786
rect 27495 33749 27505 33813
rect 27569 33749 28315 33813
rect 28379 33749 28389 33813
rect 19245 33682 19255 33746
rect 19319 33682 23143 33746
rect 23207 33682 23217 33746
rect -27089 33493 -26990 33498
rect -21540 33551 -21434 33575
rect -21540 33487 -21518 33551
rect -21454 33487 -21434 33551
rect -21540 33466 -21434 33487
rect -6958 33179 -6874 33184
rect -15149 33115 -15139 33179
rect -15075 33115 -6948 33179
rect -6884 33115 -6874 33179
rect -6958 33110 -6874 33115
rect -27094 32899 -26995 32904
rect -27094 32365 -27084 32899
rect -27005 32365 -26995 32899
rect -27094 32360 -26995 32365
rect 7354 32352 7438 32357
rect 5307 32345 5391 32350
rect 5121 32281 5317 32345
rect 5381 32281 5391 32345
rect 7354 32288 7364 32352
rect 7428 32288 7607 32352
rect 7354 32283 7438 32288
rect 5307 32276 5391 32281
rect 4964 31452 5028 32173
rect 7702 31452 7766 32173
rect 7942 31811 8053 31841
rect 7942 31747 7965 31811
rect 8029 31747 8053 31811
rect 7942 31723 8053 31747
rect 4964 31375 5028 31388
rect 7702 31375 7766 31388
rect 11337 31327 11347 31391
rect 11411 31327 13831 31391
rect 13895 31327 13905 31391
rect 5702 31191 5766 31192
rect 3944 31123 4742 31187
rect 4941 31127 5766 31191
rect 3961 30389 4025 31123
rect 4325 30432 4440 30460
rect 4325 30368 4354 30432
rect 4418 30368 4440 30432
rect 5702 30394 5766 31127
rect 6964 31191 7028 31192
rect 6964 31127 7789 31191
rect 6964 30394 7028 31127
rect 7988 31123 8786 31187
rect 8300 30437 8415 30464
rect 4325 30342 4440 30368
rect 8300 30373 8328 30437
rect 8392 30373 8415 30437
rect 8705 30389 8769 31123
rect 11956 30708 11966 30772
rect 12030 30708 14586 30772
rect 14650 30708 14660 30772
rect 50606 30469 50842 39730
rect 52801 33632 53037 41020
rect 55146 37094 55382 41987
rect 57729 40402 57965 42541
rect 57729 40166 62907 40402
rect 55146 36858 62907 37094
rect 52801 33396 62907 33632
rect 8300 30348 8415 30373
rect 3298 30305 3418 30335
rect 3298 30241 3326 30305
rect 3390 30241 3418 30305
rect 3298 30212 3418 30241
rect 50606 30233 62907 30469
rect -12703 29752 -12619 29757
rect 1903 29752 1987 29757
rect -12703 29688 -12693 29752
rect -12629 29688 -3918 29752
rect -3854 29688 1913 29752
rect 1977 29688 1987 29752
rect -12703 29683 -12619 29688
rect 1903 29683 1987 29688
rect 3961 29389 4025 30187
rect 4328 29982 4609 30046
rect -13479 29329 -13395 29334
rect 1903 29329 1987 29334
rect -13479 29265 -13469 29329
rect -13405 29265 -5279 29329
rect -5215 29265 1913 29329
rect 1977 29265 1987 29329
rect -13479 29260 -13395 29265
rect 1903 29260 1987 29265
rect 3961 28389 4025 29187
rect 4328 28600 4392 29982
rect 5702 29394 5766 30192
rect 6964 29394 7028 30192
rect 8121 29982 8402 30046
rect 4701 28813 4765 29012
rect 4691 28808 4775 28813
rect 4691 28744 4701 28808
rect 4765 28744 4775 28808
rect 4691 28739 4775 28744
rect 4318 28595 4402 28600
rect 4318 28531 4328 28595
rect 4392 28593 4402 28595
rect 4392 28531 4579 28593
rect 4318 28529 4579 28531
rect 4318 28526 4402 28529
rect 5702 28394 5766 29192
rect 6964 28394 7028 29192
rect 7960 28851 8024 29021
rect 7950 28846 8034 28851
rect 7950 28782 7960 28846
rect 8024 28782 8034 28846
rect 7950 28777 8034 28782
rect 8338 28597 8402 29982
rect 8705 29389 8769 30187
rect 16692 29752 16811 29781
rect 16692 29688 16721 29752
rect 16785 29688 16811 29752
rect 16692 29659 16811 29688
rect 17378 29329 17506 29366
rect 17378 29265 17412 29329
rect 17476 29265 17506 29329
rect 17378 29232 17506 29265
rect 8328 28593 8412 28597
rect 8151 28592 8412 28593
rect 8151 28529 8338 28592
rect 8328 28528 8338 28529
rect 8402 28528 8412 28592
rect 8328 28523 8412 28528
rect 8705 28389 8769 29187
rect 10623 28740 10633 28804
rect 10697 28740 11966 28804
rect 12030 28740 12040 28804
rect -15722 28098 -15603 28103
rect -17645 27644 -17497 27649
rect -17645 27516 -17635 27644
rect -17507 27516 -17497 27644
rect -15722 27645 -15712 28098
rect -15613 27645 -15603 28098
rect -12399 28076 -12306 28081
rect -12399 27670 -12389 28076
rect -12316 27670 -12306 28076
rect -12399 27665 -12306 27670
rect -15722 27640 -15603 27645
rect -17645 27511 -17497 27516
rect -5309 27532 -5186 27565
rect -5309 27468 -5279 27532
rect -5215 27468 -5186 27532
rect -5309 27440 -5186 27468
rect 3961 27451 4025 28187
rect 5702 27451 5766 28192
rect -12404 27427 -12287 27432
rect -12404 27198 -12394 27427
rect -12297 27198 -12287 27427
rect 3961 27389 4764 27451
rect 3966 27387 4764 27389
rect 4966 27394 5766 27451
rect 6964 27451 7028 28192
rect 8705 27451 8769 28187
rect 6964 27394 7764 27451
rect 4966 27387 5764 27394
rect 6966 27387 7764 27394
rect 7966 27389 8769 27451
rect 7966 27387 8764 27389
rect -12404 27193 -12287 27198
rect -3948 26855 -3825 26889
rect -3948 26791 -3918 26855
rect -3854 26791 -3825 26855
rect -3948 26764 -3825 26791
rect -38200 26611 -34846 26616
rect -38200 26514 -38190 26611
rect -34856 26514 -34846 26611
rect -38200 26509 -34846 26514
rect -12406 26486 -12291 26491
rect -17645 26415 -17497 26420
rect -17645 26287 -17635 26415
rect -17507 26287 -17497 26415
rect -17645 26282 -17497 26287
rect -15735 26281 -15626 26286
rect -15735 26044 -15725 26281
rect -15636 26044 -15626 26281
rect -12406 26057 -12396 26486
rect -12301 26057 -12291 26486
rect 4966 26402 5030 27200
rect 7700 26402 7764 27200
rect 11337 26286 11347 26350
rect 11411 26286 11837 26350
rect 11901 26286 11911 26350
rect -12406 26052 -12291 26057
rect -15735 26039 -15626 26044
rect 19861 26009 19945 26014
rect 13840 25945 13850 26009
rect 13914 25945 19871 26009
rect 19935 25945 25879 26009
rect 25943 25945 25950 26009
rect 19861 25940 19945 25945
rect -12394 25823 -12311 25828
rect -19098 25571 -19088 25804
rect -18855 25571 -15505 25804
rect -13999 25664 -13915 25669
rect -13999 25600 -13989 25664
rect -13925 25600 -12544 25664
rect -13999 25595 -13915 25600
rect -18560 25570 -18327 25571
rect -25459 25482 -25359 25487
rect -40603 25171 -40347 25176
rect -57094 24935 -40593 25171
rect -40357 24935 -40347 25171
rect -25459 25175 -25449 25482
rect -25369 25175 -25359 25482
rect -25459 25170 -25359 25175
rect -15738 25447 -15505 25571
rect -15738 25018 -15727 25447
rect -15632 25018 -15505 25447
rect -12608 25419 -12544 25600
rect -12394 25604 -12384 25823
rect -12321 25604 -12311 25823
rect -12394 25599 -12311 25604
rect -12177 25600 -11324 25664
rect -11260 25600 -11250 25664
rect -12177 25419 -12113 25600
rect 19863 25598 19947 25603
rect 13256 25534 13266 25598
rect 13330 25534 19873 25598
rect 19937 25534 26463 25598
rect 26527 25534 26537 25598
rect 19863 25529 19947 25534
rect -12608 25355 -12113 25419
rect -15738 25011 -15505 25018
rect -17645 25002 -17497 25007
rect -40603 24930 -40347 24935
rect -25462 24945 -25355 24950
rect -25462 24714 -25452 24945
rect -25365 24714 -25355 24945
rect -17645 24874 -17635 25002
rect -17507 24874 -17497 25002
rect -17645 24869 -17497 24874
rect -14420 24872 -14336 24877
rect -14420 24808 -14410 24872
rect -14346 24808 -11977 24872
rect -11913 24808 -11903 24872
rect -14420 24803 -14336 24808
rect 7591 24784 7601 24848
rect 7665 24784 15230 24848
rect 15294 24784 15304 24848
rect -25462 24709 -25355 24714
rect -12403 24712 -12318 24717
rect -12403 24458 -12393 24712
rect -12328 24458 -12318 24712
rect -12403 24453 -12318 24458
rect 5705 24594 5793 24599
rect -12408 24239 -12306 24244
rect -12408 24003 -12398 24239
rect -12316 24003 -12306 24239
rect 5705 24186 5715 24594
rect 5783 24186 5793 24594
rect 7058 24592 7142 24597
rect 7256 24592 7266 24593
rect 7058 24528 7068 24592
rect 7132 24529 7266 24592
rect 7330 24529 7340 24593
rect 7132 24528 7290 24529
rect 7058 24523 7142 24528
rect 8119 24466 8129 24530
rect 8193 24466 15990 24530
rect 16054 24466 16064 24530
rect 5705 24181 5793 24186
rect 11073 24138 11080 24202
rect 11144 24138 19929 24202
rect -12408 23998 -12306 24003
rect -11334 23823 -11324 23887
rect -11260 23823 7266 23887
rect 7330 23823 19255 23887
rect 19319 23823 19329 23887
rect -17645 23773 -17497 23778
rect -17645 23645 -17635 23773
rect -17507 23645 -17497 23773
rect -17645 23640 -17497 23645
rect 7081 23652 7165 23657
rect -15735 23637 -15648 23642
rect -38192 23605 -34842 23610
rect -38192 23503 -38182 23605
rect -34852 23503 -34842 23605
rect -38192 23498 -34842 23503
rect -15735 23405 -15725 23637
rect -15658 23405 -15648 23637
rect 7081 23588 7091 23652
rect 7155 23588 7165 23652
rect 7081 23583 7165 23588
rect 7091 23518 7155 23583
rect -11987 23454 -11977 23518
rect -11913 23454 18252 23518
rect 18316 23454 18326 23518
rect -15735 23400 -15648 23405
rect 8777 23356 8953 23361
rect -12399 23277 -12309 23282
rect -12399 22857 -12389 23277
rect -12319 22857 -12309 23277
rect 8777 23246 8787 23356
rect 8943 23246 8953 23356
rect 8777 23241 8953 23246
rect 19865 23210 19929 24138
rect 42846 24174 46200 24179
rect 42846 24065 42856 24174
rect 46190 24065 46200 24174
rect 42846 24060 46200 24065
rect 36045 24018 36148 24038
rect 36045 23954 36066 24018
rect 36130 23954 36148 24018
rect 36045 23934 36148 23954
rect 35126 23866 35241 23893
rect 35126 23802 35152 23866
rect 35216 23802 35241 23866
rect 35126 23772 35241 23802
rect 39336 23714 39430 23719
rect 37809 23611 37902 23616
rect 37809 23492 37819 23611
rect 37892 23492 37902 23611
rect 37809 23487 37902 23492
rect 39336 23493 39346 23714
rect 39420 23493 39430 23714
rect 39336 23488 39430 23493
rect 2540 23063 2624 23068
rect 4770 23063 4780 23159
rect 2540 22999 2550 23063
rect 2614 22999 4780 23063
rect 2540 22994 2624 22999
rect 4770 22919 4780 22999
rect 5243 23063 5253 23159
rect 12578 23146 12588 23210
rect 12652 23146 27111 23210
rect 27175 23146 27186 23210
rect 39325 23200 39431 23205
rect 37809 23194 37915 23199
rect 10192 23063 10276 23068
rect 5243 22999 5718 23063
rect 5782 22999 10202 23063
rect 10266 22999 10276 23063
rect 5243 22919 5253 22999
rect 10192 22994 10276 22999
rect 11836 22916 11900 22979
rect 37809 22946 37819 23194
rect 37905 22946 37915 23194
rect 39325 22952 39335 23200
rect 39421 22952 39431 23200
rect 39325 22947 39431 22952
rect 37809 22941 37915 22946
rect 11827 22915 11837 22916
rect -12399 22852 -12309 22857
rect 11466 22851 11476 22915
rect 11540 22852 11837 22915
rect 11901 22915 11911 22916
rect 11901 22852 14589 22915
rect 11540 22851 14589 22852
rect -12762 22724 -12087 22777
rect -16609 22660 -16599 22724
rect -16535 22713 8129 22724
rect -16535 22660 -12687 22713
rect -12151 22660 8129 22713
rect 8193 22660 8203 22724
rect -12401 22624 -12313 22629
rect -12401 22399 -12391 22624
rect -12323 22399 -12313 22624
rect -12401 22394 -12313 22399
rect -17046 22209 7601 22273
rect 7665 22209 7675 22273
rect -17046 21097 -16982 22209
rect 14525 22091 14589 22851
rect 15481 22851 16400 22915
rect 15481 22091 15545 22851
rect 14525 22027 15545 22091
rect 16336 22084 16400 22851
rect 17405 22851 18389 22915
rect 17405 22084 17469 22851
rect 18325 22493 18389 22851
rect 18900 22851 19930 22915
rect 18900 22493 18964 22851
rect 18325 22429 18964 22493
rect 16336 22020 17469 22084
rect 19866 21655 19930 22851
rect 35090 22790 35290 22795
rect 36904 22790 36914 22815
rect 35090 22610 35100 22790
rect 35280 22730 36914 22790
rect 35280 22668 35760 22730
rect 36021 22668 36914 22730
rect 35280 22610 36914 22668
rect 35090 22605 35290 22610
rect 36904 22579 36914 22610
rect 37156 22579 37166 22815
rect 47546 22734 47802 22739
rect 47546 22498 47556 22734
rect 47792 22498 62907 22734
rect 47546 22493 47802 22498
rect 39336 22388 39430 22393
rect 37816 22280 37906 22285
rect 37816 22151 37826 22280
rect 37896 22151 37906 22280
rect 39336 22167 39346 22388
rect 39420 22167 39430 22388
rect 39336 22162 39430 22167
rect 37816 22146 37906 22151
rect 39331 21834 39437 21839
rect 37804 21823 37909 21828
rect -981 21625 -897 21630
rect 6297 21625 6381 21630
rect -981 21561 -971 21625
rect -907 21561 6307 21625
rect 6371 21561 6381 21625
rect 12062 21591 12072 21655
rect 12136 21591 27657 21655
rect 27721 21591 27731 21655
rect 37804 21621 37814 21823
rect 37899 21621 37909 21823
rect 37804 21616 37909 21621
rect -981 21556 -897 21561
rect 6297 21556 6381 21561
rect 35126 21585 35244 21615
rect 35126 21521 35152 21585
rect 35216 21521 35244 21585
rect 39331 21586 39341 21834
rect 39427 21586 39437 21834
rect 39331 21581 39437 21586
rect 35126 21488 35244 21521
rect 35457 21379 35564 21402
rect 35457 21315 35477 21379
rect 35541 21315 35564 21379
rect 35457 21293 35564 21315
rect 42844 21178 46198 21183
rect -27920 21033 6374 21097
rect 42844 21069 42854 21178
rect 46188 21069 46198 21178
rect 42844 21064 46198 21069
rect -38178 19065 -34851 19070
rect -38178 18987 -38168 19065
rect -34861 18987 -34851 19065
rect -38178 18982 -34851 18987
rect -40606 17630 -40350 17635
rect -57094 17394 -40596 17630
rect -40360 17394 -40350 17630
rect -40606 17389 -40350 17394
rect -38184 16075 -34842 16080
rect -38184 15987 -38174 16075
rect -34852 15987 -34842 16075
rect -38184 15982 -34842 15987
rect -27920 15446 -27856 21033
rect 6310 20962 6374 21033
rect 14678 21027 14762 21032
rect 12926 20963 12936 21027
rect 13000 20963 14688 21027
rect 14752 20963 14762 21027
rect 6300 20957 6384 20962
rect 14678 20958 14762 20963
rect 6300 20893 6310 20957
rect 6374 20893 6384 20957
rect 6300 20888 6384 20893
rect -981 20715 -897 20720
rect -24170 20651 -971 20715
rect -907 20651 -897 20715
rect -25462 17922 -25377 17927
rect -25462 17627 -25452 17922
rect -25387 17627 -25377 17922
rect -25462 17622 -25377 17627
rect -25460 17404 -25368 17409
rect -25460 17169 -25450 17404
rect -25378 17169 -25368 17404
rect -25460 17164 -25368 17169
rect -24170 16254 -24106 20651
rect -16609 20587 -16599 20651
rect -16535 20587 -16525 20651
rect -981 20646 -897 20651
rect -7442 20270 11080 20334
rect 11144 20270 11154 20334
rect -12387 17968 -12259 17999
rect -12387 17904 -12355 17968
rect -12291 17904 -12259 17968
rect -12387 17870 -12259 17904
rect -10445 17157 -10321 17194
rect -10445 17093 -10416 17157
rect -10352 17093 -10321 17157
rect -10445 17061 -10321 17093
rect -10425 16288 -10341 16293
rect -24180 16249 -24096 16254
rect -24180 16185 -24170 16249
rect -24106 16185 -24096 16249
rect -18719 16203 -17699 16267
rect -16119 16203 -15099 16267
rect -13519 16203 -12499 16267
rect -10785 16224 -10415 16288
rect -10351 16224 -10341 16288
rect -10425 16219 -10341 16224
rect -24180 16180 -24096 16185
rect -27930 15441 -27846 15446
rect -27930 15377 -27920 15441
rect -27856 15377 -27846 15441
rect -27930 15372 -27846 15377
rect -19071 14880 -19007 15900
rect -12197 14873 -12133 15893
rect -15965 14472 -15232 14536
rect -25527 14446 -25434 14451
rect -25527 14157 -25517 14446
rect -25444 14157 -25434 14446
rect -25527 14152 -25434 14157
rect -13074 14141 -12990 14146
rect -18240 14073 -18139 14097
rect -13331 14077 -13064 14141
rect -13000 14077 -12990 14141
rect -18240 14009 -18223 14073
rect -18159 14009 -18139 14073
rect -13074 14072 -12990 14077
rect -18240 13986 -18139 14009
rect -25528 13925 -25436 13930
rect -25528 13690 -25518 13925
rect -25446 13690 -25436 13925
rect -25528 13685 -25436 13690
rect -19071 12280 -19007 13300
rect -12197 12273 -12133 13293
rect -18722 11937 -17702 12001
rect -16122 11937 -15102 12001
rect -13522 11937 -12502 12001
rect -10999 10223 -10881 10250
rect -13969 10181 -13846 10211
rect -13969 10117 -13941 10181
rect -13877 10117 -13846 10181
rect -10999 10159 -10970 10223
rect -10906 10159 -10881 10223
rect -10999 10138 -10881 10159
rect -13969 10089 -13846 10117
rect -7442 9819 -7378 20270
rect -6759 19739 11476 19803
rect 11540 19739 11550 19803
rect -6759 10646 -6695 19739
rect 41 19513 125 19518
rect -2825 19449 -2815 19513
rect -2751 19449 51 19513
rect 115 19449 125 19513
rect -5289 18979 -5279 19043
rect -5215 18979 -5205 19043
rect -3928 18979 -3918 19043
rect -3854 18979 -3844 19043
rect -5279 18871 -5215 18979
rect -5279 18807 -4725 18871
rect -3918 18870 -3854 18979
rect -5815 15708 -5690 15744
rect -5815 15644 -5786 15708
rect -5722 15644 -5690 15708
rect -5815 15613 -5690 15644
rect -4789 14637 -4725 18807
rect -4448 18806 -3854 18870
rect -4789 14573 -4552 14637
rect -4912 14446 -4822 14451
rect -4912 14236 -4902 14446
rect -4832 14236 -4822 14446
rect -4912 14231 -4822 14236
rect -4914 14003 -4850 14011
rect -4927 13998 -4823 14003
rect -4927 13706 -4917 13998
rect -4833 13706 -4823 13998
rect -4927 13701 -4823 13706
rect -4914 13279 -4850 13701
rect -5014 13215 -4850 13279
rect -5717 10838 -5391 10843
rect -5014 10838 -4950 13215
rect -4616 12380 -4552 14573
rect -6172 10833 -5927 10838
rect -6172 10758 -6162 10833
rect -5937 10758 -5927 10833
rect -5735 10774 -5707 10838
rect -6172 10753 -5927 10758
rect -5717 10751 -5707 10774
rect -5401 10774 -4950 10838
rect -5401 10751 -5391 10774
rect -5717 10746 -5391 10751
rect -6759 10582 -6092 10646
rect -6156 10209 -6092 10582
rect -6166 10204 -6082 10209
rect -6166 10140 -6156 10204
rect -6092 10140 -6082 10204
rect -6166 10135 -6082 10140
rect -5371 10204 -5287 10209
rect -5371 10140 -5361 10204
rect -5297 10140 -5287 10204
rect -5371 10135 -5287 10140
rect -5361 9819 -5297 10135
rect -7442 9755 -5297 9819
rect -6177 9592 -5919 9597
rect -6177 9513 -6167 9592
rect -5929 9513 -5919 9592
rect -6177 9508 -5919 9513
rect -5718 9595 -5389 9600
rect -5718 9509 -5708 9595
rect -5399 9572 -5389 9595
rect -5014 9572 -4950 10774
rect -4789 12316 -4552 12380
rect -4789 10238 -4725 12316
rect -4448 10238 -4384 18806
rect -2815 18299 -2751 19449
rect 41 19444 125 19449
rect 23667 19382 23776 19404
rect 23667 19318 23689 19382
rect 23753 19318 23776 19382
rect 14657 19278 14771 19303
rect 23667 19292 23776 19318
rect -766 19212 -682 19217
rect -2408 19148 -2398 19212
rect -2334 19148 -756 19212
rect -692 19148 -682 19212
rect 14657 19214 14686 19278
rect 14750 19214 14771 19278
rect 14657 19183 14771 19214
rect -766 19143 -682 19148
rect 4847 19173 5204 19178
rect 3051 19106 3135 19111
rect 4847 19106 4857 19173
rect 3051 19042 3061 19106
rect 3125 19042 4857 19106
rect 3051 19037 3135 19042
rect 4847 19027 4857 19042
rect 5194 19106 5204 19173
rect 7075 19106 7159 19111
rect 8971 19106 9055 19111
rect 5194 19042 7085 19106
rect 7149 19042 8981 19106
rect 9045 19042 9089 19106
rect 10203 19058 10327 19083
rect 5194 19027 5204 19042
rect 7075 19037 7159 19042
rect 8971 19037 9055 19042
rect 4847 19022 5204 19027
rect 10203 18994 10232 19058
rect 10296 18994 10327 19058
rect 10203 18968 10327 18994
rect 20928 19062 21079 19106
rect 20928 18998 20971 19062
rect 21035 18998 21079 19062
rect 20928 18951 21079 18998
rect 5697 18910 5781 18915
rect 7696 18910 7780 18915
rect -1514 18846 -1504 18910
rect -1440 18846 5707 18910
rect 5771 18846 7706 18910
rect 7770 18846 7780 18910
rect 5697 18841 5781 18846
rect 7696 18841 7780 18846
rect 8239 18718 8373 18758
rect 4889 18651 4973 18656
rect 6887 18651 6971 18656
rect -1143 18587 -1133 18651
rect -1069 18587 4899 18651
rect 4963 18587 6897 18651
rect 6961 18587 6971 18651
rect 8239 18654 8280 18718
rect 8344 18654 8373 18718
rect 13564 18688 13648 18693
rect 8239 18617 8373 18654
rect 12920 18624 12930 18688
rect 12994 18624 13574 18688
rect 13638 18624 13648 18688
rect 13564 18619 13648 18624
rect 4889 18582 4973 18587
rect 6887 18582 6971 18587
rect 14105 18507 14115 18571
rect 14179 18507 14189 18571
rect 25604 18507 25614 18571
rect 25678 18507 25688 18571
rect 3697 18312 3781 18317
rect 9696 18312 9780 18317
rect -3509 18235 -2751 18299
rect -690 18248 -680 18312
rect -616 18248 3707 18312
rect 3771 18248 9706 18312
rect 9770 18248 9780 18312
rect 3697 18243 3781 18248
rect 9696 18243 9780 18248
rect -3509 16205 -3445 18235
rect 2888 18031 2972 18036
rect 8889 18031 8973 18036
rect -294 17967 -284 18031
rect -220 17967 2898 18031
rect 2962 17967 8899 18031
rect 8963 17967 8973 18031
rect 2888 17962 2972 17967
rect 8889 17962 8973 17967
rect -3221 17624 -3211 17864
rect -2748 17772 -2738 17864
rect 223 17772 307 17777
rect -2748 17708 233 17772
rect 297 17708 307 17772
rect -2748 17624 -2738 17708
rect 223 17703 307 17708
rect 14358 17699 14368 17763
rect 14432 17699 14442 17763
rect 25351 17700 25361 17764
rect 25425 17700 25435 17764
rect 14659 17549 14776 17576
rect -831 17525 -747 17530
rect -847 17461 -821 17525
rect -757 17461 981 17525
rect 1045 17461 1077 17525
rect 14659 17485 14689 17549
rect 14753 17485 14776 17549
rect -831 17456 -747 17461
rect 14659 17455 14776 17485
rect 23665 17552 23778 17575
rect 23665 17488 23689 17552
rect 23753 17488 23778 17552
rect 23665 17458 23778 17488
rect 4268 17289 4387 17313
rect 4268 17225 4295 17289
rect 4359 17225 4387 17289
rect 4268 17194 4387 17225
rect 6200 17289 6319 17314
rect 6200 17225 6227 17289
rect 6291 17225 6319 17289
rect 6200 17195 6319 17225
rect 13593 17083 13677 17088
rect 12946 17019 12956 17083
rect 13020 17019 13603 17083
rect 13667 17019 13677 17083
rect 13593 17014 13677 17019
rect 18 16446 11149 16451
rect 18 16413 251 16446
rect -2932 16252 251 16413
rect 18 16238 251 16252
rect 11139 16238 11149 16446
rect 18 16233 11149 16238
rect -3519 16141 -3509 16205
rect -3445 16141 -3435 16205
rect 18 16189 248 16233
rect -3018 15454 -2934 15459
rect -3938 15390 -3928 15454
rect -3864 15390 -3008 15454
rect -2944 15390 -2934 15454
rect -3018 15385 -2934 15390
rect -3154 14998 -3051 15003
rect -3154 14719 -3144 14998
rect -3061 14719 -3051 14998
rect -3154 14714 -3051 14719
rect -3033 14644 -2949 14649
rect -3519 14580 -3509 14644
rect -3445 14580 -3023 14644
rect -2959 14580 -2949 14644
rect -3033 14575 -2949 14580
rect 18 13993 28 16189
rect -2956 13832 28 13993
rect -2608 13137 -2524 13142
rect -2608 13073 -2598 13137
rect -2534 13073 -2524 13137
rect -2608 13068 -2524 13073
rect -1818 13133 -1715 13138
rect -2895 12328 -2811 12333
rect -2895 12264 -2885 12328
rect -2821 12264 -2811 12328
rect -2895 12259 -2811 12264
rect -4799 10233 -4715 10238
rect -4799 10169 -4789 10233
rect -4725 10169 -4715 10233
rect -4799 10164 -4715 10169
rect -4458 10233 -4374 10238
rect -4458 10169 -4448 10233
rect -4384 10169 -4374 10233
rect -4458 10164 -4374 10169
rect -5399 9509 -4950 9572
rect -5718 9508 -4950 9509
rect -5718 9504 -5389 9508
rect -5014 8707 -4950 9508
rect -5014 8643 -3185 8707
rect -3121 8643 -3111 8707
rect -18719 8403 -17699 8467
rect -16119 8403 -15099 8467
rect -13519 8403 -12499 8467
rect -19071 7080 -19007 8100
rect -12197 7073 -12133 8093
rect -2885 7532 -2821 12259
rect -2598 8340 -2534 13068
rect -1818 12726 -1808 13133
rect -1725 12726 -1715 13133
rect -1818 12721 -1715 12726
rect -1508 12409 -1424 12414
rect -1508 12345 -1498 12409
rect -1434 12345 -1424 12409
rect -1508 12340 -1424 12345
rect -1936 11535 -1852 11540
rect -1936 11471 -1926 11535
rect -1862 11471 -1852 11535
rect -1936 11466 -1852 11471
rect -1769 11529 -1683 11534
rect -2222 10729 -2138 10734
rect -2222 10665 -2212 10729
rect -2148 10665 -2138 10729
rect -2222 10660 -2138 10665
rect -2212 9134 -2148 10660
rect -1926 9942 -1862 11466
rect -1769 11140 -1759 11529
rect -1693 11140 -1683 11529
rect -1769 11135 -1683 11140
rect -1498 10788 -1434 12340
rect -1508 10783 -1424 10788
rect -1508 10719 -1498 10783
rect -1434 10719 -1424 10783
rect -1508 10714 -1424 10719
rect -1936 9937 -1852 9942
rect -1936 9873 -1926 9937
rect -1862 9873 -1852 9937
rect -1936 9868 -1852 9873
rect -1769 9930 -1685 9935
rect -2222 9129 -2138 9134
rect -2222 9065 -2212 9129
rect -2148 9065 -2138 9129
rect -2222 9060 -2138 9065
rect -2608 8335 -2524 8340
rect -2608 8271 -2598 8335
rect -2534 8271 -2524 8335
rect -2608 8266 -2524 8271
rect -2895 7527 -2811 7532
rect -2895 7463 -2885 7527
rect -2821 7463 -2811 7527
rect -2895 7458 -2811 7463
rect -7224 7243 -6741 7248
rect -7224 7003 -7214 7243
rect -6751 7003 -6741 7243
rect -7224 6998 -6741 7003
rect -25531 6669 -25436 6674
rect -15965 6672 -15232 6736
rect -4927 6695 -4826 6700
rect -25531 6408 -25521 6669
rect -25446 6408 -25436 6669
rect -25531 6403 -25436 6408
rect -4927 6392 -4917 6695
rect -4836 6649 -4826 6695
rect -4836 6585 -3184 6649
rect -3120 6585 -3110 6649
rect -4836 6392 -4826 6585
rect -4927 6387 -4826 6392
rect -18271 6303 -18171 6328
rect -13085 6313 -13001 6318
rect -18271 6239 -18251 6303
rect -18187 6239 -18171 6303
rect -13326 6249 -13075 6313
rect -13011 6249 -13001 6313
rect -13085 6244 -13001 6249
rect -18271 6217 -18171 6239
rect -25532 6174 -25437 6179
rect -25532 5929 -25522 6174
rect -25447 5929 -25437 6174
rect -4917 6163 -4831 6168
rect -4917 5950 -4907 6163
rect -4841 5950 -4831 6163
rect -3060 6042 -2976 6047
rect -3938 5978 -3928 6042
rect -3864 5978 -3050 6042
rect -2986 5978 -2976 6042
rect -3060 5973 -2976 5978
rect -4917 5945 -4831 5950
rect -25532 5924 -25437 5929
rect -3203 5577 -3100 5582
rect -19071 4480 -19007 5500
rect -12197 4473 -12133 5493
rect -10766 5052 -10702 5314
rect -3203 5296 -3193 5577
rect -3110 5296 -3100 5577
rect -3203 5291 -3100 5296
rect -3038 5233 -2954 5238
rect -3519 5169 -3509 5233
rect -3445 5169 -3435 5233
rect -3038 5169 -3028 5233
rect -2964 5169 -2954 5233
rect -10776 5047 -10692 5052
rect -10776 4983 -10766 5047
rect -10702 4983 -10692 5047
rect -10776 4978 -10692 4983
rect -3509 4978 -3445 5169
rect -3038 5164 -2954 5169
rect -3031 4978 -2967 5164
rect -3509 4914 -2967 4978
rect -18722 4137 -17702 4201
rect -16122 4137 -15102 4201
rect -13522 4137 -12502 4201
rect -2885 -4979 -2821 7458
rect -2598 -4516 -2534 8266
rect -2212 -3981 -2148 9060
rect -1926 -3509 -1862 9868
rect -1769 9532 -1759 9930
rect -1695 9532 -1685 9930
rect -1769 9527 -1685 9532
rect -1498 9130 -1434 10714
rect 18 10640 28 13832
rect 187 16184 248 16189
rect 11229 16184 11409 16189
rect 187 10640 197 16184
rect 5468 14599 5666 14604
rect 5468 14421 5478 14599
rect 5656 14421 5666 14599
rect 11229 14426 11239 16184
rect 11399 15269 11409 16184
rect 23644 15788 23786 15820
rect 14650 15753 14786 15785
rect 14650 15689 14685 15753
rect 14749 15689 14786 15753
rect 14650 15653 14786 15689
rect 23644 15724 23686 15788
rect 23750 15724 23786 15788
rect 23644 15685 23786 15724
rect 20897 15496 21018 15526
rect 20897 15432 20928 15496
rect 20992 15432 21018 15496
rect 20897 15400 21018 15432
rect 11399 15228 13084 15269
rect 14680 15228 14764 15233
rect 11399 15164 12973 15228
rect 13037 15164 14690 15228
rect 14754 15164 14764 15228
rect 11399 15113 13084 15164
rect 14680 15159 14764 15164
rect 11399 14426 11409 15113
rect 11229 14421 11409 14426
rect 5468 14416 5666 14421
rect 23664 13997 23769 14018
rect 14650 13965 14778 13997
rect 11247 13954 11394 13959
rect 11247 13572 11257 13954
rect 11246 13426 11257 13572
rect 11247 12990 11257 13426
rect 11384 13572 11394 13954
rect 14650 13901 14685 13965
rect 14749 13901 14778 13965
rect 23664 13933 23686 13997
rect 23750 13933 23769 13997
rect 23664 13909 23769 13933
rect 14650 13860 14778 13901
rect 11384 13528 13075 13572
rect 13626 13528 13710 13533
rect 11384 13464 13003 13528
rect 13067 13464 13636 13528
rect 13700 13464 13710 13528
rect 11384 13426 13075 13464
rect 13626 13459 13710 13464
rect 11384 12990 11394 13426
rect 14105 13107 14115 13171
rect 14179 13107 14189 13171
rect 11247 12985 11394 12990
rect 14358 12299 14368 12363
rect 14432 12299 14442 12363
rect 14675 12180 14789 12202
rect 11233 12129 11408 12134
rect 4620 11980 4818 11985
rect 4620 11802 4630 11980
rect 4808 11802 4818 11980
rect 4620 11797 4818 11802
rect 11233 11316 11243 12129
rect 11398 11724 11408 12129
rect 14675 12116 14702 12180
rect 14766 12116 14789 12180
rect 14675 12087 14789 12116
rect 23667 12190 23779 12214
rect 23667 12126 23691 12190
rect 23755 12126 23779 12190
rect 23667 12098 23779 12126
rect 20945 11906 21080 11947
rect 20945 11842 20985 11906
rect 21049 11842 21080 11906
rect 20945 11804 21080 11842
rect 11398 11676 13124 11724
rect 13689 11676 13773 11681
rect 11398 11612 13001 11676
rect 13065 11612 13699 11676
rect 13763 11612 13773 11676
rect 11398 11560 13124 11612
rect 13689 11607 13773 11612
rect 11398 11316 11408 11560
rect 11233 11311 11408 11316
rect 18 10635 197 10640
rect 6473 10537 11228 10542
rect 6473 10356 6483 10537
rect 11218 10356 11228 10537
rect 6473 10351 11228 10356
rect 14666 10383 14780 10406
rect 14666 10319 14691 10383
rect 14755 10319 14780 10383
rect 14666 10290 14780 10319
rect 23664 10380 23783 10410
rect 23664 10316 23691 10380
rect 23755 10316 23783 10380
rect 23664 10286 23783 10316
rect 13866 10150 21128 10155
rect 362 10144 1822 10149
rect 362 10003 372 10144
rect 1812 10003 1822 10144
rect 362 9998 1822 10003
rect 5717 10135 11732 10140
rect 5717 9990 5727 10135
rect 11722 9990 11732 10135
rect 5717 9985 11732 9990
rect 13866 9993 13876 10150
rect 21118 9993 21128 10150
rect 13866 9988 21128 9993
rect 19 9830 222 9835
rect -1508 9125 -1424 9130
rect -1508 9061 -1498 9125
rect -1434 9061 -1424 9125
rect -1508 9056 -1424 9061
rect -1768 8330 -1680 8335
rect -1768 7930 -1758 8330
rect -1690 7930 -1680 8330
rect -1768 7925 -1680 7930
rect -1498 7591 -1434 9056
rect -1508 7586 -1424 7591
rect -1508 7522 -1498 7586
rect -1434 7522 -1424 7586
rect -1508 7517 -1424 7522
rect -1498 7263 -1434 7517
rect -1508 7258 -1424 7263
rect -1508 6974 -1498 7258
rect -1434 6974 -1424 7258
rect -1508 6969 -1424 6974
rect -1498 6456 -1434 6969
rect -1508 6451 -1424 6456
rect -1508 6387 -1498 6451
rect -1434 6387 -1424 6451
rect -1508 6382 -1424 6387
rect 19 5570 29 9830
rect 212 5570 222 9830
rect 36043 9154 36151 9176
rect 36043 9090 36066 9154
rect 36130 9090 36151 9154
rect 36043 9064 36151 9090
rect 36888 8705 36898 8792
rect 34644 8641 36898 8705
rect 17636 8451 17834 8456
rect 4669 8366 4867 8371
rect 4669 8188 4679 8366
rect 4857 8188 4867 8366
rect 17636 8273 17646 8451
rect 17824 8273 17834 8451
rect 17636 8268 17834 8273
rect 34644 8336 34708 8641
rect 35459 8531 35583 8563
rect 36888 8556 36898 8641
rect 37140 8556 37150 8792
rect 35459 8467 35489 8531
rect 35553 8467 35583 8531
rect 35459 8436 35583 8467
rect 36604 8469 36720 8498
rect 36604 8405 36631 8469
rect 36695 8405 36720 8469
rect 36604 8377 36720 8405
rect 34644 8288 35088 8336
rect 34644 8283 35098 8288
rect 34644 8272 35024 8283
rect 4669 8183 4867 8188
rect 21240 7514 21427 7519
rect 13340 6491 13538 6496
rect 4669 6366 4867 6371
rect 4669 6188 4679 6366
rect 4857 6188 4867 6366
rect 13340 6313 13350 6491
rect 13528 6313 13538 6491
rect 13340 6308 13538 6313
rect 17636 6451 17834 6456
rect 17636 6273 17646 6451
rect 17824 6273 17834 6451
rect 17636 6268 17834 6273
rect 4669 6183 4867 6188
rect 19 5565 222 5570
rect 16091 5088 16289 5093
rect 16091 4910 16101 5088
rect 16279 4910 16289 5088
rect 16091 4905 16289 4910
rect 19091 5088 19289 5093
rect 19091 4910 19101 5088
rect 19279 4910 19289 5088
rect 19091 4905 19289 4910
rect 21240 4540 21250 7514
rect 21417 4540 21427 7514
rect 21240 4535 21427 4540
rect 34644 7013 34708 8272
rect 35014 8219 35024 8272
rect 35088 8219 35098 8283
rect 35014 8214 35098 8219
rect 40011 8121 40269 8135
rect 38558 8038 39142 8083
rect 36007 7881 36581 7896
rect 36007 7814 36301 7881
rect 36532 7814 36581 7881
rect 38558 7892 38575 8038
rect 38645 7913 39142 8038
rect 40011 7933 40100 8121
rect 40181 7933 40269 8121
rect 40011 7913 40269 7933
rect 38645 7892 40721 7913
rect 38558 7843 40721 7892
rect 36007 7800 36581 7814
rect 35008 7223 35127 7253
rect 35008 7159 35028 7223
rect 35092 7188 35127 7223
rect 36007 7188 36103 7800
rect 38902 7673 40721 7843
rect 38558 7563 38659 7568
rect 38558 7375 38568 7563
rect 38649 7375 38659 7563
rect 38558 7370 38659 7375
rect 36338 7337 36971 7349
rect 36338 7275 36362 7337
rect 36531 7275 36971 7337
rect 36338 7253 36971 7275
rect 37067 7253 37077 7349
rect 35092 7159 36103 7188
rect 35008 7124 36103 7159
rect 35008 7123 35127 7124
rect 34644 6959 35091 7013
rect 34644 6954 35101 6959
rect 34644 6949 35027 6954
rect 34644 5623 34708 6949
rect 35017 6890 35027 6949
rect 35091 6890 35101 6954
rect 35017 6885 35101 6890
rect 36007 6816 36103 7124
rect 36007 6800 36442 6816
rect 36007 6795 36447 6800
rect 36007 6721 36352 6795
rect 36437 6721 36447 6795
rect 38902 6765 39142 7673
rect 40077 7576 40178 7581
rect 40077 7388 40087 7576
rect 40168 7388 40178 7576
rect 40077 7383 40178 7388
rect 40481 7170 40721 7673
rect 42592 7232 45933 7237
rect 40481 6930 40801 7170
rect 41264 6930 41274 7170
rect 42592 7143 42602 7232
rect 45923 7143 45933 7232
rect 42592 7138 45933 7143
rect 40481 6797 40721 6930
rect 36007 6720 36447 6721
rect 36342 6716 36447 6720
rect 35000 5885 35108 5908
rect 35000 5821 35027 5885
rect 35091 5866 35108 5885
rect 35091 5821 35644 5866
rect 35000 5802 35644 5821
rect 35000 5796 35108 5802
rect 35580 5714 35644 5802
rect 36346 5727 36442 6716
rect 38541 6707 39142 6765
rect 38541 6582 38571 6707
rect 38649 6582 39142 6707
rect 38541 6525 39142 6582
rect 40076 6785 40721 6797
rect 40076 6597 40092 6785
rect 40173 6597 40721 6785
rect 40076 6557 40721 6597
rect 36961 6265 37077 6270
rect 36961 6169 36971 6265
rect 37067 6169 37077 6265
rect 36961 6164 37077 6169
rect 38553 6232 38654 6237
rect 38553 6044 38563 6232
rect 38644 6044 38654 6232
rect 38553 6039 38654 6044
rect 35934 5714 36442 5727
rect 35580 5707 36442 5714
rect 35580 5650 35970 5707
rect 35934 5644 35970 5650
rect 36149 5644 36442 5707
rect 35934 5631 36442 5644
rect 34644 5567 35088 5623
rect 34644 5562 35098 5567
rect 34644 5559 35024 5562
rect 4669 4366 4867 4371
rect 4669 4188 4679 4366
rect 4857 4188 4867 4366
rect 34644 4288 34708 5559
rect 35014 5498 35024 5559
rect 35088 5498 35098 5562
rect 35014 5493 35098 5498
rect 35934 4727 36030 5631
rect 38902 5395 39142 6525
rect 40082 6229 40183 6234
rect 40082 6041 40092 6229
rect 40173 6041 40183 6229
rect 40082 6036 40183 6041
rect 40481 5416 40721 6557
rect 47463 5800 47719 5805
rect 47463 5564 47473 5800
rect 47709 5564 62907 5800
rect 47463 5559 47719 5564
rect 38561 5322 39142 5395
rect 38561 5187 38574 5322
rect 38648 5187 39142 5322
rect 36498 5162 36971 5177
rect 36498 5092 36514 5162
rect 36734 5092 36971 5162
rect 36498 5081 36971 5092
rect 37067 5081 37077 5177
rect 38561 5155 39142 5187
rect 40088 5405 40721 5416
rect 40088 5217 40109 5405
rect 40190 5217 40721 5405
rect 40088 5176 40721 5217
rect 38552 4879 38653 4884
rect 35934 4633 36445 4727
rect 38552 4691 38562 4879
rect 38643 4691 38653 4879
rect 38552 4686 38653 4691
rect 35934 4631 36537 4633
rect 36349 4613 36537 4631
rect 36349 4555 36364 4613
rect 36509 4555 36537 4613
rect 36349 4537 36537 4555
rect 35014 4492 35119 4516
rect 35014 4428 35035 4492
rect 35099 4480 35119 4492
rect 36349 4480 36445 4537
rect 35099 4428 36445 4480
rect 35014 4416 36445 4428
rect 35014 4403 35119 4416
rect 34644 4224 35088 4288
rect 4669 4183 4867 4188
rect 35014 4192 35088 4224
rect 35014 4187 35098 4192
rect 35014 4123 35024 4187
rect 35088 4123 35098 4187
rect 35014 4118 35098 4123
rect 36349 3627 36445 4416
rect 36962 4089 37078 4094
rect 36962 3993 36972 4089
rect 37068 3993 37078 4089
rect 36962 3988 37078 3993
rect 38902 3986 39142 5155
rect 40082 4857 40183 4862
rect 40082 4669 40092 4857
rect 40173 4669 40183 4857
rect 40082 4664 40183 4669
rect 40481 4267 40721 5176
rect 38548 3934 39142 3986
rect 38548 3781 38572 3934
rect 38651 3818 39142 3934
rect 40015 4026 40255 4037
rect 40015 3838 40099 4026
rect 40180 3838 40255 4026
rect 40015 3818 40255 3838
rect 40481 4027 40799 4267
rect 41262 4027 41272 4267
rect 42589 4233 45969 4238
rect 42589 4144 42599 4233
rect 45959 4144 45969 4233
rect 42589 4139 45969 4144
rect 40481 3818 40721 4027
rect 38651 3781 40721 3818
rect 38548 3746 40721 3781
rect 36349 3536 36448 3627
rect 38902 3578 40721 3746
rect 36349 3531 36496 3536
rect 36349 3459 36359 3531
rect 36486 3459 36496 3531
rect 36349 3454 36496 3459
rect 38555 3479 38656 3484
rect 35005 3122 35116 3144
rect 35005 3058 35031 3122
rect 35095 3113 35116 3122
rect 36359 3113 36423 3454
rect 38555 3291 38565 3479
rect 38646 3291 38656 3479
rect 38555 3286 38656 3291
rect 40079 3473 40180 3478
rect 40079 3285 40089 3473
rect 40170 3285 40180 3473
rect 40079 3280 40180 3285
rect 35095 3058 36423 3113
rect 35005 3049 36423 3058
rect 35005 3029 35116 3049
rect 40481 3045 40721 3578
rect 18 2773 200 2778
rect 18 359 28 2773
rect 190 359 200 2773
rect 12197 2773 12395 2778
rect 12197 2595 12207 2773
rect 12385 2595 12395 2773
rect 12197 2590 12395 2595
rect 4669 2366 4867 2371
rect 4669 2188 4679 2366
rect 4857 2188 4867 2366
rect 4669 2183 4867 2188
rect 36043 2214 36151 2236
rect 36043 2150 36066 2214
rect 36130 2150 36151 2214
rect 21233 2139 21429 2144
rect 21233 1288 21243 2139
rect 21419 1288 21429 2139
rect 36043 2124 36151 2150
rect 36888 1765 36898 1852
rect 21233 1283 21429 1288
rect 34644 1701 36898 1765
rect 34644 1396 34708 1701
rect 35459 1591 35583 1623
rect 36888 1616 36898 1701
rect 37140 1616 37150 1852
rect 35459 1527 35489 1591
rect 35553 1527 35583 1591
rect 35459 1496 35583 1527
rect 36604 1529 36720 1558
rect 36604 1465 36631 1529
rect 36695 1465 36720 1529
rect 36604 1437 36720 1465
rect 34644 1348 35088 1396
rect 34644 1343 35098 1348
rect 34644 1332 35024 1343
rect 18 354 200 359
rect 312 232 21117 237
rect 312 67 322 232
rect 21107 67 21117 232
rect 312 62 21117 67
rect 34644 73 34708 1332
rect 35014 1279 35024 1332
rect 35088 1279 35098 1343
rect 35014 1274 35098 1279
rect 40011 1181 40269 1195
rect 38558 1098 39142 1143
rect 36007 941 36581 956
rect 36007 874 36301 941
rect 36532 874 36581 941
rect 38558 952 38575 1098
rect 38645 973 39142 1098
rect 40011 993 40100 1181
rect 40181 993 40269 1181
rect 40011 973 40269 993
rect 38645 952 40721 973
rect 38558 903 40721 952
rect 36007 860 36581 874
rect 35008 283 35127 313
rect 35008 219 35028 283
rect 35092 248 35127 283
rect 36007 248 36103 860
rect 38902 733 40721 903
rect 38558 623 38659 628
rect 38558 435 38568 623
rect 38649 435 38659 623
rect 38558 430 38659 435
rect 36338 397 36971 409
rect 36338 335 36362 397
rect 36531 335 36971 397
rect 36338 313 36971 335
rect 37067 313 37077 409
rect 35092 219 36103 248
rect 35008 184 36103 219
rect 35008 183 35127 184
rect 34644 19 35091 73
rect 34644 14 35101 19
rect 34644 9 35027 14
rect 34644 -1317 34708 9
rect 35017 -50 35027 9
rect 35091 -50 35101 14
rect 35017 -55 35101 -50
rect 36007 -124 36103 184
rect 36007 -140 36442 -124
rect 36007 -145 36447 -140
rect 36007 -219 36352 -145
rect 36437 -219 36447 -145
rect 38902 -175 39142 733
rect 40077 636 40178 641
rect 40077 448 40087 636
rect 40168 448 40178 636
rect 40077 443 40178 448
rect 40481 230 40721 733
rect 42589 309 45940 314
rect 40481 -10 40801 230
rect 41264 -10 41274 230
rect 42589 199 42599 309
rect 45930 199 45940 309
rect 42589 194 45940 199
rect 40481 -143 40721 -10
rect 36007 -220 36447 -219
rect 36342 -224 36447 -220
rect 35000 -1055 35108 -1032
rect 35000 -1119 35027 -1055
rect 35091 -1074 35108 -1055
rect 35091 -1119 35644 -1074
rect 35000 -1138 35644 -1119
rect 35000 -1144 35108 -1138
rect 35580 -1226 35644 -1138
rect 36346 -1213 36442 -224
rect 38541 -233 39142 -175
rect 38541 -358 38571 -233
rect 38649 -358 39142 -233
rect 38541 -415 39142 -358
rect 40076 -155 40721 -143
rect 40076 -343 40092 -155
rect 40173 -343 40721 -155
rect 40076 -383 40721 -343
rect 36961 -675 37077 -670
rect 36961 -771 36971 -675
rect 37067 -771 37077 -675
rect 36961 -776 37077 -771
rect 38553 -708 38654 -703
rect 38553 -896 38563 -708
rect 38644 -896 38654 -708
rect 38553 -901 38654 -896
rect 35934 -1226 36442 -1213
rect 35580 -1233 36442 -1226
rect 35580 -1290 35970 -1233
rect 35934 -1296 35970 -1290
rect 36149 -1296 36442 -1233
rect 35934 -1309 36442 -1296
rect 34644 -1373 35088 -1317
rect 34644 -1378 35098 -1373
rect 34644 -1381 35024 -1378
rect 34644 -2652 34708 -1381
rect 35014 -1442 35024 -1381
rect 35088 -1442 35098 -1378
rect 35014 -1447 35098 -1442
rect 35934 -2213 36030 -1309
rect 38902 -1545 39142 -415
rect 40082 -711 40183 -706
rect 40082 -899 40092 -711
rect 40173 -899 40183 -711
rect 40082 -904 40183 -899
rect 40481 -1524 40721 -383
rect 47479 -1140 47735 -1135
rect 47479 -1376 47489 -1140
rect 47725 -1376 62907 -1140
rect 47479 -1381 47735 -1376
rect 38561 -1618 39142 -1545
rect 38561 -1753 38574 -1618
rect 38648 -1753 39142 -1618
rect 36498 -1778 36971 -1763
rect 36498 -1848 36514 -1778
rect 36734 -1848 36971 -1778
rect 36498 -1859 36971 -1848
rect 37067 -1859 37077 -1763
rect 38561 -1785 39142 -1753
rect 40088 -1535 40721 -1524
rect 40088 -1723 40109 -1535
rect 40190 -1723 40721 -1535
rect 40088 -1764 40721 -1723
rect 38552 -2061 38653 -2056
rect 35934 -2307 36445 -2213
rect 38552 -2249 38562 -2061
rect 38643 -2249 38653 -2061
rect 38552 -2254 38653 -2249
rect 35934 -2309 36537 -2307
rect 36349 -2327 36537 -2309
rect 36349 -2385 36364 -2327
rect 36509 -2385 36537 -2327
rect 36349 -2403 36537 -2385
rect 35014 -2448 35119 -2424
rect 35014 -2512 35035 -2448
rect 35099 -2460 35119 -2448
rect 36349 -2460 36445 -2403
rect 35099 -2512 36445 -2460
rect 35014 -2524 36445 -2512
rect 35014 -2537 35119 -2524
rect 34644 -2716 35088 -2652
rect 35014 -2748 35088 -2716
rect 35014 -2753 35098 -2748
rect 35014 -2817 35024 -2753
rect 35088 -2817 35098 -2753
rect 35014 -2822 35098 -2817
rect 36349 -3313 36445 -2524
rect 36962 -2851 37078 -2846
rect 36962 -2947 36972 -2851
rect 37068 -2947 37078 -2851
rect 36962 -2952 37078 -2947
rect 38902 -2954 39142 -1785
rect 40082 -2083 40183 -2078
rect 40082 -2271 40092 -2083
rect 40173 -2271 40183 -2083
rect 40082 -2276 40183 -2271
rect 40481 -2673 40721 -1764
rect 38548 -3006 39142 -2954
rect 38548 -3159 38572 -3006
rect 38651 -3122 39142 -3006
rect 40015 -2914 40255 -2903
rect 40015 -3102 40099 -2914
rect 40180 -3102 40255 -2914
rect 40015 -3122 40255 -3102
rect 40481 -2913 40799 -2673
rect 41262 -2913 41272 -2673
rect 42577 -2708 45943 -2703
rect 42577 -2796 42587 -2708
rect 45933 -2796 45943 -2708
rect 42577 -2801 45943 -2796
rect 40481 -3122 40721 -2913
rect 38651 -3159 40721 -3122
rect 38548 -3194 40721 -3159
rect 36349 -3404 36448 -3313
rect 38902 -3362 40721 -3194
rect 36349 -3409 36496 -3404
rect 36349 -3481 36359 -3409
rect 36486 -3481 36496 -3409
rect 36349 -3486 36496 -3481
rect 38555 -3461 38656 -3456
rect -1926 -3573 21202 -3509
rect 21266 -3573 21276 -3509
rect 35005 -3818 35116 -3796
rect 35005 -3882 35031 -3818
rect 35095 -3827 35116 -3818
rect 36359 -3827 36423 -3486
rect 38555 -3649 38565 -3461
rect 38646 -3649 38656 -3461
rect 38555 -3654 38656 -3649
rect 40079 -3467 40180 -3462
rect 40079 -3655 40089 -3467
rect 40170 -3655 40180 -3467
rect 40079 -3660 40180 -3655
rect 35095 -3882 36423 -3827
rect 35005 -3891 36423 -3882
rect 35005 -3911 35116 -3891
rect 40481 -3895 40721 -3362
rect -2212 -4045 21202 -3981
rect 21266 -4045 21276 -3981
rect -2598 -4580 21202 -4516
rect 21266 -4580 21276 -4516
rect -2885 -5043 21202 -4979
rect 21266 -5043 21276 -4979
rect -3605 -6822 -3493 -6817
rect -3605 -10130 -3595 -6822
rect -3503 -10130 -3493 -6822
rect -3605 -10135 -3493 -10130
rect -610 -6825 -476 -6820
rect -610 -10140 -600 -6825
rect -486 -10140 -476 -6825
rect -610 -10145 -476 -10140
rect -2189 -12082 -1933 -12077
rect -2189 -12318 -2179 -12082
rect -1943 -12318 -1933 -12082
rect -2189 -12323 -1933 -12318
rect -2179 -18865 -1943 -12323
rect -2179 -19101 -885 -18865
rect -1121 -24022 -885 -19101
<< via3 >>
rect -16849 73398 -16748 76723
rect -13848 73404 -13747 76729
rect 11143 73392 11271 76732
rect 14144 73405 14272 76745
rect -16664 71738 -16600 71802
rect -15486 71734 -15422 71798
rect -15269 71741 -15205 71805
rect -14135 71738 -14071 71802
rect -16554 70234 -16490 70298
rect -15440 70220 -15376 70284
rect -15227 70221 -15163 70285
rect -14063 70221 -13999 70285
rect 36631 69270 36695 69334
rect 36065 68676 36131 68742
rect -15963 68105 -15890 68261
rect -15422 68166 -15358 68515
rect -14879 68108 -14806 68264
rect 35476 68016 35542 68082
rect -16577 67549 -16513 67613
rect -15422 67543 -15358 67607
rect -14304 67554 -14240 67618
rect -13096 66705 -13032 66769
rect -8073 66705 -8009 66769
rect -12315 66382 -12251 66446
rect -7266 66382 -7202 66446
rect -11305 65949 -11241 66013
rect -2673 65949 -2609 66013
rect -10536 65696 -10472 65760
rect -1866 65696 -1802 65760
rect -8073 65265 -8009 65329
rect -2673 65265 -2609 65329
rect -7266 65012 -7202 65076
rect -1866 65012 -1802 65076
rect 17430 64169 17496 64743
rect 23958 64169 24024 64743
rect 31574 64169 31640 64743
rect -11071 63205 -10737 63557
rect -10187 63338 -10123 63402
rect -9884 63338 -9442 63402
rect -8073 63340 -7631 63404
rect -6278 63336 -5836 63400
rect -4479 63334 -4037 63398
rect -2688 63338 -2246 63402
rect -886 63334 -444 63398
rect -6939 62966 -6699 63206
rect 757 62992 1287 63232
rect 17975 62166 18041 62740
rect 19063 62166 19129 62740
rect 21239 62166 21305 62740
rect 22327 62166 22393 62740
rect 23415 62166 23481 62740
rect 24503 62166 24569 62740
rect 25591 62166 25657 62740
rect 26679 62166 26745 62740
rect 28855 62166 28921 62740
rect 29943 62166 30009 62740
rect 31031 62166 31097 62740
rect -8557 54531 -8493 54595
rect -6866 54532 -6802 54596
rect -5161 54531 -5097 54595
rect -3365 54531 -3301 54595
rect -1536 54531 -1472 54595
rect -9704 54339 -9462 54403
rect -7909 54338 -7667 54402
rect -6109 54340 -5867 54404
rect -4311 54339 -4069 54403
rect -2513 54340 -2271 54404
rect -710 54339 -468 54403
rect 176 54340 240 54404
rect -7265 54019 -7201 54083
rect -1865 54019 -1801 54083
rect -8073 53766 -8009 53830
rect -2673 53766 -2609 53830
rect -10536 53338 -10472 53402
rect -1865 53338 -1801 53402
rect -11305 53082 -11241 53146
rect -2673 53082 -2609 53146
rect 347 53121 519 60827
rect 5410 58752 5588 58930
rect 2047 57297 2225 57475
rect 4047 57297 4225 57475
rect 5410 55752 5588 55930
rect 4007 53001 4185 53179
rect -12315 52649 -12251 52713
rect -7265 52649 -7201 52713
rect -13096 52326 -13032 52390
rect -8073 52326 -8009 52390
rect 7725 51858 7903 52036
rect -8854 51014 -8770 51249
rect -7722 51183 -7658 51247
rect -5688 50883 -3888 51066
rect -3362 50896 -2536 51074
rect -1655 50886 -765 51064
rect -8874 50378 -8780 50791
rect -8480 50377 -8416 50441
rect -8480 50008 -8416 50072
rect -27070 49656 -26726 49720
rect -7722 49360 -7658 49424
rect -25984 49114 -25640 49178
rect -5932 47776 -5748 50720
rect -78 47752 121 50774
rect 10177 47617 10551 60836
rect 17430 60169 17496 60743
rect 18518 60169 18584 60743
rect 19606 60169 19672 60743
rect 20694 60169 20760 60743
rect 21782 60169 21848 60743
rect 22870 60169 22936 60743
rect 23958 60169 24024 60743
rect 25046 60169 25112 60743
rect 26134 60169 26200 60743
rect 27222 60169 27288 60743
rect 28310 60169 28376 60743
rect 29398 60169 29464 60743
rect 30486 60169 30552 60743
rect 31574 60169 31640 60743
rect 17975 58166 18041 58740
rect 19063 58166 19129 58740
rect 20151 58166 20217 58740
rect 21239 58166 21305 58740
rect 22327 58166 22393 58740
rect 23415 58166 23481 58740
rect 24503 58166 24569 58740
rect 25591 58166 25657 58740
rect 26679 58166 26745 58740
rect 27767 58166 27833 58740
rect 28855 58166 28921 58740
rect 29943 58166 30009 58740
rect 31031 58166 31097 58740
rect 17430 56169 17496 56743
rect 18518 56169 18584 56743
rect 19606 56169 19672 56743
rect 20694 56169 20760 56743
rect 21782 56169 21848 56743
rect 22870 56169 22936 56743
rect 23958 56169 24024 56743
rect 25046 56169 25112 56743
rect 26134 56169 26200 56743
rect 27222 56169 27288 56743
rect 28310 56169 28376 56743
rect 29398 56169 29464 56743
rect 30486 56169 30552 56743
rect 31574 56169 31640 56743
rect 17975 54166 18041 54740
rect 19063 54166 19129 54740
rect 20151 54166 20217 54740
rect 21239 54166 21305 54740
rect 22327 54166 22393 54740
rect 23415 54166 23481 54740
rect 24503 54166 24569 54740
rect 25591 54166 25657 54740
rect 26679 54166 26745 54740
rect 27767 54166 27833 54740
rect 28855 54166 28921 54740
rect 29943 54166 30009 54740
rect 31031 54166 31097 54740
rect 17430 52169 17496 52743
rect 18518 52169 18584 52743
rect 19606 52169 19672 52743
rect 20694 52169 20760 52743
rect 21782 52169 21848 52743
rect 22870 52169 22936 52743
rect 23958 52169 24024 52743
rect 25046 52169 25112 52743
rect 26134 52169 26200 52743
rect 27222 52169 27288 52743
rect 28310 52169 28376 52743
rect 29398 52169 29464 52743
rect 30486 52169 30552 52743
rect 31574 52169 31640 52743
rect 17975 50166 18041 50740
rect 20151 50166 20217 50740
rect 21239 50166 21305 50740
rect 23415 50166 23481 50740
rect 24503 50166 24569 50740
rect 25591 50166 25657 50740
rect 27767 50166 27833 50740
rect 28855 50166 28921 50740
rect 31031 50166 31097 50740
rect 17430 48169 17496 48743
rect 18518 48169 18584 48743
rect 19606 48169 19672 48743
rect 20694 48169 20760 48743
rect 21782 48169 21848 48743
rect 22870 48169 22936 48743
rect 23958 48169 24024 48743
rect 29398 48169 29464 48743
rect 30486 48169 30552 48743
rect 31574 48169 31640 48743
rect -11361 47192 -11297 47256
rect -6411 47192 -6347 47256
rect -27087 42779 -26990 43313
rect -27082 41002 -26995 42169
rect -27077 39476 -26990 40643
rect -31812 38827 -31748 39166
rect -31811 38141 -31747 38613
rect -29614 38349 -29150 38413
rect -27082 38232 -26998 39120
rect -10487 46569 -10423 46633
rect -6411 46569 -6347 46633
rect -13469 42997 -13405 43061
rect -9208 42997 -9144 43061
rect -12693 42334 -12629 42398
rect -10069 42334 -10005 42398
rect -21475 42099 -21411 42163
rect -5924 39819 -5722 46274
rect 17975 46166 18041 46740
rect 19063 46166 19129 46740
rect 20151 46166 20217 46740
rect 21239 46166 21305 46740
rect 22327 46166 22393 46740
rect 24503 46166 24569 46740
rect 25591 46166 25657 46740
rect 26679 46166 26745 46740
rect 27767 46166 27833 46740
rect 28855 46166 28921 46740
rect 29943 46166 30009 46740
rect 31031 46166 31097 46740
rect -4101 45129 -3923 45307
rect -1482 44281 -1304 44459
rect 344 44318 558 45844
rect 2132 44330 2310 44508
rect 4132 44330 4310 44508
rect 6132 44330 6310 44508
rect 8132 44330 8310 44508
rect 352 39855 512 41383
rect 10180 39867 10551 46128
rect 18245 45684 18309 45748
rect 18791 45684 18855 45748
rect 19337 45675 19401 45739
rect 19882 45674 19946 45738
rect 21517 45684 21581 45748
rect 22051 45671 22115 45735
rect 22598 45677 22662 45741
rect 23143 45677 23207 45741
rect 25863 45674 25927 45738
rect 26406 45678 26470 45742
rect 26948 45672 27012 45736
rect 27505 45663 27569 45727
rect 29129 45674 29193 45738
rect 29673 45667 29737 45731
rect 30223 45671 30287 45735
rect 30756 45671 30820 45735
rect 18791 45008 18855 45072
rect 44754 45007 45306 45074
rect 25863 44827 25927 44891
rect 18245 44637 18309 44701
rect 26406 44462 26470 44526
rect 41516 44462 41874 44527
rect 22598 43858 22662 43922
rect 44766 43854 45293 43925
rect 30756 43677 30820 43741
rect 23143 43487 23207 43551
rect 30222 43311 30286 43375
rect 41514 43312 41872 43377
rect 19882 41318 19946 41382
rect 44756 41312 45283 41383
rect 26948 41137 27012 41201
rect 19337 40947 19401 41011
rect 27505 40772 27569 40836
rect 41432 40771 41790 40836
rect 21517 40048 21581 40112
rect 44756 40042 45283 40113
rect 29673 39867 29737 39931
rect -5684 39666 -148 39846
rect 22051 39677 22115 39741
rect -29652 37259 -29143 37323
rect -27079 36465 -26995 37353
rect -27077 34985 -26996 36160
rect -18883 36124 -18807 39537
rect 29129 39502 29193 39566
rect 41430 39502 41788 39567
rect -11713 38726 -11649 38790
rect -4713 38726 -4649 38790
rect -10905 38383 -10841 38447
rect -4123 38383 -4059 38447
rect 2513 38642 2595 38881
rect -7722 37835 -7658 37899
rect -2398 37835 -2334 37899
rect -760 37835 -696 37899
rect 1473 37835 1537 37899
rect -8480 37307 -8416 37371
rect -2815 37307 -2751 37371
rect -760 37306 -696 37370
rect 2515 37996 2614 38420
rect 13831 38372 13895 38436
rect 18245 38372 18309 38436
rect 25863 38354 25927 38418
rect 32414 38354 32478 38418
rect 14586 37797 14650 37861
rect 18791 37797 18855 37861
rect 26406 37774 26470 37838
rect 31824 37774 31888 37838
rect 1996 37306 2060 37370
rect 15230 37246 15294 37310
rect 19337 37246 19401 37310
rect 30756 37165 30820 37229
rect 31231 37165 31295 37229
rect 2168 36898 2232 37149
rect 2169 36250 2233 36668
rect 15990 36664 16054 36728
rect 19882 36664 19946 36728
rect 30222 36529 30286 36593
rect 30584 36529 30648 36593
rect 3582 36030 3811 36094
rect -9208 35877 -9144 35941
rect 5055 36018 5351 36104
rect 5574 36027 5801 36097
rect 3121 35553 3240 35672
rect 6936 36020 7157 36089
rect 9575 36023 9802 36091
rect 16721 35986 16785 36050
rect 21517 35986 21581 36050
rect 29673 35906 29737 35970
rect 29990 35906 30054 35970
rect 7503 35522 7622 35641
rect 9070 35531 9189 35650
rect -10069 35287 -10005 35351
rect 17412 35279 17476 35343
rect 22051 35279 22115 35343
rect 29129 35194 29193 35258
rect 29407 35194 29471 35258
rect -27079 33498 -27000 34691
rect -13395 34612 -13331 34676
rect 18252 34519 18316 34583
rect 22598 34519 22662 34583
rect 26948 34458 27012 34522
rect 28828 34458 28892 34522
rect -4713 34131 -4649 34195
rect -4123 33786 -4059 33850
rect 27505 33749 27569 33813
rect 28315 33749 28379 33813
rect 19255 33682 19319 33746
rect 23143 33682 23207 33746
rect -21518 33487 -21454 33551
rect -15139 33115 -15075 33179
rect -27084 32365 -27005 32899
rect 7965 31747 8029 31811
rect 11347 31327 11411 31391
rect 13831 31327 13895 31391
rect 4354 30368 4418 30432
rect 8328 30373 8392 30437
rect 11966 30708 12030 30772
rect 14586 30708 14650 30772
rect 3326 30241 3390 30305
rect -3918 29688 -3854 29752
rect -5279 29265 -5215 29329
rect 16721 29688 16785 29752
rect 17412 29265 17476 29329
rect 10633 28740 10697 28804
rect 11966 28740 12030 28804
rect -17635 27516 -17507 27644
rect -15712 27645 -15613 28098
rect -12389 27670 -12316 28076
rect -5279 27468 -5215 27532
rect -12394 27198 -12297 27427
rect -3918 26791 -3854 26855
rect -38190 26514 -34856 26611
rect -17635 26287 -17507 26415
rect -15725 26044 -15636 26281
rect -12396 26057 -12301 26486
rect 11347 26286 11411 26350
rect 11837 26286 11901 26350
rect 13850 25945 13914 26009
rect 25879 25945 25943 26009
rect -19088 25571 -18855 25804
rect -25449 25175 -25369 25482
rect -11324 25600 -11260 25664
rect 13266 25534 13330 25598
rect 26463 25534 26527 25598
rect -25452 24714 -25365 24945
rect -17635 24874 -17507 25002
rect -11977 24808 -11913 24872
rect 7601 24784 7665 24848
rect 15230 24784 15294 24848
rect -12393 24458 -12328 24712
rect -12398 24003 -12316 24239
rect 5715 24186 5783 24594
rect 7266 24529 7330 24593
rect 8129 24466 8193 24530
rect 15990 24466 16054 24530
rect 11080 24138 11144 24202
rect -11324 23823 -11260 23887
rect 7266 23823 7330 23887
rect 19255 23823 19319 23887
rect -17635 23645 -17507 23773
rect -38182 23503 -34852 23605
rect -15725 23405 -15658 23637
rect -11977 23454 -11913 23518
rect 18252 23454 18316 23518
rect -12389 22857 -12319 23277
rect 8787 23246 8943 23356
rect 42856 24065 46190 24174
rect 36066 23954 36130 24018
rect 35152 23802 35216 23866
rect 37819 23492 37892 23611
rect 39346 23493 39420 23714
rect 4780 22919 5243 23159
rect 12588 23146 12652 23210
rect 27111 23146 27175 23210
rect 5718 22999 5782 23063
rect 37819 22946 37905 23194
rect 39335 22952 39421 23200
rect 11476 22851 11540 22915
rect 11837 22852 11901 22916
rect -16599 22660 -16535 22724
rect 8129 22660 8193 22724
rect -12391 22399 -12323 22624
rect 7601 22209 7665 22273
rect 36914 22579 37156 22815
rect 37826 22151 37896 22280
rect 39346 22167 39420 22388
rect 12072 21591 12136 21655
rect 27657 21591 27721 21655
rect 37814 21621 37899 21823
rect 35152 21521 35216 21585
rect 39341 21586 39427 21834
rect 35477 21315 35541 21379
rect 42854 21069 46188 21178
rect -38168 18987 -34861 19065
rect -38174 15987 -34852 16075
rect 12936 20963 13000 21027
rect -25452 17627 -25387 17922
rect -25450 17169 -25378 17404
rect -16599 20587 -16535 20651
rect 11080 20270 11144 20334
rect -12355 17904 -12291 17968
rect -10416 17093 -10352 17157
rect -25517 14157 -25444 14446
rect -18223 14009 -18159 14073
rect -25518 13690 -25446 13925
rect -13941 10117 -13877 10181
rect -10970 10159 -10906 10223
rect 11476 19739 11540 19803
rect -2815 19449 -2751 19513
rect -5279 18979 -5215 19043
rect -3918 18979 -3854 19043
rect -5786 15644 -5722 15708
rect -4902 14236 -4832 14446
rect -6162 10758 -5937 10833
rect -6167 9513 -5929 9592
rect 23689 19318 23753 19382
rect -2398 19148 -2334 19212
rect 14686 19214 14750 19278
rect 4857 19027 5194 19173
rect 10232 18994 10296 19058
rect 20971 18998 21035 19062
rect -1504 18846 -1440 18910
rect -1133 18587 -1069 18651
rect 8280 18654 8344 18718
rect 12930 18624 12994 18688
rect 14115 18507 14179 18571
rect 25614 18507 25678 18571
rect -680 18248 -616 18312
rect -284 17967 -220 18031
rect -3211 17624 -2748 17864
rect 14368 17699 14432 17763
rect 25361 17700 25425 17764
rect 981 17461 1045 17525
rect 14689 17485 14753 17549
rect 23689 17488 23753 17552
rect 4295 17225 4359 17289
rect 6227 17225 6291 17289
rect 12956 17019 13020 17083
rect 251 16238 11139 16446
rect -3509 16141 -3445 16205
rect -3928 15390 -3864 15454
rect -3144 14719 -3061 14998
rect -3509 14580 -3445 14644
rect -3185 8643 -3121 8707
rect -1808 12726 -1725 13133
rect -1759 11140 -1693 11529
rect -7214 7003 -6751 7243
rect -25521 6408 -25446 6669
rect -3184 6585 -3120 6649
rect -18251 6239 -18187 6303
rect -25522 5929 -25447 6174
rect -4907 5950 -4841 6163
rect -3928 5978 -3864 6042
rect -3193 5296 -3110 5577
rect -3509 5169 -3445 5233
rect -1759 9532 -1695 9930
rect 5478 14421 5656 14599
rect 14685 15689 14749 15753
rect 23686 15724 23750 15788
rect 20928 15432 20992 15496
rect 12973 15164 13037 15228
rect 14685 13901 14749 13965
rect 23686 13933 23750 13997
rect 13003 13464 13067 13528
rect 14115 13107 14179 13171
rect 14368 12299 14432 12363
rect 4630 11802 4808 11980
rect 14702 12116 14766 12180
rect 23691 12126 23755 12190
rect 20985 11842 21049 11906
rect 13001 11612 13065 11676
rect 6483 10356 11218 10537
rect 14691 10319 14755 10383
rect 23691 10316 23755 10380
rect 372 10003 1812 10144
rect 5727 9990 11722 10135
rect 13876 9993 21118 10150
rect -1758 7930 -1690 8330
rect 29 5570 212 9830
rect 36066 9090 36130 9154
rect 4679 8188 4857 8366
rect 17646 8273 17824 8451
rect 36898 8556 37140 8792
rect 35489 8467 35553 8531
rect 36631 8405 36695 8469
rect 4679 6188 4857 6366
rect 13350 6313 13528 6491
rect 17646 6273 17824 6451
rect 16101 4910 16279 5088
rect 19101 4910 19279 5088
rect 21250 4540 21417 7514
rect 35028 7159 35092 7223
rect 38568 7375 38649 7563
rect 36971 7253 37067 7349
rect 40087 7388 40168 7576
rect 40801 6930 41264 7170
rect 42602 7143 45923 7232
rect 35027 5821 35091 5885
rect 36971 6169 37067 6265
rect 38563 6044 38644 6232
rect 4679 4188 4857 4366
rect 40092 6041 40173 6229
rect 36971 5081 37067 5177
rect 38562 4691 38643 4879
rect 35035 4428 35099 4492
rect 36972 3993 37068 4089
rect 40092 4669 40173 4857
rect 40799 4027 41262 4267
rect 42599 4144 45959 4233
rect 35031 3058 35095 3122
rect 38565 3291 38646 3479
rect 40089 3285 40170 3473
rect 28 359 190 2773
rect 12207 2595 12385 2773
rect 4679 2188 4857 2366
rect 36066 2150 36130 2214
rect 21243 1288 21419 2139
rect 36898 1616 37140 1852
rect 35489 1527 35553 1591
rect 36631 1465 36695 1529
rect 322 67 21107 232
rect 35028 219 35092 283
rect 38568 435 38649 623
rect 36971 313 37067 409
rect 40087 448 40168 636
rect 40801 -10 41264 230
rect 42599 199 45930 309
rect 35027 -1119 35091 -1055
rect 36971 -771 37067 -675
rect 38563 -896 38644 -708
rect 40092 -899 40173 -711
rect 36971 -1859 37067 -1763
rect 38562 -2249 38643 -2061
rect 35035 -2512 35099 -2448
rect 36972 -2947 37068 -2851
rect 40092 -2271 40173 -2083
rect 40799 -2913 41262 -2673
rect 42587 -2796 45933 -2708
rect 21202 -3573 21266 -3509
rect 35031 -3882 35095 -3818
rect 38565 -3649 38646 -3461
rect 40089 -3655 40170 -3467
rect 21202 -4045 21266 -3981
rect 21202 -4580 21266 -4516
rect 21202 -5043 21266 -4979
rect -3595 -10130 -3503 -6822
rect -600 -10140 -486 -6825
<< metal4 >>
rect -57093 86442 -55093 88442
rect -53093 86442 -43285 88442
rect -42665 86442 -35285 88442
rect -34665 86442 -27285 88442
rect -26665 86442 -19285 88442
rect -18665 86442 -11285 88442
rect -10665 86442 -3285 88442
rect -2665 86442 4715 88442
rect 5335 86442 12715 88442
rect 13335 86442 20715 88442
rect 21335 86442 28715 88442
rect 29335 86442 36715 88442
rect 37335 86442 44715 88442
rect 45335 86442 54907 88442
rect 56907 86442 62907 88442
rect -57093 82442 -51093 84442
rect -49093 82442 -39285 84442
rect -38665 82442 -31285 84442
rect -30665 82442 -23285 84442
rect -22665 82442 -15285 84442
rect -14665 82442 -7285 84442
rect -6665 82442 715 84442
rect 1335 82442 8715 84442
rect 9335 82442 16715 84442
rect 17335 82442 24715 84442
rect 25335 82442 32715 84442
rect 33335 82442 40715 84442
rect 41335 82442 48715 84442
rect 49335 82442 58907 84442
rect 60907 82442 62907 84442
rect -16930 76723 -16690 76806
rect -16930 75068 -16849 76723
rect -18711 74828 -16849 75068
rect -16930 73398 -16849 74828
rect -16748 73398 -16690 76723
rect -13914 76729 -13674 76891
rect -13914 75253 -13848 76729
rect -14713 75013 -13848 75253
rect -16930 72559 -16690 73398
rect -13914 73404 -13848 75013
rect -13747 73404 -13674 76729
rect 11083 76732 11323 76878
rect 11083 75172 11143 76732
rect 11082 74932 11143 75172
rect -13914 73242 -13674 73404
rect 11083 73392 11143 74932
rect 11271 75172 11323 76732
rect 14083 76745 14323 76876
rect 11271 74932 12758 75172
rect 11271 73392 11323 74932
rect 11083 73244 11323 73392
rect 14083 73405 14144 76745
rect 14272 75164 14323 76745
rect 14272 74924 16757 75164
rect 14272 73405 14323 74924
rect 14083 73232 14323 73405
rect -16930 72495 -14071 72559
rect -16665 71802 -16599 71803
rect -16665 71738 -16664 71802
rect -16600 71738 -16599 71802
rect -15486 71799 -15422 72495
rect -15270 71805 -15204 71806
rect -16665 71737 -16599 71738
rect -15487 71798 -15421 71799
rect -16664 70898 -16600 71737
rect -15487 71734 -15486 71798
rect -15422 71734 -15421 71798
rect -15270 71741 -15269 71805
rect -15205 71741 -15204 71805
rect -14135 71803 -14071 72495
rect -15270 71740 -15204 71741
rect -14136 71802 -14070 71803
rect -15487 71733 -15421 71734
rect -15269 70994 -15205 71740
rect -14136 71738 -14135 71802
rect -14071 71738 -14070 71802
rect -14136 71737 -14070 71738
rect -15269 70898 -15242 70994
rect -16664 70834 -15242 70898
rect -16664 70303 -16600 70834
rect -16664 70298 -16489 70303
rect -18711 70143 -18665 70237
rect -16664 70234 -16554 70298
rect -16490 70234 -16489 70298
rect -15227 70286 -15163 70754
rect -15228 70285 -15162 70286
rect -16555 70233 -16489 70234
rect -15441 70284 -15375 70285
rect -15441 70220 -15440 70284
rect -15376 70220 -15375 70284
rect -15228 70221 -15227 70285
rect -15163 70221 -15162 70285
rect -15228 70220 -15162 70221
rect -14064 70285 -13998 70286
rect -14064 70221 -14063 70285
rect -13999 70221 -13998 70285
rect -14064 70220 -13998 70221
rect -15441 70219 -15375 70220
rect -15440 70143 -15376 70219
rect -14063 70143 -13999 70220
rect -18711 70079 -13999 70143
rect -18711 69997 -18665 70079
rect 36630 69334 36696 69335
rect 36630 69270 36631 69334
rect 36695 69270 36696 69334
rect 36630 69258 36696 69270
rect -16577 68743 -15239 68807
rect -16577 67614 -16513 68743
rect -15962 68262 -15898 68743
rect -14709 68743 -14240 68807
rect -15422 68516 -15358 68542
rect -15423 68515 -15357 68516
rect -15964 68261 -15889 68262
rect -15964 68105 -15963 68261
rect -15890 68105 -15889 68261
rect -15423 68166 -15422 68515
rect -15358 68166 -15357 68515
rect -14874 68265 -14810 68675
rect -15423 68165 -15357 68166
rect -14880 68264 -14805 68265
rect -15964 68104 -15889 68105
rect -16578 67613 -16512 67614
rect -16578 67549 -16577 67613
rect -16513 67549 -16512 67613
rect -15422 67608 -15358 68165
rect -14880 68108 -14879 68264
rect -14806 68108 -14805 68264
rect -14880 68107 -14805 68108
rect -14304 67619 -14240 68743
rect 36064 68742 36132 68743
rect 36064 68676 36065 68742
rect 36131 68676 36132 68742
rect 36064 68675 36132 68676
rect 36065 68638 36131 68675
rect 35475 68082 35543 68083
rect 35475 68016 35476 68082
rect 35542 68016 35543 68082
rect 35475 68015 35543 68016
rect -14305 67618 -14239 67619
rect -16578 67548 -16512 67549
rect -15423 67607 -15357 67608
rect -15423 67543 -15422 67607
rect -15358 67543 -15357 67607
rect -14305 67554 -14304 67618
rect -14240 67554 -14239 67618
rect -14305 67553 -14239 67554
rect -15423 67542 -15357 67543
rect -15422 67030 -15358 67542
rect -18715 66966 -15358 67030
rect -13096 66770 -13032 66772
rect -13097 66769 -13031 66770
rect -13097 66705 -13096 66769
rect -13032 66705 -13031 66769
rect -13097 66704 -13031 66705
rect -8074 66769 -8008 66770
rect -8074 66705 -8073 66769
rect -8009 66705 -8008 66769
rect -8074 66704 -8008 66705
rect -13096 59581 -13032 66704
rect -12316 66446 -12250 66447
rect -12316 66382 -12315 66446
rect -12251 66382 -12250 66446
rect -12316 66381 -12250 66382
rect -12315 59581 -12251 66381
rect -11305 66014 -11241 66018
rect -11306 66013 -11240 66014
rect -11306 65949 -11305 66013
rect -11241 65949 -11240 66013
rect -11306 65948 -11240 65949
rect -11305 59581 -11241 65948
rect -10536 65761 -10472 65768
rect -10537 65760 -10471 65761
rect -10537 65696 -10536 65760
rect -10472 65696 -10471 65760
rect -10537 65695 -10471 65696
rect -11072 63557 -10736 63558
rect -11072 63205 -11071 63557
rect -10737 63205 -10736 63557
rect -11072 63204 -10736 63205
rect -10536 59581 -10472 65695
rect -8073 65330 -8009 66704
rect -7267 66446 -7201 66447
rect -7267 66382 -7266 66446
rect -7202 66382 -7201 66446
rect -7267 66381 -7201 66382
rect -8074 65329 -8008 65330
rect -8074 65265 -8073 65329
rect -8009 65265 -8008 65329
rect -8074 65264 -8008 65265
rect -7266 65077 -7202 66381
rect -2674 66013 -2608 66014
rect -2674 65949 -2673 66013
rect -2609 65949 -2608 66013
rect -2674 65948 -2608 65949
rect -2673 65330 -2609 65948
rect -1867 65760 -1801 65761
rect -1867 65696 -1866 65760
rect -1802 65696 -1801 65760
rect -1867 65695 -1801 65696
rect -2674 65329 -2608 65330
rect -2674 65265 -2673 65329
rect -2609 65265 -2599 65329
rect -2674 65264 -2608 65265
rect -1866 65077 -1802 65695
rect -7267 65076 -7201 65077
rect -7267 65012 -7266 65076
rect -7202 65012 -7201 65076
rect -7267 65011 -7201 65012
rect -1867 65076 -1801 65077
rect -1867 65012 -1866 65076
rect -1802 65012 -1791 65076
rect -1867 65011 -1801 65012
rect 16717 64743 33332 64767
rect 16717 64169 17430 64743
rect 17496 64719 23958 64743
rect 17496 64191 20763 64719
rect 21288 64191 23958 64719
rect 17496 64169 23958 64191
rect 24024 64725 31574 64743
rect 24024 64197 28757 64725
rect 29282 64197 31574 64725
rect 24024 64169 31574 64197
rect 31640 64169 33332 64743
rect 16717 64147 33332 64169
rect -8074 63404 -7630 63405
rect -10188 63402 -10122 63403
rect -9885 63402 -9441 63403
rect -8074 63402 -8073 63404
rect -10188 63338 -10187 63402
rect -10123 63338 -9884 63402
rect -9442 63340 -8073 63402
rect -7631 63402 -7630 63404
rect -7631 63400 -3241 63402
rect -7631 63340 -6278 63400
rect -9442 63338 -6278 63340
rect -10188 63337 -10122 63338
rect -9885 63337 -9441 63338
rect -6279 63336 -6278 63338
rect -5836 63398 -3241 63400
rect -5836 63338 -4479 63398
rect -5836 63336 -5835 63338
rect -6279 63335 -5835 63336
rect -4480 63334 -4479 63338
rect -4037 63338 -3241 63398
rect -4037 63334 -4036 63338
rect -4480 63333 -4036 63334
rect -6940 63206 -6698 63207
rect -6940 62966 -6939 63206
rect -6699 62966 -6698 63206
rect -2711 63402 -2245 63403
rect -2711 63338 -2688 63402
rect -2246 63398 243 63402
rect -2246 63338 -886 63398
rect -2711 63337 -2245 63338
rect -887 63334 -886 63338
rect -444 63338 243 63398
rect -444 63334 -443 63338
rect -887 63333 -443 63334
rect 756 63232 1288 63233
rect 756 62992 757 63232
rect 1287 62992 1288 63232
rect 756 62991 1288 62992
rect -6940 62965 -6698 62966
rect 16715 62740 33227 62767
rect 16715 62728 17975 62740
rect 16715 62200 16766 62728
rect 17291 62200 17975 62728
rect 16715 62166 17975 62200
rect 18041 62166 19063 62740
rect 19129 62166 21239 62740
rect 21305 62166 22327 62740
rect 22393 62166 23415 62740
rect 23481 62166 24503 62740
rect 24569 62721 25591 62740
rect 24569 62193 24762 62721
rect 25287 62193 25591 62721
rect 24569 62166 25591 62193
rect 25657 62166 26679 62740
rect 26745 62166 28855 62740
rect 28921 62166 29943 62740
rect 30009 62166 31031 62740
rect 31097 62717 33227 62740
rect 31097 62189 32765 62717
rect 31097 62166 33227 62189
rect 16715 62147 33227 62166
rect -13469 59517 -13032 59581
rect -26125 49178 -23234 49223
rect -26125 49114 -25984 49178
rect -25640 49114 -23234 49178
rect -26125 48983 -23234 49114
rect -27162 43313 -26922 43373
rect -27162 43156 -27087 43313
rect -26990 43156 -26922 43313
rect -13469 43062 -13405 59517
rect -13096 52391 -13032 59517
rect -12693 59517 -12251 59581
rect -13097 52390 -13031 52391
rect -13097 52326 -13096 52390
rect -13032 52326 -13031 52390
rect -13097 52325 -13031 52326
rect -13470 43061 -13404 43062
rect -13470 42997 -13469 43061
rect -13405 42997 -13404 43061
rect -13470 42996 -13404 42997
rect -13469 42992 -13405 42996
rect -27162 42779 -27087 42916
rect -26990 42779 -26922 42916
rect -27162 42169 -26922 42779
rect -12693 42399 -12629 59517
rect -12315 52714 -12251 59517
rect -11713 59517 -11241 59581
rect -12316 52713 -12250 52714
rect -12316 52649 -12315 52713
rect -12251 52649 -12250 52713
rect -12316 52648 -12250 52649
rect -11713 44606 -11649 59517
rect -11305 53147 -11241 59517
rect -10905 59517 -10472 59581
rect -11306 53146 -11240 53147
rect -11306 53082 -11305 53146
rect -11241 53082 -11240 53146
rect -11306 53081 -11240 53082
rect -11362 47256 -11296 47257
rect -11362 47192 -11361 47256
rect -11297 47192 -11296 47256
rect -11362 47191 -11296 47192
rect -11361 44606 -11297 47191
rect -11713 44542 -11297 44606
rect -10905 44619 -10841 59517
rect -10536 53403 -10472 59517
rect 344 60827 640 60887
rect -6865 54597 -6801 54706
rect -6867 54596 -6801 54597
rect -8558 54595 -8492 54596
rect -6867 54595 -6866 54596
rect -8558 54531 -8557 54595
rect -8493 54532 -6866 54595
rect -6802 54595 -6801 54596
rect -5162 54595 -5096 54596
rect -3366 54595 -3300 54596
rect -1537 54595 -1471 54596
rect -6802 54532 -5161 54595
rect -8493 54531 -5161 54532
rect -5097 54531 -3365 54595
rect -3301 54531 -1536 54595
rect -1472 54531 240 54595
rect -8558 54530 -8492 54531
rect -5162 54530 -5096 54531
rect -3366 54530 -3300 54531
rect -1537 54530 -1471 54531
rect -6110 54404 -5866 54405
rect -9705 54403 -9461 54404
rect -6110 54403 -6109 54404
rect -9731 54339 -9704 54403
rect -9462 54402 -6109 54403
rect -9462 54339 -7909 54402
rect -9705 54338 -9461 54339
rect -7910 54338 -7909 54339
rect -7667 54340 -6109 54402
rect -5867 54403 -5866 54404
rect -4312 54403 -4068 54404
rect -5867 54340 -4311 54403
rect -7667 54339 -4311 54340
rect -4069 54339 -3237 54403
rect -7667 54338 -7666 54339
rect -4312 54338 -4068 54339
rect -7910 54337 -7666 54338
rect 176 54405 240 54531
rect -2514 54404 -2270 54405
rect 175 54404 241 54405
rect -2514 54403 -2513 54404
rect -2707 54340 -2513 54403
rect -2271 54403 -2270 54404
rect -711 54403 -467 54404
rect -2271 54340 -710 54403
rect -2707 54339 -710 54340
rect -468 54339 -467 54403
rect 175 54340 176 54404
rect 240 54340 241 54404
rect 175 54339 241 54340
rect -711 54338 -467 54339
rect -7266 54083 -7200 54084
rect -7266 54019 -7265 54083
rect -7201 54019 -7200 54083
rect -7266 54018 -7200 54019
rect -1866 54083 -1800 54084
rect -1866 54019 -1865 54083
rect -1801 54019 -1791 54083
rect -1866 54018 -1800 54019
rect -8074 53830 -8008 53831
rect -8074 53766 -8073 53830
rect -8009 53766 -8008 53830
rect -8074 53765 -8008 53766
rect -10537 53402 -10471 53403
rect -10537 53338 -10536 53402
rect -10472 53338 -10471 53402
rect -10537 53337 -10471 53338
rect -8073 52391 -8009 53765
rect -7265 52714 -7201 54018
rect -2674 53830 -2608 53831
rect -2674 53766 -2673 53830
rect -2609 53766 -2599 53830
rect -2674 53765 -2608 53766
rect -2673 53147 -2609 53765
rect -1865 53403 -1801 54018
rect -1866 53402 -1800 53403
rect -1866 53338 -1865 53402
rect -1801 53338 -1800 53402
rect 344 53400 347 60827
rect -1866 53337 -1800 53338
rect -2674 53146 -2608 53147
rect -2674 53082 -2673 53146
rect -2609 53082 -2608 53146
rect 338 53121 347 53400
rect 519 60125 640 60827
rect 10176 60836 10552 60837
rect 519 60124 768 60125
rect 519 59884 756 60124
rect 10176 60113 10177 60836
rect 519 57511 640 59884
rect 9291 59873 10177 60113
rect 5390 58930 5630 59104
rect 5390 58752 5410 58930
rect 5588 58752 5630 58930
rect 5390 57511 5630 58752
rect 519 57475 5630 57511
rect 519 57297 2047 57475
rect 2225 57297 4047 57475
rect 4225 57297 5630 57475
rect 519 57271 5630 57297
rect 519 56750 640 57271
rect 519 56749 668 56750
rect 519 56509 756 56749
rect 519 56508 668 56509
rect 519 53400 640 56508
rect 5390 55930 5630 57271
rect 10176 56738 10177 59873
rect 9290 56498 10177 56738
rect 5390 55752 5410 55930
rect 5588 55752 5630 55930
rect 5390 55603 5630 55752
rect 519 53399 671 53400
rect 519 53374 1315 53399
rect 519 53134 756 53374
rect 1286 53345 1315 53374
rect 10176 53363 10177 56498
rect 1286 53179 4187 53345
rect 1286 53167 4007 53179
rect 1286 53134 1315 53167
rect 519 53121 1315 53134
rect 338 53104 1315 53121
rect -2674 53081 -2608 53082
rect 4006 53001 4007 53167
rect 4185 53001 4187 53179
rect 9290 53123 10177 53363
rect 4006 53000 4187 53001
rect -7266 52713 -7200 52714
rect -7266 52649 -7265 52713
rect -7201 52649 -7200 52713
rect -7266 52648 -7200 52649
rect -8074 52390 -8008 52391
rect -8074 52326 -8073 52390
rect -8009 52326 -8008 52390
rect -8074 52325 -8008 52326
rect 4009 52033 4187 53000
rect 7724 52036 7904 52037
rect 7724 52033 7725 52036
rect 4009 51858 7725 52033
rect 7903 52033 7904 52036
rect 10176 52033 10177 53123
rect 7903 51858 10177 52033
rect 4009 51855 10177 51858
rect -9010 51461 -7237 51701
rect -9010 51250 -8770 51461
rect -9010 51249 -8769 51250
rect -9010 51014 -8854 51249
rect -8770 51014 -8769 51249
rect -7723 51247 -7657 51248
rect -7723 51183 -7722 51247
rect -7658 51183 -7657 51247
rect -7723 51182 -7657 51183
rect -8855 51013 -8769 51014
rect -8875 50791 -8777 50792
rect -8875 50378 -8874 50791
rect -8780 50378 -8777 50791
rect -8875 50377 -8777 50378
rect -8481 50441 -8415 50442
rect -8481 50377 -8480 50441
rect -8416 50377 -8415 50441
rect -8481 50376 -8415 50377
rect -8480 50073 -8416 50376
rect -8481 50072 -8415 50073
rect -8481 50008 -8480 50072
rect -8416 50008 -8415 50072
rect -8481 50007 -8415 50008
rect -10488 46633 -10422 46634
rect -10488 46569 -10487 46633
rect -10423 46569 -10422 46633
rect -10488 46568 -10422 46569
rect -10487 44619 -10423 46568
rect -10905 44555 -10423 44619
rect -12694 42398 -12628 42399
rect -12694 42334 -12693 42398
rect -12629 42334 -12628 42398
rect -12694 42333 -12628 42334
rect -12693 42328 -12629 42333
rect -27162 41002 -27082 42169
rect -26995 41002 -26922 42169
rect -21476 42163 -21410 42164
rect -21476 42099 -21475 42163
rect -21411 42099 -17680 42163
rect -21476 42098 -21410 42099
rect -27162 40643 -26922 41002
rect -27162 39950 -27077 40643
rect -26990 39950 -26922 40643
rect -17744 39824 -17680 42099
rect -17744 39760 -17097 39824
rect -27162 39476 -27077 39710
rect -26990 39476 -26922 39710
rect -31813 39166 -31747 39167
rect -31813 38827 -31812 39166
rect -31748 39023 -31747 39166
rect -27162 39120 -26922 39476
rect -31748 38959 -30945 39023
rect -31748 38827 -31747 38959
rect -31813 38826 -31747 38827
rect -31812 38613 -31746 38614
rect -31812 38415 -31811 38613
rect -34755 38351 -31811 38415
rect -31812 38141 -31811 38351
rect -31747 38141 -31746 38613
rect -31009 38509 -30945 38959
rect -29615 38413 -29149 38414
rect -30743 38349 -29614 38413
rect -29150 38349 -29149 38413
rect -29615 38348 -29149 38349
rect -31812 38140 -31746 38141
rect -27162 38232 -27082 39120
rect -26998 38232 -26922 39120
rect -27162 37353 -26922 38232
rect -18956 39537 -18716 39689
rect -18956 37904 -18883 39537
rect -22729 37664 -18883 37904
rect -29653 37323 -29142 37324
rect -30755 37259 -29652 37323
rect -29143 37259 -29142 37323
rect -29653 37258 -29142 37259
rect -27162 36465 -27079 37353
rect -26995 36465 -26922 37353
rect -27162 36160 -26922 36465
rect -27162 35881 -27077 36160
rect -26996 35881 -26922 36160
rect -18956 36124 -18883 37664
rect -18807 36124 -18716 39537
rect -11713 38791 -11649 44542
rect -11714 38790 -11648 38791
rect -13395 38783 -13331 38784
rect -14898 38719 -13331 38783
rect -11714 38726 -11713 38790
rect -11649 38726 -11648 38790
rect -11714 38725 -11648 38726
rect -11713 38724 -11649 38725
rect -18956 35957 -18716 36124
rect -17743 36329 -17006 36393
rect -27162 34985 -27077 35641
rect -26996 34985 -26922 35641
rect -27162 34691 -26922 34985
rect -27162 33498 -27079 34691
rect -27000 33498 -26922 34691
rect -27162 32899 -26922 33498
rect -21519 33551 -21453 33552
rect -17743 33551 -17679 36329
rect -21519 33487 -21518 33551
rect -21454 33487 -17679 33551
rect -21519 33486 -21453 33487
rect -15139 33180 -15075 35346
rect -13395 34677 -13331 38719
rect -10905 38448 -10841 44555
rect -9209 43061 -9143 43062
rect -9209 42997 -9208 43061
rect -9144 42997 -9143 43061
rect -9209 42996 -9143 42997
rect -10070 42398 -10004 42399
rect -10070 42334 -10069 42398
rect -10005 42334 -10004 42398
rect -10070 42333 -10004 42334
rect -10906 38447 -10840 38448
rect -10906 38383 -10905 38447
rect -10841 38383 -10840 38447
rect -10906 38382 -10840 38383
rect -10905 38376 -10841 38382
rect -10069 35352 -10005 42333
rect -9208 35942 -9144 42996
rect -8480 37372 -8416 50007
rect -7722 49425 -7658 51182
rect -5972 51121 -5695 51124
rect -5972 51101 139 51121
rect -5972 51074 -3231 51101
rect -2701 51074 139 51101
rect -5972 51066 -3362 51074
rect -5972 50883 -5688 51066
rect -3888 50896 -3362 51066
rect -2536 51064 139 51074
rect -2536 50896 -1655 51064
rect -3888 50883 -3231 50896
rect -5972 50861 -3231 50883
rect -2701 50886 -1655 50896
rect -765 50886 139 51064
rect -2701 50861 139 50886
rect -5972 50845 139 50861
rect -5972 50720 -5695 50845
rect -7723 49424 -7657 49425
rect -7723 49360 -7722 49424
rect -7658 49360 -7657 49424
rect -7723 49359 -7657 49360
rect -7722 37900 -7658 49359
rect -5972 47776 -5932 50720
rect -5748 48791 -5695 50720
rect -138 50774 139 50845
rect -138 48791 -78 50774
rect -5748 48773 -78 48791
rect -5748 48533 -3237 48773
rect -2707 48533 -78 48773
rect -5748 48514 -78 48533
rect -5748 47776 -5695 48514
rect -5972 47688 -5695 47776
rect -138 47752 -78 48514
rect 121 47752 139 50774
rect 600 49999 1298 50017
rect 600 49759 756 49999
rect 1286 49759 1298 49999
rect 10176 49988 10177 51855
rect 600 49722 1298 49759
rect 9290 49748 10177 49988
rect -138 47715 139 47752
rect 10176 47617 10177 49748
rect 10551 47617 10552 60836
rect 16717 60743 33332 60767
rect 16717 60169 17430 60743
rect 17496 60169 18518 60743
rect 18584 60169 19606 60743
rect 19672 60169 20694 60743
rect 20760 60719 21782 60743
rect 20760 60191 20763 60719
rect 21288 60191 21782 60719
rect 20760 60169 21782 60191
rect 21848 60169 22870 60743
rect 22936 60169 23958 60743
rect 24024 60169 25046 60743
rect 25112 60169 26134 60743
rect 26200 60169 27222 60743
rect 27288 60169 28310 60743
rect 28376 60725 29398 60743
rect 28376 60197 28757 60725
rect 29282 60197 29398 60725
rect 28376 60169 29398 60197
rect 29464 60169 30486 60743
rect 30552 60169 31574 60743
rect 31640 60169 33332 60743
rect 16717 60147 33332 60169
rect 16715 58740 33227 58767
rect 16715 58728 17975 58740
rect 16715 58200 16766 58728
rect 17291 58200 17975 58728
rect 16715 58166 17975 58200
rect 18041 58166 19063 58740
rect 19129 58166 20151 58740
rect 20217 58166 21239 58740
rect 21305 58166 22327 58740
rect 22393 58166 23415 58740
rect 23481 58166 24503 58740
rect 24569 58721 25591 58740
rect 24569 58193 24762 58721
rect 25287 58193 25591 58721
rect 24569 58166 25591 58193
rect 25657 58166 26679 58740
rect 26745 58166 27767 58740
rect 27833 58166 28855 58740
rect 28921 58166 29943 58740
rect 30009 58166 31031 58740
rect 31097 58717 33227 58740
rect 31097 58189 32765 58717
rect 31097 58166 33227 58189
rect 16715 58147 33227 58166
rect 16717 56743 33332 56767
rect 16717 56169 17430 56743
rect 17496 56169 18518 56743
rect 18584 56169 19606 56743
rect 19672 56169 20694 56743
rect 20760 56719 21782 56743
rect 20760 56191 20763 56719
rect 21288 56191 21782 56719
rect 20760 56169 21782 56191
rect 21848 56169 22870 56743
rect 22936 56169 23958 56743
rect 24024 56169 25046 56743
rect 25112 56169 26134 56743
rect 26200 56169 27222 56743
rect 27288 56169 28310 56743
rect 28376 56725 29398 56743
rect 28376 56197 28757 56725
rect 29282 56197 29398 56725
rect 28376 56169 29398 56197
rect 29464 56169 30486 56743
rect 30552 56169 31574 56743
rect 31640 56169 33332 56743
rect 16717 56147 33332 56169
rect 16715 54740 33227 54767
rect 16715 54728 17975 54740
rect 16715 54200 16766 54728
rect 17291 54200 17975 54728
rect 16715 54166 17975 54200
rect 18041 54166 19063 54740
rect 19129 54166 20151 54740
rect 20217 54166 21239 54740
rect 21305 54166 22327 54740
rect 22393 54166 23415 54740
rect 23481 54166 24503 54740
rect 24569 54721 25591 54740
rect 24569 54193 24762 54721
rect 25287 54193 25591 54721
rect 24569 54166 25591 54193
rect 25657 54166 26679 54740
rect 26745 54166 27767 54740
rect 27833 54166 28855 54740
rect 28921 54166 29943 54740
rect 30009 54166 31031 54740
rect 31097 54717 33227 54740
rect 31097 54189 32765 54717
rect 31097 54166 33227 54189
rect 16715 54147 33227 54166
rect 16717 52743 33332 52767
rect 16717 52169 17430 52743
rect 17496 52169 18518 52743
rect 18584 52169 19606 52743
rect 19672 52169 20694 52743
rect 20760 52719 21782 52743
rect 20760 52191 20763 52719
rect 21288 52191 21782 52719
rect 20760 52169 21782 52191
rect 21848 52169 22870 52743
rect 22936 52169 23958 52743
rect 24024 52169 25046 52743
rect 25112 52169 26134 52743
rect 26200 52169 27222 52743
rect 27288 52169 28310 52743
rect 28376 52725 29398 52743
rect 28376 52197 28757 52725
rect 29282 52197 29398 52725
rect 28376 52169 29398 52197
rect 29464 52169 30486 52743
rect 30552 52169 31574 52743
rect 31640 52169 33332 52743
rect 16717 52147 33332 52169
rect 16715 50740 33227 50767
rect 16715 50728 17975 50740
rect 16715 50200 16766 50728
rect 17291 50200 17975 50728
rect 16715 50166 17975 50200
rect 18041 50166 20151 50740
rect 20217 50166 21239 50740
rect 21305 50166 23415 50740
rect 23481 50166 24503 50740
rect 24569 50721 25591 50740
rect 24569 50193 24762 50721
rect 25287 50193 25591 50721
rect 24569 50166 25591 50193
rect 25657 50166 27767 50740
rect 27833 50166 28855 50740
rect 28921 50166 31031 50740
rect 31097 50717 33227 50740
rect 31097 50189 32765 50717
rect 31097 50166 33227 50189
rect 16715 50147 33227 50166
rect 16717 48743 33332 48767
rect 16717 48169 17430 48743
rect 17496 48169 18518 48743
rect 18584 48169 19606 48743
rect 19672 48169 20694 48743
rect 20760 48719 21782 48743
rect 20760 48191 20763 48719
rect 21288 48191 21782 48719
rect 20760 48169 21782 48191
rect 21848 48169 22870 48743
rect 22936 48169 23958 48743
rect 24024 48725 29398 48743
rect 24024 48197 28757 48725
rect 29282 48197 29398 48725
rect 24024 48169 29398 48197
rect 29464 48169 30486 48743
rect 30552 48169 31574 48743
rect 31640 48169 33332 48743
rect 16717 48147 33332 48169
rect 10176 47616 10552 47617
rect -6412 47256 -6346 47257
rect -6412 47192 -6411 47256
rect -6347 47192 12030 47256
rect -6412 47191 -6346 47192
rect -6412 46633 -6346 46634
rect -6412 46569 -6411 46633
rect -6347 46569 11411 46633
rect -6412 46568 -6346 46569
rect -5972 46274 -5674 46319
rect -5972 39819 -5924 46274
rect -5722 45377 -5674 46274
rect 10179 46128 10552 46129
rect 330 45844 619 45964
rect -5722 45355 -1240 45377
rect -5722 45307 -3248 45355
rect -5722 45129 -4101 45307
rect -3923 45129 -3248 45307
rect -5722 45115 -3248 45129
rect -2718 45115 -1240 45355
rect -5722 45079 -1240 45115
rect -5722 39891 -5674 45079
rect -1538 44459 -1240 45079
rect -1538 44281 -1482 44459
rect -1304 44281 -1240 44459
rect -1538 44206 -1240 44281
rect 330 44318 344 45844
rect 558 44544 619 45844
rect 10179 44544 10180 46128
rect 558 44514 10180 44544
rect 558 44318 752 44514
rect 330 44274 752 44318
rect 1282 44508 10180 44514
rect 1282 44330 2132 44508
rect 2310 44330 4132 44508
rect 4310 44330 6132 44508
rect 6310 44330 8132 44508
rect 8310 44330 10180 44508
rect 1282 44274 10180 44330
rect 330 44255 10180 44274
rect 10179 43238 10180 44255
rect 9290 42998 10180 43238
rect 325 41383 565 41411
rect -5722 39886 -135 39891
rect -5722 39846 -3233 39886
rect -2703 39846 -135 39886
rect -5722 39819 -5684 39846
rect -5972 39748 -5684 39819
rect -5713 39666 -5684 39748
rect -148 39666 -135 39846
rect 325 39855 352 41383
rect 512 40868 565 41383
rect 512 40629 762 40868
rect 512 40628 928 40629
rect 512 39855 565 40628
rect 10179 39867 10180 42998
rect 10551 39867 10552 46128
rect 10179 39866 10552 39867
rect 325 39810 565 39855
rect -5713 39646 -3233 39666
rect -2703 39646 -135 39666
rect -5713 39636 -135 39646
rect 1286 39286 2638 39350
rect 2512 38881 2638 39286
rect -4714 38790 -4648 38791
rect -4714 38726 -4713 38790
rect -4649 38726 -4648 38790
rect -4714 38725 -4648 38726
rect -7723 37899 -7657 37900
rect -7723 37835 -7722 37899
rect -7658 37835 -7657 37899
rect -7723 37834 -7657 37835
rect -8481 37371 -8415 37372
rect -8481 37307 -8480 37371
rect -8416 37307 -8415 37371
rect -8481 37306 -8415 37307
rect -9209 35941 -9143 35942
rect -9209 35877 -9208 35941
rect -9144 35877 -9143 35941
rect -9209 35876 -9143 35877
rect -10070 35351 -10004 35352
rect -10070 35287 -10069 35351
rect -10005 35287 -10004 35351
rect -10070 35286 -10004 35287
rect -13396 34676 -13330 34677
rect -13396 34612 -13395 34676
rect -13331 34612 -13330 34676
rect -13396 34611 -13330 34612
rect -4713 34196 -4649 38725
rect 2512 38642 2513 38881
rect 2595 38642 2638 38881
rect 2512 38632 2638 38642
rect -4124 38447 -4058 38448
rect -4124 38383 -4123 38447
rect -4059 38383 -4058 38447
rect -4124 38382 -4058 38383
rect 2514 38420 2640 38422
rect -4714 34195 -4648 34196
rect -4714 34131 -4713 34195
rect -4649 34131 -4648 34195
rect -4714 34130 -4648 34131
rect -4123 33851 -4059 38382
rect 2514 37996 2515 38420
rect 2614 37996 2640 38420
rect 2514 37971 2640 37996
rect 2514 37907 4761 37971
rect -2398 37900 -2334 37901
rect -2399 37899 -2333 37900
rect -761 37899 -695 37900
rect 1472 37899 1538 37900
rect -2399 37835 -2398 37899
rect -2334 37835 -2333 37899
rect -777 37835 -760 37899
rect -696 37835 1473 37899
rect 1537 37835 1569 37899
rect 2514 37875 2614 37907
rect -2399 37834 -2333 37835
rect -761 37834 -695 37835
rect 1472 37834 1538 37835
rect -2815 37372 -2751 37375
rect -2816 37371 -2750 37372
rect -2816 37307 -2815 37371
rect -2751 37307 -2750 37371
rect -2816 37306 -2750 37307
rect -4124 33850 -4058 33851
rect -4124 33786 -4123 33850
rect -4059 33786 -4058 33850
rect -4124 33785 -4058 33786
rect -15140 33179 -15074 33180
rect -15140 33115 -15139 33179
rect -15075 33115 -15074 33179
rect -15140 33114 -15074 33115
rect -27162 32767 -27084 32899
rect -27005 32767 -26922 32899
rect -27162 32365 -27084 32527
rect -27005 32365 -26922 32527
rect -27162 32329 -26922 32365
rect -3919 29752 -3853 29753
rect -3919 29688 -3918 29752
rect -3854 29688 -3853 29752
rect -3919 29687 -3853 29688
rect -5279 29330 -5215 29332
rect -5280 29329 -5214 29330
rect -5280 29265 -5279 29329
rect -5215 29265 -5214 29329
rect -5280 29264 -5214 29265
rect -15741 28708 -15500 28709
rect -18708 28468 -15500 28708
rect -17700 27644 -17460 28468
rect -17700 27516 -17635 27644
rect -17507 27516 -17460 27644
rect -15741 28098 -15500 28468
rect -15741 27645 -15712 28098
rect -15613 27645 -15500 28098
rect -12394 28076 -12266 28089
rect -12394 27670 -12389 28076
rect -12316 28003 -12266 28076
rect -12316 27875 -11237 28003
rect -12316 27670 -12266 27875
rect -12394 27658 -12266 27670
rect -15741 27619 -15500 27645
rect -17700 27461 -17460 27516
rect -12386 27428 -12258 27461
rect -12395 27427 -12258 27428
rect -12395 27388 -12394 27427
rect -14704 27260 -12394 27388
rect -12395 27198 -12394 27260
rect -12297 27388 -12258 27427
rect -12297 27260 -12247 27388
rect -12297 27198 -12258 27260
rect -12395 27197 -12258 27198
rect -12386 27188 -12258 27197
rect -35224 26612 -34761 26668
rect -38191 26611 -34761 26612
rect -38191 26514 -38190 26611
rect -34856 26514 -34761 26611
rect -38191 26513 -34855 26514
rect -12422 26486 -12294 26493
rect -17691 26415 -17458 26461
rect -17691 26287 -17635 26415
rect -17507 26287 -17458 26415
rect -17691 25810 -17458 26287
rect -15742 26281 -15509 26354
rect -15742 26044 -15725 26281
rect -15636 26044 -15509 26281
rect -12422 26057 -12396 26486
rect -12301 26330 -12294 26486
rect -11717 26330 -11589 27875
rect -5279 27533 -5215 29264
rect -5280 27532 -5214 27533
rect -5280 27468 -5279 27532
rect -5215 27468 -5214 27532
rect -5280 27467 -5214 27468
rect -12301 26202 -11589 26330
rect -12301 26057 -12294 26202
rect -12422 26053 -12294 26057
rect -15742 25810 -15509 26044
rect -17691 25578 -15238 25810
rect -12383 25765 -12255 25856
rect -14708 25637 -12255 25765
rect -12383 25595 -12255 25637
rect -17691 25577 -14847 25578
rect -25450 25482 -25368 25483
rect -25450 25433 -25449 25482
rect -26698 25305 -25449 25433
rect -25450 25175 -25449 25305
rect -25369 25433 -25368 25482
rect -25369 25305 -25316 25433
rect -25369 25175 -25368 25305
rect -25450 25174 -25368 25175
rect -17691 25002 -17458 25577
rect -11717 25313 -11589 26202
rect -11324 25665 -11260 25666
rect -11325 25664 -11259 25665
rect -11325 25600 -11324 25664
rect -11260 25600 -11259 25664
rect -11325 25599 -11259 25600
rect -25453 24945 -25364 24946
rect -25453 24714 -25452 24945
rect -25365 24893 -25364 24945
rect -25365 24765 -23236 24893
rect -25365 24714 -25364 24765
rect -25453 24713 -25364 24714
rect -17691 24874 -17635 25002
rect -17507 24874 -17458 25002
rect -17691 24811 -17458 24874
rect -12398 25185 -11589 25313
rect -12398 24712 -12270 25185
rect -11978 24872 -11912 24873
rect -11978 24808 -11977 24872
rect -11913 24808 -11912 24872
rect -11978 24807 -11912 24808
rect -12398 24458 -12393 24712
rect -12328 24458 -12270 24712
rect -12398 24441 -12270 24458
rect -12434 24239 -12306 24264
rect -12434 24003 -12398 24239
rect -12316 24003 -12306 24239
rect -17692 23773 -17452 23854
rect -17692 23731 -17635 23773
rect -18811 23730 -17635 23731
rect -38742 23605 -34770 23710
rect -38742 23503 -38182 23605
rect -34852 23503 -34770 23605
rect -38742 23474 -34770 23503
rect -18709 23645 -17635 23730
rect -17507 23645 -17452 23773
rect -18709 23491 -17452 23645
rect -15726 23637 -15493 23639
rect -15726 23405 -15725 23637
rect -15658 23405 -15237 23637
rect -15726 23404 -15237 23405
rect -12434 23592 -12306 24003
rect -14707 23464 -12306 23592
rect -11977 23519 -11913 24807
rect -11324 23888 -11260 25599
rect -11325 23887 -11259 23888
rect -11325 23823 -11324 23887
rect -11260 23823 -11259 23887
rect -11325 23822 -11259 23823
rect -11978 23518 -11912 23519
rect -16600 22724 -16534 22725
rect -16600 22660 -16599 22724
rect -16535 22660 -16534 22724
rect -16600 22659 -16534 22660
rect -16599 20652 -16535 22659
rect -13885 22584 -13757 23464
rect -11978 23454 -11977 23518
rect -11913 23454 -11912 23518
rect -11978 23453 -11912 23454
rect -11977 23442 -11913 23453
rect -12390 23277 -12318 23278
rect -12390 22857 -12389 23277
rect -12319 23108 -12258 23277
rect -12319 22980 -11246 23108
rect -12319 22857 -12258 22980
rect -12390 22856 -12258 22857
rect -12386 22837 -12258 22856
rect -12400 22624 -12272 22651
rect -12400 22584 -12391 22624
rect -13885 22456 -12391 22584
rect -12400 22399 -12391 22456
rect -12323 22399 -12272 22624
rect -12400 22350 -12272 22399
rect -16600 20651 -16534 20652
rect -16600 20587 -16599 20651
rect -16535 20587 -16534 20651
rect -16600 20586 -16534 20587
rect -38169 19065 -35218 19066
rect -38169 18987 -38168 19065
rect -5279 19044 -5215 27467
rect -3918 26856 -3854 29687
rect -3919 26855 -3853 26856
rect -3919 26791 -3918 26855
rect -3854 26791 -3853 26855
rect -3919 26790 -3853 26791
rect -3918 19044 -3854 26790
rect -2815 19514 -2751 37306
rect -2816 19513 -2750 19514
rect -2816 19449 -2815 19513
rect -2751 19449 -2750 19513
rect -2816 19448 -2750 19449
rect -2398 19213 -2334 37834
rect -761 37370 -695 37371
rect 1995 37370 2061 37371
rect -761 37306 -760 37370
rect -696 37306 1996 37370
rect 2060 37306 2094 37370
rect -761 37305 -695 37306
rect 1995 37305 2061 37306
rect 2167 37149 2233 37150
rect 2167 36996 2168 37149
rect 1287 36932 2168 36996
rect 2167 36898 2168 36932
rect 2232 36898 2233 37149
rect 2167 36897 2233 36898
rect 2169 36669 2233 36680
rect 2168 36668 2234 36669
rect 2168 36250 2169 36668
rect 2233 36567 2234 36668
rect 2233 36503 4768 36567
rect 2233 36250 2234 36503
rect 2168 36249 2234 36250
rect 3664 36095 3783 36115
rect 5179 36105 5243 36420
rect 5054 36104 5352 36105
rect 3581 36094 3812 36095
rect 3581 36030 3582 36094
rect 3811 36030 3812 36094
rect 3581 36029 3812 36030
rect 3664 35957 3783 36029
rect 5054 36018 5055 36104
rect 5351 36018 5352 36104
rect 5629 36098 5748 36115
rect 5573 36097 5802 36098
rect 5573 36027 5574 36097
rect 5801 36027 5802 36097
rect 6981 36090 7100 36125
rect 9645 36092 9764 36100
rect 9574 36091 9803 36092
rect 5573 36026 5802 36027
rect 6935 36089 7158 36090
rect 5054 36017 5352 36018
rect 5629 35957 5748 36026
rect 6935 36020 6936 36089
rect 7157 36020 7158 36089
rect 6935 36019 7158 36020
rect 6981 35957 7100 36019
rect 1304 35838 8758 35957
rect 9574 36023 9575 36091
rect 9802 36023 9803 36091
rect 9574 36022 9803 36023
rect 9645 35957 9764 36022
rect 9288 35838 9764 35957
rect 3120 35672 3241 35673
rect 3120 35553 3121 35672
rect 3240 35553 3241 35672
rect 9069 35650 9190 35651
rect 3120 35552 3241 35553
rect 7502 35641 7623 35642
rect 3121 35418 3240 35552
rect 7502 35522 7503 35641
rect 7622 35522 7623 35641
rect 9069 35531 9070 35650
rect 9189 35531 9190 35650
rect 9069 35530 9190 35531
rect 7502 35521 7623 35522
rect 3046 35299 4774 35418
rect 7503 35418 7622 35521
rect 9070 35418 9189 35530
rect 5304 35299 9189 35418
rect 4701 31450 4765 32172
rect 7965 31812 8029 32172
rect 7964 31811 8030 31812
rect 7964 31747 7965 31811
rect 8029 31747 8030 31811
rect 7964 31746 8030 31747
rect 3944 31386 4765 31450
rect 4941 31390 5739 31454
rect 6991 31390 7789 31454
rect 7965 31450 8029 31746
rect 4701 31372 4765 31386
rect 7965 31386 8786 31450
rect 11347 31392 11411 46569
rect 11346 31391 11412 31392
rect 7965 31372 8029 31386
rect 11346 31327 11347 31391
rect 11411 31327 11412 31391
rect 11346 31326 11412 31327
rect 3698 30389 3762 31187
rect 4353 30432 4419 30433
rect 4353 30368 4354 30432
rect 4418 30368 4705 30432
rect 5965 30394 6029 31192
rect 6701 30394 6765 31192
rect 8327 30437 8393 30438
rect 8028 30373 8328 30437
rect 8392 30373 8393 30437
rect 8968 30389 9032 31187
rect 8327 30372 8393 30373
rect 4353 30367 4419 30368
rect 3325 30305 3391 30306
rect 3325 30241 3326 30305
rect 3390 30241 3743 30305
rect 3325 30240 3391 30241
rect 3698 29389 3762 30187
rect 4701 29396 4765 30194
rect 5965 29394 6029 30192
rect 6701 29394 6765 30192
rect 7965 29396 8029 30194
rect 8968 29389 9032 30187
rect 3698 28389 3762 29167
rect 4967 28378 5031 29176
rect 5965 28394 6029 29192
rect 6701 28394 6765 29192
rect 7699 28378 7763 29176
rect 8968 28389 9032 29187
rect 10632 28804 10698 28805
rect 10632 28740 10633 28804
rect 10697 28740 10698 28804
rect 10632 28739 10698 28740
rect 3698 27389 3762 28187
rect 5965 27394 6029 28192
rect 6701 27394 6765 28192
rect 8968 27389 9032 28187
rect 4703 27188 4767 27200
rect 7963 27188 8027 27200
rect 3966 27124 4767 27188
rect 4966 27124 5764 27188
rect 6966 27124 7764 27188
rect 7963 27124 8764 27188
rect 4703 26402 4767 27124
rect 7963 26402 8027 27124
rect 7600 24848 7666 24849
rect 7600 24784 7601 24848
rect 7665 24784 7666 24848
rect 7600 24783 7666 24784
rect 5718 24595 5782 24717
rect 5714 24594 5784 24595
rect 5714 24186 5715 24594
rect 5783 24186 5784 24594
rect 7265 24593 7331 24594
rect 7265 24529 7266 24593
rect 7330 24529 7331 24593
rect 7265 24528 7331 24529
rect 5714 24185 5784 24186
rect 4779 23159 5244 23160
rect 4779 22919 4780 23159
rect 5243 22919 5244 23159
rect 5718 23064 5782 24185
rect 7266 23888 7330 24528
rect 7265 23887 7331 23888
rect 7265 23823 7266 23887
rect 7330 23823 7331 23887
rect 7265 23822 7331 23823
rect 5717 23063 5783 23064
rect 5717 22999 5718 23063
rect 5782 22999 5783 23063
rect 5717 22998 5783 22999
rect 4779 22918 5244 22919
rect 7601 22274 7665 24783
rect 8128 24530 8194 24531
rect 8128 24466 8129 24530
rect 8193 24466 8194 24530
rect 8128 24465 8194 24466
rect 8129 22725 8193 24465
rect 8786 23246 8787 23255
rect 8943 23246 8944 23255
rect 8786 23245 8944 23246
rect 8128 22724 8194 22725
rect 8128 22660 8129 22724
rect 8193 22660 8194 22724
rect 8128 22659 8194 22660
rect 8129 22651 8193 22659
rect 7600 22273 7666 22274
rect 7600 22209 7601 22273
rect 7665 22209 7666 22273
rect 7600 22208 7666 22209
rect 10633 20950 10697 28739
rect 11347 26351 11411 31326
rect 11966 30773 12030 47192
rect 16715 46740 33227 46767
rect 16715 46728 17975 46740
rect 16715 46200 16766 46728
rect 17291 46200 17975 46728
rect 16715 46166 17975 46200
rect 18041 46166 19063 46740
rect 19129 46166 20151 46740
rect 20217 46166 21239 46740
rect 21305 46166 22327 46740
rect 22393 46166 24503 46740
rect 24569 46721 25591 46740
rect 24569 46193 24762 46721
rect 25287 46193 25591 46721
rect 24569 46166 25591 46193
rect 25657 46166 26679 46740
rect 26745 46166 27767 46740
rect 27833 46166 28855 46740
rect 28921 46166 29943 46740
rect 30009 46166 31031 46740
rect 31097 46717 33227 46740
rect 31097 46189 32765 46717
rect 31097 46166 33227 46189
rect 16715 46147 33227 46166
rect 18244 45748 18310 45749
rect 18244 45684 18245 45748
rect 18309 45684 18310 45748
rect 18244 45683 18310 45684
rect 18790 45748 18856 45749
rect 18790 45684 18791 45748
rect 18855 45684 18856 45748
rect 21516 45748 21582 45749
rect 18790 45683 18856 45684
rect 19336 45739 19402 45740
rect 18245 44702 18309 45683
rect 18791 45073 18855 45683
rect 19336 45675 19337 45739
rect 19401 45675 19402 45739
rect 19336 45674 19402 45675
rect 19881 45738 19947 45739
rect 19881 45674 19882 45738
rect 19946 45674 19947 45738
rect 21516 45684 21517 45748
rect 21581 45684 21582 45748
rect 26405 45742 26471 45743
rect 22597 45741 22663 45742
rect 21516 45683 21582 45684
rect 22050 45735 22116 45736
rect 18790 45072 18856 45073
rect 18790 45008 18791 45072
rect 18855 45008 18856 45072
rect 18790 45007 18856 45008
rect 18244 44701 18310 44702
rect 18244 44637 18245 44701
rect 18309 44637 18310 44701
rect 18244 44636 18310 44637
rect 18245 38437 18309 44636
rect 13830 38436 13896 38437
rect 13830 38372 13831 38436
rect 13895 38372 13896 38436
rect 13830 38371 13896 38372
rect 18244 38436 18310 38437
rect 18244 38372 18245 38436
rect 18309 38372 18310 38436
rect 18244 38371 18310 38372
rect 13831 31392 13895 38371
rect 18791 37862 18855 45007
rect 19337 41012 19401 45674
rect 19881 45673 19947 45674
rect 19882 41383 19946 45673
rect 19881 41382 19947 41383
rect 19881 41318 19882 41382
rect 19946 41318 19947 41382
rect 19881 41317 19947 41318
rect 19336 41011 19402 41012
rect 19336 40947 19337 41011
rect 19401 40947 19402 41011
rect 19336 40946 19402 40947
rect 14585 37861 14651 37862
rect 14585 37797 14586 37861
rect 14650 37797 14651 37861
rect 14585 37796 14651 37797
rect 18790 37861 18856 37862
rect 18790 37797 18791 37861
rect 18855 37797 18856 37861
rect 18790 37796 18856 37797
rect 13830 31391 13896 31392
rect 13830 31327 13831 31391
rect 13895 31327 13896 31391
rect 13830 31326 13896 31327
rect 14586 30773 14650 37796
rect 19337 37311 19401 40946
rect 15229 37310 15295 37311
rect 15229 37246 15230 37310
rect 15294 37246 15295 37310
rect 15229 37245 15295 37246
rect 19336 37310 19402 37311
rect 19336 37246 19337 37310
rect 19401 37246 19402 37310
rect 19336 37245 19402 37246
rect 11965 30772 12031 30773
rect 11965 30708 11966 30772
rect 12030 30708 12031 30772
rect 11965 30707 12031 30708
rect 14585 30772 14651 30773
rect 14585 30708 14586 30772
rect 14650 30708 14651 30772
rect 14585 30707 14651 30708
rect 11966 28805 12030 30707
rect 11965 28804 12031 28805
rect 11965 28740 11966 28804
rect 12030 28740 12031 28804
rect 11965 28739 12031 28740
rect 11966 28734 12030 28739
rect 11346 26350 11412 26351
rect 11346 26286 11347 26350
rect 11411 26286 11412 26350
rect 11346 26285 11412 26286
rect 11836 26350 11902 26351
rect 11836 26286 11837 26350
rect 11901 26286 11902 26350
rect 11836 26285 11902 26286
rect 11347 26280 11411 26285
rect 11080 24203 11144 24209
rect 11079 24202 11145 24203
rect 11079 24138 11080 24202
rect 11144 24138 11145 24202
rect 11079 24137 11145 24138
rect 10632 20886 10698 20950
rect 11080 20886 11144 24137
rect 11837 22917 11901 26285
rect 13849 26009 13915 26010
rect 13849 25945 13850 26009
rect 13914 25945 13915 26009
rect 13849 25944 13915 25945
rect 13265 25598 13331 25599
rect 13265 25534 13266 25598
rect 13330 25534 13331 25598
rect 13265 25533 13331 25534
rect 12588 23211 12652 23220
rect 12587 23210 12653 23211
rect 12587 23146 12588 23210
rect 12652 23146 12653 23210
rect 12587 23145 12653 23146
rect 11836 22916 11902 22917
rect 11475 22915 11541 22916
rect 11475 22851 11476 22915
rect 11540 22851 11541 22915
rect 11836 22852 11837 22916
rect 11901 22852 11902 22916
rect 11836 22851 11902 22852
rect 11475 22850 11541 22851
rect 10632 20820 11144 20886
rect 11080 20335 11144 20820
rect 11079 20334 11145 20335
rect 11079 20270 11080 20334
rect 11144 20270 11145 20334
rect 11079 20269 11145 20270
rect 11476 19804 11540 22850
rect 12072 21656 12136 21664
rect 12071 21655 12137 21656
rect 12071 21591 12072 21655
rect 12136 21591 12137 21655
rect 12071 21590 12137 21591
rect 11475 19803 11541 19804
rect 11475 19739 11476 19803
rect 11540 19739 11541 19803
rect 11475 19738 11541 19739
rect -2399 19212 -2333 19213
rect -2399 19148 -2398 19212
rect -2334 19148 -2333 19212
rect -2399 19147 -2333 19148
rect -5280 19043 -5214 19044
rect -34861 18987 -34860 18993
rect -38169 18986 -34860 18987
rect -5280 18979 -5279 19043
rect -5215 18979 -5214 19043
rect -5280 18978 -5214 18979
rect -3919 19043 -3853 19044
rect -3919 18979 -3918 19043
rect -3854 18979 -3853 19043
rect -3919 18978 -3853 18979
rect -12356 17968 -12290 17969
rect -25453 17922 -25386 17923
rect -25453 17913 -25452 17922
rect -26708 17785 -25452 17913
rect -25453 17627 -25452 17785
rect -25387 17913 -25386 17922
rect -25387 17785 -25378 17913
rect -12356 17904 -12355 17968
rect -12291 17904 -12290 17968
rect -12356 17903 -12290 17904
rect -25387 17627 -25386 17785
rect -25453 17626 -25386 17627
rect -12355 17495 -12291 17903
rect -3212 17864 -2747 17865
rect -3212 17624 -3211 17864
rect -2748 17624 -2747 17864
rect -3212 17623 -2747 17624
rect -25451 17404 -25377 17405
rect -25451 17336 -25450 17404
rect -25454 17208 -25450 17336
rect -25451 17169 -25450 17208
rect -25378 17336 -25377 17404
rect -25378 17208 -24738 17336
rect -25378 17169 -25377 17208
rect -25451 17168 -25377 17169
rect -38741 16076 -34857 16078
rect -38741 16075 -34851 16076
rect -38741 15987 -38174 16075
rect -34852 15987 -34851 16075
rect -38741 15986 -34851 15987
rect -38741 15984 -34857 15986
rect -24866 15445 -24738 17208
rect -18719 17145 -17699 17209
rect -16119 17145 -15099 17209
rect -13519 17145 -12499 17209
rect -10417 17157 -10351 17158
rect -10912 17093 -10416 17157
rect -10352 17093 -10351 17157
rect -10417 17092 -10351 17093
rect -2398 16989 -2334 19147
rect 10231 19058 10297 19059
rect 10231 18994 10232 19058
rect 10296 18994 10297 19058
rect 10231 18993 10297 18994
rect -1505 18910 -1439 18911
rect -1505 18846 -1504 18910
rect -1440 18846 -1439 18910
rect -1505 18845 -1439 18846
rect -3928 16925 -2334 16989
rect -24866 15317 -23253 15445
rect -25518 14446 -25443 14447
rect -25518 14425 -25517 14446
rect -26701 14297 -25517 14425
rect -25518 14157 -25517 14297
rect -25444 14425 -25443 14446
rect -25444 14297 -25414 14425
rect -25444 14157 -25443 14297
rect -25518 14156 -25443 14157
rect -25519 13925 -25445 13926
rect -25519 13874 -25518 13925
rect -25520 13746 -25518 13874
rect -25519 13690 -25518 13746
rect -25446 13874 -25445 13925
rect -24866 13874 -24738 15317
rect -20013 14880 -19949 15900
rect -11255 14873 -11191 15893
rect -5787 15708 -5721 15709
rect -6755 15644 -5786 15708
rect -5722 15644 -5721 15708
rect -5787 15643 -5721 15644
rect -3928 15455 -3864 16925
rect -3510 16205 -3444 16206
rect -3510 16141 -3509 16205
rect -3445 16141 -3444 16205
rect -3510 16140 -3444 16141
rect -3929 15454 -3863 15455
rect -3929 15390 -3928 15454
rect -3864 15390 -3863 15454
rect -3929 15389 -3863 15390
rect -4903 14446 -4831 14447
rect -4903 14345 -4902 14446
rect -6758 14281 -4902 14345
rect -4903 14236 -4902 14281
rect -4832 14345 -4831 14446
rect -4832 14281 -4828 14345
rect -4832 14236 -4831 14281
rect -4903 14235 -4831 14236
rect -18224 14073 -18158 14074
rect -18224 14009 -18223 14073
rect -18159 14009 -17732 14073
rect -18224 14008 -18158 14009
rect -25446 13746 -24738 13874
rect -25446 13690 -25445 13746
rect -25519 13689 -25445 13690
rect -16124 13625 -15104 13689
rect -20013 12280 -19949 13300
rect -11255 12273 -11191 13293
rect -18722 10995 -17702 11059
rect -16122 10995 -15102 11059
rect -13522 10995 -12502 11059
rect -6163 10833 -5936 10834
rect -6163 10832 -6162 10833
rect -6758 10768 -6162 10832
rect -6163 10758 -6162 10768
rect -5937 10832 -5936 10833
rect -5937 10768 -5929 10832
rect -5937 10758 -5936 10768
rect -6163 10757 -5936 10758
rect -10971 10223 -10905 10224
rect -13942 10181 -13876 10182
rect -13942 10117 -13941 10181
rect -13877 10117 -13876 10181
rect -10971 10159 -10970 10223
rect -10906 10159 -10905 10223
rect -10971 10158 -10905 10159
rect -13942 10116 -13876 10117
rect -13941 9700 -13877 10116
rect -10970 9696 -10906 10158
rect -6168 9592 -5928 9593
rect -6168 9572 -6167 9592
rect -6748 9513 -6167 9572
rect -5929 9572 -5928 9592
rect -5929 9513 -5909 9572
rect -6748 9508 -5909 9513
rect -18719 9345 -17699 9409
rect -16119 9345 -15099 9409
rect -13519 9345 -12499 9409
rect -20013 7080 -19949 8100
rect -11255 7073 -11191 8093
rect -7215 7243 -6750 7244
rect -7215 7003 -7214 7243
rect -6751 7003 -6750 7243
rect -7215 7002 -6750 7003
rect -25522 6669 -25445 6670
rect -25522 6646 -25521 6669
rect -26709 6518 -25521 6646
rect -25522 6408 -25521 6518
rect -25446 6646 -25445 6669
rect -25446 6518 -25404 6646
rect -25446 6408 -25445 6518
rect -25522 6407 -25445 6408
rect -18252 6303 -18186 6304
rect -18252 6239 -18251 6303
rect -18187 6239 -17700 6303
rect -18252 6238 -18186 6239
rect -25523 6174 -25446 6175
rect -25523 5929 -25522 6174
rect -25447 6141 -25446 6174
rect -4911 6164 -4847 6176
rect -4911 6163 -4840 6164
rect -25447 5929 -25388 6141
rect -25523 5928 -25388 5929
rect -25516 4984 -25388 5928
rect -4911 5950 -4907 6163
rect -4841 5950 -4840 6163
rect -3928 6043 -3864 15389
rect -3509 14645 -3445 16140
rect -3134 14999 -3070 15001
rect -3145 14998 -3060 14999
rect -3145 14719 -3144 14998
rect -3061 14719 -3060 14998
rect -3145 14718 -3060 14719
rect -3510 14644 -3444 14645
rect -3510 14580 -3509 14644
rect -3445 14580 -3444 14644
rect -3510 14579 -3444 14580
rect -3929 6042 -3863 6043
rect -3929 5978 -3928 6042
rect -3864 5978 -3863 6042
rect -3929 5977 -3863 5978
rect -3928 5973 -3864 5977
rect -4911 5949 -4840 5950
rect -16124 5825 -15104 5889
rect -4911 5670 -4847 5949
rect -6748 5606 -4847 5670
rect -25516 4856 -23232 4984
rect -20013 4480 -19949 5500
rect -11255 4473 -11191 5493
rect -3509 5234 -3445 14579
rect -3134 14048 -3070 14718
rect -2736 13878 -2305 13942
rect -2369 12955 -2305 13878
rect -1809 13133 -1724 13134
rect -1809 12955 -1808 13133
rect -2369 12891 -1808 12955
rect -2369 11390 -2305 12891
rect -1809 12726 -1808 12891
rect -1725 12726 -1724 13133
rect -1809 12725 -1724 12726
rect -1760 11529 -1692 11530
rect -1760 11390 -1759 11529
rect -2369 11326 -1759 11390
rect -1760 11140 -1759 11326
rect -1693 11140 -1692 11529
rect -1760 11139 -1692 11140
rect -1760 9930 -1694 9931
rect -1760 9775 -1759 9930
rect -2390 9711 -1759 9775
rect -2390 8710 -2326 9711
rect -1760 9532 -1759 9711
rect -1695 9532 -1694 9930
rect -1760 9531 -1694 9532
rect -2738 8646 -2326 8710
rect -2390 8179 -2326 8646
rect -1759 8330 -1689 8331
rect -1759 8179 -1758 8330
rect -2390 8115 -1758 8179
rect -1759 7930 -1758 8115
rect -1690 7930 -1689 8330
rect -1759 7929 -1689 7930
rect -2736 6587 -2335 6651
rect -3194 5577 -3109 5578
rect -3194 5411 -3193 5577
rect -3201 5347 -3193 5411
rect -3194 5296 -3193 5347
rect -3110 5411 -3109 5577
rect -2399 5411 -2335 6587
rect -3110 5347 -2335 5411
rect -3110 5296 -3109 5347
rect -3194 5295 -3109 5296
rect -3510 5233 -3444 5234
rect -3510 5169 -3509 5233
rect -3445 5169 -3444 5233
rect -3510 5168 -3444 5169
rect -18722 3195 -17702 3259
rect -16122 3195 -15102 3259
rect -13522 3195 -12502 3259
rect -1504 -3060 -1440 18845
rect 8279 18718 8345 18719
rect 8279 18654 8280 18718
rect 8344 18654 8345 18718
rect 8279 18653 8345 18654
rect -1134 18651 -1068 18652
rect -1134 18587 -1133 18651
rect -1069 18587 -1068 18651
rect -1134 18586 -1068 18587
rect -1133 -2703 -1069 18586
rect -681 18312 -615 18313
rect -681 18248 -680 18312
rect -616 18248 -615 18312
rect -681 18247 -615 18248
rect -680 -2288 -616 18247
rect -285 18031 -219 18032
rect -285 17967 -284 18031
rect -220 17967 -219 18031
rect -285 17966 -219 17967
rect -284 -1862 -220 17966
rect 4294 17289 4360 17290
rect 6226 17289 6292 17290
rect 8280 17289 8344 18653
rect 4294 17225 4295 17289
rect 4359 17225 6227 17289
rect 6291 17225 8789 17289
rect 4294 17224 4360 17225
rect 6226 17224 6292 17225
rect 10232 17289 10296 18993
rect 9252 17225 10296 17289
rect 250 16446 4794 16447
rect 5256 16446 11140 16447
rect 250 16238 251 16446
rect 11139 16238 11140 16446
rect 250 16237 4792 16238
rect 5256 16237 11140 16238
rect 5477 14599 5657 14600
rect 5477 14598 5478 14599
rect 5257 14421 5478 14598
rect 5656 14598 5657 14599
rect 5656 14421 5667 14598
rect 5257 14420 5667 14421
rect 12072 12363 12136 21590
rect 12588 13171 12652 23145
rect 13266 17763 13330 25533
rect 13850 18571 13914 25944
rect 15230 24849 15294 37245
rect 19882 36729 19946 41317
rect 21517 40113 21581 45683
rect 22050 45671 22051 45735
rect 22115 45671 22116 45735
rect 22597 45677 22598 45741
rect 22662 45677 22663 45741
rect 22597 45676 22663 45677
rect 23142 45741 23208 45742
rect 23142 45677 23143 45741
rect 23207 45677 23208 45741
rect 23142 45676 23208 45677
rect 25862 45738 25928 45739
rect 22050 45670 22116 45671
rect 21516 40112 21582 40113
rect 21516 40048 21517 40112
rect 21581 40048 21582 40112
rect 21516 40047 21582 40048
rect 15989 36728 16055 36729
rect 15989 36664 15990 36728
rect 16054 36664 16055 36728
rect 15989 36663 16055 36664
rect 19881 36728 19947 36729
rect 19881 36664 19882 36728
rect 19946 36664 19947 36728
rect 19881 36663 19947 36664
rect 15229 24848 15295 24849
rect 15229 24784 15230 24848
rect 15294 24784 15295 24848
rect 15229 24783 15295 24784
rect 15990 24531 16054 36663
rect 21517 36051 21581 40047
rect 22051 39742 22115 45670
rect 22598 43923 22662 45676
rect 22597 43922 22663 43923
rect 22597 43858 22598 43922
rect 22662 43858 22663 43922
rect 22597 43857 22663 43858
rect 22050 39741 22116 39742
rect 22050 39677 22051 39741
rect 22115 39677 22116 39741
rect 22050 39676 22116 39677
rect 16720 36050 16786 36051
rect 16720 35986 16721 36050
rect 16785 35986 16786 36050
rect 16720 35985 16786 35986
rect 21516 36050 21582 36051
rect 21516 35986 21517 36050
rect 21581 35986 21582 36050
rect 21516 35985 21582 35986
rect 16721 29753 16785 35985
rect 22051 35344 22115 39676
rect 17411 35343 17477 35344
rect 17411 35279 17412 35343
rect 17476 35279 17477 35343
rect 17411 35278 17477 35279
rect 22050 35343 22116 35344
rect 22050 35279 22051 35343
rect 22115 35279 22116 35343
rect 22050 35278 22116 35279
rect 16720 29752 16786 29753
rect 16720 29688 16721 29752
rect 16785 29688 16786 29752
rect 16720 29687 16786 29688
rect 17412 29330 17476 35278
rect 22598 34584 22662 43857
rect 23143 43552 23207 45676
rect 25862 45674 25863 45738
rect 25927 45674 25928 45738
rect 26405 45678 26406 45742
rect 26470 45678 26471 45742
rect 29128 45738 29194 45739
rect 26405 45677 26471 45678
rect 26947 45736 27013 45737
rect 25862 45673 25928 45674
rect 25863 44892 25927 45673
rect 25862 44891 25928 44892
rect 25862 44827 25863 44891
rect 25927 44827 25928 44891
rect 25862 44826 25928 44827
rect 23142 43551 23208 43552
rect 23142 43487 23143 43551
rect 23207 43487 23208 43551
rect 23142 43486 23208 43487
rect 18251 34583 18317 34584
rect 18251 34519 18252 34583
rect 18316 34519 18317 34583
rect 18251 34518 18317 34519
rect 22597 34583 22663 34584
rect 22597 34519 22598 34583
rect 22662 34519 22663 34583
rect 22597 34518 22663 34519
rect 17411 29329 17477 29330
rect 17411 29265 17412 29329
rect 17476 29265 17477 29329
rect 17411 29264 17477 29265
rect 17412 29261 17476 29264
rect 15989 24530 16055 24531
rect 15989 24466 15990 24530
rect 16054 24466 16055 24530
rect 15989 24465 16055 24466
rect 18252 23519 18316 34518
rect 23143 33747 23207 43486
rect 25863 38419 25927 44826
rect 26406 44527 26470 45677
rect 26947 45672 26948 45736
rect 27012 45672 27013 45736
rect 26947 45671 27013 45672
rect 27504 45727 27570 45728
rect 26405 44526 26471 44527
rect 26405 44462 26406 44526
rect 26470 44462 26471 44526
rect 26405 44461 26471 44462
rect 25862 38418 25928 38419
rect 25862 38354 25863 38418
rect 25927 38354 25928 38418
rect 25862 38353 25928 38354
rect 26406 37839 26470 44461
rect 26948 41202 27012 45671
rect 27504 45663 27505 45727
rect 27569 45663 27570 45727
rect 29128 45674 29129 45738
rect 29193 45674 29194 45738
rect 30222 45735 30288 45736
rect 29128 45673 29194 45674
rect 29672 45731 29738 45732
rect 27504 45662 27570 45663
rect 26947 41201 27013 41202
rect 26947 41137 26948 41201
rect 27012 41137 27013 41201
rect 26947 41136 27013 41137
rect 26405 37838 26471 37839
rect 26405 37774 26406 37838
rect 26470 37774 26471 37838
rect 26405 37773 26471 37774
rect 26948 34523 27012 41136
rect 27505 40837 27569 45662
rect 27504 40836 27570 40837
rect 27504 40772 27505 40836
rect 27569 40772 27570 40836
rect 27504 40771 27570 40772
rect 26947 34522 27013 34523
rect 26947 34458 26948 34522
rect 27012 34458 27013 34522
rect 26947 34457 27013 34458
rect 27505 33814 27569 40771
rect 29129 39567 29193 45673
rect 29672 45667 29673 45731
rect 29737 45667 29738 45731
rect 29672 45666 29738 45667
rect 30222 45671 30223 45735
rect 30287 45671 30288 45735
rect 30222 45670 30288 45671
rect 30755 45735 30821 45736
rect 30755 45671 30756 45735
rect 30820 45671 30821 45735
rect 30755 45670 30821 45671
rect 29673 39932 29737 45666
rect 30222 43376 30286 45670
rect 30756 43742 30820 45670
rect 30755 43741 30821 43742
rect 30755 43677 30756 43741
rect 30820 43677 30821 43741
rect 30755 43676 30821 43677
rect 30221 43375 30287 43376
rect 30221 43311 30222 43375
rect 30286 43311 30287 43375
rect 30221 43310 30287 43311
rect 29672 39931 29738 39932
rect 29672 39867 29673 39931
rect 29737 39867 29738 39931
rect 29672 39866 29738 39867
rect 29128 39566 29194 39567
rect 29128 39502 29129 39566
rect 29193 39502 29194 39566
rect 29128 39501 29194 39502
rect 29129 35259 29193 39501
rect 29673 35971 29737 39866
rect 30222 36594 30286 43310
rect 30756 37230 30820 43676
rect 32413 38418 32479 38419
rect 32413 38354 32414 38418
rect 32478 38354 32479 38418
rect 32413 38353 32479 38354
rect 31823 37838 31889 37839
rect 31823 37774 31824 37838
rect 31888 37774 31889 37838
rect 31823 37773 31889 37774
rect 30755 37229 30821 37230
rect 30755 37165 30756 37229
rect 30820 37165 30821 37229
rect 30755 37164 30821 37165
rect 31230 37229 31296 37230
rect 31230 37165 31231 37229
rect 31295 37165 31296 37229
rect 31230 37164 31296 37165
rect 30221 36593 30287 36594
rect 30221 36529 30222 36593
rect 30286 36529 30287 36593
rect 30221 36528 30287 36529
rect 30583 36593 30649 36594
rect 30583 36529 30584 36593
rect 30648 36529 30649 36593
rect 30583 36528 30649 36529
rect 29672 35970 29738 35971
rect 29672 35906 29673 35970
rect 29737 35906 29738 35970
rect 29672 35905 29738 35906
rect 29989 35970 30055 35971
rect 29989 35906 29990 35970
rect 30054 35906 30055 35970
rect 29989 35905 30055 35906
rect 29128 35258 29194 35259
rect 29128 35194 29129 35258
rect 29193 35194 29194 35258
rect 29128 35193 29194 35194
rect 29406 35258 29472 35259
rect 29406 35194 29407 35258
rect 29471 35194 29472 35258
rect 29406 35193 29472 35194
rect 28827 34522 28893 34523
rect 28827 34458 28828 34522
rect 28892 34458 28893 34522
rect 28827 34457 28893 34458
rect 27504 33813 27570 33814
rect 27504 33749 27505 33813
rect 27569 33749 27570 33813
rect 27504 33748 27570 33749
rect 28314 33813 28380 33814
rect 28314 33749 28315 33813
rect 28379 33749 28380 33813
rect 28314 33748 28380 33749
rect 19254 33746 19320 33747
rect 19254 33682 19255 33746
rect 19319 33682 19320 33746
rect 19254 33681 19320 33682
rect 23142 33746 23208 33747
rect 23142 33682 23143 33746
rect 23207 33682 23208 33746
rect 23142 33681 23208 33682
rect 19255 23888 19319 33681
rect 25878 26009 25944 26010
rect 25878 25945 25879 26009
rect 25943 25945 25944 26009
rect 25878 25944 25944 25945
rect 19254 23887 19320 23888
rect 19254 23823 19255 23887
rect 19319 23823 19320 23887
rect 19254 23822 19320 23823
rect 18251 23518 18317 23519
rect 18251 23454 18252 23518
rect 18316 23454 18317 23518
rect 18251 23453 18317 23454
rect 23688 19382 23754 19383
rect 23688 19318 23689 19382
rect 23753 19318 23754 19382
rect 23688 19317 23754 19318
rect 14685 19278 14751 19279
rect 14685 19214 14686 19278
rect 14750 19214 14751 19278
rect 14685 19213 14751 19214
rect 14686 19095 14750 19213
rect 14686 19094 14753 19095
rect 14686 19030 16889 19094
rect 14114 18571 14180 18572
rect 13850 18507 14115 18571
rect 14179 18507 14180 18571
rect 14114 18506 14180 18507
rect 14367 17763 14433 17764
rect 13266 17699 14368 17763
rect 14432 17699 14433 17763
rect 14367 17698 14433 17699
rect 14689 17550 14753 19030
rect 23689 19083 23753 19317
rect 23689 19019 24903 19083
rect 23689 17553 23753 19019
rect 25613 18571 25679 18572
rect 25879 18571 25943 25944
rect 26462 25598 26528 25599
rect 26462 25534 26463 25598
rect 26527 25534 26528 25598
rect 26462 25533 26528 25534
rect 25613 18507 25614 18571
rect 25678 18507 25943 18571
rect 25613 18506 25679 18507
rect 25360 17764 25426 17765
rect 26463 17764 26527 25533
rect 27111 23211 27175 23222
rect 27110 23210 27176 23211
rect 27110 23146 27111 23210
rect 27175 23146 27176 23210
rect 27110 23145 27176 23146
rect 25360 17700 25361 17764
rect 25425 17700 26527 17764
rect 25360 17699 25426 17700
rect 23688 17552 23754 17553
rect 14688 17549 14754 17550
rect 14688 17485 14689 17549
rect 14753 17485 14754 17549
rect 23688 17488 23689 17552
rect 23753 17488 23754 17552
rect 23688 17487 23754 17488
rect 14688 17484 14754 17485
rect 23685 15788 23751 15789
rect 14686 15754 14824 15781
rect 14684 15753 14824 15754
rect 14684 15689 14685 15753
rect 14749 15689 14824 15753
rect 23685 15724 23686 15788
rect 23750 15724 23751 15788
rect 23685 15723 23751 15724
rect 14684 15688 14824 15689
rect 14685 15524 14824 15688
rect 14685 15423 16797 15524
rect 14685 13966 14824 15423
rect 23686 15473 23750 15723
rect 23686 15409 24905 15473
rect 23686 13998 23750 15409
rect 14684 13965 14824 13966
rect 14684 13901 14685 13965
rect 14749 13901 14824 13965
rect 23685 13997 23751 13998
rect 23685 13933 23686 13997
rect 23750 13933 23751 13997
rect 23685 13932 23751 13933
rect 14684 13900 14824 13901
rect 14114 13171 14180 13172
rect 12588 13107 14115 13171
rect 14179 13107 14180 13171
rect 14114 13106 14180 13107
rect 14367 12363 14433 12364
rect 12072 12299 14368 12363
rect 14432 12299 14433 12363
rect 14367 12298 14433 12299
rect 14685 12180 14824 13900
rect 27111 13171 27175 23145
rect 27657 21656 27721 21665
rect 27656 21655 27722 21656
rect 27656 21591 27657 21655
rect 27721 21591 27722 21655
rect 27656 21590 27722 21591
rect 25678 13107 27175 13171
rect 27657 12364 27721 21590
rect 25425 12300 27721 12364
rect 14685 12116 14702 12180
rect 14766 12116 14824 12180
rect 23690 12190 23756 12191
rect 23690 12126 23691 12190
rect 23755 12126 23756 12190
rect 23690 12125 23756 12126
rect 4629 11980 4783 11981
rect 4629 11802 4630 11980
rect 4629 11801 4783 11802
rect 10804 10538 12783 10617
rect 6482 10537 12783 10538
rect 6482 10356 6483 10537
rect 11218 10439 12783 10537
rect 11218 10356 11338 10439
rect 13246 10439 13289 10617
rect 6482 10355 11338 10356
rect 10804 10326 11338 10355
rect 14685 10383 14824 12116
rect 23691 11890 23755 12125
rect 23691 11826 24893 11890
rect 14685 10350 14691 10383
rect 14690 10319 14691 10350
rect 14755 10350 14824 10383
rect 23691 10381 23755 11826
rect 23690 10380 23756 10381
rect 14755 10319 14756 10350
rect 14690 10318 14756 10319
rect 23690 10316 23691 10380
rect 23755 10316 23756 10380
rect 23690 10315 23756 10316
rect 13875 10150 21119 10151
rect 371 10144 792 10145
rect 1255 10144 1813 10145
rect 371 10003 372 10144
rect 1812 10003 1813 10144
rect 371 10002 792 10003
rect 1255 10002 1813 10003
rect 4603 10136 6206 10143
rect 4603 10135 11723 10136
rect 4603 9990 5727 10135
rect 11722 9990 11723 10135
rect 13875 9993 13876 10150
rect 21118 9993 21119 10150
rect 13875 9992 16808 9993
rect 4603 9989 8768 9990
rect 28 9830 213 9831
rect 28 5570 29 9830
rect 212 7975 213 9830
rect 4603 9829 6206 9989
rect 9231 9989 11723 9990
rect 4603 8366 4917 9829
rect 14204 9590 14475 9992
rect 17271 9992 21119 9993
rect 4603 8188 4679 8366
rect 4857 8188 4917 8366
rect 212 7960 1288 7975
rect 212 7720 805 7960
rect 1268 7720 1288 7960
rect 212 7696 1288 7720
rect 212 5570 213 7696
rect 28 5569 213 5570
rect 4603 6366 4917 8188
rect 4603 6188 4679 6366
rect 4857 6188 4917 6366
rect 13303 9319 14475 9590
rect 13303 6491 13574 9319
rect 13303 6313 13350 6491
rect 13528 6313 13574 6491
rect 13303 6266 13574 6313
rect 17605 8451 17876 9992
rect 17605 8273 17646 8451
rect 17824 8273 17876 8451
rect 17605 6451 17876 8273
rect 17605 6273 17646 6451
rect 17824 6273 17876 6451
rect 4603 4366 4917 6188
rect 17605 5138 17876 6273
rect 21249 7514 21418 7515
rect 21249 5846 21250 7514
rect 21239 5552 21250 5846
rect 16014 5088 19356 5138
rect 16014 4910 16101 5088
rect 16279 4910 19101 5088
rect 19279 4910 19356 5088
rect 16014 4867 19356 4910
rect 21249 4540 21250 5552
rect 21417 5846 21418 7514
rect 21417 5552 24797 5846
rect 21417 4540 21418 5552
rect 25260 5552 25309 5846
rect 21249 4539 21418 4540
rect 4603 4188 4679 4366
rect 4857 4188 4917 4366
rect 27 2773 191 2774
rect 27 359 28 2773
rect 190 2308 191 2773
rect 4603 2366 4917 4188
rect 190 2273 1289 2308
rect 190 2033 778 2273
rect 1241 2033 1289 2273
rect 190 2012 1289 2033
rect 4603 2188 4679 2366
rect 4857 2188 4917 2366
rect 190 359 191 2012
rect 27 358 191 359
rect 321 232 794 233
rect 4603 233 4917 2188
rect 12169 2773 12420 2815
rect 12169 2595 12207 2773
rect 12385 2595 12420 2773
rect 1257 232 8814 233
rect 12169 233 12420 2595
rect 21242 2139 21420 2140
rect 21242 1649 21243 2139
rect 21228 1336 21243 1649
rect 21242 1288 21243 1336
rect 21419 1649 21420 2139
rect 21419 1606 25325 1649
rect 21419 1366 24796 1606
rect 25259 1366 25325 1606
rect 21419 1336 25325 1366
rect 21419 1288 21420 1336
rect 21242 1287 21420 1288
rect 9277 232 16791 233
rect 17254 232 21108 233
rect 321 67 322 232
rect 21107 67 21108 232
rect 321 66 21108 67
rect 28315 -1862 28379 33748
rect -284 -1926 28379 -1862
rect 28828 -2288 28892 34457
rect -680 -2352 28892 -2288
rect 29407 -2703 29471 35193
rect -1133 -2767 29471 -2703
rect 29990 -3060 30054 35905
rect -1504 -3124 30054 -3060
rect 21201 -3509 21267 -3508
rect 30584 -3509 30648 36528
rect 21201 -3573 21202 -3509
rect 21266 -3573 30648 -3509
rect 21201 -3574 21267 -3573
rect 21201 -3981 21267 -3980
rect 31231 -3981 31295 37164
rect 21201 -4045 21202 -3981
rect 21266 -4045 31295 -3981
rect 21201 -4046 21267 -4045
rect 21201 -4516 21267 -4515
rect 31824 -4516 31888 37773
rect 21201 -4580 21202 -4516
rect 21266 -4580 31888 -4516
rect 21201 -4581 21267 -4580
rect 21201 -4979 21267 -4978
rect 32414 -4979 32478 38353
rect 33254 23984 35216 24048
rect 35152 23867 35216 23984
rect 35151 23866 35217 23867
rect 35151 23802 35152 23866
rect 35216 23802 35217 23866
rect 35151 23801 35217 23802
rect 35151 21585 35217 21586
rect 33253 21521 35152 21585
rect 35216 21521 35217 21585
rect 35151 21520 35217 21521
rect 35477 21380 35541 68015
rect 36066 24019 36130 68638
rect 36065 24018 36131 24019
rect 36065 23954 36066 24018
rect 36130 23954 36131 24018
rect 36065 23953 36131 23954
rect 35476 21379 35542 21380
rect 35476 21315 35477 21379
rect 35541 21315 35542 21379
rect 35476 21314 35542 21315
rect 35477 8532 35541 21314
rect 36066 9155 36130 23953
rect 36065 9154 36131 9155
rect 36065 9090 36066 9154
rect 36130 9090 36131 9154
rect 36065 9089 36131 9090
rect 35477 8531 35554 8532
rect 35477 8467 35489 8531
rect 35553 8467 35554 8531
rect 35477 8466 35554 8467
rect 35027 7223 35093 7224
rect 33256 7159 35028 7223
rect 35092 7159 35093 7223
rect 35027 7158 35093 7159
rect 35026 5885 35092 5886
rect 33247 5821 35027 5885
rect 35091 5821 35092 5885
rect 35026 5820 35092 5821
rect 35034 4492 35100 4493
rect 33253 4428 35035 4492
rect 35099 4428 35100 4492
rect 35034 4427 35100 4428
rect 35030 3122 35096 3123
rect 33249 3058 35031 3122
rect 35095 3058 35096 3122
rect 35030 3057 35096 3058
rect 35477 1592 35541 8466
rect 36066 2215 36130 9089
rect 36631 8470 36695 69258
rect 44736 45174 45324 45179
rect 44736 45074 44795 45174
rect 45258 45074 45324 45174
rect 44736 45007 44754 45074
rect 45306 45007 45324 45074
rect 44736 44934 44795 45007
rect 45258 44934 45324 45007
rect 44736 44931 45324 44934
rect 41587 44528 41827 44551
rect 41515 44527 41875 44528
rect 41515 44462 41516 44527
rect 41874 44462 41875 44527
rect 41515 44461 41875 44462
rect 41587 44304 41827 44461
rect 41263 44064 41827 44304
rect 41587 43378 41827 44064
rect 44765 43925 44795 43926
rect 45258 43925 45294 43926
rect 44765 43854 44766 43925
rect 45293 43854 45294 43925
rect 44765 43853 44795 43854
rect 45258 43853 45294 43854
rect 41513 43377 41873 43378
rect 41513 43312 41514 43377
rect 41872 43312 41873 43377
rect 41513 43311 41873 43312
rect 41587 43295 41827 43311
rect 44755 41383 44779 41384
rect 45242 41383 45284 41384
rect 44755 41312 44756 41383
rect 45283 41312 45284 41383
rect 44755 41311 44779 41312
rect 45242 41311 45284 41312
rect 41494 40837 41734 40855
rect 41431 40836 41791 40837
rect 41431 40771 41432 40836
rect 41790 40771 41791 40836
rect 41431 40770 41791 40771
rect 41494 40559 41734 40770
rect 41271 40319 41734 40559
rect 41494 39568 41734 40319
rect 44755 40113 44772 40114
rect 45235 40113 45284 40114
rect 44755 40042 44756 40113
rect 45283 40042 45284 40113
rect 44755 40041 44772 40042
rect 45235 40041 45284 40042
rect 41429 39567 41789 39568
rect 41429 39502 41430 39567
rect 41788 39502 41789 39567
rect 41429 39501 41789 39502
rect 41494 39483 41734 39501
rect 42785 24174 44801 24252
rect 45264 24174 46299 24252
rect 42785 24065 42856 24174
rect 46190 24065 46299 24174
rect 42785 24012 44801 24065
rect 45264 24012 46299 24065
rect 37661 23714 40175 23728
rect 37661 23611 39346 23714
rect 37661 23492 37819 23611
rect 37892 23493 39346 23611
rect 39420 23493 40175 23714
rect 37892 23492 40175 23493
rect 37661 23488 40175 23492
rect 39334 23200 39422 23201
rect 37818 23194 37906 23195
rect 37818 23190 37819 23194
rect 37274 22954 37819 23190
rect 37274 22816 37510 22954
rect 37818 22946 37819 22954
rect 37905 23190 37906 23194
rect 39334 23190 39335 23200
rect 37905 22954 39335 23190
rect 37905 22946 37906 22954
rect 39334 22952 39335 22954
rect 39421 23190 39422 23200
rect 39421 22954 39497 23190
rect 39421 22952 39422 22954
rect 39334 22951 39422 22952
rect 37818 22945 37906 22946
rect 36913 22815 37510 22816
rect 36913 22579 36914 22815
rect 37156 22580 37510 22815
rect 37156 22579 37157 22580
rect 36913 22578 37157 22579
rect 37274 21827 37510 22580
rect 39935 22732 40175 23488
rect 39935 22492 40801 22732
rect 39935 22402 40175 22492
rect 37732 22388 40175 22402
rect 37732 22280 39346 22388
rect 37732 22162 37826 22280
rect 37825 22151 37826 22162
rect 37896 22167 39346 22280
rect 39420 22167 40175 22388
rect 37896 22162 40175 22167
rect 37896 22151 37897 22162
rect 37825 22150 37897 22151
rect 39340 21834 39428 21835
rect 39340 21827 39341 21834
rect 37274 21823 39341 21827
rect 37274 21621 37814 21823
rect 37899 21621 39341 21823
rect 37274 21591 39341 21621
rect 39340 21586 39341 21591
rect 39427 21827 39428 21834
rect 39427 21591 39497 21827
rect 39427 21586 39428 21591
rect 39340 21585 39428 21586
rect 42729 21178 48791 21244
rect 42729 21069 42854 21178
rect 46188 21069 48791 21178
rect 42729 21005 48791 21069
rect 42729 21004 49031 21005
rect 36630 8469 36696 8470
rect 36630 8405 36631 8469
rect 36695 8405 36696 8469
rect 36630 8404 36696 8405
rect 36065 2214 36131 2215
rect 36065 2150 36066 2214
rect 36130 2150 36131 2214
rect 36065 2149 36131 2150
rect 36066 2136 36130 2149
rect 35477 1591 35554 1592
rect 35477 1527 35489 1591
rect 35553 1527 35554 1591
rect 36631 1530 36695 8404
rect 36971 7350 37067 8537
rect 37895 7593 38131 8554
rect 37895 7563 38667 7593
rect 37895 7375 38568 7563
rect 38649 7375 38667 7563
rect 37895 7357 38667 7375
rect 39402 7590 39638 8553
rect 39402 7576 40189 7590
rect 39402 7388 40087 7576
rect 40168 7388 40189 7576
rect 36970 7349 37068 7350
rect 36970 7253 36971 7349
rect 37067 7253 37068 7349
rect 36970 7252 37068 7253
rect 36971 6525 37067 7252
rect 37895 7138 38131 7357
rect 37894 6902 38131 7138
rect 37895 6525 38131 6902
rect 39402 7354 40189 7388
rect 39402 6525 39638 7354
rect 42601 7232 44796 7233
rect 45259 7232 45924 7233
rect 40800 7170 41265 7171
rect 40800 6930 40801 7170
rect 41264 6930 41265 7170
rect 42601 7143 42602 7232
rect 45923 7143 45924 7232
rect 42601 7142 45924 7143
rect 40800 6929 41265 6930
rect 37180 6289 39638 6525
rect 36970 6265 37068 6289
rect 36970 6169 36971 6265
rect 37067 6169 37068 6265
rect 36970 6168 37068 6169
rect 36971 5178 37067 6168
rect 36970 5177 37068 5178
rect 36970 5109 36971 5177
rect 37067 5109 37068 5177
rect 37895 5109 38131 6289
rect 38562 6232 38646 6289
rect 38562 6044 38563 6232
rect 38644 6205 38646 6232
rect 39402 6275 39638 6289
rect 39402 6229 40175 6275
rect 38644 6044 38645 6205
rect 38562 6043 38645 6044
rect 39402 6041 40092 6229
rect 40173 6041 40175 6229
rect 39402 6039 40175 6041
rect 39402 5109 39638 6039
rect 37141 4879 39638 5109
rect 37141 4873 38562 4879
rect 36971 4090 37067 4873
rect 36971 4089 37069 4090
rect 36971 3993 36972 4089
rect 37068 3993 37069 4089
rect 36971 3992 37069 3993
rect 36971 2832 37067 3992
rect 37895 3500 38131 4873
rect 38561 4691 38562 4873
rect 38643 4873 39638 4879
rect 38643 4691 38644 4873
rect 38561 4690 38644 4691
rect 39402 4857 40189 4873
rect 39402 4669 40092 4857
rect 40173 4669 40189 4857
rect 39402 4637 40189 4669
rect 39402 3503 39638 4637
rect 40798 4267 41263 4268
rect 40798 4027 40799 4267
rect 41262 4233 46002 4267
rect 41262 4144 42599 4233
rect 45959 4144 46002 4233
rect 41262 4027 46002 4144
rect 40798 4026 41263 4027
rect 37895 3480 38646 3500
rect 37895 3479 38647 3480
rect 37895 3291 38565 3479
rect 38646 3291 38647 3479
rect 37895 3290 38647 3291
rect 39402 3473 40187 3503
rect 37895 3264 38646 3290
rect 39402 3285 40089 3473
rect 40170 3285 40187 3473
rect 39402 3267 40187 3285
rect 37895 2750 38131 3264
rect 39402 2820 39638 3267
rect 35477 1526 35554 1527
rect 36630 1529 36696 1530
rect 35477 1493 35541 1526
rect 36630 1465 36631 1529
rect 36695 1465 36696 1529
rect 36630 1464 36696 1465
rect 36631 1436 36695 1464
rect 36971 410 37067 1597
rect 37895 653 38131 1614
rect 37895 623 38667 653
rect 37895 435 38568 623
rect 38649 435 38667 623
rect 37895 417 38667 435
rect 39402 650 39638 1613
rect 39402 636 40189 650
rect 39402 448 40087 636
rect 40168 448 40189 636
rect 36970 409 37068 410
rect 36970 313 36971 409
rect 37067 313 37068 409
rect 36970 312 37068 313
rect 35027 283 35093 284
rect 33256 219 35028 283
rect 35092 219 35093 283
rect 35027 218 35093 219
rect 36971 -415 37067 312
rect 37895 198 38131 417
rect 37894 -38 38131 198
rect 37895 -415 38131 -38
rect 39402 414 40189 448
rect 39402 -415 39638 414
rect 42598 309 44799 310
rect 45262 309 45931 310
rect 40800 230 41265 231
rect 40800 -10 40801 230
rect 41264 -10 41265 230
rect 42598 199 42599 309
rect 45930 199 45931 309
rect 42598 198 45931 199
rect 40800 -11 41265 -10
rect 37180 -651 39638 -415
rect 36970 -675 37068 -651
rect 36970 -771 36971 -675
rect 37067 -771 37068 -675
rect 36970 -772 37068 -771
rect 35026 -1055 35092 -1054
rect 33247 -1119 35027 -1055
rect 35091 -1119 35092 -1055
rect 35026 -1120 35092 -1119
rect 36971 -1762 37067 -772
rect 36970 -1763 37068 -1762
rect 36970 -1831 36971 -1763
rect 37067 -1831 37068 -1763
rect 37895 -1831 38131 -651
rect 38562 -708 38646 -651
rect 38562 -896 38563 -708
rect 38644 -735 38646 -708
rect 39402 -665 39638 -651
rect 39402 -711 40175 -665
rect 38644 -896 38645 -735
rect 38562 -897 38645 -896
rect 39402 -899 40092 -711
rect 40173 -899 40175 -711
rect 39402 -901 40175 -899
rect 39402 -1831 39638 -901
rect 37141 -2061 39638 -1831
rect 37141 -2067 38562 -2061
rect 35034 -2448 35100 -2447
rect 33253 -2512 35035 -2448
rect 35099 -2512 35100 -2448
rect 35034 -2513 35100 -2512
rect 36971 -2850 37067 -2067
rect 36971 -2851 37069 -2850
rect 36971 -2947 36972 -2851
rect 37068 -2947 37069 -2851
rect 36971 -2948 37069 -2947
rect 35030 -3818 35096 -3817
rect 33249 -3882 35031 -3818
rect 35095 -3882 35096 -3818
rect 35030 -3883 35096 -3882
rect 36971 -4108 37067 -2948
rect 37895 -3440 38131 -2067
rect 38561 -2249 38562 -2067
rect 38643 -2067 39638 -2061
rect 38643 -2249 38644 -2067
rect 38561 -2250 38644 -2249
rect 39402 -2083 40189 -2067
rect 39402 -2271 40092 -2083
rect 40173 -2271 40189 -2083
rect 39402 -2303 40189 -2271
rect 39402 -3437 39638 -2303
rect 40798 -2673 41263 -2672
rect 40798 -2680 40799 -2673
rect 41262 -2680 41517 -2673
rect 41262 -2708 46063 -2680
rect 41262 -2796 42587 -2708
rect 45933 -2796 46063 -2708
rect 41262 -2913 46063 -2796
rect 41248 -2920 46063 -2913
rect 37895 -3460 38646 -3440
rect 37895 -3461 38647 -3460
rect 37895 -3649 38565 -3461
rect 38646 -3649 38647 -3461
rect 37895 -3650 38647 -3649
rect 39402 -3467 40187 -3437
rect 37895 -3676 38646 -3650
rect 39402 -3655 40089 -3467
rect 40170 -3655 40187 -3467
rect 39402 -3673 40187 -3655
rect 37895 -4190 38131 -3676
rect 39402 -4120 39638 -3673
rect 21201 -5043 21202 -4979
rect 21266 -5043 32478 -4979
rect 21201 -5044 21267 -5043
rect -2735 -6413 -487 -6173
rect -3596 -6822 -3502 -6821
rect -3596 -8276 -3595 -6822
rect -6741 -8516 -3595 -8276
rect -3596 -10130 -3595 -8516
rect -3503 -8276 -3502 -6822
rect -600 -6824 -487 -6413
rect -601 -6825 -485 -6824
rect -3503 -8516 -3494 -8276
rect -3503 -10130 -3502 -8516
rect -3596 -10131 -3502 -10130
rect -601 -10140 -600 -6825
rect -486 -10140 -485 -6825
rect -601 -10141 -485 -10140
rect -57093 -18021 -55093 -16021
rect -53093 -18021 -43285 -16021
rect -42665 -18021 -35285 -16021
rect -34665 -18021 -27285 -16021
rect -26665 -18021 -19285 -16021
rect -18665 -18021 -11285 -16021
rect -10665 -18021 -3285 -16021
rect -2665 -18021 4715 -16021
rect 5335 -18021 12715 -16021
rect 13335 -18021 20715 -16021
rect 21335 -18021 28715 -16021
rect 29335 -18021 36715 -16021
rect 37335 -18021 44715 -16021
rect 45335 -18021 54907 -16021
rect 56907 -18021 62907 -16021
rect -57093 -22021 -51093 -20021
rect -49093 -22021 -39285 -20021
rect -38665 -22021 -31285 -20021
rect -30665 -22021 -23285 -20021
rect -22665 -22021 -15285 -20021
rect -14665 -22021 -7285 -20021
rect -6665 -22021 715 -20021
rect 1335 -22021 8715 -20021
rect 9335 -22021 16715 -20021
rect 17335 -22021 24715 -20021
rect 25335 -22021 32715 -20021
rect 33335 -22021 40715 -20021
rect 41335 -22021 48715 -20021
rect 49335 -22021 58907 -20021
rect 60907 -22021 62907 -20021
<< via4 >>
rect -55093 86442 -53093 88442
rect -43285 86442 -42665 88442
rect -35285 86442 -34665 88442
rect -27285 86442 -26665 88442
rect -19285 86442 -18665 88442
rect -11285 86442 -10665 88442
rect -3285 86442 -2665 88442
rect 4715 86442 5335 88442
rect 12715 86442 13335 88442
rect 20715 86442 21335 88442
rect 28715 86442 29335 88442
rect 36715 86442 37335 88442
rect 44715 86442 45335 88442
rect 54907 86442 56907 88442
rect -51093 82442 -49093 84442
rect -39285 82442 -38665 84442
rect -31285 82442 -30665 84442
rect -23285 82442 -22665 84442
rect -15285 82442 -14665 84442
rect -7285 82442 -6665 84442
rect 715 82442 1335 84442
rect 8715 82442 9335 84442
rect 16715 82442 17335 84442
rect 24715 82442 25335 84442
rect 32715 82442 33335 84442
rect 40715 82442 41335 84442
rect 48715 82442 49335 84442
rect 58907 82442 60907 84442
rect -19241 74828 -18711 75068
rect -15243 75013 -14713 75253
rect 12758 74932 13288 75172
rect 16757 74924 17287 75164
rect -15242 70754 -14712 70994
rect -19241 69997 -18711 70237
rect -15239 68675 -14709 68915
rect -19245 66882 -18715 67122
rect -11071 63205 -10737 63557
rect 20763 64191 21288 64719
rect 28757 64197 29282 64725
rect -6939 62966 -6699 63206
rect -3241 63171 -2711 63411
rect 757 62992 1287 63232
rect 16766 62200 17291 62728
rect 24762 62193 25287 62721
rect 32765 62189 33290 62717
rect -19238 50450 -18708 50690
rect -27236 49720 -26706 49826
rect -27236 49656 -27070 49720
rect -27070 49656 -26726 49720
rect -26726 49656 -26706 49720
rect -27236 49586 -26706 49656
rect -23234 48983 -22704 49223
rect -27162 42916 -27087 43156
rect -27087 42916 -26990 43156
rect -26990 42916 -26709 43156
rect -6978 54706 -6706 55397
rect -3237 54182 -2707 54422
rect 756 59884 1286 60124
rect 8761 59873 9291 60113
rect 756 56509 1286 56749
rect 8760 56498 9290 56738
rect 756 53134 1286 53374
rect 8760 53123 9290 53363
rect -7237 51461 -6707 51701
rect -27162 39710 -27077 39950
rect -27077 39710 -26990 39950
rect -26990 39710 -26699 39950
rect -35218 38258 -34755 38498
rect -31206 38269 -30743 38509
rect -31218 37171 -30755 37411
rect -23192 37540 -22729 38013
rect -27162 35641 -27077 35881
rect -27077 35641 -26996 35881
rect -26996 35641 -26699 35881
rect -3231 51074 -2701 51101
rect -3231 50896 -2701 51074
rect -3231 50861 -2701 50896
rect -3237 48533 -2707 48773
rect 756 49759 1286 49999
rect 8760 49748 9290 49988
rect 20763 60191 21288 60719
rect 28757 60197 29282 60725
rect 16766 58200 17291 58728
rect 24762 58193 25287 58721
rect 32765 58189 33290 58717
rect 20763 56191 21288 56719
rect 28757 56197 29282 56725
rect 16766 54200 17291 54728
rect 24762 54193 25287 54721
rect 32765 54189 33290 54717
rect 20763 52191 21288 52719
rect 28757 52197 29282 52725
rect 16766 50200 17291 50728
rect 24762 50193 25287 50721
rect 32765 50189 33290 50717
rect 20763 48191 21288 48719
rect 28757 48197 29282 48725
rect -3248 45115 -2718 45355
rect 752 44274 1282 44514
rect 8760 42998 9290 43238
rect -3233 39846 -2703 39886
rect -3233 39666 -2703 39846
rect 762 40629 1292 40869
rect -3233 39646 -2703 39666
rect 756 39200 1286 39440
rect -27162 32527 -27084 32767
rect -27084 32527 -27005 32767
rect -27005 32527 -26704 32767
rect -19238 28468 -18708 28708
rect -15234 27203 -14704 27443
rect -35224 26668 -34761 26908
rect -11237 27815 -10707 28055
rect -19246 25804 -18716 25810
rect -19246 25571 -19088 25804
rect -19088 25571 -18855 25804
rect -18855 25571 -18716 25804
rect -19246 25570 -18716 25571
rect -15238 25578 -14708 25818
rect -27228 25274 -26698 25514
rect -23236 24677 -22706 24917
rect -39205 23474 -38742 23714
rect -19239 23490 -18709 23730
rect -15237 23399 -14707 23639
rect -11246 22914 -10716 23154
rect -35218 19065 -34755 19233
rect -35218 18993 -34861 19065
rect -34861 18993 -34755 19065
rect 4761 37813 5291 38053
rect 757 36855 1287 37095
rect 4768 36420 5298 36660
rect 774 35776 1304 36016
rect 8758 35788 9288 36028
rect 4774 35242 5304 35482
rect 4780 22919 5243 23159
rect 8774 23356 9237 23495
rect 8774 23255 8787 23356
rect 8787 23255 8943 23356
rect 8943 23255 9237 23356
rect 16766 46200 17291 46728
rect 24762 46193 25287 46721
rect 32765 46189 33290 46717
rect 4797 19173 5260 19233
rect -27238 17723 -26708 17963
rect -3211 17624 -2748 17864
rect -39204 15960 -38741 16200
rect 4797 19027 4857 19173
rect 4857 19027 5194 19173
rect 5194 19027 5260 19173
rect 4797 18993 5260 19027
rect -27231 14237 -26701 14477
rect -23253 15250 -22723 15490
rect -7218 15572 -6755 15812
rect -3201 16210 -2738 16450
rect -7221 14212 -6758 14452
rect -7221 10672 -6758 10912
rect -7211 9422 -6748 9662
rect -7214 7003 -6751 7243
rect -27239 6470 -26709 6710
rect -7211 5524 -6748 5764
rect -23232 4804 -22702 5044
rect -3199 13808 -2736 14048
rect -3201 8707 -2738 8802
rect -3201 8643 -3185 8707
rect -3185 8643 -3121 8707
rect -3121 8643 -2738 8707
rect -3201 8562 -2738 8643
rect -3199 6649 -2736 6743
rect -3199 6585 -3184 6649
rect -3184 6585 -3120 6649
rect -3120 6585 -2736 6649
rect -3199 6503 -2736 6585
rect 789 17525 1252 17618
rect 789 17461 981 17525
rect 981 17461 1045 17525
rect 1045 17461 1252 17525
rect 789 17378 1252 17461
rect 8789 17163 9252 17403
rect 4794 16446 5256 16746
rect 4794 16430 5256 16446
rect 4792 16238 5256 16430
rect 4792 16190 5256 16238
rect 4794 15884 5256 16190
rect 4794 14381 5257 14621
rect 12861 21027 13103 21097
rect 12861 20963 12936 21027
rect 12936 20963 13000 21027
rect 13000 20963 13103 21027
rect 12861 20855 13103 20963
rect 12849 18688 13091 18796
rect 12849 18624 12930 18688
rect 12930 18624 12994 18688
rect 12994 18624 13091 18688
rect 12849 18554 13091 18624
rect 16889 18946 17131 19188
rect 20893 19062 21135 19161
rect 20893 18998 20971 19062
rect 20971 18998 21035 19062
rect 21035 18998 21135 19062
rect 20893 18919 21135 18998
rect 24903 18914 25145 19156
rect 12843 17083 13085 17191
rect 12843 17019 12956 17083
rect 12956 17019 13020 17083
rect 13020 17019 13085 17083
rect 12843 16949 13085 17019
rect 12862 15228 13104 15320
rect 12862 15164 12973 15228
rect 12973 15164 13037 15228
rect 13037 15164 13104 15228
rect 12862 15078 13104 15164
rect 16797 15353 17039 15595
rect 20836 15496 21078 15590
rect 20836 15432 20928 15496
rect 20928 15432 20992 15496
rect 20992 15432 21078 15496
rect 20836 15348 21078 15432
rect 24905 15321 25147 15563
rect 12884 13528 13126 13619
rect 12884 13464 13003 13528
rect 13003 13464 13067 13528
rect 13067 13464 13126 13528
rect 12884 13377 13126 13464
rect 4783 11980 5246 12013
rect 4783 11802 4808 11980
rect 4808 11802 5246 11980
rect 4783 11773 5246 11802
rect 12897 11676 13139 11764
rect 12897 11612 13001 11676
rect 13001 11612 13065 11676
rect 13065 11612 13139 11676
rect 12897 11522 13139 11612
rect 12783 10413 13246 10653
rect 20890 11906 21132 12002
rect 20890 11842 20985 11906
rect 20985 11842 21049 11906
rect 21049 11842 21132 11906
rect 20890 11760 21132 11842
rect 24893 11730 25135 11972
rect 792 10144 1255 10149
rect 792 10003 1255 10144
rect 792 9909 1255 10003
rect 8768 9990 9231 10124
rect 16808 9993 17271 10139
rect 8768 9884 9231 9990
rect 16808 9899 17271 9993
rect 805 7720 1268 7960
rect 24797 5410 25260 5982
rect 778 2033 1241 2273
rect 794 232 1257 325
rect 8814 232 9277 337
rect 24796 1366 25259 1606
rect 16791 232 17254 325
rect 794 85 1257 232
rect 8814 97 9277 232
rect 16791 85 17254 232
rect 32791 23894 33254 24134
rect 32790 21434 33253 21674
rect 32793 7053 33256 7293
rect 32784 5753 33247 5993
rect 32790 4338 33253 4578
rect 32786 2965 33249 3205
rect 44795 45074 45258 45174
rect 44795 45007 45258 45074
rect 44795 44934 45258 45007
rect 40800 44064 41263 44304
rect 44795 43925 45258 44013
rect 44795 43854 45258 43925
rect 44795 43773 45258 43854
rect 44779 41383 45242 41504
rect 44779 41312 45242 41383
rect 44779 41264 45242 41312
rect 40808 40319 41271 40559
rect 44772 40113 45235 40193
rect 44772 40042 45235 40113
rect 44772 39953 45235 40042
rect 44801 24174 45264 24252
rect 44801 24065 45264 24174
rect 44801 24012 45264 24065
rect 36914 22579 37156 22815
rect 40801 22492 41264 22732
rect 48791 21005 49254 21245
rect 36881 8792 37155 8810
rect 36881 8556 36898 8792
rect 36898 8556 37140 8792
rect 37140 8556 37155 8792
rect 36881 8537 37155 8556
rect 44796 7232 45259 7446
rect 40801 6930 41264 7170
rect 44796 7206 45259 7232
rect 36938 6289 37180 6525
rect 36899 5081 36971 5109
rect 36971 5081 37067 5109
rect 37067 5081 37141 5109
rect 36899 4873 37141 5081
rect 40799 4027 41262 4267
rect 36889 2559 37163 2832
rect 36881 1852 37155 1870
rect 36881 1616 36898 1852
rect 36898 1616 37140 1852
rect 37140 1616 37155 1852
rect 36881 1597 37155 1616
rect 32793 113 33256 353
rect 44799 309 45262 521
rect 40801 -10 41264 230
rect 44799 281 45262 309
rect 36938 -651 37180 -415
rect 32784 -1187 33247 -947
rect 36899 -1859 36971 -1831
rect 36971 -1859 37067 -1831
rect 37067 -1859 37141 -1831
rect 36899 -2067 37141 -1859
rect 32790 -2602 33253 -2362
rect 32786 -3975 33249 -3735
rect 40785 -2913 40799 -2680
rect 40799 -2913 41262 -2673
rect 40785 -2920 41248 -2913
rect 36889 -4381 37163 -4108
rect -3198 -6413 -2735 -6173
rect -7204 -8516 -6741 -8276
rect -55093 -18021 -53093 -16021
rect -43285 -18021 -42665 -16021
rect -35285 -18021 -34665 -16021
rect -27285 -18021 -26665 -16021
rect -19285 -18021 -18665 -16021
rect -11285 -18021 -10665 -16021
rect -3285 -18021 -2665 -16021
rect 4715 -18021 5335 -16021
rect 12715 -18021 13335 -16021
rect 20715 -18021 21335 -16021
rect 28715 -18021 29335 -16021
rect 36715 -18021 37335 -16021
rect 44715 -18021 45335 -16021
rect 54907 -18021 56907 -16021
rect -51093 -22021 -49093 -20021
rect -39285 -22021 -38665 -20021
rect -31285 -22021 -30665 -20021
rect -23285 -22021 -22665 -20021
rect -15285 -22021 -14665 -20021
rect -7285 -22021 -6665 -20021
rect 715 -22021 1335 -20021
rect 8715 -22021 9335 -20021
rect 16715 -22021 17335 -20021
rect 24715 -22021 25335 -20021
rect 32715 -22021 33335 -20021
rect 40715 -22021 41335 -20021
rect 48715 -22021 49335 -20021
rect 58907 -22021 60907 -20021
<< metal5 >>
rect -55093 88466 -53093 90442
rect -55117 88442 -53069 88466
rect -55117 86442 -55093 88442
rect -53093 86442 -53069 88442
rect -55117 86418 -53069 86442
rect -55093 -15997 -53093 86418
rect -51093 84466 -49093 90441
rect 54907 88466 56907 90441
rect -43309 88442 -42641 88466
rect -43309 86442 -43285 88442
rect -42665 86442 -42641 88442
rect -43309 86418 -42641 86442
rect -51117 84442 -49069 84466
rect -51117 82442 -51093 84442
rect -49093 82442 -49069 84442
rect -51117 82418 -49069 82442
rect -55117 -16021 -53069 -15997
rect -55117 -18021 -55093 -16021
rect -53093 -18021 -53069 -16021
rect -55117 -18045 -53069 -18021
rect -55093 -24021 -53093 -18045
rect -51093 -19997 -49093 82418
rect -43285 -15997 -42665 86418
rect -39285 84466 -38665 88466
rect -35309 88442 -34641 88466
rect -35309 86442 -35285 88442
rect -34665 86442 -34641 88442
rect -35309 86418 -34641 86442
rect -39309 84442 -38641 84466
rect -39309 82442 -39285 84442
rect -38665 82442 -38641 84442
rect -39309 82418 -38641 82442
rect -39285 23714 -38665 82418
rect -39285 23474 -39205 23714
rect -38742 23474 -38665 23714
rect -39285 16200 -38665 23474
rect -39285 15960 -39204 16200
rect -38741 15960 -38665 16200
rect -43309 -16021 -42641 -15997
rect -43309 -18021 -43285 -16021
rect -42665 -18021 -42641 -16021
rect -43309 -18045 -42641 -18021
rect -51117 -20021 -49069 -19997
rect -51117 -22021 -51093 -20021
rect -49093 -22021 -49069 -20021
rect -51117 -22045 -49069 -22021
rect -43285 -22045 -42665 -18045
rect -39285 -19997 -38665 15960
rect -35285 38498 -34665 86418
rect -31285 84466 -30665 88466
rect -27309 88442 -26641 88466
rect -27309 86442 -27285 88442
rect -26665 86442 -26641 88442
rect -27309 86418 -26641 86442
rect -31309 84442 -30641 84466
rect -31309 82442 -31285 84442
rect -30665 82442 -30641 84442
rect -31309 82418 -30641 82442
rect -35285 38258 -35218 38498
rect -34755 38258 -34665 38498
rect -35285 26908 -34665 38258
rect -35285 26668 -35224 26908
rect -34761 26668 -34665 26908
rect -35285 19233 -34665 26668
rect -35285 18993 -35218 19233
rect -34755 18993 -34665 19233
rect -35285 -15997 -34665 18993
rect -31285 38509 -30665 82418
rect -31285 38269 -31206 38509
rect -30743 38269 -30665 38509
rect -31285 37411 -30665 38269
rect -31285 37171 -31218 37411
rect -30755 37171 -30665 37411
rect -35309 -16021 -34641 -15997
rect -35309 -18021 -35285 -16021
rect -34665 -18021 -34641 -16021
rect -35309 -18045 -34641 -18021
rect -39309 -20021 -38641 -19997
rect -39309 -22021 -39285 -20021
rect -38665 -22021 -38641 -20021
rect -39309 -22045 -38641 -22021
rect -35285 -22045 -34665 -18045
rect -31285 -19997 -30665 37171
rect -27285 49826 -26665 86418
rect -23285 84466 -22665 88466
rect -19309 88442 -18641 88466
rect -19309 86442 -19285 88442
rect -18665 86442 -18641 88442
rect -19309 86418 -18641 86442
rect -23309 84442 -22641 84466
rect -23309 82442 -23285 84442
rect -22665 82442 -22641 84442
rect -23309 82418 -22641 82442
rect -27285 49586 -27236 49826
rect -26706 49586 -26665 49826
rect -27285 43156 -26665 49586
rect -27285 42916 -27162 43156
rect -26709 42916 -26665 43156
rect -27285 39950 -26665 42916
rect -27285 39710 -27162 39950
rect -26699 39710 -26665 39950
rect -27285 35881 -26665 39710
rect -27285 35641 -27162 35881
rect -26699 35641 -26665 35881
rect -27285 32767 -26665 35641
rect -27285 32527 -27162 32767
rect -26704 32527 -26665 32767
rect -27285 25514 -26665 32527
rect -27285 25274 -27228 25514
rect -26698 25274 -26665 25514
rect -27285 17963 -26665 25274
rect -27285 17723 -27238 17963
rect -26708 17723 -26665 17963
rect -27285 14477 -26665 17723
rect -27285 14237 -27231 14477
rect -26701 14237 -26665 14477
rect -27285 6710 -26665 14237
rect -27285 6470 -27239 6710
rect -26709 6470 -26665 6710
rect -27285 -15997 -26665 6470
rect -23285 49223 -22665 82418
rect -23285 48983 -23234 49223
rect -22704 48983 -22665 49223
rect -23285 38013 -22665 48983
rect -23285 37540 -23192 38013
rect -22729 37540 -22665 38013
rect -23285 24917 -22665 37540
rect -23285 24677 -23236 24917
rect -22706 24677 -22665 24917
rect -23285 15490 -22665 24677
rect -23285 15250 -23253 15490
rect -22723 15250 -22665 15490
rect -23285 5044 -22665 15250
rect -23285 4804 -23232 5044
rect -22702 4804 -22665 5044
rect -27309 -16021 -26641 -15997
rect -27309 -18021 -27285 -16021
rect -26665 -18021 -26641 -16021
rect -27309 -18045 -26641 -18021
rect -31309 -20021 -30641 -19997
rect -31309 -22021 -31285 -20021
rect -30665 -22021 -30641 -20021
rect -31309 -22045 -30641 -22021
rect -27285 -22045 -26665 -18045
rect -23285 -19997 -22665 4804
rect -19285 75068 -18665 86418
rect -15285 84466 -14665 88466
rect -11309 88442 -10641 88466
rect -11309 86442 -11285 88442
rect -10665 86442 -10641 88442
rect -11309 86418 -10641 86442
rect -15309 84442 -14641 84466
rect -15309 82442 -15285 84442
rect -14665 82442 -14641 84442
rect -15309 82418 -14641 82442
rect -19285 74828 -19241 75068
rect -18711 74828 -18665 75068
rect -19285 70237 -18665 74828
rect -19285 69997 -19241 70237
rect -18711 69997 -18665 70237
rect -19285 67122 -18665 69997
rect -19285 66882 -19245 67122
rect -18715 66882 -18665 67122
rect -19285 50690 -18665 66882
rect -19285 50450 -19238 50690
rect -18708 50450 -18665 50690
rect -19285 28708 -18665 50450
rect -19285 28468 -19238 28708
rect -18708 28468 -18665 28708
rect -19285 25810 -18665 28468
rect -19285 25570 -19246 25810
rect -18716 25570 -18665 25810
rect -19285 23730 -18665 25570
rect -19285 23490 -19239 23730
rect -18709 23490 -18665 23730
rect -19285 -15997 -18665 23490
rect -15285 75253 -14665 82418
rect -15285 75013 -15243 75253
rect -14713 75013 -14665 75253
rect -15285 70994 -14665 75013
rect -15285 70754 -15242 70994
rect -14712 70754 -14665 70994
rect -15285 68915 -14665 70754
rect -15285 68675 -15239 68915
rect -14709 68675 -14665 68915
rect -15285 27443 -14665 68675
rect -15285 27203 -15234 27443
rect -14704 27203 -14665 27443
rect -15285 25818 -14665 27203
rect -15285 25578 -15238 25818
rect -14708 25578 -14665 25818
rect -15285 23639 -14665 25578
rect -15285 23399 -15237 23639
rect -14707 23399 -14665 23639
rect -19309 -16021 -18641 -15997
rect -19309 -18021 -19285 -16021
rect -18665 -18021 -18641 -16021
rect -19309 -18045 -18641 -18021
rect -23309 -20021 -22641 -19997
rect -23309 -22021 -23285 -20021
rect -22665 -22021 -22641 -20021
rect -23309 -22045 -22641 -22021
rect -19285 -22045 -18665 -18045
rect -15285 -19997 -14665 23399
rect -11285 63557 -10665 86418
rect -7285 84466 -6665 88466
rect -3309 88442 -2641 88466
rect -3309 86442 -3285 88442
rect -2665 86442 -2641 88442
rect -3309 86418 -2641 86442
rect -7309 84442 -6641 84466
rect -7309 82442 -7285 84442
rect -6665 82442 -6641 84442
rect -7309 82418 -6641 82442
rect -11285 63205 -11071 63557
rect -10737 63205 -10665 63557
rect -11285 28055 -10665 63205
rect -11285 27815 -11237 28055
rect -10707 27815 -10665 28055
rect -11285 23154 -10665 27815
rect -11285 22914 -11246 23154
rect -10716 22914 -10665 23154
rect -11285 -15997 -10665 22914
rect -7285 63206 -6665 82418
rect -7285 62966 -6939 63206
rect -6699 62966 -6665 63206
rect -7285 55397 -6665 62966
rect -7285 54706 -6978 55397
rect -6706 54706 -6665 55397
rect -7285 51701 -6665 54706
rect -7285 51461 -7237 51701
rect -6707 51461 -6665 51701
rect -7285 15812 -6665 51461
rect -7285 15572 -7218 15812
rect -6755 15572 -6665 15812
rect -7285 14452 -6665 15572
rect -7285 14212 -7221 14452
rect -6758 14212 -6665 14452
rect -7285 10912 -6665 14212
rect -7285 10672 -7221 10912
rect -6758 10672 -6665 10912
rect -7285 9662 -6665 10672
rect -7285 9422 -7211 9662
rect -6748 9422 -6665 9662
rect -7285 7243 -6665 9422
rect -7285 7003 -7214 7243
rect -6751 7003 -6665 7243
rect -7285 5764 -6665 7003
rect -7285 5524 -7211 5764
rect -6748 5524 -6665 5764
rect -7285 -8276 -6665 5524
rect -7285 -8516 -7204 -8276
rect -6741 -8516 -6665 -8276
rect -11309 -16021 -10641 -15997
rect -11309 -18021 -11285 -16021
rect -10665 -18021 -10641 -16021
rect -11309 -18045 -10641 -18021
rect -15309 -20021 -14641 -19997
rect -15309 -22021 -15285 -20021
rect -14665 -22021 -14641 -20021
rect -15309 -22045 -14641 -22021
rect -11285 -22045 -10665 -18045
rect -7285 -19997 -6665 -8516
rect -3285 63411 -2665 86418
rect 715 84466 1335 88466
rect 4691 88442 5359 88466
rect 4691 86442 4715 88442
rect 5335 86442 5359 88442
rect 4691 86418 5359 86442
rect 691 84442 1359 84466
rect 691 82442 715 84442
rect 1335 82442 1359 84442
rect 691 82418 1359 82442
rect -3285 63171 -3241 63411
rect -2711 63171 -2665 63411
rect -3285 54422 -2665 63171
rect -3285 54182 -3237 54422
rect -2707 54182 -2665 54422
rect -3285 51101 -2665 54182
rect -3285 50861 -3231 51101
rect -2701 50861 -2665 51101
rect -3285 48773 -2665 50861
rect -3285 48533 -3237 48773
rect -2707 48533 -2665 48773
rect -3285 45355 -2665 48533
rect -3285 45115 -3248 45355
rect -2718 45115 -2665 45355
rect -3285 39886 -2665 45115
rect -3285 39646 -3233 39886
rect -2703 39646 -2665 39886
rect -3285 17864 -2665 39646
rect -3285 17624 -3211 17864
rect -2748 17624 -2665 17864
rect -3285 16450 -2665 17624
rect -3285 16210 -3201 16450
rect -2738 16210 -2665 16450
rect -3285 14048 -2665 16210
rect -3285 13808 -3199 14048
rect -2736 13808 -2665 14048
rect -3285 8802 -2665 13808
rect -3285 8562 -3201 8802
rect -2738 8562 -2665 8802
rect -3285 6743 -2665 8562
rect -3285 6503 -3199 6743
rect -2736 6503 -2665 6743
rect -3285 -6173 -2665 6503
rect -3285 -6413 -3198 -6173
rect -2735 -6413 -2665 -6173
rect -3285 -15997 -2665 -6413
rect 715 63232 1335 82418
rect 715 62992 757 63232
rect 1287 62992 1335 63232
rect 715 60124 1335 62992
rect 715 59884 756 60124
rect 1286 59884 1335 60124
rect 715 56749 1335 59884
rect 715 56509 756 56749
rect 1286 56509 1335 56749
rect 715 53374 1335 56509
rect 715 53134 756 53374
rect 1286 53134 1335 53374
rect 715 49999 1335 53134
rect 715 49759 756 49999
rect 1286 49759 1335 49999
rect 715 44514 1335 49759
rect 715 44274 752 44514
rect 1282 44274 1335 44514
rect 715 40869 1335 44274
rect 715 40629 762 40869
rect 1292 40629 1335 40869
rect 715 39440 1335 40629
rect 715 39200 756 39440
rect 1286 39200 1335 39440
rect 715 37095 1335 39200
rect 715 36855 757 37095
rect 1287 36855 1335 37095
rect 715 36016 1335 36855
rect 715 35776 774 36016
rect 1304 35776 1335 36016
rect 715 17618 1335 35776
rect 715 17378 789 17618
rect 1252 17378 1335 17618
rect 715 10149 1335 17378
rect 715 9909 792 10149
rect 1255 9909 1335 10149
rect 715 7960 1335 9909
rect 715 7720 805 7960
rect 1268 7720 1335 7960
rect 715 2273 1335 7720
rect 715 2033 778 2273
rect 1241 2033 1335 2273
rect 715 325 1335 2033
rect 715 85 794 325
rect 1257 85 1335 325
rect -3309 -16021 -2641 -15997
rect -3309 -18021 -3285 -16021
rect -2665 -18021 -2641 -16021
rect -3309 -18045 -2641 -18021
rect -7309 -20021 -6641 -19997
rect -7309 -22021 -7285 -20021
rect -6665 -22021 -6641 -20021
rect -7309 -22045 -6641 -22021
rect -3285 -22045 -2665 -18045
rect 715 -19997 1335 85
rect 4715 38053 5335 86418
rect 8715 84466 9335 88466
rect 12691 88442 13359 88466
rect 12691 86442 12715 88442
rect 13335 86442 13359 88442
rect 12691 86418 13359 86442
rect 8691 84442 9359 84466
rect 8691 82442 8715 84442
rect 9335 82442 9359 84442
rect 8691 82418 9359 82442
rect 4715 37813 4761 38053
rect 5291 37813 5335 38053
rect 4715 36660 5335 37813
rect 4715 36420 4768 36660
rect 5298 36420 5335 36660
rect 4715 35482 5335 36420
rect 4715 35242 4774 35482
rect 5304 35242 5335 35482
rect 4715 23159 5335 35242
rect 4715 22919 4780 23159
rect 5243 22919 5335 23159
rect 4715 19233 5335 22919
rect 4715 18993 4797 19233
rect 5260 18993 5335 19233
rect 4715 16746 5335 18993
rect 4715 16430 4794 16746
rect 4715 16190 4792 16430
rect 4715 15884 4794 16190
rect 5256 15884 5335 16746
rect 4715 14621 5335 15884
rect 4715 14381 4794 14621
rect 5257 14381 5335 14621
rect 4715 12013 5335 14381
rect 4715 11773 4783 12013
rect 5246 11773 5335 12013
rect 4715 -15997 5335 11773
rect 8715 60113 9335 82418
rect 8715 59873 8761 60113
rect 9291 59873 9335 60113
rect 8715 56738 9335 59873
rect 8715 56498 8760 56738
rect 9290 56498 9335 56738
rect 8715 53363 9335 56498
rect 8715 53123 8760 53363
rect 9290 53123 9335 53363
rect 8715 49988 9335 53123
rect 8715 49748 8760 49988
rect 9290 49748 9335 49988
rect 8715 43238 9335 49748
rect 8715 42998 8760 43238
rect 9290 42998 9335 43238
rect 8715 36028 9335 42998
rect 8715 35788 8758 36028
rect 9288 35788 9335 36028
rect 8715 23495 9335 35788
rect 8715 23255 8774 23495
rect 9237 23255 9335 23495
rect 8715 17403 9335 23255
rect 8715 17163 8789 17403
rect 9252 17163 9335 17403
rect 8715 10124 9335 17163
rect 8715 9884 8768 10124
rect 9231 9884 9335 10124
rect 8715 337 9335 9884
rect 8715 97 8814 337
rect 9277 97 9335 337
rect 4691 -16021 5359 -15997
rect 4691 -18021 4715 -16021
rect 5335 -18021 5359 -16021
rect 4691 -18045 5359 -18021
rect 691 -20021 1359 -19997
rect 691 -22021 715 -20021
rect 1335 -22021 1359 -20021
rect 691 -22045 1359 -22021
rect 4715 -22045 5335 -18045
rect 8715 -19997 9335 97
rect 12715 75172 13335 86418
rect 16715 84466 17335 88466
rect 20691 88442 21359 88466
rect 20691 86442 20715 88442
rect 21335 86442 21359 88442
rect 20691 86418 21359 86442
rect 16691 84442 17359 84466
rect 16691 82442 16715 84442
rect 17335 82442 17359 84442
rect 16691 82418 17359 82442
rect 12715 74932 12758 75172
rect 13288 74932 13335 75172
rect 12715 21097 13335 74932
rect 12715 20855 12861 21097
rect 13103 20855 13335 21097
rect 12715 18796 13335 20855
rect 12715 18554 12849 18796
rect 13091 18554 13335 18796
rect 12715 17191 13335 18554
rect 12715 16949 12843 17191
rect 13085 16949 13335 17191
rect 12715 15320 13335 16949
rect 12715 15078 12862 15320
rect 13104 15078 13335 15320
rect 12715 13619 13335 15078
rect 12715 13377 12884 13619
rect 13126 13377 13335 13619
rect 12715 11764 13335 13377
rect 12715 11522 12897 11764
rect 13139 11522 13335 11764
rect 12715 10653 13335 11522
rect 12715 10413 12783 10653
rect 13246 10413 13335 10653
rect 12715 -15997 13335 10413
rect 16715 75164 17335 82418
rect 16715 74924 16757 75164
rect 17287 74924 17335 75164
rect 16715 62728 17335 74924
rect 16715 62200 16766 62728
rect 17291 62200 17335 62728
rect 16715 58728 17335 62200
rect 16715 58200 16766 58728
rect 17291 58200 17335 58728
rect 16715 54728 17335 58200
rect 16715 54200 16766 54728
rect 17291 54200 17335 54728
rect 16715 50728 17335 54200
rect 16715 50200 16766 50728
rect 17291 50200 17335 50728
rect 16715 46728 17335 50200
rect 16715 46200 16766 46728
rect 17291 46200 17335 46728
rect 16715 19188 17335 46200
rect 16715 18946 16889 19188
rect 17131 18946 17335 19188
rect 16715 15595 17335 18946
rect 16715 15353 16797 15595
rect 17039 15353 17335 15595
rect 16715 10139 17335 15353
rect 16715 9899 16808 10139
rect 17271 9899 17335 10139
rect 16715 325 17335 9899
rect 16715 85 16791 325
rect 17254 85 17335 325
rect 12691 -16021 13359 -15997
rect 12691 -18021 12715 -16021
rect 13335 -18021 13359 -16021
rect 12691 -18045 13359 -18021
rect 8691 -20021 9359 -19997
rect 8691 -22021 8715 -20021
rect 9335 -22021 9359 -20021
rect 8691 -22045 9359 -22021
rect 12715 -22045 13335 -18045
rect 16715 -19997 17335 85
rect 20715 64719 21335 86418
rect 24715 84466 25335 88466
rect 28691 88442 29359 88466
rect 28691 86442 28715 88442
rect 29335 86442 29359 88442
rect 28691 86418 29359 86442
rect 24691 84442 25359 84466
rect 24691 82442 24715 84442
rect 25335 82442 25359 84442
rect 24691 82418 25359 82442
rect 20715 64191 20763 64719
rect 21288 64191 21335 64719
rect 20715 60719 21335 64191
rect 20715 60191 20763 60719
rect 21288 60191 21335 60719
rect 20715 56719 21335 60191
rect 20715 56191 20763 56719
rect 21288 56191 21335 56719
rect 20715 52719 21335 56191
rect 20715 52191 20763 52719
rect 21288 52191 21335 52719
rect 20715 48719 21335 52191
rect 20715 48191 20763 48719
rect 21288 48191 21335 48719
rect 20715 19161 21335 48191
rect 20715 18919 20893 19161
rect 21135 18919 21335 19161
rect 20715 15590 21335 18919
rect 20715 15348 20836 15590
rect 21078 15348 21335 15590
rect 20715 12002 21335 15348
rect 20715 11760 20890 12002
rect 21132 11760 21335 12002
rect 20715 -15997 21335 11760
rect 24715 62721 25335 82418
rect 24715 62193 24762 62721
rect 25287 62193 25335 62721
rect 24715 58721 25335 62193
rect 24715 58193 24762 58721
rect 25287 58193 25335 58721
rect 24715 54721 25335 58193
rect 24715 54193 24762 54721
rect 25287 54193 25335 54721
rect 24715 50721 25335 54193
rect 24715 50193 24762 50721
rect 25287 50193 25335 50721
rect 24715 46721 25335 50193
rect 24715 46193 24762 46721
rect 25287 46193 25335 46721
rect 24715 19156 25335 46193
rect 24715 18914 24903 19156
rect 25145 18914 25335 19156
rect 24715 15563 25335 18914
rect 24715 15321 24905 15563
rect 25147 15321 25335 15563
rect 24715 11972 25335 15321
rect 24715 11730 24893 11972
rect 25135 11730 25335 11972
rect 24715 5982 25335 11730
rect 24715 5410 24797 5982
rect 25260 5410 25335 5982
rect 24715 1606 25335 5410
rect 24715 1366 24796 1606
rect 25259 1366 25335 1606
rect 20691 -16021 21359 -15997
rect 20691 -18021 20715 -16021
rect 21335 -18021 21359 -16021
rect 20691 -18045 21359 -18021
rect 16691 -20021 17359 -19997
rect 16691 -22021 16715 -20021
rect 17335 -22021 17359 -20021
rect 16691 -22045 17359 -22021
rect 20715 -22045 21335 -18045
rect 24715 -19997 25335 1366
rect 28715 64725 29335 86418
rect 32715 84466 33335 88466
rect 36691 88442 37359 88466
rect 36691 86442 36715 88442
rect 37335 86442 37359 88442
rect 36691 86418 37359 86442
rect 32691 84442 33359 84466
rect 32691 82442 32715 84442
rect 33335 82442 33359 84442
rect 32691 82418 33359 82442
rect 28715 64197 28757 64725
rect 29282 64197 29335 64725
rect 28715 60725 29335 64197
rect 28715 60197 28757 60725
rect 29282 60197 29335 60725
rect 28715 56725 29335 60197
rect 28715 56197 28757 56725
rect 29282 56197 29335 56725
rect 28715 52725 29335 56197
rect 28715 52197 28757 52725
rect 29282 52197 29335 52725
rect 28715 48725 29335 52197
rect 28715 48197 28757 48725
rect 29282 48197 29335 48725
rect 28715 -15997 29335 48197
rect 32715 62717 33335 82418
rect 32715 62189 32765 62717
rect 33290 62189 33335 62717
rect 32715 58717 33335 62189
rect 32715 58189 32765 58717
rect 33290 58189 33335 58717
rect 32715 54717 33335 58189
rect 32715 54189 32765 54717
rect 33290 54189 33335 54717
rect 32715 50717 33335 54189
rect 32715 50189 32765 50717
rect 33290 50189 33335 50717
rect 32715 46717 33335 50189
rect 32715 46189 32765 46717
rect 33290 46189 33335 46717
rect 32715 24134 33335 46189
rect 32715 23894 32791 24134
rect 33254 23894 33335 24134
rect 32715 21674 33335 23894
rect 32715 21434 32790 21674
rect 33253 21434 33335 21674
rect 32715 7293 33335 21434
rect 32715 7053 32793 7293
rect 33256 7053 33335 7293
rect 32715 5993 33335 7053
rect 32715 5753 32784 5993
rect 33247 5753 33335 5993
rect 32715 4578 33335 5753
rect 32715 4338 32790 4578
rect 33253 4338 33335 4578
rect 32715 3205 33335 4338
rect 32715 2965 32786 3205
rect 33249 2965 33335 3205
rect 32715 353 33335 2965
rect 32715 113 32793 353
rect 33256 113 33335 353
rect 32715 -947 33335 113
rect 32715 -1187 32784 -947
rect 33247 -1187 33335 -947
rect 32715 -2362 33335 -1187
rect 32715 -2602 32790 -2362
rect 33253 -2602 33335 -2362
rect 32715 -3735 33335 -2602
rect 32715 -3975 32786 -3735
rect 33249 -3975 33335 -3735
rect 28691 -16021 29359 -15997
rect 28691 -18021 28715 -16021
rect 29335 -18021 29359 -16021
rect 28691 -18045 29359 -18021
rect 24691 -20021 25359 -19997
rect 24691 -22021 24715 -20021
rect 25335 -22021 25359 -20021
rect 24691 -22045 25359 -22021
rect 28715 -22045 29335 -18045
rect 32715 -19997 33335 -3975
rect 36715 22815 37335 86418
rect 40715 84466 41335 88466
rect 44691 88442 45359 88466
rect 44691 86442 44715 88442
rect 45335 86442 45359 88442
rect 44691 86418 45359 86442
rect 40691 84442 41359 84466
rect 40691 82442 40715 84442
rect 41335 82442 41359 84442
rect 40691 82418 41359 82442
rect 36715 22579 36914 22815
rect 37156 22579 37335 22815
rect 36715 8810 37335 22579
rect 36715 8537 36881 8810
rect 37155 8537 37335 8810
rect 36715 6525 37335 8537
rect 36715 6289 36938 6525
rect 37180 6289 37335 6525
rect 36715 5109 37335 6289
rect 36715 4873 36899 5109
rect 37141 4873 37335 5109
rect 36715 2832 37335 4873
rect 36715 2559 36889 2832
rect 37163 2559 37335 2832
rect 36715 1870 37335 2559
rect 36715 1597 36881 1870
rect 37155 1597 37335 1870
rect 36715 -415 37335 1597
rect 36715 -651 36938 -415
rect 37180 -651 37335 -415
rect 36715 -1831 37335 -651
rect 36715 -2067 36899 -1831
rect 37141 -2067 37335 -1831
rect 36715 -4108 37335 -2067
rect 36715 -4381 36889 -4108
rect 37163 -4381 37335 -4108
rect 36715 -15997 37335 -4381
rect 40715 44304 41335 82418
rect 40715 44064 40800 44304
rect 41263 44064 41335 44304
rect 40715 40559 41335 44064
rect 40715 40319 40808 40559
rect 41271 40319 41335 40559
rect 40715 22732 41335 40319
rect 40715 22492 40801 22732
rect 41264 22492 41335 22732
rect 40715 7170 41335 22492
rect 40715 6930 40801 7170
rect 41264 6930 41335 7170
rect 40715 4267 41335 6930
rect 40715 4027 40799 4267
rect 41262 4027 41335 4267
rect 40715 230 41335 4027
rect 40715 -10 40801 230
rect 41264 -10 41335 230
rect 40715 -2673 41335 -10
rect 40715 -2680 40799 -2673
rect 40715 -2920 40785 -2680
rect 41262 -2913 41335 -2673
rect 41248 -2920 41335 -2913
rect 36691 -16021 37359 -15997
rect 36691 -18021 36715 -16021
rect 37335 -18021 37359 -16021
rect 36691 -18045 37359 -18021
rect 32691 -20021 33359 -19997
rect 32691 -22021 32715 -20021
rect 33335 -22021 33359 -20021
rect 32691 -22045 33359 -22021
rect 36715 -22045 37335 -18045
rect 40715 -19997 41335 -2920
rect 44715 45174 45335 86418
rect 48715 84466 49335 88466
rect 54883 88442 56931 88466
rect 54883 86442 54907 88442
rect 56907 86442 56931 88442
rect 54883 86418 56931 86442
rect 48691 84442 49359 84466
rect 48691 82442 48715 84442
rect 49335 82442 49359 84442
rect 48691 82418 49359 82442
rect 44715 44934 44795 45174
rect 45258 44934 45335 45174
rect 44715 44013 45335 44934
rect 44715 43773 44795 44013
rect 45258 43773 45335 44013
rect 44715 41504 45335 43773
rect 44715 41264 44779 41504
rect 45242 41264 45335 41504
rect 44715 40193 45335 41264
rect 44715 39953 44772 40193
rect 45235 39953 45335 40193
rect 44715 24252 45335 39953
rect 44715 24012 44801 24252
rect 45264 24012 45335 24252
rect 44715 7446 45335 24012
rect 44715 7206 44796 7446
rect 45259 7206 45335 7446
rect 44715 521 45335 7206
rect 44715 281 44799 521
rect 45262 281 45335 521
rect 44715 -15997 45335 281
rect 48715 21245 49335 82418
rect 48715 21005 48791 21245
rect 49254 21005 49335 21245
rect 44691 -16021 45359 -15997
rect 44691 -18021 44715 -16021
rect 45335 -18021 45359 -16021
rect 44691 -18045 45359 -18021
rect 40691 -20021 41359 -19997
rect 40691 -22021 40715 -20021
rect 41335 -22021 41359 -20021
rect 40691 -22045 41359 -22021
rect 44715 -22045 45335 -18045
rect 48715 -19997 49335 21005
rect 54907 -15997 56907 86418
rect 58907 84466 60907 90441
rect 58883 84442 60931 84466
rect 58883 82442 58907 84442
rect 60907 82442 60931 84442
rect 58883 82418 60931 82442
rect 54883 -16021 56931 -15997
rect 54883 -18021 54907 -16021
rect 56907 -18021 56931 -16021
rect 54883 -18045 56931 -18021
rect 48691 -20021 49359 -19997
rect 48691 -22021 48715 -20021
rect 49335 -22021 49359 -20021
rect 48691 -22045 49359 -22021
rect -51093 -24021 -49093 -22045
rect 54907 -24021 56907 -18045
rect 58907 -19997 60907 82418
rect 58883 -20021 60931 -19997
rect 58883 -22021 58907 -20021
rect 60907 -22021 60931 -20021
rect 58883 -22045 60931 -22021
rect 58907 -24021 60907 -22045
use a_mux2_en  a_mux2_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/a_mux2_en
timestamp 1654408082
transform 1 0 36330 0 1 23897
box -2638 -2585 3429 115
use a_mux2_en  a_mux2_en_1
timestamp 1654408082
transform 0 -1 -16584 1 0 68726
box -2638 -2585 3429 115
use a_mux4_en  a_mux4_en_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/a_mux4_en
timestamp 1654408082
transform 1 0 37083 0 1 1386
box -3690 -5314 3456 148
use a_mux4_en  a_mux4_en_1
timestamp 1654408082
transform 1 0 37083 0 1 8326
box -3690 -5314 3456 148
use clock_v2  clock_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/clock_v2
timestamp 1654408082
transform 0 1 31620 -1 0 62637
box -3193 -14204 16946 36
use comparator_v2  comparator_v2_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/comparator_v2
timestamp 1654408082
transform 0 -1 -18981 -1 0 39564
box -3788 -193 7250 10729
use esd_cell  esd_cell_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/esd_cell
timestamp 1654408082
transform 1 0 -38260 0 1 16027
box -65 -65 3553 3095
use esd_cell  esd_cell_1
timestamp 1654408082
transform 1 0 -38260 0 1 23557
box -65 -65 3553 3095
use esd_cell  esd_cell_2
timestamp 1654408082
transform 0 -1 14206 1 0 73319
box -65 -65 3553 3095
use esd_cell  esd_cell_3
timestamp 1654408082
transform 0 1 -3548 -1 0 -6736
box -65 -65 3553 3095
use esd_cell  esd_cell_4
timestamp 1654408082
transform 0 -1 -13798 1 0 73319
box -65 -65 3553 3095
use esd_cell  esd_cell_5
timestamp 1654408082
transform 1 0 42777 0 1 21122
box -65 -65 3553 3095
use esd_cell  esd_cell_6
timestamp 1654408082
transform 1 0 42522 0 1 -2751
box -65 -65 3553 3095
use esd_cell  esd_cell_7
timestamp 1654408082
transform 1 0 42522 0 1 4189
box -65 -65 3553 3095
use onebit_dac  onebit_dac_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/onebit_dac
timestamp 1654408082
transform 1 0 -17091 0 1 24436
box -313 -1154 1895 1114
use onebit_dac  onebit_dac_1
timestamp 1654408082
transform 1 0 -17086 0 1 27078
box -313 -1154 1895 1114
use ota  ota_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/ota
timestamp 1654408082
transform 1 0 7664 0 1 17642
box -7664 -17642 18422 2891
use ota  ota_1
timestamp 1654408082
transform 0 -1 -7144 1 0 47315
box -7664 -17642 18422 2891
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_0
timestamp 1654408082
transform 0 1 9865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_1
timestamp 1654408082
transform 0 1 9865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_2
timestamp 1654408082
transform 0 1 9865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_3
timestamp 1654408082
transform 0 1 9865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_4
timestamp 1654408082
transform 0 1 9865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_5
timestamp 1654408082
transform 0 1 9865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_6
timestamp 1654408082
transform 0 1 9865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_7
timestamp 1654408082
transform 0 1 9865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_8
timestamp 1654408082
transform 0 1 8865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_9
timestamp 1654408082
transform 0 1 8865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_10
timestamp 1654408082
transform 0 1 8865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_11
timestamp 1654408082
transform 0 1 8865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_12
timestamp 1654408082
transform 0 1 8865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_13
timestamp 1654408082
transform 0 1 8865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_14
timestamp 1654408082
transform 0 1 8865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_15
timestamp 1654408082
transform 0 1 8865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_16
timestamp 1654408082
transform 0 1 8865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_17
timestamp 1654408082
transform 0 1 7865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_18
timestamp 1654408082
transform 0 1 7865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_19
timestamp 1654408082
transform 0 1 7865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_20
timestamp 1654408082
transform 0 1 7865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_21
timestamp 1654408082
transform 0 1 7865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_22
timestamp 1654408082
transform 0 1 7865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_23
timestamp 1654408082
transform 0 1 7865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_24
timestamp 1654408082
transform 0 1 7865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_25
timestamp 1654408082
transform 0 1 7865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_26
timestamp 1654408082
transform 0 1 6865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_27
timestamp 1654408082
transform 0 1 6865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_28
timestamp 1654408082
transform 0 1 6865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_29
timestamp 1654408082
transform 0 1 6865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_30
timestamp 1654408082
transform 0 1 6865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_31
timestamp 1654408082
transform 0 1 6865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_32
timestamp 1654408082
transform 0 1 6865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_33
timestamp 1654408082
transform 0 1 6865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_34
timestamp 1654408082
transform 0 1 6865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_35
timestamp 1654408082
transform 0 -1 3865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_36
timestamp 1654408082
transform 0 -1 3865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_37
timestamp 1654408082
transform 0 -1 2865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_38
timestamp 1654408082
transform 0 -1 2865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_39
timestamp 1654408082
transform 0 -1 3865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_40
timestamp 1654408082
transform 0 -1 3865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_41
timestamp 1654408082
transform 0 -1 2865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_42
timestamp 1654408082
transform 0 -1 2865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_43
timestamp 1654408082
transform 0 -1 3865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_44
timestamp 1654408082
transform 0 -1 3865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_45
timestamp 1654408082
transform 0 -1 2865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_46
timestamp 1654408082
transform 0 -1 2865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_47
timestamp 1654408082
transform 0 -1 3865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_48
timestamp 1654408082
transform 0 -1 3865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_49
timestamp 1654408082
transform 0 -1 2865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_50
timestamp 1654408082
transform 0 -1 2865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_51
timestamp 1654408082
transform 0 -1 3865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_52
timestamp 1654408082
transform 0 -1 2865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_53
timestamp 1654408082
transform 0 -1 5865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_54
timestamp 1654408082
transform 0 -1 4865 -1 0 26238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_55
timestamp 1654408082
transform 0 -1 5865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_56
timestamp 1654408082
transform 0 -1 4865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_57
timestamp 1654408082
transform 0 -1 5865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_58
timestamp 1654408082
transform 0 -1 4865 -1 0 28238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_59
timestamp 1654408082
transform 0 -1 5865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_60
timestamp 1654408082
transform 0 -1 4865 -1 0 27238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_61
timestamp 1654408082
transform 0 -1 5865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_62
timestamp 1654408082
transform 0 -1 5865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_63
timestamp 1654408082
transform 0 -1 4865 -1 0 30238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_64
timestamp 1654408082
transform 0 -1 4865 -1 0 29238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_65
timestamp 1654408082
transform 0 -1 5865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_66
timestamp 1654408082
transform 0 -1 5865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_67
timestamp 1654408082
transform 0 -1 4865 -1 0 32238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_68
timestamp 1654408082
transform 0 -1 4865 -1 0 31238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_69
timestamp 1654408082
transform 0 -1 5865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_70
timestamp 1654408082
transform 0 1 9865 -1 0 25238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_71
timestamp 1654408082
transform 0 -1 4865 -1 0 33238
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_0
timestamp 1654408082
transform 1 0 -9068 0 1 19276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_1
timestamp 1654408082
transform 1 0 -9068 0 1 16676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_2
timestamp 1654408082
transform 1 0 -9068 0 1 14076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_3
timestamp 1654408082
transform 1 0 -9068 0 1 11476
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_4
timestamp 1654408082
transform 1 0 -9068 0 1 8876
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_5
timestamp 1654408082
transform 1 0 -19468 0 1 3676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_6
timestamp 1654408082
transform 1 0 -11668 0 1 11476
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_7
timestamp 1654408082
transform 1 0 -11668 0 1 14076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_8
timestamp 1654408082
transform 1 0 -11668 0 1 16676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_9
timestamp 1654408082
transform 1 0 -11668 0 1 19276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_10
timestamp 1654408082
transform 1 0 -16868 0 1 3676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_11
timestamp 1654408082
transform 1 0 -14268 0 1 11476
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_12
timestamp 1654408082
transform 1 0 -14268 0 1 14076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_13
timestamp 1654408082
transform 1 0 -14268 0 1 16676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_14
timestamp 1654408082
transform 1 0 -14268 0 1 19276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_15
timestamp 1654408082
transform 1 0 -11668 0 1 3676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_16
timestamp 1654408082
transform 1 0 -16868 0 1 11476
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_17
timestamp 1654408082
transform 1 0 -16868 0 1 14076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_18
timestamp 1654408082
transform 1 0 -16868 0 1 16676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_19
timestamp 1654408082
transform 1 0 -16868 0 1 19276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_20
timestamp 1654408082
transform 1 0 -14268 0 1 3676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_21
timestamp 1654408082
transform 1 0 -19468 0 1 11476
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_22
timestamp 1654408082
transform 1 0 -19468 0 1 14076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_23
timestamp 1654408082
transform 1 0 -19468 0 1 16676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_24
timestamp 1654408082
transform 1 0 -19468 0 1 19276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_25
timestamp 1654408082
transform 1 0 -22068 0 1 8876
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_26
timestamp 1654408082
transform 1 0 -22068 0 1 11476
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_27
timestamp 1654408082
transform 1 0 -22068 0 1 14076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_28
timestamp 1654408082
transform 1 0 -22068 0 1 16676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_29
timestamp 1654408082
transform 1 0 -22068 0 1 19276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_30
timestamp 1654408082
transform 1 0 -16868 0 1 8876
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_31
timestamp 1654408082
transform 1 0 -19468 0 1 8876
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_32
timestamp 1654408082
transform 1 0 -16868 0 1 6276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_33
timestamp 1654408082
transform 1 0 -19468 0 1 6276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_34
timestamp 1654408082
transform 1 0 -11668 0 1 8876
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_35
timestamp 1654408082
transform 1 0 -14268 0 1 8876
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_36
timestamp 1654408082
transform 1 0 -11668 0 1 6276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_37
timestamp 1654408082
transform 1 0 -14268 0 1 6276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_38
timestamp 1654408082
transform 1 0 -22068 0 1 6276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_39
timestamp 1654408082
transform 1 0 -9068 0 1 6276
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_40
timestamp 1654408082
transform 1 0 -22068 0 1 3676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_41
timestamp 1654408082
transform 1 0 -9068 0 1 3676
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_42
timestamp 1654408082
transform 1 0 -22068 0 1 1076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_43
timestamp 1654408082
transform 1 0 -9068 0 1 1076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_44
timestamp 1654408082
transform 1 0 -19468 0 1 1076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_45
timestamp 1654408082
transform 1 0 -16868 0 1 1076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_46
timestamp 1654408082
transform 1 0 -14268 0 1 1076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_47
timestamp 1654408082
transform 1 0 -11668 0 1 1076
box -1030 -980 976 980
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_0
timestamp 1654408082
transform 1 0 -15946 0 -1 36367
box -1310 -1260 1210 1260
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_1
timestamp 1654408082
transform 1 0 -15946 0 -1 39777
box -1310 -1260 1210 1260
use sky130_fd_pr__nfet_01v8_CFEPS5  sky130_fd_pr__nfet_01v8_CFEPS5_0
timestamp 1654408082
transform 1 0 -31520 0 -1 38989
box -311 -274 311 274
use sky130_fd_pr__pfet_01v8_XAYTAL  sky130_fd_pr__pfet_01v8_XAYTAL_0
timestamp 1654408082
transform 1 0 -31520 0 -1 38389
box -311 -319 311 319
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654408082
transform 1 0 -26628 0 1 49146
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1654408082
transform 1 0 42422 0 1 39535
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_2
timestamp 1654408082
transform 1 0 42422 0 1 40805
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_3
timestamp 1654408082
transform 1 0 42422 0 1 43345
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_4
timestamp 1654408082
transform 1 0 42422 0 1 44495
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654408082
transform 1 0 43158 0 1 39535
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1654408082
transform 1 0 43158 0 1 40805
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_2
timestamp 1654408082
transform 1 0 43158 0 1 43345
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_3
timestamp 1654408082
transform 1 0 43158 0 1 44495
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654408082
transform 1 0 -27088 0 1 49146
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1654408082
transform 1 0 -25892 0 1 49146
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1654408082
transform 1 0 41962 0 1 39535
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1654408082
transform 1 0 45458 0 1 39535
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1654408082
transform 1 0 41962 0 1 40805
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1654408082
transform 1 0 45458 0 1 40805
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1654408082
transform 1 0 41962 0 1 43345
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1654408082
transform 1 0 45458 0 1 43345
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1654408082
transform 1 0 41962 0 1 44495
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1654408082
transform 1 0 45458 0 1 44495
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654408082
transform 1 0 39938 0 1 39535
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_1
timestamp 1654408082
transform 1 0 39938 0 1 40805
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_2
timestamp 1654408082
transform 1 0 39938 0 1 43345
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_3
timestamp 1654408082
transform 1 0 39938 0 1 44495
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654408082
transform 1 0 -25984 0 1 49146
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1654408082
transform 1 0 -26720 0 1 49146
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1654408082
transform 1 0 43066 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1654408082
transform 1 0 42330 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1654408082
transform 1 0 45366 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1654408082
transform 1 0 41870 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1654408082
transform 1 0 39846 0 1 39535
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1654408082
transform 1 0 39846 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1654408082
transform 1 0 43066 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1654408082
transform 1 0 42330 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1654408082
transform 1 0 41870 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1654408082
transform 1 0 45366 0 1 40805
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1654408082
transform 1 0 39846 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1654408082
transform 1 0 43066 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1654408082
transform 1 0 42330 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1654408082
transform 1 0 41870 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1654408082
transform 1 0 45366 0 1 43345
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1654408082
transform 1 0 39846 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1654408082
transform 1 0 43066 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1654408082
transform 1 0 42330 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1654408082
transform 1 0 41870 0 1 44495
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1654408082
transform 1 0 45366 0 1 44495
box -38 -48 130 592
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/transmission_gate
timestamp 1654408082
transform 1 0 -26675 0 1 13627
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1654408082
transform 1 0 -6071 0 -1 14526
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1654408082
transform 1 0 -26675 0 1 5859
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1654408082
transform 1 0 -2967 0 1 12195
box -216 -51 1283 1063
use transmission_gate  transmission_gate_4
timestamp 1654408082
transform 1 0 -2967 0 1 10595
box -216 -51 1283 1063
use transmission_gate  transmission_gate_5
timestamp 1654408082
transform 1 0 -2967 0 1 8995
box -216 -51 1283 1063
use transmission_gate  transmission_gate_6
timestamp 1654408082
transform 1 0 -2967 0 1 7395
box -216 -51 1283 1063
use transmission_gate  transmission_gate_7
timestamp 1654408082
transform 1 0 -6071 0 1 5869
box -216 -51 1283 1063
use transmission_gate  transmission_gate_8
timestamp 1654408082
transform 0 1 -6231 -1 0 11991
box -216 -51 1283 1063
use transmission_gate  transmission_gate_9
timestamp 1654408082
transform 0 1 -6231 1 0 8354
box -216 -51 1283 1063
use transmission_gate  transmission_gate_10
timestamp 1654408082
transform -1 0 -1901 0 -1 15522
box -216 -51 1283 1063
use transmission_gate  transmission_gate_11
timestamp 1654408082
transform -1 0 -1903 0 -1 6110
box -216 -51 1283 1063
use transmission_gate  transmission_gate_12
timestamp 1654408082
transform 0 -1 3839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_13
timestamp 1654408082
transform 0 -1 5839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_14
timestamp 1654408082
transform 0 -1 7839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_15
timestamp 1654408082
transform 0 -1 9839 1 0 17833
box -216 -51 1283 1063
use transmission_gate  transmission_gate_16
timestamp 1654408082
transform 0 1 -826 -1 0 18922
box -216 -51 1283 1063
use transmission_gate  transmission_gate_17
timestamp 1654408082
transform 0 -1 3845 1 0 22174
box -216 -51 1283 1063
use transmission_gate  transmission_gate_18
timestamp 1654408082
transform 0 1 9022 1 0 22174
box -216 -51 1283 1063
use transmission_gate  transmission_gate_19
timestamp 1654408082
transform -1 0 6948 0 1 23654
box -216 -51 1283 1063
use transmission_gate  transmission_gate_20
timestamp 1654408082
transform 0 -1 3873 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_21
timestamp 1654408082
transform 0 -1 5873 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_22
timestamp 1654408082
transform 0 1 6861 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_23
timestamp 1654408082
transform 0 -1 9873 1 0 34868
box -216 -51 1283 1063
use transmission_gate  transmission_gate_24
timestamp 1654408082
transform 1 0 1359 0 -1 38947
box -216 -51 1283 1063
use transmission_gate  transmission_gate_25
timestamp 1654408082
transform 1 0 1007 0 -1 37197
box -216 -51 1283 1063
use transmission_gate  transmission_gate_26
timestamp 1654408082
transform -1 0 -7618 0 -1 51315
box -216 -51 1283 1063
use transmission_gate  transmission_gate_27
timestamp 1654408082
transform 1 0 -13548 0 1 27131
box -216 -51 1283 1063
use transmission_gate  transmission_gate_28
timestamp 1654408082
transform 1 0 -13548 0 1 25531
box -216 -51 1283 1063
use transmission_gate  transmission_gate_29
timestamp 1654408082
transform 1 0 -13548 0 1 23931
box -216 -51 1283 1063
use transmission_gate  transmission_gate_30
timestamp 1654408082
transform 1 0 -13548 0 1 22331
box -216 -51 1283 1063
use transmission_gate  transmission_gate_31
timestamp 1654408082
transform 1 0 -26607 0 1 24644
box -216 -51 1283 1063
use transmission_gate  transmission_gate_32
timestamp 1654408082
transform 1 0 -26607 0 1 17101
box -216 -51 1283 1063
<< labels >>
flabel metal1 40521 5685 40521 5685 1 FreeSans 400 0 0 0 out
flabel metal1 40521 -1255 40521 -1255 1 FreeSans 400 0 0 0 out
flabel metal3 -56975 25027 -56975 25027 1 FreeSans 16000 0 0 0 ip
flabel metal3 -57006 17492 -57006 17492 1 FreeSans 16000 0 0 0 in
flabel metal3 -56866 37447 -56866 37447 1 FreeSans 16000 0 0 0 op
flabel metal3 -56957 50045 -56957 50045 1 FreeSans 16000 0 0 0 rst_n
flabel metal3 -16863 90254 -16863 90254 1 FreeSans 16000 0 0 0 a_probe_1
flabel metal3 11101 90277 11101 90277 1 FreeSans 16000 0 0 0 i_bias_2
flabel metal3 23035 90264 23035 90264 1 FreeSans 16000 0 0 0 clk
flabel metal3 62718 76068 62718 76068 1 FreeSans 16000 0 0 0 a_mod_grp_ctrl_1
flabel metal3 62776 68706 62776 68706 1 FreeSans 16000 0 0 0 a_mod_grp_ctrl_0
flabel metal3 62776 61266 62776 61266 1 FreeSans 16000 0 0 0 debug
flabel metal3 62793 55222 62793 55222 1 FreeSans 16000 0 0 0 d_clk_grp_1_ctrl_0
flabel metal3 62783 50992 62783 50992 1 FreeSans 16000 0 0 0 d_clk_grp_1_ctrl_1
flabel metal3 62738 47250 62738 47250 1 FreeSans 16000 0 0 0 d_probe_0
flabel metal3 62730 43660 62730 43660 1 FreeSans 16000 0 0 0 d_probe_1
flabel metal3 62755 33541 62755 33541 1 FreeSans 16000 0 0 0 d_probe_2
flabel metal3 62821 30323 62821 30323 1 FreeSans 16000 0 0 0 d_probe_3
flabel metal3 62686 40251 62686 40251 1 FreeSans 16000 0 0 0 d_clk_grp_2_ctrl_0
flabel metal3 62811 36995 62811 36995 1 FreeSans 16000 0 0 0 d_clk_grp_2_ctrl_1
flabel metal3 62769 22636 62769 22636 1 FreeSans 16000 0 0 0 a_probe_0
flabel metal3 62810 5693 62810 5693 1 FreeSans 16000 0 0 0 a_probe_2
flabel metal3 62725 -1241 62725 -1241 1 FreeSans 16000 0 0 0 a_probe_3
flabel metal3 -998 -23902 -998 -23902 1 FreeSans 16000 0 0 0 i_bias_1
flabel metal5 -54092 90092 -54092 90092 1 FreeSans 16000 0 0 0 VDD
flabel metal5 -50052 90052 -50052 90052 1 FreeSans 16000 0 0 0 VSS
flabel metal5 55900 90138 55900 90138 1 FreeSans 16000 0 0 0 VDD
flabel metal5 59914 90094 59914 90094 1 FreeSans 16000 0 0 0 VSS
flabel metal5 -54102 -23638 -54102 -23638 1 FreeSans 16000 0 0 0 VDD
flabel metal5 -50108 -23638 -50108 -23638 1 FreeSans 16000 0 0 0 VSS
flabel metal5 55928 -23634 55928 -23634 1 FreeSans 16000 0 0 0 VDD
flabel metal5 59912 -23508 59912 -23508 1 FreeSans 16000 0 0 0 VSS
<< end >>
