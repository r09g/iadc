magic
tech sky130A
magscale 1 2
timestamp 1652659422
<< nwell >>
rect -647 -356 647 294
<< pmos >>
rect -447 -137 -417 137
rect -351 -137 -321 137
rect -255 -137 -225 137
rect -159 -137 -129 137
rect -63 -137 -33 137
rect 33 -137 63 137
rect 129 -137 159 137
rect 225 -137 255 137
rect 321 -137 351 137
rect 417 -137 447 137
<< pdiff >>
rect -509 125 -447 137
rect -509 -125 -497 125
rect -463 -125 -447 125
rect -509 -137 -447 -125
rect -417 125 -351 137
rect -417 -125 -401 125
rect -367 -125 -351 125
rect -417 -137 -351 -125
rect -321 125 -255 137
rect -321 -125 -305 125
rect -271 -125 -255 125
rect -321 -137 -255 -125
rect -225 125 -159 137
rect -225 -125 -209 125
rect -175 -125 -159 125
rect -225 -137 -159 -125
rect -129 125 -63 137
rect -129 -125 -113 125
rect -79 -125 -63 125
rect -129 -137 -63 -125
rect -33 125 33 137
rect -33 -125 -17 125
rect 17 -125 33 125
rect -33 -137 33 -125
rect 63 125 129 137
rect 63 -125 79 125
rect 113 -125 129 125
rect 63 -137 129 -125
rect 159 125 225 137
rect 159 -125 175 125
rect 209 -125 225 125
rect 159 -137 225 -125
rect 255 125 321 137
rect 255 -125 271 125
rect 305 -125 321 125
rect 255 -137 321 -125
rect 351 125 417 137
rect 351 -125 367 125
rect 401 -125 417 125
rect 351 -137 417 -125
rect 447 125 509 137
rect 447 -125 463 125
rect 497 -125 509 125
rect 447 -137 509 -125
<< pdiffc >>
rect -497 -125 -463 125
rect -401 -125 -367 125
rect -305 -125 -271 125
rect -209 -125 -175 125
rect -113 -125 -79 125
rect -17 -125 17 125
rect 79 -125 113 125
rect 175 -125 209 125
rect 271 -125 305 125
rect 367 -125 401 125
rect 463 -125 497 125
<< nsubdiff >>
rect -611 224 -515 258
rect 515 224 611 258
rect -611 162 -577 224
rect 577 162 611 224
rect -611 -286 -577 -224
rect 577 -286 611 -224
rect -611 -320 -515 -286
rect 515 -320 611 -286
<< nsubdiffcont >>
rect -515 224 515 258
rect -611 -224 -577 162
rect 577 -224 611 162
rect -515 -320 515 -286
<< poly >>
rect -447 137 -417 163
rect -351 137 -321 163
rect -255 137 -225 163
rect -159 137 -129 163
rect -63 137 -33 163
rect 33 137 63 163
rect 129 137 159 163
rect 225 137 255 163
rect 321 137 351 163
rect 417 137 447 163
rect -447 -168 -417 -137
rect -351 -168 -321 -137
rect -255 -168 -225 -137
rect -159 -168 -129 -137
rect -63 -168 -33 -137
rect 33 -168 63 -137
rect 129 -168 159 -137
rect 225 -168 255 -137
rect 321 -168 351 -137
rect 417 -168 447 -137
rect -513 -184 513 -168
rect -513 -218 -497 -184
rect -463 -218 -305 -184
rect -271 -218 -113 -184
rect -79 -218 79 -184
rect 113 -218 271 -184
rect 305 -218 463 -184
rect 497 -218 513 -184
rect -513 -234 513 -218
<< polycont >>
rect -497 -218 -463 -184
rect -305 -218 -271 -184
rect -113 -218 -79 -184
rect 79 -218 113 -184
rect 271 -218 305 -184
rect 463 -218 497 -184
<< locali >>
rect -611 224 -515 258
rect 515 224 611 258
rect -611 162 -577 224
rect 577 162 611 224
rect -497 125 -463 141
rect -497 -141 -463 -125
rect -401 125 -367 141
rect -401 -141 -367 -125
rect -305 125 -271 141
rect -305 -141 -271 -125
rect -209 125 -175 141
rect -209 -141 -175 -125
rect -113 125 -79 141
rect -113 -141 -79 -125
rect -17 125 17 141
rect -17 -141 17 -125
rect 79 125 113 141
rect 79 -141 113 -125
rect 175 125 209 141
rect 175 -141 209 -125
rect 271 125 305 141
rect 271 -141 305 -125
rect 367 125 401 141
rect 367 -141 401 -125
rect 463 125 497 141
rect 463 -141 497 -125
rect -513 -218 -497 -184
rect -463 -218 -447 -184
rect -321 -218 -305 -184
rect -271 -218 -255 -184
rect -129 -218 -113 -184
rect -79 -218 -63 -184
rect 63 -218 79 -184
rect 113 -218 129 -184
rect 255 -218 271 -184
rect 305 -218 321 -184
rect 447 -218 463 -184
rect 497 -218 513 -184
rect -611 -286 -577 -224
rect 577 -286 611 -224
rect -611 -320 -515 -286
rect 515 -320 611 -286
<< viali >>
rect -497 -125 -463 125
rect -401 -125 -367 125
rect -305 -125 -271 125
rect -209 -125 -175 125
rect -113 -125 -79 125
rect -17 -125 17 125
rect 79 -125 113 125
rect 175 -125 209 125
rect 271 -125 305 125
rect 367 -125 401 125
rect 463 -125 497 125
rect -497 -218 -463 -184
rect -305 -218 -271 -184
rect -113 -218 -79 -184
rect 79 -218 113 -184
rect 271 -218 305 -184
rect 463 -218 497 -184
<< metal1 >>
rect -503 125 -457 137
rect -503 -125 -497 125
rect -463 -125 -457 125
rect -503 -137 -457 -125
rect -407 125 -361 137
rect -407 -125 -401 125
rect -367 -125 -361 125
rect -407 -137 -361 -125
rect -311 125 -265 137
rect -311 -125 -305 125
rect -271 -125 -265 125
rect -311 -137 -265 -125
rect -215 125 -169 137
rect -215 -125 -209 125
rect -175 -125 -169 125
rect -215 -137 -169 -125
rect -119 125 -73 137
rect -119 -125 -113 125
rect -79 -125 -73 125
rect -119 -137 -73 -125
rect -23 125 23 137
rect -23 -125 -17 125
rect 17 -125 23 125
rect -23 -137 23 -125
rect 73 125 119 137
rect 73 -125 79 125
rect 113 -125 119 125
rect 73 -137 119 -125
rect 169 125 215 137
rect 169 -125 175 125
rect 209 -125 215 125
rect 169 -137 215 -125
rect 265 125 311 137
rect 265 -125 271 125
rect 305 -125 311 125
rect 265 -137 311 -125
rect 361 125 407 137
rect 361 -125 367 125
rect 401 -125 407 125
rect 361 -137 407 -125
rect 457 125 503 137
rect 457 -125 463 125
rect 497 -125 503 125
rect 457 -137 503 -125
rect -513 -184 -447 -176
rect -513 -218 -497 -184
rect -463 -218 -447 -184
rect -513 -227 -447 -218
rect -321 -184 -255 -176
rect -321 -218 -305 -184
rect -271 -218 -255 -184
rect -321 -227 -255 -218
rect -129 -184 -63 -176
rect -129 -218 -113 -184
rect -79 -218 -63 -184
rect -129 -227 -63 -218
rect 63 -184 129 -176
rect 63 -218 79 -184
rect 113 -218 129 -184
rect 63 -227 129 -218
rect 255 -184 321 -176
rect 255 -218 271 -184
rect 305 -218 321 -184
rect 255 -227 321 -218
rect 447 -184 513 -176
rect 447 -218 463 -184
rect 497 -218 513 -184
rect 447 -227 513 -218
<< properties >>
string FIXED_BBOX -594 -303 594 303
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.37 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
