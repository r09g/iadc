* NGSPICE file created from digital_filter.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 Y A VGND VPWR VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPWR VGND VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_16 Y A VGND VPWR VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_1 X A1 B1 A2 VGND VPWR VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__fa_2 COUT SUM A B CIN VGND VPWR VNB VPB
X0 a_1171_369# CIN a_1086_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND CIN a_829_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1086_47# SUM VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 COUT a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_829_369# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR CIN a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_473_371# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X7 a_294_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A a_473_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X9 a_829_369# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_829_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_829_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_473_371# CIN a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X13 a_473_47# CIN a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_473_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR a_1086_47# SUM VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_80_21# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 COUT a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 SUM a_1086_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_80_21# B a_289_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X20 a_80_21# B a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A a_473_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 SUM a_1086_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR a_80_21# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_289_371# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X25 a_1194_47# CIN a_1086_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1086_47# a_80_21# a_829_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND A a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1266_371# B a_1171_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X29 VPWR A a_1266_371# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X30 a_1266_47# B a_1194_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1086_47# a_80_21# a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_1 C B Y D A VPWR VGND VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinvlp_2 VGND VPWR Y A VNB VPB
X0 Y A a_150_67# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X2 a_150_67# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__sdlclkp_4 SCE CLK GCLK GATE VGND VPWR VNB VPB
X0 a_257_147# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_109_369# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_315# a_287_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_287_413# a_257_147# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 VPWR a_257_147# a_257_243# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_257_147# a_257_243# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_465_315# a_383_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1127_47# a_465_315# a_1045_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_287_413# a_257_243# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_383_413# a_257_147# a_287_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND CLK a_1127_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_257_147# CLK VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_47# GATE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VPWR CLK a_1045_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1045_47# a_465_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_395_47# a_257_243# a_287_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VGND a_465_315# a_395_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND SCE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_465_315# a_287_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 Y A VPWR VGND VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__nand3_1 Y A C B VGND VPWR VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__ha_2 VGND VPWR A COUT SUM B VNB VPB
X0 VPWR A a_342_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_766_47# B a_342_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B a_389_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 COUT a_342_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_342_199# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_468_369# B a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# a_342_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_389_47# a_342_199# a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_389_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 COUT a_342_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_342_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_79_21# SUM VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR a_79_21# SUM VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_342_199# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 SUM a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A a_468_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 SUM a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 B1 Y A2 VPWR VGND VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_0 VPWR VGND X B A VNB VPB
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__nor3_1 C Y A B VGND VPWR VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1 B X A VPWR VGND VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt digital_filter clk rst_n sclk cs_n data_in data_out[11] data_out[10] data_out[9]
+ data_out[8] data_out[7] data_out[6] data_out[5] data_out[4] data_out[3] data_out[2]
+ data_out[1] data_out[0] new_data serial_data_out VSS VDD
Xsky130_fd_sc_hd__decap_6_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_7 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__fa_2_6/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_42 sky130_fd_sc_hd__dfxtp_1_42/Q sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_24/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_20 data_out[4] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__o21a_1_3/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_31 sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_3/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_64 sky130_fd_sc_hd__nor2_1_1/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_29/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_53 sky130_fd_sc_hd__fa_2_6/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_13/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_4 sky130_fd_sc_hd__dfxtp_1_4/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_2/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_9 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__fa_2_3/B
+ sky130_fd_sc_hd__nor2_1_6/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_6_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_8 sky130_fd_sc_hd__nor2_1_6/A sky130_fd_sc_hd__fa_2_4/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_43 sky130_fd_sc_hd__o21a_1_2/A2 sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_23/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_32 sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_4/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_10 sky130_fd_sc_hd__a22o_1_7/B1 sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_8/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_21 data_out[5] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__dfxtp_1_44/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_54 sky130_fd_sc_hd__fa_2_7/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_12/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_5 sky130_fd_sc_hd__dfxtp_1_5/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_3/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__a22o_1_0 data_out[11] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_0/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_3/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_6_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_9 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__fa_2_2/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_22 data_out[6] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__o21a_1_2/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_33 sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_5/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_44 sky130_fd_sc_hd__dfxtp_1_44/Q sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_21/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_11 sky130_fd_sc_hd__a22o_1_8/B1 sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_9/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_55 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_11/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_6 sky130_fd_sc_hd__dfxtp_1_6/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_4/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__a22o_1_1 data_out[10] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_1/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_4/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_6_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__dfxtp_1_23 data_out[7] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__dfxtp_1_42/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_34 sky130_fd_sc_hd__ha_2_2/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_6/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_56 sky130_fd_sc_hd__fa_2_1/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_36/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_12 sky130_fd_sc_hd__a22o_1_9/B1 sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_10/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_45 sky130_fd_sc_hd__o21a_1_3/A2 sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_22/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_7 sky130_fd_sc_hd__dfxtp_1_7/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_5/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a22o_1_2 data_out[9] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_2/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_5/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_16_0 sky130_fd_sc_hd__dfxtp_1_1/CLK sky130_fd_sc_hd__clkinv_4_1/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__decap_6_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__dfxtp_1_24 data_out[8] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__o21a_1_1/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_57 sky130_fd_sc_hd__fa_2_0/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_37/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_46 sky130_fd_sc_hd__o21a_1_4/A2 sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_20/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_35 sky130_fd_sc_hd__ha_2_1/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_7/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_13 sky130_fd_sc_hd__dfxtp_1_13/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_11/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_8 sky130_fd_sc_hd__dfxtp_1_8/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_6/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a22o_1_3 data_out[8] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_3/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_6/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_6_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__o21a_1_0 sky130_fd_sc_hd__o21a_1_0/X sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__xnor2_1_0/B sky130_fd_sc_hd__o21a_1_0/A2 VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_25 data_out[9] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__dfxtp_1_40/Q
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_58 sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_35/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_47 sky130_fd_sc_hd__fa_2_0/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_19/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_36 sky130_fd_sc_hd__ha_2_0/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_8/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_14 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__o21ai_1_0/A1 VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_9 sky130_fd_sc_hd__dfxtp_1_9/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_7/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a22o_1_4 data_out[7] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_4/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_7/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__fa_2_0 sky130_fd_sc_hd__o21a_1_4/A1 sky130_fd_sc_hd__fa_2_0/SUM
+ sky130_fd_sc_hd__fa_2_0/A sky130_fd_sc_hd__fa_2_0/B sky130_fd_sc_hd__fa_2_0/CIN
+ VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__nand4_1_0 sky130_fd_sc_hd__ha_2_2/A sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__nor3_1_0/C
+ sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__ha_2_6/B VDD VSS VSS VDD sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__clkinvlp_2_0 VSS VDD sky130_fd_sc_hd__nor2_1_4/A sky130_fd_sc_hd__dfxtp_1_44/Q
+ VSS VDD sky130_fd_sc_hd__clkinvlp_2
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_0/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_6_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__o21a_1_1 sky130_fd_sc_hd__o21a_1_1/X sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__o21a_1_1/A2 VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__xnor2_1_0 VSS VDD sky130_fd_sc_hd__xnor2_1_0/B sky130_fd_sc_hd__xnor2_1_0/Y
+ sky130_fd_sc_hd__xnor2_1_0/A VSS VDD sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_26 data_out[10] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__o21a_1_0/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_59 sky130_fd_sc_hd__fa_2_3/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_34/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_48 sky130_fd_sc_hd__fa_2_1/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_18/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_15 sky130_fd_sc_hd__o21ai_1_0/A1 sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sclk VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_37 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_9/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__clkinv_4_0/A sky130_fd_sc_hd__clkinv_4_1/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__fa_2_1 sky130_fd_sc_hd__fa_2_0/CIN sky130_fd_sc_hd__fa_2_1/SUM sky130_fd_sc_hd__fa_2_1/A
+ sky130_fd_sc_hd__fa_2_1/B sky130_fd_sc_hd__fa_2_1/CIN VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_5 data_out[6] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_5/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_8/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__o21a_1_2 sky130_fd_sc_hd__o21a_1_2/X sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__o21a_1_2/A2 VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_38 sky130_fd_sc_hd__o21a_1_0/A2 sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_28/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__xnor2_1_1 VSS VDD sky130_fd_sc_hd__xnor2_1_1/B sky130_fd_sc_hd__xnor2_1_1/Y
+ sky130_fd_sc_hd__fa_2_0/B VSS VDD sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_49 sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_17/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_27 data_out[11] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__xnor2_1_0/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_16 data_out[0] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__fa_2_2/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_1/Y
+ VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__fa_2_2 sky130_fd_sc_hd__fa_2_1/CIN sky130_fd_sc_hd__fa_2_2/SUM sky130_fd_sc_hd__fa_2_2/A
+ sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__fa_2_2/CIN VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_6 data_out[5] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_6/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_9/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__nor2_1_2/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__o21a_1_3 sky130_fd_sc_hd__o21a_1_3/X sky130_fd_sc_hd__o21a_1_3/A1
+ sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__o21a_1_3/A2 VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_39 sky130_fd_sc_hd__xnor2_1_0/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_27/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_28 new_data sky130_fd_sc_hd__dfxtp_1_1/CLK sky130_fd_sc_hd__and2_0_1/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_17 data_out[1] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__fa_2_1/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_3 sky130_fd_sc_hd__fa_2_2/CIN sky130_fd_sc_hd__fa_2_3/SUM sky130_fd_sc_hd__fa_2_3/A
+ sky130_fd_sc_hd__fa_2_3/B sky130_fd_sc_hd__fa_2_3/CIN VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_7 data_out[4] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_7/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__a22o_1_7/B1 VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_1_10 sky130_fd_sc_hd__nor2_1_6/B sky130_fd_sc_hd__fa_2_5/B
+ sky130_fd_sc_hd__nor2_1_7/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_4_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__nor2_1_3/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__sdlclkp_4_0 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__clkinv_4_1/A
+ sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__o21ai_1_0/Y VSS VDD VSS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__decap_3_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_29 sky130_fd_sc_hd__ha_2_6/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_0/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_18 data_out[2] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__fa_2_0/A
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21a_1_4 sky130_fd_sc_hd__o21a_1_4/X sky130_fd_sc_hd__o21a_1_4/A1
+ sky130_fd_sc_hd__o21a_1_4/B1 sky130_fd_sc_hd__o21a_1_4/A2 VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__a22o_1_8 data_out[3] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_8/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__a22o_1_8/B1 VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__fa_2_4 sky130_fd_sc_hd__fa_2_3/CIN sky130_fd_sc_hd__fa_2_4/SUM sky130_fd_sc_hd__fa_2_4/A
+ sky130_fd_sc_hd__fa_2_4/B sky130_fd_sc_hd__fa_2_4/CIN VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_10 data_out[1] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_10/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__dfxtp_1_13/Q VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_2_0 sky130_fd_sc_hd__clkinv_4_0/A clk VDD VSS VSS VDD sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__decap_4_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__sdlclkp_4_1 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__clkinv_4_1/A
+ sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__and2_0_1/X VSS VDD VSS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__nor2_1_4/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_5 sky130_fd_sc_hd__o21a_1_5/X sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__xnor2_1_1/B sky130_fd_sc_hd__fa_2_1/B VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_19 data_out[3] sky130_fd_sc_hd__dfxtp_1_27/CLK sky130_fd_sc_hd__o21a_1_4/A2
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_5 sky130_fd_sc_hd__fa_2_4/CIN sky130_fd_sc_hd__fa_2_5/SUM sky130_fd_sc_hd__fa_2_5/A
+ sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_5/CIN VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_9 data_out[2] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_9/X
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__a22o_1_9/B1 VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_11 data_out[0] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_11/X
+ sky130_fd_sc_hd__nand2_1_0/B serial_data_out VDD VSS VSS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__nor2_1_5/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_6 sky130_fd_sc_hd__o21a_1_6/X sky130_fd_sc_hd__nor2_1_6/Y
+ sky130_fd_sc_hd__nor2_1_5/B sky130_fd_sc_hd__fa_2_3/B VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__fa_2_6 sky130_fd_sc_hd__fa_2_5/CIN sky130_fd_sc_hd__fa_2_6/SUM sky130_fd_sc_hd__fa_2_6/A
+ sky130_fd_sc_hd__fa_2_6/B sky130_fd_sc_hd__fa_2_6/CIN VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_4_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_6 sky130_fd_sc_hd__nor2_1_6/B sky130_fd_sc_hd__nor2_1_6/Y
+ sky130_fd_sc_hd__nor2_1_6/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_7 sky130_fd_sc_hd__o21a_1_7/X sky130_fd_sc_hd__nor2_1_7/Y
+ sky130_fd_sc_hd__nor2_1_6/B sky130_fd_sc_hd__fa_2_5/B VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__fa_2_7 sky130_fd_sc_hd__fa_2_6/CIN sky130_fd_sc_hd__fa_2_7/SUM sky130_fd_sc_hd__fa_2_7/A
+ sky130_fd_sc_hd__fa_2_7/B sky130_fd_sc_hd__nor2_1_0/A VSS VDD VSS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__o21ai_1_0 VSS VDD sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__o21ai_1_0/A1
+ sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__o21ai_1_0/Y VSS VDD sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__decap_4_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_7 sky130_fd_sc_hd__nor2_1_7/B sky130_fd_sc_hd__nor2_1_7/Y
+ sky130_fd_sc_hd__nor2_1_7/A VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_8 sky130_fd_sc_hd__o21a_1_8/X sky130_fd_sc_hd__o21a_1_8/A1
+ sky130_fd_sc_hd__nor2_1_7/B sky130_fd_sc_hd__fa_2_7/B VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_4_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_9 sky130_fd_sc_hd__o21a_1_9/X data_in sky130_fd_sc_hd__o21a_1_9/B1
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD VSS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__decap_4_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_4_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_4_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand3_1_0 sky130_fd_sc_hd__nor3_1_0/B sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__ha_2_1/A VSS VDD VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_4_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand3_1_1 sky130_fd_sc_hd__nor2_1_4/B sky130_fd_sc_hd__o21a_1_4/A1
+ sky130_fd_sc_hd__o21a_1_3/A2 sky130_fd_sc_hd__o21a_1_4/A2 VSS VDD VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__nand3_1_2 sky130_fd_sc_hd__nor2_1_7/B data_in sky130_fd_sc_hd__fa_2_7/B
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD VSS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__diode_2_0 sclk VSS VDD VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__ha_2_0 VSS VDD sky130_fd_sc_hd__ha_2_0/A sky130_fd_sc_hd__xor2_1_0/A
+ sky130_fd_sc_hd__ha_2_0/SUM sky130_fd_sc_hd__ha_2_0/B VSS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__ha_2_1 VSS VDD sky130_fd_sc_hd__ha_2_1/A sky130_fd_sc_hd__ha_2_0/B
+ sky130_fd_sc_hd__ha_2_1/SUM sky130_fd_sc_hd__ha_2_1/B VSS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__ha_2_2 VSS VDD sky130_fd_sc_hd__ha_2_2/A sky130_fd_sc_hd__ha_2_1/B
+ sky130_fd_sc_hd__ha_2_2/SUM sky130_fd_sc_hd__ha_2_2/B VSS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_0 sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__nor2_1_2/Y
+ sky130_fd_sc_hd__and2_0_26/A sky130_fd_sc_hd__nor2_1_2/B VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_30 VDD VSS sky130_fd_sc_hd__and2_0_30/X rst_n sky130_fd_sc_hd__o21a_1_8/X
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_3 VSS VDD sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__ha_2_2/B
+ sky130_fd_sc_hd__ha_2_3/SUM sky130_fd_sc_hd__ha_2_3/B VSS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_1 sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__nor2_1_3/Y
+ sky130_fd_sc_hd__and2_0_24/A sky130_fd_sc_hd__nor2_1_3/B VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_31 VDD VSS sky130_fd_sc_hd__and2_0_31/X rst_n sky130_fd_sc_hd__and2_0_31/A
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_20 VDD VSS sky130_fd_sc_hd__and2_0_20/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__o21a_1_4/X VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_4 VSS VDD sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__ha_2_3/B
+ sky130_fd_sc_hd__ha_2_4/SUM sky130_fd_sc_hd__ha_2_4/B VSS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_2 sky130_fd_sc_hd__nor2_1_4/A sky130_fd_sc_hd__nor2_1_4/Y
+ sky130_fd_sc_hd__and2_0_21/A sky130_fd_sc_hd__nor2_1_4/B VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_21 VDD VSS sky130_fd_sc_hd__and2_0_21/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__and2_0_21/A VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_32 VDD VSS sky130_fd_sc_hd__and2_0_32/X rst_n sky130_fd_sc_hd__o21a_1_7/X
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_10 VDD VSS sky130_fd_sc_hd__nor2_1_0/A sky130_fd_sc_hd__nor2_1_1/B
+ sky130_fd_sc_hd__nor2_1_1/A VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_5 VSS VDD sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__ha_2_4/B
+ sky130_fd_sc_hd__ha_2_5/SUM sky130_fd_sc_hd__ha_2_5/B VSS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_3 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__nor2_1_5/Y
+ sky130_fd_sc_hd__and2_0_35/A sky130_fd_sc_hd__nor2_1_5/B VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_33 VDD VSS sky130_fd_sc_hd__and2_0_33/X rst_n sky130_fd_sc_hd__and2_0_33/A
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__and2_0_11 VDD VSS sky130_fd_sc_hd__and2_0_11/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__nor2_1_0/Y VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_22 VDD VSS sky130_fd_sc_hd__and2_0_22/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__o21a_1_3/X VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_6 VSS VDD sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__ha_2_5/B
+ sky130_fd_sc_hd__ha_2_6/SUM sky130_fd_sc_hd__ha_2_6/B VSS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__conb_1_0 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_0/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_4 sky130_fd_sc_hd__nor2_1_6/A sky130_fd_sc_hd__nor2_1_6/Y
+ sky130_fd_sc_hd__and2_0_33/A sky130_fd_sc_hd__nor2_1_6/B VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_23 VDD VSS sky130_fd_sc_hd__and2_0_23/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__o21a_1_2/X VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_34 VDD VSS sky130_fd_sc_hd__and2_0_34/X rst_n sky130_fd_sc_hd__o21a_1_6/X
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_12 VDD VSS sky130_fd_sc_hd__and2_0_12/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_7/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_1 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_1/HI
+ VDD VSS VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__and2_0_0 VDD VSS sky130_fd_sc_hd__and2_0_0/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__and2_0_0/A VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_8_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_5 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nor2_1_7/Y
+ sky130_fd_sc_hd__and2_0_31/A sky130_fd_sc_hd__nor2_1_7/B VDD VSS VSS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_24 VDD VSS sky130_fd_sc_hd__and2_0_24/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__and2_0_24/A VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_35 VDD VSS sky130_fd_sc_hd__and2_0_35/X rst_n sky130_fd_sc_hd__and2_0_35/A
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_13 VDD VSS sky130_fd_sc_hd__and2_0_13/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_6/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_1_0/B
+ sky130_fd_sc_hd__nand2_1_0/A VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_1 VDD VSS sky130_fd_sc_hd__and2_0_1/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__nor3_1_0/Y VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_8_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_6_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_25 VDD VSS sky130_fd_sc_hd__and2_0_25/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__o21a_1_1/X VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_36 VDD VSS sky130_fd_sc_hd__and2_0_36/X rst_n sky130_fd_sc_hd__o21a_1_5/X
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_14 VDD VSS sky130_fd_sc_hd__and2_0_14/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_5/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__and2_0_2 VDD VSS sky130_fd_sc_hd__and2_0_2/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__ha_2_6/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand2_1_1/Y new_data cs_n VSS VDD VSS
+ VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_6_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_26 VDD VSS sky130_fd_sc_hd__and2_0_26/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__and2_0_26/A VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_37 VDD VSS sky130_fd_sc_hd__and2_0_37/X rst_n sky130_fd_sc_hd__xnor2_1_1/Y
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_15 VDD VSS sky130_fd_sc_hd__and2_0_15/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_4/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__nand2_1_0/B cs_n VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__ha_2_0/A
+ sky130_fd_sc_hd__ha_2_4/A VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_3 VDD VSS sky130_fd_sc_hd__and2_0_3/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__ha_2_5/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_6_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__nand2_1_1/Y
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__and2_0_27 VDD VSS sky130_fd_sc_hd__and2_0_27/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__xnor2_1_0/Y VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_16 VDD VSS sky130_fd_sc_hd__and2_0_16/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_3/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_8_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__o21a_1_4/B1 sky130_fd_sc_hd__o21a_1_4/A2
+ sky130_fd_sc_hd__o21a_1_4/A1 VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_4 VDD VSS sky130_fd_sc_hd__and2_0_4/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__ha_2_4/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor3_1_0 sky130_fd_sc_hd__nor3_1_0/C sky130_fd_sc_hd__nor3_1_0/Y
+ sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__nor3_1_0/B VSS VDD VSS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__decap_6_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__and2_0_0/A sky130_fd_sc_hd__ha_2_6/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_28 VDD VSS sky130_fd_sc_hd__and2_0_28/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__o21a_1_0/X VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_17 VDD VSS sky130_fd_sc_hd__and2_0_17/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_2/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__and2_0_5 VDD VSS sky130_fd_sc_hd__and2_0_5/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__ha_2_3/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__xnor2_1_0/B sky130_fd_sc_hd__o21a_1_0/A2
+ sky130_fd_sc_hd__nor2_1_2/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_6_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_29 VDD VSS sky130_fd_sc_hd__and2_0_29/X rst_n sky130_fd_sc_hd__o21a_1_9/X
+ VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_18 VDD VSS sky130_fd_sc_hd__and2_0_18/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_1/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__o21a_1_3/A1 sky130_fd_sc_hd__o21a_1_4/B1
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_60 sky130_fd_sc_hd__fa_2_4/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_33/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_0 sky130_fd_sc_hd__and2_0_9/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__dfxtp_1_1/Q VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__nand2_1_5 sky130_fd_sc_hd__nor2_1_2/B sky130_fd_sc_hd__o21a_1_1/A2
+ sky130_fd_sc_hd__nor2_1_3/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_6 VDD VSS sky130_fd_sc_hd__and2_0_6/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__ha_2_2/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_6_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__dfxtp_1_42/Q
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_19 VDD VSS sky130_fd_sc_hd__and2_0_19/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ sky130_fd_sc_hd__fa_2_0/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_61 sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_32/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_50 sky130_fd_sc_hd__fa_2_3/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_16/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_1 sky130_fd_sc_hd__dfxtp_1_1/Q sky130_fd_sc_hd__dfxtp_1_1/CLK
+ rst_n VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__nand2_1_6 sky130_fd_sc_hd__nor2_1_3/B sky130_fd_sc_hd__o21a_1_2/A2
+ sky130_fd_sc_hd__nor2_1_4/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_7 VDD VSS sky130_fd_sc_hd__and2_0_7/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__ha_2_1/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor2_1_0 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/X
+ sky130_fd_sc_hd__xor2_1_0/A VDD VSS VSS VDD sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_6_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__dfxtp_1_40/Q
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_40 sky130_fd_sc_hd__dfxtp_1_40/Q sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_26/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_62 sky130_fd_sc_hd__fa_2_6/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_31/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_51 sky130_fd_sc_hd__fa_2_4/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_15/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_2 serial_data_out sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_0/X
+ VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_7 sky130_fd_sc_hd__o21a_1_9/B1 sky130_fd_sc_hd__nor2_1_1/A
+ data_in VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_8 VDD VSS sky130_fd_sc_hd__and2_0_8/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__ha_2_0/SUM VSS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_6_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_6 sky130_fd_sc_hd__o21a_1_8/A1 sky130_fd_sc_hd__o21a_1_9/B1
+ VSS VDD VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_41 sky130_fd_sc_hd__o21a_1_1/A2 sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_25/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_30 sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_2/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_63 sky130_fd_sc_hd__fa_2_7/B sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_30/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_52 sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__dfxtp_1_1/CLK
+ sky130_fd_sc_hd__and2_0_14/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_3 sky130_fd_sc_hd__dfxtp_1_3/Q sky130_fd_sc_hd__dfxtp_1_9/CLK
+ sky130_fd_sc_hd__a22o_1_1/X VDD VSS VSS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_8 sky130_fd_sc_hd__xnor2_1_1/B sky130_fd_sc_hd__fa_2_1/B
+ sky130_fd_sc_hd__nor2_1_5/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_9 VDD VSS sky130_fd_sc_hd__and2_0_9/X sky130_fd_sc_hd__and2_0_9/B
+ sky130_fd_sc_hd__xor2_1_0/X VSS VDD sky130_fd_sc_hd__and2_0
.ends

