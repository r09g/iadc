magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< nwell >>
rect -1489 -241 1489 241
<< pmoslvt >>
rect -1395 -140 -1275 140
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
rect 1275 -140 1395 140
<< pdiff >>
rect -1453 128 -1395 140
rect -1453 -128 -1441 128
rect -1407 -128 -1395 128
rect -1453 -140 -1395 -128
rect -1275 128 -1217 140
rect -1275 -128 -1263 128
rect -1229 -128 -1217 128
rect -1275 -140 -1217 -128
rect -1097 128 -1039 140
rect -1097 -128 -1085 128
rect -1051 -128 -1039 128
rect -1097 -140 -1039 -128
rect -919 128 -861 140
rect -919 -128 -907 128
rect -873 -128 -861 128
rect -919 -140 -861 -128
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
rect 861 128 919 140
rect 861 -128 873 128
rect 907 -128 919 128
rect 861 -140 919 -128
rect 1039 128 1097 140
rect 1039 -128 1051 128
rect 1085 -128 1097 128
rect 1039 -140 1097 -128
rect 1217 128 1275 140
rect 1217 -128 1229 128
rect 1263 -128 1275 128
rect 1217 -140 1275 -128
rect 1395 128 1453 140
rect 1395 -128 1407 128
rect 1441 -128 1453 128
rect 1395 -140 1453 -128
<< pdiffc >>
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
<< poly >>
rect -1373 221 -1297 237
rect -1373 205 -1357 221
rect -1395 187 -1357 205
rect -1313 205 -1297 221
rect -1195 221 -1119 237
rect -1195 205 -1179 221
rect -1313 187 -1275 205
rect -1395 140 -1275 187
rect -1217 187 -1179 205
rect -1135 205 -1119 221
rect -1017 221 -941 237
rect -1017 205 -1001 221
rect -1135 187 -1097 205
rect -1217 140 -1097 187
rect -1039 187 -1001 205
rect -957 205 -941 221
rect -839 221 -763 237
rect -839 205 -823 221
rect -957 187 -919 205
rect -1039 140 -919 187
rect -861 187 -823 205
rect -779 205 -763 221
rect -661 221 -585 237
rect -661 205 -645 221
rect -779 187 -741 205
rect -861 140 -741 187
rect -683 187 -645 205
rect -601 205 -585 221
rect -483 221 -407 237
rect -483 205 -467 221
rect -601 187 -563 205
rect -683 140 -563 187
rect -505 187 -467 205
rect -423 205 -407 221
rect -305 221 -229 237
rect -305 205 -289 221
rect -423 187 -385 205
rect -505 140 -385 187
rect -327 187 -289 205
rect -245 205 -229 221
rect -127 221 -51 237
rect -127 205 -111 221
rect -245 187 -207 205
rect -327 140 -207 187
rect -149 187 -111 205
rect -67 205 -51 221
rect 51 221 127 237
rect 51 205 67 221
rect -67 187 -29 205
rect -149 140 -29 187
rect 29 187 67 205
rect 111 205 127 221
rect 229 221 305 237
rect 229 205 245 221
rect 111 187 149 205
rect 29 140 149 187
rect 207 187 245 205
rect 289 205 305 221
rect 407 221 483 237
rect 407 205 423 221
rect 289 187 327 205
rect 207 140 327 187
rect 385 187 423 205
rect 467 205 483 221
rect 585 221 661 237
rect 585 205 601 221
rect 467 187 505 205
rect 385 140 505 187
rect 563 187 601 205
rect 645 205 661 221
rect 763 221 839 237
rect 763 205 779 221
rect 645 187 683 205
rect 563 140 683 187
rect 741 187 779 205
rect 823 205 839 221
rect 941 221 1017 237
rect 941 205 957 221
rect 823 187 861 205
rect 741 140 861 187
rect 919 187 957 205
rect 1001 205 1017 221
rect 1119 221 1195 237
rect 1119 205 1135 221
rect 1001 187 1039 205
rect 919 140 1039 187
rect 1097 187 1135 205
rect 1179 205 1195 221
rect 1297 221 1373 237
rect 1297 205 1313 221
rect 1179 187 1217 205
rect 1097 140 1217 187
rect 1275 187 1313 205
rect 1357 205 1373 221
rect 1357 187 1395 205
rect 1275 140 1395 187
rect -1395 -187 -1275 -140
rect -1395 -205 -1357 -187
rect -1373 -221 -1357 -205
rect -1313 -205 -1275 -187
rect -1217 -187 -1097 -140
rect -1217 -205 -1179 -187
rect -1313 -221 -1297 -205
rect -1373 -237 -1297 -221
rect -1195 -221 -1179 -205
rect -1135 -205 -1097 -187
rect -1039 -187 -919 -140
rect -1039 -205 -1001 -187
rect -1135 -221 -1119 -205
rect -1195 -237 -1119 -221
rect -1017 -221 -1001 -205
rect -957 -205 -919 -187
rect -861 -187 -741 -140
rect -861 -205 -823 -187
rect -957 -221 -941 -205
rect -1017 -237 -941 -221
rect -839 -221 -823 -205
rect -779 -205 -741 -187
rect -683 -187 -563 -140
rect -683 -205 -645 -187
rect -779 -221 -763 -205
rect -839 -237 -763 -221
rect -661 -221 -645 -205
rect -601 -205 -563 -187
rect -505 -187 -385 -140
rect -505 -205 -467 -187
rect -601 -221 -585 -205
rect -661 -237 -585 -221
rect -483 -221 -467 -205
rect -423 -205 -385 -187
rect -327 -187 -207 -140
rect -327 -205 -289 -187
rect -423 -221 -407 -205
rect -483 -237 -407 -221
rect -305 -221 -289 -205
rect -245 -205 -207 -187
rect -149 -187 -29 -140
rect -149 -205 -111 -187
rect -245 -221 -229 -205
rect -305 -237 -229 -221
rect -127 -221 -111 -205
rect -67 -205 -29 -187
rect 29 -187 149 -140
rect 29 -205 67 -187
rect -67 -221 -51 -205
rect -127 -237 -51 -221
rect 51 -221 67 -205
rect 111 -205 149 -187
rect 207 -187 327 -140
rect 207 -205 245 -187
rect 111 -221 127 -205
rect 51 -237 127 -221
rect 229 -221 245 -205
rect 289 -205 327 -187
rect 385 -187 505 -140
rect 385 -205 423 -187
rect 289 -221 305 -205
rect 229 -237 305 -221
rect 407 -221 423 -205
rect 467 -205 505 -187
rect 563 -187 683 -140
rect 563 -205 601 -187
rect 467 -221 483 -205
rect 407 -237 483 -221
rect 585 -221 601 -205
rect 645 -205 683 -187
rect 741 -187 861 -140
rect 741 -205 779 -187
rect 645 -221 661 -205
rect 585 -237 661 -221
rect 763 -221 779 -205
rect 823 -205 861 -187
rect 919 -187 1039 -140
rect 919 -205 957 -187
rect 823 -221 839 -205
rect 763 -237 839 -221
rect 941 -221 957 -205
rect 1001 -205 1039 -187
rect 1097 -187 1217 -140
rect 1097 -205 1135 -187
rect 1001 -221 1017 -205
rect 941 -237 1017 -221
rect 1119 -221 1135 -205
rect 1179 -205 1217 -187
rect 1275 -187 1395 -140
rect 1275 -205 1313 -187
rect 1179 -221 1195 -205
rect 1119 -237 1195 -221
rect 1297 -221 1313 -205
rect 1357 -205 1395 -187
rect 1357 -221 1373 -205
rect 1297 -237 1373 -221
<< polycont >>
rect -1357 187 -1313 221
rect -1179 187 -1135 221
rect -1001 187 -957 221
rect -823 187 -779 221
rect -645 187 -601 221
rect -467 187 -423 221
rect -289 187 -245 221
rect -111 187 -67 221
rect 67 187 111 221
rect 245 187 289 221
rect 423 187 467 221
rect 601 187 645 221
rect 779 187 823 221
rect 957 187 1001 221
rect 1135 187 1179 221
rect 1313 187 1357 221
rect -1357 -221 -1313 -187
rect -1179 -221 -1135 -187
rect -1001 -221 -957 -187
rect -823 -221 -779 -187
rect -645 -221 -601 -187
rect -467 -221 -423 -187
rect -289 -221 -245 -187
rect -111 -221 -67 -187
rect 67 -221 111 -187
rect 245 -221 289 -187
rect 423 -221 467 -187
rect 601 -221 645 -187
rect 779 -221 823 -187
rect 957 -221 1001 -187
rect 1135 -221 1179 -187
rect 1313 -221 1357 -187
<< locali >>
rect -1373 187 -1357 221
rect -1313 187 -1297 221
rect -1195 187 -1179 221
rect -1135 187 -1119 221
rect -1017 187 -1001 221
rect -957 187 -941 221
rect -839 187 -823 221
rect -779 187 -763 221
rect -661 187 -645 221
rect -601 187 -585 221
rect -483 187 -467 221
rect -423 187 -407 221
rect -305 187 -289 221
rect -245 187 -229 221
rect -127 187 -111 221
rect -67 187 -51 221
rect 51 187 67 221
rect 111 187 127 221
rect 229 187 245 221
rect 289 187 305 221
rect 407 187 423 221
rect 467 187 483 221
rect 585 187 601 221
rect 645 187 661 221
rect 763 187 779 221
rect 823 187 839 221
rect 941 187 957 221
rect 1001 187 1017 221
rect 1119 187 1135 221
rect 1179 187 1195 221
rect 1297 187 1313 221
rect 1357 187 1373 221
rect -1441 128 -1407 144
rect -1441 -144 -1407 -128
rect -1263 128 -1229 144
rect -1263 -144 -1229 -128
rect -1085 128 -1051 144
rect -1085 -144 -1051 -128
rect -907 128 -873 144
rect -907 -144 -873 -128
rect -729 128 -695 144
rect -729 -144 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 144
rect 695 -144 729 -128
rect 873 128 907 144
rect 873 -144 907 -128
rect 1051 128 1085 144
rect 1051 -144 1085 -128
rect 1229 128 1263 144
rect 1229 -144 1263 -128
rect 1407 128 1441 144
rect 1407 -144 1441 -128
rect -1373 -221 -1357 -187
rect -1313 -221 -1297 -187
rect -1195 -221 -1179 -187
rect -1135 -221 -1119 -187
rect -1017 -221 -1001 -187
rect -957 -221 -941 -187
rect -839 -221 -823 -187
rect -779 -221 -763 -187
rect -661 -221 -645 -187
rect -601 -221 -585 -187
rect -483 -221 -467 -187
rect -423 -221 -407 -187
rect -305 -221 -289 -187
rect -245 -221 -229 -187
rect -127 -221 -111 -187
rect -67 -221 -51 -187
rect 51 -221 67 -187
rect 111 -221 127 -187
rect 229 -221 245 -187
rect 289 -221 305 -187
rect 407 -221 423 -187
rect 467 -221 483 -187
rect 585 -221 601 -187
rect 645 -221 661 -187
rect 763 -221 779 -187
rect 823 -221 839 -187
rect 941 -221 957 -187
rect 1001 -221 1017 -187
rect 1119 -221 1135 -187
rect 1179 -221 1195 -187
rect 1297 -221 1313 -187
rect 1357 -221 1373 -187
<< viali >>
rect -1357 187 -1313 221
rect -1179 187 -1135 221
rect -1001 187 -957 221
rect -823 187 -779 221
rect -645 187 -601 221
rect -467 187 -423 221
rect -289 187 -245 221
rect -111 187 -67 221
rect 67 187 111 221
rect 245 187 289 221
rect 423 187 467 221
rect 601 187 645 221
rect 779 187 823 221
rect 957 187 1001 221
rect 1135 187 1179 221
rect 1313 187 1357 221
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
rect -1357 -221 -1313 -187
rect -1179 -221 -1135 -187
rect -1001 -221 -957 -187
rect -823 -221 -779 -187
rect -645 -221 -601 -187
rect -467 -221 -423 -187
rect -289 -221 -245 -187
rect -111 -221 -67 -187
rect 67 -221 111 -187
rect 245 -221 289 -187
rect 423 -221 467 -187
rect 601 -221 645 -187
rect 779 -221 823 -187
rect 957 -221 1001 -187
rect 1135 -221 1179 -187
rect 1313 -221 1357 -187
<< metal1 >>
rect -1373 221 -1297 237
rect -1373 187 -1357 221
rect -1313 187 -1297 221
rect -1373 181 -1297 187
rect -1195 221 -1119 237
rect -1195 187 -1179 221
rect -1135 187 -1119 221
rect -1195 181 -1119 187
rect -1017 221 -941 237
rect -1017 187 -1001 221
rect -957 187 -941 221
rect -1017 181 -941 187
rect -839 221 -763 237
rect -839 187 -823 221
rect -779 187 -763 221
rect -839 181 -763 187
rect -661 221 -585 237
rect -661 187 -645 221
rect -601 187 -585 221
rect -661 181 -585 187
rect -483 221 -407 237
rect -483 187 -467 221
rect -423 187 -407 221
rect -483 181 -407 187
rect -305 221 -229 237
rect -305 187 -289 221
rect -245 187 -229 221
rect -305 181 -229 187
rect -127 221 -51 237
rect -127 187 -111 221
rect -67 187 -51 221
rect -127 181 -51 187
rect 51 221 127 237
rect 51 187 67 221
rect 111 187 127 221
rect 51 181 127 187
rect 229 221 305 237
rect 229 187 245 221
rect 289 187 305 221
rect 229 181 305 187
rect 407 221 483 237
rect 407 187 423 221
rect 467 187 483 221
rect 407 181 483 187
rect 585 221 661 237
rect 585 187 601 221
rect 645 187 661 221
rect 585 181 661 187
rect 763 221 839 237
rect 763 187 779 221
rect 823 187 839 221
rect 763 181 839 187
rect 941 221 1017 237
rect 941 187 957 221
rect 1001 187 1017 221
rect 941 181 1017 187
rect 1119 221 1195 237
rect 1119 187 1135 221
rect 1179 187 1195 221
rect 1119 181 1195 187
rect 1297 221 1373 237
rect 1297 187 1313 221
rect 1357 187 1373 221
rect 1297 181 1373 187
rect -1447 128 -1401 140
rect -1447 -128 -1441 128
rect -1407 -128 -1401 128
rect -1447 -140 -1401 -128
rect -1269 128 -1223 140
rect -1269 -128 -1263 128
rect -1229 -128 -1223 128
rect -1269 -140 -1223 -128
rect -1091 128 -1045 140
rect -1091 -128 -1085 128
rect -1051 -128 -1045 128
rect -1091 -140 -1045 -128
rect -913 128 -867 140
rect -913 -128 -907 128
rect -873 -128 -867 128
rect -913 -140 -867 -128
rect -735 128 -689 140
rect -735 -128 -729 128
rect -695 -128 -689 128
rect -735 -140 -689 -128
rect -557 128 -511 140
rect -557 -128 -551 128
rect -517 -128 -511 128
rect -557 -140 -511 -128
rect -379 128 -333 140
rect -379 -128 -373 128
rect -339 -128 -333 128
rect -379 -140 -333 -128
rect -201 128 -155 140
rect -201 -128 -195 128
rect -161 -128 -155 128
rect -201 -140 -155 -128
rect -23 128 23 140
rect -23 -128 -17 128
rect 17 -128 23 128
rect -23 -140 23 -128
rect 155 128 201 140
rect 155 -128 161 128
rect 195 -128 201 128
rect 155 -140 201 -128
rect 333 128 379 140
rect 333 -128 339 128
rect 373 -128 379 128
rect 333 -140 379 -128
rect 511 128 557 140
rect 511 -128 517 128
rect 551 -128 557 128
rect 511 -140 557 -128
rect 689 128 735 140
rect 689 -128 695 128
rect 729 -128 735 128
rect 689 -140 735 -128
rect 867 128 913 140
rect 867 -128 873 128
rect 907 -128 913 128
rect 867 -140 913 -128
rect 1045 128 1091 140
rect 1045 -128 1051 128
rect 1085 -128 1091 128
rect 1045 -140 1091 -128
rect 1223 128 1269 140
rect 1223 -128 1229 128
rect 1263 -128 1269 128
rect 1223 -140 1269 -128
rect 1401 128 1447 140
rect 1401 -128 1407 128
rect 1441 -128 1447 128
rect 1401 -140 1447 -128
rect -1373 -187 -1297 -181
rect -1373 -221 -1357 -187
rect -1313 -221 -1297 -187
rect -1373 -237 -1297 -221
rect -1195 -187 -1119 -181
rect -1195 -221 -1179 -187
rect -1135 -221 -1119 -187
rect -1195 -237 -1119 -221
rect -1017 -187 -941 -181
rect -1017 -221 -1001 -187
rect -957 -221 -941 -187
rect -1017 -237 -941 -221
rect -839 -187 -763 -181
rect -839 -221 -823 -187
rect -779 -221 -763 -187
rect -839 -237 -763 -221
rect -661 -187 -585 -181
rect -661 -221 -645 -187
rect -601 -221 -585 -187
rect -661 -237 -585 -221
rect -483 -187 -407 -181
rect -483 -221 -467 -187
rect -423 -221 -407 -187
rect -483 -237 -407 -221
rect -305 -187 -229 -181
rect -305 -221 -289 -187
rect -245 -221 -229 -187
rect -305 -237 -229 -221
rect -127 -187 -51 -181
rect -127 -221 -111 -187
rect -67 -221 -51 -187
rect -127 -237 -51 -221
rect 51 -187 127 -181
rect 51 -221 67 -187
rect 111 -221 127 -187
rect 51 -237 127 -221
rect 229 -187 305 -181
rect 229 -221 245 -187
rect 289 -221 305 -187
rect 229 -237 305 -221
rect 407 -187 483 -181
rect 407 -221 423 -187
rect 467 -221 483 -187
rect 407 -237 483 -221
rect 585 -187 661 -181
rect 585 -221 601 -187
rect 645 -221 661 -187
rect 585 -237 661 -221
rect 763 -187 839 -181
rect 763 -221 779 -187
rect 823 -221 839 -187
rect 763 -237 839 -221
rect 941 -187 1017 -181
rect 941 -221 957 -187
rect 1001 -221 1017 -187
rect 941 -237 1017 -221
rect 1119 -187 1195 -181
rect 1119 -221 1135 -187
rect 1179 -221 1195 -187
rect 1119 -237 1195 -221
rect 1297 -187 1373 -181
rect 1297 -221 1313 -187
rect 1357 -221 1373 -187
rect 1297 -237 1373 -221
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 16 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
