* NGSPICE file created from comparator_v2.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_VCQUSW a_n810_n632# a_1802_n632# a_n4080_n100# a_2640_n100#
+ a_2010_n100# a_3852_131# a_n3750_n632# a_n3120_n632# a_3600_n632# a_2594_n401# a_n88_n632#
+ a_n2866_n401# a_n2912_n100# a_n718_n632# a_n556_n729# a_2548_n100# a_n182_n100#
+ a_n3658_n632# a_n3028_n632# a_n3496_n729# a_2012_n632# a_2642_n632# a_n1140_n100#
+ a_n1770_n100# a_n1398_n197# a_2172_131# a_n812_n100# a_n4128_131# a_3224_n729# a_n766_n401#
+ a_3480_n100# a_n3122_n100# a_n3752_n100# a_240_n632# a_870_n632# a_n2448_131# a_3388_n100#
+ a_3434_n401# a_n3706_n401# a_3482_n632# a_492_131# a_1500_n632# a_4064_n729# a_n1650_n632#
+ a_n1020_n632# a_n768_131# a_n2238_n197# a_n1558_n632# a_n2610_n100# a_n1396_n729#
+ w_n4520_n851# a_750_n100# a_120_n100# a_1124_n729# a_n2490_n632# a_2340_n632# a_2970_n632#
+ a_1380_n100# a_658_n100# a_n510_n100# a_n1022_n100# a_n1652_n100# a_n138_n197# a_1288_n100#
+ a_n3450_n100# a_n3078_n197# a_n2398_n632# a_122_n632# a_752_n632# a_1334_n401# a_74_n401#
+ a_702_n197# a_1382_n632# a_n1606_n401# a_1962_n197# a_3012_131# a_n390_n632# a_1918_n100#
+ a_28_n100# a_3180_n632# a_n2492_n100# a_1332_131# a_n2236_n729# a_n298_n632# a_3810_n632#
+ a_2850_n100# a_2220_n100# a_n3960_n632# a_n3330_n632# a_2174_n401# a_n1608_131#
+ a_n928_n632# a_n2446_n401# a_n136_n729# a_n3868_n632# a_n3238_n632# a_2758_n100#
+ a_2128_n100# a_n392_n100# a_n3076_n729# a_2802_n197# a_2222_n632# a_2852_n632# a_n1350_n100#
+ a_n1980_n100# a_n4170_n632# a_4020_n632# a_n346_n401# a_3690_n100# a_3060_n100#
+ a_n3332_n100# a_n3962_n100# a_2592_131# a_450_n632# a_n3286_n401# a_3598_n100# a_n4078_n632#
+ a_1080_n632# a_3014_n401# a_n2868_131# a_3062_n632# a_3692_n632# a_n2190_n100# a_3642_n197#
+ a_n1860_n632# a_n1230_n632# a_1710_n632# a_n4172_n100# a_n2820_n100# a_n1768_n632#
+ a_n1138_n632# a_n1188_131# a_704_n729# a_n4126_n401# a_960_n100# a_330_n100# a_1964_n729#
+ a_1590_n100# a_282_n197# a_n2070_n632# a_2550_n632# a_n90_n100# a_n978_n197# a_n1186_n401#
+ a_868_n100# a_238_n100# a_n720_n100# a_n1232_n100# a_n1862_n100# a_914_n401# a_1498_n100#
+ a_n3030_n100# a_n3660_n100# a_n2700_n632# a_332_n632# a_962_n632# a_1542_n197# a_1592_n632#
+ a_n3918_n197# a_n2608_n632# a_3390_n632# a_n2072_n100# a_3432_131# a_n600_n632#
+ a_1752_131# a_2804_n729# a_n3540_n632# a_2430_n100# a_n2702_n100# a_n3708_131# a_n508_n632#
+ a_n2026_n401# a_2382_n197# a_2968_n100# a_2338_n100# a_n976_n729# a_n3448_n632#
+ a_n1560_n100# a_2432_n632# a_3644_n729# a_3270_n100# a_n602_n100# a_n2028_131# a_n3916_n729#
+ a_n3542_n100# a_660_n632# a_n1818_n197# a_3178_n100# a_1290_n632# a_3900_n100# a_3854_n401#
+ a_3222_n197# a_3272_n632# a_n348_131# a_30_n632# a_3808_n100# a_n1440_n632# a_1920_n632#
+ a_284_n729# a_n2658_n197# a_3902_n632# a_n2400_n100# a_n1978_n632# a_n1348_n632#
+ a_n3288_131# a_4110_n100# a_494_n401# a_540_n100# a_4062_n197# a_4018_n100# a_1544_n729#
+ a_n2280_n632# a_2130_n632# a_2760_n632# a_1170_n100# a_72_131# a_n300_n100# a_n930_n100#
+ a_n1442_n100# a_n558_n197# a_n1816_n729# a_448_n100# a_n3240_n100# a_n3870_n100#
+ a_n3498_n197# a_n2188_n632# a_4112_n632# a_1078_n100# a_1754_n401# a_1800_n100#
+ a_n2910_n632# a_542_n632# a_1122_n197# a_n180_n632# a_1172_n632# a_2384_n729# a_n2818_n632#
+ a_1708_n100# a_912_131# VSUBS a_n2656_n729# a_n2282_n100#
X0 a_n90_n100# a_n138_n197# a_n182_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X1 a_330_n100# a_282_n197# a_238_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2 a_n3868_n632# a_n3916_n729# a_n3960_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X3 a_n1348_n632# a_n1396_n729# a_n1440_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X4 a_n3450_n100# a_n3498_n197# a_n3542_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X5 a_3480_n100# a_3432_131# a_3388_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X6 a_3062_n632# a_3014_n401# a_2970_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X7 a_542_n632# a_494_n401# a_450_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X8 a_2432_n632# a_2384_n729# a_2340_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X9 a_n1770_n100# a_n1818_n197# a_n1862_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X10 a_1800_n100# a_1752_131# a_1708_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X11 a_n508_n632# a_n556_n729# a_n600_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X12 a_1592_n632# a_1544_n729# a_1500_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X13 a_2222_n632# a_2174_n401# a_2130_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X14 a_540_n100# a_492_131# a_448_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X15 a_2220_n100# a_2172_131# a_2128_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X16 a_n3660_n100# a_n3708_131# a_n3752_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X17 a_n300_n100# a_n348_131# a_n392_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X18 a_3690_n100# a_3642_n197# a_3598_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X19 a_n3028_n632# a_n3076_n729# a_n3120_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X20 a_n2398_n632# a_n2446_n401# a_n2490_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X21 a_4110_n100# a_4062_n197# a_4018_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X22 a_n1558_n632# a_n1606_n401# a_n1650_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X23 a_n1980_n100# a_n2028_131# a_n2072_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X24 a_2010_n100# a_1962_n197# a_1918_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X25 a_3272_n632# a_3224_n729# a_3180_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X26 a_n510_n100# a_n558_n197# a_n602_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X27 a_750_n100# a_702_n197# a_658_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X28 a_752_n632# a_704_n729# a_660_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X29 a_2642_n632# a_2594_n401# a_2550_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X30 a_n3870_n100# a_n3918_n197# a_n3962_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X31 a_3900_n100# a_3852_131# a_3808_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X32 a_n4078_n632# a_n4126_n401# a_n4170_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X33 a_n718_n632# a_n766_n401# a_n810_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X34 a_1802_n632# a_1754_n401# a_1710_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X35 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=2.48e+12p pd=2.096e+07u as=0p ps=0u w=1e+06u l=150000u
X36 a_n3238_n632# a_n3286_n401# a_n3330_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X37 a_n2608_n632# a_n2656_n729# a_n2700_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X38 a_n2190_n100# a_n2238_n197# a_n2282_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X39 a_n720_n100# a_n768_131# a_n812_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X40 a_960_n100# a_912_131# a_868_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X41 a_n1768_n632# a_n1816_n729# a_n1860_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X42 a_4112_n632# a_4064_n729# a_4020_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X43 a_n4080_n100# a_n4128_131# a_n4172_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X44 a_2852_n632# a_2804_n729# a_2760_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X45 a_3482_n632# a_3434_n401# a_3390_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X46 a_962_n632# a_914_n401# a_870_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X47 a_n2400_n100# a_n2448_131# a_n2492_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X48 a_2430_n100# a_2382_n197# a_2338_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X49 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n928_n632# a_n976_n729# a_n1020_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X51 a_122_n632# a_74_n401# a_30_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X52 a_2012_n632# a_1964_n729# a_1920_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X53 a_n3448_n632# a_n3496_n729# a_n3540_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X54 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_n930_n100# a_n978_n197# a_n1022_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X56 a_n2818_n632# a_n2866_n401# a_n2910_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X57 a_n1140_n100# a_n1188_131# a_n1232_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X58 a_1170_n100# a_1122_n197# a_1078_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X59 a_n88_n632# a_n136_n729# a_n180_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X60 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_n2610_n100# a_n2658_n197# a_n2702_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X62 a_2640_n100# a_2592_131# a_2548_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X63 a_1172_n632# a_1124_n729# a_1080_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X64 a_3692_n632# a_3644_n729# a_3600_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X65 a_n3030_n100# a_n3078_n197# a_n3122_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X66 a_3060_n100# a_3012_131# a_2968_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X67 a_n1978_n632# a_n2026_n401# a_n2070_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X68 a_n3658_n632# a_n3706_n401# a_n3750_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X69 a_n1138_n632# a_n1186_n401# a_n1230_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X70 a_n1350_n100# a_n1398_n197# a_n1442_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X71 a_1380_n100# a_1332_131# a_1288_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X72 a_n2820_n100# a_n2868_131# a_n2912_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X73 a_2850_n100# a_2802_n197# a_2758_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X74 a_332_n632# a_284_n729# a_240_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X75 a_n3240_n100# a_n3288_131# a_n3332_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X76 a_3270_n100# a_3222_n197# a_3178_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X77 a_n298_n632# a_n346_n401# a_n390_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X78 a_1382_n632# a_1334_n401# a_1290_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X79 a_3902_n632# a_3854_n401# a_3810_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X80 a_n1560_n100# a_n1608_131# a_n1652_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X81 a_120_n100# a_72_131# a_28_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X82 a_1590_n100# a_1542_n197# a_1498_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X83 a_n2188_n632# a_n2236_n729# a_n2280_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
C0 w_n4520_n851# a_3642_n197# 0.09fF
C1 a_n508_n632# a_n1020_n632# 0.01fF
C2 a_n180_n632# a_n1348_n632# 0.01fF
C3 a_n390_n632# a_n1138_n632# 0.01fF
C4 a_n88_n632# a_n1440_n632# 0.00fF
C5 a_n600_n632# a_n928_n632# 0.02fF
C6 a_n298_n632# a_n1230_n632# 0.01fF
C7 a_240_n632# a_n508_n632# 0.01fF
C8 a_n182_n100# a_540_n100# 0.01fF
C9 a_3692_n632# a_3644_n729# 0.00fF
C10 a_3224_n729# a_3270_n100# 0.00fF
C11 a_n2072_n100# w_n4520_n851# 0.02fF
C12 a_n2448_131# a_n1398_n197# 0.00fF
C13 a_n810_n632# w_n4520_n851# 0.01fF
C14 a_n4078_n632# a_n3960_n632# 0.07fF
C15 a_n4170_n632# a_n3868_n632# 0.02fF
C16 a_1710_n632# w_n4520_n851# 0.01fF
C17 a_2970_n632# a_3692_n632# 0.01fF
C18 a_2852_n632# a_3810_n632# 0.01fF
C19 a_2760_n632# a_3902_n632# 0.01fF
C20 a_n2282_n100# a_n1442_n100# 0.01fF
C21 a_n2400_n100# a_n1350_n100# 0.01fF
C22 a_n2190_n100# a_n2236_n729# 0.00fF
C23 a_n4128_131# a_n4170_n632# 0.00fF
C24 a_n558_n197# a_n602_n100# 0.00fF
C25 a_n1768_n632# a_n1440_n632# 0.02fF
C26 a_n1650_n632# a_n1558_n632# 0.09fF
C27 a_492_131# a_448_n100# 0.00fF
C28 a_3060_n100# w_n4520_n851# 0.03fF
C29 a_n1980_n100# a_n3450_n100# 0.00fF
C30 a_870_n632# a_n600_n632# 0.00fF
C31 a_n2070_n632# a_n1020_n632# 0.01fF
C32 a_n1860_n632# a_n1230_n632# 0.01fF
C33 a_n1818_n197# a_n3078_n197# 0.00fF
C34 a_n2188_n632# a_n928_n632# 0.00fF
C35 a_n1978_n632# a_n1138_n632# 0.01fF
C36 a_870_n632# a_1920_n632# 0.01fF
C37 a_4020_n632# a_3062_n632# 0.01fF
C38 a_n1818_n197# a_n768_131# 0.00fF
C39 a_2430_n100# a_2548_n100# 0.07fF
C40 a_2338_n100# a_2640_n100# 0.02fF
C41 a_120_n100# a_n1442_n100# 0.00fF
C42 a_n346_n401# a_n1186_n401# 0.01fF
C43 a_n1442_n100# a_n720_n100# 0.01fF
C44 a_n1140_n100# a_n1022_n100# 0.07fF
C45 a_n1232_n100# a_n930_n100# 0.02fF
C46 a_n1350_n100# a_n812_n100# 0.01fF
C47 a_1708_n100# a_868_n100# 0.01fF
C48 a_3222_n197# a_1752_131# 0.00fF
C49 a_4020_n632# a_4064_n729# 0.00fF
C50 w_n4520_n851# a_n2398_n632# 0.01fF
C51 w_n4520_n851# a_2432_n632# 0.01fF
C52 a_3224_n729# a_3854_n401# 0.00fF
C53 a_332_n632# a_n718_n632# 0.01fF
C54 a_3644_n729# a_3434_n401# 0.00fF
C55 a_n1186_n401# a_n766_n401# 0.01fF
C56 a_332_n632# a_1802_n632# 0.00fF
C57 a_n392_n100# a_658_n100# 0.01fF
C58 a_1918_n100# a_2128_n100# 0.03fF
C59 a_1800_n100# a_2220_n100# 0.02fF
C60 a_3012_131# a_2382_n197# 0.00fF
C61 a_2220_n100# a_3388_n100# 0.01fF
C62 a_2128_n100# a_3480_n100# 0.00fF
C63 a_2010_n100# a_3598_n100# 0.00fF
C64 a_n3330_n632# a_n2398_n632# 0.01fF
C65 a_n3448_n632# a_n2280_n632# 0.01fF
C66 a_n3658_n632# a_n2070_n632# 0.00fF
C67 a_448_n100# a_n1022_n100# 0.00fF
C68 a_n3028_n632# a_n2700_n632# 0.02fF
C69 a_3480_n100# a_3690_n100# 0.03fF
C70 a_3388_n100# a_3808_n100# 0.02fF
C71 a_3270_n100# a_3900_n100# 0.01fF
C72 a_n3120_n632# a_n2608_n632# 0.01fF
C73 a_n3540_n632# a_n2188_n632# 0.00fF
C74 a_n3238_n632# a_n2490_n632# 0.01fF
C75 a_1122_n197# a_1078_n100# 0.00fF
C76 a_2172_131# a_1752_131# 0.01fF
C77 a_2592_131# a_1332_131# 0.00fF
C78 a_n2190_n100# a_n1560_n100# 0.01fF
C79 a_n2072_n100# a_n1652_n100# 0.02fF
C80 a_n1980_n100# a_n1770_n100# 0.03fF
C81 a_4112_n632# a_2970_n632# 0.01fF
C82 a_n3708_131# a_n3498_n197# 0.00fF
C83 a_1754_n401# a_2384_n729# 0.00fF
C84 a_2594_n401# a_1544_n729# 0.00fF
C85 a_2174_n401# a_1964_n729# 0.00fF
C86 a_n348_131# a_n1398_n197# 0.00fF
C87 a_238_n100# w_n4520_n851# 0.02fF
C88 a_3432_131# a_4062_n197# 0.00fF
C89 a_n810_n632# a_n390_n632# 0.02fF
C90 a_n718_n632# a_n508_n632# 0.03fF
C91 a_1382_n632# a_n88_n632# 0.00fF
C92 a_1802_n632# a_2012_n632# 0.03fF
C93 a_n1980_n100# a_n510_n100# 0.00fF
C94 a_n1560_n100# a_n602_n100# 0.01fF
C95 a_1172_n632# a_1500_n632# 0.02fF
C96 a_n2820_n100# a_n2492_n100# 0.02fF
C97 a_n2702_n100# a_n2610_n100# 0.09fF
C98 a_962_n632# a_1710_n632# 0.01fF
C99 a_238_n100# a_330_n100# 0.09fF
C100 a_960_n100# a_1170_n100# 0.03fF
C101 a_1918_n100# w_n4520_n851# 0.02fF
C102 a_2338_n100# a_1170_n100# 0.01fF
C103 a_2430_n100# a_1078_n100# 0.00fF
C104 w_n4520_n851# a_3480_n100# 0.04fF
C105 a_1500_n632# a_3062_n632# 0.00fF
C106 a_n3030_n100# a_n3870_n100# 0.01fF
C107 a_n3122_n100# a_n3752_n100# 0.01fF
C108 a_n2702_n100# a_n4172_n100# 0.00fF
C109 a_n3240_n100# a_n3660_n100# 0.02fF
C110 a_n3332_n100# a_n3542_n100# 0.03fF
C111 a_n2912_n100# a_n3962_n100# 0.01fF
C112 a_n2820_n100# a_n4080_n100# 0.00fF
C113 a_3644_n729# a_2384_n729# 0.00fF
C114 a_1918_n100# a_330_n100# 0.00fF
C115 a_1498_n100# a_960_n100# 0.01fF
C116 a_1498_n100# a_2338_n100# 0.01fF
C117 a_1380_n100# a_2430_n100# 0.01fF
C118 a_n4128_131# a_n3288_131# 0.01fF
C119 w_n4520_n851# a_n928_n632# 0.01fF
C120 a_450_n632# a_1592_n632# 0.01fF
C121 a_n2238_n197# a_n1818_n197# 0.01fF
C122 a_3900_n100# a_3854_n401# 0.00fF
C123 a_448_n100# a_1078_n100# 0.01fF
C124 a_540_n100# a_960_n100# 0.02fF
C125 a_n182_n100# a_120_n100# 0.02fF
C126 a_658_n100# a_868_n100# 0.03fF
C127 a_n300_n100# a_n602_n100# 0.02fF
C128 a_n182_n100# a_n720_n100# 0.01fF
C129 a_n90_n100# a_n812_n100# 0.01fF
C130 a_n3868_n632# a_n2818_n632# 0.01fF
C131 a_n3750_n632# a_n2910_n632# 0.01fF
C132 a_2174_n401# a_2222_n632# 0.00fF
C133 a_2172_131# a_702_n197# 0.00fF
C134 a_n2910_n632# a_n1348_n632# 0.00fF
C135 a_n2818_n632# a_n1440_n632# 0.00fF
C136 a_n2868_131# a_n2866_n401# 0.01fF
C137 a_n810_n632# a_n1978_n632# 0.01fF
C138 a_n718_n632# a_n2070_n632# 0.00fF
C139 a_n600_n632# a_n2188_n632# 0.00fF
C140 a_1380_n100# a_448_n100# 0.01fF
C141 a_282_n197# a_1122_n197# 0.01fF
C142 a_1802_n632# a_2760_n632# 0.01fF
C143 a_1710_n632# a_2852_n632# 0.01fF
C144 a_2012_n632# a_2550_n632# 0.01fF
C145 a_1592_n632# a_2970_n632# 0.00fF
C146 a_1920_n632# a_2642_n632# 0.01fF
C147 a_122_n632# a_n88_n632# 0.03fF
C148 a_962_n632# a_2432_n632# 0.00fF
C149 a_1172_n632# a_2222_n632# 0.01fF
C150 a_n2868_131# a_n2658_n197# 0.00fF
C151 a_704_n729# a_1544_n729# 0.01fF
C152 a_2222_n632# a_3062_n632# 0.01fF
C153 a_2130_n632# a_3180_n632# 0.01fF
C154 a_n2190_n100# a_n3030_n100# 0.01fF
C155 a_n1862_n100# a_n3332_n100# 0.00fF
C156 a_n2072_n100# a_n3122_n100# 0.01fF
C157 a_n2400_n100# a_n2820_n100# 0.02fF
C158 a_n1980_n100# a_n3240_n100# 0.00fF
C159 a_n2282_n100# a_n2912_n100# 0.01fF
C160 w_n4520_n851# a_914_n401# 0.10fF
C161 a_2968_n100# a_2970_n632# 0.00fF
C162 w_n4520_n851# a_n3540_n632# 0.03fF
C163 w_n4520_n851# a_n3496_n729# 0.12fF
C164 a_n3540_n632# a_n3330_n632# 0.03fF
C165 a_n3658_n632# a_n3238_n632# 0.02fF
C166 a_n4170_n632# a_n2700_n632# 0.00fF
C167 a_1080_n632# a_1500_n632# 0.02fF
C168 a_870_n632# w_n4520_n851# 0.01fF
C169 a_n2700_n632# a_n1768_n632# 0.01fF
C170 w_n4520_n851# a_n4126_n401# 0.12fF
C171 a_1800_n100# a_1752_131# 0.00fF
C172 w_n4520_n851# a_n3542_n100# 0.04fF
C173 a_1962_n197# a_492_131# 0.00fF
C174 a_1800_n100# a_1754_n401# 0.00fF
C175 a_n2492_n100# a_n1140_n100# 0.00fF
C176 a_n2610_n100# a_n1022_n100# 0.00fF
C177 a_n3448_n632# a_n3450_n100# 0.00fF
C178 a_n2490_n632# a_n1860_n632# 0.01fF
C179 a_n2398_n632# a_n1978_n632# 0.02fF
C180 a_1122_n197# a_2382_n197# 0.00fF
C181 a_1542_n197# a_1962_n197# 0.01fF
C182 a_n2280_n632# a_n2070_n632# 0.03fF
C183 a_n3496_n729# a_n2656_n729# 0.01fF
C184 a_2550_n632# a_2760_n632# 0.03fF
C185 a_752_n632# a_n180_n632# 0.01fF
C186 a_2432_n632# a_2852_n632# 0.02fF
C187 a_2340_n632# a_2970_n632# 0.01fF
C188 a_n3286_n401# a_n3496_n729# 0.00fF
C189 a_2010_n100# a_2012_n632# 0.00fF
C190 a_n2866_n401# a_n3916_n729# 0.00fF
C191 a_n3706_n401# a_n3076_n729# 0.00fF
C192 a_n4126_n401# a_n2656_n729# 0.00fF
C193 a_752_n632# a_1172_n632# 0.02fF
C194 a_n90_n100# a_1288_n100# 0.00fF
C195 a_542_n632# a_1382_n632# 0.01fF
C196 a_n392_n100# a_238_n100# 0.01fF
C197 a_n4126_n401# a_n3286_n401# 0.01fF
C198 a_28_n100# a_n1022_n100# 0.01fF
C199 a_3272_n632# a_3600_n632# 0.02fF
C200 a_3180_n632# a_3692_n632# 0.01fF
C201 a_3390_n632# a_3482_n632# 0.09fF
C202 a_3062_n632# a_3810_n632# 0.01fF
C203 a_2220_n100# a_3178_n100# 0.01fF
C204 a_2128_n100# a_750_n100# 0.00fF
C205 a_3178_n100# a_3808_n100# 0.01fF
C206 a_3060_n100# a_3900_n100# 0.01fF
C207 a_2968_n100# a_4018_n100# 0.01fF
C208 a_2850_n100# a_4110_n100# 0.00fF
C209 a_240_n632# a_284_n729# 0.00fF
C210 a_n88_n632# a_n1230_n632# 0.01fF
C211 a_n390_n632# a_n928_n632# 0.01fF
C212 a_n298_n632# a_n1020_n632# 0.01fF
C213 a_n180_n632# a_n1138_n632# 0.01fF
C214 a_240_n632# a_n298_n632# 0.01fF
C215 a_n3288_131# a_n3708_131# 0.01fF
C216 a_1080_n632# a_2222_n632# 0.01fF
C217 a_n1608_131# a_n978_n197# 0.00fF
C218 a_n978_n197# a_n976_n729# 0.01fF
C219 a_n1862_n100# w_n4520_n851# 0.02fF
C220 a_2430_n100# a_2382_n197# 0.00fF
C221 a_n1608_131# w_n4520_n851# 0.12fF
C222 w_n4520_n851# a_n976_n729# 0.12fF
C223 a_n600_n632# w_n4520_n851# 0.01fF
C224 a_914_n401# a_1334_n401# 0.01fF
C225 a_n4078_n632# a_n3750_n632# 0.02fF
C226 a_n3960_n632# a_n3868_n632# 0.09fF
C227 a_1920_n632# w_n4520_n851# 0.01fF
C228 a_2970_n632# a_3902_n632# 0.01fF
C229 a_914_n401# a_n136_n729# 0.00fF
C230 a_n346_n401# a_1124_n729# 0.00fF
C231 a_542_n632# a_2130_n632# 0.00fF
C232 a_n2072_n100# a_n1442_n100# 0.01fF
C233 a_n2190_n100# a_n1350_n100# 0.01fF
C234 a_n2282_n100# a_n1232_n100# 0.01fF
C235 a_n2400_n100# a_n1140_n100# 0.00fF
C236 a_450_n632# a_n1020_n632# 0.00fF
C237 a_n1558_n632# a_n1440_n632# 0.07fF
C238 a_n1650_n632# a_n1348_n632# 0.02fF
C239 a_n1768_n632# a_n1230_n632# 0.01fF
C240 a_240_n632# a_450_n632# 0.03fF
C241 a_122_n632# a_542_n632# 0.02fF
C242 a_2594_n401# a_3434_n401# 0.01fF
C243 a_962_n632# a_914_n401# 0.00fF
C244 w_n4520_n851# a_750_n100# 0.02fF
C245 a_1122_n197# a_912_131# 0.00fF
C246 a_n2072_n100# a_n2028_131# 0.00fF
C247 a_870_n632# a_n390_n632# 0.00fF
C248 a_n1978_n632# a_n928_n632# 0.01fF
C249 a_n1860_n632# a_n1020_n632# 0.01fF
C250 a_n346_n401# a_74_n401# 0.01fF
C251 a_4112_n632# a_3180_n632# 0.01fF
C252 a_4020_n632# a_3272_n632# 0.01fF
C253 a_330_n100# a_750_n100# 0.02fF
C254 a_238_n100# a_868_n100# 0.01fF
C255 a_120_n100# a_960_n100# 0.01fF
C256 a_28_n100# a_1078_n100# 0.01fF
C257 a_752_n632# a_1080_n632# 0.02fF
C258 a_870_n632# a_962_n632# 0.09fF
C259 a_2548_n100# a_2640_n100# 0.09fF
C260 a_2430_n100# a_2758_n100# 0.02fF
C261 a_2338_n100# a_2850_n100# 0.01fF
C262 a_n2448_131# a_n2658_n197# 0.00fF
C263 a_120_n100# a_n1232_n100# 0.00fF
C264 a_74_n401# a_n766_n401# 0.01fF
C265 a_n1022_n100# a_n930_n100# 0.09fF
C266 a_n1140_n100# a_n812_n100# 0.02fF
C267 a_n1232_n100# a_n720_n100# 0.01fF
C268 a_n1350_n100# a_n602_n100# 0.01fF
C269 a_1918_n100# a_868_n100# 0.01fF
C270 a_1380_n100# a_28_n100# 0.00fF
C271 w_n4520_n851# a_n2188_n632# 0.01fF
C272 a_30_n632# a_n1440_n632# 0.00fF
C273 w_n4520_n851# a_2642_n632# 0.02fF
C274 a_332_n632# a_n508_n632# 0.01fF
C275 a_4064_n729# a_3854_n401# 0.00fF
C276 a_2010_n100# a_2220_n100# 0.03fF
C277 a_n182_n100# a_658_n100# 0.01fF
C278 a_3012_131# a_3222_n197# 0.00fF
C279 a_2220_n100# a_3598_n100# 0.00fF
C280 a_2128_n100# a_3690_n100# 0.00fF
C281 a_n3540_n632# a_n1978_n632# 0.00fF
C282 a_n3330_n632# a_n2188_n632# 0.01fF
C283 a_n3238_n632# a_n2280_n632# 0.01fF
C284 a_n3448_n632# a_n2070_n632# 0.00fF
C285 a_448_n100# a_n812_n100# 0.00fF
C286 a_3598_n100# a_3808_n100# 0.03fF
C287 a_3480_n100# a_3900_n100# 0.02fF
C288 a_3388_n100# a_4018_n100# 0.01fF
C289 a_3270_n100# a_4110_n100# 0.01fF
C290 a_n2818_n632# a_n2700_n632# 0.07fF
C291 a_n3120_n632# a_n2398_n632# 0.01fF
C292 a_n2910_n632# a_n2608_n632# 0.02fF
C293 a_n3028_n632# a_n2490_n632# 0.01fF
C294 a_n1188_131# a_n1140_n100# 0.00fF
C295 a_n1980_n100# a_n1560_n100# 0.02fF
C296 a_n1862_n100# a_n1652_n100# 0.03fF
C297 a_n1186_n401# a_n1188_131# 0.01fF
C298 a_n4128_131# a_n4172_n100# 0.00fF
C299 a_n1652_n100# a_n1608_131# 0.00fF
C300 a_n2280_n632# a_n2236_n729# 0.00fF
C301 a_3012_131# a_2172_131# 0.01fF
C302 a_3014_n401# a_1964_n729# 0.00fF
C303 a_2594_n401# a_2384_n729# 0.00fF
C304 a_n2446_n401# a_n2398_n632# 0.00fF
C305 a_n3332_n100# w_n4520_n851# 0.03fF
C306 a_1498_n100# a_1542_n197# 0.00fF
C307 a_3222_n197# a_3180_n632# 0.00fF
C308 a_n348_131# a_n558_n197# 0.00fF
C309 a_n976_n729# a_n136_n729# 0.01fF
C310 a_492_131# a_540_n100# 0.00fF
C311 a_1802_n632# a_1754_n401# 0.00fF
C312 w_n4520_n851# a_n3918_n197# 0.11fF
C313 a_n508_n632# a_n556_n729# 0.00fF
C314 a_n3332_n100# a_n3330_n632# 0.00fF
C315 a_n810_n632# a_n180_n632# 0.01fF
C316 a_n718_n632# a_n298_n632# 0.02fF
C317 a_n600_n632# a_n390_n632# 0.03fF
C318 a_n1862_n100# a_n392_n100# 0.00fF
C319 a_2968_n100# a_3012_131# 0.00fF
C320 a_n1770_n100# a_n510_n100# 0.00fF
C321 a_962_n632# a_n600_n632# 0.00fF
C322 a_n2610_n100# a_n2492_n100# 0.07fF
C323 a_962_n632# a_1920_n632# 0.01fF
C324 a_1172_n632# a_1710_n632# 0.01fF
C325 a_2128_n100# w_n4520_n851# 0.02fF
C326 a_2430_n100# a_1288_n100# 0.01fF
C327 a_2548_n100# a_1170_n100# 0.00fF
C328 a_2640_n100# a_1078_n100# 0.00fF
C329 w_n4520_n851# a_3690_n100# 0.04fF
C330 a_1710_n632# a_3062_n632# 0.00fF
C331 a_1592_n632# a_3180_n632# 0.00fF
C332 a_4020_n632# a_4062_n197# 0.00fF
C333 a_n510_n100# a_n556_n729# 0.00fF
C334 a_n348_131# a_72_131# 0.01fF
C335 a_n3122_n100# a_n3542_n100# 0.02fF
C336 a_n3030_n100# a_n3660_n100# 0.01fF
C337 a_n768_131# a_n720_n100# 0.00fF
C338 a_n2610_n100# a_n4080_n100# 0.00fF
C339 a_n2912_n100# a_n3752_n100# 0.01fF
C340 a_n2820_n100# a_n3870_n100# 0.01fF
C341 a_n3240_n100# a_n3450_n100# 0.03fF
C342 a_n2702_n100# a_n3962_n100# 0.00fF
C343 a_n508_n632# a_n510_n100# 0.00fF
C344 a_870_n632# a_868_n100# 0.00fF
C345 a_1708_n100# a_960_n100# 0.01fF
C346 a_n4172_n100# a_n4080_n100# 0.09fF
C347 a_3060_n100# a_3062_n632# 0.00fF
C348 a_1708_n100# a_2338_n100# 0.01fF
C349 a_1590_n100# a_2430_n100# 0.01fF
C350 a_1498_n100# a_2548_n100# 0.01fF
C351 a_1380_n100# a_2640_n100# 0.00fF
C352 a_2338_n100# a_3270_n100# 0.01fF
C353 a_450_n632# a_n718_n632# 0.01fF
C354 a_450_n632# a_1802_n632# 0.00fF
C355 a_448_n100# a_1288_n100# 0.01fF
C356 a_n1398_n197# a_n558_n197# 0.01fF
C357 a_n392_n100# a_750_n100# 0.01fF
C358 a_3432_131# a_2382_n197# 0.00fF
C359 a_n90_n100# a_n602_n100# 0.01fF
C360 a_540_n100# a_n1022_n100# 0.00fF
C361 a_2592_131# a_1752_131# 0.01fF
C362 a_n2818_n632# a_n1230_n632# 0.00fF
C363 w_n4520_n851# a_n978_n197# 0.10fF
C364 a_1590_n100# a_448_n100# 0.01fF
C365 a_n508_n632# a_n2070_n632# 0.00fF
C366 a_n718_n632# a_n1860_n632# 0.01fF
C367 a_n600_n632# a_n1978_n632# 0.00fF
C368 a_1802_n632# a_2970_n632# 0.01fF
C369 a_1920_n632# a_2852_n632# 0.01fF
C370 a_2012_n632# a_2760_n632# 0.01fF
C371 a_1172_n632# a_2432_n632# 0.00fF
C372 a_n1186_n401# a_n1230_n632# 0.00fF
C373 a_2222_n632# a_3272_n632# 0.01fF
C374 a_72_131# a_n1398_n197# 0.00fF
C375 a_2130_n632# a_3390_n632# 0.00fF
C376 a_2432_n632# a_3062_n632# 0.01fF
C377 a_2340_n632# a_3180_n632# 0.01fF
C378 a_2802_n197# a_4062_n197# 0.00fF
C379 a_n2282_n100# a_n2702_n100# 0.02fF
C380 a_n1770_n100# a_n3240_n100# 0.00fF
C381 a_n2190_n100# a_n2820_n100# 0.01fF
C382 a_n1862_n100# a_n3122_n100# 0.00fF
C383 a_n1980_n100# a_n3030_n100# 0.01fF
C384 a_n2400_n100# a_n2610_n100# 0.03fF
C385 a_n2072_n100# a_n2912_n100# 0.01fF
C386 w_n4520_n851# a_n3330_n632# 0.03fF
C387 a_330_n100# w_n4520_n851# 0.02fF
C388 a_72_131# a_1332_131# 0.00fF
C389 a_3852_131# a_4062_n197# 0.00fF
C390 a_1382_n632# a_30_n632# 0.00fF
C391 w_n4520_n851# a_n2656_n729# 0.12fF
C392 a_n2282_n100# a_n2238_n197# 0.00fF
C393 a_n3448_n632# a_n3238_n632# 0.03fF
C394 a_n3540_n632# a_n3120_n632# 0.02fF
C395 a_n4078_n632# a_n2608_n632# 0.00fF
C396 a_n3658_n632# a_n3028_n632# 0.01fF
C397 a_n3960_n632# a_n2700_n632# 0.00fF
C398 a_2760_n632# a_2804_n729# 0.00fF
C399 a_1080_n632# a_1710_n632# 0.01fF
C400 a_1078_n100# a_1170_n100# 0.09fF
C401 a_n2490_n632# a_n1768_n632# 0.01fF
C402 w_n4520_n851# a_n3286_n401# 0.10fF
C403 a_n2700_n632# a_n1558_n632# 0.01fF
C404 a_n2608_n632# a_n1650_n632# 0.01fF
C405 a_n2658_n197# a_n1398_n197# 0.00fF
C406 a_n3286_n401# a_n3330_n632# 0.00fF
C407 a_1380_n100# a_1170_n100# 0.03fF
C408 a_1498_n100# a_1078_n100# 0.02fF
C409 a_n2492_n100# a_n930_n100# 0.00fF
C410 a_1962_n197# a_2382_n197# 0.01fF
C411 a_n2188_n632# a_n1978_n632# 0.03fF
C412 a_n2280_n632# a_n1860_n632# 0.02fF
C413 a_1542_n197# a_2802_n197# 0.00fF
C414 a_n3076_n729# a_n2236_n729# 0.01fF
C415 a_2550_n632# a_2970_n632# 0.02fF
C416 a_2642_n632# a_2852_n632# 0.03fF
C417 a_n2868_131# a_n3498_n197# 0.00fF
C418 a_n2866_n401# a_n3076_n729# 0.00fF
C419 a_n3706_n401# a_n2236_n729# 0.00fF
C420 a_n3286_n401# a_n2656_n729# 0.00fF
C421 a_n2446_n401# a_n3496_n729# 0.00fF
C422 a_542_n632# a_1592_n632# 0.01fF
C423 a_540_n100# a_1078_n100# 0.01fF
C424 a_n182_n100# a_238_n100# 0.02fF
C425 a_658_n100# a_960_n100# 0.02fF
C426 a_750_n100# a_868_n100# 0.07fF
C427 a_n3706_n401# a_n2866_n401# 0.01fF
C428 a_n300_n100# a_n348_131# 0.00fF
C429 a_28_n100# a_n812_n100# 0.01fF
C430 a_3180_n632# a_3902_n632# 0.01fF
C431 a_3482_n632# a_3600_n632# 0.07fF
C432 a_1380_n100# a_1498_n100# 0.07fF
C433 a_3390_n632# a_3692_n632# 0.02fF
C434 a_3272_n632# a_3810_n632# 0.01fF
C435 a_2172_131# a_1122_n197# 0.00fF
C436 a_3272_n632# a_3270_n100# 0.00fF
C437 a_3178_n100# a_4018_n100# 0.01fF
C438 a_3060_n100# a_4110_n100# 0.01fF
C439 a_1380_n100# a_540_n100# 0.01fF
C440 a_1500_n632# a_1542_n197# 0.00fF
C441 a_n180_n632# a_n928_n632# 0.01fF
C442 a_n88_n632# a_n1020_n632# 0.01fF
C443 a_122_n632# a_30_n632# 0.09fF
C444 a_240_n632# a_n88_n632# 0.02fF
C445 a_1332_131# a_1752_131# 0.01fF
C446 a_1080_n632# a_2432_n632# 0.00fF
C447 a_n1608_131# a_n138_n197# 0.00fF
C448 a_1124_n729# a_1544_n729# 0.01fF
C449 a_n558_n197# a_n556_n729# 0.01fF
C450 a_n1818_n197# a_n1188_131# 0.00fF
C451 a_n1652_n100# w_n4520_n851# 0.02fF
C452 w_n4520_n851# a_1334_n401# 0.10fF
C453 w_n4520_n851# a_n136_n729# 0.12fF
C454 a_n348_131# a_702_n197# 0.00fF
C455 a_n390_n632# w_n4520_n851# 0.01fF
C456 a_914_n401# a_2174_n401# 0.00fF
C457 a_n3868_n632# a_n3750_n632# 0.07fF
C458 a_962_n632# w_n4520_n851# 0.01fF
C459 a_1290_n632# a_1382_n632# 0.09fF
C460 a_74_n401# a_1544_n729# 0.00fF
C461 a_2430_n100# a_2384_n729# 0.00fF
C462 a_n2190_n100# a_n1140_n100# 0.01fF
C463 a_n2282_n100# a_n1022_n100# 0.00fF
C464 a_n2400_n100# a_n930_n100# 0.00fF
C465 a_n1980_n100# a_n1350_n100# 0.01fF
C466 a_n1862_n100# a_n1442_n100# 0.02fF
C467 a_n3332_n100# a_n3122_n100# 0.03fF
C468 a_n2072_n100# a_n1232_n100# 0.01fF
C469 a_n1558_n632# a_n1230_n632# 0.02fF
C470 a_n510_n100# a_n558_n197# 0.00fF
C471 a_n1768_n632# a_n1020_n632# 0.01fF
C472 a_n1440_n632# a_n1348_n632# 0.09fF
C473 a_n1650_n632# a_n1138_n632# 0.01fF
C474 a_n1980_n100# a_n2026_n401# 0.00fF
C475 a_3014_n401# a_3854_n401# 0.01fF
C476 a_n1816_n729# a_n976_n729# 0.01fF
C477 a_1962_n197# a_912_131# 0.00fF
C478 a_n392_n100# w_n4520_n851# 0.02fF
C479 a_n2446_n401# a_n976_n729# 0.00fF
C480 a_870_n632# a_n180_n632# 0.01fF
C481 a_4112_n632# a_3390_n632# 0.01fF
C482 w_n4520_n851# a_3224_n729# 0.12fF
C483 a_4020_n632# a_3482_n632# 0.01fF
C484 a_28_n100# a_1288_n100# 0.00fF
C485 a_n2028_131# a_n1608_131# 0.01fF
C486 a_2338_n100# a_3060_n100# 0.01fF
C487 a_2430_n100# a_2968_n100# 0.01fF
C488 a_2548_n100# a_2850_n100# 0.02fF
C489 a_2640_n100# a_2758_n100# 0.07fF
C490 a_660_n632# a_1382_n632# 0.01fF
C491 a_870_n632# a_1172_n632# 0.02fF
C492 a_n392_n100# a_330_n100# 0.01fF
C493 a_3390_n632# a_3434_n401# 0.00fF
C494 a_120_n100# a_n1022_n100# 0.01fF
C495 a_n2868_131# a_n2820_n100# 0.00fF
C496 a_n4170_n632# a_n3658_n632# 0.01fF
C497 a_n930_n100# a_n812_n100# 0.07fF
C498 a_n1022_n100# a_n720_n100# 0.02fF
C499 a_n1140_n100# a_n602_n100# 0.01fF
C500 a_2128_n100# a_868_n100# 0.00fF
C501 a_1590_n100# a_28_n100# 0.00fF
C502 a_332_n632# a_284_n729# 0.00fF
C503 a_n766_n401# a_n720_n100# 0.00fF
C504 a_30_n632# a_n1230_n632# 0.00fF
C505 w_n4520_n851# a_n1978_n632# 0.01fF
C506 w_n4520_n851# a_2852_n632# 0.03fF
C507 a_702_n197# a_1332_131# 0.00fF
C508 a_332_n632# a_n298_n632# 0.01fF
C509 a_1290_n632# a_2130_n632# 0.01fF
C510 a_492_131# a_494_n401# 0.01fF
C511 a_122_n632# a_1290_n632# 0.01fF
C512 a_2220_n100# a_3808_n100# 0.00fF
C513 a_448_n100# a_n602_n100# 0.01fF
C514 a_3690_n100# a_3900_n100# 0.03fF
C515 a_3598_n100# a_4018_n100# 0.02fF
C516 a_3480_n100# a_4110_n100# 0.01fF
C517 a_n3028_n632# a_n2280_n632# 0.01fF
C518 a_n2818_n632# a_n2490_n632# 0.02fF
C519 a_n2910_n632# a_n2398_n632# 0.01fF
C520 a_n3448_n632# a_n1860_n632# 0.00fF
C521 a_n3330_n632# a_n1978_n632# 0.00fF
C522 a_n3238_n632# a_n2070_n632# 0.01fF
C523 a_n3120_n632# a_n2188_n632# 0.01fF
C524 a_n1770_n100# a_n1560_n100# 0.03fF
C525 a_122_n632# a_74_n401# 0.00fF
C526 a_1334_n401# a_n136_n729# 0.00fF
C527 a_n3122_n100# w_n4520_n851# 0.03fF
C528 a_660_n632# a_2130_n632# 0.00fF
C529 a_542_n632# a_n1020_n632# 0.00fF
C530 a_n2448_131# a_n3498_n197# 0.00fF
C531 a_n556_n729# a_284_n729# 0.01fF
C532 a_240_n632# a_542_n632# 0.02fF
C533 a_332_n632# a_450_n632# 0.07fF
C534 a_122_n632# a_660_n632# 0.01fF
C535 a_3432_131# a_3434_n401# 0.01fF
C536 a_n810_n632# a_n768_131# 0.00fF
C537 a_1290_n632# a_1288_n100# 0.00fF
C538 w_n4520_n851# a_868_n100# 0.02fF
C539 a_n3240_n100# a_n3238_n632# 0.00fF
C540 a_n508_n632# a_n298_n632# 0.03fF
C541 a_n718_n632# a_n88_n632# 0.01fF
C542 a_n600_n632# a_n180_n632# 0.02fF
C543 a_n1770_n100# a_n300_n100# 0.00fF
C544 a_n1560_n100# a_n510_n100# 0.01fF
C545 a_n1652_n100# a_n392_n100# 0.00fF
C546 a_962_n632# a_n390_n632# 0.00fF
C547 a_3060_n100# a_3014_n401# 0.00fF
C548 a_1172_n632# a_1920_n632# 0.01fF
C549 a_n3030_n100# a_n3076_n729# 0.00fF
C550 a_n346_n401# a_494_n401# 0.01fF
C551 a_330_n100# a_868_n100# 0.01fF
C552 a_238_n100# a_960_n100# 0.01fF
C553 a_120_n100# a_1078_n100# 0.01fF
C554 a_2640_n100# a_1288_n100# 0.00fF
C555 a_2758_n100# a_1170_n100# 0.00fF
C556 a_870_n632# a_1080_n632# 0.03fF
C557 w_n4520_n851# a_3900_n100# 0.06fF
C558 a_n2868_131# a_n3288_131# 0.01fF
C559 a_1710_n632# a_3272_n632# 0.00fF
C560 a_1802_n632# a_3180_n632# 0.00fF
C561 a_1920_n632# a_3062_n632# 0.01fF
C562 a_n3708_131# a_n3750_n632# 0.00fF
C563 a_n2610_n100# a_n3870_n100# 0.00fF
C564 a_n2702_n100# a_n3752_n100# 0.01fF
C565 a_n2912_n100# a_n3542_n100# 0.01fF
C566 a_n2492_n100# a_n3962_n100# 0.00fF
C567 a_n2820_n100# a_n3660_n100# 0.01fF
C568 a_n3030_n100# a_n3450_n100# 0.02fF
C569 a_238_n100# a_n1232_n100# 0.00fF
C570 a_n390_n632# a_n392_n100# 0.00fF
C571 a_494_n401# a_n766_n401# 0.00fF
C572 a_1754_n401# a_2804_n729# 0.00fF
C573 a_1918_n100# a_960_n100# 0.01fF
C574 a_1918_n100# a_2338_n100# 0.02fF
C575 a_1800_n100# a_2430_n100# 0.01fF
C576 a_1708_n100# a_2548_n100# 0.01fF
C577 a_1590_n100# a_2640_n100# 0.01fF
C578 a_3178_n100# a_3180_n632# 0.00fF
C579 a_1498_n100# a_2758_n100# 0.00fF
C580 a_1380_n100# a_2850_n100# 0.00fF
C581 a_n4172_n100# a_n3870_n100# 0.02fF
C582 a_n4080_n100# a_n3962_n100# 0.07fF
C583 a_1380_n100# a_120_n100# 0.00fF
C584 a_2548_n100# a_3270_n100# 0.01fF
C585 a_2430_n100# a_3388_n100# 0.01fF
C586 a_2338_n100# a_3480_n100# 0.01fF
C587 a_450_n632# a_n508_n632# 0.01fF
C588 a_n810_n632# a_n1650_n632# 0.01fF
C589 a_n718_n632# a_n1768_n632# 0.01fF
C590 a_450_n632# a_2012_n632# 0.00fF
C591 a_n978_n197# a_n138_n197# 0.01fF
C592 a_n182_n100# a_750_n100# 0.01fF
C593 a_3432_131# a_3222_n197# 0.00fF
C594 a_n510_n100# a_n300_n100# 0.03fF
C595 a_540_n100# a_n812_n100# 0.00fF
C596 a_2594_n401# a_2550_n632# 0.00fF
C597 w_n4520_n851# a_n138_n197# 0.10fF
C598 a_n508_n632# a_n1860_n632# 0.00fF
C599 a_n390_n632# a_n1978_n632# 0.00fF
C600 a_1800_n100# a_448_n100# 0.00fF
C601 a_2012_n632# a_2970_n632# 0.01fF
C602 a_3432_131# a_2172_131# 0.00fF
C603 a_3012_131# a_2592_131# 0.01fF
C604 a_2592_131# a_2594_n401# 0.01fF
C605 a_1172_n632# a_2642_n632# 0.00fF
C606 a_2804_n729# a_3644_n729# 0.01fF
C607 a_2550_n632# a_3180_n632# 0.01fF
C608 a_2432_n632# a_3272_n632# 0.01fF
C609 a_2340_n632# a_3390_n632# 0.01fF
C610 a_2642_n632# a_3062_n632# 0.02fF
C611 a_2130_n632# a_3600_n632# 0.00fF
C612 a_2222_n632# a_3482_n632# 0.00fF
C613 a_72_131# a_n558_n197# 0.00fF
C614 a_3642_n197# a_4062_n197# 0.01fF
C615 a_n2072_n100# a_n2702_n100# 0.01fF
C616 a_n2282_n100# a_n2492_n100# 0.03fF
C617 a_n2190_n100# a_n2610_n100# 0.02fF
C618 a_n1652_n100# a_n3122_n100# 0.00fF
C619 a_n1770_n100# a_n3030_n100# 0.00fF
C620 a_n1862_n100# a_n2912_n100# 0.01fF
C621 a_n1980_n100# a_n2820_n100# 0.01fF
C622 a_n1398_n197# a_n1350_n100# 0.00fF
C623 w_n4520_n851# a_n3120_n632# 0.03fF
C624 a_n1398_n197# a_n1396_n729# 0.01fF
C625 a_n2400_n100# a_n3962_n100# 0.00fF
C626 a_1592_n632# a_30_n632# 0.00fF
C627 w_n4520_n851# a_n1442_n100# 0.02fF
C628 w_n4520_n851# a_n1816_n729# 0.12fF
C629 a_n3448_n632# a_n3028_n632# 0.02fF
C630 a_n3658_n632# a_n2818_n632# 0.01fF
C631 a_n3960_n632# a_n2490_n632# 0.00fF
C632 a_n3868_n632# a_n2608_n632# 0.00fF
C633 a_n3330_n632# a_n3120_n632# 0.03fF
C634 a_n3750_n632# a_n2700_n632# 0.01fF
C635 a_n3540_n632# a_n2910_n632# 0.01fF
C636 a_914_n401# a_960_n100# 0.00fF
C637 a_1080_n632# a_1920_n632# 0.01fF
C638 a_1170_n100# a_1288_n100# 0.07fF
C639 a_n2608_n632# a_n1440_n632# 0.01fF
C640 a_n2398_n632# a_n1650_n632# 0.01fF
C641 a_n2280_n632# a_n1768_n632# 0.01fF
C642 a_n2490_n632# a_n1558_n632# 0.01fF
C643 a_n2700_n632# a_n1348_n632# 0.00fF
C644 w_n4520_n851# a_n2446_n401# 0.10fF
C645 a_n2028_131# a_n978_n197# 0.00fF
C646 a_122_n632# a_n1348_n632# 0.00fF
C647 a_n3028_n632# a_n3076_n729# 0.00fF
C648 a_n2028_131# w_n4520_n851# 0.12fF
C649 a_1498_n100# a_1288_n100# 0.03fF
C650 a_1590_n100# a_1170_n100# 0.02fF
C651 a_1708_n100# a_1078_n100# 0.01fF
C652 a_2382_n197# a_2802_n197# 0.01fF
C653 a_n2070_n632# a_n1860_n632# 0.03fF
C654 a_1962_n197# a_3222_n197# 0.00fF
C655 a_n2656_n729# a_n1816_n729# 0.01fF
C656 a_2760_n632# a_2970_n632# 0.03fF
C657 a_n3286_n401# a_n1816_n729# 0.00fF
C658 a_n2026_n401# a_n3076_n729# 0.00fF
C659 a_n2866_n401# a_n2236_n729# 0.00fF
C660 a_n2446_n401# a_n2656_n729# 0.00fF
C661 a_542_n632# a_n718_n632# 0.00fF
C662 a_542_n632# a_1802_n632# 0.00fF
C663 a_540_n100# a_1288_n100# 0.01fF
C664 a_n3286_n401# a_n2446_n401# 0.01fF
C665 a_n392_n100# a_868_n100# 0.00fF
C666 a_3852_131# a_2382_n197# 0.00fF
C667 a_28_n100# a_n602_n100# 0.01fF
C668 a_1498_n100# a_1590_n100# 0.09fF
C669 a_1380_n100# a_1708_n100# 0.02fF
C670 a_3482_n632# a_3810_n632# 0.02fF
C671 a_3600_n632# a_3692_n632# 0.09fF
C672 a_3390_n632# a_3902_n632# 0.01fF
C673 a_3390_n632# a_3388_n100# 0.00fF
C674 a_2172_131# a_1962_n197# 0.00fF
C675 a_n2400_n100# a_n2282_n100# 0.07fF
C676 a_1590_n100# a_540_n100# 0.01fF
C677 a_1080_n632# a_2642_n632# 0.00fF
C678 a_1544_n729# a_1964_n729# 0.01fF
C679 a_1124_n729# a_2384_n729# 0.00fF
C680 a_n138_n197# a_n136_n729# 0.01fF
C681 a_2758_n100# a_2802_n197# 0.00fF
C682 w_n4520_n851# a_2174_n401# 0.10fF
C683 a_n2448_131# a_n3288_131# 0.01fF
C684 a_1500_n632# a_1544_n729# 0.00fF
C685 a_n180_n632# w_n4520_n851# 0.01fF
C686 a_1290_n632# a_1592_n632# 0.02fF
C687 a_1172_n632# w_n4520_n851# 0.01fF
C688 a_1382_n632# a_1500_n632# 0.07fF
C689 a_n1652_n100# a_n1442_n100# 0.03fF
C690 a_n1862_n100# a_n1232_n100# 0.01fF
C691 a_n2072_n100# a_n1022_n100# 0.01fF
C692 a_n2190_n100# a_n930_n100# 0.00fF
C693 a_n2282_n100# a_n812_n100# 0.00fF
C694 a_n1770_n100# a_n1350_n100# 0.02fF
C695 a_n1980_n100# a_n1140_n100# 0.01fF
C696 a_n3332_n100# a_n2912_n100# 0.02fF
C697 a_n3240_n100# a_n3030_n100# 0.03fF
C698 a_n1440_n632# a_n1138_n632# 0.02fF
C699 a_n1348_n632# a_n1230_n632# 0.07fF
C700 a_n1558_n632# a_n1020_n632# 0.01fF
C701 a_n1650_n632# a_n928_n632# 0.01fF
C702 w_n4520_n851# a_3062_n632# 0.03fF
C703 a_n1396_n729# a_n556_n729# 0.01fF
C704 a_3432_131# a_3388_n100# 0.00fF
C705 a_n182_n100# w_n4520_n851# 0.02fF
C706 a_n1608_131# a_n1606_n401# 0.01fF
C707 a_n2026_n401# a_n556_n729# 0.00fF
C708 a_n1606_n401# a_n976_n729# 0.00fF
C709 a_n3498_n197# a_n3450_n100# 0.00fF
C710 a_n810_n632# a_n766_n401# 0.00fF
C711 w_n4520_n851# a_4064_n729# 0.11fF
C712 a_4112_n632# a_3600_n632# 0.01fF
C713 a_4020_n632# a_3692_n632# 0.02fF
C714 a_660_n632# a_1592_n632# 0.01fF
C715 a_2640_n100# a_2968_n100# 0.02fF
C716 a_2548_n100# a_3060_n100# 0.01fF
C717 a_2430_n100# a_3178_n100# 0.01fF
C718 a_2758_n100# a_2850_n100# 0.09fF
C719 a_n182_n100# a_330_n100# 0.01fF
C720 a_658_n100# a_1078_n100# 0.02fF
C721 a_750_n100# a_960_n100# 0.03fF
C722 a_2338_n100# a_750_n100# 0.00fF
C723 a_120_n100# a_n812_n100# 0.01fF
C724 a_n392_n100# a_n1442_n100# 0.01fF
C725 a_n510_n100# a_n1350_n100# 0.01fF
C726 a_2592_131# a_1122_n197# 0.00fF
C727 a_702_n197# a_n558_n197# 0.00fF
C728 a_n812_n100# a_n720_n100# 0.09fF
C729 a_n930_n100# a_n602_n100# 0.02fF
C730 a_n3960_n632# a_n3658_n632# 0.02fF
C731 a_n4078_n632# a_n3540_n632# 0.01fF
C732 a_n4170_n632# a_n3448_n632# 0.01fF
C733 a_1380_n100# a_658_n100# 0.01fF
C734 a_30_n632# a_n1020_n632# 0.01fF
C735 a_n3960_n632# a_n3916_n729# 0.00fF
C736 a_332_n632# a_n88_n632# 0.02fF
C737 a_240_n632# a_30_n632# 0.03fF
C738 a_1382_n632# a_2222_n632# 0.01fF
C739 a_1290_n632# a_2340_n632# 0.01fF
C740 a_1500_n632# a_2130_n632# 0.01fF
C741 a_n2868_131# a_n1818_n197# 0.00fF
C742 a_n4126_n401# a_n4078_n632# 0.00fF
C743 a_122_n632# a_1500_n632# 0.00fF
C744 a_n3120_n632# a_n1978_n632# 0.01fF
C745 a_n2910_n632# a_n2188_n632# 0.01fF
C746 a_3808_n100# a_4018_n100# 0.03fF
C747 a_3690_n100# a_4110_n100# 0.02fF
C748 a_n3028_n632# a_n2070_n632# 0.01fF
C749 a_n3238_n632# a_n1860_n632# 0.00fF
C750 a_n2818_n632# a_n2280_n632# 0.01fF
C751 a_1754_n401# a_1752_131# 0.01fF
C752 a_n348_131# a_1122_n197# 0.00fF
C753 a_72_131# a_702_n197# 0.00fF
C754 a_122_n632# a_120_n100# 0.00fF
C755 a_1334_n401# a_2174_n401# 0.01fF
C756 a_n2026_n401# a_n2070_n632# 0.00fF
C757 a_n1608_131# a_n3078_n197# 0.00fF
C758 a_1754_n401# a_284_n729# 0.00fF
C759 a_n2912_n100# w_n4520_n851# 0.03fF
C760 a_1080_n632# w_n4520_n851# 0.01fF
C761 a_494_n401# a_1544_n729# 0.00fF
C762 a_n1608_131# a_n768_131# 0.01fF
C763 a_n180_n632# a_n136_n729# 0.00fF
C764 a_n3122_n100# a_n3120_n632# 0.00fF
C765 a_4020_n632# a_4112_n632# 0.09fF
C766 a_n390_n632# a_n180_n632# 0.03fF
C767 a_n508_n632# a_n88_n632# 0.02fF
C768 a_n1652_n100# a_n182_n100# 0.00fF
C769 a_n1560_n100# a_n300_n100# 0.00fF
C770 a_962_n632# a_n180_n632# 0.01fF
C771 a_1172_n632# a_n390_n632# 0.00fF
C772 a_n2700_n632# a_n2608_n632# 0.09fF
C773 a_2130_n632# a_2222_n632# 0.09fF
C774 a_2850_n100# a_1288_n100# 0.00fF
C775 a_752_n632# a_1382_n632# 0.01fF
C776 a_962_n632# a_1172_n632# 0.03fF
C777 a_120_n100# a_1288_n100# 0.01fF
C778 w_n4520_n851# a_4110_n100# 0.14fF
C779 a_2012_n632# a_3180_n632# 0.01fF
C780 a_1802_n632# a_3390_n632# 0.00fF
C781 a_1920_n632# a_3272_n632# 0.00fF
C782 a_n2610_n100# a_n3660_n100# 0.01fF
C783 a_n2820_n100# a_n3450_n100# 0.01fF
C784 a_238_n100# a_n1022_n100# 0.00fF
C785 a_n2492_n100# a_n3752_n100# 0.00fF
C786 a_n2702_n100# a_n3542_n100# 0.01fF
C787 a_n1770_n100# a_n1768_n632# 0.00fF
C788 a_n298_n632# a_n300_n100# 0.00fF
C789 a_2594_n401# a_2804_n729# 0.00fF
C790 a_2174_n401# a_3224_n729# 0.00fF
C791 a_2128_n100# a_960_n100# 0.01fF
C792 a_n1608_131# a_n1650_n632# 0.00fF
C793 a_n3962_n100# a_n3870_n100# 0.09fF
C794 a_n4080_n100# a_n3752_n100# 0.02fF
C795 a_n4172_n100# a_n3660_n100# 0.01fF
C796 a_1498_n100# a_2968_n100# 0.00fF
C797 a_1590_n100# a_2850_n100# 0.00fF
C798 a_2128_n100# a_2338_n100# 0.03fF
C799 a_2010_n100# a_2430_n100# 0.02fF
C800 a_1918_n100# a_2548_n100# 0.01fF
C801 a_1800_n100# a_2640_n100# 0.01fF
C802 a_1708_n100# a_2758_n100# 0.01fF
C803 a_1590_n100# a_120_n100# 0.00fF
C804 a_2640_n100# a_3388_n100# 0.01fF
C805 a_2548_n100# a_3480_n100# 0.01fF
C806 a_2430_n100# a_3598_n100# 0.01fF
C807 a_2338_n100# a_3690_n100# 0.00fF
C808 a_2758_n100# a_3270_n100# 0.01fF
C809 a_1122_n197# a_1332_131# 0.00fF
C810 a_702_n197# a_1752_131# 0.00fF
C811 a_450_n632# a_n298_n632# 0.01fF
C812 a_n508_n632# a_n1768_n632# 0.00fF
C813 a_n810_n632# a_n1440_n632# 0.01fF
C814 a_n600_n632# a_n1650_n632# 0.01fF
C815 a_n718_n632# a_n1558_n632# 0.01fF
C816 a_240_n632# a_1290_n632# 0.01fF
C817 a_n392_n100# a_n182_n100# 0.03fF
C818 a_n510_n100# a_n90_n100# 0.02fF
C819 a_540_n100# a_n602_n100# 0.01fF
C820 a_2010_n100# a_448_n100# 0.00fF
C821 a_n298_n632# a_n1860_n632# 0.00fF
C822 a_3224_n729# a_4064_n729# 0.01fF
C823 a_752_n632# a_2130_n632# 0.00fF
C824 a_2340_n632# a_3600_n632# 0.00fF
C825 a_2432_n632# a_3482_n632# 0.01fF
C826 a_2852_n632# a_3062_n632# 0.03fF
C827 a_2550_n632# a_3390_n632# 0.01fF
C828 a_2642_n632# a_3272_n632# 0.01fF
C829 a_2222_n632# a_3692_n632# 0.00fF
C830 a_2760_n632# a_3180_n632# 0.02fF
C831 a_n556_n729# a_704_n729# 0.00fF
C832 a_332_n632# a_542_n632# 0.03fF
C833 a_122_n632# a_752_n632# 0.01fF
C834 a_240_n632# a_660_n632# 0.02fF
C835 a_n2072_n100# a_n2492_n100# 0.02fF
C836 a_n1862_n100# a_n2702_n100# 0.01fF
C837 a_n1652_n100# a_n2912_n100# 0.00fF
C838 a_n1770_n100# a_n2820_n100# 0.01fF
C839 a_n1980_n100# a_n2610_n100# 0.01fF
C840 a_n1560_n100# a_n3030_n100# 0.00fF
C841 w_n4520_n851# a_n2910_n632# 0.03fF
C842 a_3434_n401# a_1964_n729# 0.00fF
C843 w_n4520_n851# a_960_n100# 0.02fF
C844 a_2338_n100# w_n4520_n851# 0.02fF
C845 a_n3708_131# a_n3752_n100# 0.00fF
C846 a_n2400_n100# a_n3752_n100# 0.00fF
C847 a_n2282_n100# a_n3870_n100# 0.00fF
C848 a_n718_n632# a_30_n632# 0.01fF
C849 w_n4520_n851# a_n1232_n100# 0.02fF
C850 a_n3918_n197# a_n3078_n197# 0.01fF
C851 a_n3868_n632# a_n2398_n632# 0.00fF
C852 a_1080_n632# a_n390_n632# 0.00fF
C853 a_n3238_n632# a_n3028_n632# 0.03fF
C854 a_n3330_n632# a_n2910_n632# 0.02fF
C855 a_n3448_n632# a_n2818_n632# 0.01fF
C856 a_n3750_n632# a_n2490_n632# 0.00fF
C857 a_n346_n401# a_914_n401# 0.00fF
C858 w_n4520_n851# a_n1606_n401# 0.10fF
C859 a_n2280_n632# a_n1558_n632# 0.01fF
C860 a_n2700_n632# a_n1138_n632# 0.00fF
C861 a_n2490_n632# a_n1348_n632# 0.01fF
C862 a_n2188_n632# a_n1650_n632# 0.01fF
C863 a_n2398_n632# a_n1440_n632# 0.01fF
C864 a_n2608_n632# a_n1230_n632# 0.00fF
C865 a_n2070_n632# a_n1768_n632# 0.02fF
C866 a_n1608_131# a_n2238_n197# 0.00fF
C867 a_330_n100# a_960_n100# 0.01fF
C868 a_238_n100# a_1078_n100# 0.01fF
C869 a_962_n632# a_1080_n632# 0.07fF
C870 a_122_n632# a_n1138_n632# 0.00fF
C871 a_330_n100# a_n1232_n100# 0.00fF
C872 a_n2448_131# a_n1818_n197# 0.00fF
C873 a_1708_n100# a_1288_n100# 0.02fF
C874 a_1800_n100# a_1170_n100# 0.01fF
C875 a_1918_n100# a_1078_n100# 0.01fF
C876 a_1380_n100# a_238_n100# 0.01fF
C877 a_2802_n197# a_3222_n197# 0.01fF
C878 a_2382_n197# a_3642_n197# 0.00fF
C879 a_n2236_n729# a_n1396_n729# 0.01fF
C880 a_n2446_n401# a_n1816_n729# 0.00fF
C881 a_n2026_n401# a_n2236_n729# 0.00fF
C882 a_n1606_n401# a_n2656_n729# 0.00fF
C883 a_n2866_n401# a_n1396_n729# 0.00fF
C884 a_542_n632# a_n508_n632# 0.01fF
C885 a_542_n632# a_2012_n632# 0.00fF
C886 a_n182_n100# a_868_n100# 0.01fF
C887 a_n2866_n401# a_n2026_n401# 0.01fF
C888 a_3852_131# a_3222_n197# 0.00fF
C889 a_3692_n632# a_3810_n632# 0.07fF
C890 a_1590_n100# a_1708_n100# 0.07fF
C891 a_1498_n100# a_1800_n100# 0.02fF
C892 a_1380_n100# a_1918_n100# 0.01fF
C893 a_3600_n632# a_3902_n632# 0.02fF
C894 a_658_n100# a_n812_n100# 0.00fF
C895 a_3482_n632# a_3480_n100# 0.00fF
C896 a_2172_131# a_2802_n197# 0.00fF
C897 a_n2400_n100# a_n2072_n100# 0.02fF
C898 a_n2282_n100# a_n2190_n100# 0.09fF
C899 a_1800_n100# a_540_n100# 0.00fF
C900 a_3432_131# a_2592_131# 0.01fF
C901 a_1964_n729# a_2384_n729# 0.01fF
C902 a_n768_131# a_n978_n197# 0.00fF
C903 w_n4520_n851# a_3014_n401# 0.10fF
C904 a_n180_n632# a_n138_n197# 0.00fF
C905 w_n4520_n851# a_n3078_n197# 0.10fF
C906 w_n4520_n851# a_n768_131# 0.12fF
C907 a_1500_n632# a_1592_n632# 0.09fF
C908 a_1382_n632# a_1710_n632# 0.02fF
C909 a_1290_n632# a_1802_n632# 0.01fF
C910 a_n2190_n100# a_n720_n100# 0.00fF
C911 a_n1770_n100# a_n1140_n100# 0.01fF
C912 a_n1980_n100# a_n930_n100# 0.01fF
C913 a_n1560_n100# a_n1350_n100# 0.03fF
C914 a_n1862_n100# a_n1022_n100# 0.01fF
C915 a_n1652_n100# a_n1232_n100# 0.02fF
C916 a_n2072_n100# a_n812_n100# 0.00fF
C917 a_n3240_n100# a_n2820_n100# 0.02fF
C918 a_n3332_n100# a_n2702_n100# 0.01fF
C919 a_n3122_n100# a_n2912_n100# 0.03fF
C920 a_n346_n401# a_n976_n729# 0.00fF
C921 a_n182_n100# a_n138_n197# 0.00fF
C922 a_n1348_n632# a_n1020_n632# 0.02fF
C923 a_n1440_n632# a_n928_n632# 0.01fF
C924 a_n1230_n632# a_n1138_n632# 0.09fF
C925 w_n4520_n851# a_3272_n632# 0.03fF
C926 a_240_n632# a_n1348_n632# 0.00fF
C927 a_238_n100# a_282_n197# 0.00fF
C928 a_962_n632# a_960_n100# 0.00fF
C929 a_n766_n401# a_n976_n729# 0.00fF
C930 a_n1606_n401# a_n136_n729# 0.00fF
C931 a_n1186_n401# a_n556_n729# 0.00fF
C932 a_n810_n632# a_n812_n100# 0.00fF
C933 a_4020_n632# a_3902_n632# 0.07fF
C934 w_n4520_n851# a_n4078_n632# 0.08fF
C935 a_4112_n632# a_3810_n632# 0.02fF
C936 a_660_n632# a_n718_n632# 0.00fF
C937 a_n2658_n197# a_n3498_n197# 0.01fF
C938 a_660_n632# a_1802_n632# 0.01fF
C939 a_2758_n100# a_3060_n100# 0.02fF
C940 a_2850_n100# a_2968_n100# 0.07fF
C941 a_2640_n100# a_3178_n100# 0.01fF
C942 a_658_n100# a_1288_n100# 0.01fF
C943 w_n4520_n851# a_n1650_n632# 0.01fF
C944 a_n392_n100# a_960_n100# 0.00fF
C945 a_n348_131# a_n1818_n197# 0.00fF
C946 a_120_n100# a_n602_n100# 0.01fF
C947 a_n2400_n100# a_n2398_n632# 0.00fF
C948 a_2592_131# a_1962_n197# 0.00fF
C949 a_n182_n100# a_n1442_n100# 0.00fF
C950 a_n510_n100# a_n1140_n100# 0.01fF
C951 a_n392_n100# a_n1232_n100# 0.01fF
C952 a_n300_n100# a_n1350_n100# 0.01fF
C953 a_n4170_n632# a_n3238_n632# 0.01fF
C954 a_n3750_n632# a_n3658_n632# 0.09fF
C955 a_n720_n100# a_n602_n100# 0.07fF
C956 a_n3960_n632# a_n3448_n632# 0.01fF
C957 a_n3868_n632# a_n3540_n632# 0.02fF
C958 a_n4078_n632# a_n3330_n632# 0.01fF
C959 a_n3238_n632# a_n1768_n632# 0.00fF
C960 a_1590_n100# a_658_n100# 0.01fF
C961 a_1290_n632# a_2550_n632# 0.00fF
C962 a_1500_n632# a_2340_n632# 0.01fF
C963 a_1382_n632# a_2432_n632# 0.01fF
C964 a_1710_n632# a_2130_n632# 0.02fF
C965 a_1592_n632# a_2222_n632# 0.01fF
C966 a_122_n632# a_n810_n632# 0.01fF
C967 a_122_n632# a_1710_n632# 0.00fF
C968 a_n510_n100# a_448_n100# 0.01fF
C969 a_3900_n100# a_4110_n100# 0.03fF
C970 a_n2818_n632# a_n2070_n632# 0.01fF
C971 a_n3028_n632# a_n1860_n632# 0.01fF
C972 a_n2910_n632# a_n1978_n632# 0.01fF
C973 a_3012_131# a_1752_131# 0.00fF
C974 a_n4128_131# a_n4126_n401# 0.01fF
C975 a_n3288_131# a_n3240_n100# 0.00fF
C976 a_1754_n401# a_2594_n401# 0.01fF
C977 a_n2702_n100# w_n4520_n851# 0.02fF
C978 a_2010_n100# a_1962_n197# 0.00fF
C979 a_2640_n100# a_2592_131# 0.00fF
C980 a_3222_n197# a_3270_n100# 0.00fF
C981 a_n2238_n197# a_n978_n197# 0.00fF
C982 a_n1818_n197# a_n1398_n197# 0.01fF
C983 w_n4520_n851# a_4062_n197# 0.10fF
C984 a_n3030_n100# a_n3028_n632# 0.00fF
C985 w_n4520_n851# a_n2238_n197# 0.10fF
C986 a_n298_n632# a_n88_n632# 0.03fF
C987 a_n1560_n100# a_n90_n100# 0.00fF
C988 a_1172_n632# a_n180_n632# 0.00fF
C989 a_n2912_n100# a_n1442_n100# 0.00fF
C990 a_n2700_n632# a_n2398_n632# 0.02fF
C991 a_n2608_n632# a_n2490_n632# 0.07fF
C992 a_3434_n401# a_3854_n401# 0.01fF
C993 a_2130_n632# a_2432_n632# 0.02fF
C994 a_2222_n632# a_2340_n632# 0.07fF
C995 a_752_n632# a_1592_n632# 0.01fF
C996 a_750_n100# a_1078_n100# 0.02fF
C997 a_868_n100# a_960_n100# 0.09fF
C998 a_n2820_n100# a_n2866_n401# 0.00fF
C999 a_1920_n632# a_3482_n632# 0.00fF
C1000 a_2012_n632# a_3390_n632# 0.00fF
C1001 a_2338_n100# a_868_n100# 0.00fF
C1002 a_492_131# a_n978_n197# 0.00fF
C1003 a_n2492_n100# a_n3542_n100# 0.01fF
C1004 a_n2610_n100# a_n3450_n100# 0.01fF
C1005 a_238_n100# a_n812_n100# 0.01fF
C1006 a_n1652_n100# a_n1650_n632# 0.00fF
C1007 a_n180_n632# a_n182_n100# 0.00fF
C1008 a_2594_n401# a_3644_n729# 0.00fF
C1009 a_3014_n401# a_3224_n729# 0.00fF
C1010 a_n4126_n401# a_n4080_n100# 0.00fF
C1011 a_n3870_n100# a_n3752_n100# 0.07fF
C1012 a_n4172_n100# a_n3450_n100# 0.01fF
C1013 a_n3962_n100# a_n3660_n100# 0.02fF
C1014 a_n4080_n100# a_n3542_n100# 0.01fF
C1015 a_2220_n100# a_2430_n100# 0.03fF
C1016 a_2128_n100# a_2548_n100# 0.02fF
C1017 a_2010_n100# a_2640_n100# 0.01fF
C1018 w_n4520_n851# a_492_131# 0.12fF
C1019 a_1918_n100# a_2758_n100# 0.01fF
C1020 a_1800_n100# a_2850_n100# 0.01fF
C1021 a_1708_n100# a_2968_n100# 0.00fF
C1022 a_1590_n100# a_3060_n100# 0.00fF
C1023 a_2758_n100# a_3480_n100# 0.01fF
C1024 a_2968_n100# a_3270_n100# 0.02fF
C1025 a_2850_n100# a_3388_n100# 0.01fF
C1026 a_1380_n100# a_750_n100# 0.01fF
C1027 a_2640_n100# a_3598_n100# 0.01fF
C1028 a_2548_n100# a_3690_n100# 0.01fF
C1029 a_2430_n100# a_3808_n100# 0.00fF
C1030 a_2338_n100# a_3900_n100# 0.00fF
C1031 a_1962_n197# a_1332_131# 0.00fF
C1032 w_n4520_n851# a_1542_n197# 0.10fF
C1033 a_450_n632# a_n88_n632# 0.01fF
C1034 a_332_n632# a_30_n632# 0.02fF
C1035 a_n600_n632# a_n1440_n632# 0.01fF
C1036 a_n390_n632# a_n1650_n632# 0.00fF
C1037 a_n298_n632# a_n1768_n632# 0.00fF
C1038 a_n718_n632# a_n1348_n632# 0.01fF
C1039 a_n508_n632# a_n1558_n632# 0.01fF
C1040 a_n810_n632# a_n1230_n632# 0.02fF
C1041 a_240_n632# a_1500_n632# 0.00fF
C1042 a_n300_n100# a_n90_n100# 0.03fF
C1043 a_3012_131# a_2970_n632# 0.00fF
C1044 a_3272_n632# a_3224_n729# 0.00fF
C1045 a_72_131# a_1122_n197# 0.00fF
C1046 a_1754_n401# a_704_n729# 0.00fF
C1047 a_1290_n632# a_1332_131# 0.00fF
C1048 a_914_n401# a_1544_n729# 0.00fF
C1049 a_752_n632# a_2340_n632# 0.00fF
C1050 a_2432_n632# a_3692_n632# 0.00fF
C1051 a_2970_n632# a_3180_n632# 0.03fF
C1052 a_2642_n632# a_3482_n632# 0.01fF
C1053 a_2852_n632# a_3272_n632# 0.02fF
C1054 a_2340_n632# a_3810_n632# 0.00fF
C1055 a_2760_n632# a_3390_n632# 0.01fF
C1056 a_2550_n632# a_3600_n632# 0.01fF
C1057 a_284_n729# a_704_n729# 0.01fF
C1058 a_n1770_n100# a_n2610_n100# 0.01fF
C1059 a_n1862_n100# a_n2492_n100# 0.01fF
C1060 a_n1560_n100# a_n2820_n100# 0.00fF
C1061 a_n1652_n100# a_n2702_n100# 0.01fF
C1062 a_n978_n197# a_n1022_n100# 0.00fF
C1063 w_n4520_n851# a_n346_n401# 0.10fF
C1064 a_n3122_n100# a_n3078_n197# 0.00fF
C1065 a_3854_n401# a_2384_n729# 0.00fF
C1066 a_2548_n100# w_n4520_n851# 0.02fF
C1067 a_n2400_n100# a_n3542_n100# 0.01fF
C1068 a_n2190_n100# a_n3752_n100# 0.00fF
C1069 a_n508_n632# a_30_n632# 0.01fF
C1070 a_n2282_n100# a_n3660_n100# 0.00fF
C1071 w_n4520_n851# a_n1022_n100# 0.02fF
C1072 a_n1770_n100# a_n1818_n197# 0.00fF
C1073 a_n3120_n632# a_n2910_n632# 0.03fF
C1074 a_n3750_n632# a_n2280_n632# 0.00fF
C1075 a_1080_n632# a_n180_n632# 0.00fF
C1076 a_n3238_n632# a_n2818_n632# 0.02fF
C1077 a_n2398_n632# a_n1230_n632# 0.01fF
C1078 w_n4520_n851# a_n766_n401# 0.10fF
C1079 a_n2070_n632# a_n1558_n632# 0.01fF
C1080 a_n2608_n632# a_n1020_n632# 0.00fF
C1081 a_n2490_n632# a_n1138_n632# 0.00fF
C1082 a_n1978_n632# a_n1650_n632# 0.02fF
C1083 a_n2280_n632# a_n1348_n632# 0.01fF
C1084 a_n2188_n632# a_n1440_n632# 0.01fF
C1085 a_n1860_n632# a_n1768_n632# 0.09fF
C1086 a_870_n632# a_1382_n632# 0.01fF
C1087 a_238_n100# a_1288_n100# 0.01fF
C1088 a_1080_n632# a_1172_n632# 0.09fF
C1089 a_122_n632# a_n928_n632# 0.01fF
C1090 a_n3288_131# a_n2658_n197# 0.00fF
C1091 a_330_n100# a_n1022_n100# 0.00fF
C1092 a_n2866_n401# a_n2818_n632# 0.00fF
C1093 a_n1442_n100# a_n1232_n100# 0.03fF
C1094 a_1918_n100# a_1288_n100# 0.01fF
C1095 a_2010_n100# a_1170_n100# 0.01fF
C1096 a_2128_n100# a_1078_n100# 0.01fF
C1097 a_3222_n197# a_3642_n197# 0.01fF
C1098 a_n1350_n100# a_n1396_n729# 0.00fF
C1099 a_1590_n100# a_238_n100# 0.00fF
C1100 a_1122_n197# a_1752_131# 0.00fF
C1101 a_n2026_n401# a_n1396_n729# 0.00fF
C1102 a_542_n632# a_n298_n632# 0.01fF
C1103 a_n1186_n401# a_n2236_n729# 0.00fF
C1104 a_n1606_n401# a_n1816_n729# 0.00fF
C1105 a_n2446_n401# a_n1606_n401# 0.01fF
C1106 a_332_n632# a_1290_n632# 0.01fF
C1107 a_912_131# a_914_n401# 0.01fF
C1108 a_n510_n100# a_28_n100# 0.01fF
C1109 a_3810_n632# a_3902_n632# 0.09fF
C1110 a_1708_n100# a_1800_n100# 0.09fF
C1111 a_1590_n100# a_1918_n100# 0.02fF
C1112 a_1498_n100# a_2010_n100# 0.01fF
C1113 a_1380_n100# a_2128_n100# 0.01fF
C1114 a_658_n100# a_n602_n100# 0.00fF
C1115 a_2172_131# a_3642_n197# 0.00fF
C1116 a_1800_n100# a_3270_n100# 0.00fF
C1117 a_3600_n632# a_3598_n100# 0.00fF
C1118 a_3270_n100# a_3388_n100# 0.07fF
C1119 a_n3540_n632# a_n2700_n632# 0.01fF
C1120 a_n3658_n632# a_n2608_n632# 0.01fF
C1121 a_702_n197# a_704_n729# 0.01fF
C1122 a_n2282_n100# a_n1980_n100# 0.02fF
C1123 a_n2190_n100# a_n2072_n100# 0.07fF
C1124 a_n2400_n100# a_n1862_n100# 0.01fF
C1125 a_2010_n100# a_540_n100# 0.00fF
C1126 a_n4128_131# a_n3918_n197# 0.00fF
C1127 a_870_n632# a_912_131# 0.00fF
C1128 a_4020_n632# a_2550_n632# 0.00fF
C1129 a_870_n632# a_2130_n632# 0.00fF
C1130 a_4064_n729# a_4110_n100# 0.00fF
C1131 a_n768_131# a_n138_n197# 0.00fF
C1132 a_240_n632# a_752_n632# 0.01fF
C1133 a_122_n632# a_870_n632# 0.01fF
C1134 a_332_n632# a_660_n632# 0.02fF
C1135 a_450_n632# a_542_n632# 0.09fF
C1136 w_n4520_n851# a_1078_n100# 0.02fF
C1137 a_n3078_n197# a_n3120_n632# 0.00fF
C1138 a_1382_n632# a_1920_n632# 0.01fF
C1139 a_1290_n632# a_2012_n632# 0.01fF
C1140 a_1500_n632# a_1802_n632# 0.02fF
C1141 a_1592_n632# a_1710_n632# 0.07fF
C1142 a_n1862_n100# a_n812_n100# 0.01fF
C1143 a_n1652_n100# a_n1022_n100# 0.01fF
C1144 a_n3030_n100# a_n2820_n100# 0.03fF
C1145 a_n2072_n100# a_n602_n100# 0.00fF
C1146 a_n3332_n100# a_n2492_n100# 0.01fF
C1147 a_n3240_n100# a_n2610_n100# 0.01fF
C1148 a_n1770_n100# a_n930_n100# 0.01fF
C1149 a_n1980_n100# a_n720_n100# 0.00fF
C1150 a_330_n100# a_1078_n100# 0.01fF
C1151 a_n3122_n100# a_n2702_n100# 0.02fF
C1152 a_n1560_n100# a_n1140_n100# 0.02fF
C1153 a_n1138_n632# a_n1020_n632# 0.07fF
C1154 a_n1230_n632# a_n928_n632# 0.02fF
C1155 a_74_n401# a_n556_n729# 0.00fF
C1156 a_n346_n401# a_n136_n729# 0.00fF
C1157 w_n4520_n851# a_3482_n632# 0.03fF
C1158 a_1380_n100# w_n4520_n851# 0.02fF
C1159 a_240_n632# a_n1138_n632# 0.00fF
C1160 a_n390_n632# a_n346_n401# 0.00fF
C1161 a_n3332_n100# a_n4080_n100# 0.01fF
C1162 a_n3240_n100# a_n4172_n100# 0.01fF
C1163 a_n766_n401# a_n136_n729# 0.00fF
C1164 a_n1186_n401# a_284_n729# 0.00fF
C1165 a_n718_n632# a_n720_n100# 0.00fF
C1166 a_1380_n100# a_330_n100# 0.01fF
C1167 a_702_n197# a_1122_n197# 0.01fF
C1168 a_n2028_131# a_n3078_n197# 0.00fF
C1169 w_n4520_n851# a_n3868_n632# 0.05fF
C1170 a_660_n632# a_n508_n632# 0.01fF
C1171 a_660_n632# a_2012_n632# 0.00fF
C1172 a_2968_n100# a_3060_n100# 0.09fF
C1173 a_2850_n100# a_3178_n100# 0.02fF
C1174 w_n4520_n851# a_n1440_n632# 0.01fF
C1175 a_3902_n632# a_3854_n401# 0.00fF
C1176 a_n182_n100# a_960_n100# 0.01fF
C1177 a_n1608_131# a_n1188_131# 0.01fF
C1178 a_n2028_131# a_n768_131# 0.00fF
C1179 a_3480_n100# a_3434_n401# 0.00fF
C1180 a_n4128_131# w_n4520_n851# 0.14fF
C1181 a_n2282_n100# a_n2280_n632# 0.00fF
C1182 a_750_n100# a_n812_n100# 0.00fF
C1183 a_2592_131# a_2802_n197# 0.00fF
C1184 a_n510_n100# a_n930_n100# 0.02fF
C1185 a_n392_n100# a_n1022_n100# 0.01fF
C1186 a_n300_n100# a_n1140_n100# 0.01fF
C1187 a_n182_n100# a_n1232_n100# 0.01fF
C1188 a_n90_n100# a_n1350_n100# 0.00fF
C1189 a_n3960_n632# a_n3238_n632# 0.01fF
C1190 a_n4170_n632# a_n3028_n632# 0.01fF
C1191 a_n3868_n632# a_n3330_n632# 0.01fF
C1192 a_n4078_n632# a_n3120_n632# 0.01fF
C1193 a_n3750_n632# a_n3448_n632# 0.02fF
C1194 a_2432_n632# a_2384_n729# 0.00fF
C1195 a_n3120_n632# a_n1650_n632# 0.00fF
C1196 a_n3028_n632# a_n1768_n632# 0.00fF
C1197 a_1800_n100# a_658_n100# 0.01fF
C1198 a_3852_131# a_2592_131# 0.00fF
C1199 a_1592_n632# a_2432_n632# 0.01fF
C1200 a_1290_n632# a_2760_n632# 0.00fF
C1201 a_1802_n632# a_2222_n632# 0.02fF
C1202 a_1382_n632# a_2642_n632# 0.00fF
C1203 a_1500_n632# a_2550_n632# 0.01fF
C1204 a_1920_n632# a_2130_n632# 0.03fF
C1205 a_1710_n632# a_2340_n632# 0.01fF
C1206 a_122_n632# a_n600_n632# 0.01fF
C1207 a_n3706_n401# a_n3750_n632# 0.00fF
C1208 a_n300_n100# a_448_n100# 0.01fF
C1209 a_n2818_n632# a_n1860_n632# 0.01fF
C1210 a_n2400_n100# a_n3332_n100# 0.01fF
C1211 a_282_n197# a_n978_n197# 0.00fF
C1212 a_450_n632# a_448_n100# 0.00fF
C1213 a_n3708_131# a_n3918_n197# 0.00fF
C1214 a_2174_n401# a_3014_n401# 0.01fF
C1215 w_n4520_n851# a_282_n197# 0.10fF
C1216 a_n2492_n100# w_n4520_n851# 0.02fF
C1217 a_n1818_n197# a_n558_n197# 0.00fF
C1218 w_n4520_n851# a_n4080_n100# 0.08fF
C1219 a_30_n632# a_72_131# 0.00fF
C1220 a_n2912_n100# a_n2910_n632# 0.00fF
C1221 a_330_n100# a_282_n197# 0.00fF
C1222 a_3014_n401# a_3062_n632# 0.00fF
C1223 a_1380_n100# a_1334_n401# 0.00fF
C1224 a_2010_n100# a_1964_n729# 0.00fF
C1225 a_n2702_n100# a_n1442_n100# 0.00fF
C1226 a_n2820_n100# a_n1350_n100# 0.00fF
C1227 a_n2608_n632# a_n2280_n632# 0.02fF
C1228 a_n2490_n632# a_n2398_n632# 0.09fF
C1229 a_n2700_n632# a_n2188_n632# 0.01fF
C1230 a_2340_n632# a_2432_n632# 0.09fF
C1231 a_2222_n632# a_2550_n632# 0.02fF
C1232 a_2130_n632# a_2642_n632# 0.01fF
C1233 a_752_n632# a_n718_n632# 0.00fF
C1234 a_752_n632# a_1802_n632# 0.01fF
C1235 a_750_n100# a_1288_n100# 0.01fF
C1236 a_2012_n632# a_3600_n632# 0.00fF
C1237 a_n392_n100# a_1078_n100# 0.00fF
C1238 a_492_131# a_n138_n197# 0.00fF
C1239 a_28_n100# a_72_131# 0.00fF
C1240 a_238_n100# a_n602_n100# 0.01fF
C1241 a_n1560_n100# a_n1558_n632# 0.00fF
C1242 a_n88_n632# a_n90_n100# 0.00fF
C1243 a_3014_n401# a_4064_n729# 0.00fF
C1244 a_3062_n632# a_3272_n632# 0.03fF
C1245 a_n2610_n100# a_n2658_n197# 0.00fF
C1246 a_n3962_n100# a_n3450_n100# 0.01fF
C1247 a_n3870_n100# a_n3542_n100# 0.02fF
C1248 a_n3752_n100# a_n3660_n100# 0.09fF
C1249 a_2220_n100# a_2640_n100# 0.02fF
C1250 a_2128_n100# a_2758_n100# 0.01fF
C1251 a_2010_n100# a_2850_n100# 0.01fF
C1252 a_1918_n100# a_2968_n100# 0.01fF
C1253 a_1800_n100# a_3060_n100# 0.00fF
C1254 a_1708_n100# a_3178_n100# 0.00fF
C1255 a_1590_n100# a_750_n100# 0.01fF
C1256 a_2640_n100# a_3808_n100# 0.01fF
C1257 a_2548_n100# a_3900_n100# 0.00fF
C1258 a_2430_n100# a_4018_n100# 0.00fF
C1259 a_2758_n100# a_3690_n100# 0.01fF
C1260 a_3178_n100# a_3270_n100# 0.09fF
C1261 a_3060_n100# a_3388_n100# 0.02fF
C1262 a_2968_n100# a_3480_n100# 0.01fF
C1263 a_2850_n100# a_3598_n100# 0.01fF
C1264 w_n4520_n851# a_2382_n197# 0.10fF
C1265 a_2802_n197# a_1332_131# 0.00fF
C1266 a_n718_n632# a_n1138_n632# 0.02fF
C1267 a_n298_n632# a_n1558_n632# 0.00fF
C1268 a_n600_n632# a_n1230_n632# 0.01fF
C1269 a_n508_n632# a_n1348_n632# 0.01fF
C1270 a_n180_n632# a_n1650_n632# 0.00fF
C1271 a_n810_n632# a_n1020_n632# 0.03fF
C1272 a_n390_n632# a_n1440_n632# 0.01fF
C1273 a_240_n632# a_n810_n632# 0.01fF
C1274 a_240_n632# a_1710_n632# 0.00fF
C1275 a_n2028_131# a_n2238_n197# 0.00fF
C1276 a_n2658_n197# a_n1818_n197# 0.01fF
C1277 a_n510_n100# a_540_n100# 0.01fF
C1278 a_n3708_131# w_n4520_n851# 0.13fF
C1279 a_n2400_n100# w_n4520_n851# 0.02fF
C1280 w_n4520_n851# a_1544_n729# 0.12fF
C1281 a_914_n401# a_2384_n729# 0.00fF
C1282 a_1382_n632# w_n4520_n851# 0.01fF
C1283 a_2550_n632# a_3810_n632# 0.00fF
C1284 a_2760_n632# a_3600_n632# 0.01fF
C1285 a_2128_n100# a_2130_n632# 0.00fF
C1286 a_2432_n632# a_3902_n632# 0.00fF
C1287 a_2852_n632# a_3482_n632# 0.01fF
C1288 a_2970_n632# a_3390_n632# 0.02fF
C1289 a_2642_n632# a_3692_n632# 0.01fF
C1290 a_n1560_n100# a_n2610_n100# 0.01fF
C1291 a_n1652_n100# a_n2492_n100# 0.01fF
C1292 a_2758_n100# w_n4520_n851# 0.02fF
C1293 a_n2282_n100# a_n3450_n100# 0.01fF
C1294 a_n2190_n100# a_n3542_n100# 0.00fF
C1295 a_n2072_n100# a_n3660_n100# 0.00fF
C1296 a_n298_n632# a_30_n632# 0.02fF
C1297 w_n4520_n851# a_n812_n100# 0.02fF
C1298 a_n1560_n100# a_28_n100# 0.00fF
C1299 a_n3028_n632# a_n2818_n632# 0.03fF
C1300 a_n1978_n632# a_n1440_n632# 0.01fF
C1301 a_n2070_n632# a_n1348_n632# 0.01fF
C1302 a_n2280_n632# a_n1138_n632# 0.01fF
C1303 a_n2188_n632# a_n1230_n632# 0.01fF
C1304 a_n1860_n632# a_n1558_n632# 0.02fF
C1305 a_n2490_n632# a_n928_n632# 0.00fF
C1306 a_n2398_n632# a_n1020_n632# 0.00fF
C1307 a_870_n632# a_1592_n632# 0.01fF
C1308 a_868_n100# a_1078_n100# 0.03fF
C1309 a_72_131# a_74_n401# 0.01fF
C1310 a_2338_n100# a_960_n100# 0.00fF
C1311 a_n1188_131# a_n978_n197# 0.00fF
C1312 a_330_n100# a_n812_n100# 0.01fF
C1313 a_n346_n401# a_n1816_n729# 0.00fF
C1314 a_n1350_n100# a_n1140_n100# 0.03fF
C1315 a_2128_n100# a_1288_n100# 0.01fF
C1316 a_2220_n100# a_1170_n100# 0.01fF
C1317 w_n4520_n851# a_n1188_131# 0.12fF
C1318 a_n1442_n100# a_n1022_n100# 0.02fF
C1319 w_n4520_n851# a_912_131# 0.12fF
C1320 a_1800_n100# a_238_n100# 0.00fF
C1321 a_1380_n100# a_868_n100# 0.01fF
C1322 a_1962_n197# a_1752_131# 0.00fF
C1323 a_542_n632# a_n88_n632# 0.01fF
C1324 a_n1186_n401# a_n1396_n729# 0.00fF
C1325 a_450_n632# a_30_n632# 0.02fF
C1326 a_n766_n401# a_n1816_n729# 0.00fF
C1327 w_n4520_n851# a_n2700_n632# 0.02fF
C1328 w_n4520_n851# a_2130_n632# 0.01fF
C1329 a_n2026_n401# a_n1186_n401# 0.01fF
C1330 a_122_n632# w_n4520_n851# 0.01fF
C1331 a_332_n632# a_1500_n632# 0.01fF
C1332 a_n300_n100# a_28_n100# 0.02fF
C1333 a_1800_n100# a_1918_n100# 0.07fF
C1334 a_1708_n100# a_2010_n100# 0.02fF
C1335 a_1590_n100# a_2128_n100# 0.01fF
C1336 a_1498_n100# a_2220_n100# 0.01fF
C1337 a_2010_n100# a_3270_n100# 0.00fF
C1338 a_1918_n100# a_3388_n100# 0.00fF
C1339 a_3692_n632# a_3690_n100# 0.00fF
C1340 a_4064_n729# a_4062_n197# 0.01fF
C1341 a_n3658_n632# a_n2398_n632# 0.00fF
C1342 a_3388_n100# a_3480_n100# 0.09fF
C1343 a_3270_n100# a_3598_n100# 0.02fF
C1344 a_n3330_n632# a_n2700_n632# 0.01fF
C1345 a_n3540_n632# a_n2490_n632# 0.01fF
C1346 a_n3448_n632# a_n2608_n632# 0.01fF
C1347 a_n2190_n100# a_n1862_n100# 0.02fF
C1348 a_n2400_n100# a_n1652_n100# 0.01fF
C1349 a_n2072_n100# a_n1980_n100# 0.09fF
C1350 a_n2282_n100# a_n1770_n100# 0.01fF
C1351 a_240_n632# a_238_n100# 0.00fF
C1352 a_4112_n632# a_2642_n632# 0.00fF
C1353 a_4020_n632# a_2760_n632# 0.00fF
C1354 a_n2700_n632# a_n2656_n729# 0.00fF
C1355 a_1334_n401# a_1544_n729# 0.00fF
C1356 a_1754_n401# a_1124_n729# 0.00fF
C1357 a_870_n632# a_2340_n632# 0.00fF
C1358 a_n3288_131# a_n3498_n197# 0.00fF
C1359 a_284_n729# a_1124_n729# 0.01fF
C1360 a_n1818_n197# a_n1860_n632# 0.00fF
C1361 a_1382_n632# a_1334_n401# 0.00fF
C1362 w_n4520_n851# a_1288_n100# 0.02fF
C1363 a_2012_n632# a_1964_n729# 0.00fF
C1364 a_n810_n632# a_n718_n632# 0.09fF
C1365 a_1290_n632# a_n298_n632# 0.00fF
C1366 a_1592_n632# a_1920_n632# 0.02fF
C1367 a_1500_n632# a_2012_n632# 0.01fF
C1368 a_1710_n632# a_1802_n632# 0.09fF
C1369 a_2802_n197# a_2804_n729# 0.01fF
C1370 a_n1770_n100# a_n720_n100# 0.01fF
C1371 a_n1560_n100# a_n930_n100# 0.01fF
C1372 a_n1862_n100# a_n602_n100# 0.00fF
C1373 a_n1652_n100# a_n812_n100# 0.01fF
C1374 a_330_n100# a_1288_n100# 0.01fF
C1375 a_n2912_n100# a_n2702_n100# 0.03fF
C1376 a_n3030_n100# a_n2610_n100# 0.02fF
C1377 a_n3122_n100# a_n2492_n100# 0.01fF
C1378 a_74_n401# a_284_n729# 0.00fF
C1379 a_962_n632# a_1382_n632# 0.02fF
C1380 a_n1020_n632# a_n928_n632# 0.09fF
C1381 a_1590_n100# w_n4520_n851# 0.02fF
C1382 w_n4520_n851# a_3692_n632# 0.04fF
C1383 a_240_n632# a_n928_n632# 0.01fF
C1384 a_n3030_n100# a_n4172_n100# 0.01fF
C1385 a_n3122_n100# a_n4080_n100# 0.01fF
C1386 a_n3332_n100# a_n3870_n100# 0.01fF
C1387 a_n3240_n100# a_n3962_n100# 0.01fF
C1388 a_2804_n729# a_1964_n729# 0.01fF
C1389 a_n600_n632# a_n602_n100# 0.00fF
C1390 a_1590_n100# a_330_n100# 0.00fF
C1391 a_n3918_n197# a_n3870_n100# 0.00fF
C1392 a_2802_n197# a_2760_n632# 0.00fF
C1393 a_702_n197# a_1962_n197# 0.00fF
C1394 a_660_n632# a_n298_n632# 0.01fF
C1395 a_3060_n100# a_3178_n100# 0.07fF
C1396 w_n4520_n851# a_n1230_n632# 0.01fF
C1397 a_450_n632# a_1290_n632# 0.01fF
C1398 a_n510_n100# a_120_n100# 0.01fF
C1399 a_n2190_n100# a_n2188_n632# 0.00fF
C1400 a_750_n100# a_n602_n100# 0.00fF
C1401 a_2592_131# a_3642_n197# 0.00fF
C1402 a_n510_n100# a_n720_n100# 0.03fF
C1403 a_n392_n100# a_n812_n100# 0.02fF
C1404 a_n300_n100# a_n930_n100# 0.01fF
C1405 a_n182_n100# a_n1022_n100# 0.01fF
C1406 a_n90_n100# a_n1140_n100# 0.01fF
C1407 a_n3750_n632# a_n3238_n632# 0.01fF
C1408 a_n4078_n632# a_n2910_n632# 0.01fF
C1409 a_n4170_n632# a_n2818_n632# 0.00fF
C1410 a_n3868_n632# a_n3120_n632# 0.01fF
C1411 a_n3960_n632# a_n3028_n632# 0.01fF
C1412 a_4110_n100# a_4062_n197# 0.00fF
C1413 a_n3028_n632# a_n1558_n632# 0.00fF
C1414 a_n2910_n632# a_n1650_n632# 0.00fF
C1415 a_n2818_n632# a_n1768_n632# 0.01fF
C1416 a_2850_n100# a_2804_n729# 0.00fF
C1417 a_2010_n100# a_658_n100# 0.00fF
C1418 a_n810_n632# a_n2280_n632# 0.00fF
C1419 a_1500_n632# a_2760_n632# 0.00fF
C1420 a_1920_n632# a_2340_n632# 0.02fF
C1421 a_2012_n632# a_2222_n632# 0.03fF
C1422 a_1592_n632# a_2642_n632# 0.01fF
C1423 a_1382_n632# a_2852_n632# 0.00fF
C1424 a_1710_n632# a_2550_n632# 0.01fF
C1425 a_1802_n632# a_2432_n632# 0.01fF
C1426 a_n1440_n632# a_n1442_n100# 0.00fF
C1427 a_122_n632# a_n390_n632# 0.01fF
C1428 a_962_n632# a_2130_n632# 0.01fF
C1429 a_n90_n100# a_448_n100# 0.01fF
C1430 a_n1606_n401# a_n1650_n632# 0.00fF
C1431 a_240_n632# a_870_n632# 0.01fF
C1432 a_122_n632# a_962_n632# 0.01fF
C1433 a_332_n632# a_752_n632# 0.02fF
C1434 a_450_n632# a_660_n632# 0.03fF
C1435 a_n2400_n100# a_n3122_n100# 0.01fF
C1436 a_n2190_n100# a_n3332_n100# 0.01fF
C1437 a_n2282_n100# a_n3240_n100# 0.01fF
C1438 a_282_n197# a_n138_n197# 0.01fF
C1439 a_4112_n632# w_n4520_n851# 0.14fF
C1440 w_n4520_n851# a_3434_n401# 0.09fF
C1441 a_n3658_n632# a_n3540_n632# 0.07fF
C1442 a_660_n632# a_702_n197# 0.00fF
C1443 a_3642_n197# a_3598_n100# 0.00fF
C1444 a_494_n401# a_n556_n729# 0.00fF
C1445 a_332_n632# a_n1138_n632# 0.00fF
C1446 w_n4520_n851# a_n3870_n100# 0.05fF
C1447 a_n2820_n100# a_n2818_n632# 0.00fF
C1448 a_3852_131# a_3808_n100# 0.00fF
C1449 a_2128_n100# a_2172_131# 0.00fF
C1450 a_n2610_n100# a_n1350_n100# 0.00fF
C1451 a_n2702_n100# a_n1232_n100# 0.00fF
C1452 a_n2492_n100# a_n1442_n100# 0.01fF
C1453 a_n2490_n632# a_n2188_n632# 0.02fF
C1454 a_n2608_n632# a_n2070_n632# 0.01fF
C1455 a_n2398_n632# a_n2280_n632# 0.07fF
C1456 a_n2700_n632# a_n1978_n632# 0.01fF
C1457 a_n3916_n729# a_n3496_n729# 0.01fF
C1458 a_2340_n632# a_2642_n632# 0.02fF
C1459 a_2130_n632# a_2852_n632# 0.01fF
C1460 a_2222_n632# a_2760_n632# 0.01fF
C1461 a_2432_n632# a_2550_n632# 0.07fF
C1462 a_752_n632# a_n508_n632# 0.00fF
C1463 a_752_n632# a_2012_n632# 0.00fF
C1464 a_n2868_131# a_n1608_131# 0.00fF
C1465 a_n4126_n401# a_n3916_n729# 0.00fF
C1466 a_n182_n100# a_1078_n100# 0.00fF
C1467 a_n300_n100# a_1170_n100# 0.00fF
C1468 a_28_n100# a_n1350_n100# 0.00fF
C1469 a_3062_n632# a_3482_n632# 0.02fF
C1470 a_3180_n632# a_3390_n632# 0.03fF
C1471 a_n3752_n100# a_n3450_n100# 0.02fF
C1472 a_2220_n100# a_2850_n100# 0.01fF
C1473 a_2128_n100# a_2968_n100# 0.01fF
C1474 a_2010_n100# a_3060_n100# 0.01fF
C1475 a_1918_n100# a_3178_n100# 0.00fF
C1476 a_n3660_n100# a_n3542_n100# 0.07fF
C1477 a_n1020_n632# a_n976_n729# 0.00fF
C1478 a_2758_n100# a_3900_n100# 0.01fF
C1479 a_3178_n100# a_3480_n100# 0.02fF
C1480 a_3060_n100# a_3598_n100# 0.01fF
C1481 a_2968_n100# a_3690_n100# 0.01fF
C1482 a_2850_n100# a_3808_n100# 0.01fF
C1483 a_1800_n100# a_750_n100# 0.01fF
C1484 a_2640_n100# a_4018_n100# 0.00fF
C1485 a_2548_n100# a_4110_n100# 0.00fF
C1486 a_1380_n100# a_n182_n100# 0.00fF
C1487 w_n4520_n851# a_3222_n197# 0.10fF
C1488 a_n180_n632# a_n1440_n632# 0.00fF
C1489 a_n390_n632# a_n1230_n632# 0.01fF
C1490 a_n600_n632# a_n1020_n632# 0.02fF
C1491 a_n88_n632# a_n1558_n632# 0.00fF
C1492 a_n298_n632# a_n1348_n632# 0.01fF
C1493 a_n718_n632# a_n928_n632# 0.03fF
C1494 a_n508_n632# a_n1138_n632# 0.01fF
C1495 a_240_n632# a_n600_n632# 0.01fF
C1496 a_3600_n632# a_3644_n729# 0.00fF
C1497 a_n300_n100# a_540_n100# 0.01fF
C1498 a_912_131# a_868_n100# 0.00fF
C1499 a_n2190_n100# w_n4520_n851# 0.02fF
C1500 w_n4520_n851# a_2384_n729# 0.12fF
C1501 w_n4520_n851# a_2172_131# 0.12fF
C1502 a_3012_131# a_3432_131# 0.01fF
C1503 a_1592_n632# w_n4520_n851# 0.01fF
C1504 a_n4170_n632# a_n3960_n632# 0.03fF
C1505 a_2760_n632# a_3810_n632# 0.01fF
C1506 a_2970_n632# a_3600_n632# 0.01fF
C1507 a_2642_n632# a_3902_n632# 0.00fF
C1508 a_2852_n632# a_3692_n632# 0.01fF
C1509 a_2220_n100# a_2222_n632# 0.00fF
C1510 a_n2400_n100# a_n1442_n100# 0.01fF
C1511 a_n1768_n632# a_n1558_n632# 0.03fF
C1512 a_n2400_n100# a_n2446_n401# 0.00fF
C1513 a_2968_n100# w_n4520_n851# 0.03fF
C1514 a_n1980_n100# a_n3542_n100# 0.00fF
C1515 a_n2072_n100# a_n3450_n100# 0.00fF
C1516 a_1080_n632# a_1078_n100# 0.00fF
C1517 a_n88_n632# a_30_n632# 0.07fF
C1518 w_n4520_n851# a_n602_n100# 0.02fF
C1519 a_n2188_n632# a_n1020_n632# 0.01fF
C1520 a_n2280_n632# a_n928_n632# 0.00fF
C1521 a_n1860_n632# a_n1348_n632# 0.01fF
C1522 a_870_n632# a_n718_n632# 0.00fF
C1523 a_n1978_n632# a_n1230_n632# 0.01fF
C1524 a_n2070_n632# a_n1138_n632# 0.01fF
C1525 a_n2238_n197# a_n3078_n197# 0.01fF
C1526 a_870_n632# a_1802_n632# 0.01fF
C1527 a_868_n100# a_1288_n100# 0.02fF
C1528 a_2548_n100# a_960_n100# 0.00fF
C1529 a_n1188_131# a_n138_n197# 0.00fF
C1530 a_2338_n100# a_2548_n100# 0.03fF
C1531 a_n2238_n197# a_n768_131# 0.00fF
C1532 a_120_n100# a_72_131# 0.00fF
C1533 a_912_131# a_n138_n197# 0.00fF
C1534 a_330_n100# a_n602_n100# 0.01fF
C1535 a_74_n401# a_n1396_n729# 0.00fF
C1536 a_n346_n401# a_n1606_n401# 0.00fF
C1537 a_n1442_n100# a_n812_n100# 0.01fF
C1538 a_n1232_n100# a_n1022_n100# 0.03fF
C1539 a_n1350_n100# a_n930_n100# 0.02fF
C1540 a_1590_n100# a_868_n100# 0.01fF
C1541 a_n1186_n401# a_n1140_n100# 0.00fF
C1542 a_2802_n197# a_1752_131# 0.00fF
C1543 w_n4520_n851# a_n2490_n632# 0.01fF
C1544 a_n2868_131# a_n3918_n197# 0.00fF
C1545 w_n4520_n851# a_2340_n632# 0.01fF
C1546 a_3224_n729# a_3434_n401# 0.00fF
C1547 a_2804_n729# a_3854_n401# 0.00fF
C1548 a_332_n632# a_n810_n632# 0.01fF
C1549 a_n1606_n401# a_n766_n401# 0.01fF
C1550 a_332_n632# a_1710_n632# 0.00fF
C1551 a_n90_n100# a_28_n100# 0.07fF
C1552 a_n510_n100# a_658_n100# 0.01fF
C1553 a_1918_n100# a_2010_n100# 0.09fF
C1554 a_1800_n100# a_2128_n100# 0.02fF
C1555 a_1708_n100# a_2220_n100# 0.01fF
C1556 a_3012_131# a_1962_n197# 0.00fF
C1557 a_492_131# a_n768_131# 0.00fF
C1558 a_3810_n632# a_3808_n100# 0.00fF
C1559 a_2220_n100# a_3270_n100# 0.01fF
C1560 a_2128_n100# a_3388_n100# 0.00fF
C1561 a_2010_n100# a_3480_n100# 0.00fF
C1562 a_n4170_n632# a_n4172_n100# 0.00fF
C1563 a_448_n100# a_n1140_n100# 0.00fF
C1564 a_n3120_n632# a_n2700_n632# 0.02fF
C1565 a_n3658_n632# a_n2188_n632# 0.00fF
C1566 a_n3238_n632# a_n2608_n632# 0.01fF
C1567 a_n3330_n632# a_n2490_n632# 0.01fF
C1568 a_n3540_n632# a_n2280_n632# 0.00fF
C1569 a_n3448_n632# a_n2398_n632# 0.01fF
C1570 a_3480_n100# a_3598_n100# 0.07fF
C1571 a_3388_n100# a_3690_n100# 0.02fF
C1572 a_3270_n100# a_3808_n100# 0.01fF
C1573 a_n2282_n100# a_n1560_n100# 0.01fF
C1574 a_n2190_n100# a_n1652_n100# 0.01fF
C1575 a_n1980_n100# a_n1862_n100# 0.07fF
C1576 a_n2072_n100# a_n1770_n100# 0.02fF
C1577 a_4020_n632# a_2970_n632# 0.01fF
C1578 a_4112_n632# a_2852_n632# 0.00fF
C1579 a_1754_n401# a_1964_n729# 0.00fF
C1580 a_2594_n401# a_1124_n729# 0.00fF
C1581 a_2174_n401# a_1544_n729# 0.00fF
C1582 a_1334_n401# a_2384_n729# 0.00fF
C1583 a_n2028_131# a_n1188_131# 0.01fF
C1584 a_n2448_131# a_n1608_131# 0.01fF
C1585 a_n810_n632# a_n508_n632# 0.02fF
C1586 a_n718_n632# a_n600_n632# 0.07fF
C1587 a_1290_n632# a_n88_n632# 0.00fF
C1588 a_1382_n632# a_n180_n632# 0.00fF
C1589 a_1710_n632# a_2012_n632# 0.02fF
C1590 a_1802_n632# a_1920_n632# 0.07fF
C1591 a_3222_n197# a_3224_n729# 0.01fF
C1592 a_n2072_n100# a_n510_n100# 0.00fF
C1593 a_n1652_n100# a_n602_n100# 0.01fF
C1594 a_2640_n100# a_2594_n401# 0.00fF
C1595 a_n1560_n100# a_n720_n100# 0.01fF
C1596 a_n2820_n100# a_n2610_n100# 0.03fF
C1597 a_962_n632# a_1592_n632# 0.01fF
C1598 a_n2912_n100# a_n2492_n100# 0.02fF
C1599 a_1172_n632# a_1382_n632# 0.03fF
C1600 a_960_n100# a_1078_n100# 0.07fF
C1601 a_1800_n100# w_n4520_n851# 0.02fF
C1602 a_2338_n100# a_1078_n100# 0.00fF
C1603 w_n4520_n851# a_3902_n632# 0.06fF
C1604 w_n4520_n851# a_3388_n100# 0.03fF
C1605 a_n3918_n197# a_n3916_n729# 0.01fF
C1606 a_n2912_n100# a_n4080_n100# 0.01fF
C1607 a_n3122_n100# a_n3870_n100# 0.01fF
C1608 a_n3240_n100# a_n3752_n100# 0.01fF
C1609 a_n2820_n100# a_n4172_n100# 0.00fF
C1610 a_n3030_n100# a_n3962_n100# 0.01fF
C1611 a_n3332_n100# a_n3660_n100# 0.02fF
C1612 a_n2868_131# w_n4520_n851# 0.12fF
C1613 a_3224_n729# a_2384_n729# 0.01fF
C1614 a_n978_n197# a_n1020_n632# 0.00fF
C1615 a_n766_n401# a_n768_131# 0.01fF
C1616 a_1800_n100# a_330_n100# 0.00fF
C1617 a_1380_n100# a_960_n100# 0.02fF
C1618 a_1380_n100# a_2338_n100# 0.01fF
C1619 a_660_n632# a_n88_n632# 0.01fF
C1620 a_542_n632# a_30_n632# 0.01fF
C1621 a_4020_n632# a_4018_n100# 0.00fF
C1622 w_n4520_n851# a_n1020_n632# 0.01fF
C1623 a_450_n632# a_1500_n632# 0.01fF
C1624 a_240_n632# w_n4520_n851# 0.01fF
C1625 a_n300_n100# a_120_n100# 0.02fF
C1626 a_n2072_n100# a_n2070_n632# 0.00fF
C1627 a_n392_n100# a_n602_n100# 0.03fF
C1628 a_n300_n100# a_n720_n100# 0.02fF
C1629 a_n182_n100# a_n812_n100# 0.01fF
C1630 a_n90_n100# a_n930_n100# 0.01fF
C1631 a_n3750_n632# a_n3028_n632# 0.01fF
C1632 a_n3960_n632# a_n2818_n632# 0.01fF
C1633 a_n3868_n632# a_n2910_n632# 0.01fF
C1634 a_2174_n401# a_2130_n632# 0.00fF
C1635 a_n2910_n632# a_n1440_n632# 0.00fF
C1636 a_n2818_n632# a_n1558_n632# 0.00fF
C1637 a_2220_n100# a_658_n100# 0.00fF
C1638 a_n718_n632# a_n2188_n632# 0.00fF
C1639 a_n810_n632# a_n2070_n632# 0.00fF
C1640 a_1500_n632# a_2970_n632# 0.00fF
C1641 a_2012_n632# a_2432_n632# 0.02fF
C1642 a_1802_n632# a_2642_n632# 0.01fF
C1643 a_1920_n632# a_2550_n632# 0.01fF
C1644 a_1592_n632# a_2852_n632# 0.00fF
C1645 a_1710_n632# a_2760_n632# 0.01fF
C1646 a_n1348_n632# a_n1350_n100# 0.00fF
C1647 a_122_n632# a_n180_n632# 0.02fF
C1648 a_n1348_n632# a_n1396_n729# 0.00fF
C1649 a_962_n632# a_2340_n632# 0.00fF
C1650 a_1172_n632# a_2130_n632# 0.01fF
C1651 a_704_n729# a_1124_n729# 0.01fF
C1652 a_122_n632# a_1172_n632# 0.01fF
C1653 a_2130_n632# a_3062_n632# 0.01fF
C1654 a_n2282_n100# a_n3030_n100# 0.01fF
C1655 a_n2190_n100# a_n3122_n100# 0.01fF
C1656 a_n1980_n100# a_n3332_n100# 0.00fF
C1657 a_n2400_n100# a_n2912_n100# 0.01fF
C1658 a_n2072_n100# a_n3240_n100# 0.01fF
C1659 w_n4520_n851# a_n3658_n632# 0.04fF
C1660 a_494_n401# a_1754_n401# 0.00fF
C1661 w_n4520_n851# a_n3916_n729# 0.13fF
C1662 a_n3540_n632# a_n3448_n632# 0.09fF
C1663 a_n3658_n632# a_n3330_n632# 0.02fF
C1664 a_1080_n632# a_1382_n632# 0.02fF
C1665 a_74_n401# a_704_n729# 0.00fF
C1666 a_494_n401# a_284_n729# 0.00fF
C1667 a_1708_n100# a_1752_131# 0.00fF
C1668 a_332_n632# a_n928_n632# 0.00fF
C1669 a_n1608_131# a_n348_131# 0.00fF
C1670 a_n2448_131# a_n3918_n197# 0.00fF
C1671 a_n3288_131# a_n1818_n197# 0.00fF
C1672 w_n4520_n851# a_n3660_n100# 0.04fF
C1673 a_n3448_n632# a_n3496_n729# 0.00fF
C1674 a_1542_n197# a_492_131# 0.00fF
C1675 a_660_n632# a_704_n729# 0.00fF
C1676 a_1122_n197# a_1962_n197# 0.01fF
C1677 a_n2398_n632# a_n2070_n632# 0.02fF
C1678 a_n2492_n100# a_n1232_n100# 0.00fF
C1679 a_n2608_n632# a_n1860_n632# 0.01fF
C1680 a_n2490_n632# a_n1978_n632# 0.01fF
C1681 a_n2610_n100# a_n1140_n100# 0.00fF
C1682 a_n2280_n632# a_n2188_n632# 0.09fF
C1683 a_n3496_n729# a_n3076_n729# 0.01fF
C1684 a_n3916_n729# a_n2656_n729# 0.00fF
C1685 a_2222_n632# a_2970_n632# 0.01fF
C1686 a_2432_n632# a_2760_n632# 0.02fF
C1687 a_752_n632# a_n298_n632# 0.01fF
C1688 a_2340_n632# a_2852_n632# 0.01fF
C1689 a_2550_n632# a_2642_n632# 0.09fF
C1690 a_n3286_n401# a_n3916_n729# 0.00fF
C1691 a_n4126_n401# a_n3076_n729# 0.00fF
C1692 a_n3706_n401# a_n3496_n729# 0.00fF
C1693 a_n90_n100# a_1170_n100# 0.00fF
C1694 a_n182_n100# a_1288_n100# 0.00fF
C1695 a_542_n632# a_1290_n632# 0.01fF
C1696 a_n510_n100# a_238_n100# 0.01fF
C1697 a_n3496_n729# a_n3450_n100# 0.00fF
C1698 a_n4126_n401# a_n3706_n401# 0.01fF
C1699 a_868_n100# a_n602_n100# 0.00fF
C1700 a_28_n100# a_n1140_n100# 0.01fF
C1701 a_3180_n632# a_3600_n632# 0.02fF
C1702 a_3062_n632# a_3692_n632# 0.01fF
C1703 a_3272_n632# a_3482_n632# 0.03fF
C1704 a_1122_n197# a_1124_n729# 0.01fF
C1705 a_n3542_n100# a_n3450_n100# 0.09fF
C1706 a_2220_n100# a_3060_n100# 0.01fF
C1707 a_2128_n100# a_3178_n100# 0.01fF
C1708 a_450_n632# a_494_n401# 0.00fF
C1709 a_2010_n100# a_750_n100# 0.00fF
C1710 a_2758_n100# a_4110_n100# 0.00fF
C1711 a_3178_n100# a_3690_n100# 0.01fF
C1712 a_3060_n100# a_3808_n100# 0.01fF
C1713 a_2968_n100# a_3900_n100# 0.01fF
C1714 a_2850_n100# a_4018_n100# 0.01fF
C1715 a_n4128_131# a_n3078_n197# 0.00fF
C1716 a_1498_n100# a_n90_n100# 0.00fF
C1717 a_n390_n632# a_n1020_n632# 0.01fF
C1718 a_n88_n632# a_n1348_n632# 0.00fF
C1719 a_n298_n632# a_n1138_n632# 0.01fF
C1720 a_n180_n632# a_n1230_n632# 0.01fF
C1721 a_n508_n632# a_n928_n632# 0.02fF
C1722 a_240_n632# a_n390_n632# 0.01fF
C1723 a_1080_n632# a_2130_n632# 0.01fF
C1724 a_n1608_131# a_n1398_n197# 0.00fF
C1725 a_240_n632# a_962_n632# 0.01fF
C1726 a_122_n632# a_1080_n632# 0.01fF
C1727 a_28_n100# a_448_n100# 0.02fF
C1728 a_n90_n100# a_540_n100# 0.01fF
C1729 a_332_n632# a_870_n632# 0.01fF
C1730 a_450_n632# a_752_n632# 0.02fF
C1731 a_542_n632# a_660_n632# 0.07fF
C1732 a_n1980_n100# w_n4520_n851# 0.02fF
C1733 a_n2448_131# a_n978_n197# 0.00fF
C1734 a_2338_n100# a_2382_n197# 0.00fF
C1735 a_n2448_131# w_n4520_n851# 0.12fF
C1736 a_n718_n632# w_n4520_n851# 0.01fF
C1737 a_n4078_n632# a_n3868_n632# 0.03fF
C1738 a_1802_n632# w_n4520_n851# 0.01fF
C1739 a_n4170_n632# a_n3750_n632# 0.02fF
C1740 a_2852_n632# a_3902_n632# 0.01fF
C1741 a_2970_n632# a_3810_n632# 0.01fF
C1742 a_914_n401# a_n556_n729# 0.00fF
C1743 a_n2190_n100# a_n1442_n100# 0.01fF
C1744 a_n2282_n100# a_n1350_n100# 0.01fF
C1745 a_n2400_n100# a_n1232_n100# 0.01fF
C1746 a_450_n632# a_n1138_n632# 0.00fF
C1747 a_n1650_n632# a_n1440_n632# 0.03fF
C1748 a_n1768_n632# a_n1348_n632# 0.02fF
C1749 a_2174_n401# a_3434_n401# 0.00fF
C1750 a_3178_n100# w_n4520_n851# 0.03fF
C1751 a_3432_131# a_3390_n632# 0.00fF
C1752 a_282_n197# a_n768_131# 0.00fF
C1753 a_n1862_n100# a_n3450_n100# 0.00fF
C1754 a_n1978_n632# a_n1020_n632# 0.01fF
C1755 a_870_n632# a_n508_n632# 0.00fF
C1756 a_n2070_n632# a_n928_n632# 0.01fF
C1757 a_n1860_n632# a_n1138_n632# 0.01fF
C1758 a_870_n632# a_2012_n632# 0.01fF
C1759 a_4020_n632# a_3180_n632# 0.01fF
C1760 a_4112_n632# a_3062_n632# 0.01fF
C1761 a_2430_n100# a_2640_n100# 0.03fF
C1762 a_2338_n100# a_2758_n100# 0.02fF
C1763 a_120_n100# a_n1350_n100# 0.00fF
C1764 a_n1350_n100# a_n720_n100# 0.01fF
C1765 a_n1232_n100# a_n812_n100# 0.02fF
C1766 a_n1140_n100# a_n930_n100# 0.03fF
C1767 a_74_n401# a_n1186_n401# 0.00fF
C1768 a_n346_n401# a_n766_n401# 0.01fF
C1769 a_n1442_n100# a_n602_n100# 0.01fF
C1770 a_1800_n100# a_868_n100# 0.01fF
C1771 a_4112_n632# a_4064_n729# 0.00fF
C1772 w_n4520_n851# a_n2280_n632# 0.01fF
C1773 a_30_n632# a_n1558_n632# 0.00fF
C1774 w_n4520_n851# a_2550_n632# 0.01fF
C1775 a_3644_n729# a_3854_n401# 0.00fF
C1776 a_4064_n729# a_3434_n401# 0.00fF
C1777 a_332_n632# a_n600_n632# 0.01fF
C1778 a_332_n632# a_1920_n632# 0.00fF
C1779 a_912_131# a_960_n100# 0.00fF
C1780 a_n300_n100# a_658_n100# 0.01fF
C1781 a_3012_131# a_2802_n197# 0.00fF
C1782 a_2010_n100# a_2128_n100# 0.07fF
C1783 a_1918_n100# a_2220_n100# 0.02fF
C1784 a_2220_n100# a_3480_n100# 0.00fF
C1785 a_2128_n100# a_3598_n100# 0.00fF
C1786 a_3902_n632# a_3900_n100# 0.00fF
C1787 a_n4078_n632# a_n4080_n100# 0.00fF
C1788 a_n3028_n632# a_n2608_n632# 0.02fF
C1789 a_448_n100# a_n930_n100# 0.00fF
C1790 a_3598_n100# a_3690_n100# 0.09fF
C1791 a_3480_n100# a_3808_n100# 0.02fF
C1792 a_3388_n100# a_3900_n100# 0.01fF
C1793 a_3270_n100# a_4018_n100# 0.01fF
C1794 a_n3448_n632# a_n2188_n632# 0.00fF
C1795 a_n3540_n632# a_n2070_n632# 0.00fF
C1796 a_n3238_n632# a_n2398_n632# 0.01fF
C1797 a_n3330_n632# a_n2280_n632# 0.01fF
C1798 a_n2910_n632# a_n2700_n632# 0.03fF
C1799 a_n3120_n632# a_n2490_n632# 0.01fF
C1800 a_n1188_131# a_n1232_n100# 0.00fF
C1801 a_1122_n197# a_1170_n100# 0.00fF
C1802 w_n4520_n851# a_2592_131# 0.12fF
C1803 a_n1862_n100# a_n1770_n100# 0.09fF
C1804 a_n1980_n100# a_n1652_n100# 0.02fF
C1805 a_n2072_n100# a_n1560_n100# 0.01fF
C1806 a_n3708_131# a_n3078_n197# 0.00fF
C1807 a_542_n632# a_540_n100# 0.00fF
C1808 a_3012_131# a_3852_131# 0.01fF
C1809 a_3014_n401# a_1544_n729# 0.00fF
C1810 a_1710_n632# a_1752_131# 0.00fF
C1811 a_2594_n401# a_1964_n729# 0.00fF
C1812 a_2174_n401# a_2384_n729# 0.00fF
C1813 a_2172_131# a_2174_n401# 0.01fF
C1814 a_n2446_n401# a_n2490_n632# 0.00fF
C1815 a_n348_131# a_n978_n197# 0.00fF
C1816 a_n976_n729# a_n556_n729# 0.01fF
C1817 a_1710_n632# a_1754_n401# 0.00fF
C1818 a_n600_n632# a_n556_n729# 0.00fF
C1819 a_702_n197# a_658_n100# 0.00fF
C1820 w_n4520_n851# a_n348_131# 0.12fF
C1821 a_n810_n632# a_n298_n632# 0.01fF
C1822 a_n718_n632# a_n390_n632# 0.02fF
C1823 a_n600_n632# a_n508_n632# 0.09fF
C1824 a_1500_n632# a_n88_n632# 0.00fF
C1825 a_1920_n632# a_2012_n632# 0.09fF
C1826 a_3642_n197# a_3644_n729# 0.01fF
C1827 a_n1980_n100# a_n392_n100# 0.00fF
C1828 a_n1862_n100# a_n510_n100# 0.00fF
C1829 a_n2702_n100# a_n2492_n100# 0.03fF
C1830 a_1172_n632# a_1592_n632# 0.02fF
C1831 a_962_n632# a_1802_n632# 0.01fF
C1832 a_2010_n100# w_n4520_n851# 0.02fF
C1833 a_960_n100# a_1288_n100# 0.02fF
C1834 a_2338_n100# a_1288_n100# 0.01fF
C1835 a_2430_n100# a_1170_n100# 0.00fF
C1836 a_2548_n100# a_1078_n100# 0.00fF
C1837 w_n4520_n851# a_3598_n100# 0.04fF
C1838 a_1592_n632# a_3062_n632# 0.00fF
C1839 a_n768_131# a_n812_n100# 0.00fF
C1840 a_n2610_n100# a_n4172_n100# 0.00fF
C1841 a_n2702_n100# a_n4080_n100# 0.00fF
C1842 a_n2820_n100# a_n3962_n100# 0.01fF
C1843 a_n3332_n100# a_n3450_n100# 0.07fF
C1844 a_n3122_n100# a_n3660_n100# 0.01fF
C1845 a_n3240_n100# a_n3542_n100# 0.02fF
C1846 a_n3030_n100# a_n3752_n100# 0.01fF
C1847 a_30_n632# a_28_n100# 0.00fF
C1848 a_n2912_n100# a_n3870_n100# 0.01fF
C1849 a_1590_n100# a_960_n100# 0.01fF
C1850 a_1590_n100# a_2338_n100# 0.01fF
C1851 a_1498_n100# a_2430_n100# 0.01fF
C1852 a_1380_n100# a_2548_n100# 0.01fF
C1853 a_4112_n632# a_4110_n100# 0.00fF
C1854 a_450_n632# a_n810_n632# 0.00fF
C1855 a_450_n632# a_1710_n632# 0.00fF
C1856 a_448_n100# a_1170_n100# 0.01fF
C1857 a_n90_n100# a_120_n100# 0.03fF
C1858 a_n1398_n197# a_n978_n197# 0.01fF
C1859 a_n1980_n100# a_n1978_n632# 0.00fF
C1860 a_n510_n100# a_750_n100# 0.00fF
C1861 a_n1188_131# a_n768_131# 0.01fF
C1862 a_3432_131# a_1962_n197# 0.00fF
C1863 a_n182_n100# a_n602_n100# 0.02fF
C1864 a_n90_n100# a_n720_n100# 0.01fF
C1865 a_n3750_n632# a_n2818_n632# 0.01fF
C1866 a_n2818_n632# a_n1348_n632# 0.00fF
C1867 w_n4520_n851# a_n1398_n197# 0.10fF
C1868 a_282_n197# a_492_131# 0.00fF
C1869 a_n600_n632# a_n2070_n632# 0.00fF
C1870 a_n810_n632# a_n1860_n632# 0.01fF
C1871 a_n718_n632# a_n1978_n632# 0.00fF
C1872 a_1498_n100# a_448_n100# 0.01fF
C1873 a_282_n197# a_1542_n197# 0.00fF
C1874 a_1920_n632# a_2760_n632# 0.01fF
C1875 a_1710_n632# a_2970_n632# 0.00fF
C1876 a_n1230_n632# a_n1232_n100# 0.00fF
C1877 a_2012_n632# a_2642_n632# 0.01fF
C1878 a_1802_n632# a_2852_n632# 0.01fF
C1879 w_n4520_n851# a_1332_131# 0.12fF
C1880 a_962_n632# a_2550_n632# 0.00fF
C1881 a_1172_n632# a_2340_n632# 0.01fF
C1882 a_n2868_131# a_n2028_131# 0.01fF
C1883 a_704_n729# a_1964_n729# 0.00fF
C1884 a_448_n100# a_540_n100# 0.09fF
C1885 a_2340_n632# a_3062_n632# 0.01fF
C1886 a_2222_n632# a_3180_n632# 0.01fF
C1887 a_2130_n632# a_3272_n632# 0.01fF
C1888 a_n1980_n100# a_n3122_n100# 0.01fF
C1889 a_n2072_n100# a_n3030_n100# 0.01fF
C1890 a_n1862_n100# a_n3240_n100# 0.00fF
C1891 a_n2282_n100# a_n2820_n100# 0.01fF
C1892 a_n2400_n100# a_n2702_n100# 0.02fF
C1893 a_n1770_n100# a_n3332_n100# 0.00fF
C1894 a_n2190_n100# a_n2912_n100# 0.01fF
C1895 w_n4520_n851# a_n3448_n632# 0.03fF
C1896 a_1290_n632# a_30_n632# 0.00fF
C1897 a_n3708_131# a_n2238_n197# 0.00fF
C1898 w_n4520_n851# a_n3076_n729# 0.12fF
C1899 a_n3540_n632# a_n3238_n632# 0.02fF
C1900 a_n4078_n632# a_n2700_n632# 0.00fF
C1901 a_n3448_n632# a_n3330_n632# 0.07fF
C1902 a_n3658_n632# a_n3120_n632# 0.01fF
C1903 a_n4170_n632# a_n2608_n632# 0.00fF
C1904 a_1080_n632# a_1592_n632# 0.01fF
C1905 w_n4520_n851# a_n3706_n401# 0.10fF
C1906 a_n2608_n632# a_n1768_n632# 0.01fF
C1907 a_n2700_n632# a_n1650_n632# 0.01fF
C1908 w_n4520_n851# a_n3450_n100# 0.03fF
C1909 a_30_n632# a_74_n401# 0.00fF
C1910 a_n390_n632# a_n348_131# 0.00fF
C1911 a_1380_n100# a_1078_n100# 0.02fF
C1912 a_n2492_n100# a_n1022_n100# 0.00fF
C1913 a_n2398_n632# a_n1860_n632# 0.01fF
C1914 a_n2280_n632# a_n1978_n632# 0.02fF
C1915 a_1542_n197# a_2382_n197# 0.01fF
C1916 a_n2188_n632# a_n2070_n632# 0.07fF
C1917 a_n3076_n729# a_n2656_n729# 0.01fF
C1918 a_n3496_n729# a_n2236_n729# 0.00fF
C1919 a_2642_n632# a_2760_n632# 0.07fF
C1920 a_2432_n632# a_2970_n632# 0.01fF
C1921 a_2550_n632# a_2852_n632# 0.02fF
C1922 a_752_n632# a_n88_n632# 0.01fF
C1923 a_660_n632# a_30_n632# 0.01fF
C1924 a_n3286_n401# a_n3076_n729# 0.00fF
C1925 a_n3706_n401# a_n2656_n729# 0.00fF
C1926 a_n2866_n401# a_n3496_n729# 0.00fF
C1927 a_n2446_n401# a_n3916_n729# 0.00fF
C1928 a_332_n632# w_n4520_n851# 0.01fF
C1929 a_542_n632# a_1500_n632# 0.01fF
C1930 a_n300_n100# a_238_n100# 0.01fF
C1931 a_n4126_n401# a_n2866_n401# 0.00fF
C1932 a_n3706_n401# a_n3286_n401# 0.01fF
C1933 a_n392_n100# a_n348_131# 0.00fF
C1934 a_28_n100# a_n930_n100# 0.01fF
C1935 a_3390_n632# a_3600_n632# 0.03fF
C1936 a_3062_n632# a_3902_n632# 0.01fF
C1937 a_3180_n632# a_3810_n632# 0.01fF
C1938 a_3272_n632# a_3692_n632# 0.02fF
C1939 a_1542_n197# a_1544_n729# 0.01fF
C1940 a_332_n632# a_330_n100# 0.00fF
C1941 a_2220_n100# a_750_n100# 0.00fF
C1942 a_3178_n100# a_3900_n100# 0.01fF
C1943 a_3060_n100# a_4018_n100# 0.01fF
C1944 a_2968_n100# a_4110_n100# 0.01fF
C1945 a_n298_n632# a_n928_n632# 0.01fF
C1946 a_n180_n632# a_n1020_n632# 0.01fF
C1947 a_n88_n632# a_n1138_n632# 0.01fF
C1948 a_n2702_n100# a_n2700_n632# 0.00fF
C1949 a_240_n632# a_n180_n632# 0.02fF
C1950 a_1080_n632# a_2340_n632# 0.00fF
C1951 a_n1608_131# a_n558_n197# 0.00fF
C1952 a_240_n632# a_1172_n632# 0.01fF
C1953 a_n2238_n197# a_n1188_131# 0.00fF
C1954 a_n1770_n100# w_n4520_n851# 0.02fF
C1955 a_n600_n632# a_n558_n197# 0.00fF
C1956 a_1334_n401# a_1332_131# 0.01fF
C1957 w_n4520_n851# a_n556_n729# 0.12fF
C1958 a_n508_n632# w_n4520_n851# 0.01fF
C1959 a_2012_n632# w_n4520_n851# 0.01fF
C1960 a_914_n401# a_1754_n401# 0.01fF
C1961 a_n3960_n632# a_n3750_n632# 0.03fF
C1962 a_74_n401# a_1124_n729# 0.00fF
C1963 a_494_n401# a_704_n729# 0.00fF
C1964 a_914_n401# a_284_n729# 0.00fF
C1965 a_n2282_n100# a_n1140_n100# 0.01fF
C1966 a_n2400_n100# a_n1022_n100# 0.00fF
C1967 a_n3332_n100# a_n3240_n100# 0.09fF
C1968 a_n2072_n100# a_n1350_n100# 0.01fF
C1969 a_n2190_n100# a_n1232_n100# 0.01fF
C1970 a_n1980_n100# a_n1442_n100# 0.01fF
C1971 a_450_n632# a_n928_n632# 0.00fF
C1972 a_n1768_n632# a_n1138_n632# 0.01fF
C1973 a_n1558_n632# a_n1348_n632# 0.03fF
C1974 a_n1650_n632# a_n1230_n632# 0.02fF
C1975 a_492_131# a_912_131# 0.01fF
C1976 a_3014_n401# a_3434_n401# 0.01fF
C1977 a_2594_n401# a_3854_n401# 0.00fF
C1978 a_n2236_n729# a_n976_n729# 0.00fF
C1979 a_1542_n197# a_912_131# 0.00fF
C1980 a_n510_n100# w_n4520_n851# 0.02fF
C1981 a_752_n632# a_704_n729# 0.00fF
C1982 a_n2448_131# a_n2446_n401# 0.01fF
C1983 a_n1980_n100# a_n2028_131# 0.00fF
C1984 a_n1860_n632# a_n928_n632# 0.01fF
C1985 a_870_n632# a_n298_n632# 0.01fF
C1986 a_4020_n632# a_3390_n632# 0.01fF
C1987 a_4112_n632# a_3272_n632# 0.01fF
C1988 w_n4520_n851# a_2804_n729# 0.12fF
C1989 a_28_n100# a_1170_n100# 0.01fF
C1990 a_2548_n100# a_2758_n100# 0.03fF
C1991 a_2430_n100# a_2850_n100# 0.02fF
C1992 a_2338_n100# a_2968_n100# 0.01fF
C1993 a_660_n632# a_1290_n632# 0.01fF
C1994 a_n1608_131# a_n2658_n197# 0.00fF
C1995 a_n510_n100# a_330_n100# 0.01fF
C1996 a_960_n100# a_n602_n100# 0.00fF
C1997 a_n2448_131# a_n2028_131# 0.01fF
C1998 a_120_n100# a_n1140_n100# 0.00fF
C1999 a_n2868_131# a_n2912_n100# 0.00fF
C2000 a_n1022_n100# a_n812_n100# 0.03fF
C2001 a_n1140_n100# a_n720_n100# 0.02fF
C2002 a_n1232_n100# a_n602_n100# 0.01fF
C2003 a_542_n632# a_494_n401# 0.00fF
C2004 a_2010_n100# a_868_n100# 0.01fF
C2005 a_1498_n100# a_28_n100# 0.00fF
C2006 w_n4520_n851# a_n2070_n632# 0.01fF
C2007 a_30_n632# a_n1348_n632# 0.00fF
C2008 w_n4520_n851# a_2760_n632# 0.02fF
C2009 a_332_n632# a_n390_n632# 0.01fF
C2010 a_120_n100# a_448_n100# 0.02fF
C2011 a_28_n100# a_540_n100# 0.01fF
C2012 a_n90_n100# a_658_n100# 0.01fF
C2013 a_332_n632# a_962_n632# 0.01fF
C2014 a_2128_n100# a_2220_n100# 0.09fF
C2015 a_450_n632# a_870_n632# 0.02fF
C2016 a_3012_131# a_3642_n197# 0.00fF
C2017 a_542_n632# a_752_n632# 0.03fF
C2018 a_240_n632# a_1080_n632# 0.01fF
C2019 a_2220_n100# a_3690_n100# 0.00fF
C2020 a_n3960_n632# a_n3962_n100# 0.00fF
C2021 a_n3330_n632# a_n2070_n632# 0.00fF
C2022 a_n3120_n632# a_n2280_n632# 0.01fF
C2023 a_n2910_n632# a_n2490_n632# 0.02fF
C2024 a_n2818_n632# a_n2608_n632# 0.03fF
C2025 a_n3028_n632# a_n2398_n632# 0.01fF
C2026 a_n3448_n632# a_n1978_n632# 0.00fF
C2027 a_448_n100# a_n720_n100# 0.01fF
C2028 a_3690_n100# a_3808_n100# 0.07fF
C2029 a_3598_n100# a_3900_n100# 0.02fF
C2030 a_3480_n100# a_4018_n100# 0.01fF
C2031 a_3388_n100# a_4110_n100# 0.01fF
C2032 a_n3238_n632# a_n2188_n632# 0.01fF
C2033 a_n1770_n100# a_n1652_n100# 0.07fF
C2034 a_n1862_n100# a_n1560_n100# 0.02fF
C2035 a_2338_n100# a_2340_n632# 0.00fF
C2036 a_n4128_131# a_n4080_n100# 0.00fF
C2037 a_n1560_n100# a_n1608_131# 0.00fF
C2038 a_n2188_n632# a_n2236_n729# 0.00fF
C2039 a_3014_n401# a_2384_n729# 0.00fF
C2040 a_n3240_n100# w_n4520_n851# 0.03fF
C2041 a_1590_n100# a_1542_n197# 0.00fF
C2042 a_1170_n100# a_1124_n729# 0.00fF
C2043 a_n348_131# a_n138_n197# 0.00fF
C2044 a_n556_n729# a_n136_n729# 0.01fF
C2045 a_n976_n729# a_284_n729# 0.00fF
C2046 a_n600_n632# a_n298_n632# 0.02fF
C2047 a_n508_n632# a_n390_n632# 0.07fF
C2048 a_n810_n632# a_n88_n632# 0.01fF
C2049 a_n718_n632# a_n180_n632# 0.01fF
C2050 a_3060_n100# a_3012_131# 0.00fF
C2051 a_n1862_n100# a_n300_n100# 0.00fF
C2052 a_n1652_n100# a_n510_n100# 0.01fF
C2053 a_n1770_n100# a_n392_n100# 0.00fF
C2054 a_962_n632# a_n508_n632# 0.00fF
C2055 a_1172_n632# a_1802_n632# 0.01fF
C2056 a_962_n632# a_2012_n632# 0.01fF
C2057 a_2220_n100# w_n4520_n851# 0.02fF
C2058 a_2548_n100# a_1288_n100# 0.00fF
C2059 a_2640_n100# a_1170_n100# 0.00fF
C2060 a_n3240_n100# a_n3286_n401# 0.00fF
C2061 w_n4520_n851# a_3808_n100# 0.05fF
C2062 a_1380_n100# a_1382_n632# 0.00fF
C2063 a_1710_n632# a_3180_n632# 0.00fF
C2064 a_1802_n632# a_3062_n632# 0.00fF
C2065 a_n2912_n100# a_n3660_n100# 0.01fF
C2066 a_n3122_n100# a_n3450_n100# 0.02fF
C2067 a_n2820_n100# a_n3752_n100# 0.01fF
C2068 a_n2492_n100# a_n4080_n100# 0.00fF
C2069 a_n3030_n100# a_n3542_n100# 0.01fF
C2070 a_n2702_n100# a_n3870_n100# 0.01fF
C2071 a_n2610_n100# a_n3962_n100# 0.00fF
C2072 a_238_n100# a_n1350_n100# 0.00fF
C2073 a_1334_n401# a_2804_n729# 0.00fF
C2074 a_n4128_131# a_n3708_131# 0.01fF
C2075 a_1800_n100# a_960_n100# 0.01fF
C2076 a_1380_n100# a_2758_n100# 0.00fF
C2077 a_n4172_n100# a_n3962_n100# 0.03fF
C2078 a_1800_n100# a_2338_n100# 0.01fF
C2079 a_1708_n100# a_2430_n100# 0.01fF
C2080 a_1590_n100# a_2548_n100# 0.01fF
C2081 a_1498_n100# a_2640_n100# 0.01fF
C2082 a_2430_n100# a_3270_n100# 0.01fF
C2083 a_2338_n100# a_3388_n100# 0.01fF
C2084 a_n2868_131# a_n2910_n632# 0.00fF
C2085 a_450_n632# a_n600_n632# 0.01fF
C2086 a_n2658_n197# a_n3918_n197# 0.00fF
C2087 a_n810_n632# a_n1768_n632# 0.01fF
C2088 a_450_n632# a_1920_n632# 0.00fF
C2089 a_n978_n197# a_n558_n197# 0.01fF
C2090 a_n1398_n197# a_n138_n197# 0.00fF
C2091 a_n1862_n100# a_n1860_n632# 0.00fF
C2092 a_n300_n100# a_750_n100# 0.01fF
C2093 a_3432_131# a_2802_n197# 0.00fF
C2094 a_n510_n100# a_n392_n100# 0.07fF
C2095 a_540_n100# a_n930_n100# 0.00fF
C2096 a_1332_131# a_n138_n197# 0.00fF
C2097 w_n4520_n851# a_n558_n197# 0.10fF
C2098 a_3432_131# a_3852_131# 0.01fF
C2099 a_n600_n632# a_n1860_n632# 0.00fF
C2100 a_n508_n632# a_n1978_n632# 0.00fF
C2101 a_1708_n100# a_448_n100# 0.00fF
C2102 a_2012_n632# a_2852_n632# 0.01fF
C2103 a_1920_n632# a_2970_n632# 0.01fF
C2104 a_n1138_n632# a_n1140_n100# 0.00fF
C2105 a_1172_n632# a_2550_n632# 0.00fF
C2106 a_n1186_n401# a_n1138_n632# 0.00fF
C2107 a_2804_n729# a_3224_n729# 0.01fF
C2108 a_2222_n632# a_3390_n632# 0.01fF
C2109 a_2130_n632# a_3482_n632# 0.00fF
C2110 a_2432_n632# a_3180_n632# 0.01fF
C2111 a_2550_n632# a_3062_n632# 0.01fF
C2112 a_2340_n632# a_3272_n632# 0.01fF
C2113 a_72_131# a_n978_n197# 0.00fF
C2114 a_3222_n197# a_4062_n197# 0.01fF
C2115 a_n2190_n100# a_n2702_n100# 0.01fF
C2116 a_n2282_n100# a_n2610_n100# 0.02fF
C2117 a_n1770_n100# a_n3122_n100# 0.00fF
C2118 a_n1862_n100# a_n3030_n100# 0.01fF
C2119 a_n1980_n100# a_n2912_n100# 0.01fF
C2120 a_n2072_n100# a_n2820_n100# 0.01fF
C2121 a_n1652_n100# a_n3240_n100# 0.00fF
C2122 a_n2400_n100# a_n2492_n100# 0.09fF
C2123 a_n1398_n197# a_n1442_n100# 0.00fF
C2124 w_n4520_n851# a_n3238_n632# 0.03fF
C2125 a_702_n197# a_750_n100# 0.00fF
C2126 w_n4520_n851# a_72_131# 0.12fF
C2127 a_1500_n632# a_30_n632# 0.00fF
C2128 w_n4520_n851# a_n2236_n729# 0.12fF
C2129 a_n2190_n100# a_n2238_n197# 0.00fF
C2130 a_n4078_n632# a_n2490_n632# 0.00fF
C2131 a_n3448_n632# a_n3120_n632# 0.02fF
C2132 a_n3540_n632# a_n3028_n632# 0.01fF
C2133 a_n3658_n632# a_n2910_n632# 0.01fF
C2134 a_n3868_n632# a_n2700_n632# 0.01fF
C2135 a_n3330_n632# a_n3238_n632# 0.09fF
C2136 a_n3960_n632# a_n2608_n632# 0.00fF
C2137 a_2852_n632# a_2804_n729# 0.00fF
C2138 a_1080_n632# a_1802_n632# 0.01fF
C2139 a_1078_n100# a_1288_n100# 0.03fF
C2140 a_n2700_n632# a_n1440_n632# 0.00fF
C2141 w_n4520_n851# a_n2866_n401# 0.10fF
C2142 a_n2490_n632# a_n1650_n632# 0.01fF
C2143 a_n2398_n632# a_n1768_n632# 0.01fF
C2144 a_n2608_n632# a_n1558_n632# 0.01fF
C2145 a_n2028_131# a_n1398_n197# 0.00fF
C2146 a_122_n632# a_n1440_n632# 0.00fF
C2147 a_n3120_n632# a_n3076_n729# 0.00fF
C2148 w_n4520_n851# a_n2658_n197# 0.10fF
C2149 a_n3286_n401# a_n3238_n632# 0.00fF
C2150 a_1380_n100# a_1288_n100# 0.09fF
C2151 a_1498_n100# a_1170_n100# 0.02fF
C2152 a_1590_n100# a_1078_n100# 0.01fF
C2153 a_n2188_n632# a_n1860_n632# 0.02fF
C2154 a_n2070_n632# a_n1978_n632# 0.09fF
C2155 a_1962_n197# a_2802_n197# 0.01fF
C2156 a_n3076_n729# a_n1816_n729# 0.00fF
C2157 a_n2656_n729# a_n2236_n729# 0.01fF
C2158 a_2642_n632# a_2970_n632# 0.02fF
C2159 a_2760_n632# a_2852_n632# 0.09fF
C2160 a_n2868_131# a_n3078_n197# 0.00fF
C2161 a_542_n632# a_n810_n632# 0.00fF
C2162 a_n2446_n401# a_n3076_n729# 0.00fF
C2163 a_n3286_n401# a_n2236_n729# 0.00fF
C2164 a_n2866_n401# a_n2656_n729# 0.00fF
C2165 a_n2026_n401# a_n3496_n729# 0.00fF
C2166 a_542_n632# a_1710_n632# 0.01fF
C2167 a_540_n100# a_1170_n100# 0.01fF
C2168 a_28_n100# a_120_n100# 0.09fF
C2169 a_n90_n100# a_238_n100# 0.02fF
C2170 a_n3286_n401# a_n2866_n401# 0.01fF
C2171 a_n3706_n401# a_n2446_n401# 0.00fF
C2172 a_n510_n100# a_868_n100# 0.00fF
C2173 a_1380_n100# a_1590_n100# 0.03fF
C2174 a_28_n100# a_n720_n100# 0.01fF
C2175 a_3272_n632# a_3902_n632# 0.01fF
C2176 a_3482_n632# a_3692_n632# 0.03fF
C2177 a_3390_n632# a_3810_n632# 0.02fF
C2178 a_1962_n197# a_1964_n729# 0.01fF
C2179 a_2172_131# a_1542_n197# 0.00fF
C2180 a_n2658_n197# a_n2656_n729# 0.01fF
C2181 a_282_n197# a_n1188_131# 0.00fF
C2182 a_282_n197# a_912_131# 0.00fF
C2183 a_3178_n100# a_4110_n100# 0.01fF
C2184 a_1498_n100# a_540_n100# 0.01fF
C2185 a_n88_n632# a_n928_n632# 0.01fF
C2186 a_n2610_n100# a_n2608_n632# 0.00fF
C2187 w_n4520_n851# a_1752_131# 0.12fF
C2188 a_1080_n632# a_2550_n632# 0.00fF
C2189 a_1124_n729# a_1964_n729# 0.01fF
C2190 a_448_n100# a_658_n100# 0.03fF
C2191 a_n1560_n100# w_n4520_n851# 0.02fF
C2192 a_3644_n729# a_3690_n100# 0.00fF
C2193 w_n4520_n851# a_1754_n401# 0.10fF
C2194 w_n4520_n851# a_284_n729# 0.12fF
C2195 a_n298_n632# w_n4520_n851# 0.01fF
C2196 a_n3498_n197# a_n3540_n632# 0.00fF
C2197 a_1290_n632# a_1500_n632# 0.03fF
C2198 a_n1862_n100# a_n1350_n100# 0.01fF
C2199 a_n2072_n100# a_n1140_n100# 0.01fF
C2200 a_n1770_n100# a_n1442_n100# 0.02fF
C2201 a_n2190_n100# a_n1022_n100# 0.01fF
C2202 a_n2282_n100# a_n930_n100# 0.00fF
C2203 a_n2400_n100# a_n812_n100# 0.00fF
C2204 a_n1980_n100# a_n1232_n100# 0.01fF
C2205 a_n3332_n100# a_n3030_n100# 0.02fF
C2206 a_330_n100# a_284_n729# 0.00fF
C2207 a_n3240_n100# a_n3122_n100# 0.07fF
C2208 a_n1770_n100# a_n1816_n729# 0.00fF
C2209 a_n1768_n632# a_n928_n632# 0.01fF
C2210 a_n1650_n632# a_n1020_n632# 0.01fF
C2211 a_n1440_n632# a_n1230_n632# 0.03fF
C2212 a_n1558_n632# a_n1138_n632# 0.02fF
C2213 a_n3498_n197# a_n3496_n729# 0.01fF
C2214 a_n1396_n729# a_n976_n729# 0.01fF
C2215 a_n1816_n729# a_n556_n729# 0.00fF
C2216 a_2382_n197# a_912_131# 0.00fF
C2217 a_n300_n100# w_n4520_n851# 0.02fF
C2218 a_n2026_n401# a_n976_n729# 0.00fF
C2219 a_n3498_n197# a_n3542_n100# 0.00fF
C2220 a_752_n632# a_30_n632# 0.01fF
C2221 a_870_n632# a_n88_n632# 0.01fF
C2222 w_n4520_n851# a_3644_n729# 0.10fF
C2223 a_4020_n632# a_3600_n632# 0.02fF
C2224 a_4112_n632# a_3482_n632# 0.01fF
C2225 a_120_n100# a_74_n401# 0.00fF
C2226 a_2640_n100# a_2850_n100# 0.03fF
C2227 a_2548_n100# a_2968_n100# 0.02fF
C2228 a_2430_n100# a_3060_n100# 0.01fF
C2229 a_2338_n100# a_3178_n100# 0.01fF
C2230 a_660_n632# a_1500_n632# 0.01fF
C2231 a_450_n632# w_n4520_n851# 0.01fF
C2232 a_n300_n100# a_330_n100# 0.01fF
C2233 a_3482_n632# a_3434_n401# 0.00fF
C2234 a_120_n100# a_n930_n100# 0.01fF
C2235 a_n510_n100# a_n1442_n100# 0.01fF
C2236 a_n930_n100# a_n720_n100# 0.03fF
C2237 a_n1022_n100# a_n602_n100# 0.02fF
C2238 a_n4078_n632# a_n3658_n632# 0.02fF
C2239 a_n4170_n632# a_n3540_n632# 0.01fF
C2240 a_2220_n100# a_868_n100# 0.00fF
C2241 w_n4520_n851# a_n1860_n632# 0.01fF
C2242 a_30_n632# a_n1138_n632# 0.01fF
C2243 w_n4520_n851# a_2970_n632# 0.03fF
C2244 w_n4520_n851# a_702_n197# 0.10fF
C2245 a_332_n632# a_n180_n632# 0.01fF
C2246 a_1290_n632# a_2222_n632# 0.01fF
C2247 a_1382_n632# a_2130_n632# 0.01fF
C2248 a_n2868_131# a_n2238_n197# 0.00fF
C2249 a_n4126_n401# a_n4170_n632# 0.00fF
C2250 a_122_n632# a_1382_n632# 0.00fF
C2251 a_332_n632# a_1172_n632# 0.01fF
C2252 a_n3868_n632# a_n3870_n100# 0.00fF
C2253 a_n2910_n632# a_n2280_n632# 0.01fF
C2254 a_n3330_n632# a_n1860_n632# 0.00fF
C2255 a_n3238_n632# a_n1978_n632# 0.00fF
C2256 a_n2818_n632# a_n2398_n632# 0.02fF
C2257 a_3808_n100# a_3900_n100# 0.09fF
C2258 a_3690_n100# a_4018_n100# 0.02fF
C2259 a_3598_n100# a_4110_n100# 0.01fF
C2260 a_n3120_n632# a_n2070_n632# 0.01fF
C2261 a_n3028_n632# a_n2188_n632# 0.01fF
C2262 a_n1652_n100# a_n1560_n100# 0.09fF
C2263 a_2430_n100# a_2432_n632# 0.00fF
C2264 a_1334_n401# a_1754_n401# 0.01fF
C2265 a_494_n401# a_1124_n729# 0.00fF
C2266 a_914_n401# a_704_n729# 0.00fF
C2267 a_n3030_n100# w_n4520_n851# 0.03fF
C2268 a_1334_n401# a_284_n729# 0.00fF
C2269 a_660_n632# a_2222_n632# 0.00fF
C2270 a_542_n632# a_n928_n632# 0.00fF
C2271 a_n2448_131# a_n3078_n197# 0.00fF
C2272 a_n136_n729# a_284_n729# 0.01fF
C2273 a_n2028_131# a_n2070_n632# 0.00fF
C2274 a_n600_n632# a_n88_n632# 0.01fF
C2275 a_1590_n100# a_1544_n729# 0.00fF
C2276 a_n390_n632# a_n298_n632# 0.09fF
C2277 a_n508_n632# a_n180_n632# 0.02fF
C2278 a_n1770_n100# a_n182_n100# 0.00fF
C2279 a_n1560_n100# a_n392_n100# 0.01fF
C2280 a_n1652_n100# a_n300_n100# 0.00fF
C2281 a_962_n632# a_n298_n632# 0.00fF
C2282 a_74_n401# a_494_n401# 0.01fF
C2283 a_1172_n632# a_2012_n632# 0.01fF
C2284 a_2758_n100# a_1288_n100# 0.00fF
C2285 a_120_n100# a_1170_n100# 0.01fF
C2286 a_752_n632# a_1290_n632# 0.01fF
C2287 w_n4520_n851# a_4018_n100# 0.08fF
C2288 a_1498_n100# a_1500_n632# 0.00fF
C2289 a_2012_n632# a_3062_n632# 0.01fF
C2290 a_1920_n632# a_3180_n632# 0.00fF
C2291 a_1802_n632# a_3272_n632# 0.00fF
C2292 a_n2492_n100# a_n3870_n100# 0.00fF
C2293 a_n2702_n100# a_n3660_n100# 0.01fF
C2294 a_n2820_n100# a_n3542_n100# 0.01fF
C2295 a_238_n100# a_n1140_n100# 0.00fF
C2296 a_n2912_n100# a_n3450_n100# 0.01fF
C2297 a_n2610_n100# a_n3752_n100# 0.01fF
C2298 a_2174_n401# a_2804_n729# 0.00fF
C2299 a_1754_n401# a_3224_n729# 0.00fF
C2300 a_2010_n100# a_960_n100# 0.01fF
C2301 a_n4172_n100# a_n3752_n100# 0.02fF
C2302 a_2010_n100# a_2338_n100# 0.02fF
C2303 a_1918_n100# a_2430_n100# 0.01fF
C2304 a_1800_n100# a_2548_n100# 0.01fF
C2305 a_1708_n100# a_2640_n100# 0.01fF
C2306 a_1590_n100# a_2758_n100# 0.01fF
C2307 a_1498_n100# a_2850_n100# 0.00fF
C2308 a_1380_n100# a_2968_n100# 0.00fF
C2309 a_n4080_n100# a_n3870_n100# 0.03fF
C2310 a_1498_n100# a_120_n100# 0.00fF
C2311 a_2640_n100# a_3270_n100# 0.01fF
C2312 a_2548_n100# a_3388_n100# 0.01fF
C2313 a_2430_n100# a_3480_n100# 0.01fF
C2314 a_2338_n100# a_3598_n100# 0.00fF
C2315 a_450_n632# a_n390_n632# 0.01fF
C2316 a_n810_n632# a_n1558_n632# 0.01fF
C2317 a_n600_n632# a_n1768_n632# 0.01fF
C2318 a_n718_n632# a_n1650_n632# 0.01fF
C2319 a_n558_n197# a_n138_n197# 0.01fF
C2320 a_28_n100# a_658_n100# 0.01fF
C2321 a_n90_n100# a_750_n100# 0.01fF
C2322 a_238_n100# a_448_n100# 0.03fF
C2323 a_120_n100# a_540_n100# 0.02fF
C2324 a_450_n632# a_962_n632# 0.01fF
C2325 a_542_n632# a_870_n632# 0.02fF
C2326 a_660_n632# a_752_n632# 0.09fF
C2327 a_3432_131# a_3642_n197# 0.00fF
C2328 a_332_n632# a_1080_n632# 0.01fF
C2329 a_n392_n100# a_n300_n100# 0.09fF
C2330 a_n510_n100# a_n182_n100# 0.02fF
C2331 a_540_n100# a_n720_n100# 0.00fF
C2332 a_2594_n401# a_2642_n632# 0.00fF
C2333 a_n390_n632# a_n1860_n632# 0.00fF
C2334 a_1918_n100# a_448_n100# 0.00fF
C2335 a_n1020_n632# a_n1022_n100# 0.00fF
C2336 a_1172_n632# a_2760_n632# 0.00fF
C2337 a_3224_n729# a_3644_n729# 0.01fF
C2338 a_2804_n729# a_4064_n729# 0.00fF
C2339 a_2130_n632# a_3692_n632# 0.00fF
C2340 a_2760_n632# a_3062_n632# 0.02fF
C2341 a_2432_n632# a_3390_n632# 0.01fF
C2342 a_2222_n632# a_3600_n632# 0.00fF
C2343 a_2642_n632# a_3180_n632# 0.01fF
C2344 a_2340_n632# a_3482_n632# 0.01fF
C2345 a_2550_n632# a_3272_n632# 0.01fF
C2346 a_72_131# a_n138_n197# 0.00fF
C2347 a_n1652_n100# a_n3030_n100# 0.00fF
C2348 a_n1770_n100# a_n2912_n100# 0.01fF
C2349 a_n1862_n100# a_n2820_n100# 0.01fF
C2350 a_n2190_n100# a_n2492_n100# 0.02fF
C2351 a_n2072_n100# a_n2610_n100# 0.01fF
C2352 a_n1560_n100# a_n3122_n100# 0.00fF
C2353 a_n1980_n100# a_n2702_n100# 0.01fF
C2354 w_n4520_n851# a_n3028_n632# 0.03fF
C2355 a_n2400_n100# a_n3870_n100# 0.00fF
C2356 a_n1188_131# a_n1230_n632# 0.00fF
C2357 a_n810_n632# a_30_n632# 0.01fF
C2358 w_n4520_n851# a_n1350_n100# 0.02fF
C2359 a_n3918_n197# a_n3498_n197# 0.01fF
C2360 w_n4520_n851# a_n1396_n729# 0.12fF
C2361 a_n3960_n632# a_n2398_n632# 0.00fF
C2362 a_n3868_n632# a_n2490_n632# 0.00fF
C2363 a_n3238_n632# a_n3120_n632# 0.07fF
C2364 a_1080_n632# a_n508_n632# 0.00fF
C2365 a_n3330_n632# a_n3028_n632# 0.02fF
C2366 a_n3448_n632# a_n2910_n632# 0.01fF
C2367 a_n3540_n632# a_n2818_n632# 0.01fF
C2368 a_n3750_n632# a_n2608_n632# 0.01fF
C2369 a_1080_n632# a_2012_n632# 0.01fF
C2370 a_n2280_n632# a_n1650_n632# 0.01fF
C2371 a_n2398_n632# a_n1558_n632# 0.01fF
C2372 a_n2608_n632# a_n1348_n632# 0.00fF
C2373 a_n2700_n632# a_n1230_n632# 0.00fF
C2374 a_n2490_n632# a_n1440_n632# 0.01fF
C2375 a_n2188_n632# a_n1768_n632# 0.02fF
C2376 w_n4520_n851# a_n2026_n401# 0.10fF
C2377 a_n2028_131# a_n558_n197# 0.00fF
C2378 a_750_n100# a_704_n729# 0.00fF
C2379 a_122_n632# a_n1230_n632# 0.00fF
C2380 a_n348_131# a_n768_131# 0.01fF
C2381 a_n2448_131# a_n2238_n197# 0.00fF
C2382 a_2220_n100# a_2174_n401# 0.00fF
C2383 a_1590_n100# a_1288_n100# 0.02fF
C2384 a_1708_n100# a_1170_n100# 0.01fF
C2385 a_1800_n100# a_1078_n100# 0.01fF
C2386 a_n1978_n632# a_n1860_n632# 0.07fF
C2387 a_2382_n197# a_3222_n197# 0.01fF
C2388 a_n2656_n729# a_n1396_n729# 0.00fF
C2389 a_n2236_n729# a_n1816_n729# 0.01fF
C2390 a_2852_n632# a_2970_n632# 0.07fF
C2391 a_n2446_n401# a_n2236_n729# 0.00fF
C2392 a_n2026_n401# a_n2656_n729# 0.00fF
C2393 a_n1606_n401# a_n3076_n729# 0.00fF
C2394 a_n2866_n401# a_n1816_n729# 0.00fF
C2395 a_542_n632# a_n600_n632# 0.01fF
C2396 a_494_n401# a_540_n100# 0.00fF
C2397 a_542_n632# a_1920_n632# 0.00fF
C2398 a_n3286_n401# a_n2026_n401# 0.00fF
C2399 a_n2866_n401# a_n2446_n401# 0.01fF
C2400 a_n300_n100# a_868_n100# 0.01fF
C2401 a_3852_131# a_2802_n197# 0.00fF
C2402 a_3482_n632# a_3902_n632# 0.02fF
C2403 a_3600_n632# a_3810_n632# 0.03fF
C2404 a_1498_n100# a_1708_n100# 0.03fF
C2405 a_1380_n100# a_1800_n100# 0.02fF
C2406 a_658_n100# a_n930_n100# 0.00fF
C2407 a_2172_131# a_2382_n197# 0.00fF
C2408 a_2382_n197# a_2384_n729# 0.01fF
C2409 a_n2400_n100# a_n2190_n100# 0.03fF
C2410 a_660_n632# a_658_n100# 0.00fF
C2411 a_1708_n100# a_540_n100# 0.01fF
C2412 a_n2492_n100# a_n2490_n632# 0.00fF
C2413 a_1544_n729# a_2384_n729# 0.01fF
C2414 a_n2028_131# a_n2658_n197# 0.00fF
C2415 a_n768_131# a_n1398_n197# 0.00fF
C2416 a_3012_131# w_n4520_n851# 0.13fF
C2417 w_n4520_n851# a_2594_n401# 0.10fF
C2418 w_n4520_n851# a_n3498_n197# 0.11fF
C2419 a_2850_n100# a_2802_n197# 0.00fF
C2420 a_n2238_n197# a_n2280_n632# 0.00fF
C2421 a_1592_n632# a_1544_n729# 0.00fF
C2422 a_n2868_131# a_n4128_131# 0.00fF
C2423 a_n88_n632# w_n4520_n851# 0.01fF
C2424 a_2592_131# a_4062_n197# 0.00fF
C2425 a_1290_n632# a_1710_n632# 0.02fF
C2426 a_1382_n632# a_1592_n632# 0.03fF
C2427 a_n1770_n100# a_n1232_n100# 0.01fF
C2428 a_n1980_n100# a_n1022_n100# 0.01fF
C2429 a_n1862_n100# a_n1140_n100# 0.01fF
C2430 a_n1652_n100# a_n1350_n100# 0.02fF
C2431 a_n2072_n100# a_n930_n100# 0.01fF
C2432 a_n2190_n100# a_n812_n100# 0.00fF
C2433 a_n2282_n100# a_n720_n100# 0.00fF
C2434 a_n1560_n100# a_n1442_n100# 0.07fF
C2435 a_n3240_n100# a_n2912_n100# 0.02fF
C2436 a_n3332_n100# a_n2820_n100# 0.01fF
C2437 a_n3122_n100# a_n3030_n100# 0.09fF
C2438 a_n1348_n632# a_n1138_n632# 0.03fF
C2439 a_n1440_n632# a_n1020_n632# 0.02fF
C2440 a_n1558_n632# a_n928_n632# 0.01fF
C2441 w_n4520_n851# a_3180_n632# 0.03fF
C2442 a_n3078_n197# a_n3076_n729# 0.01fF
C2443 a_n1396_n729# a_n136_n729# 0.00fF
C2444 a_3432_131# a_3480_n100# 0.00fF
C2445 a_n90_n100# w_n4520_n851# 0.02fF
C2446 a_n1186_n401# a_n976_n729# 0.00fF
C2447 a_n1606_n401# a_n556_n729# 0.00fF
C2448 a_2382_n197# a_2340_n632# 0.00fF
C2449 a_n718_n632# a_n766_n401# 0.00fF
C2450 a_660_n632# a_n810_n632# 0.00fF
C2451 a_4112_n632# a_3692_n632# 0.02fF
C2452 a_4020_n632# a_3810_n632# 0.03fF
C2453 w_n4520_n851# a_n4170_n632# 0.14fF
C2454 a_660_n632# a_1710_n632# 0.01fF
C2455 a_2758_n100# a_2968_n100# 0.03fF
C2456 a_2640_n100# a_3060_n100# 0.02fF
C2457 a_2548_n100# a_3178_n100# 0.01fF
C2458 a_658_n100# a_1170_n100# 0.01fF
C2459 w_n4520_n851# a_n1768_n632# 0.01fF
C2460 a_28_n100# a_238_n100# 0.03fF
C2461 a_n90_n100# a_330_n100# 0.02fF
C2462 a_2172_131# a_912_131# 0.00fF
C2463 a_n510_n100# a_960_n100# 0.00fF
C2464 a_120_n100# a_n720_n100# 0.01fF
C2465 a_2592_131# a_1542_n197# 0.00fF
C2466 a_n300_n100# a_n1442_n100# 0.01fF
C2467 a_n510_n100# a_n1232_n100# 0.01fF
C2468 a_n392_n100# a_n1350_n100# 0.01fF
C2469 a_n3868_n632# a_n3658_n632# 0.03fF
C2470 a_n4078_n632# a_n3448_n632# 0.01fF
C2471 a_n4170_n632# a_n3330_n632# 0.01fF
C2472 a_702_n197# a_n138_n197# 0.01fF
C2473 a_n3960_n632# a_n3540_n632# 0.02fF
C2474 a_n812_n100# a_n602_n100# 0.03fF
C2475 a_2172_131# a_2130_n632# 0.00fF
C2476 a_n3330_n632# a_n1768_n632# 0.00fF
C2477 a_1498_n100# a_658_n100# 0.01fF
C2478 a_30_n632# a_n928_n632# 0.01fF
C2479 a_n3868_n632# a_n3916_n729# 0.00fF
C2480 a_1592_n632# a_2130_n632# 0.01fF
C2481 a_1500_n632# a_2222_n632# 0.01fF
C2482 a_1382_n632# a_2340_n632# 0.01fF
C2483 a_1290_n632# a_2432_n632# 0.01fF
C2484 a_240_n632# a_282_n197# 0.00fF
C2485 a_122_n632# a_1592_n632# 0.00fF
C2486 a_540_n100# a_658_n100# 0.07fF
C2487 a_448_n100# a_750_n100# 0.02fF
C2488 a_n3750_n632# a_n3752_n100# 0.00fF
C2489 a_n3028_n632# a_n1978_n632# 0.01fF
C2490 a_n2818_n632# a_n2188_n632# 0.01fF
C2491 a_n2910_n632# a_n2070_n632# 0.01fF
C2492 a_n3120_n632# a_n1860_n632# 0.00fF
C2493 a_3900_n100# a_4018_n100# 0.07fF
C2494 a_3808_n100# a_4110_n100# 0.02fF
C2495 a_n348_131# a_492_131# 0.01fF
C2496 a_2548_n100# a_2550_n632# 0.00fF
C2497 w_n4520_n851# a_704_n729# 0.12fF
C2498 a_n1860_n632# a_n1816_n729# 0.00fF
C2499 a_n3288_131# a_n3332_n100# 0.00fF
C2500 a_1754_n401# a_2174_n401# 0.01fF
C2501 a_1334_n401# a_2594_n401# 0.00fF
C2502 a_n2026_n401# a_n1978_n632# 0.00fF
C2503 a_n2820_n100# w_n4520_n851# 0.02fF
C2504 a_3642_n197# a_3600_n632# 0.00fF
C2505 a_1918_n100# a_1962_n197# 0.00fF
C2506 a_494_n401# a_1964_n729# 0.00fF
C2507 a_2548_n100# a_2592_131# 0.00fF
C2508 a_n3288_131# a_n3918_n197# 0.00fF
C2509 a_n2238_n197# a_n1398_n197# 0.01fF
C2510 a_n88_n632# a_n136_n729# 0.00fF
C2511 a_3852_131# a_3810_n632# 0.00fF
C2512 a_n298_n632# a_n180_n632# 0.07fF
C2513 a_n390_n632# a_n88_n632# 0.02fF
C2514 a_n2868_131# a_n3708_131# 0.01fF
C2515 a_n1652_n100# a_n90_n100# 0.00fF
C2516 a_962_n632# a_n88_n632# 0.01fF
C2517 a_1172_n632# a_n298_n632# 0.00fF
C2518 a_n1560_n100# a_n182_n100# 0.00fF
C2519 a_870_n632# a_30_n632# 0.01fF
C2520 a_n3030_n100# a_n1442_n100# 0.00fF
C2521 a_n2700_n632# a_n2490_n632# 0.03fF
C2522 a_2130_n632# a_2340_n632# 0.03fF
C2523 a_752_n632# a_1500_n632# 0.01fF
C2524 a_542_n632# w_n4520_n851# 0.01fF
C2525 a_2012_n632# a_3272_n632# 0.00fF
C2526 a_1920_n632# a_3390_n632# 0.00fF
C2527 a_1590_n100# a_1592_n632# 0.00fF
C2528 a_n348_131# a_n346_n401# 0.01fF
C2529 a_n90_n100# a_n136_n729# 0.00fF
C2530 a_n2492_n100# a_n3660_n100# 0.01fF
C2531 a_n2702_n100# a_n3450_n100# 0.01fF
C2532 a_n2610_n100# a_n3542_n100# 0.01fF
C2533 a_238_n100# a_n930_n100# 0.01fF
C2534 a_2174_n401# a_3644_n729# 0.00fF
C2535 a_2594_n401# a_3224_n729# 0.00fF
C2536 a_3014_n401# a_2804_n729# 0.00fF
C2537 a_2220_n100# a_960_n100# 0.00fF
C2538 a_n3962_n100# a_n3752_n100# 0.03fF
C2539 a_n4080_n100# a_n3660_n100# 0.02fF
C2540 a_n4172_n100# a_n3542_n100# 0.01fF
C2541 a_1800_n100# a_2758_n100# 0.01fF
C2542 a_1708_n100# a_2850_n100# 0.01fF
C2543 a_1590_n100# a_2968_n100# 0.00fF
C2544 a_1498_n100# a_3060_n100# 0.00fF
C2545 a_492_131# a_1332_131# 0.01fF
C2546 a_1708_n100# a_120_n100# 0.00fF
C2547 a_2220_n100# a_2338_n100# 0.07fF
C2548 a_2128_n100# a_2430_n100# 0.02fF
C2549 a_2010_n100# a_2548_n100# 0.01fF
C2550 a_1918_n100# a_2640_n100# 0.01fF
C2551 a_2640_n100# a_3480_n100# 0.01fF
C2552 a_2548_n100# a_3598_n100# 0.01fF
C2553 a_2430_n100# a_3690_n100# 0.00fF
C2554 a_2338_n100# a_3808_n100# 0.00fF
C2555 a_2758_n100# a_3388_n100# 0.01fF
C2556 a_2850_n100# a_3270_n100# 0.02fF
C2557 w_n4520_n851# a_1122_n197# 0.10fF
C2558 a_1542_n197# a_1332_131# 0.00fF
C2559 a_450_n632# a_n180_n632# 0.01fF
C2560 a_n718_n632# a_n1440_n632# 0.01fF
C2561 a_n600_n632# a_n1558_n632# 0.01fF
C2562 a_n508_n632# a_n1650_n632# 0.01fF
C2563 a_n810_n632# a_n1348_n632# 0.01fF
C2564 a_n390_n632# a_n1768_n632# 0.00fF
C2565 a_450_n632# a_1172_n632# 0.01fF
C2566 a_240_n632# a_1382_n632# 0.01fF
C2567 a_n300_n100# a_n182_n100# 0.07fF
C2568 a_n392_n100# a_n90_n100# 0.02fF
C2569 a_3180_n632# a_3224_n729# 0.00fF
C2570 a_n3288_131# w_n4520_n851# 0.13fF
C2571 a_n928_n632# a_n930_n100# 0.00fF
C2572 a_1334_n401# a_704_n729# 0.00fF
C2573 a_914_n401# a_1124_n729# 0.00fF
C2574 a_3644_n729# a_4064_n729# 0.01fF
C2575 a_752_n632# a_2222_n632# 0.00fF
C2576 a_2852_n632# a_3180_n632# 0.02fF
C2577 a_2970_n632# a_3062_n632# 0.09fF
C2578 a_2550_n632# a_3482_n632# 0.01fF
C2579 a_2340_n632# a_3692_n632# 0.00fF
C2580 a_2642_n632# a_3390_n632# 0.01fF
C2581 a_2222_n632# a_3810_n632# 0.00fF
C2582 a_660_n632# a_n928_n632# 0.00fF
C2583 a_2432_n632# a_3600_n632# 0.01fF
C2584 a_2760_n632# a_3272_n632# 0.01fF
C2585 a_n136_n729# a_704_n729# 0.01fF
C2586 a_n3288_131# a_n3330_n632# 0.00fF
C2587 a_n1770_n100# a_n2702_n100# 0.01fF
C2588 a_3852_131# a_3854_n401# 0.01fF
C2589 a_n1862_n100# a_n2610_n100# 0.01fF
C2590 a_n1652_n100# a_n2820_n100# 0.01fF
C2591 a_n1560_n100# a_n2912_n100# 0.00fF
C2592 a_n1980_n100# a_n2492_n100# 0.01fF
C2593 w_n4520_n851# a_n2818_n632# 0.02fF
C2594 a_3434_n401# a_2384_n729# 0.00fF
C2595 a_2430_n100# w_n4520_n851# 0.02fF
C2596 a_n3708_131# a_n3660_n100# 0.00fF
C2597 a_n2282_n100# a_n3752_n100# 0.00fF
C2598 a_n600_n632# a_30_n632# 0.01fF
C2599 a_n2400_n100# a_n3660_n100# 0.00fF
C2600 a_n2448_131# a_n2492_n100# 0.00fF
C2601 w_n4520_n851# a_n1140_n100# 0.02fF
C2602 a_n3288_131# a_n3286_n401# 0.01fF
C2603 a_n1862_n100# a_n1818_n197# 0.00fF
C2604 a_n3238_n632# a_n2910_n632# 0.02fF
C2605 a_n3330_n632# a_n2818_n632# 0.01fF
C2606 a_n3120_n632# a_n3028_n632# 0.09fF
C2607 a_n3750_n632# a_n2398_n632# 0.00fF
C2608 a_n3868_n632# a_n2280_n632# 0.00fF
C2609 a_1080_n632# a_n298_n632# 0.00fF
C2610 a_74_n401# a_914_n401# 0.01fF
C2611 a_n2608_n632# a_n1138_n632# 0.00fF
C2612 a_n2398_n632# a_n1348_n632# 0.01fF
C2613 a_n1978_n632# a_n1768_n632# 0.03fF
C2614 a_n2280_n632# a_n1440_n632# 0.01fF
C2615 a_n2490_n632# a_n1230_n632# 0.00fF
C2616 w_n4520_n851# a_n1186_n401# 0.10fF
C2617 a_n2070_n632# a_n1650_n632# 0.02fF
C2618 a_n2188_n632# a_n1558_n632# 0.01fF
C2619 a_n1608_131# a_n1818_n197# 0.00fF
C2620 a_870_n632# a_1290_n632# 0.02fF
C2621 a_238_n100# a_1170_n100# 0.01fF
C2622 a_122_n632# a_n1020_n632# 0.01fF
C2623 a_122_n632# a_240_n632# 0.07fF
C2624 a_330_n100# a_n1140_n100# 0.00fF
C2625 a_n2866_n401# a_n2910_n632# 0.00fF
C2626 w_n4520_n851# a_448_n100# 0.02fF
C2627 a_n1442_n100# a_n1350_n100# 0.09fF
C2628 a_1800_n100# a_1288_n100# 0.01fF
C2629 a_1918_n100# a_1170_n100# 0.01fF
C2630 a_2010_n100# a_1078_n100# 0.01fF
C2631 a_2802_n197# a_3642_n197# 0.01fF
C2632 a_1498_n100# a_238_n100# 0.00fF
C2633 a_n1816_n729# a_n1396_n729# 0.01fF
C2634 a_n2026_n401# a_n1816_n729# 0.00fF
C2635 a_n1186_n401# a_n2656_n729# 0.00fF
C2636 a_542_n632# a_n390_n632# 0.01fF
C2637 a_n1606_n401# a_n2236_n729# 0.00fF
C2638 a_n2446_n401# a_n1396_n729# 0.00fF
C2639 a_542_n632# a_962_n632# 0.02fF
C2640 a_330_n100# a_448_n100# 0.07fF
C2641 a_238_n100# a_540_n100# 0.02fF
C2642 a_n2866_n401# a_n1606_n401# 0.00fF
C2643 a_660_n632# a_870_n632# 0.03fF
C2644 a_120_n100# a_658_n100# 0.01fF
C2645 a_28_n100# a_750_n100# 0.01fF
C2646 a_n90_n100# a_868_n100# 0.01fF
C2647 a_450_n632# a_1080_n632# 0.01fF
C2648 a_3852_131# a_3642_n197# 0.00fF
C2649 a_n2446_n401# a_n2026_n401# 0.01fF
C2650 a_1590_n100# a_1800_n100# 0.03fF
C2651 a_1498_n100# a_1918_n100# 0.02fF
C2652 a_1380_n100# a_2010_n100# 0.01fF
C2653 a_3692_n632# a_3902_n632# 0.03fF
C2654 a_658_n100# a_n720_n100# 0.00fF
C2655 a_1708_n100# a_3270_n100# 0.00fF
C2656 a_2172_131# a_3222_n197# 0.00fF
C2657 a_n3918_n197# a_n3960_n632# 0.00fF
C2658 a_n3658_n632# a_n2700_n632# 0.01fF
C2659 a_n2028_131# a_n2026_n401# 0.01fF
C2660 a_n2400_n100# a_n1980_n100# 0.02fF
C2661 a_n2282_n100# a_n2072_n100# 0.03fF
C2662 a_1918_n100# a_540_n100# 0.00fF
C2663 a_4020_n632# a_2432_n632# 0.00fF
C2664 a_1920_n632# a_1962_n197# 0.00fF
C2665 a_n2448_131# a_n3708_131# 0.00fF
C2666 a_n2448_131# a_n2400_n100# 0.00fF
C2667 a_n768_131# a_n558_n197# 0.00fF
C2668 a_1500_n632# a_1710_n632# 0.03fF
C2669 a_1382_n632# a_1802_n632# 0.02fF
C2670 a_1290_n632# a_1920_n632# 0.01fF
C2671 a_n2072_n100# a_n720_n100# 0.00fF
C2672 a_n2190_n100# a_n602_n100# 0.00fF
C2673 a_n1770_n100# a_n1022_n100# 0.01fF
C2674 a_n1980_n100# a_n812_n100# 0.01fF
C2675 a_n1560_n100# a_n1232_n100# 0.02fF
C2676 a_n1862_n100# a_n930_n100# 0.01fF
C2677 a_n1652_n100# a_n1140_n100# 0.01fF
C2678 a_n3332_n100# a_n2610_n100# 0.01fF
C2679 a_n3240_n100# a_n2702_n100# 0.01fF
C2680 a_n3030_n100# a_n2912_n100# 0.07fF
C2681 a_n3122_n100# a_n2820_n100# 0.02fF
C2682 a_n1230_n632# a_n1020_n632# 0.03fF
C2683 a_n346_n401# a_n556_n729# 0.00fF
C2684 a_n1348_n632# a_n928_n632# 0.02fF
C2685 a_74_n401# a_n976_n729# 0.00fF
C2686 a_n90_n100# a_n138_n197# 0.00fF
C2687 w_n4520_n851# a_3390_n632# 0.03fF
C2688 a_1380_n100# a_1332_131# 0.00fF
C2689 a_72_131# a_n768_131# 0.01fF
C2690 a_240_n632# a_n1230_n632# 0.00fF
C2691 a_n1560_n100# a_n1606_n401# 0.00fF
C2692 a_n930_n100# a_n976_n729# 0.00fF
C2693 a_n3332_n100# a_n4172_n100# 0.01fF
C2694 a_n348_131# a_282_n197# 0.00fF
C2695 a_n1186_n401# a_n136_n729# 0.00fF
C2696 a_n766_n401# a_n556_n729# 0.00fF
C2697 a_n1398_n197# a_n1440_n632# 0.00fF
C2698 a_4112_n632# a_3902_n632# 0.03fF
C2699 a_n2028_131# a_n3498_n197# 0.00fF
C2700 w_n4520_n851# a_n3960_n632# 0.06fF
C2701 a_660_n632# a_n600_n632# 0.00fF
C2702 a_n2658_n197# a_n3078_n197# 0.01fF
C2703 a_660_n632# a_1920_n632# 0.00fF
C2704 a_2758_n100# a_3178_n100# 0.02fF
C2705 a_2850_n100# a_3060_n100# 0.03fF
C2706 a_3810_n632# a_3854_n401# 0.00fF
C2707 w_n4520_n851# a_n1558_n632# 0.01fF
C2708 a_n300_n100# a_960_n100# 0.00fF
C2709 a_n2448_131# a_n1188_131# 0.00fF
C2710 a_2592_131# a_2382_n197# 0.00fF
C2711 a_n510_n100# a_n1022_n100# 0.01fF
C2712 a_n392_n100# a_n1140_n100# 0.01fF
C2713 a_n300_n100# a_n1232_n100# 0.01fF
C2714 a_n182_n100# a_n1350_n100# 0.01fF
C2715 a_n90_n100# a_n1442_n100# 0.00fF
C2716 a_n4170_n632# a_n3120_n632# 0.01fF
C2717 a_n3750_n632# a_n3540_n632# 0.03fF
C2718 a_n3960_n632# a_n3330_n632# 0.01fF
C2719 a_n3868_n632# a_n3448_n632# 0.02fF
C2720 a_n4078_n632# a_n3238_n632# 0.01fF
C2721 a_2340_n632# a_2384_n729# 0.00fF
C2722 a_n3238_n632# a_n1650_n632# 0.00fF
C2723 a_n3120_n632# a_n1768_n632# 0.00fF
C2724 a_1708_n100# a_658_n100# 0.01fF
C2725 a_1710_n632# a_2222_n632# 0.01fF
C2726 a_1592_n632# a_2340_n632# 0.01fF
C2727 a_1382_n632# a_2550_n632# 0.01fF
C2728 a_1500_n632# a_2432_n632# 0.01fF
C2729 a_1802_n632# a_2130_n632# 0.02fF
C2730 a_1290_n632# a_2642_n632# 0.00fF
C2731 a_122_n632# a_n718_n632# 0.01fF
C2732 a_n1768_n632# a_n1816_n729# 0.00fF
C2733 a_n392_n100# a_448_n100# 0.01fF
C2734 a_4018_n100# a_4110_n100# 0.09fF
C2735 a_n2910_n632# a_n1860_n632# 0.01fF
C2736 a_n2818_n632# a_n1978_n632# 0.01fF
C2737 a_3432_131# w_n4520_n851# 0.12fF
C2738 a_2640_n100# a_2642_n632# 0.00fF
C2739 a_30_n632# w_n4520_n851# 0.01fF
C2740 a_1754_n401# a_3014_n401# 0.00fF
C2741 a_2174_n401# a_2594_n401# 0.01fF
C2742 a_282_n197# a_1332_131# 0.00fF
C2743 a_n2610_n100# w_n4520_n851# 0.02fF
C2744 a_n1818_n197# a_n978_n197# 0.01fF
C2745 w_n4520_n851# a_n4172_n100# 0.14fF
C2746 w_n4520_n851# a_n1818_n197# 0.10fF
C2747 a_28_n100# w_n4520_n851# 0.02fF
C2748 a_n180_n632# a_n88_n632# 0.09fF
C2749 a_n2820_n100# a_n1442_n100# 0.00fF
C2750 a_1172_n632# a_n88_n632# 0.00fF
C2751 a_n2912_n100# a_n1350_n100# 0.00fF
C2752 a_n2700_n632# a_n2280_n632# 0.02fF
C2753 a_n2608_n632# a_n2398_n632# 0.03fF
C2754 a_n2610_n100# a_n2656_n729# 0.00fF
C2755 a_2130_n632# a_2550_n632# 0.02fF
C2756 a_2222_n632# a_2432_n632# 0.03fF
C2757 a_752_n632# a_n810_n632# 0.00fF
C2758 a_752_n632# a_1710_n632# 0.01fF
C2759 a_750_n100# a_1170_n100# 0.02fF
C2760 a_120_n100# a_238_n100# 0.07fF
C2761 a_28_n100# a_330_n100# 0.02fF
C2762 a_2012_n632# a_3482_n632# 0.00fF
C2763 a_1708_n100# a_1710_n632# 0.00fF
C2764 a_2430_n100# a_868_n100# 0.00fF
C2765 a_n510_n100# a_1078_n100# 0.00fF
C2766 a_492_131# a_n558_n197# 0.00fF
C2767 a_n2492_n100# a_n3450_n100# 0.01fF
C2768 a_n3916_n729# a_n3870_n100# 0.00fF
C2769 a_238_n100# a_n720_n100# 0.01fF
C2770 a_3014_n401# a_3644_n729# 0.00fF
C2771 a_2594_n401# a_4064_n729# 0.00fF
C2772 a_1122_n197# a_n138_n197# 0.00fF
C2773 a_n2238_n197# a_n2236_n729# 0.01fF
C2774 a_3062_n632# a_3180_n632# 0.07fF
C2775 a_n2702_n100# a_n2658_n197# 0.00fF
C2776 a_n3962_n100# a_n3542_n100# 0.02fF
C2777 a_n4080_n100# a_n3450_n100# 0.01fF
C2778 a_n3870_n100# a_n3660_n100# 0.03fF
C2779 a_2220_n100# a_2548_n100# 0.02fF
C2780 a_2128_n100# a_2640_n100# 0.01fF
C2781 a_2010_n100# a_2758_n100# 0.01fF
C2782 a_1918_n100# a_2850_n100# 0.01fF
C2783 a_1800_n100# a_2968_n100# 0.01fF
C2784 a_1708_n100# a_3060_n100# 0.00fF
C2785 a_1590_n100# a_3178_n100# 0.00fF
C2786 a_2430_n100# a_3900_n100# 0.00fF
C2787 a_2548_n100# a_3808_n100# 0.00fF
C2788 a_2640_n100# a_3690_n100# 0.01fF
C2789 a_2758_n100# a_3598_n100# 0.01fF
C2790 a_3060_n100# a_3270_n100# 0.03fF
C2791 a_2968_n100# a_3388_n100# 0.02fF
C2792 a_2850_n100# a_3480_n100# 0.01fF
C2793 a_1498_n100# a_750_n100# 0.01fF
C2794 a_2382_n197# a_1332_131# 0.00fF
C2795 w_n4520_n851# a_1962_n197# 0.10fF
C2796 a_n298_n632# a_n1650_n632# 0.00fF
C2797 a_n508_n632# a_n1440_n632# 0.01fF
C2798 a_n180_n632# a_n1768_n632# 0.00fF
C2799 a_n810_n632# a_n1138_n632# 0.02fF
C2800 a_n390_n632# a_n1558_n632# 0.01fF
C2801 a_n600_n632# a_n1348_n632# 0.01fF
C2802 a_n718_n632# a_n1230_n632# 0.01fF
C2803 a_240_n632# a_1592_n632# 0.00fF
C2804 a_540_n100# a_750_n100# 0.03fF
C2805 a_448_n100# a_868_n100# 0.02fF
C2806 a_n2658_n197# a_n2238_n197# 0.01fF
C2807 a_n182_n100# a_n90_n100# 0.09fF
C2808 a_n348_131# a_n1188_131# 0.01fF
C2809 a_3014_n401# a_2970_n632# 0.00fF
C2810 a_n348_131# a_912_131# 0.00fF
C2811 a_72_131# a_492_131# 0.01fF
C2812 w_n4520_n851# a_1124_n729# 0.12fF
C2813 a_702_n197# a_n768_131# 0.00fF
C2814 a_72_131# a_1542_n197# 0.00fF
C2815 a_2174_n401# a_704_n729# 0.00fF
C2816 a_914_n401# a_1964_n729# 0.00fF
C2817 a_1290_n632# w_n4520_n851# 0.01fF
C2818 a_2550_n632# a_3692_n632# 0.01fF
C2819 a_2432_n632# a_3810_n632# 0.00fF
C2820 a_2852_n632# a_3390_n632# 0.01fF
C2821 a_2970_n632# a_3272_n632# 0.02fF
C2822 a_2760_n632# a_3482_n632# 0.01fF
C2823 a_2642_n632# a_3600_n632# 0.01fF
C2824 a_2340_n632# a_3902_n632# 0.00fF
C2825 a_n1652_n100# a_n2610_n100# 0.01fF
C2826 a_n1770_n100# a_n2492_n100# 0.01fF
C2827 a_n1560_n100# a_n2702_n100# 0.01fF
C2828 a_n978_n197# a_n930_n100# 0.00fF
C2829 a_n3708_131# a_n3706_n401# 0.01fF
C2830 a_n3030_n100# a_n3078_n197# 0.00fF
C2831 w_n4520_n851# a_74_n401# 0.10fF
C2832 a_2640_n100# w_n4520_n851# 0.02fF
C2833 a_n2400_n100# a_n3450_n100# 0.01fF
C2834 a_n390_n632# a_30_n632# 0.02fF
C2835 a_n2282_n100# a_n3542_n100# 0.00fF
C2836 a_n2190_n100# a_n3660_n100# 0.00fF
C2837 w_n4520_n851# a_n930_n100# 0.02fF
C2838 a_n3028_n632# a_n2910_n632# 0.07fF
C2839 a_1080_n632# a_n88_n632# 0.01fF
C2840 a_n3750_n632# a_n2188_n632# 0.00fF
C2841 a_962_n632# a_30_n632# 0.01fF
C2842 a_n3120_n632# a_n2818_n632# 0.02fF
C2843 a_n2490_n632# a_n1020_n632# 0.00fF
C2844 a_n2188_n632# a_n1348_n632# 0.01fF
C2845 a_n1860_n632# a_n1650_n632# 0.03fF
C2846 a_n2398_n632# a_n1138_n632# 0.00fF
C2847 a_n2070_n632# a_n1440_n632# 0.01fF
C2848 a_n1978_n632# a_n1558_n632# 0.02fF
C2849 a_n2280_n632# a_n1230_n632# 0.01fF
C2850 a_870_n632# a_1500_n632# 0.01fF
C2851 a_660_n632# w_n4520_n851# 0.01fF
C2852 a_n1188_131# a_n1398_n197# 0.00fF
C2853 a_n3288_131# a_n2028_131# 0.00fF
C2854 a_330_n100# a_n930_n100# 0.00fF
C2855 a_2010_n100# a_1288_n100# 0.01fF
C2856 a_2128_n100# a_1170_n100# 0.01fF
C2857 a_2220_n100# a_1078_n100# 0.01fF
C2858 a_n1442_n100# a_n1140_n100# 0.02fF
C2859 a_n1350_n100# a_n1232_n100# 0.07fF
C2860 a_912_131# a_1332_131# 0.01fF
C2861 a_1708_n100# a_238_n100# 0.00fF
C2862 a_492_131# a_1752_131# 0.00fF
C2863 a_1542_n197# a_1752_131# 0.00fF
C2864 a_n766_n401# a_n2236_n729# 0.00fF
C2865 a_n1606_n401# a_n1396_n729# 0.00fF
C2866 a_n1186_n401# a_n1816_n729# 0.00fF
C2867 a_542_n632# a_n180_n632# 0.01fF
C2868 a_n2446_n401# a_n1186_n401# 0.00fF
C2869 a_n2026_n401# a_n1606_n401# 0.01fF
C2870 a_542_n632# a_1172_n632# 0.01fF
C2871 a_332_n632# a_1382_n632# 0.01fF
C2872 a_n392_n100# a_28_n100# 0.02fF
C2873 a_1708_n100# a_1918_n100# 0.03fF
C2874 a_1590_n100# a_2010_n100# 0.02fF
C2875 a_1498_n100# a_2128_n100# 0.01fF
C2876 a_1380_n100# a_2220_n100# 0.01fF
C2877 a_1918_n100# a_3270_n100# 0.00fF
C2878 a_1800_n100# a_3388_n100# 0.00fF
C2879 a_n3540_n632# a_n2608_n632# 0.01fF
C2880 a_n3658_n632# a_n2490_n632# 0.01fF
C2881 a_3270_n100# a_3480_n100# 0.03fF
C2882 a_n3448_n632# a_n2700_n632# 0.01fF
C2883 a_n2190_n100# a_n1980_n100# 0.03fF
C2884 a_n2400_n100# a_n1770_n100# 0.01fF
C2885 a_n2282_n100# a_n1862_n100# 0.02fF
C2886 a_2128_n100# a_540_n100# 0.00fF
C2887 a_4020_n632# a_2642_n632# 0.00fF
C2888 a_4112_n632# a_2550_n632# 0.00fF
C2889 a_1334_n401# a_1124_n729# 0.00fF
C2890 a_870_n632# a_2222_n632# 0.00fF
C2891 a_n136_n729# a_1124_n729# 0.00fF
C2892 a_3178_n100# a_3222_n197# 0.00fF
C2893 a_1290_n632# a_1334_n401# 0.00fF
C2894 a_1920_n632# a_1964_n729# 0.00fF
C2895 w_n4520_n851# a_1170_n100# 0.02fF
C2896 a_1332_131# a_1288_n100# 0.00fF
C2897 a_450_n632# a_492_131# 0.00fF
C2898 a_1592_n632# a_1802_n632# 0.03fF
C2899 a_74_n401# a_1334_n401# 0.00fF
C2900 a_1382_n632# a_2012_n632# 0.01fF
C2901 a_494_n401# a_914_n401# 0.01fF
C2902 a_1500_n632# a_1920_n632# 0.02fF
C2903 a_n2912_n100# a_n2820_n100# 0.09fF
C2904 a_330_n100# a_1170_n100# 0.01fF
C2905 a_n1980_n100# a_n602_n100# 0.00fF
C2906 a_n1560_n100# a_n1022_n100# 0.01fF
C2907 a_n1862_n100# a_n720_n100# 0.01fF
C2908 a_n3240_n100# a_n2492_n100# 0.01fF
C2909 a_n1652_n100# a_n930_n100# 0.01fF
C2910 a_n3030_n100# a_n2702_n100# 0.02fF
C2911 a_n1770_n100# a_n812_n100# 0.01fF
C2912 a_n3122_n100# a_n2610_n100# 0.01fF
C2913 a_962_n632# a_1290_n632# 0.02fF
C2914 a_74_n401# a_n136_n729# 0.00fF
C2915 a_n346_n401# a_284_n729# 0.00fF
C2916 a_n1138_n632# a_n928_n632# 0.03fF
C2917 a_1498_n100# w_n4520_n851# 0.02fF
C2918 w_n4520_n851# a_3600_n632# 0.04fF
C2919 a_240_n632# a_n1020_n632# 0.00fF
C2920 a_122_n632# a_332_n632# 0.03fF
C2921 a_n298_n632# a_n346_n401# 0.00fF
C2922 a_n3240_n100# a_n4080_n100# 0.01fF
C2923 a_n3122_n100# a_n4172_n100# 0.01fF
C2924 a_n3332_n100# a_n3962_n100# 0.01fF
C2925 w_n4520_n851# a_540_n100# 0.02fF
C2926 a_n766_n401# a_284_n729# 0.00fF
C2927 a_702_n197# a_492_131# 0.00fF
C2928 a_2804_n729# a_1544_n729# 0.00fF
C2929 a_1498_n100# a_330_n100# 0.01fF
C2930 a_n3918_n197# a_n3962_n100# 0.00fF
C2931 a_702_n197# a_1542_n197# 0.01fF
C2932 a_660_n632# a_n390_n632# 0.01fF
C2933 w_n4520_n851# a_n3750_n632# 0.04fF
C2934 a_2968_n100# a_3178_n100# 0.03fF
C2935 w_n4520_n851# a_n1348_n632# 0.01fF
C2936 a_330_n100# a_540_n100# 0.03fF
C2937 a_238_n100# a_658_n100# 0.02fF
C2938 a_120_n100# a_750_n100# 0.01fF
C2939 a_28_n100# a_868_n100# 0.01fF
C2940 a_n90_n100# a_960_n100# 0.01fF
C2941 a_n300_n100# a_n346_n401# 0.00fF
C2942 a_752_n632# a_870_n632# 0.07fF
C2943 a_542_n632# a_1080_n632# 0.01fF
C2944 a_660_n632# a_962_n632# 0.02fF
C2945 a_750_n100# a_n720_n100# 0.00fF
C2946 a_2592_131# a_3222_n197# 0.00fF
C2947 a_n510_n100# a_n812_n100# 0.02fF
C2948 a_n392_n100# a_n930_n100# 0.01fF
C2949 a_n300_n100# a_n1022_n100# 0.01fF
C2950 a_n182_n100# a_n1140_n100# 0.01fF
C2951 a_n90_n100# a_n1232_n100# 0.01fF
C2952 a_n3960_n632# a_n3120_n632# 0.01fF
C2953 a_n3750_n632# a_n3330_n632# 0.02fF
C2954 a_n4078_n632# a_n3028_n632# 0.01fF
C2955 a_n4170_n632# a_n2910_n632# 0.00fF
C2956 a_n3868_n632# a_n3238_n632# 0.01fF
C2957 a_4018_n100# a_4062_n197# 0.00fF
C2958 a_n3028_n632# a_n1650_n632# 0.00fF
C2959 a_n3120_n632# a_n1558_n632# 0.00fF
C2960 a_n2910_n632# a_n1768_n632# 0.01fF
C2961 a_n2448_131# a_n2490_n632# 0.00fF
C2962 a_1918_n100# a_658_n100# 0.00fF
C2963 a_n810_n632# a_n2398_n632# 0.00fF
C2964 a_1802_n632# a_2340_n632# 0.01fF
C2965 a_1592_n632# a_2550_n632# 0.01fF
C2966 a_1920_n632# a_2222_n632# 0.02fF
C2967 a_2012_n632# a_2130_n632# 0.07fF
C2968 a_1290_n632# a_2852_n632# 0.00fF
C2969 a_1710_n632# a_2432_n632# 0.01fF
C2970 a_1500_n632# a_2642_n632# 0.01fF
C2971 a_1382_n632# a_2760_n632# 0.00fF
C2972 a_1080_n632# a_1122_n197# 0.00fF
C2973 a_122_n632# a_n508_n632# 0.01fF
C2974 a_2172_131# a_2592_131# 0.01fF
C2975 a_n182_n100# a_448_n100# 0.01fF
C2976 a_n2400_n100# a_n3240_n100# 0.01fF
C2977 a_n2282_n100# a_n3332_n100# 0.01fF
C2978 a_2758_n100# a_2760_n632# 0.00fF
C2979 a_282_n197# a_n558_n197# 0.01fF
C2980 a_3012_131# a_3014_n401# 0.01fF
C2981 a_4020_n632# w_n4520_n851# 0.08fF
C2982 a_2594_n401# a_3014_n401# 0.01fF
C2983 a_n3498_n197# a_n3078_n197# 0.01fF
C2984 a_n4128_131# a_n2658_n197# 0.00fF
C2985 a_494_n401# a_n976_n729# 0.00fF
C2986 a_332_n632# a_n1230_n632# 0.00fF
C2987 w_n4520_n851# a_n3962_n100# 0.06fF
C2988 a_72_131# a_282_n197# 0.00fF
C2989 a_n2702_n100# a_n1350_n100# 0.00fF
C2990 a_n3658_n632# a_n3660_n100# 0.00fF
C2991 a_n2610_n100# a_n1442_n100# 0.01fF
C2992 a_n2820_n100# a_n1232_n100# 0.00fF
C2993 a_n2700_n632# a_n2070_n632# 0.01fF
C2994 a_n2608_n632# a_n2188_n632# 0.02fF
C2995 a_n2490_n632# a_n2280_n632# 0.03fF
C2996 a_2130_n632# a_2760_n632# 0.01fF
C2997 a_2340_n632# a_2550_n632# 0.03fF
C2998 a_2222_n632# a_2642_n632# 0.02fF
C2999 a_752_n632# a_n600_n632# 0.00fF
C3000 a_752_n632# a_1920_n632# 0.01fF
C3001 a_1800_n100# a_1802_n632# 0.00fF
C3002 a_n300_n100# a_1078_n100# 0.00fF
C3003 a_n392_n100# a_1170_n100# 0.00fF
C3004 a_n2868_131# a_n2448_131# 0.01fF
C3005 a_28_n100# a_n1442_n100# 0.00fF
C3006 a_3062_n632# a_3390_n632# 0.02fF
C3007 a_3180_n632# a_3272_n632# 0.09fF
C3008 a_n1818_n197# a_n1816_n729# 0.01fF
C3009 a_n3752_n100# a_n3542_n100# 0.03fF
C3010 a_2220_n100# a_2758_n100# 0.01fF
C3011 a_2128_n100# a_2850_n100# 0.01fF
C3012 a_2010_n100# a_2968_n100# 0.01fF
C3013 a_1918_n100# a_3060_n100# 0.01fF
C3014 a_1800_n100# a_3178_n100# 0.00fF
C3015 a_n3870_n100# a_n3450_n100# 0.02fF
C3016 a_752_n632# a_750_n100# 0.00fF
C3017 a_1708_n100# a_750_n100# 0.01fF
C3018 a_2640_n100# a_3900_n100# 0.00fF
C3019 a_2548_n100# a_4018_n100# 0.00fF
C3020 a_2758_n100# a_3808_n100# 0.01fF
C3021 a_3178_n100# a_3388_n100# 0.03fF
C3022 a_3060_n100# a_3480_n100# 0.02fF
C3023 a_2968_n100# a_3598_n100# 0.01fF
C3024 a_2850_n100# a_3690_n100# 0.01fF
C3025 w_n4520_n851# a_2802_n197# 0.10fF
C3026 a_n390_n632# a_n1348_n632# 0.01fF
C3027 a_n810_n632# a_n928_n632# 0.07fF
C3028 a_n88_n632# a_n1650_n632# 0.00fF
C3029 a_n298_n632# a_n1440_n632# 0.01fF
C3030 a_n718_n632# a_n1020_n632# 0.02fF
C3031 a_n508_n632# a_n1230_n632# 0.01fF
C3032 a_n180_n632# a_n1558_n632# 0.00fF
C3033 a_n600_n632# a_n1138_n632# 0.01fF
C3034 a_240_n632# a_n718_n632# 0.01fF
C3035 a_n2028_131# a_n1818_n197# 0.00fF
C3036 a_240_n632# a_1802_n632# 0.00fF
C3037 a_n392_n100# a_540_n100# 0.01fF
C3038 a_n2282_n100# w_n4520_n851# 0.02fF
C3039 a_3852_131# w_n4520_n851# 0.11fF
C3040 a_2172_131# a_1332_131# 0.01fF
C3041 w_n4520_n851# a_1964_n729# 0.12fF
C3042 a_282_n197# a_1752_131# 0.00fF
C3043 a_1500_n632# w_n4520_n851# 0.01fF
C3044 a_n4170_n632# a_n4078_n632# 0.09fF
C3045 a_2760_n632# a_3692_n632# 0.01fF
C3046 a_2852_n632# a_3600_n632# 0.01fF
C3047 a_2550_n632# a_3902_n632# 0.00fF
C3048 a_2970_n632# a_3482_n632# 0.01fF
C3049 a_2642_n632# a_3810_n632# 0.01fF
C3050 a_n1560_n100# a_n2492_n100# 0.01fF
C3051 a_n1768_n632# a_n1650_n632# 0.07fF
C3052 a_120_n100# w_n4520_n851# 0.02fF
C3053 a_282_n197# a_284_n729# 0.01fF
C3054 a_2850_n100# w_n4520_n851# 0.03fF
C3055 a_n2072_n100# a_n3542_n100# 0.00fF
C3056 a_n2190_n100# a_n3450_n100# 0.00fF
C3057 a_n180_n632# a_30_n632# 0.03fF
C3058 a_3012_131# a_4062_n197# 0.00fF
C3059 w_n4520_n851# a_n720_n100# 0.02fF
C3060 a_n2910_n632# a_n2818_n632# 0.09fF
C3061 a_1172_n632# a_30_n632# 0.01fF
C3062 a_n3708_131# a_n2658_n197# 0.00fF
C3063 a_n2070_n632# a_n1230_n632# 0.01fF
C3064 a_n2398_n632# a_n928_n632# 0.00fF
C3065 a_n1978_n632# a_n1348_n632# 0.01fF
C3066 a_n2280_n632# a_n1020_n632# 0.00fF
C3067 a_n2188_n632# a_n1138_n632# 0.01fF
C3068 a_n1860_n632# a_n1440_n632# 0.02fF
C3069 a_n2238_n197# a_n3498_n197# 0.00fF
C3070 a_870_n632# a_1710_n632# 0.01fF
C3071 a_120_n100# a_330_n100# 0.03fF
C3072 a_868_n100# a_1170_n100# 0.02fF
C3073 a_2430_n100# a_960_n100# 0.00fF
C3074 a_n1188_131# a_n558_n197# 0.00fF
C3075 a_2338_n100# a_2430_n100# 0.09fF
C3076 a_912_131# a_n558_n197# 0.00fF
C3077 a_330_n100# a_n720_n100# 0.01fF
C3078 a_n346_n401# a_n1396_n729# 0.00fF
C3079 a_n1442_n100# a_n930_n100# 0.01fF
C3080 a_n1232_n100# a_n1140_n100# 0.09fF
C3081 a_n1350_n100# a_n1022_n100# 0.02fF
C3082 a_2220_n100# a_1288_n100# 0.01fF
C3083 a_1498_n100# a_868_n100# 0.01fF
C3084 a_n766_n401# a_n1396_n729# 0.00fF
C3085 a_2382_n197# a_1752_131# 0.00fF
C3086 w_n4520_n851# a_n2608_n632# 0.01fF
C3087 w_n4520_n851# a_2222_n632# 0.01fF
C3088 a_2804_n729# a_3434_n401# 0.00fF
C3089 a_n1606_n401# a_n1186_n401# 0.01fF
C3090 a_n2026_n401# a_n766_n401# 0.00fF
C3091 a_332_n632# a_1592_n632# 0.00fF
C3092 a_n182_n100# a_28_n100# 0.03fF
C3093 a_658_n100# a_750_n100# 0.09fF
C3094 a_540_n100# a_868_n100# 0.02fF
C3095 a_448_n100# a_960_n100# 0.01fF
C3096 a_1800_n100# a_2010_n100# 0.03fF
C3097 a_1708_n100# a_2128_n100# 0.02fF
C3098 a_1590_n100# a_2220_n100# 0.01fF
C3099 a_3012_131# a_1542_n197# 0.00fF
C3100 a_72_131# a_n1188_131# 0.00fF
C3101 a_72_131# a_912_131# 0.01fF
C3102 a_1918_n100# a_3480_n100# 0.00fF
C3103 a_2010_n100# a_3388_n100# 0.00fF
C3104 a_2128_n100# a_3270_n100# 0.01fF
C3105 a_n3238_n632# a_n2700_n632# 0.01fF
C3106 a_n3330_n632# a_n2608_n632# 0.01fF
C3107 a_n3448_n632# a_n2490_n632# 0.01fF
C3108 a_n3540_n632# a_n2398_n632# 0.01fF
C3109 a_n3658_n632# a_n2280_n632# 0.00fF
C3110 a_3388_n100# a_3598_n100# 0.03fF
C3111 a_3270_n100# a_3690_n100# 0.02fF
C3112 a_n2072_n100# a_n1862_n100# 0.03fF
C3113 a_n2400_n100# a_n1560_n100# 0.01fF
C3114 a_n2282_n100# a_n1652_n100# 0.01fF
C3115 a_n2190_n100# a_n1770_n100# 0.02fF
C3116 a_4020_n632# a_2852_n632# 0.01fF
C3117 a_4112_n632# a_2760_n632# 0.00fF
C3118 a_n2608_n632# a_n2656_n729# 0.00fF
C3119 a_282_n197# a_702_n197# 0.01fF
C3120 a_1334_n401# a_1964_n729# 0.00fF
C3121 a_2174_n401# a_1124_n729# 0.00fF
C3122 a_1754_n401# a_1544_n729# 0.00fF
C3123 a_870_n632# a_2432_n632# 0.00fF
C3124 a_284_n729# a_1544_n729# 0.00fF
C3125 a_n3288_131# a_n3078_n197# 0.00fF
C3126 a_n2658_n197# a_n1188_131# 0.00fF
C3127 w_n4520_n851# a_494_n401# 0.10fF
C3128 a_n2658_n197# a_n2700_n632# 0.00fF
C3129 a_1172_n632# a_1124_n729# 0.00fF
C3130 a_n810_n632# a_n600_n632# 0.03fF
C3131 a_1080_n632# a_30_n632# 0.01fF
C3132 a_1290_n632# a_n180_n632# 0.00fF
C3133 a_1710_n632# a_1920_n632# 0.03fF
C3134 a_1592_n632# a_2012_n632# 0.02fF
C3135 a_n1770_n100# a_n602_n100# 0.01fF
C3136 a_n1560_n100# a_n812_n100# 0.01fF
C3137 a_n1652_n100# a_n720_n100# 0.01fF
C3138 a_n2820_n100# a_n2702_n100# 0.07fF
C3139 a_n2912_n100# a_n2610_n100# 0.02fF
C3140 a_n3030_n100# a_n2492_n100# 0.01fF
C3141 a_n2868_131# a_n1398_n197# 0.00fF
C3142 a_1172_n632# a_1290_n632# 0.07fF
C3143 a_752_n632# w_n4520_n851# 0.01fF
C3144 a_962_n632# a_1500_n632# 0.01fF
C3145 a_1708_n100# w_n4520_n851# 0.02fF
C3146 w_n4520_n851# a_3810_n632# 0.05fF
C3147 w_n4520_n851# a_3270_n100# 0.03fF
C3148 a_n3122_n100# a_n3962_n100# 0.01fF
C3149 a_n3030_n100# a_n4080_n100# 0.01fF
C3150 a_n3332_n100# a_n3752_n100# 0.02fF
C3151 a_n3240_n100# a_n3870_n100# 0.01fF
C3152 a_n2912_n100# a_n4172_n100# 0.00fF
C3153 a_2804_n729# a_2384_n729# 0.01fF
C3154 a_3224_n729# a_1964_n729# 0.00fF
C3155 a_912_131# a_1752_131# 0.01fF
C3156 a_1708_n100# a_330_n100# 0.00fF
C3157 a_660_n632# a_n180_n632# 0.01fF
C3158 w_n4520_n851# a_n1138_n632# 0.01fF
C3159 a_660_n632# a_1172_n632# 0.01fF
C3160 a_450_n632# a_1382_n632# 0.01fF
C3161 a_n392_n100# a_120_n100# 0.01fF
C3162 a_n90_n100# a_n1022_n100# 0.01fF
C3163 a_n182_n100# a_n930_n100# 0.01fF
C3164 a_n300_n100# a_n812_n100# 0.01fF
C3165 a_n392_n100# a_n720_n100# 0.02fF
C3166 a_n510_n100# a_n602_n100# 0.09fF
C3167 a_n4078_n632# a_n2818_n632# 0.00fF
C3168 a_n3750_n632# a_n3120_n632# 0.01fF
C3169 a_n3960_n632# a_n2910_n632# 0.01fF
C3170 a_n3868_n632# a_n3028_n632# 0.01fF
C3171 a_n3028_n632# a_n1440_n632# 0.00fF
C3172 a_n2818_n632# a_n1650_n632# 0.01fF
C3173 a_n2910_n632# a_n1558_n632# 0.00fF
C3174 a_2128_n100# a_658_n100# 0.00fF
C3175 a_n718_n632# a_n2280_n632# 0.00fF
C3176 a_n810_n632# a_n2188_n632# 0.00fF
C3177 a_1382_n632# a_2970_n632# 0.00fF
C3178 a_1500_n632# a_2852_n632# 0.00fF
C3179 a_1592_n632# a_2760_n632# 0.01fF
C3180 a_1710_n632# a_2642_n632# 0.01fF
C3181 a_2012_n632# a_2340_n632# 0.02fF
C3182 a_1920_n632# a_2432_n632# 0.01fF
C3183 a_1802_n632# a_2550_n632# 0.01fF
C3184 a_n1440_n632# a_n1396_n729# 0.00fF
C3185 a_122_n632# a_n298_n632# 0.02fF
C3186 a_962_n632# a_2222_n632# 0.00fF
C3187 a_n1606_n401# a_n1558_n632# 0.00fF
C3188 a_n2282_n100# a_n3122_n100# 0.01fF
C3189 a_n2072_n100# a_n3332_n100# 0.00fF
C3190 a_n2400_n100# a_n3030_n100# 0.01fF
C3191 a_n2190_n100# a_n3240_n100# 0.01fF
C3192 a_2850_n100# a_2852_n632# 0.00fF
C3193 a_1080_n632# a_1124_n729# 0.00fF
C3194 w_n4520_n851# a_3854_n401# 0.08fF
C3195 a_494_n401# a_1334_n401# 0.01fF
C3196 a_n3658_n632# a_n3448_n632# 0.03fF
C3197 a_3642_n197# a_3690_n100# 0.00fF
C3198 a_494_n401# a_n136_n729# 0.00fF
C3199 a_n346_n401# a_704_n729# 0.00fF
C3200 a_1080_n632# a_1290_n632# 0.03fF
C3201 a_332_n632# a_n1020_n632# 0.00fF
C3202 a_240_n632# a_332_n632# 0.09fF
C3203 a_n3288_131# a_n2238_n197# 0.00fF
C3204 a_122_n632# a_450_n632# 0.02fF
C3205 w_n4520_n851# a_n3752_n100# 0.04fF
C3206 a_n3540_n632# a_n3496_n729# 0.00fF
C3207 a_3852_131# a_3900_n100# 0.00fF
C3208 a_870_n632# a_914_n401# 0.00fF
C3209 a_1172_n632# a_1170_n100# 0.00fF
C3210 w_n4520_n851# a_658_n100# 0.02fF
C3211 a_2220_n100# a_2172_131# 0.00fF
C3212 a_1122_n197# a_492_131# 0.00fF
C3213 a_702_n197# a_912_131# 0.00fF
C3214 a_n766_n401# a_704_n729# 0.00fF
C3215 a_n3706_n401# a_n3658_n632# 0.00fF
C3216 a_n2492_n100# a_n1350_n100# 0.01fF
C3217 a_n3540_n632# a_n3542_n100# 0.00fF
C3218 a_n2610_n100# a_n1232_n100# 0.00fF
C3219 a_n2702_n100# a_n1140_n100# 0.00fF
C3220 a_1122_n197# a_1542_n197# 0.01fF
C3221 a_n2398_n632# a_n2188_n632# 0.03fF
C3222 a_n2490_n632# a_n2070_n632# 0.02fF
C3223 a_n2700_n632# a_n1860_n632# 0.01fF
C3224 a_n2608_n632# a_n1978_n632# 0.01fF
C3225 a_n3916_n729# a_n3076_n729# 0.01fF
C3226 a_2222_n632# a_2852_n632# 0.01fF
C3227 a_2130_n632# a_2970_n632# 0.01fF
C3228 a_2340_n632# a_2760_n632# 0.02fF
C3229 a_2432_n632# a_2642_n632# 0.03fF
C3230 a_752_n632# a_n390_n632# 0.01fF
C3231 a_n3706_n401# a_n3916_n729# 0.00fF
C3232 a_1918_n100# a_1920_n632# 0.00fF
C3233 a_n4126_n401# a_n3496_n729# 0.00fF
C3234 a_660_n632# a_1080_n632# 0.02fF
C3235 a_752_n632# a_962_n632# 0.03fF
C3236 a_330_n100# a_658_n100# 0.02fF
C3237 a_238_n100# a_750_n100# 0.01fF
C3238 a_120_n100# a_868_n100# 0.01fF
C3239 a_28_n100# a_960_n100# 0.01fF
C3240 a_n90_n100# a_1078_n100# 0.01fF
C3241 a_n182_n100# a_1170_n100# 0.00fF
C3242 a_n300_n100# a_1288_n100# 0.00fF
C3243 a_868_n100# a_n720_n100# 0.00fF
C3244 a_28_n100# a_n1232_n100# 0.00fF
C3245 a_3272_n632# a_3390_n632# 0.07fF
C3246 a_3062_n632# a_3600_n632# 0.01fF
C3247 a_3180_n632# a_3482_n632# 0.02fF
C3248 a_n3706_n401# a_n3660_n100# 0.00fF
C3249 a_2592_131# a_2550_n632# 0.00fF
C3250 a_n3660_n100# a_n3450_n100# 0.03fF
C3251 a_2220_n100# a_2968_n100# 0.01fF
C3252 a_2128_n100# a_3060_n100# 0.01fF
C3253 a_2010_n100# a_3178_n100# 0.01fF
C3254 a_1918_n100# a_750_n100# 0.01fF
C3255 a_n928_n632# a_n976_n729# 0.00fF
C3256 a_n4128_131# a_n3498_n197# 0.00fF
C3257 a_2758_n100# a_4018_n100# 0.00fF
C3258 a_3178_n100# a_3598_n100# 0.02fF
C3259 a_3060_n100# a_3690_n100# 0.01fF
C3260 a_2968_n100# a_3808_n100# 0.01fF
C3261 a_2850_n100# a_3900_n100# 0.01fF
C3262 a_2640_n100# a_4110_n100# 0.00fF
C3263 a_1380_n100# a_n90_n100# 0.00fF
C3264 w_n4520_n851# VSUBS 31.73fF
.ends

.subckt latch_pmos_pair sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n632#
+ VSUBS sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100#
Xsky130_fd_pr__pfet_01v8_VCQUSW_0 sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131# VSUBS sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100# sky130_fd_pr__pfet_01v8_VCQUSW
C0 sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851# VSUBS 31.73fF
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VPWR Y VNB VPB a_27_47#
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 VPWR VPB 0.43fF
C1 B a_27_47# 0.33fF
C2 B A 0.16fF
C3 B VPB 0.21fF
C4 Y VPWR 1.44fF
C5 B Y 0.30fF
C6 a_27_47# VGND 0.77fF
C7 A VGND 0.08fF
C8 B VPWR 0.12fF
C9 Y VGND 0.13fF
C10 VPWR VGND 0.12fF
C11 B VGND 0.10fF
C12 A a_27_47# 0.10fF
C13 A VPB 0.18fF
C14 Y a_27_47# 0.41fF
C15 Y A 0.35fF
C16 Y VPB 0.02fF
C17 VPWR a_27_47# 0.07fF
C18 VPWR A 0.09fF
C19 VGND VNB 0.48fF
C20 Y VNB 0.01fF
C21 VPWR VNB 0.18fF
C22 A VNB 0.26fF
C23 B VNB 0.30fF
C24 VPB VNB 0.87fF
C25 a_27_47# VNB 0.06fF
.ends

.subckt sky130_fd_pr__pfet_01v8_VCG74W a_543_n100# a_159_n100# a_n609_n100# a_495_n197#
+ a_n705_n100# a_255_n100# a_n657_n197# a_n369_131# a_351_n100# a_n417_n100# a_n801_n100#
+ a_303_n197# a_n129_n100# a_n513_n100# a_n465_n197# a_n561_131# a_63_n100# a_n225_n100#
+ a_399_131# a_111_n197# a_n321_n100# a_n273_n197# a_15_131# a_n753_131# a_639_n100#
+ w_n1031_n319# a_591_131# a_207_131# a_735_n100# a_n33_n100# a_687_n197# a_447_n100#
+ a_n81_n197# a_n177_131# VSUBS
X0 a_63_n100# a_15_131# a_n33_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n129_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_255_n100# a_207_131# a_159_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_351_n100# a_303_n197# a_255_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_543_n100# a_495_n197# a_447_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 w_n1031_n319# w_n1031_n319# a_735_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=5.24e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6 a_159_n100# a_111_n197# a_63_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_447_n100# a_399_131# a_351_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_639_n100# a_591_131# a_543_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_735_n100# a_687_n197# a_639_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n801_n100# w_n1031_n319# w_n1031_n319# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_n513_n100# a_n561_131# a_n609_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X12 a_n321_n100# a_n369_131# a_n417_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_n225_n100# a_n273_n197# a_n321_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_n705_n100# a_n753_131# a_n801_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_n609_n100# a_n657_n197# a_n705_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n417_n100# a_n465_n197# a_n513_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n129_n100# a_n177_131# a_n225_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_63_n100# a_n513_n100# 0.01fF
C1 a_735_n100# a_n513_n100# 0.00fF
C2 a_207_131# a_687_n197# 0.00fF
C3 a_303_n197# a_n273_n197# 0.01fF
C4 a_159_n100# a_n513_n100# 0.01fF
C5 a_n177_131# a_687_n197# 0.00fF
C6 a_n561_131# a_687_n197# 0.00fF
C7 a_n129_n100# a_n513_n100# 0.02fF
C8 a_n705_n100# a_n609_n100# 0.09fF
C9 a_n753_131# a_n369_131# 0.01fF
C10 a_399_131# a_207_131# 0.04fF
C11 a_495_n197# w_n1031_n319# 0.11fF
C12 a_n753_131# a_n81_n197# 0.00fF
C13 a_399_131# a_n561_131# 0.01fF
C14 a_n177_131# a_399_131# 0.01fF
C15 a_n33_n100# a_n705_n100# 0.01fF
C16 a_63_n100# w_n1031_n319# 0.04fF
C17 a_735_n100# w_n1031_n319# 0.15fF
C18 a_351_n100# a_447_n100# 0.09fF
C19 a_159_n100# w_n1031_n319# 0.04fF
C20 a_n609_n100# a_n657_n197# 0.00fF
C21 a_n129_n100# w_n1031_n319# 0.04fF
C22 a_591_131# a_207_131# 0.01fF
C23 a_n225_n100# a_63_n100# 0.02fF
C24 a_n225_n100# a_735_n100# 0.01fF
C25 a_591_131# a_n177_131# 0.01fF
C26 a_591_131# a_n561_131# 0.00fF
C27 a_159_n100# a_n225_n100# 0.02fF
C28 a_n129_n100# a_n225_n100# 0.09fF
C29 a_351_n100# a_n609_n100# 0.01fF
C30 a_207_131# a_n657_n197# 0.00fF
C31 a_n417_n100# a_n705_n100# 0.02fF
C32 a_n561_131# a_n657_n197# 0.01fF
C33 a_n177_131# a_n657_n197# 0.00fF
C34 a_15_131# a_495_n197# 0.00fF
C35 a_n513_n100# a_n705_n100# 0.04fF
C36 a_447_n100# a_n801_n100# 0.00fF
C37 a_n33_n100# a_351_n100# 0.02fF
C38 a_303_n197# a_207_131# 0.01fF
C39 a_63_n100# a_15_131# 0.00fF
C40 a_687_n197# w_n1031_n319# 0.13fF
C41 a_n177_131# a_303_n197# 0.00fF
C42 a_303_n197# a_n561_131# 0.00fF
C43 a_495_n197# a_111_n197# 0.01fF
C44 a_399_131# w_n1031_n319# 0.12fF
C45 a_n801_n100# a_n609_n100# 0.04fF
C46 a_63_n100# a_111_n197# 0.00fF
C47 a_351_n100# a_n417_n100# 0.01fF
C48 a_n705_n100# w_n1031_n319# 0.08fF
C49 a_n321_n100# a_63_n100# 0.02fF
C50 a_159_n100# a_111_n197# 0.00fF
C51 a_735_n100# a_n321_n100# 0.01fF
C52 a_543_n100# a_447_n100# 0.09fF
C53 a_159_n100# a_n321_n100# 0.01fF
C54 a_63_n100# a_255_n100# 0.04fF
C55 a_n129_n100# a_n321_n100# 0.04fF
C56 a_735_n100# a_255_n100# 0.01fF
C57 a_n33_n100# a_n801_n100# 0.01fF
C58 a_591_131# w_n1031_n319# 0.12fF
C59 a_159_n100# a_255_n100# 0.09fF
C60 a_n225_n100# a_n705_n100# 0.01fF
C61 a_351_n100# a_n513_n100# 0.01fF
C62 a_n129_n100# a_255_n100# 0.02fF
C63 a_15_131# a_687_n197# 0.00fF
C64 a_n369_131# a_495_n197# 0.00fF
C65 a_543_n100# a_n609_n100# 0.01fF
C66 a_n81_n197# a_495_n197# 0.01fF
C67 a_n657_n197# w_n1031_n319# 0.16fF
C68 a_399_131# a_15_131# 0.01fF
C69 a_n417_n100# a_n801_n100# 0.02fF
C70 a_687_n197# a_111_n197# 0.01fF
C71 a_351_n100# w_n1031_n319# 0.05fF
C72 a_n33_n100# a_543_n100# 0.01fF
C73 a_303_n197# w_n1031_n319# 0.11fF
C74 a_n129_n100# a_n81_n197# 0.00fF
C75 a_n801_n100# a_n513_n100# 0.02fF
C76 a_399_131# a_111_n197# 0.00fF
C77 a_591_131# a_15_131# 0.01fF
C78 a_n225_n100# a_351_n100# 0.01fF
C79 a_543_n100# a_n417_n100# 0.01fF
C80 a_n321_n100# a_n705_n100# 0.02fF
C81 a_15_131# a_n657_n197# 0.00fF
C82 a_591_131# a_111_n197# 0.00fF
C83 a_n369_131# a_687_n197# 0.00fF
C84 a_n705_n100# a_255_n100# 0.01fF
C85 a_n81_n197# a_687_n197# 0.01fF
C86 a_n801_n100# w_n1031_n319# 0.15fF
C87 a_n273_n197# a_n465_n197# 0.04fF
C88 a_543_n100# a_n513_n100# 0.01fF
C89 a_639_n100# a_63_n100# 0.01fF
C90 a_303_n197# a_15_131# 0.00fF
C91 a_639_n100# a_735_n100# 0.09fF
C92 a_399_131# a_n369_131# 0.01fF
C93 a_639_n100# a_159_n100# 0.01fF
C94 a_n657_n197# a_111_n197# 0.01fF
C95 a_399_131# a_n81_n197# 0.00fF
C96 a_639_n100# a_n129_n100# 0.01fF
C97 a_n225_n100# a_n801_n100# 0.01fF
C98 a_303_n197# a_111_n197# 0.04fF
C99 a_543_n100# w_n1031_n319# 0.06fF
C100 a_351_n100# a_n321_n100# 0.01fF
C101 a_n753_131# a_495_n197# 0.00fF
C102 a_591_131# a_n369_131# 0.01fF
C103 a_591_131# a_n81_n197# 0.00fF
C104 a_351_n100# a_255_n100# 0.09fF
C105 a_303_n197# a_255_n100# 0.00fF
C106 a_543_n100# a_n225_n100# 0.01fF
C107 a_n369_131# a_n657_n197# 0.00fF
C108 a_n81_n197# a_n657_n197# 0.01fF
C109 a_639_n100# a_687_n197# 0.00fF
C110 a_303_n197# a_n369_131# 0.00fF
C111 a_303_n197# a_n81_n197# 0.01fF
C112 a_207_131# a_n465_n197# 0.00fF
C113 a_n321_n100# a_n801_n100# 0.01fF
C114 a_639_n100# a_n705_n100# 0.00fF
C115 a_n561_131# a_n465_n197# 0.01fF
C116 a_n177_131# a_n465_n197# 0.00fF
C117 a_n801_n100# a_255_n100# 0.01fF
C118 a_591_131# a_639_n100# 0.00fF
C119 a_n753_131# a_687_n197# 0.00fF
C120 a_n273_n197# a_207_131# 0.00fF
C121 a_n417_n100# a_n465_n197# 0.00fF
C122 a_n273_n197# a_n561_131# 0.00fF
C123 a_n177_131# a_n273_n197# 0.01fF
C124 a_399_131# a_n753_131# 0.00fF
C125 a_447_n100# a_n609_n100# 0.01fF
C126 a_543_n100# a_n321_n100# 0.01fF
C127 a_543_n100# a_255_n100# 0.02fF
C128 a_n513_n100# a_n465_n197# 0.00fF
C129 a_n753_131# a_n705_n100# 0.00fF
C130 a_639_n100# a_351_n100# 0.02fF
C131 a_n33_n100# a_447_n100# 0.01fF
C132 a_591_131# a_n753_131# 0.00fF
C133 a_n753_131# a_n657_n197# 0.01fF
C134 a_n465_n197# w_n1031_n319# 0.14fF
C135 a_n33_n100# a_n609_n100# 0.01fF
C136 a_n561_131# a_n609_n100# 0.00fF
C137 a_n417_n100# a_447_n100# 0.01fF
C138 a_639_n100# a_n801_n100# 0.00fF
C139 a_303_n197# a_n753_131# 0.00fF
C140 a_735_n100# a_63_n100# 0.01fF
C141 a_159_n100# a_63_n100# 0.09fF
C142 a_447_n100# a_n513_n100# 0.01fF
C143 a_n273_n197# w_n1031_n319# 0.13fF
C144 a_n177_131# a_207_131# 0.01fF
C145 a_207_131# a_n561_131# 0.01fF
C146 a_159_n100# a_735_n100# 0.01fF
C147 a_n129_n100# a_63_n100# 0.04fF
C148 a_n129_n100# a_735_n100# 0.01fF
C149 a_n417_n100# a_n609_n100# 0.04fF
C150 a_n177_131# a_n561_131# 0.01fF
C151 a_n129_n100# a_159_n100# 0.02fF
C152 a_n225_n100# a_n273_n197# 0.00fF
C153 a_n513_n100# a_n609_n100# 0.09fF
C154 a_15_131# a_n465_n197# 0.00fF
C155 a_n33_n100# a_n417_n100# 0.02fF
C156 a_639_n100# a_543_n100# 0.09fF
C157 a_447_n100# w_n1031_n319# 0.05fF
C158 a_495_n197# a_687_n197# 0.04fF
C159 a_n753_131# a_n801_n100# 0.00fF
C160 a_n33_n100# a_n513_n100# 0.01fF
C161 a_735_n100# a_687_n197# 0.00fF
C162 a_n225_n100# a_447_n100# 0.01fF
C163 a_n465_n197# a_111_n197# 0.01fF
C164 a_n513_n100# a_n561_131# 0.00fF
C165 a_399_131# a_495_n197# 0.01fF
C166 a_n273_n197# a_15_131# 0.00fF
C167 a_n609_n100# w_n1031_n319# 0.06fF
C168 a_n225_n100# a_n609_n100# 0.02fF
C169 a_63_n100# a_n705_n100# 0.01fF
C170 a_591_131# a_495_n197# 0.01fF
C171 a_n273_n197# a_111_n197# 0.01fF
C172 a_735_n100# a_n705_n100# 0.00fF
C173 a_n417_n100# a_n513_n100# 0.09fF
C174 a_n33_n100# w_n1031_n319# 0.04fF
C175 a_207_131# w_n1031_n319# 0.12fF
C176 a_159_n100# a_n705_n100# 0.01fF
C177 a_n321_n100# a_n273_n197# 0.00fF
C178 a_n177_131# w_n1031_n319# 0.13fF
C179 a_n561_131# w_n1031_n319# 0.14fF
C180 a_n129_n100# a_n705_n100# 0.01fF
C181 a_n369_131# a_n465_n197# 0.01fF
C182 a_495_n197# a_n657_n197# 0.00fF
C183 a_n33_n100# a_n225_n100# 0.04fF
C184 a_n81_n197# a_n465_n197# 0.01fF
C185 a_n177_131# a_n225_n100# 0.00fF
C186 a_n417_n100# w_n1031_n319# 0.05fF
C187 a_303_n197# a_495_n197# 0.04fF
C188 a_399_131# a_687_n197# 0.00fF
C189 a_n321_n100# a_447_n100# 0.01fF
C190 a_n273_n197# a_n369_131# 0.01fF
C191 a_n273_n197# a_n81_n197# 0.04fF
C192 a_447_n100# a_255_n100# 0.04fF
C193 a_351_n100# a_63_n100# 0.02fF
C194 a_351_n100# a_735_n100# 0.02fF
C195 a_n225_n100# a_n417_n100# 0.04fF
C196 a_n513_n100# w_n1031_n319# 0.05fF
C197 a_15_131# a_207_131# 0.04fF
C198 a_n33_n100# a_15_131# 0.00fF
C199 a_159_n100# a_351_n100# 0.04fF
C200 a_n129_n100# a_351_n100# 0.01fF
C201 a_15_131# a_n561_131# 0.01fF
C202 a_n177_131# a_15_131# 0.04fF
C203 a_n321_n100# a_n609_n100# 0.02fF
C204 a_591_131# a_687_n197# 0.01fF
C205 a_n225_n100# a_n513_n100# 0.02fF
C206 a_255_n100# a_n609_n100# 0.01fF
C207 a_207_131# a_111_n197# 0.01fF
C208 a_591_131# a_399_131# 0.04fF
C209 a_n657_n197# a_687_n197# 0.00fF
C210 a_n561_131# a_111_n197# 0.00fF
C211 a_n177_131# a_111_n197# 0.00fF
C212 a_n33_n100# a_n321_n100# 0.02fF
C213 a_63_n100# a_n801_n100# 0.01fF
C214 a_n33_n100# a_255_n100# 0.02fF
C215 a_207_131# a_255_n100# 0.00fF
C216 a_735_n100# a_n801_n100# 0.00fF
C217 a_399_131# a_n657_n197# 0.00fF
C218 a_159_n100# a_n801_n100# 0.01fF
C219 a_n225_n100# w_n1031_n319# 0.04fF
C220 a_303_n197# a_687_n197# 0.01fF
C221 a_n129_n100# a_n801_n100# 0.01fF
C222 a_n705_n100# a_n657_n197# 0.00fF
C223 a_n417_n100# a_n321_n100# 0.09fF
C224 a_399_131# a_351_n100# 0.00fF
C225 a_303_n197# a_399_131# 0.01fF
C226 a_543_n100# a_495_n197# 0.00fF
C227 a_n369_131# a_207_131# 0.01fF
C228 a_n753_131# a_n465_n197# 0.00fF
C229 a_591_131# a_n657_n197# 0.00fF
C230 a_n33_n100# a_n81_n197# 0.00fF
C231 a_207_131# a_n81_n197# 0.00fF
C232 a_n417_n100# a_255_n100# 0.01fF
C233 a_n177_131# a_n369_131# 0.04fF
C234 a_n369_131# a_n561_131# 0.04fF
C235 a_351_n100# a_n705_n100# 0.01fF
C236 a_n561_131# a_n81_n197# 0.00fF
C237 a_543_n100# a_63_n100# 0.01fF
C238 a_n177_131# a_n81_n197# 0.01fF
C239 a_543_n100# a_735_n100# 0.04fF
C240 a_n321_n100# a_n513_n100# 0.04fF
C241 a_15_131# w_n1031_n319# 0.12fF
C242 a_543_n100# a_159_n100# 0.02fF
C243 a_639_n100# a_447_n100# 0.04fF
C244 a_n129_n100# a_543_n100# 0.01fF
C245 a_n513_n100# a_255_n100# 0.01fF
C246 a_591_131# a_303_n197# 0.00fF
C247 a_n753_131# a_n273_n197# 0.00fF
C248 a_n417_n100# a_n369_131# 0.00fF
C249 a_303_n197# a_n657_n197# 0.01fF
C250 w_n1031_n319# a_111_n197# 0.12fF
C251 a_639_n100# a_n609_n100# 0.00fF
C252 a_n321_n100# w_n1031_n319# 0.05fF
C253 a_n801_n100# a_n705_n100# 0.09fF
C254 a_255_n100# w_n1031_n319# 0.05fF
C255 a_303_n197# a_351_n100# 0.00fF
C256 a_n225_n100# a_n321_n100# 0.09fF
C257 a_n33_n100# a_639_n100# 0.01fF
C258 a_n225_n100# a_255_n100# 0.01fF
C259 a_n369_131# w_n1031_n319# 0.13fF
C260 a_n81_n197# w_n1031_n319# 0.13fF
C261 a_543_n100# a_n705_n100# 0.00fF
C262 a_15_131# a_111_n197# 0.01fF
C263 a_639_n100# a_n417_n100# 0.01fF
C264 a_351_n100# a_n801_n100# 0.01fF
C265 a_591_131# a_543_n100# 0.00fF
C266 a_n753_131# a_207_131# 0.01fF
C267 a_639_n100# a_n513_n100# 0.01fF
C268 a_n753_131# a_n561_131# 0.04fF
C269 a_n177_131# a_n753_131# 0.01fF
C270 a_495_n197# a_n465_n197# 0.01fF
C271 a_15_131# a_n369_131# 0.01fF
C272 a_15_131# a_n81_n197# 0.01fF
C273 a_n321_n100# a_255_n100# 0.01fF
C274 a_543_n100# a_351_n100# 0.04fF
C275 a_639_n100# w_n1031_n319# 0.08fF
C276 a_n273_n197# a_495_n197# 0.01fF
C277 a_n369_131# a_111_n197# 0.00fF
C278 a_n81_n197# a_111_n197# 0.04fF
C279 a_639_n100# a_n225_n100# 0.01fF
C280 a_n321_n100# a_n369_131# 0.00fF
C281 a_447_n100# a_495_n197# 0.00fF
C282 a_543_n100# a_n801_n100# 0.00fF
C283 a_n465_n197# a_687_n197# 0.00fF
C284 a_n753_131# w_n1031_n319# 0.17fF
C285 a_447_n100# a_63_n100# 0.02fF
C286 a_735_n100# a_447_n100# 0.02fF
C287 a_159_n100# a_447_n100# 0.02fF
C288 a_n369_131# a_n81_n197# 0.00fF
C289 a_399_131# a_n465_n197# 0.00fF
C290 a_n129_n100# a_447_n100# 0.01fF
C291 a_n273_n197# a_687_n197# 0.01fF
C292 a_63_n100# a_n609_n100# 0.01fF
C293 a_735_n100# a_n609_n100# 0.00fF
C294 a_159_n100# a_n609_n100# 0.01fF
C295 a_207_131# a_495_n197# 0.00fF
C296 a_639_n100# a_n321_n100# 0.01fF
C297 a_n129_n100# a_n609_n100# 0.01fF
C298 a_591_131# a_n465_n197# 0.00fF
C299 a_399_131# a_n273_n197# 0.00fF
C300 a_n561_131# a_495_n197# 0.00fF
C301 a_n177_131# a_495_n197# 0.00fF
C302 a_639_n100# a_255_n100# 0.02fF
C303 a_n33_n100# a_63_n100# 0.09fF
C304 a_n753_131# a_15_131# 0.01fF
C305 a_n33_n100# a_735_n100# 0.01fF
C306 a_n33_n100# a_159_n100# 0.04fF
C307 a_159_n100# a_207_131# 0.00fF
C308 a_n657_n197# a_n465_n197# 0.04fF
C309 a_n33_n100# a_n129_n100# 0.09fF
C310 a_n129_n100# a_n177_131# 0.00fF
C311 a_591_131# a_n273_n197# 0.00fF
C312 a_399_131# a_447_n100# 0.00fF
C313 a_n753_131# a_111_n197# 0.00fF
C314 a_303_n197# a_n465_n197# 0.01fF
C315 a_n417_n100# a_63_n100# 0.01fF
C316 a_735_n100# a_n417_n100# 0.01fF
C317 a_n273_n197# a_n657_n197# 0.01fF
C318 a_447_n100# a_n705_n100# 0.01fF
C319 a_159_n100# a_n417_n100# 0.01fF
C320 a_n129_n100# a_n417_n100# 0.02fF
C321 w_n1031_n319# VSUBS 3.95fF
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6625e+11p ps=3.78e+06u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
C0 VPWR X 0.30fF
C1 a_27_47# X 0.26fF
C2 VPWR a_27_47# 0.24fF
C3 VPB X 0.00fF
C4 VPWR VPB 0.24fF
C5 VPB a_27_47# 0.12fF
C6 A X 0.01fF
C7 VGND X 0.19fF
C8 VPWR A 0.02fF
C9 VPWR VGND 0.06fF
C10 A a_27_47# 0.21fF
C11 VGND a_27_47# 0.19fF
C12 A VPB 0.10fF
C13 A VGND 0.02fF
C14 VGND VNB 0.28fF
C15 X VNB 0.00fF
C16 VPWR VNB 0.08fF
C17 A VNB 0.13fF
C18 VPB VNB 0.43fF
C19 a_27_47# VNB 0.15fF
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
C0 VGND VPWR 3.03fF
C1 VPB VPWR 0.47fF
C2 VGND VPB 0.87fF
C3 VPWR VNB 1.33fF
C4 VGND VNB 0.77fF
C5 VPB VNB 1.14fF
.ends

.subckt precharge_pmos sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131#
+ VSUBS
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ VSUBS sky130_fd_pr__pfet_01v8_VCG74W
C0 sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319# VSUBS 3.95fF
.ends

.subckt current_tail a_543_n100# a_159_n100# a_n609_n100# a_n1569_n100# a_n705_n100#
+ a_255_n100# a_1407_n100# a_351_n100# a_n417_n100# a_n801_n100# a_1503_n100# a_1119_n100#
+ a_n1377_n100# a_n129_n100# a_n513_n100# a_1215_n100# a_63_n100# a_n1089_n100# a_n1473_n100#
+ a_n225_n100# a_1311_n100# a_927_n100# a_n1185_n100# a_n321_n100# a_1023_n100# a_639_n100#
+ a_n1281_n100# a_735_n100# a_n33_n100# a_n897_n100# a_831_n100# a_447_n100# a_n1521_122#
+ a_n993_n100# a_n1763_n274#
X0 a_n801_n100# a_n1521_122# a_n897_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n513_n100# a_n1521_122# a_n609_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n321_n100# a_n1521_122# a_n417_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_n225_n100# a_n1521_122# a_n321_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_n897_n100# a_n1521_122# a_n993_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 a_n705_n100# a_n1521_122# a_n801_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_n609_n100# a_n1521_122# a_n705_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n417_n100# a_n1521_122# a_n513_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n129_n100# a_n1521_122# a_n225_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_63_n100# a_n1521_122# a_n33_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_927_n100# a_n1521_122# a_831_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11 a_1023_n100# a_n1521_122# a_927_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_n1569_n100# a_n1763_n274# a_n1763_n274# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=6.2e+11p ps=5.24e+06u w=1e+06u l=150000u
X13 a_1119_n100# a_n1521_122# a_1023_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_1215_n100# a_n1521_122# a_1119_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_1311_n100# a_n1521_122# a_1215_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_1407_n100# a_n1521_122# a_1311_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17 a_1503_n100# a_n1521_122# a_1407_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1763_n274# a_n1763_n274# a_1503_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n33_n100# a_n1521_122# a_n129_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_351_n100# a_n1521_122# a_255_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X21 a_159_n100# a_n1521_122# a_63_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22 a_255_n100# a_n1521_122# a_159_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_447_n100# a_n1521_122# a_351_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X24 a_543_n100# a_n1521_122# a_447_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X25 a_639_n100# a_n1521_122# a_543_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X26 a_735_n100# a_n1521_122# a_639_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_831_n100# a_n1521_122# a_735_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n1473_n100# a_n1521_122# a_n1569_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X29 a_n1377_n100# a_n1521_122# a_n1473_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X30 a_n1281_n100# a_n1521_122# a_n1377_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X31 a_n1185_n100# a_n1521_122# a_n1281_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X32 a_n1089_n100# a_n1521_122# a_n1185_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X33 a_n993_n100# a_n1521_122# a_n1089_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_1311_n100# a_735_n100# 0.01fF
C1 a_n609_n100# a_n321_n100# 0.02fF
C2 a_63_n100# a_n897_n100# 0.01fF
C3 a_n129_n100# a_n1185_n100# 0.01fF
C4 a_n513_n100# a_735_n100# 0.00fF
C5 a_n609_n100# a_831_n100# 0.00fF
C6 a_639_n100# a_735_n100# 0.09fF
C7 a_1023_n100# a_n129_n100# 0.01fF
C8 a_1119_n100# a_n225_n100# 0.00fF
C9 a_n1569_n100# a_n1185_n100# 0.02fF
C10 a_n705_n100# a_n225_n100# 0.01fF
C11 a_1503_n100# a_63_n100# 0.00fF
C12 a_n705_n100# a_n1521_122# 0.03fF
C13 a_n225_n100# a_447_n100# 0.01fF
C14 a_255_n100# a_n1281_n100# 0.00fF
C15 a_447_n100# a_n1521_122# 0.03fF
C16 a_n417_n100# a_n897_n100# 0.01fF
C17 a_n321_n100# a_63_n100# 0.02fF
C18 a_63_n100# a_831_n100# 0.01fF
C19 a_159_n100# a_735_n100# 0.01fF
C20 a_1311_n100# a_255_n100# 0.01fF
C21 a_927_n100# a_543_n100# 0.02fF
C22 a_1215_n100# a_351_n100# 0.01fF
C23 a_1407_n100# a_1311_n100# 0.09fF
C24 a_n513_n100# a_255_n100# 0.01fF
C25 a_255_n100# a_639_n100# 0.02fF
C26 a_1407_n100# a_639_n100# 0.01fF
C27 a_n33_n100# a_n1473_n100# 0.00fF
C28 a_255_n100# a_n993_n100# 0.00fF
C29 a_n417_n100# a_n321_n100# 0.09fF
C30 a_n129_n100# a_n1089_n100# 0.01fF
C31 a_n417_n100# a_831_n100# 0.00fF
C32 a_1119_n100# a_n33_n100# 0.01fF
C33 a_n1281_n100# a_n801_n100# 0.01fF
C34 a_1215_n100# a_n225_n100# 0.00fF
C35 a_n1569_n100# a_n1089_n100# 0.01fF
C36 a_1215_n100# a_n1521_122# 0.03fF
C37 a_n705_n100# a_n33_n100# 0.01fF
C38 a_n705_n100# a_n1473_n100# 0.01fF
C39 a_159_n100# a_255_n100# 0.09fF
C40 a_n129_n100# a_543_n100# 0.01fF
C41 a_n33_n100# a_447_n100# 0.01fF
C42 a_1407_n100# a_159_n100# 0.00fF
C43 a_351_n100# a_n1281_n100# 0.00fF
C44 a_n1185_n100# a_n1089_n100# 0.09fF
C45 a_n513_n100# a_n801_n100# 0.02fF
C46 a_639_n100# a_n801_n100# 0.00fF
C47 a_735_n100# a_n897_n100# 0.00fF
C48 a_927_n100# a_n609_n100# 0.00fF
C49 a_1119_n100# a_447_n100# 0.01fF
C50 a_1023_n100# a_543_n100# 0.01fF
C51 a_1311_n100# a_351_n100# 0.01fF
C52 a_n993_n100# a_n801_n100# 0.04fF
C53 a_1503_n100# a_735_n100# 0.01fF
C54 a_n705_n100# a_447_n100# 0.01fF
C55 a_n513_n100# a_351_n100# 0.01fF
C56 a_351_n100# a_639_n100# 0.02fF
C57 a_n129_n100# a_n1377_n100# 0.00fF
C58 a_n225_n100# a_n1281_n100# 0.01fF
C59 a_n1569_n100# a_n1377_n100# 0.04fF
C60 a_n1521_122# a_n1281_n100# 0.03fF
C61 a_351_n100# a_n993_n100# 0.00fF
C62 a_159_n100# a_n801_n100# 0.01fF
C63 a_n321_n100# a_735_n100# 0.01fF
C64 a_735_n100# a_831_n100# 0.09fF
C65 a_927_n100# a_63_n100# 0.01fF
C66 a_1311_n100# a_n225_n100# 0.00fF
C67 a_1215_n100# a_n33_n100# 0.00fF
C68 a_n1377_n100# a_n1185_n100# 0.04fF
C69 a_n513_n100# a_n225_n100# 0.02fF
C70 a_255_n100# a_n897_n100# 0.01fF
C71 a_n609_n100# a_n129_n100# 0.01fF
C72 a_n225_n100# a_639_n100# 0.01fF
C73 a_n609_n100# a_n1569_n100# 0.01fF
C74 a_n513_n100# a_n1521_122# 0.03fF
C75 a_639_n100# a_n1521_122# 0.03fF
C76 a_159_n100# a_351_n100# 0.04fF
C77 a_1503_n100# a_255_n100# 0.00fF
C78 a_n225_n100# a_n993_n100# 0.01fF
C79 a_1407_n100# a_1503_n100# 0.09fF
C80 a_1119_n100# a_1215_n100# 0.09fF
C81 a_n609_n100# a_n1185_n100# 0.01fF
C82 a_927_n100# a_n417_n100# 0.00fF
C83 a_1023_n100# a_n609_n100# 0.00fF
C84 a_543_n100# a_n1089_n100# 0.00fF
C85 a_1215_n100# a_447_n100# 0.01fF
C86 a_n321_n100# a_255_n100# 0.01fF
C87 a_n129_n100# a_63_n100# 0.04fF
C88 a_n225_n100# a_159_n100# 0.02fF
C89 a_255_n100# a_831_n100# 0.01fF
C90 a_63_n100# a_n1569_n100# 0.00fF
C91 a_1407_n100# a_831_n100# 0.01fF
C92 a_n33_n100# a_n1281_n100# 0.00fF
C93 a_n1473_n100# a_n1281_n100# 0.04fF
C94 a_n897_n100# a_n801_n100# 0.09fF
C95 a_63_n100# a_n1185_n100# 0.00fF
C96 a_1023_n100# a_63_n100# 0.01fF
C97 a_1311_n100# a_n33_n100# 0.00fF
C98 a_n1377_n100# a_n1089_n100# 0.02fF
C99 a_351_n100# a_n897_n100# 0.00fF
C100 a_n513_n100# a_n33_n100# 0.01fF
C101 a_n417_n100# a_n129_n100# 0.02fF
C102 a_n33_n100# a_639_n100# 0.01fF
C103 a_n513_n100# a_n1473_n100# 0.01fF
C104 a_n705_n100# a_n1281_n100# 0.01fF
C105 a_n417_n100# a_n1569_n100# 0.01fF
C106 a_1503_n100# a_351_n100# 0.01fF
C107 a_n33_n100# a_n993_n100# 0.01fF
C108 a_n1473_n100# a_n993_n100# 0.01fF
C109 a_1119_n100# a_1311_n100# 0.04fF
C110 a_n321_n100# a_n801_n100# 0.01fF
C111 a_n417_n100# a_n1185_n100# 0.01fF
C112 a_831_n100# a_n801_n100# 0.00fF
C113 a_n609_n100# a_n1089_n100# 0.01fF
C114 a_1119_n100# a_n513_n100# 0.00fF
C115 a_1023_n100# a_n417_n100# 0.00fF
C116 a_927_n100# a_735_n100# 0.04fF
C117 a_1119_n100# a_639_n100# 0.01fF
C118 a_1311_n100# a_447_n100# 0.01fF
C119 a_n225_n100# a_n897_n100# 0.01fF
C120 a_n705_n100# a_n513_n100# 0.04fF
C121 a_n705_n100# a_639_n100# 0.00fF
C122 a_n1521_122# a_n897_n100# 0.03fF
C123 a_n609_n100# a_543_n100# 0.01fF
C124 a_n513_n100# a_447_n100# 0.01fF
C125 a_n321_n100# a_351_n100# 0.01fF
C126 a_n33_n100# a_159_n100# 0.04fF
C127 a_351_n100# a_831_n100# 0.01fF
C128 a_447_n100# a_639_n100# 0.04fF
C129 a_159_n100# a_n1473_n100# 0.00fF
C130 a_n705_n100# a_n993_n100# 0.02fF
C131 a_447_n100# a_n993_n100# 0.00fF
C132 a_63_n100# a_n1089_n100# 0.01fF
C133 a_1119_n100# a_159_n100# 0.01fF
C134 a_n321_n100# a_n225_n100# 0.09fF
C135 a_n705_n100# a_159_n100# 0.01fF
C136 a_n225_n100# a_831_n100# 0.01fF
C137 a_n129_n100# a_735_n100# 0.01fF
C138 a_n321_n100# a_n1521_122# 0.03fF
C139 a_927_n100# a_255_n100# 0.01fF
C140 a_n609_n100# a_n1377_n100# 0.01fF
C141 a_831_n100# a_n1521_122# 0.03fF
C142 a_1407_n100# a_927_n100# 0.01fF
C143 a_63_n100# a_543_n100# 0.01fF
C144 a_159_n100# a_447_n100# 0.02fF
C145 a_1215_n100# a_1311_n100# 0.09fF
C146 a_n417_n100# a_n1089_n100# 0.01fF
C147 a_1023_n100# a_735_n100# 0.02fF
C148 a_1215_n100# a_639_n100# 0.01fF
C149 a_n33_n100# a_n897_n100# 0.01fF
C150 a_n1473_n100# a_n897_n100# 0.01fF
C151 a_n417_n100# a_543_n100# 0.01fF
C152 a_63_n100# a_n1377_n100# 0.00fF
C153 a_1503_n100# a_n33_n100# 0.00fF
C154 a_n129_n100# a_255_n100# 0.02fF
C155 a_1407_n100# a_n129_n100# 0.00fF
C156 a_1215_n100# a_159_n100# 0.01fF
C157 a_n705_n100# a_n897_n100# 0.04fF
C158 a_1503_n100# a_1119_n100# 0.02fF
C159 a_n321_n100# a_n33_n100# 0.02fF
C160 a_447_n100# a_n897_n100# 0.00fF
C161 a_n609_n100# a_63_n100# 0.01fF
C162 a_n33_n100# a_831_n100# 0.01fF
C163 a_255_n100# a_n1185_n100# 0.00fF
C164 a_n513_n100# a_n1281_n100# 0.01fF
C165 a_n321_n100# a_n1473_n100# 0.01fF
C166 a_927_n100# a_351_n100# 0.01fF
C167 a_n417_n100# a_n1377_n100# 0.01fF
C168 a_1023_n100# a_255_n100# 0.01fF
C169 a_1407_n100# a_1023_n100# 0.02fF
C170 a_1503_n100# a_447_n100# 0.01fF
C171 a_n1281_n100# a_n993_n100# 0.02fF
C172 a_1119_n100# a_n321_n100# 0.00fF
C173 a_1119_n100# a_831_n100# 0.02fF
C174 a_1311_n100# a_639_n100# 0.01fF
C175 a_n609_n100# a_n417_n100# 0.04fF
C176 a_n705_n100# a_n321_n100# 0.02fF
C177 a_n129_n100# a_n801_n100# 0.01fF
C178 a_n705_n100# a_831_n100# 0.00fF
C179 a_n513_n100# a_639_n100# 0.01fF
C180 a_927_n100# a_n225_n100# 0.01fF
C181 a_n1569_n100# a_n801_n100# 0.01fF
C182 a_n321_n100# a_447_n100# 0.01fF
C183 a_543_n100# a_735_n100# 0.04fF
C184 a_447_n100# a_831_n100# 0.02fF
C185 a_159_n100# a_n1281_n100# 0.00fF
C186 a_n513_n100# a_n993_n100# 0.01fF
C187 a_639_n100# a_n993_n100# 0.00fF
C188 a_n129_n100# a_351_n100# 0.01fF
C189 a_n1185_n100# a_n801_n100# 0.02fF
C190 a_1311_n100# a_159_n100# 0.01fF
C191 a_1503_n100# a_1215_n100# 0.02fF
C192 a_n513_n100# a_159_n100# 0.01fF
C193 a_n417_n100# a_63_n100# 0.01fF
C194 a_351_n100# a_n1185_n100# 0.00fF
C195 a_255_n100# a_n1089_n100# 0.00fF
C196 a_159_n100# a_639_n100# 0.01fF
C197 a_1023_n100# a_351_n100# 0.01fF
C198 a_159_n100# a_n993_n100# 0.01fF
C199 a_n225_n100# a_n129_n100# 0.09fF
C200 a_n129_n100# a_n1521_122# 0.03fF
C201 a_n225_n100# a_n1569_n100# 0.00fF
C202 a_255_n100# a_543_n100# 0.02fF
C203 a_1407_n100# a_543_n100# 0.01fF
C204 a_1215_n100# a_n321_n100# 0.00fF
C205 a_1215_n100# a_831_n100# 0.02fF
C206 a_n609_n100# a_735_n100# 0.00fF
C207 a_n225_n100# a_n1185_n100# 0.01fF
C208 a_1023_n100# a_n225_n100# 0.00fF
C209 a_927_n100# a_n33_n100# 0.01fF
C210 a_n1281_n100# a_n897_n100# 0.02fF
C211 a_1023_n100# a_n1521_122# 0.03fF
C212 a_255_n100# a_n1377_n100# 0.00fF
C213 a_n1089_n100# a_n801_n100# 0.02fF
C214 a_927_n100# a_1119_n100# 0.04fF
C215 a_n513_n100# a_n897_n100# 0.02fF
C216 a_639_n100# a_n897_n100# 0.00fF
C217 a_1503_n100# a_1311_n100# 0.04fF
C218 a_927_n100# a_n705_n100# 0.00fF
C219 a_543_n100# a_n801_n100# 0.00fF
C220 a_351_n100# a_n1089_n100# 0.00fF
C221 a_63_n100# a_735_n100# 0.01fF
C222 a_n321_n100# a_n1281_n100# 0.01fF
C223 a_927_n100# a_447_n100# 0.01fF
C224 a_n993_n100# a_n897_n100# 0.09fF
C225 a_1503_n100# a_639_n100# 0.01fF
C226 a_n129_n100# a_n33_n100# 0.09fF
C227 a_n609_n100# a_255_n100# 0.01fF
C228 a_n129_n100# a_n1473_n100# 0.00fF
C229 a_n33_n100# a_n1569_n100# 0.00fF
C230 a_351_n100# a_543_n100# 0.04fF
C231 a_n1569_n100# a_n1473_n100# 0.09fF
C232 a_1311_n100# a_n321_n100# 0.00fF
C233 a_1311_n100# a_831_n100# 0.01fF
C234 a_159_n100# a_n897_n100# 0.01fF
C235 a_n513_n100# a_n321_n100# 0.04fF
C236 a_n225_n100# a_n1089_n100# 0.01fF
C237 a_n417_n100# a_735_n100# 0.01fF
C238 a_n321_n100# a_639_n100# 0.01fF
C239 a_n513_n100# a_831_n100# 0.00fF
C240 a_n33_n100# a_n1185_n100# 0.01fF
C241 a_639_n100# a_831_n100# 0.04fF
C242 a_1119_n100# a_n129_n100# 0.00fF
C243 a_1023_n100# a_n33_n100# 0.01fF
C244 a_n1377_n100# a_n801_n100# 0.01fF
C245 a_n1521_122# a_n1089_n100# 0.03fF
C246 a_n1473_n100# a_n1185_n100# 0.02fF
C247 a_1503_n100# a_159_n100# 0.00fF
C248 a_n705_n100# a_n129_n100# 0.01fF
C249 a_n321_n100# a_n993_n100# 0.01fF
C250 a_n705_n100# a_n1569_n100# 0.01fF
C251 a_n225_n100# a_543_n100# 0.01fF
C252 a_63_n100# a_255_n100# 0.04fF
C253 a_n129_n100# a_447_n100# 0.01fF
C254 a_1407_n100# a_63_n100# 0.00fF
C255 a_1023_n100# a_1119_n100# 0.09fF
C256 a_927_n100# a_1215_n100# 0.02fF
C257 a_n609_n100# a_n801_n100# 0.04fF
C258 a_n705_n100# a_n1185_n100# 0.01fF
C259 a_n321_n100# a_159_n100# 0.01fF
C260 a_447_n100# a_n1185_n100# 0.00fF
C261 a_159_n100# a_831_n100# 0.01fF
C262 a_1023_n100# a_447_n100# 0.01fF
C263 a_n417_n100# a_255_n100# 0.01fF
C264 a_n609_n100# a_351_n100# 0.01fF
C265 a_n225_n100# a_n1377_n100# 0.01fF
C266 a_63_n100# a_n801_n100# 0.01fF
C267 a_n33_n100# a_n1089_n100# 0.01fF
C268 a_1215_n100# a_n129_n100# 0.00fF
C269 a_n1473_n100# a_n1089_n100# 0.02fF
C270 a_n609_n100# a_n225_n100# 0.02fF
C271 a_63_n100# a_351_n100# 0.02fF
C272 a_n33_n100# a_543_n100# 0.01fF
C273 a_1023_n100# a_1215_n100# 0.04fF
C274 a_927_n100# a_1311_n100# 0.02fF
C275 a_n417_n100# a_n801_n100# 0.02fF
C276 a_n321_n100# a_n897_n100# 0.01fF
C277 a_n705_n100# a_n1089_n100# 0.02fF
C278 a_927_n100# a_n513_n100# 0.00fF
C279 a_927_n100# a_639_n100# 0.02fF
C280 a_447_n100# a_n1089_n100# 0.00fF
C281 a_1119_n100# a_543_n100# 0.01fF
C282 a_1503_n100# a_831_n100# 0.01fF
C283 a_n705_n100# a_543_n100# 0.00fF
C284 a_n417_n100# a_351_n100# 0.01fF
C285 a_n225_n100# a_63_n100# 0.02fF
C286 a_255_n100# a_735_n100# 0.01fF
C287 a_1407_n100# a_735_n100# 0.01fF
C288 a_n33_n100# a_n1377_n100# 0.00fF
C289 a_n129_n100# a_n1281_n100# 0.01fF
C290 a_63_n100# a_n1521_122# 0.03fF
C291 a_447_n100# a_543_n100# 0.09fF
C292 a_n1569_n100# a_n1281_n100# 0.02fF
C293 a_n1473_n100# a_n1377_n100# 0.09fF
C294 a_n321_n100# a_831_n100# 0.01fF
C295 a_927_n100# a_159_n100# 0.01fF
C296 a_1311_n100# a_n129_n100# 0.00fF
C297 a_n1281_n100# a_n1185_n100# 0.09fF
C298 a_n417_n100# a_n225_n100# 0.04fF
C299 a_n513_n100# a_n129_n100# 0.02fF
C300 a_n609_n100# a_n33_n100# 0.01fF
C301 a_n129_n100# a_639_n100# 0.01fF
C302 a_n705_n100# a_n1377_n100# 0.01fF
C303 a_n609_n100# a_n1473_n100# 0.01fF
C304 a_n513_n100# a_n1569_n100# 0.01fF
C305 a_n129_n100# a_n993_n100# 0.01fF
C306 a_n1569_n100# a_n993_n100# 0.01fF
C307 a_1023_n100# a_1311_n100# 0.02fF
C308 a_1407_n100# a_255_n100# 0.01fF
C309 a_735_n100# a_n801_n100# 0.00fF
C310 a_n513_n100# a_n1185_n100# 0.01fF
C311 a_1023_n100# a_n513_n100# 0.00fF
C312 a_1023_n100# a_639_n100# 0.02fF
C313 a_1215_n100# a_543_n100# 0.01fF
C314 a_n705_n100# a_n609_n100# 0.09fF
C315 a_n1185_n100# a_n993_n100# 0.04fF
C316 a_n609_n100# a_447_n100# 0.01fF
C317 a_n129_n100# a_159_n100# 0.02fF
C318 a_n33_n100# a_63_n100# 0.09fF
C319 a_351_n100# a_735_n100# 0.02fF
C320 a_63_n100# a_n1473_n100# 0.00fF
C321 a_159_n100# a_n1185_n100# 0.00fF
C322 a_1023_n100# a_159_n100# 0.01fF
C323 a_1119_n100# a_63_n100# 0.01fF
C324 a_n1281_n100# a_n1089_n100# 0.04fF
C325 a_1503_n100# a_927_n100# 0.01fF
C326 a_n705_n100# a_63_n100# 0.01fF
C327 a_255_n100# a_n801_n100# 0.01fF
C328 a_n417_n100# a_n33_n100# 0.02fF
C329 a_n225_n100# a_735_n100# 0.01fF
C330 a_n417_n100# a_n1473_n100# 0.01fF
C331 a_63_n100# a_447_n100# 0.02fF
C332 a_255_n100# a_351_n100# 0.09fF
C333 a_1407_n100# a_351_n100# 0.01fF
C334 a_n513_n100# a_n1089_n100# 0.01fF
C335 a_1119_n100# a_n417_n100# 0.00fF
C336 a_927_n100# a_n321_n100# 0.00fF
C337 a_927_n100# a_831_n100# 0.09fF
C338 a_1311_n100# a_543_n100# 0.01fF
C339 a_n129_n100# a_n897_n100# 0.01fF
C340 a_n705_n100# a_n417_n100# 0.02fF
C341 a_n1089_n100# a_n993_n100# 0.09fF
C342 a_n1569_n100# a_n897_n100# 0.01fF
C343 a_n417_n100# a_447_n100# 0.01fF
C344 a_n513_n100# a_543_n100# 0.01fF
C345 a_543_n100# a_639_n100# 0.09fF
C346 a_1503_n100# a_n129_n100# 0.00fF
C347 a_n1377_n100# a_n1281_n100# 0.09fF
C348 a_543_n100# a_n993_n100# 0.00fF
C349 a_n225_n100# a_255_n100# 0.01fF
C350 a_1407_n100# a_n225_n100# 0.00fF
C351 a_255_n100# a_n1521_122# 0.03fF
C352 a_1407_n100# a_n1521_122# 0.03fF
C353 a_n1185_n100# a_n897_n100# 0.02fF
C354 a_159_n100# a_n1089_n100# 0.00fF
C355 a_1215_n100# a_63_n100# 0.01fF
C356 a_1503_n100# a_1023_n100# 0.01fF
C357 a_n321_n100# a_n129_n100# 0.04fF
C358 a_351_n100# a_n801_n100# 0.01fF
C359 a_n129_n100# a_831_n100# 0.01fF
C360 a_n33_n100# a_735_n100# 0.01fF
C361 a_n609_n100# a_n1281_n100# 0.01fF
C362 a_n321_n100# a_n1569_n100# 0.00fF
C363 a_n513_n100# a_n1377_n100# 0.01fF
C364 a_159_n100# a_543_n100# 0.02fF
C365 a_n1377_n100# a_n993_n100# 0.02fF
C366 a_n321_n100# a_n1185_n100# 0.01fF
C367 a_1215_n100# a_n417_n100# 0.00fF
C368 a_1023_n100# a_n321_n100# 0.00fF
C369 a_1023_n100# a_831_n100# 0.04fF
C370 a_1119_n100# a_735_n100# 0.02fF
C371 a_n609_n100# a_n513_n100# 0.09fF
C372 a_n225_n100# a_n801_n100# 0.01fF
C373 a_n609_n100# a_639_n100# 0.00fF
C374 a_n705_n100# a_735_n100# 0.00fF
C375 a_447_n100# a_735_n100# 0.02fF
C376 a_63_n100# a_n1281_n100# 0.00fF
C377 a_159_n100# a_n1377_n100# 0.00fF
C378 a_n609_n100# a_n993_n100# 0.02fF
C379 a_n225_n100# a_351_n100# 0.01fF
C380 a_n33_n100# a_255_n100# 0.02fF
C381 a_1407_n100# a_n33_n100# 0.00fF
C382 a_n1089_n100# a_n897_n100# 0.04fF
C383 a_1311_n100# a_63_n100# 0.00fF
C384 a_543_n100# a_n897_n100# 0.00fF
C385 a_n609_n100# a_159_n100# 0.01fF
C386 a_n513_n100# a_63_n100# 0.01fF
C387 a_63_n100# a_639_n100# 0.01fF
C388 a_n417_n100# a_n1281_n100# 0.01fF
C389 a_1119_n100# a_255_n100# 0.01fF
C390 a_1407_n100# a_1119_n100# 0.02fF
C391 a_1503_n100# a_543_n100# 0.01fF
C392 a_63_n100# a_n993_n100# 0.01fF
C393 a_n705_n100# a_255_n100# 0.01fF
C394 a_255_n100# a_447_n100# 0.04fF
C395 a_1407_n100# a_447_n100# 0.01fF
C396 a_n321_n100# a_n1089_n100# 0.01fF
C397 a_1215_n100# a_735_n100# 0.01fF
C398 a_n513_n100# a_n417_n100# 0.09fF
C399 a_n33_n100# a_n801_n100# 0.01fF
C400 a_n417_n100# a_639_n100# 0.01fF
C401 a_n1377_n100# a_n897_n100# 0.01fF
C402 a_927_n100# a_n129_n100# 0.01fF
C403 a_n1473_n100# a_n801_n100# 0.01fF
C404 a_63_n100# a_159_n100# 0.09fF
C405 a_n321_n100# a_543_n100# 0.01fF
C406 a_543_n100# a_831_n100# 0.02fF
C407 a_n417_n100# a_n993_n100# 0.01fF
C408 a_n33_n100# a_351_n100# 0.02fF
C409 a_927_n100# a_1023_n100# 0.09fF
C410 a_n705_n100# a_n801_n100# 0.09fF
C411 a_n609_n100# a_n897_n100# 0.02fF
C412 a_447_n100# a_n801_n100# 0.00fF
C413 a_n417_n100# a_159_n100# 0.01fF
C414 a_1215_n100# a_255_n100# 0.01fF
C415 a_1119_n100# a_351_n100# 0.01fF
C416 a_n321_n100# a_n1377_n100# 0.01fF
C417 a_1407_n100# a_1215_n100# 0.04fF
C418 a_n225_n100# a_n33_n100# 0.04fF
C419 a_n705_n100# a_351_n100# 0.01fF
C420 a_n129_n100# a_n1569_n100# 0.00fF
C421 a_n225_n100# a_n1473_n100# 0.00fF
C422 a_n1521_122# a_n1473_n100# 0.03fF
C423 a_351_n100# a_447_n100# 0.09fF
C424 a_1503_n100# a_n1763_n274# 0.14fF
C425 a_1407_n100# a_n1763_n274# 0.07fF
C426 a_1311_n100# a_n1763_n274# 0.06fF
C427 a_1215_n100# a_n1763_n274# 0.05fF
C428 a_1119_n100# a_n1763_n274# 0.04fF
C429 a_1023_n100# a_n1763_n274# 0.04fF
C430 a_927_n100# a_n1763_n274# 0.03fF
C431 a_831_n100# a_n1763_n274# 0.03fF
C432 a_735_n100# a_n1763_n274# 0.03fF
C433 a_639_n100# a_n1763_n274# 0.03fF
C434 a_543_n100# a_n1763_n274# 0.03fF
C435 a_447_n100# a_n1763_n274# 0.03fF
C436 a_351_n100# a_n1763_n274# 0.03fF
C437 a_255_n100# a_n1763_n274# 0.03fF
C438 a_159_n100# a_n1763_n274# 0.03fF
C439 a_63_n100# a_n1763_n274# 0.02fF
C440 a_n33_n100# a_n1763_n274# 0.03fF
C441 a_n129_n100# a_n1763_n274# 0.02fF
C442 a_n225_n100# a_n1763_n274# 0.03fF
C443 a_n321_n100# a_n1763_n274# 0.03fF
C444 a_n417_n100# a_n1763_n274# 0.03fF
C445 a_n513_n100# a_n1763_n274# 0.03fF
C446 a_n609_n100# a_n1763_n274# 0.03fF
C447 a_n705_n100# a_n1763_n274# 0.03fF
C448 a_n801_n100# a_n1763_n274# 0.03fF
C449 a_n897_n100# a_n1763_n274# 0.03fF
C450 a_n993_n100# a_n1763_n274# 0.03fF
C451 a_n1089_n100# a_n1763_n274# 0.04fF
C452 a_n1185_n100# a_n1763_n274# 0.04fF
C453 a_n1281_n100# a_n1763_n274# 0.05fF
C454 a_n1377_n100# a_n1763_n274# 0.06fF
C455 a_n1473_n100# a_n1763_n274# 0.08fF
C456 a_n1569_n100# a_n1763_n274# 0.15fF
C457 a_n1521_122# a_n1763_n274# 3.88fF
.ends

.subckt sky130_fd_pr__nfet_01v8_J3WY8C a_n4080_n100# a_n1188_122# a_282_n188# a_n978_n188#
+ a_1542_n188# a_n3918_n188# a_3432_122# a_1752_122# a_n3708_122# a_2382_n188# a_4228_n100#
+ a_n2028_122# a_n1818_n188# a_3222_n188# a_n348_122# a_n2658_n188# a_n3288_122# a_4062_n188#
+ a_72_122# a_n558_n188# a_n3498_n188# a_1122_n188# a_912_122# a_n4172_n100# a_3852_122#
+ a_n1398_n188# a_2172_122# a_n4128_122# a_n2448_122# a_492_122# a_n768_122# a_n2238_n188#
+ a_n138_n188# a_n3078_n188# a_1962_n188# a_702_n188# a_3012_122# a_1332_122# a_n1608_122#
+ a_n4382_n100# a_2802_n188# a_2592_122# a_3642_n188# a_n2868_122# VSUBS
X0 a_n4080_n100# a_n1398_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=1.24e+13p pd=1.048e+08u as=1.24e+13p ps=1.048e+08u w=1e+06u l=150000u
X1 a_n4080_n100# a_1332_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n4080_n100# a_n2868_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n4080_n100# a_2802_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n4080_n100# a_n3288_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n4080_n100# a_3222_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n4080_n100# a_72_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n4080_n100# a_n1608_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n4080_n100# a_1542_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n4080_n100# a_n138_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n4080_n100# a_282_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n4080_n100# a_n3498_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n4080_n100# a_3432_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n4080_n100# a_n1818_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n4080_n100# a_1752_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n4080_n100# a_492_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n4080_n100# a_2172_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n4080_n100# a_n3708_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n4080_n100# a_n348_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n4080_n100# a_3642_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n4080_n100# a_4062_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_n4080_n100# a_n2028_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n4080_n100# a_1962_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_n4080_n100# a_702_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_n4080_n100# a_n3918_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n4080_n100# a_n558_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n4080_n100# a_3852_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_4228_n100# a_4228_n100# a_4228_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X28 a_n4080_n100# a_n2238_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_n4080_n100# a_n768_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_n4080_n100# a_912_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n4080_n100# a_n4128_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_n4080_n100# a_n2448_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_n4080_n100# a_2382_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_n4080_n100# a_n978_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n4382_n100# a_n4382_n100# a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X36 a_n4080_n100# a_n1188_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_n4080_n100# a_1122_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n4080_n100# a_n2658_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_n4080_n100# a_2592_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_n4080_n100# a_n3078_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_n4080_n100# a_3012_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_3432_122# a_n4172_n100# 0.06fF
C1 a_1542_n188# a_n4172_n100# 0.02fF
C2 a_n4128_122# a_n4080_n100# 0.02fF
C3 a_2802_n188# a_n4172_n100# 0.02fF
C4 a_3852_122# a_n4172_n100# 0.06fF
C5 a_72_122# a_n4172_n100# 0.06fF
C6 a_n1188_122# a_n2658_n188# 0.00fF
C7 a_n138_n188# a_n1398_n188# 0.00fF
C8 a_702_n188# a_1332_122# 0.00fF
C9 a_n1608_122# a_n4080_n100# 0.02fF
C10 a_n348_122# a_n138_n188# 0.00fF
C11 a_n4172_n100# a_1332_122# 0.06fF
C12 a_2382_n188# a_2592_122# 0.00fF
C13 a_1122_n188# a_702_n188# 0.01fF
C14 a_n4172_n100# a_n2028_122# 0.06fF
C15 a_1542_n188# a_912_122# 0.00fF
C16 a_n3708_122# a_n2448_122# 0.00fF
C17 a_n3498_n188# a_n2658_n188# 0.01fF
C18 a_n1188_122# a_n4080_n100# 0.02fF
C19 a_72_122# a_912_122# 0.01fF
C20 a_3642_n188# a_3432_122# 0.00fF
C21 a_1122_n188# a_n4172_n100# 0.02fF
C22 a_282_n188# a_n768_122# 0.00fF
C23 a_n2868_122# a_n2448_122# 0.01fF
C24 a_2802_n188# a_3642_n188# 0.01fF
C25 a_n1398_n188# a_n2868_122# 0.00fF
C26 a_3852_122# a_3642_n188# 0.00fF
C27 a_n2028_122# a_n2238_n188# 0.00fF
C28 a_2382_n188# a_n4080_n100# 0.06fF
C29 a_72_122# a_n558_n188# 0.00fF
C30 a_n1398_n188# a_n1818_n188# 0.01fF
C31 a_n2448_122# a_n1818_n188# 0.00fF
C32 a_912_122# a_1332_122# 0.01fF
C33 a_n4128_122# a_n4172_n100# 0.06fF
C34 a_n3498_n188# a_n4080_n100# 0.06fF
C35 a_3222_n188# a_2382_n188# 0.01fF
C36 a_n348_122# a_n1818_n188# 0.00fF
C37 a_1122_n188# a_912_122# 0.00fF
C38 a_n558_n188# a_n2028_122# 0.00fF
C39 a_1542_n188# a_1752_122# 0.00fF
C40 a_2802_n188# a_1752_122# 0.00fF
C41 a_n4172_n100# a_n1608_122# 0.06fF
C42 a_n768_122# a_n4080_n100# 0.02fF
C43 a_72_122# a_n138_n188# 0.00fF
C44 a_n3918_n188# a_n2448_122# 0.00fF
C45 a_n3288_122# a_n2028_122# 0.00fF
C46 a_4228_n100# a_3432_122# 0.00fF
C47 a_n978_n188# a_n2448_122# 0.00fF
C48 a_n1188_122# a_n4172_n100# 0.06fF
C49 a_1962_n188# a_2592_122# 0.00fF
C50 a_n978_n188# a_n1398_n188# 0.01fF
C51 a_492_122# a_n348_122# 0.01fF
C52 a_n2238_n188# a_n1608_122# 0.00fF
C53 a_2802_n188# a_4228_n100# 0.00fF
C54 a_3432_122# a_3012_122# 0.01fF
C55 a_n138_n188# a_1332_122# 0.00fF
C56 a_3852_122# a_4228_n100# 0.01fF
C57 a_1332_122# a_1752_122# 0.01fF
C58 a_1542_n188# a_3012_122# 0.00fF
C59 a_2382_n188# a_n4172_n100# 0.02fF
C60 a_2802_n188# a_3012_122# 0.00fF
C61 a_n4128_122# a_n4382_n100# 0.00fF
C62 a_3852_122# a_3012_122# 0.01fF
C63 a_n978_n188# a_n348_122# 0.00fF
C64 a_n1188_122# a_n2238_n188# 0.00fF
C65 a_1962_n188# a_n4080_n100# 0.06fF
C66 a_1122_n188# a_n138_n188# 0.00fF
C67 a_1122_n188# a_1752_122# 0.00fF
C68 a_n4128_122# a_n3288_122# 0.01fF
C69 a_n3498_n188# a_n4172_n100# 0.02fF
C70 a_n558_n188# a_n1608_122# 0.00fF
C71 a_702_n188# a_n768_122# 0.00fF
C72 a_3222_n188# a_1962_n188# 0.00fF
C73 a_2382_n188# a_912_122# 0.00fF
C74 a_n2868_122# a_n2028_122# 0.01fF
C75 a_n1188_122# a_n558_n188# 0.00fF
C76 a_n3498_n188# a_n2238_n188# 0.00fF
C77 a_n4172_n100# a_n768_122# 0.06fF
C78 a_3642_n188# a_2382_n188# 0.00fF
C79 a_492_122# a_1542_n188# 0.00fF
C80 a_n2028_122# a_n1818_n188# 0.00fF
C81 a_492_122# a_72_122# 0.01fF
C82 a_n2238_n188# a_n768_122# 0.00fF
C83 a_n138_n188# a_n1608_122# 0.00fF
C84 a_n4128_122# a_n3708_122# 0.01fF
C85 a_1962_n188# a_702_n188# 0.00fF
C86 a_72_122# a_n978_n188# 0.00fF
C87 a_n4382_n100# a_n3498_n188# 0.00fF
C88 a_n4128_122# a_n2868_122# 0.00fF
C89 a_n1188_122# a_n138_n188# 0.00fF
C90 a_492_122# a_1332_122# 0.01fF
C91 a_1962_n188# a_n4172_n100# 0.02fF
C92 a_2172_122# a_3432_122# 0.00fF
C93 a_n3288_122# a_n3498_n188# 0.00fF
C94 a_2172_122# a_1542_n188# 0.00fF
C95 a_2172_122# a_2802_n188# 0.00fF
C96 a_2382_n188# a_1752_122# 0.00fF
C97 a_n558_n188# a_n768_122# 0.00fF
C98 a_492_122# a_1122_n188# 0.00fF
C99 a_n978_n188# a_n2028_122# 0.00fF
C100 a_n2868_122# a_n1608_122# 0.00fF
C101 a_n3078_n188# a_n2658_n188# 0.01fF
C102 a_n1398_n188# a_n2448_122# 0.00fF
C103 a_n1608_122# a_n1818_n188# 0.00fF
C104 a_2172_122# a_1332_122# 0.01fF
C105 a_1962_n188# a_912_122# 0.00fF
C106 a_2382_n188# a_3012_122# 0.00fF
C107 a_n4128_122# a_n3918_n188# 0.00fF
C108 a_n348_122# a_n1398_n188# 0.00fF
C109 a_n1188_122# a_n1818_n188# 0.00fF
C110 a_n138_n188# a_n768_122# 0.00fF
C111 a_n3078_n188# a_n4080_n100# 0.06fF
C112 a_2172_122# a_1122_n188# 0.00fF
C113 a_n3708_122# a_n3498_n188# 0.00fF
C114 a_n3498_n188# a_n2868_122# 0.00fF
C115 a_n978_n188# a_n1608_122# 0.00fF
C116 a_282_n188# a_n4080_n100# 0.06fF
C117 a_1962_n188# a_1752_122# 0.00fF
C118 a_n978_n188# a_n1188_122# 0.00fF
C119 a_n1818_n188# a_n768_122# 0.00fF
C120 a_n2658_n188# a_n4080_n100# 0.06fF
C121 a_2592_122# a_n4080_n100# 0.02fF
C122 a_72_122# a_n1398_n188# 0.00fF
C123 a_n3918_n188# a_n3498_n188# 0.01fF
C124 a_n4172_n100# a_n3078_n188# 0.02fF
C125 a_1962_n188# a_3012_122# 0.00fF
C126 a_72_122# a_n348_122# 0.01fF
C127 a_2172_122# a_2382_n188# 0.00fF
C128 a_3222_n188# a_2592_122# 0.00fF
C129 a_492_122# a_n768_122# 0.00fF
C130 a_n2448_122# a_n2028_122# 0.01fF
C131 a_n3078_n188# a_n2238_n188# 0.01fF
C132 a_n1398_n188# a_n2028_122# 0.00fF
C133 a_702_n188# a_282_n188# 0.01fF
C134 a_n978_n188# a_n768_122# 0.00fF
C135 a_282_n188# a_n4172_n100# 0.02fF
C136 a_3222_n188# a_n4080_n100# 0.06fF
C137 a_4062_n188# a_2592_122# 0.00fF
C138 a_1122_n188# a_n348_122# 0.00fF
C139 a_n4172_n100# a_n2658_n188# 0.02fF
C140 a_492_122# a_1962_n188# 0.00fF
C141 a_n4382_n100# a_n3078_n188# 0.00fF
C142 a_2592_122# a_n4172_n100# 0.06fF
C143 a_2802_n188# a_3432_122# 0.00fF
C144 a_3852_122# a_3432_122# 0.01fF
C145 a_2802_n188# a_1542_n188# 0.00fF
C146 a_n3288_122# a_n3078_n188# 0.00fF
C147 a_4062_n188# a_n4080_n100# 0.06fF
C148 a_72_122# a_1542_n188# 0.00fF
C149 a_282_n188# a_912_122# 0.00fF
C150 a_n2658_n188# a_n2238_n188# 0.01fF
C151 a_3852_122# a_2802_n188# 0.00fF
C152 a_702_n188# a_n4080_n100# 0.06fF
C153 a_n1398_n188# a_n1608_122# 0.00fF
C154 a_n2448_122# a_n1608_122# 0.01fF
C155 a_n4172_n100# a_n4080_n100# 15.77fF
C156 a_282_n188# a_n558_n188# 0.01fF
C157 a_3222_n188# a_4062_n188# 0.01fF
C158 a_1542_n188# a_1332_122# 0.00fF
C159 a_2172_122# a_1962_n188# 0.00fF
C160 a_2802_n188# a_1332_122# 0.00fF
C161 a_n348_122# a_n1608_122# 0.00fF
C162 a_n1188_122# a_n1398_n188# 0.00fF
C163 a_n1188_122# a_n2448_122# 0.00fF
C164 a_72_122# a_1332_122# 0.00fF
C165 a_n2238_n188# a_n4080_n100# 0.06fF
C166 a_3222_n188# a_n4172_n100# 0.02fF
C167 a_n4382_n100# a_n2658_n188# 0.00fF
C168 a_1122_n188# a_1542_n188# 0.01fF
C169 a_3642_n188# a_2592_122# 0.00fF
C170 a_n348_122# a_n1188_122# 0.01fF
C171 a_72_122# a_1122_n188# 0.00fF
C172 a_n3708_122# a_n3078_n188# 0.00fF
C173 a_n3288_122# a_n2658_n188# 0.00fF
C174 a_912_122# a_n4080_n100# 0.02fF
C175 a_282_n188# a_n138_n188# 0.01fF
C176 a_282_n188# a_1752_122# 0.00fF
C177 a_n2868_122# a_n3078_n188# 0.00fF
C178 a_n3498_n188# a_n2448_122# 0.00fF
C179 a_3642_n188# a_n4080_n100# 0.06fF
C180 a_n558_n188# a_n4080_n100# 0.06fF
C181 a_1122_n188# a_1332_122# 0.00fF
C182 a_4062_n188# a_n4172_n100# 0.02fF
C183 a_n4382_n100# a_n4080_n100# 0.14fF
C184 a_702_n188# a_n4172_n100# 0.02fF
C185 a_n3078_n188# a_n1818_n188# 0.00fF
C186 a_n1398_n188# a_n768_122# 0.00fF
C187 a_2592_122# a_1752_122# 0.01fF
C188 a_n3288_122# a_n4080_n100# 0.02fF
C189 a_3222_n188# a_3642_n188# 0.01fF
C190 a_n348_122# a_n768_122# 0.01fF
C191 a_n3708_122# a_n2658_n188# 0.00fF
C192 a_n4172_n100# a_n2238_n188# 0.02fF
C193 a_4228_n100# a_2592_122# 0.00fF
C194 a_n138_n188# a_n4080_n100# 0.06fF
C195 a_n4080_n100# a_1752_122# 0.02fF
C196 a_702_n188# a_912_122# 0.00fF
C197 a_n3918_n188# a_n3078_n188# 0.01fF
C198 a_n2868_122# a_n2658_n188# 0.00fF
C199 a_72_122# a_n1188_122# 0.00fF
C200 a_2382_n188# a_3432_122# 0.00fF
C201 a_2592_122# a_3012_122# 0.01fF
C202 a_3642_n188# a_4062_n188# 0.01fF
C203 a_2382_n188# a_1542_n188# 0.01fF
C204 a_912_122# a_n4172_n100# 0.06fF
C205 a_2802_n188# a_2382_n188# 0.01fF
C206 a_702_n188# a_n558_n188# 0.00fF
C207 a_3852_122# a_2382_n188# 0.00fF
C208 a_n2028_122# a_n1608_122# 0.01fF
C209 a_n2658_n188# a_n1818_n188# 0.01fF
C210 a_3222_n188# a_1752_122# 0.00fF
C211 a_4228_n100# a_n4080_n100# 0.21fF
C212 a_n3708_122# a_n4080_n100# 0.02fF
C213 a_3642_n188# a_n4172_n100# 0.02fF
C214 a_n558_n188# a_n4172_n100# 0.02fF
C215 a_3012_122# a_n4080_n100# 0.02fF
C216 a_n4382_n100# a_n4172_n100# 0.21fF
C217 a_n1188_122# a_n2028_122# 0.01fF
C218 a_492_122# a_282_n188# 0.00fF
C219 a_n2868_122# a_n4080_n100# 0.02fF
C220 a_2382_n188# a_1332_122# 0.00fF
C221 a_3222_n188# a_4228_n100# 0.00fF
C222 a_n3288_122# a_n4172_n100# 0.06fF
C223 a_n978_n188# a_282_n188# 0.00fF
C224 a_n1818_n188# a_n4080_n100# 0.06fF
C225 a_3222_n188# a_3012_122# 0.00fF
C226 a_n3918_n188# a_n2658_n188# 0.00fF
C227 a_702_n188# a_n138_n188# 0.01fF
C228 a_702_n188# a_1752_122# 0.00fF
C229 a_1122_n188# a_2382_n188# 0.00fF
C230 a_72_122# a_n768_122# 0.01fF
C231 a_n3498_n188# a_n2028_122# 0.00fF
C232 a_n3288_122# a_n2238_n188# 0.00fF
C233 a_n558_n188# a_912_122# 0.00fF
C234 a_n138_n188# a_n4172_n100# 0.02fF
C235 a_n4172_n100# a_1752_122# 0.06fF
C236 a_4062_n188# a_4228_n100# 0.00fF
C237 a_4062_n188# a_3012_122# 0.00fF
C238 a_492_122# a_n4080_n100# 0.02fF
C239 a_n3918_n188# a_n4080_n100# 0.06fF
C240 a_n2028_122# a_n768_122# 0.00fF
C241 a_1962_n188# a_3432_122# 0.00fF
C242 a_1962_n188# a_1542_n188# 0.01fF
C243 a_4228_n100# a_n4172_n100# 0.14fF
C244 a_n3708_122# a_n4172_n100# 0.06fF
C245 a_1962_n188# a_2802_n188# 0.01fF
C246 a_n1188_122# a_n1608_122# 0.01fF
C247 a_2172_122# a_2592_122# 0.01fF
C248 a_n978_n188# a_n4080_n100# 0.06fF
C249 a_n4172_n100# a_3012_122# 0.06fF
C250 a_n4128_122# a_n3498_n188# 0.00fF
C251 a_n4382_n100# a_n3288_122# 0.00fF
C252 a_n138_n188# a_912_122# 0.00fF
C253 a_912_122# a_1752_122# 0.01fF
C254 a_n2868_122# a_n4172_n100# 0.06fF
C255 a_n3708_122# a_n2238_n188# 0.00fF
C256 a_n558_n188# a_n138_n188# 0.01fF
C257 a_n4172_n100# a_n1818_n188# 0.02fF
C258 a_1962_n188# a_1332_122# 0.00fF
C259 a_2172_122# a_n4080_n100# 0.02fF
C260 a_n2868_122# a_n2238_n188# 0.00fF
C261 a_n3078_n188# a_n2448_122# 0.00fF
C262 a_1122_n188# a_1962_n188# 0.01fF
C263 a_n2238_n188# a_n1818_n188# 0.01fF
C264 a_3642_n188# a_4228_n100# 0.00fF
C265 a_492_122# a_702_n188# 0.00fF
C266 a_3222_n188# a_2172_122# 0.00fF
C267 a_n1608_122# a_n768_122# 0.01fF
C268 a_3642_n188# a_3012_122# 0.00fF
C269 a_n4382_n100# a_n3708_122# 0.00fF
C270 a_492_122# a_n4172_n100# 0.06fF
C271 a_n3918_n188# a_n4172_n100# 0.02fF
C272 a_n3708_122# a_n3288_122# 0.01fF
C273 a_n4382_n100# a_n2868_122# 0.00fF
C274 a_n1188_122# a_n768_122# 0.01fF
C275 a_n978_n188# a_n4172_n100# 0.02fF
C276 a_n558_n188# a_n1818_n188# 0.00fF
C277 a_n3288_122# a_n2868_122# 0.01fF
C278 a_2172_122# a_702_n188# 0.00fF
C279 a_n348_122# a_282_n188# 0.00fF
C280 a_n1398_n188# a_n2658_n188# 0.00fF
C281 a_n978_n188# a_n2238_n188# 0.00fF
C282 a_n2448_122# a_n2658_n188# 0.00fF
C283 a_n3288_122# a_n1818_n188# 0.00fF
C284 a_2172_122# a_n4172_n100# 0.06fF
C285 a_3012_122# a_1752_122# 0.00fF
C286 a_492_122# a_912_122# 0.01fF
C287 a_492_122# a_n558_n188# 0.00fF
C288 a_n4382_n100# a_n3918_n188# 0.01fF
C289 a_4228_n100# a_3012_122# 0.00fF
C290 a_1962_n188# a_2382_n188# 0.01fF
C291 a_n978_n188# a_n558_n188# 0.01fF
C292 a_n2448_122# a_n4080_n100# 0.02fF
C293 a_n1398_n188# a_n4080_n100# 0.06fF
C294 a_n3708_122# a_n2868_122# 0.01fF
C295 a_n3918_n188# a_n3288_122# 0.00fF
C296 a_2172_122# a_912_122# 0.00fF
C297 a_n348_122# a_n4080_n100# 0.02fF
C298 a_2172_122# a_3642_n188# 0.00fF
C299 a_492_122# a_n138_n188# 0.00fF
C300 a_492_122# a_1752_122# 0.00fF
C301 a_1542_n188# a_282_n188# 0.00fF
C302 a_n2868_122# a_n1818_n188# 0.00fF
C303 a_n3078_n188# a_n2028_122# 0.00fF
C304 a_72_122# a_282_n188# 0.00fF
C305 a_n978_n188# a_n138_n188# 0.01fF
C306 a_2592_122# a_3432_122# 0.01fF
C307 a_n3708_122# a_n3918_n188# 0.00fF
C308 a_1542_n188# a_2592_122# 0.00fF
C309 a_282_n188# a_1332_122# 0.00fF
C310 a_2802_n188# a_2592_122# 0.00fF
C311 a_3852_122# a_2592_122# 0.00fF
C312 a_2172_122# a_1752_122# 0.01fF
C313 a_n4128_122# a_n3078_n188# 0.00fF
C314 a_n3918_n188# a_n2868_122# 0.00fF
C315 a_n4172_n100# a_n2448_122# 0.06fF
C316 a_n1398_n188# a_n4172_n100# 0.02fF
C317 a_702_n188# a_n348_122# 0.00fF
C318 a_3432_122# a_n4080_n100# 0.02fF
C319 a_1122_n188# a_282_n188# 0.01fF
C320 a_1542_n188# a_n4080_n100# 0.06fF
C321 a_n2658_n188# a_n2028_122# 0.00fF
C322 a_2802_n188# a_n4080_n100# 0.06fF
C323 a_2592_122# a_1332_122# 0.00fF
C324 a_3852_122# a_n4080_n100# 0.02fF
C325 a_n348_122# a_n4172_n100# 0.06fF
C326 a_72_122# a_n4080_n100# 0.02fF
C327 a_n3078_n188# a_n1608_122# 0.00fF
C328 a_n1398_n188# a_n2238_n188# 0.01fF
C329 a_n978_n188# a_n1818_n188# 0.01fF
C330 a_n2448_122# a_n2238_n188# 0.00fF
C331 a_2172_122# a_3012_122# 0.01fF
C332 a_3222_n188# a_3432_122# 0.00fF
C333 a_1122_n188# a_2592_122# 0.00fF
C334 a_3222_n188# a_2802_n188# 0.01fF
C335 a_3222_n188# a_3852_122# 0.00fF
C336 a_1332_122# a_n4080_n100# 0.02fF
C337 a_n2028_122# a_n4080_n100# 0.02fF
C338 a_n4128_122# a_n2658_n188# 0.00fF
C339 a_n348_122# a_912_122# 0.00fF
C340 a_n558_n188# a_n1398_n188# 0.01fF
C341 a_1122_n188# a_n4080_n100# 0.06fF
C342 a_492_122# a_n978_n188# 0.00fF
C343 a_4062_n188# a_3432_122# 0.00fF
C344 a_702_n188# a_1542_n188# 0.01fF
C345 a_2802_n188# a_4062_n188# 0.00fF
C346 a_n348_122# a_n558_n188# 0.00fF
C347 a_3852_122# a_4062_n188# 0.00fF
C348 a_n3288_122# a_n2448_122# 0.01fF
C349 a_n3498_n188# a_n3078_n188# 0.01fF
C350 a_n1188_122# a_282_n188# 0.00fF
C351 a_n2658_n188# a_n1608_122# 0.00fF
C352 a_72_122# a_702_n188# 0.00fF
C353 a_n4080_n100# VSUBS 1.08fF
C354 a_n4172_n100# VSUBS 1.03fF
C355 a_4062_n188# VSUBS 0.11fF
C356 a_4228_n100# VSUBS 0.17fF
C357 a_3642_n188# VSUBS 0.10fF
C358 a_3852_122# VSUBS 0.09fF
C359 a_3222_n188# VSUBS 0.11fF
C360 a_3432_122# VSUBS 0.11fF
C361 a_2802_n188# VSUBS 0.12fF
C362 a_3012_122# VSUBS 0.11fF
C363 a_2382_n188# VSUBS 0.12fF
C364 a_2592_122# VSUBS 0.12fF
C365 a_1962_n188# VSUBS 0.12fF
C366 a_2172_122# VSUBS 0.12fF
C367 a_1542_n188# VSUBS 0.12fF
C368 a_1752_122# VSUBS 0.12fF
C369 a_1122_n188# VSUBS 0.12fF
C370 a_1332_122# VSUBS 0.12fF
C371 a_702_n188# VSUBS 0.12fF
C372 a_912_122# VSUBS 0.12fF
C373 a_282_n188# VSUBS 0.12fF
C374 a_492_122# VSUBS 0.12fF
C375 a_n138_n188# VSUBS 0.12fF
C376 a_72_122# VSUBS 0.12fF
C377 a_n558_n188# VSUBS 0.12fF
C378 a_n348_122# VSUBS 0.12fF
C379 a_n978_n188# VSUBS 0.12fF
C380 a_n768_122# VSUBS 0.12fF
C381 a_n1398_n188# VSUBS 0.12fF
C382 a_n1188_122# VSUBS 0.12fF
C383 a_n1818_n188# VSUBS 0.12fF
C384 a_n1608_122# VSUBS 0.12fF
C385 a_n2238_n188# VSUBS 0.12fF
C386 a_n2028_122# VSUBS 0.12fF
C387 a_n2658_n188# VSUBS 0.12fF
C388 a_n2448_122# VSUBS 0.12fF
C389 a_n3078_n188# VSUBS 0.12fF
C390 a_n2868_122# VSUBS 0.12fF
C391 a_n3498_n188# VSUBS 0.12fF
C392 a_n3288_122# VSUBS 0.12fF
C393 a_n3918_n188# VSUBS 0.12fF
C394 a_n3708_122# VSUBS 0.12fF
C395 a_n4382_n100# VSUBS 0.20fF
C396 a_n4128_122# VSUBS 0.13fF
.ends

.subckt latch_nmos_pair sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
C0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C2 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C5 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C6 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C7 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.02fF
C8 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.02fF
C9 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C10 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C11 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C12 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C13 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C14 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C15 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C16 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C17 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 1.18fF
C18 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C19 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C20 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C21 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.01fF
C22 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C23 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C24 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.57fF
C25 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C26 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C27 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C28 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C29 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C30 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C31 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C32 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C33 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C34 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C35 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C36 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C37 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C38 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C39 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.02fF
C40 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# -0.00fF
C41 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C42 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C43 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C44 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C45 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C46 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C47 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.02fF
C48 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C49 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C50 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C51 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C52 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C53 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C54 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C55 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C56 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C57 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C58 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C59 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C60 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C61 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.02fF
C62 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C63 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C64 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C65 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C66 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C67 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C68 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C69 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C70 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C71 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# -0.00fF
C72 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.02fF
C73 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C74 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C75 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C76 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C77 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C78 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C79 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C80 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C81 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C82 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C83 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C84 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C85 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C86 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C87 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C88 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C89 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C90 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C91 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C92 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C93 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C94 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.02fF
C95 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C96 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C97 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.02fF
C98 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.02fF
C99 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C100 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C101 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# -0.00fF
C102 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C103 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C104 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.02fF
C105 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C106 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C107 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# -0.00fF
C108 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C109 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C110 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C111 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C112 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.01fF
C113 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.02fF
C114 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.02fF
C115 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C117 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C118 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C119 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C121 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C122 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C123 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.02fF
C125 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C126 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# -0.00fF
C127 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C128 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C129 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C130 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.02fF
C131 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C132 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C133 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.02fF
C134 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C135 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C136 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C137 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C138 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C139 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C140 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C141 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C142 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C143 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C144 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C145 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# -0.00fF
C146 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.17fF
C147 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C148 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.02fF
C149 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C150 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.02fF
C151 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C152 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C153 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C154 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C155 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C156 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.31fF
C157 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C158 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C159 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C160 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C161 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C162 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C163 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C164 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C165 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C166 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C167 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C168 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C169 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C170 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C171 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C172 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C173 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C174 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C175 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C176 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C177 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C178 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C180 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C181 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.02fF
C182 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C183 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C184 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C186 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C187 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C189 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C190 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C191 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C192 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.02fF
C193 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C194 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C195 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.02fF
C196 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C197 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C201 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C202 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C203 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C204 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C206 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C207 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C208 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.02fF
C209 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C210 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C211 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C212 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C213 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.02fF
C214 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C215 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.01fF
C216 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C217 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.02fF
C218 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C219 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.02fF
C220 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C221 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C222 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C223 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C224 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# -0.00fF
C225 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C226 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C227 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C228 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C229 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C230 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C231 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C232 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C233 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C234 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C235 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.42fF
C236 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C237 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C238 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C239 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C240 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C241 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C242 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C243 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C244 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C245 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C246 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C247 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C249 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C250 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C251 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C252 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C253 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C254 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C255 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C256 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C257 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C258 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C259 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C260 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C261 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# -0.00fF
C262 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C263 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C264 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C265 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C266 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C267 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C268 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C269 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C270 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C271 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C272 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C273 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C274 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C275 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.42fF
C276 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C277 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C278 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C279 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C280 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C281 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C282 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.01fF
C283 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C284 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C285 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# -0.00fF
C286 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C287 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C288 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C289 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C290 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C291 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C292 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C293 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C294 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C295 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# -0.00fF
C296 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# -0.00fF
C297 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C298 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C299 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C300 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C301 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C302 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.02fF
C303 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# -0.00fF
C304 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C305 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C306 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C307 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C308 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C309 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C310 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C311 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C312 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C313 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C314 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C315 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C316 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C317 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C318 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C319 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C320 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C321 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C322 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C323 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C324 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C325 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C326 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C327 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C328 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.02fF
C329 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C330 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C331 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C332 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C333 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C334 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C335 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C336 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C337 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C338 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C339 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C340 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C341 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C342 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C343 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C344 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C345 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C346 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C347 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C348 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C349 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C350 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C351 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.01fF
C352 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C353 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C354 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C355 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C356 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C357 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C358 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.02fF
C359 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C360 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.01fF
C361 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C362 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.02fF
C363 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C364 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C365 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C366 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C367 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C368 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C369 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C370 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C371 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.02fF
C372 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C373 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C374 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C375 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C376 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C377 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C378 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C379 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C380 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C381 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C382 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C383 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C384 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C385 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C386 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C387 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C388 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C389 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C390 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# -0.00fF
C391 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C392 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C393 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C394 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C395 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C396 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C397 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C398 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C399 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C400 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C401 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C402 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C405 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C406 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C407 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C408 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C409 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C410 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C411 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C412 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C413 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C414 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C415 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C416 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C417 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C418 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.02fF
C419 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.02fF
C420 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C421 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C422 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C423 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# -0.00fF
C424 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C425 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C426 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C427 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C428 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.02fF
C429 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C430 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C431 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C432 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# -0.00fF
C433 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C434 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C435 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C436 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.02fF
C437 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C438 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C439 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C440 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.02fF
C441 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.01fF
C442 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C443 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C444 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C445 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C446 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C447 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C448 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C449 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C450 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C451 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# -0.00fF
C452 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C453 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.02fF
C454 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C455 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C457 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C458 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C459 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C460 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C461 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C462 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C463 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C464 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C465 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.02fF
C466 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C467 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C468 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C469 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C470 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C471 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C472 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C473 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C474 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C475 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C476 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C477 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C478 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C479 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C480 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C481 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C483 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C484 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C485 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C486 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C487 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C488 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C489 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C490 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C491 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C492 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C493 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C494 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C495 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C496 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C497 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# -0.00fF
C498 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C499 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.00fF
C500 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C501 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C502 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C503 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C504 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C505 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C506 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C507 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C508 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# -0.00fF
C509 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.30fF
C510 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C511 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C512 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C513 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C514 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C515 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C516 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C517 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C518 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C519 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.02fF
C520 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C521 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C522 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C523 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.02fF
C524 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C525 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.02fF
C526 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C527 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C528 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C529 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C530 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C531 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C532 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C533 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C534 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C535 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.00fF
C536 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# -0.00fF
C537 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C538 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C539 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C540 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C541 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C542 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C543 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C544 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.01fF
C545 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C546 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C547 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C548 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.01fF
C549 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C550 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C551 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C552 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C553 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C554 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C555 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C556 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C557 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C558 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C559 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C560 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.44fF
C561 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# -0.00fF
C563 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C564 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C565 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C566 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C567 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.02fF
C568 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.01fF
C569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C570 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C571 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C572 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C574 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C575 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C577 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C578 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C579 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C580 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C581 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C582 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.02fF
C583 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C584 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C585 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C586 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.02fF
C587 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C588 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C589 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C590 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C591 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C592 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C593 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C594 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C595 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C596 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C597 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C598 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C599 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C600 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C601 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C602 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C603 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C604 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C605 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C606 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C607 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C608 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C609 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C611 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.02fF
C612 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C613 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C614 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C615 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C616 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.02fF
C617 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C618 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C619 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C620 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C621 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.02fF
C623 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C624 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C625 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C626 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C627 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C628 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C629 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C630 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# -0.00fF
C631 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.02fF
C632 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C633 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C634 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C635 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C636 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C637 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C638 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C639 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C640 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.01fF
C642 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C643 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C644 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C645 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C646 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C647 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C649 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.02fF
C650 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C651 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C652 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C653 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C654 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C655 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C656 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C657 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C658 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C659 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# -0.00fF
C660 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C661 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C662 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C663 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C664 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C665 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C666 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C667 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 1.18fF
C668 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C669 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C670 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C671 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C672 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C673 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C674 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C675 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C676 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C677 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C678 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C679 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C680 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.02fF
C681 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C683 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C684 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C685 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C686 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C687 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C688 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C689 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C690 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C691 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C692 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C693 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C694 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C695 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C696 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C697 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C698 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C699 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C700 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C701 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 1.18fF
C702 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C703 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C704 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C705 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C706 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C707 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C708 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C709 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# -0.00fF
C710 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C711 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C712 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C713 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C714 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C715 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C716 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C717 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C718 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C719 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C720 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C721 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C722 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C724 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C725 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C726 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C727 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C728 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C729 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C730 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C731 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C732 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C733 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C734 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C735 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C736 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C737 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C738 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C739 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.02fF
C740 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.01fF
C741 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C742 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C743 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C744 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C745 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C746 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C747 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# -0.00fF
C748 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C749 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C750 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C751 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C752 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C753 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C754 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C755 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C756 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C757 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C758 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C759 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C760 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C761 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.02fF
C762 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C763 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C764 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C765 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C766 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C767 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C768 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C769 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C770 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C771 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C772 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C773 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C774 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C775 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C776 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C777 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C778 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C779 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C780 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C781 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C782 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# -0.00fF
C783 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C784 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C785 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C786 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C787 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C788 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C789 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C790 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C791 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C792 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C793 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C794 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C795 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C796 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C797 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C798 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C799 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C800 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# -0.00fF
C801 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C802 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C803 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C804 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C805 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C806 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C807 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C808 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C809 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C810 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C811 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C812 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C813 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C814 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.02fF
C815 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C816 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C817 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C818 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C819 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C820 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C821 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C822 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C823 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C824 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# -0.00fF
C825 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C826 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C827 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C828 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.02fF
C829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C830 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C831 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# -0.01fF
C832 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.02fF
C833 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C834 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C835 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C836 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C837 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C838 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C839 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C840 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C841 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C842 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C843 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.02fF
C844 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C845 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C846 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C847 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C848 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.02fF
C849 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C850 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C851 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C852 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C853 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C854 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C855 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C856 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C857 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.01fF
C858 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C859 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C860 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C861 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C862 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C863 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C864 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.02fF
C865 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# -0.00fF
C866 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C867 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C868 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C869 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C870 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C871 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C872 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C873 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C874 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C875 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C876 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C877 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C878 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# -0.00fF
C879 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C880 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C881 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C882 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C883 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C884 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C885 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C886 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C887 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C888 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C889 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.02fF
C890 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C891 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.02fF
C892 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.02fF
C893 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.02fF
C894 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C895 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.02fF
C896 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C897 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C898 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C899 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C900 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.02fF
C901 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C902 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C903 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C904 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C905 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C906 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C907 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C908 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C909 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C910 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C911 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C912 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C913 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C914 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C915 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C916 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C917 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C918 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C919 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C920 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C921 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# -0.01fF
C922 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C923 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C924 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C925 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C926 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C927 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C928 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C929 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C930 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C931 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C932 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C933 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C934 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C935 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C936 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C937 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C938 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C939 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C940 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C941 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C942 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C943 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C944 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C945 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C946 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C947 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C948 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C949 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C950 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C951 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C952 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.01fF
C953 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C954 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.01fF
C955 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.02fF
C956 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C957 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C958 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C959 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# -0.00fF
C960 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C961 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C962 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C963 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C964 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C965 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C966 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C967 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C968 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C969 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.02fF
C970 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C971 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.31fF
C972 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C973 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# -0.00fF
C974 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C975 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C976 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C977 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.01fF
C978 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C979 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C980 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C981 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C982 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C983 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.93fF
C984 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C985 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C986 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C987 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# -0.01fF
C988 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C989 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C990 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C991 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C992 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C993 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C994 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C995 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C996 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C997 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C998 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C999 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C1000 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1001 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1002 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1003 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C1004 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C1005 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1006 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1007 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1008 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1009 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1010 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.02fF
C1011 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1012 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1013 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C1014 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1015 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1016 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C1017 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1018 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1019 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1020 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1021 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.01fF
C1022 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1023 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1024 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.24fF
C1025 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C1026 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# -0.00fF
C1027 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1028 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1029 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C1030 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1031 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1032 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1033 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C1034 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1035 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.02fF
C1036 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1037 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1038 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C1039 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# -0.00fF
C1040 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1041 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1042 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C1043 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1044 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1045 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1046 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C1047 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1048 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C1049 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C1050 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.01fF
C1051 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.02fF
C1052 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1053 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1054 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1055 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1056 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C1057 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.02fF
C1058 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1060 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1061 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1062 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1063 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C1064 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1065 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1066 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C1067 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1068 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1069 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.02fF
C1070 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1072 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C1073 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C1074 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1075 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C1076 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.02fF
C1077 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C1078 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1079 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1080 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1081 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1082 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C1083 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1084 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1085 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1086 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C1087 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1088 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1089 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C1090 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C1091 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1092 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1093 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C1094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C1095 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1096 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C1097 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1098 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1099 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1100 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1101 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1102 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1103 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1104 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# -0.00fF
C1105 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1106 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1107 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1108 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C1109 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1111 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1112 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.02fF
C1113 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1114 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C1116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1117 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1118 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# -0.00fF
C1119 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.42fF
C1120 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1121 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1122 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1123 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1124 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1125 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C1126 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1127 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1128 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1130 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# -0.00fF
C1132 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1133 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1134 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1135 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.02fF
C1136 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C1137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1138 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# -0.01fF
C1139 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C1140 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1142 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1143 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1144 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1146 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C1147 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C1148 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C1149 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1150 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1151 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1152 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C1153 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1154 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1155 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1156 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1157 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1158 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.57fF
C1159 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C1160 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1161 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1162 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1163 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1164 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1165 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1166 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C1167 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1168 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1169 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1170 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C1171 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1172 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# -0.00fF
C1173 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.02fF
C1174 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1175 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1176 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C1177 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1178 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C1179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# -0.00fF
C1180 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1181 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1182 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C1183 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1184 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1185 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# -0.00fF
C1186 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1187 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1189 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C1190 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C1191 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C1192 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C1193 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1194 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1195 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1196 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.02fF
C1197 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C1200 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1201 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C1202 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1203 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1204 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1205 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C1206 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1207 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1208 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1209 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1210 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1211 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C1212 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1213 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1214 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1215 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C1216 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C1217 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.44fF
C1218 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1219 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1220 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1221 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1222 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1223 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1224 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1225 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1226 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.76fF
C1227 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1228 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1229 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1230 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1231 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1232 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1233 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1234 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1235 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1236 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1237 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1238 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# -0.00fF
C1239 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C1240 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C1241 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C1242 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1243 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1244 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.01fF
C1245 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1246 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# -0.00fF
C1247 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1248 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C1249 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1250 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1251 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1252 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C1253 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C1254 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1255 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# -0.00fF
C1256 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1257 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1258 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.93fF
C1259 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1260 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.01fF
C1261 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1262 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1263 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1264 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.02fF
C1265 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.42fF
C1266 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1267 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C1268 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# -0.00fF
C1269 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1270 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C1271 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1272 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# -0.00fF
C1273 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.93fF
C1274 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C1275 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1276 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C1277 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1278 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1279 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1280 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1281 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.02fF
C1282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1283 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1284 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1285 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1286 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1287 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1288 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1289 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1290 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1291 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1292 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1293 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1294 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1295 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C1296 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C1297 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# -0.00fF
C1298 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C1299 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1300 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C1301 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1302 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C1303 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1304 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1305 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C1306 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C1307 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1308 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C1309 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1310 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1311 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1312 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C1313 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# -0.00fF
C1314 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1315 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1316 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.02fF
C1317 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1318 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.02fF
C1319 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1320 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1321 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1322 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1323 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C1324 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.02fF
C1325 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1326 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1327 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C1328 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1329 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.02fF
C1330 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1331 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1332 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.02fF
C1333 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1334 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C1335 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.02fF
C1336 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1337 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1338 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1339 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1340 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1341 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1342 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1343 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1344 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C1345 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1346 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C1347 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.02fF
C1348 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1349 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.01fF
C1350 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1351 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1352 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1353 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1354 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.01fF
C1355 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C1356 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C1357 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1358 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1359 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1360 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1361 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1362 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1363 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1364 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C1365 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C1366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C1367 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C1368 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1369 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C1370 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C1371 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1372 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1373 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C1374 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1375 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1376 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C1377 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C1378 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1379 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C1380 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1381 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1382 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1383 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C1384 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# -0.00fF
C1385 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# -0.01fF
C1386 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1387 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.02fF
C1388 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1389 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C1390 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1391 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.02fF
C1392 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1393 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C1394 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1395 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1396 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1397 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1398 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1399 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C1400 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1401 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.01fF
C1402 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1403 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C1405 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C1406 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1407 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1408 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1409 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# -0.00fF
C1410 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.93fF
C1411 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1412 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1413 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1414 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1415 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.02fF
C1416 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1417 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1418 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1419 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1420 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1421 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C1422 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C1423 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C1424 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1425 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C1426 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1427 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# -0.00fF
C1428 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1429 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1430 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1431 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1432 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C1433 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1434 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1435 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1436 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1437 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1438 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1439 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C1440 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1441 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C1442 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1443 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C1444 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.01fF
C1446 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1447 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1448 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1449 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C1450 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1451 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1452 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1453 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C1454 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1455 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C1457 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1458 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1459 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.02fF
C1460 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1461 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1462 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1463 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1464 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1465 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C1466 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.02fF
C1467 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1468 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.93fF
C1469 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C1470 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1471 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1472 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.01fF
C1473 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# -0.00fF
C1474 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1475 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1476 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1477 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1478 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1479 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# -0.00fF
C1480 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1481 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1483 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1484 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1485 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1486 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C1487 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1488 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1489 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C1490 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1491 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1492 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1493 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1494 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1495 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1496 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1497 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1498 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.02fF
C1499 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1500 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1501 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1502 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1503 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1504 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1505 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1506 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1507 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1508 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.02fF
C1509 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C1510 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1511 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.02fF
C1512 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C1513 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1514 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1515 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C1516 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1517 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.02fF
C1518 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1519 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.57fF
C1520 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C1521 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1522 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1523 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1524 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C1525 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1526 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C1527 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C1528 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C1529 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1530 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.01fF
C1531 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1532 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1533 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.22fF
C1534 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1535 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1536 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1537 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C1538 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C1540 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1541 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1542 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1543 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1544 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.02fF
C1545 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1546 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C1547 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1548 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# -0.00fF
C1549 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1550 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1551 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C1552 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C1553 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.02fF
C1554 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C1555 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1556 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1557 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1558 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1559 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C1560 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# VSUBS 1.08fF
C1561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# VSUBS 1.03fF
C1562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# VSUBS 0.11fF
C1563 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# VSUBS 0.17fF
C1564 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# VSUBS 0.10fF
C1565 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# VSUBS 0.09fF
C1566 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# VSUBS 0.11fF
C1567 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# VSUBS 0.11fF
C1568 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# VSUBS 0.12fF
C1569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# VSUBS 0.11fF
C1570 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# VSUBS 0.12fF
C1571 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# VSUBS 0.12fF
C1572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# VSUBS 0.12fF
C1573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# VSUBS 0.12fF
C1574 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# VSUBS 0.12fF
C1575 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# VSUBS 0.12fF
C1576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# VSUBS 0.12fF
C1577 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# VSUBS 0.12fF
C1578 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# VSUBS 0.12fF
C1579 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# VSUBS 0.12fF
C1580 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# VSUBS 0.12fF
C1581 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# VSUBS 0.12fF
C1582 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# VSUBS 0.12fF
C1583 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# VSUBS 0.12fF
C1584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# VSUBS 0.12fF
C1585 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# VSUBS 0.12fF
C1586 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# VSUBS 0.12fF
C1587 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# VSUBS 0.12fF
C1588 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# VSUBS 0.12fF
C1589 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# VSUBS 0.12fF
C1590 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# VSUBS 0.12fF
C1591 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# VSUBS 0.12fF
C1592 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# VSUBS 0.12fF
C1593 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# VSUBS 0.12fF
C1594 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# VSUBS 0.12fF
C1595 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# VSUBS 0.12fF
C1596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# VSUBS 0.12fF
C1597 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# VSUBS 0.12fF
C1598 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# VSUBS 0.12fF
C1599 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# VSUBS 0.12fF
C1600 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# VSUBS 0.12fF
C1601 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# VSUBS 0.12fF
C1602 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# VSUBS 0.20fF
C1603 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# VSUBS 0.13fF
C1604 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# VSUBS 1.08fF
C1605 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# VSUBS 1.03fF
C1606 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# VSUBS 0.11fF
C1607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# VSUBS 0.17fF
C1608 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# VSUBS 0.10fF
C1609 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# VSUBS 0.09fF
C1610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# VSUBS 0.11fF
C1611 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# VSUBS 0.11fF
C1612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# VSUBS 0.12fF
C1613 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# VSUBS 0.11fF
C1614 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# VSUBS 0.12fF
C1615 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# VSUBS 0.12fF
C1616 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# VSUBS 0.12fF
C1617 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# VSUBS 0.12fF
C1618 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# VSUBS 0.12fF
C1619 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# VSUBS 0.12fF
C1620 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# VSUBS 0.12fF
C1621 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# VSUBS 0.12fF
C1622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# VSUBS 0.12fF
C1623 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# VSUBS 0.12fF
C1624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# VSUBS 0.12fF
C1625 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# VSUBS 0.12fF
C1626 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# VSUBS 0.12fF
C1627 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# VSUBS 0.12fF
C1628 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# VSUBS 0.12fF
C1629 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# VSUBS 0.12fF
C1630 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# VSUBS 0.12fF
C1631 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# VSUBS 0.12fF
C1632 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# VSUBS 0.12fF
C1633 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# VSUBS 0.12fF
C1634 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# VSUBS 0.12fF
C1635 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# VSUBS 0.12fF
C1636 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# VSUBS 0.12fF
C1637 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# VSUBS 0.12fF
C1638 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# VSUBS 0.12fF
C1639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# VSUBS 0.12fF
C1640 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# VSUBS 0.12fF
C1641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# VSUBS 0.12fF
C1642 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# VSUBS 0.12fF
C1643 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# VSUBS 0.12fF
C1644 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# VSUBS 0.12fF
C1645 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# VSUBS 0.12fF
C1646 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# VSUBS 0.20fF
C1647 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# VSUBS 0.13fF
C1648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# VSUBS 1.08fF
C1649 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# VSUBS 1.03fF
C1650 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# VSUBS 0.11fF
C1651 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# VSUBS 0.17fF
C1652 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# VSUBS 0.10fF
C1653 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# VSUBS 0.09fF
C1654 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# VSUBS 0.11fF
C1655 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# VSUBS 0.11fF
C1656 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# VSUBS 0.12fF
C1657 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# VSUBS 0.11fF
C1658 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# VSUBS 0.12fF
C1659 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# VSUBS 0.12fF
C1660 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# VSUBS 0.12fF
C1661 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# VSUBS 0.12fF
C1662 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# VSUBS 0.12fF
C1663 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# VSUBS 0.12fF
C1664 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# VSUBS 0.12fF
C1665 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# VSUBS 0.12fF
C1666 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# VSUBS 0.12fF
C1667 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# VSUBS 0.12fF
C1668 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# VSUBS 0.12fF
C1669 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# VSUBS 0.12fF
C1670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# VSUBS 0.12fF
C1671 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# VSUBS 0.12fF
C1672 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# VSUBS 0.12fF
C1673 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# VSUBS 0.12fF
C1674 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# VSUBS 0.12fF
C1675 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# VSUBS 0.12fF
C1676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# VSUBS 0.12fF
C1677 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# VSUBS 0.12fF
C1678 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# VSUBS 0.12fF
C1679 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# VSUBS 0.12fF
C1680 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# VSUBS 0.12fF
C1681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# VSUBS 0.12fF
C1682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# VSUBS 0.12fF
C1683 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# VSUBS 0.12fF
C1684 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# VSUBS 0.12fF
C1685 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# VSUBS 0.12fF
C1686 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# VSUBS 0.12fF
C1687 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# VSUBS 0.12fF
C1688 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# VSUBS 0.12fF
C1689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# VSUBS 0.12fF
C1690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# VSUBS 0.20fF
C1691 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# VSUBS 0.13fF
C1692 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# VSUBS 1.08fF
C1693 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# VSUBS 1.03fF
C1694 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# VSUBS 0.11fF
C1695 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# VSUBS 0.17fF
C1696 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# VSUBS 0.10fF
C1697 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# VSUBS 0.09fF
C1698 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# VSUBS 0.11fF
C1699 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# VSUBS 0.11fF
C1700 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# VSUBS 0.12fF
C1701 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# VSUBS 0.11fF
C1702 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# VSUBS 0.12fF
C1703 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# VSUBS 0.12fF
C1704 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# VSUBS 0.12fF
C1705 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# VSUBS 0.12fF
C1706 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# VSUBS 0.12fF
C1707 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# VSUBS 0.12fF
C1708 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# VSUBS 0.12fF
C1709 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# VSUBS 0.12fF
C1710 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# VSUBS 0.12fF
C1711 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# VSUBS 0.12fF
C1712 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# VSUBS 0.12fF
C1713 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# VSUBS 0.12fF
C1714 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# VSUBS 0.12fF
C1715 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# VSUBS 0.12fF
C1716 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# VSUBS 0.12fF
C1717 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# VSUBS 0.12fF
C1718 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# VSUBS 0.12fF
C1719 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# VSUBS 0.12fF
C1720 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# VSUBS 0.12fF
C1721 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# VSUBS 0.12fF
C1722 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# VSUBS 0.12fF
C1723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# VSUBS 0.12fF
C1724 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# VSUBS 0.12fF
C1725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# VSUBS 0.12fF
C1726 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# VSUBS 0.12fF
C1727 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# VSUBS 0.12fF
C1728 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# VSUBS 0.12fF
C1729 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# VSUBS 0.12fF
C1730 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# VSUBS 0.12fF
C1731 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# VSUBS 0.12fF
C1732 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# VSUBS 0.12fF
C1733 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# VSUBS 0.12fF
C1734 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# VSUBS 0.20fF
C1735 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# VSUBS 0.13fF
.ends

.subckt input_diff_pair sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_4 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_5 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_6 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_7 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
C0 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# -0.00fF
C2 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C4 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C5 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C6 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.01fF
C7 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# -0.00fF
C8 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C9 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C10 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C11 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C12 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# 0.01fF
C13 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C14 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C15 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.02fF
C16 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C17 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.02fF
C18 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C19 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C20 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C21 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C22 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.31fF
C23 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.02fF
C24 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.02fF
C25 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C26 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C27 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C28 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C29 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C30 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C31 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C32 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C33 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C34 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C35 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C36 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C37 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C38 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C39 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C40 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C41 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C42 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C43 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C44 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# -0.00fF
C45 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C46 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C47 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C48 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.02fF
C49 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.01fF
C50 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# -0.00fF
C51 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C52 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C53 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# 0.02fF
C54 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C55 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C56 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C57 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C58 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.01fF
C59 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C60 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C61 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.02fF
C62 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C63 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C64 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C65 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C66 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C67 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C68 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C69 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.02fF
C70 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C71 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C72 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C73 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C74 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C75 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C76 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C77 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.93fF
C78 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C79 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.42fF
C80 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C81 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C82 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C83 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C84 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# -0.00fF
C85 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C86 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C87 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C88 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C89 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C90 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C91 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C92 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C93 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C94 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C95 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C96 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C97 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C98 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C99 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C100 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C101 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C102 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C103 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.00fF
C104 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C105 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C106 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C107 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C108 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C109 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C110 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C111 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C112 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C113 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C114 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C115 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C116 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C117 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C118 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C119 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C120 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C121 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.02fF
C122 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C123 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C124 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C125 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C126 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C127 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C128 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C129 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C130 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C132 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C133 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C134 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C135 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C136 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C138 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C139 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C140 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C142 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C143 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C144 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C145 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C146 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C147 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C148 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# -0.00fF
C149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C151 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C152 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C153 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C154 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C155 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C156 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C157 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C158 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.01fF
C159 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C161 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C162 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C163 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C164 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C165 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C166 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C167 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C168 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C169 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.01fF
C170 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C171 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C172 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C173 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C174 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C175 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C176 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C177 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C178 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.57fF
C179 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C180 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C181 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C182 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C183 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.93fF
C184 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.00fF
C185 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C186 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C187 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C189 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C190 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C191 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C192 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C193 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C194 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C195 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C196 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C197 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C198 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C199 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C200 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.00fF
C201 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C202 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C203 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C206 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C207 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C208 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C209 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C210 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C211 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C212 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C213 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C214 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C215 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C216 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# -0.00fF
C217 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C218 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C219 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C220 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# -0.00fF
C221 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C222 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C223 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.00fF
C224 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C225 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C226 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C227 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C228 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C229 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.02fF
C230 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C231 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.02fF
C232 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.01fF
C233 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.01fF
C234 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C235 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C236 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C237 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C238 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C239 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C240 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C241 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C242 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C243 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C244 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.02fF
C245 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C246 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.42fF
C247 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C248 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C249 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C250 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C251 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C252 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C253 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C254 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C255 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C256 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C257 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C258 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C259 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C260 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C261 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C262 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C263 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C264 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C265 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C266 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C267 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C268 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C269 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C270 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C271 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C272 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C273 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C274 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C275 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C276 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C277 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C278 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C279 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C280 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C281 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C282 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C283 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C284 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C285 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C286 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C287 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C288 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C289 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.42fF
C290 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C291 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.02fF
C292 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.00fF
C293 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C294 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C295 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.57fF
C296 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C297 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C298 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C299 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C300 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.02fF
C301 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C302 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C303 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.02fF
C304 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C305 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C306 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C307 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C308 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.01fF
C309 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C310 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# -0.00fF
C311 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.01fF
C312 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C313 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C314 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C315 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C316 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C317 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C318 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C319 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C320 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C321 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C322 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C323 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C324 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.02fF
C325 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C326 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C327 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C328 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C329 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.00fF
C330 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C331 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.02fF
C332 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.00fF
C333 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C334 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C335 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C336 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C337 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C338 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C339 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.00fF
C340 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C341 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.01fF
C342 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C343 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.93fF
C344 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C345 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.27fF
C346 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C347 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C348 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C349 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C350 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C351 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C352 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C353 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C354 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C355 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C356 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C357 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C358 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C359 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C360 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C361 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C362 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C363 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C364 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C365 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.02fF
C366 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C367 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.02fF
C368 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C369 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C370 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.01fF
C371 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C372 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.02fF
C373 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C374 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C375 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C376 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C378 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C379 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C380 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C381 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C382 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C383 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C384 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C385 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.01fF
C386 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.02fF
C387 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.02fF
C388 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C389 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C390 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C391 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C392 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C393 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C394 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C395 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C396 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.93fF
C397 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C398 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C399 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C400 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C401 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C402 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C403 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# 0.00fF
C405 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.01fF
C406 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C407 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C408 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C409 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C410 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C411 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.01fF
C412 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C413 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C414 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C415 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C416 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C417 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C418 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C419 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C420 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C421 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C422 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C423 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C424 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C425 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C426 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C427 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# -0.00fF
C428 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C429 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# -0.00fF
C430 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C431 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C432 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.01fF
C433 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.01fF
C434 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C435 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C436 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C437 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C438 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C439 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C440 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C441 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C442 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C443 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.02fF
C444 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C445 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.17fF
C446 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C447 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C448 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C449 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C450 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C451 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C452 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# -0.00fF
C453 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C454 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C455 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C456 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C457 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C458 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C459 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C460 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.27fF
C461 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C462 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C463 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C464 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.02fF
C465 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C466 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C467 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C468 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C469 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C470 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.02fF
C471 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C472 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C473 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.02fF
C474 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C475 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C476 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C477 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C478 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C479 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C480 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C481 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C482 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C483 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C484 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C485 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C486 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.30fF
C487 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C488 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# -0.00fF
C489 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C490 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C491 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C492 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C493 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C494 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C495 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C496 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C497 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C498 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C499 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C500 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.02fF
C501 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C502 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C503 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C504 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C505 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C506 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C507 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C508 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C509 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C510 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C511 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C512 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.02fF
C513 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C514 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C515 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.02fF
C516 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C517 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C518 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C519 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C520 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C521 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C522 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C523 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C524 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C525 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C526 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C527 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C528 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C529 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C530 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C531 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C532 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C533 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C534 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.00fF
C535 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# -0.00fF
C536 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C537 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C538 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C539 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# -0.00fF
C540 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C541 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.02fF
C542 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C543 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C544 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C545 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C546 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C547 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C548 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C549 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 1.18fF
C550 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C551 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C552 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C553 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C554 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C555 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# -0.00fF
C556 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C557 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C558 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C559 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.27fF
C560 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C563 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C564 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C565 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.02fF
C566 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C567 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.01fF
C568 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C569 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.02fF
C570 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C571 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C572 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C573 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C574 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C575 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C576 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C577 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C578 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C579 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C580 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C581 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C582 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C583 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C585 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.00fF
C586 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C587 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C588 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C589 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C590 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C591 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C592 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C593 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C594 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C595 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C596 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C597 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C598 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# -0.00fF
C599 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C600 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.02fF
C601 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C602 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C603 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C604 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.02fF
C605 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C606 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C608 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# -0.00fF
C609 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# -0.00fF
C610 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C611 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.02fF
C612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.02fF
C613 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.02fF
C614 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C615 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C616 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C617 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C618 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.01fF
C619 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C620 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C621 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C622 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C623 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C625 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C626 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C627 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C628 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C629 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C630 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# -0.00fF
C631 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.01fF
C632 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C633 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C634 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C635 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C636 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C637 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C638 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C640 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C641 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C642 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# -0.00fF
C643 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C644 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C645 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.02fF
C646 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C647 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.00fF
C648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C649 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C650 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# -0.00fF
C651 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C652 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C653 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C654 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C655 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C656 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C657 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C658 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C659 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C660 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C661 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C662 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C663 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.02fF
C664 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C665 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# -0.00fF
C666 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# -0.00fF
C667 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C668 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C669 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C670 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C671 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C672 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C673 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C674 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C675 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C676 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C677 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C678 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C679 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C680 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# -0.00fF
C681 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C682 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C683 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C684 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C685 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C686 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C687 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.01fF
C688 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.02fF
C689 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C690 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C691 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C692 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.02fF
C693 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C694 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C695 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C696 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C697 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C698 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C699 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C700 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C701 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.02fF
C702 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C703 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C704 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C705 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C706 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C707 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C708 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C709 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.01fF
C710 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C711 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C712 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C713 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C714 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C715 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.01fF
C716 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.93fF
C717 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C718 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# -0.00fF
C719 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C720 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C721 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C722 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C723 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.93fF
C724 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C726 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C727 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C728 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C729 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C730 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C731 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C732 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C733 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.27fF
C734 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C735 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C736 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C737 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C738 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.02fF
C739 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C740 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.01fF
C741 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C742 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.01fF
C743 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C744 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C745 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C746 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C747 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C748 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C749 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C750 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C751 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C752 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.00fF
C753 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C754 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C755 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C756 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# 0.01fF
C757 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C758 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C759 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C760 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.02fF
C761 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C762 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.01fF
C763 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# -0.01fF
C764 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C765 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C766 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C767 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C768 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C769 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C770 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C771 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.01fF
C772 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C773 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C774 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C775 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C776 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C777 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C778 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C779 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C780 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C781 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C782 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C783 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.02fF
C784 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C785 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.02fF
C786 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# -0.00fF
C787 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C788 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C789 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C790 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C791 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C792 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# -0.00fF
C793 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C794 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C795 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C796 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C797 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C798 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C799 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C800 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C801 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C802 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C803 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C804 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C805 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C806 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C807 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C808 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C809 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C810 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C811 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C812 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.01fF
C813 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C814 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C815 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C816 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.02fF
C817 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C818 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C819 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C820 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C821 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.00fF
C822 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C823 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C824 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C825 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C826 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C827 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C828 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C829 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C830 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C831 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C832 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C833 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C834 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C835 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C836 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C838 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# 0.00fF
C839 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# -0.00fF
C840 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C841 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C842 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C843 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C844 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C845 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.02fF
C846 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C847 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C848 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C849 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# -0.00fF
C850 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C851 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C852 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C853 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C854 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C855 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# -0.00fF
C856 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C857 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# -0.00fF
C858 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C859 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C860 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C861 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.02fF
C862 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C863 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C864 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C865 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.01fF
C866 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C867 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C868 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C869 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C870 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C871 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C872 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C873 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# -0.00fF
C874 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C875 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C876 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C877 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C878 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C879 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C880 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C881 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.02fF
C882 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C883 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C884 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C885 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C886 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C887 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C888 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C889 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C890 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.42fF
C891 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C892 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C893 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C894 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C896 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C897 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C898 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# -0.00fF
C899 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.02fF
C900 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C901 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C902 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C903 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C904 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C905 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C906 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C907 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C908 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C909 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.02fF
C910 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C911 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C912 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C913 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C914 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.01fF
C915 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C916 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C917 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C918 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C919 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# -0.00fF
C920 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.01fF
C921 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.02fF
C922 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C923 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.22fF
C924 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C925 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C926 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C927 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C928 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C929 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.02fF
C930 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C931 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C932 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C933 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C934 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C935 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C936 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C937 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C938 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C939 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C940 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C941 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C942 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C943 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C944 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C945 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C946 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C947 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C948 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C949 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C950 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C951 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C952 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.00fF
C953 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C954 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C955 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C956 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C957 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C958 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# -0.00fF
C959 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C960 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C961 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C962 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C963 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.02fF
C964 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.01fF
C965 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C966 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C967 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C968 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C969 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.01fF
C970 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C971 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C972 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C973 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C974 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C975 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 1.18fF
C976 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C977 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C978 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C979 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C980 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C981 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C982 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C983 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C984 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.02fF
C985 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C986 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C987 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.02fF
C988 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C989 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C990 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C991 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C992 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C993 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C994 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C995 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.02fF
C996 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C997 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# -0.01fF
C998 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C999 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C1000 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C1001 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.00fF
C1002 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1003 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C1004 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C1006 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C1007 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C1008 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.02fF
C1009 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C1010 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# 0.00fF
C1011 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1012 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1013 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C1014 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1015 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C1016 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C1017 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1018 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1019 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1020 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C1021 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C1022 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.01fF
C1023 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# -0.00fF
C1024 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1025 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1026 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C1027 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# -0.00fF
C1028 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1029 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1030 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1031 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1032 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C1033 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1034 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C1035 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1036 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C1037 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1038 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.02fF
C1039 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1040 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C1041 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1042 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C1043 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1044 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C1045 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1046 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1047 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1048 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C1049 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1050 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1051 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1052 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C1053 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C1054 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C1055 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1056 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C1057 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C1058 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C1059 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1060 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1061 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C1062 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1063 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.02fF
C1064 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C1065 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.02fF
C1066 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C1067 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C1068 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1069 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C1070 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C1071 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1072 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1073 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# -0.00fF
C1074 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C1075 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1076 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1077 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C1078 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.31fF
C1079 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1080 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C1081 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1082 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# -0.00fF
C1083 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# -0.01fF
C1084 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C1085 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C1086 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C1087 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1088 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.01fF
C1089 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1090 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1091 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1092 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1093 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1094 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1095 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C1096 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C1097 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1098 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1099 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1100 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C1101 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1102 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1103 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C1104 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C1105 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C1106 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.02fF
C1107 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1108 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C1109 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.02fF
C1110 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C1111 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1112 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1113 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.02fF
C1114 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1115 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C1116 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1117 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1118 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1119 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C1120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C1121 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1122 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C1123 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C1124 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1125 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1126 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C1127 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1128 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C1129 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.00fF
C1130 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C1131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C1132 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.44fF
C1133 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1134 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C1135 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1136 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1137 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1138 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1139 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1140 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1141 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1142 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1143 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C1144 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C1145 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C1146 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1147 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# -0.00fF
C1148 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# -0.00fF
C1149 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.01fF
C1150 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C1151 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1152 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1153 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1154 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.01fF
C1155 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C1156 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1157 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1158 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C1159 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C1160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1161 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C1162 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1163 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1164 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1165 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1166 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C1167 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1168 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C1169 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C1170 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C1171 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1172 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1173 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C1174 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1175 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C1176 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1177 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1178 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C1179 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C1180 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.02fF
C1181 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C1182 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1183 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.02fF
C1184 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.01fF
C1185 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# -0.00fF
C1186 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1187 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C1188 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.02fF
C1189 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1190 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1191 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1192 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C1193 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1194 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C1195 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1196 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.01fF
C1197 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C1198 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1199 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1200 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# -0.00fF
C1201 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1202 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.02fF
C1203 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C1204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C1205 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C1206 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1207 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C1208 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C1209 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1210 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1211 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C1212 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# -0.00fF
C1213 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1214 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1215 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C1216 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C1217 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1218 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C1219 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1220 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1221 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C1222 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1223 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.01fF
C1224 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1225 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1226 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C1227 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C1228 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1229 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1230 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C1231 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C1232 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1233 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.01fF
C1234 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.02fF
C1235 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C1236 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1237 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1238 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# -0.00fF
C1239 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1240 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1241 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C1242 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1243 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C1244 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1245 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C1246 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1247 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.02fF
C1248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1249 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# -0.00fF
C1250 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C1251 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1252 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C1253 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1254 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C1255 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C1256 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C1257 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C1258 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1259 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C1260 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C1261 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C1262 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1263 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1264 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1265 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1266 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1267 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C1268 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C1269 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1270 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1271 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.01fF
C1272 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# -0.00fF
C1273 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C1274 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1275 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.01fF
C1276 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1277 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# -0.00fF
C1278 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# -0.00fF
C1279 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1280 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.02fF
C1281 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C1282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C1283 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C1284 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1285 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.02fF
C1286 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C1287 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C1288 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1289 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C1290 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1291 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1292 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1293 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.01fF
C1294 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1295 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1296 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C1297 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C1298 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C1299 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1300 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.02fF
C1301 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# -0.00fF
C1302 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1303 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1304 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1305 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1306 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C1307 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.00fF
C1308 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C1309 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1310 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.02fF
C1311 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1312 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C1313 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.01fF
C1314 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.02fF
C1315 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C1316 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1317 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C1318 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C1319 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C1320 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C1321 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C1322 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1323 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1324 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1325 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C1326 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1327 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# -0.00fF
C1328 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1329 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C1330 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1331 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C1332 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1333 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C1334 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1335 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# -0.00fF
C1336 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# -0.00fF
C1337 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1338 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.02fF
C1339 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1340 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C1341 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1342 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C1343 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.01fF
C1344 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1345 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1346 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1347 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C1348 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1349 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1350 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C1351 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1352 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# -0.00fF
C1353 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1354 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1355 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C1356 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C1357 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1358 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C1359 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# -0.00fF
C1360 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1361 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.02fF
C1362 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1363 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1364 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C1365 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C1366 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1367 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1368 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1369 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C1370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1371 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C1372 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1373 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.01fF
C1374 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C1375 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1376 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1377 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C1378 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.01fF
C1379 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.02fF
C1380 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C1381 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C1382 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C1383 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1384 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C1385 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C1386 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1387 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C1388 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C1389 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1390 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1391 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.01fF
C1392 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1393 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1394 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.01fF
C1395 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C1396 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C1397 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1398 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1399 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C1400 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C1401 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# -0.00fF
C1402 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C1403 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1404 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1405 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C1406 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C1407 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1408 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1409 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1410 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C1411 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.00fF
C1412 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C1413 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C1414 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1415 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1416 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C1417 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C1418 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1419 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C1420 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1421 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1422 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C1423 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C1424 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C1425 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1426 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1427 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1428 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1429 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1430 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1431 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1432 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C1433 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C1434 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1435 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1436 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C1437 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.00fF
C1438 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C1439 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1440 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C1441 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1442 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1443 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# -0.01fF
C1444 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# -0.00fF
C1445 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C1446 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# -0.00fF
C1447 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# -0.00fF
C1448 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C1449 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1450 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1451 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1452 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1453 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.42fF
C1454 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1455 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1456 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1457 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C1458 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C1459 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C1460 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C1462 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C1463 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1464 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C1465 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.01fF
C1466 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# -0.00fF
C1467 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C1468 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.01fF
C1469 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1470 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C1471 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C1472 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1473 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1474 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1475 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1476 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.02fF
C1477 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1478 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.02fF
C1479 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1480 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1481 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C1482 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1483 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1484 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C1485 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1486 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.02fF
C1487 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1488 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C1489 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1490 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# 0.00fF
C1491 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# -0.01fF
C1492 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1493 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.02fF
C1494 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.57fF
C1495 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1496 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1497 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.02fF
C1498 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C1499 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C1500 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1501 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C1502 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1503 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1504 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.01fF
C1505 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C1506 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1507 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C1508 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C1509 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1510 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C1511 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.02fF
C1512 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C1513 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1514 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1515 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1516 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.01fF
C1517 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1518 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1519 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1520 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1521 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C1522 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C1523 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C1524 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.02fF
C1525 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1526 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C1527 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1528 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1529 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1530 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C1531 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.01fF
C1532 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C1533 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C1534 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C1535 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1536 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1537 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C1538 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1540 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1541 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1542 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C1543 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1544 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C1545 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.00fF
C1546 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1547 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C1548 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1549 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C1550 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.02fF
C1551 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1552 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C1553 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1554 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1555 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1556 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C1557 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C1558 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C1559 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1560 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.02fF
C1561 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1562 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1563 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.02fF
C1564 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1565 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1566 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C1567 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C1568 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.02fF
C1569 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1570 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1571 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.02fF
C1572 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C1573 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C1574 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1575 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C1576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C1577 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C1578 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C1579 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C1580 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C1581 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.02fF
C1582 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C1583 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C1584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C1585 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1586 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1587 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1588 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C1589 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C1590 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C1591 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C1592 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C1593 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C1594 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1595 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1596 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1597 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1598 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1599 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1600 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.27fF
C1601 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1602 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# -0.01fF
C1603 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C1604 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C1605 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C1606 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C1608 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1609 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C1610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1611 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1612 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C1613 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.01fF
C1614 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1615 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1616 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1617 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1618 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# -0.00fF
C1619 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C1620 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1621 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C1622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1623 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1624 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C1625 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1626 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# -0.00fF
C1627 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C1628 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C1629 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C1630 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1631 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C1632 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1633 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# -0.00fF
C1634 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C1635 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C1636 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C1637 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C1638 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1639 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1640 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C1641 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C1642 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1643 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.19fF
C1644 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1645 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.02fF
C1646 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C1647 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1648 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1649 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1650 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C1651 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.00fF
C1652 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C1653 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1654 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C1655 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C1656 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1657 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1658 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C1659 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1660 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1661 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C1662 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.02fF
C1663 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1664 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1665 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1666 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C1667 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# -0.00fF
C1668 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1669 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1670 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C1671 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C1672 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1673 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1674 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C1675 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C1676 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1677 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C1678 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# 0.00fF
C1679 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C1680 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C1682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C1683 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1684 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1685 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.27fF
C1686 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1687 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# 0.00fF
C1688 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1689 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C1690 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.01fF
C1691 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C1692 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1693 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1694 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1695 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C1696 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C1697 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.02fF
C1698 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1699 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1700 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C1701 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# -0.00fF
C1702 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1703 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.02fF
C1704 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1705 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C1706 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.01fF
C1707 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1708 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1709 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1710 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1711 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C1712 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1713 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1714 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C1715 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C1716 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1717 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1718 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1719 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1720 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1721 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1722 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1723 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1724 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1725 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C1726 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C1727 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1728 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1729 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1730 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.01fF
C1731 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1732 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.02fF
C1733 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C1734 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C1735 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1736 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C1737 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1738 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1739 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C1740 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1741 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# -0.00fF
C1742 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1743 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.02fF
C1744 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1745 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1746 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1747 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C1748 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1749 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1750 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1751 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1752 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C1753 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1754 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1755 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1756 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.01fF
C1757 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1758 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1759 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C1760 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1761 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1762 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.02fF
C1763 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1764 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1765 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1766 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C1767 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1768 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1769 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.00fF
C1770 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C1771 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1772 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C1773 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1774 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1775 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C1776 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.44fF
C1777 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.02fF
C1778 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.31fF
C1779 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C1780 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C1781 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# -0.00fF
C1782 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1783 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C1784 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1785 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C1786 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C1787 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1788 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# -0.01fF
C1789 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# -0.00fF
C1790 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1791 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1792 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.02fF
C1793 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C1794 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1795 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1796 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1797 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.01fF
C1798 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# -0.00fF
C1799 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C1800 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C1801 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C1802 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1803 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1804 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C1805 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.01fF
C1806 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1807 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C1808 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1809 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1810 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C1811 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C1812 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1813 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C1814 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1815 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1816 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1817 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C1818 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C1819 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C1820 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C1821 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1822 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C1823 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.02fF
C1824 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1825 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1826 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1827 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1828 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C1829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C1830 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1831 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1832 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C1833 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C1834 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1835 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.01fF
C1836 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C1837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1838 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C1839 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1840 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1841 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# -0.00fF
C1842 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1843 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C1844 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1845 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1846 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1847 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.00fF
C1848 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.01fF
C1849 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C1850 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1851 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C1852 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1853 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1854 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1855 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C1856 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C1857 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.01fF
C1858 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1859 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1860 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1861 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1862 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1863 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.01fF
C1864 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C1865 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C1866 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1867 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C1868 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C1869 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C1870 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C1871 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1872 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1873 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.00fF
C1874 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C1875 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C1876 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# -0.00fF
C1877 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C1878 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C1879 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1880 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1881 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# -0.00fF
C1882 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C1883 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1884 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1885 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1886 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1887 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C1888 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.57fF
C1889 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C1890 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1891 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C1892 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.01fF
C1893 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C1894 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C1895 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C1896 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C1897 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1898 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C1899 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1900 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1901 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1902 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# -0.00fF
C1903 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C1904 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C1906 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C1907 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1908 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1909 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C1910 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1911 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C1912 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C1913 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1914 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1915 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C1916 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1917 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1918 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1919 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1920 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1921 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C1922 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C1923 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C1924 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1925 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C1926 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1927 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.01fF
C1928 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1929 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C1930 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C1931 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C1932 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1933 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1934 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C1935 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C1936 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1937 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# 0.00fF
C1938 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C1939 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1940 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C1941 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C1942 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.02fF
C1943 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1944 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1945 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1946 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C1947 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C1948 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1949 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1950 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1951 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1952 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1953 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1954 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1955 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C1956 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1957 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C1958 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# -0.00fF
C1959 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1960 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.02fF
C1961 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1962 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1963 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.27fF
C1964 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# -0.00fF
C1965 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# 0.00fF
C1966 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1967 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.44fF
C1968 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C1969 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1970 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C1971 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.02fF
C1972 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1973 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1974 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.00fF
C1975 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C1976 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C1977 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C1978 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C1979 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.02fF
C1980 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C1981 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C1982 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1983 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1984 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1985 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1986 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1987 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1988 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1989 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1990 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1991 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1992 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C1993 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1994 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1995 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1996 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C1997 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# 0.01fF
C1998 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1999 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C2000 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.01fF
C2001 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.02fF
C2002 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C2003 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C2004 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2005 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C2006 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2007 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2008 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C2009 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C2010 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C2011 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2012 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.02fF
C2013 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2014 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C2015 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2016 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2017 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C2018 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.01fF
C2019 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C2020 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# -0.00fF
C2021 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2022 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2023 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C2024 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C2025 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C2026 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C2027 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2028 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2029 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2030 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C2031 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C2032 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2033 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2034 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C2035 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C2036 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2037 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# 0.00fF
C2038 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C2039 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2040 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C2041 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.01fF
C2042 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C2043 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C2044 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C2045 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C2046 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2047 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2048 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C2049 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2050 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2051 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2052 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2053 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2054 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2055 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C2056 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2057 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2058 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.02fF
C2059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.02fF
C2060 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2061 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C2062 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C2063 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.42fF
C2064 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2065 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2066 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2067 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C2068 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C2069 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2070 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C2071 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# 0.01fF
C2072 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C2073 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C2074 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C2075 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C2076 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C2077 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2078 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2079 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2080 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.27fF
C2081 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2082 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.02fF
C2083 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C2084 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2085 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.01fF
C2086 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2087 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2088 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C2089 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.02fF
C2090 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2091 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C2092 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.02fF
C2093 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C2094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2095 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2096 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2097 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2098 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2099 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2100 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2101 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# -0.00fF
C2102 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2103 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C2104 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2105 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C2106 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C2107 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2108 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2109 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C2110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2111 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.01fF
C2112 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C2113 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2114 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C2116 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# -0.00fF
C2117 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C2118 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.02fF
C2119 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C2120 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C2121 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2122 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2123 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.02fF
C2124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C2125 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C2126 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2127 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C2128 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2129 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C2130 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2131 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C2132 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# -0.00fF
C2133 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# -0.01fF
C2134 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C2135 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C2136 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C2137 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2138 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# -0.00fF
C2139 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2140 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.02fF
C2141 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C2142 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C2143 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C2144 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C2145 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.00fF
C2146 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2147 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C2148 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2149 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2150 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C2151 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.02fF
C2152 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# -0.00fF
C2153 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2154 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2155 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.01fF
C2156 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C2157 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C2158 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C2159 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C2160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2161 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2162 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2163 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2164 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2165 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.02fF
C2166 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C2167 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2168 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C2169 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C2170 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.02fF
C2171 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C2172 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C2173 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2174 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2175 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2176 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C2177 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2178 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C2179 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C2180 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2181 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2182 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C2183 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C2184 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2185 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C2186 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2187 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C2188 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C2189 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2190 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C2191 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C2192 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C2193 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2195 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2196 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C2197 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2198 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2199 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.00fF
C2200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C2201 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C2202 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.02fF
C2203 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C2204 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2205 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.01fF
C2206 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C2207 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2208 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2209 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C2210 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.01fF
C2211 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C2212 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2213 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C2214 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2215 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C2216 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C2217 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C2218 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2219 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.02fF
C2220 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.01fF
C2221 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C2222 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.00fF
C2223 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2224 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2225 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.02fF
C2226 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C2227 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2228 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2229 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C2230 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2231 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2232 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2233 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.01fF
C2234 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2235 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2236 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2237 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2238 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.02fF
C2239 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C2240 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C2241 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.01fF
C2242 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C2243 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C2244 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.01fF
C2245 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C2246 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C2247 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C2248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2249 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2250 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.01fF
C2251 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.93fF
C2252 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C2253 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C2254 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C2255 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C2256 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2257 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C2258 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2259 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C2260 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2261 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2262 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.02fF
C2263 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2264 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C2265 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2266 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.02fF
C2267 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C2268 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C2269 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C2270 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C2271 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2272 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C2273 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C2274 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2275 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2276 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C2277 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C2278 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2279 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C2280 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2281 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C2282 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C2283 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2284 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C2285 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2286 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2287 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2288 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2289 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C2290 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2291 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C2292 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2293 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2294 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2295 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C2296 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C2297 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C2298 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# -0.00fF
C2299 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# -0.00fF
C2300 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2301 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C2302 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# -0.00fF
C2303 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C2304 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C2305 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2306 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2307 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C2308 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C2309 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2310 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C2311 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.02fF
C2312 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C2313 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.02fF
C2314 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2315 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C2316 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C2317 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C2318 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C2319 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C2320 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C2321 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C2322 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2323 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.02fF
C2324 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C2325 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2326 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C2327 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C2328 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2329 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C2330 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2331 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# -0.00fF
C2332 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2333 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2334 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2335 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C2336 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C2337 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C2338 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C2339 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C2340 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2341 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.02fF
C2342 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.02fF
C2343 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2344 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# 0.00fF
C2345 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2346 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2347 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.02fF
C2348 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C2349 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C2350 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# -0.00fF
C2351 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# 0.00fF
C2352 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.02fF
C2353 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C2354 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C2355 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C2356 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2357 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C2358 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2359 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2360 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C2361 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2362 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2363 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C2364 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C2365 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# -0.00fF
C2366 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C2367 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2368 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2369 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C2371 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C2372 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2373 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2374 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C2375 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2376 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2377 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2378 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# -0.00fF
C2379 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C2380 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2381 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C2382 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2383 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C2384 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C2385 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C2386 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# -0.00fF
C2387 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2388 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C2389 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2390 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C2391 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2392 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2393 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C2394 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C2395 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2396 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2397 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2398 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2399 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2400 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C2401 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C2402 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C2403 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C2404 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2405 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C2406 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.02fF
C2407 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C2408 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2409 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C2410 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2411 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C2412 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C2413 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# -0.00fF
C2414 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C2415 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# -0.00fF
C2416 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# -0.00fF
C2417 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C2418 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2419 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.02fF
C2420 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C2421 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C2422 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# -0.00fF
C2423 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2424 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C2425 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2426 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2427 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C2428 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2429 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.01fF
C2430 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C2431 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C2432 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C2433 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2434 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C2435 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.02fF
C2436 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.01fF
C2437 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C2438 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2439 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C2440 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.02fF
C2441 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C2442 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2443 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2444 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C2445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C2446 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C2447 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C2448 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C2449 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C2450 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C2451 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.02fF
C2452 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C2453 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.02fF
C2454 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2455 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 1.18fF
C2456 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C2457 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2458 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2459 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2460 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C2461 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C2462 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C2463 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2464 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C2465 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2466 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2467 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C2468 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C2469 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C2470 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C2471 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2472 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C2473 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2474 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C2475 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2476 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2477 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C2478 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2479 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2480 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2481 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.00fF
C2482 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C2483 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C2484 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2485 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C2486 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C2487 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C2488 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C2489 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# -0.00fF
C2490 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2491 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2492 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2493 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C2494 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C2495 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C2496 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# -0.00fF
C2497 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C2498 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C2499 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2500 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C2501 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2502 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2503 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2504 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C2505 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.01fF
C2506 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C2507 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2508 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C2509 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2510 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2511 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C2512 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2513 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C2514 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2515 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2516 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C2517 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C2518 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C2519 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C2520 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C2521 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2522 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C2523 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C2524 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2525 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2526 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2527 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2528 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C2529 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2530 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2531 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C2532 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2533 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C2534 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2535 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2536 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C2537 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2538 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C2540 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C2541 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# -0.00fF
C2542 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# -0.00fF
C2543 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2544 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C2545 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2546 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C2547 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C2548 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2549 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C2550 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C2551 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2552 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2553 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C2554 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2555 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2556 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C2557 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.00fF
C2558 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.02fF
C2559 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C2560 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2561 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2562 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.31fF
C2563 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.44fF
C2564 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2565 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2566 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C2567 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C2568 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C2569 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2570 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C2571 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.02fF
C2572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2573 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2574 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C2575 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.02fF
C2576 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2577 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2578 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.31fF
C2579 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.02fF
C2580 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C2581 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C2582 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C2583 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.00fF
C2585 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.02fF
C2586 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C2587 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.02fF
C2588 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.01fF
C2589 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2590 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C2591 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# -0.00fF
C2592 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C2593 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2594 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2595 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C2597 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2598 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2599 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C2600 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C2601 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C2602 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2603 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C2604 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.02fF
C2605 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C2606 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C2607 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C2608 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2609 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2610 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2611 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C2612 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 1.18fF
C2613 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.02fF
C2614 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2615 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C2616 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2617 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C2618 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2619 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2620 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C2621 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C2622 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2623 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.02fF
C2624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# -0.00fF
C2625 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C2626 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2627 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C2628 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2629 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C2630 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C2631 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# -0.00fF
C2632 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C2633 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C2634 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C2635 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C2636 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C2637 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C2638 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C2640 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C2641 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2642 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C2643 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2644 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2645 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C2646 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2647 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.02fF
C2648 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2649 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.48fF
C2650 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C2651 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2652 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C2653 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.01fF
C2654 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C2655 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2656 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2657 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C2658 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.01fF
C2659 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2660 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C2661 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C2662 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C2663 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C2664 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.00fF
C2665 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C2666 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2667 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2668 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2669 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C2670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C2671 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C2672 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2673 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2674 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2675 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C2676 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2677 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C2678 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C2679 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2680 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C2681 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.00fF
C2682 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C2683 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2684 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2685 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.01fF
C2686 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2687 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2688 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# 0.00fF
C2689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2690 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2691 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2692 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2693 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2694 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# -0.00fF
C2695 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C2696 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C2697 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C2698 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2699 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C2700 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C2701 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C2702 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C2703 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C2704 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C2705 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.01fF
C2706 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2707 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C2708 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2709 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2710 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.02fF
C2711 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C2712 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.01fF
C2713 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2714 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C2715 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# 0.02fF
C2716 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C2717 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2718 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2719 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C2720 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# -0.00fF
C2721 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C2722 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2724 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2725 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C2726 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2727 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2728 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C2729 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2730 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2731 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C2732 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C2733 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C2734 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C2735 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2736 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2737 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2738 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C2739 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2740 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C2741 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C2742 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2743 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2744 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C2745 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C2746 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2747 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.02fF
C2748 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C2749 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C2750 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2751 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2752 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2753 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.02fF
C2754 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# -0.00fF
C2755 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2756 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2757 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C2758 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2759 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# -0.01fF
C2760 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2761 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C2762 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C2763 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2764 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.02fF
C2765 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C2766 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2767 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C2768 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2769 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C2770 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C2771 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2772 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C2773 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C2774 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2775 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C2776 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C2777 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C2778 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C2779 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C2780 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C2781 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2782 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2783 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C2784 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2785 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.02fF
C2786 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2787 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.02fF
C2788 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C2789 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C2790 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2791 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2792 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2793 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2794 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2795 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2796 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C2797 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2798 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2799 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C2800 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C2801 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C2802 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.93fF
C2803 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 1.18fF
C2804 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2805 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C2806 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.02fF
C2807 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2808 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2809 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C2810 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2811 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C2812 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# 0.02fF
C2813 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C2814 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C2815 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2816 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2817 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2818 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C2819 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2820 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# -0.00fF
C2821 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2822 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2823 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C2824 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C2825 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2826 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2827 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2828 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C2829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2830 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.01fF
C2831 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C2832 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C2833 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2834 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C2835 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2836 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C2837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C2838 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C2839 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C2840 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2841 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C2842 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C2843 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C2844 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2845 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C2846 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C2847 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2848 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2849 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C2850 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C2851 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.00fF
C2852 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C2853 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C2854 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C2855 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2856 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C2857 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C2858 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2859 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C2860 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2861 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C2862 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# -0.00fF
C2863 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C2864 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C2865 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2866 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# -0.01fF
C2867 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C2868 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C2869 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C2870 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C2871 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C2872 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2873 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2874 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C2875 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C2876 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2877 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C2878 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C2879 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C2880 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.01fF
C2881 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2882 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C2883 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.02fF
C2884 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.01fF
C2885 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C2886 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.00fF
C2887 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C2888 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C2889 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C2890 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C2891 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2892 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# -0.00fF
C2893 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.93fF
C2894 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2895 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.01fF
C2896 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2897 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2898 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C2899 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2900 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C2901 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2902 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2903 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C2904 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2905 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2906 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2907 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C2908 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C2909 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# -0.00fF
C2910 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2911 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C2912 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C2913 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C2914 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C2915 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C2916 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C2917 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# -0.00fF
C2918 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C2919 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2920 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.02fF
C2921 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C2922 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C2923 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C2924 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C2925 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2926 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C2927 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C2928 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C2929 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# -0.00fF
C2930 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C2931 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C2932 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2933 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C2934 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C2935 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2936 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2937 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C2938 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2939 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C2940 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# -0.00fF
C2941 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C2942 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.02fF
C2943 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C2944 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C2945 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C2946 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C2947 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.02fF
C2948 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2949 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2950 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C2951 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2952 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.02fF
C2953 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C2954 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C2955 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C2956 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2957 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2958 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2959 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2960 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2961 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C2962 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2963 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C2964 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C2965 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.01fF
C2966 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2967 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2968 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2969 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2970 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C2971 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# -0.00fF
C2972 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C2973 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C2974 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C2975 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2976 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.01fF
C2977 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C2978 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2979 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2980 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2981 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2982 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2983 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C2984 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C2985 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2986 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2987 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.01fF
C2988 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2989 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2990 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2991 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C2992 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2993 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C2994 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C2995 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 1.18fF
C2996 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2997 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2998 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C2999 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# -0.00fF
C3000 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3001 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.01fF
C3002 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C3003 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# -0.00fF
C3004 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.01fF
C3006 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3007 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.02fF
C3008 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# -0.00fF
C3009 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.27fF
C3010 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# 0.00fF
C3011 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# 0.00fF
C3012 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.02fF
C3013 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3014 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3015 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C3016 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3017 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C3018 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3019 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C3020 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 1.18fF
C3021 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3022 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C3023 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C3024 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3025 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C3026 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.01fF
C3027 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# -0.00fF
C3028 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.02fF
C3029 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3030 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C3031 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C3032 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C3033 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3034 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3035 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3036 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3037 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# -0.00fF
C3038 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3039 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.02fF
C3040 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.01fF
C3041 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C3042 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# -0.00fF
C3043 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C3044 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# -0.00fF
C3045 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3046 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C3047 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C3048 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C3049 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3050 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C3051 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3052 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3053 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# -0.00fF
C3054 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3055 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.19fF
C3056 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C3057 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C3058 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.93fF
C3059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C3060 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C3061 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C3062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C3063 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C3064 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3065 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C3066 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C3067 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C3068 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3069 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C3070 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C3071 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C3072 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.02fF
C3073 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.02fF
C3074 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C3075 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3076 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3077 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C3078 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3079 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3080 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3081 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C3082 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C3083 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3084 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3085 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C3086 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3087 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.01fF
C3088 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C3089 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C3090 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C3091 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C3092 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3093 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3094 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3095 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C3096 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3097 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C3098 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C3099 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.01fF
C3100 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C3101 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C3102 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C3103 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C3104 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C3105 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# -0.00fF
C3106 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C3107 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3108 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C3109 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3110 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3111 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C3112 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# -0.00fF
C3113 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3114 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C3115 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# -0.00fF
C3116 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3117 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C3118 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.01fF
C3119 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C3120 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3121 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C3122 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C3123 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C3124 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C3125 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C3126 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3127 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.01fF
C3128 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C3130 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3131 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3132 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3133 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3134 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3135 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3136 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3137 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3138 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3139 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C3140 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C3141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C3142 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C3143 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3144 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.27fF
C3145 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C3146 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C3147 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.01fF
C3148 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3149 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C3150 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.00fF
C3151 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# -0.00fF
C3152 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C3153 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3154 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3155 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3156 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3157 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C3158 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C3159 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C3160 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.02fF
C3161 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C3162 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3163 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C3164 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C3165 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3166 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3167 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3168 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3169 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3170 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3171 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C3172 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C3173 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3174 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C3175 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C3176 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3177 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.02fF
C3178 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3179 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3180 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3181 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# -0.00fF
C3182 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3183 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3184 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.00fF
C3185 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C3186 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3187 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C3188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3189 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.02fF
C3190 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3191 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3192 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# -0.00fF
C3193 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3194 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3195 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C3196 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3197 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C3198 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3199 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3200 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.01fF
C3201 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C3202 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C3203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3205 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3206 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.01fF
C3207 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3208 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C3209 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3210 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3211 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C3212 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3213 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.01fF
C3214 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C3215 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C3216 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.02fF
C3217 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C3218 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C3219 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# 0.00fF
C3220 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C3221 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.00fF
C3222 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C3223 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3224 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C3225 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3226 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C3227 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C3228 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C3229 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C3230 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C3231 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C3232 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C3233 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C3235 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3236 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C3237 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C3238 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C3239 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3240 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3241 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C3242 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C3243 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.00fF
C3244 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3245 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.02fF
C3246 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3247 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C3248 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3249 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C3250 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3251 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3252 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3253 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3254 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C3255 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.02fF
C3256 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C3257 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3258 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C3259 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# -0.00fF
C3260 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3261 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C3262 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C3263 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C3264 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C3265 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C3266 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C3267 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3268 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# 0.00fF
C3269 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C3270 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3271 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3272 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3273 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3274 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3275 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3276 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3277 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3278 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C3279 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C3280 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C3281 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C3282 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C3283 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3284 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3285 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C3286 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C3287 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3288 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3289 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3290 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3291 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3292 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3293 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3294 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C3295 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3296 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3297 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.02fF
C3298 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3299 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3300 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3301 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C3302 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C3303 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C3304 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C3305 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3306 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C3307 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3308 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C3309 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.02fF
C3310 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.02fF
C3311 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3312 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C3313 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# -0.00fF
C3314 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.01fF
C3315 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3316 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3317 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3318 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3319 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C3320 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C3321 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C3322 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3323 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3324 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.57fF
C3325 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3326 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C3327 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.02fF
C3328 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C3329 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C3330 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C3331 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C3332 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C3333 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C3334 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3335 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C3336 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C3337 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C3338 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C3339 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C3340 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3341 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C3342 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.01fF
C3343 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# 0.00fF
C3344 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3345 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3346 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C3347 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.02fF
C3348 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3349 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3350 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C3351 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C3352 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# -0.00fF
C3353 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C3354 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C3355 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C3356 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C3357 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C3358 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3359 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C3360 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C3361 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3362 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C3363 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C3364 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3365 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C3366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C3367 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3368 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C3369 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C3370 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3371 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C3372 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.02fF
C3373 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3374 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# -0.00fF
C3375 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# -0.00fF
C3376 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C3377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# -0.00fF
C3378 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3379 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C3380 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.02fF
C3381 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3382 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C3383 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3384 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C3385 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.00fF
C3386 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C3387 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3388 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.44fF
C3389 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3390 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C3391 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3392 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C3393 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C3394 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# -0.00fF
C3395 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3396 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C3397 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C3398 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C3399 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C3400 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3401 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C3402 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C3403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.02fF
C3404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C3405 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.02fF
C3406 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C3407 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3408 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.01fF
C3409 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C3410 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3411 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3412 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3413 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C3414 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3415 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3416 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.02fF
C3417 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C3418 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C3419 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C3420 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.02fF
C3421 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.02fF
C3422 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3423 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3424 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.22fF
C3425 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C3426 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3427 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C3428 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3429 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.01fF
C3430 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3431 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C3432 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C3433 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# -0.00fF
C3434 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3435 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3436 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C3437 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3438 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3439 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3440 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C3441 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# -0.01fF
C3442 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.01fF
C3443 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C3444 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C3445 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3446 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3447 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3448 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.02fF
C3449 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.01fF
C3450 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3451 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.00fF
C3452 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C3453 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# -0.00fF
C3454 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3455 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.02fF
C3456 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3457 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C3458 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3459 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C3460 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C3462 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.01fF
C3463 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C3464 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3465 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C3466 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# -0.00fF
C3467 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3468 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3469 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3470 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# -0.00fF
C3471 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# -0.00fF
C3472 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3473 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3474 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C3475 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3476 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C3477 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.00fF
C3478 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3479 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3480 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C3481 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# -0.00fF
C3482 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C3483 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.01fF
C3484 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C3485 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C3486 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3487 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3488 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3489 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3490 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C3491 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C3492 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3493 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3494 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3495 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C3496 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3497 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C3498 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C3499 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3500 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C3501 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C3502 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C3503 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3504 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.01fF
C3505 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C3506 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.00fF
C3507 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# -0.00fF
C3508 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C3509 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3510 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C3511 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C3512 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.00fF
C3513 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C3514 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3515 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C3516 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C3517 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C3518 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3519 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3520 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C3521 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C3522 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3523 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C3524 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3525 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3526 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.02fF
C3527 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3528 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3529 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.02fF
C3530 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3531 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3532 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3533 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3534 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.31fF
C3535 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3536 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3537 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3538 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C3539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C3540 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.02fF
C3541 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3542 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.02fF
C3543 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C3544 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3545 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C3546 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.02fF
C3547 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# -0.00fF
C3548 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C3549 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C3550 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.02fF
C3551 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C3552 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C3553 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3554 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# -0.00fF
C3555 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.02fF
C3556 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C3557 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C3558 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.01fF
C3559 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C3560 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C3561 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C3562 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3563 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C3564 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3565 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C3566 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.02fF
C3567 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.27fF
C3568 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C3570 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C3571 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C3573 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3574 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3575 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.02fF
C3576 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.02fF
C3577 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# -0.00fF
C3578 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3579 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.01fF
C3580 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C3581 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3582 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3583 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C3584 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3585 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3586 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3587 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C3588 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C3589 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C3590 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C3591 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3592 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3593 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C3594 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3595 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3596 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C3597 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3598 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C3599 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3600 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C3601 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C3602 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C3603 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C3604 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.02fF
C3605 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C3606 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.02fF
C3608 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C3609 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C3611 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C3612 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C3613 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.01fF
C3614 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3615 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C3616 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C3617 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C3618 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C3619 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C3620 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C3621 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C3622 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3623 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.02fF
C3624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3625 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3626 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C3627 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3628 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C3629 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C3630 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3631 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# -0.01fF
C3632 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3633 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C3634 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C3635 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C3636 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C3637 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3638 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# -0.00fF
C3639 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# -0.00fF
C3640 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C3641 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3642 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C3643 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3644 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3645 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C3646 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C3647 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3648 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3649 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3650 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C3651 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C3652 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# -0.00fF
C3653 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.27fF
C3654 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3655 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C3656 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3657 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.01fF
C3658 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C3659 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C3660 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3661 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.02fF
C3662 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3663 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3664 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C3665 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# -0.00fF
C3666 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C3667 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.02fF
C3668 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# 0.00fF
C3669 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# 0.00fF
C3670 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3671 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3672 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C3673 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.02fF
C3674 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3675 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.02fF
C3676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C3677 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C3678 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C3679 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3680 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.57fF
C3681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C3682 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C3683 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C3684 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.02fF
C3685 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C3686 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C3687 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3688 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C3689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C3690 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C3691 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C3692 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.01fF
C3693 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C3694 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.00fF
C3695 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C3696 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C3697 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C3698 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C3699 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3700 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C3701 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3702 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C3703 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C3704 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C3705 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C3706 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.01fF
C3707 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3708 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3709 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C3710 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3711 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C3712 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3713 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.02fF
C3714 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# -0.00fF
C3715 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.42fF
C3716 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# -0.00fF
C3717 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C3718 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3719 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C3720 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C3721 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.02fF
C3722 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# -0.00fF
C3723 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# -0.00fF
C3724 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.01fF
C3725 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# -0.00fF
C3726 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C3727 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3728 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.01fF
C3729 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# -0.00fF
C3730 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.02fF
C3731 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C3732 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.44fF
C3733 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3734 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3735 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C3736 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C3737 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# -0.00fF
C3738 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.01fF
C3739 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C3740 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.01fF
C3741 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3742 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3743 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C3744 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3745 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3746 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C3747 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C3748 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C3749 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3750 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3751 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C3752 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3753 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3754 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3755 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3756 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.22fF
C3757 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3758 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3759 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3760 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3761 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C3762 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C3763 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C3764 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C3765 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C3766 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.01fF
C3767 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3768 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C3769 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.01fF
C3770 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3771 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3772 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C3773 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C3774 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C3775 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C3776 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C3777 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C3778 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3779 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3780 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.01fF
C3781 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# -0.00fF
C3782 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.01fF
C3783 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C3784 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C3785 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C3786 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.01fF
C3787 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C3788 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C3789 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C3790 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C3791 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C3792 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# -0.00fF
C3793 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.02fF
C3794 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3795 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C3796 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C3797 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# -0.00fF
C3798 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C3799 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C3800 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3801 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C3802 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# -0.00fF
C3803 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C3804 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3805 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C3806 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3807 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C3808 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3809 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.02fF
C3810 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3811 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3812 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3813 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3814 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.01fF
C3815 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C3816 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3817 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.01fF
C3818 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3819 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C3820 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C3821 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C3822 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3823 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# -0.00fF
C3824 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C3825 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3826 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3827 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3828 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C3829 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C3830 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3831 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3832 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3833 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.48fF
C3834 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3835 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3836 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3837 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C3838 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C3839 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C3840 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3841 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C3842 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3843 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C3844 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3845 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.02fF
C3846 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3847 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.02fF
C3848 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C3849 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C3850 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3851 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C3852 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C3853 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3854 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C3855 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C3856 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.01fF
C3857 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C3858 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.02fF
C3859 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C3860 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C3861 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3862 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3863 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C3864 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.01fF
C3865 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3866 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C3867 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C3868 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# -0.00fF
C3869 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3870 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C3871 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C3872 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C3873 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.27fF
C3874 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C3875 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C3876 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C3877 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C3878 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3879 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# -0.00fF
C3880 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C3881 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3882 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.01fF
C3883 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3884 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C3885 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3886 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C3887 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C3888 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C3889 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C3890 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C3891 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C3892 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C3893 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C3894 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C3895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C3896 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.02fF
C3897 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3898 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3899 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C3900 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C3901 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3902 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C3903 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C3904 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# -0.00fF
C3905 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3906 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C3907 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3908 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# 0.01fF
C3909 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C3910 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3911 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3912 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.02fF
C3913 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3914 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3915 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.01fF
C3916 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C3917 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3918 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C3919 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.78fF
C3920 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C3921 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3922 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3923 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C3924 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.01fF
C3925 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.02fF
C3926 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# -0.00fF
C3927 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.02fF
C3928 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C3929 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.02fF
C3930 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C3931 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# -0.00fF
C3932 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3933 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3934 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3935 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C3936 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3937 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3938 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C3939 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C3940 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.02fF
C3941 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C3942 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# -0.00fF
C3943 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.02fF
C3944 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3945 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C3946 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3947 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3948 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C3949 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3950 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3951 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3952 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.02fF
C3953 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C3954 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.02fF
C3955 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C3956 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C3957 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C3958 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C3959 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3960 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C3961 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.02fF
C3962 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.01fF
C3963 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C3964 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.19fF
C3965 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3966 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3967 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# -0.00fF
C3968 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# -0.00fF
C3969 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3970 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C3971 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3972 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C3973 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C3974 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C3975 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C3976 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C3977 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3978 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3979 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3980 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C3981 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C3982 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C3983 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.02fF
C3984 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C3985 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C3986 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C3987 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.02fF
C3988 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3989 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.02fF
C3990 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3991 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3992 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3993 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C3994 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3995 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C3996 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C3997 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3998 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3999 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4000 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4001 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4002 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4003 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.01fF
C4004 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C4005 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4006 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4007 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4008 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C4009 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4010 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.02fF
C4011 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C4012 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C4013 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4014 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.01fF
C4015 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4016 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4017 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4018 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.01fF
C4019 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.00fF
C4020 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4021 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4022 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C4023 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C4024 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4025 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C4026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.02fF
C4027 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.02fF
C4028 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4029 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4030 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4031 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C4032 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C4033 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4034 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# -0.00fF
C4035 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4036 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C4037 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4038 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# 0.01fF
C4039 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C4040 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C4041 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4042 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# -0.00fF
C4043 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.42fF
C4044 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C4045 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.01fF
C4046 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C4047 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4048 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4049 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C4050 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C4051 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C4052 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# -0.00fF
C4053 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# -0.00fF
C4054 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4055 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4056 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# -0.00fF
C4057 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4058 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C4060 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C4061 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4062 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C4063 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4064 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4065 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4066 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C4067 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4068 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C4069 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# -0.00fF
C4070 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C4071 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C4072 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4073 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4074 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4075 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C4076 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4077 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4078 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C4079 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.02fF
C4080 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# -0.00fF
C4081 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C4082 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C4083 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.01fF
C4084 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4085 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C4086 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4087 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4088 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C4089 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.02fF
C4090 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4091 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C4092 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C4093 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C4094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C4095 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C4096 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4097 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C4098 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4099 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C4100 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C4101 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C4102 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C4103 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4104 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C4105 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C4106 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4107 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C4108 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4109 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C4110 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.01fF
C4111 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.01fF
C4112 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4113 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# -0.00fF
C4114 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4115 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# -0.00fF
C4116 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4117 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C4118 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4119 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.42fF
C4120 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C4121 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C4122 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4123 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C4124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C4125 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C4126 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.01fF
C4127 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C4128 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.01fF
C4129 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4130 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C4131 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.01fF
C4132 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4133 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C4134 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4135 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C4136 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4137 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C4138 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C4139 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4140 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C4141 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C4142 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4143 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.02fF
C4144 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4145 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.01fF
C4146 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# -0.00fF
C4147 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C4148 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C4149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C4150 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C4151 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.93fF
C4152 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4153 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C4154 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# -0.00fF
C4155 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C4156 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C4157 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.00fF
C4158 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C4159 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.02fF
C4160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4161 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.02fF
C4162 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C4163 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C4164 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4165 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4166 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.02fF
C4167 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.00fF
C4168 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C4169 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4170 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C4171 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C4172 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C4173 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# -0.00fF
C4174 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C4175 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C4176 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C4177 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# -0.00fF
C4178 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# -0.00fF
C4179 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C4180 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4181 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4182 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C4183 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4184 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4186 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C4187 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C4188 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C4189 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4190 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4191 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C4192 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C4193 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C4194 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C4195 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C4196 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C4197 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C4198 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4200 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C4201 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4202 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C4203 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4204 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4205 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C4206 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C4207 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4208 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C4209 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C4210 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.00fF
C4211 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C4212 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C4213 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.48fF
C4214 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C4215 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4216 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4217 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.00fF
C4218 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C4219 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C4220 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4221 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C4222 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4223 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4224 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# -0.00fF
C4225 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# -0.00fF
C4226 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C4227 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4228 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4229 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4230 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4231 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4232 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4233 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C4234 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C4235 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4236 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C4237 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C4238 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C4239 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C4240 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C4241 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4242 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4243 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.02fF
C4244 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C4245 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C4246 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C4247 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C4248 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C4249 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C4250 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4251 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C4252 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# -0.00fF
C4253 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4254 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4255 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4256 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4257 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4258 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.02fF
C4259 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# 0.00fF
C4260 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4261 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.00fF
C4262 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.01fF
C4263 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C4264 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.01fF
C4265 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4266 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C4267 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4268 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.02fF
C4269 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C4270 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C4271 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4272 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C4273 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4274 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.01fF
C4275 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4276 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4277 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C4278 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C4279 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4280 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4281 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# -0.00fF
C4283 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C4284 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C4285 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.01fF
C4286 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C4287 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C4288 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C4289 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4290 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4291 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C4292 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.01fF
C4293 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C4294 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.01fF
C4295 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C4296 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4297 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4298 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4299 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C4300 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4301 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4302 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.02fF
C4303 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.93fF
C4304 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4305 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4306 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4307 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4308 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# -0.00fF
C4309 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4310 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C4311 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C4312 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# -0.00fF
C4313 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C4314 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C4315 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C4316 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C4317 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C4318 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4319 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C4320 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C4321 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C4322 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# 0.00fF
C4323 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C4324 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# -0.00fF
C4325 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4326 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C4327 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C4328 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C4329 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4330 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4331 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4332 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4333 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4334 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4335 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4336 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4337 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4338 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# -0.00fF
C4339 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C4340 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# 0.00fF
C4341 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C4342 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C4343 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C4344 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C4345 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4346 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4347 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4348 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# 0.00fF
C4349 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C4350 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C4351 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C4352 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C4353 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4354 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4355 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C4356 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4357 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4358 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.02fF
C4359 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C4360 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C4361 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C4362 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C4363 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C4364 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C4365 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C4367 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C4368 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4369 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C4370 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4371 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C4372 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C4373 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4374 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4375 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# -0.01fF
C4376 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C4377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4378 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C4379 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C4380 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C4381 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C4382 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4383 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C4384 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C4385 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C4386 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4387 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# -0.00fF
C4388 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# 0.00fF
C4389 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C4390 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C4391 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# -0.00fF
C4392 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# -0.00fF
C4393 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C4394 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4395 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C4396 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C4397 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.02fF
C4398 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.02fF
C4399 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C4400 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4401 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4402 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C4404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C4405 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C4406 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C4407 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.02fF
C4408 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C4409 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# -0.00fF
C4410 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C4411 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C4412 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C4413 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C4414 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C4415 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.02fF
C4416 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C4417 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# 0.01fF
C4418 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.02fF
C4419 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C4420 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4421 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4422 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C4423 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C4424 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.02fF
C4425 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# -0.00fF
C4426 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C4427 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.01fF
C4428 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4429 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4430 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4431 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C4432 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4433 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C4434 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4435 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C4436 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C4437 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4438 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C4439 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.01fF
C4440 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C4441 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C4442 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C4443 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# 0.01fF
C4444 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C4445 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# -0.00fF
C4446 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C4447 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C4448 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4449 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C4450 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.00fF
C4451 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4452 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.01fF
C4453 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4454 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4455 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C4457 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4458 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.02fF
C4459 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.01fF
C4460 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C4461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4462 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# 0.00fF
C4463 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C4464 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C4465 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4466 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4467 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4468 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C4469 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.00fF
C4470 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C4471 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.42fF
C4472 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C4473 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C4474 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C4475 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C4476 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4477 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4478 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4479 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C4480 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C4481 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4482 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C4483 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4484 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C4485 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4486 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# -0.00fF
C4487 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.02fF
C4488 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C4489 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.01fF
C4490 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C4491 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C4492 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4493 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C4494 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.02fF
C4495 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.02fF
C4496 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4497 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C4498 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C4499 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4500 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.02fF
C4501 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4502 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C4503 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C4504 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4505 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.57fF
C4506 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C4507 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C4508 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C4509 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4510 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4511 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C4512 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4513 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C4514 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C4515 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C4516 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4517 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C4518 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C4519 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C4520 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4521 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4522 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C4523 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# 0.01fF
C4524 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4525 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C4526 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4527 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C4528 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C4529 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C4530 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C4531 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C4532 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C4533 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.01fF
C4534 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C4535 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C4536 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4537 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C4538 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C4539 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C4540 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C4541 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.01fF
C4542 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4543 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C4544 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C4545 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C4546 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4547 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4548 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.00fF
C4549 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4550 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4551 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4552 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4553 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4554 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C4555 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4556 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C4557 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C4558 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C4559 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4560 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.01fF
C4561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C4562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C4563 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# -0.01fF
C4564 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4565 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.01fF
C4566 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C4567 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C4568 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C4569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C4570 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4571 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.00fF
C4572 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.02fF
C4573 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.22fF
C4574 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C4575 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C4576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C4577 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.02fF
C4578 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# 0.00fF
C4579 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C4580 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4581 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4582 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# 0.02fF
C4583 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C4584 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C4585 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C4586 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C4587 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C4588 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4589 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C4590 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C4591 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C4592 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4593 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.00fF
C4594 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C4595 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C4596 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.01fF
C4597 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4598 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4599 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.02fF
C4600 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4601 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4602 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C4603 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4604 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4605 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C4606 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4607 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C4608 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C4609 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.24fF
C4610 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4611 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C4612 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C4613 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C4614 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.00fF
C4615 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4616 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# -0.00fF
C4617 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4618 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4619 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4620 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C4621 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C4622 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4623 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4624 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C4625 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C4626 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C4627 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C4628 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4629 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C4630 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C4631 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C4632 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.01fF
C4633 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4634 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C4635 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# -0.00fF
C4636 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4637 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C4638 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C4639 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C4640 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C4641 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C4642 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C4643 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C4644 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4645 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C4646 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4647 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4648 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4649 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4650 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4651 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4652 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4653 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.02fF
C4654 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# -0.00fF
C4655 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C4656 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C4657 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.01fF
C4658 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4659 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C4660 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.01fF
C4661 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C4662 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4663 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.02fF
C4664 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C4665 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C4666 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.19fF
C4667 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# -0.01fF
C4668 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C4669 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4671 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4672 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.02fF
C4673 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.02fF
C4674 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C4675 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C4677 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C4678 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4679 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4680 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4681 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C4682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C4683 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C4684 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# 0.00fF
C4685 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C4686 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4687 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C4688 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C4689 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C4690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C4691 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4692 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4693 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.22fF
C4694 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C4695 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4696 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.01fF
C4697 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C4698 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4699 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# 0.00fF
C4700 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4701 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# -0.00fF
C4702 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.01fF
C4703 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C4704 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C4705 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C4706 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4707 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4708 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4709 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# 0.00fF
C4710 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4711 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C4712 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C4713 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C4714 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C4715 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C4716 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C4717 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.00fF
C4718 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C4719 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4720 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4721 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C4722 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C4723 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C4724 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4726 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4727 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# -0.00fF
C4728 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C4729 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C4730 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4731 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C4732 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.02fF
C4733 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.02fF
C4734 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C4735 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C4736 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.02fF
C4737 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C4738 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4739 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4740 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4741 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# -0.00fF
C4742 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C4743 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# 0.00fF
C4744 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# 0.00fF
C4745 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# -0.00fF
C4746 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# -0.00fF
C4747 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C4748 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4749 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C4750 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.46fF
C4751 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4752 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4753 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4754 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4755 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4756 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C4757 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C4758 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4759 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4760 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C4761 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4762 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4763 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.02fF
C4764 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C4765 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C4766 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.02fF
C4767 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.02fF
C4768 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C4769 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C4770 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4771 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4772 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4773 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4774 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.00fF
C4775 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.42fF
C4776 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C4777 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C4778 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C4779 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C4780 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4781 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4782 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4783 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C4784 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C4785 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4786 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C4787 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C4788 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4789 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C4790 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C4791 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C4792 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C4793 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C4794 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C4795 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4796 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4797 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C4798 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C4799 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.01fF
C4800 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C4801 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# -0.00fF
C4802 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4803 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C4804 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C4805 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# -0.00fF
C4806 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4807 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.02fF
C4808 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4809 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.42fF
C4810 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C4811 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4812 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4813 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4814 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C4815 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4816 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C4817 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C4818 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.01fF
C4819 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4820 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4821 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.01fF
C4822 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C4823 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C4824 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C4825 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C4826 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C4827 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C4828 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C4829 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.02fF
C4830 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C4831 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4832 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4833 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C4834 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C4835 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C4836 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.02fF
C4837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C4838 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4839 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C4840 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C4841 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C4842 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.01fF
C4843 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C4844 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C4845 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.02fF
C4846 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C4847 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4848 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4849 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C4850 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4851 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4852 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4853 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C4854 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C4855 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4856 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# VSUBS 1.08fF
C4857 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# VSUBS 1.03fF
C4858 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# VSUBS 0.11fF
C4859 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# VSUBS 0.17fF
C4860 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# VSUBS 0.10fF
C4861 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# VSUBS 0.09fF
C4862 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# VSUBS 0.11fF
C4863 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# VSUBS 0.11fF
C4864 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# VSUBS 0.12fF
C4865 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# VSUBS 0.11fF
C4866 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# VSUBS 0.12fF
C4867 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# VSUBS 0.12fF
C4868 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# VSUBS 0.12fF
C4869 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# VSUBS 0.12fF
C4870 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# VSUBS 0.12fF
C4871 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# VSUBS 0.12fF
C4872 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# VSUBS 0.12fF
C4873 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# VSUBS 0.12fF
C4874 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# VSUBS 0.12fF
C4875 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# VSUBS 0.12fF
C4876 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# VSUBS 0.12fF
C4877 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# VSUBS 0.12fF
C4878 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# VSUBS 0.12fF
C4879 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# VSUBS 0.12fF
C4880 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# VSUBS 0.12fF
C4881 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# VSUBS 0.12fF
C4882 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# VSUBS 0.12fF
C4883 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# VSUBS 0.12fF
C4884 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# VSUBS 0.12fF
C4885 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# VSUBS 0.12fF
C4886 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# VSUBS 0.12fF
C4887 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# VSUBS 0.12fF
C4888 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# VSUBS 0.12fF
C4889 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# VSUBS 0.12fF
C4890 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# VSUBS 0.12fF
C4891 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# VSUBS 0.12fF
C4892 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# VSUBS 0.12fF
C4893 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# VSUBS 0.12fF
C4894 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# VSUBS 0.12fF
C4895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# VSUBS 0.12fF
C4896 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# VSUBS 0.12fF
C4897 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# VSUBS 0.12fF
C4898 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# VSUBS 0.20fF
C4899 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# VSUBS 0.13fF
C4900 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# VSUBS 1.08fF
C4901 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# VSUBS 1.03fF
C4902 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# VSUBS 0.11fF
C4903 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# VSUBS 0.17fF
C4904 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# VSUBS 0.10fF
C4905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# VSUBS 0.09fF
C4906 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# VSUBS 0.11fF
C4907 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# VSUBS 0.11fF
C4908 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# VSUBS 0.12fF
C4909 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# VSUBS 0.11fF
C4910 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# VSUBS 0.12fF
C4911 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# VSUBS 0.12fF
C4912 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# VSUBS 0.12fF
C4913 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# VSUBS 0.12fF
C4914 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# VSUBS 0.12fF
C4915 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# VSUBS 0.12fF
C4916 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# VSUBS 0.12fF
C4917 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# VSUBS 0.12fF
C4918 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# VSUBS 0.12fF
C4919 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# VSUBS 0.12fF
C4920 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# VSUBS 0.12fF
C4921 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# VSUBS 0.12fF
C4922 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# VSUBS 0.12fF
C4923 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# VSUBS 0.12fF
C4924 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# VSUBS 0.12fF
C4925 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# VSUBS 0.12fF
C4926 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# VSUBS 0.12fF
C4927 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# VSUBS 0.12fF
C4928 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# VSUBS 0.12fF
C4929 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# VSUBS 0.12fF
C4930 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# VSUBS 0.12fF
C4931 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# VSUBS 0.12fF
C4932 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# VSUBS 0.12fF
C4933 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# VSUBS 0.12fF
C4934 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# VSUBS 0.12fF
C4935 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# VSUBS 0.12fF
C4936 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# VSUBS 0.12fF
C4937 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# VSUBS 0.12fF
C4938 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# VSUBS 0.12fF
C4939 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# VSUBS 0.12fF
C4940 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# VSUBS 0.12fF
C4941 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# VSUBS 0.12fF
C4942 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# VSUBS 0.20fF
C4943 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# VSUBS 0.13fF
C4944 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# VSUBS 1.08fF
C4945 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# VSUBS 1.03fF
C4946 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# VSUBS 0.11fF
C4947 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# VSUBS 0.17fF
C4948 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# VSUBS 0.10fF
C4949 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# VSUBS 0.09fF
C4950 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# VSUBS 0.11fF
C4951 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# VSUBS 0.11fF
C4952 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# VSUBS 0.12fF
C4953 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# VSUBS 0.11fF
C4954 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# VSUBS 0.12fF
C4955 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# VSUBS 0.12fF
C4956 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# VSUBS 0.12fF
C4957 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# VSUBS 0.12fF
C4958 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# VSUBS 0.12fF
C4959 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# VSUBS 0.12fF
C4960 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# VSUBS 0.12fF
C4961 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# VSUBS 0.12fF
C4962 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# VSUBS 0.12fF
C4963 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# VSUBS 0.12fF
C4964 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# VSUBS 0.12fF
C4965 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# VSUBS 0.12fF
C4966 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# VSUBS 0.12fF
C4967 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# VSUBS 0.12fF
C4968 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# VSUBS 0.12fF
C4969 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# VSUBS 0.12fF
C4970 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# VSUBS 0.12fF
C4971 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# VSUBS 0.12fF
C4972 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# VSUBS 0.12fF
C4973 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# VSUBS 0.12fF
C4974 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# VSUBS 0.12fF
C4975 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# VSUBS 0.12fF
C4976 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# VSUBS 0.12fF
C4977 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# VSUBS 0.12fF
C4978 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# VSUBS 0.12fF
C4979 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# VSUBS 0.12fF
C4980 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# VSUBS 0.12fF
C4981 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# VSUBS 0.12fF
C4982 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# VSUBS 0.12fF
C4983 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# VSUBS 0.12fF
C4984 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# VSUBS 0.12fF
C4985 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# VSUBS 0.12fF
C4986 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# VSUBS 0.20fF
C4987 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# VSUBS 0.13fF
C4988 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# VSUBS 1.08fF
C4989 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# VSUBS 1.03fF
C4990 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# VSUBS 0.11fF
C4991 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# VSUBS 0.17fF
C4992 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# VSUBS 0.10fF
C4993 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# VSUBS 0.09fF
C4994 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# VSUBS 0.11fF
C4995 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# VSUBS 0.11fF
C4996 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# VSUBS 0.12fF
C4997 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# VSUBS 0.11fF
C4998 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# VSUBS 0.12fF
C4999 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# VSUBS 0.12fF
C5000 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# VSUBS 0.12fF
C5001 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# VSUBS 0.12fF
C5002 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# VSUBS 0.12fF
C5003 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# VSUBS 0.12fF
C5004 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# VSUBS 0.12fF
C5005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# VSUBS 0.12fF
C5006 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# VSUBS 0.12fF
C5007 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# VSUBS 0.12fF
C5008 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# VSUBS 0.12fF
C5009 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# VSUBS 0.12fF
C5010 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# VSUBS 0.12fF
C5011 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# VSUBS 0.12fF
C5012 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# VSUBS 0.12fF
C5013 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# VSUBS 0.12fF
C5014 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# VSUBS 0.12fF
C5015 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# VSUBS 0.12fF
C5016 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# VSUBS 0.12fF
C5017 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# VSUBS 0.12fF
C5018 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# VSUBS 0.12fF
C5019 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# VSUBS 0.12fF
C5020 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# VSUBS 0.12fF
C5021 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# VSUBS 0.12fF
C5022 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# VSUBS 0.12fF
C5023 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# VSUBS 0.12fF
C5024 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# VSUBS 0.12fF
C5025 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# VSUBS 0.12fF
C5026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# VSUBS 0.12fF
C5027 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# VSUBS 0.12fF
C5028 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# VSUBS 0.12fF
C5029 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# VSUBS 0.12fF
C5030 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# VSUBS 0.20fF
C5031 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# VSUBS 0.13fF
C5032 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# VSUBS 1.08fF
C5033 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# VSUBS 1.03fF
C5034 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# VSUBS 0.11fF
C5035 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# VSUBS 0.17fF
C5036 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# VSUBS 0.10fF
C5037 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# VSUBS 0.09fF
C5038 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# VSUBS 0.11fF
C5039 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# VSUBS 0.11fF
C5040 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# VSUBS 0.12fF
C5041 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# VSUBS 0.11fF
C5042 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# VSUBS 0.12fF
C5043 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# VSUBS 0.12fF
C5044 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# VSUBS 0.12fF
C5045 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# VSUBS 0.12fF
C5046 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# VSUBS 0.12fF
C5047 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# VSUBS 0.12fF
C5048 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# VSUBS 0.12fF
C5049 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# VSUBS 0.12fF
C5050 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# VSUBS 0.12fF
C5051 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# VSUBS 0.12fF
C5052 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# VSUBS 0.12fF
C5053 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# VSUBS 0.12fF
C5054 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# VSUBS 0.12fF
C5055 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# VSUBS 0.12fF
C5056 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# VSUBS 0.12fF
C5057 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# VSUBS 0.12fF
C5058 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# VSUBS 0.12fF
C5059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# VSUBS 0.12fF
C5060 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# VSUBS 0.12fF
C5061 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# VSUBS 0.12fF
C5062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# VSUBS 0.12fF
C5063 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# VSUBS 0.12fF
C5064 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# VSUBS 0.12fF
C5065 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# VSUBS 0.12fF
C5066 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# VSUBS 0.12fF
C5067 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# VSUBS 0.12fF
C5068 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# VSUBS 0.12fF
C5069 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# VSUBS 0.12fF
C5070 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# VSUBS 0.12fF
C5071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# VSUBS 0.12fF
C5072 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# VSUBS 0.12fF
C5073 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# VSUBS 0.12fF
C5074 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# VSUBS 0.20fF
C5075 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# VSUBS 0.13fF
C5076 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# VSUBS 1.08fF
C5077 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# VSUBS 1.03fF
C5078 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# VSUBS 0.11fF
C5079 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# VSUBS 0.17fF
C5080 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# VSUBS 0.10fF
C5081 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# VSUBS 0.09fF
C5082 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# VSUBS 0.11fF
C5083 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# VSUBS 0.11fF
C5084 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# VSUBS 0.12fF
C5085 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# VSUBS 0.11fF
C5086 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# VSUBS 0.12fF
C5087 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# VSUBS 0.12fF
C5088 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# VSUBS 0.12fF
C5089 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# VSUBS 0.12fF
C5090 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# VSUBS 0.12fF
C5091 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# VSUBS 0.12fF
C5092 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# VSUBS 0.12fF
C5093 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# VSUBS 0.12fF
C5094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# VSUBS 0.12fF
C5095 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# VSUBS 0.12fF
C5096 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# VSUBS 0.12fF
C5097 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# VSUBS 0.12fF
C5098 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# VSUBS 0.12fF
C5099 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# VSUBS 0.12fF
C5100 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# VSUBS 0.12fF
C5101 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# VSUBS 0.12fF
C5102 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# VSUBS 0.12fF
C5103 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# VSUBS 0.12fF
C5104 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# VSUBS 0.12fF
C5105 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# VSUBS 0.12fF
C5106 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# VSUBS 0.12fF
C5107 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# VSUBS 0.12fF
C5108 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# VSUBS 0.12fF
C5109 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# VSUBS 0.12fF
C5110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# VSUBS 0.12fF
C5111 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# VSUBS 0.12fF
C5112 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# VSUBS 0.12fF
C5113 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# VSUBS 0.12fF
C5114 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# VSUBS 0.12fF
C5115 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# VSUBS 0.12fF
C5116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# VSUBS 0.12fF
C5117 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# VSUBS 0.12fF
C5118 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# VSUBS 0.20fF
C5119 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# VSUBS 0.13fF
C5120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# VSUBS 1.08fF
C5121 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# VSUBS 1.03fF
C5122 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# VSUBS 0.11fF
C5123 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# VSUBS 0.17fF
C5124 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# VSUBS 0.10fF
C5125 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# VSUBS 0.09fF
C5126 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# VSUBS 0.11fF
C5127 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# VSUBS 0.11fF
C5128 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# VSUBS 0.12fF
C5129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# VSUBS 0.11fF
C5130 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# VSUBS 0.12fF
C5131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# VSUBS 0.12fF
C5132 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# VSUBS 0.12fF
C5133 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# VSUBS 0.12fF
C5134 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# VSUBS 0.12fF
C5135 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# VSUBS 0.12fF
C5136 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# VSUBS 0.12fF
C5137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# VSUBS 0.12fF
C5138 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# VSUBS 0.12fF
C5139 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# VSUBS 0.12fF
C5140 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# VSUBS 0.12fF
C5141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# VSUBS 0.12fF
C5142 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# VSUBS 0.12fF
C5143 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# VSUBS 0.12fF
C5144 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# VSUBS 0.12fF
C5145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# VSUBS 0.12fF
C5146 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# VSUBS 0.12fF
C5147 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# VSUBS 0.12fF
C5148 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# VSUBS 0.12fF
C5149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# VSUBS 0.12fF
C5150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# VSUBS 0.12fF
C5151 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# VSUBS 0.12fF
C5152 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# VSUBS 0.12fF
C5153 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# VSUBS 0.12fF
C5154 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# VSUBS 0.12fF
C5155 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# VSUBS 0.12fF
C5156 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# VSUBS 0.12fF
C5157 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# VSUBS 0.12fF
C5158 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# VSUBS 0.12fF
C5159 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# VSUBS 0.12fF
C5160 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# VSUBS 0.12fF
C5161 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# VSUBS 0.12fF
C5162 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# VSUBS 0.20fF
C5163 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# VSUBS 0.13fF
C5164 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# VSUBS 1.08fF
C5165 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# VSUBS 1.03fF
C5166 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# VSUBS 0.11fF
C5167 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# VSUBS 0.17fF
C5168 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# VSUBS 0.10fF
C5169 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# VSUBS 0.09fF
C5170 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# VSUBS 0.11fF
C5171 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# VSUBS 0.11fF
C5172 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# VSUBS 0.12fF
C5173 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# VSUBS 0.11fF
C5174 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# VSUBS 0.12fF
C5175 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# VSUBS 0.12fF
C5176 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# VSUBS 0.12fF
C5177 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# VSUBS 0.12fF
C5178 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# VSUBS 0.12fF
C5179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# VSUBS 0.12fF
C5180 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# VSUBS 0.12fF
C5181 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# VSUBS 0.12fF
C5182 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# VSUBS 0.12fF
C5183 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# VSUBS 0.12fF
C5184 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# VSUBS 0.12fF
C5185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# VSUBS 0.12fF
C5186 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# VSUBS 0.12fF
C5187 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# VSUBS 0.12fF
C5188 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# VSUBS 0.12fF
C5189 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# VSUBS 0.12fF
C5190 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# VSUBS 0.12fF
C5191 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# VSUBS 0.12fF
C5192 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# VSUBS 0.12fF
C5193 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# VSUBS 0.12fF
C5194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# VSUBS 0.12fF
C5195 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# VSUBS 0.12fF
C5196 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# VSUBS 0.12fF
C5197 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# VSUBS 0.12fF
C5198 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# VSUBS 0.12fF
C5199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# VSUBS 0.12fF
C5200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# VSUBS 0.12fF
C5201 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# VSUBS 0.12fF
C5202 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# VSUBS 0.12fF
C5203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# VSUBS 0.12fF
C5204 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# VSUBS 0.12fF
C5205 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# VSUBS 0.12fF
C5206 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# VSUBS 0.20fF
C5207 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# VSUBS 0.13fF
.ends

.subckt comparator_v2 clk ip in outp outn VDD VSS
Xlatch_pmos_pair_0 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD VDD VDD
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD latch_pmos_pair
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__buf_2_1/X outp VSS VDD outn VSS VDD sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__buf_2_0/X outn VSS VDD outp VSS VDD sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_pr__pfet_01v8_VCG74W_1 li_940_3458# li_940_3458# li_940_3458# clk VDD VDD
+ clk clk li_940_3458# li_940_3458# li_940_3458# clk VDD VDD clk clk VDD li_940_3458#
+ clk clk VDD clk clk clk VDD VDD clk clk li_940_3458# li_940_3458# clk VDD clk clk
+ VSS sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk VDD sky130_fd_sc_hd__buf_2_1/A clk
+ clk VDD clk clk clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ clk VDD clk clk VSS sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_sc_hd__buf_2_0 sky130_fd_sc_hd__buf_2_0/A VSS VDD sky130_fd_sc_hd__buf_2_0/X
+ VSS VDD sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_1 sky130_fd_sc_hd__buf_2_1/A VSS VDD sky130_fd_sc_hd__buf_2_1/X
+ VSS VDD sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_0 clk sky130_fd_sc_hd__buf_2_0/A clk VDD VDD clk sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A clk sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A clk clk VDD VDD clk clk clk sky130_fd_sc_hd__buf_2_0/A
+ clk clk clk clk VSS precharge_pmos
Xcurrent_tail_0 li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# VSS VSS VSS
+ li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS VSS VSS li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS li_n2324_818# li_n2324_818# VSS VSS VSS clk li_n2324_818# VSS current_tail
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_1 clk li_940_818# clk VDD VDD clk li_940_818# li_940_818# li_940_818#
+ clk li_940_818# VDD VDD clk VDD VDD clk clk li_940_818# VDD li_940_818# li_940_818#
+ clk clk VDD VDD clk clk clk li_940_818# clk clk clk clk VSS precharge_pmos
Xlatch_nmos_pair_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A latch_nmos_pair
Xinput_diff_pair_0 ip ip ip in in VSS ip in in in in VSS li_940_3458# ip ip ip in
+ ip li_n2324_818# ip ip in ip ip ip in in in ip ip ip in ip in ip in ip in in ip
+ ip VSS ip ip in ip li_n2324_818# ip ip in in in ip ip ip in in in li_940_3458# in
+ in ip ip in ip in ip ip ip VSS ip in ip ip ip in in in ip ip in in ip in VSS ip
+ in in in in in ip in li_940_818# ip ip in ip ip li_n2324_818# in in ip ip ip in
+ ip ip ip ip in in in in in in VSS ip in in ip ip ip ip ip in in ip ip in in ip li_940_818#
+ ip ip in li_n2324_818# in in in VSS ip in in ip ip ip in ip ip ip in in ip in ip
+ in ip ip ip in in in in in VSS in ip li_n2324_818# ip ip in ip ip in ip ip in ip
+ ip li_940_3458# in in ip ip ip in in in ip ip in ip ip in in in VSS ip in VSS VSS
+ in in ip ip in in ip ip ip in in ip ip li_940_3458# in ip in ip ip in li_n2324_818#
+ ip in in in in in in ip ip in in ip ip ip ip VSS ip ip ip in in in in ip ip in ip
+ ip ip in in ip ip in in ip in in li_n2324_818# in in in in ip in in ip in ip li_940_818#
+ VSS ip ip ip ip in in ip ip VSS in in in ip in in ip ip ip in in ip in in VSS in
+ in li_n2324_818# ip in in in ip ip ip ip in in ip ip li_940_818# in ip ip in in
+ in ip in ip in ip ip ip in in in ip ip ip ip in in in ip ip in in in in ip VSS VSS
+ in in ip ip in in in input_diff_pair
C0 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_1/a_27_47# 0.02fF
C1 outp sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.08fF
C2 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_1/a_27_47# 0.06fF
C3 sky130_fd_sc_hd__buf_2_0/a_27_47# outp 0.04fF
C4 sky130_fd_sc_hd__nand2_4_0/a_27_47# VDD 0.01fF
C5 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.00fF
C6 sky130_fd_sc_hd__buf_2_0/a_27_47# VDD 0.07fF
C7 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.02fF
C8 outp sky130_fd_sc_hd__buf_2_1/a_27_47# 0.02fF
C9 li_n2324_818# VDD 0.09fF
C10 li_n2324_818# sky130_fd_sc_hd__buf_2_1/A 0.95fF
C11 sky130_fd_sc_hd__buf_2_1/a_27_47# VDD 0.09fF
C12 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.03fF
C13 outp VDD 0.83fF
C14 outp sky130_fd_sc_hd__buf_2_1/A 0.05fF
C15 sky130_fd_sc_hd__nand2_4_0/a_27_47# outn 0.18fF
C16 VDD sky130_fd_sc_hd__buf_2_1/A 26.23fF
C17 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_1/X 0.05fF
C18 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.00fF
C19 sky130_fd_sc_hd__buf_2_0/a_27_47# outn 0.02fF
C20 li_n2324_818# li_940_818# 2.99fF
C21 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.01fF
C22 sky130_fd_sc_hd__buf_2_1/a_27_47# outn 0.04fF
C23 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_1/X 0.11fF
C24 outp outn 1.34fF
C25 li_n2324_818# sky130_fd_sc_hd__buf_2_0/A 1.31fF
C26 VDD li_940_818# 2.08fF
C27 li_940_818# sky130_fd_sc_hd__buf_2_1/A 21.09fF
C28 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.02fF
C29 outp sky130_fd_sc_hd__buf_2_1/X 0.03fF
C30 outp sky130_fd_sc_hd__buf_2_0/A 0.04fF
C31 sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.28fF
C32 VDD outn 0.93fF
C33 outn sky130_fd_sc_hd__buf_2_1/A 0.03fF
C34 VDD sky130_fd_sc_hd__buf_2_1/X 0.24fF
C35 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_1/A 0.09fF
C36 sky130_fd_sc_hd__buf_2_0/A VDD 30.94fF
C37 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A 76.01fF
C38 sky130_fd_sc_hd__buf_2_0/a_27_47# VSS 0.03fF
C39 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.03fF
C40 li_n2324_818# ip 48.05fF
C41 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.02fF
C42 li_n2324_818# VSS 3.07fF
C43 sky130_fd_sc_hd__buf_2_1/a_27_47# VSS 0.04fF
C44 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.01fF
C45 outp VSS 0.43fF
C46 VDD ip 0.03fF
C47 sky130_fd_sc_hd__buf_2_1/A ip 1.73fF
C48 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_0/X 0.11fF
C49 sky130_fd_sc_hd__buf_2_0/A li_940_818# 9.11fF
C50 li_n2324_818# clk 6.65fF
C51 VDD VSS 0.85fF
C52 sky130_fd_sc_hd__buf_2_1/A VSS 1.57fF
C53 outp sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.09fF
C54 outn sky130_fd_sc_hd__buf_2_1/X 0.23fF
C55 sky130_fd_sc_hd__buf_2_0/A outn 0.05fF
C56 li_940_3458# li_n2324_818# 4.64fF
C57 li_n2324_818# in 49.83fF
C58 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/X 0.06fF
C59 sky130_fd_sc_hd__nand2_4_1/a_27_47# VDD 0.02fF
C60 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.00fF
C61 clk VDD 14.94fF
C62 clk sky130_fd_sc_hd__buf_2_1/A 3.02fF
C63 outp sky130_fd_sc_hd__buf_2_0/X 0.20fF
C64 li_940_818# ip 35.81fF
C65 li_940_3458# VDD 2.17fF
C66 li_940_3458# sky130_fd_sc_hd__buf_2_1/A 9.09fF
C67 in VDD 0.01fF
C68 in sky130_fd_sc_hd__buf_2_1/A 0.67fF
C69 sky130_fd_sc_hd__buf_2_0/X VDD 0.20fF
C70 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_1/A 0.04fF
C71 li_940_818# VSS 0.96fF
C72 sky130_fd_sc_hd__buf_2_0/A ip 2.05fF
C73 outn VSS 0.55fF
C74 sky130_fd_sc_hd__buf_2_1/X VSS 0.05fF
C75 sky130_fd_sc_hd__buf_2_0/A VSS 2.10fF
C76 clk li_940_818# 4.03fF
C77 sky130_fd_sc_hd__nand2_4_1/a_27_47# outn 0.06fF
C78 li_940_3458# li_940_818# 4.44fF
C79 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_1/X 0.01fF
C80 in li_940_818# 12.98fF
C81 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.00fF
C82 clk sky130_fd_sc_hd__buf_2_0/A 3.32fF
C83 sky130_fd_sc_hd__buf_2_0/X outn 0.03fF
C84 ip VSS 2.78fF
C85 li_940_3458# sky130_fd_sc_hd__buf_2_0/A 18.81fF
C86 in sky130_fd_sc_hd__buf_2_0/A 1.07fF
C87 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_1/X 0.11fF
C88 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_0/A 0.10fF
C89 clk ip 0.62fF
C90 sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.24fF
C91 li_940_3458# ip 13.70fF
C92 in ip 30.51fF
C93 clk VSS 1.71fF
C94 li_940_3458# VSS 1.22fF
C95 in VSS 1.52fF
C96 sky130_fd_sc_hd__buf_2_0/X VSS 0.04fF
C97 li_940_3458# clk 2.08fF
C98 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.03fF
C99 in clk 0.47fF
C100 li_940_3458# in 37.79fF
C101 li_940_3458# 0 -1592.65fF
C102 li_940_818# 0 -2262.83fF
C103 outn 0 21.73fF
C104 in 0 -297.33fF
C105 li_n2324_818# 0 -3722.01fF
C106 ip 0 -420.77fF
C107 VSS 0 -70.44fF
C108 sky130_fd_sc_hd__buf_2_0/A 0 -127.11fF
C109 sky130_fd_sc_hd__buf_2_1/A 0 -211.82fF
C110 VDD 0 -582.64fF
C111 clk 0 68.21fF
C112 sky130_fd_sc_hd__buf_2_1/X 0 23.78fF
C113 sky130_fd_sc_hd__buf_2_1/a_27_47# 0 0.15fF
C114 sky130_fd_sc_hd__buf_2_0/X 0 43.25fF
C115 sky130_fd_sc_hd__buf_2_0/a_27_47# 0 0.15fF
C116 sky130_fd_sc_hd__nand2_4_1/a_27_47# 0 0.06fF
C117 outp 0 26.35fF
C118 sky130_fd_sc_hd__nand2_4_0/a_27_47# 0 0.06fF
.ends

