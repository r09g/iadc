magic
tech sky130A
magscale 1 2
timestamp 1654601900
<< error_p >>
rect -4124 181 -4066 187
rect -3704 181 -3646 187
rect -3284 181 -3226 187
rect -2864 181 -2806 187
rect -2444 181 -2386 187
rect -2024 181 -1966 187
rect -1604 181 -1546 187
rect -1184 181 -1126 187
rect -764 181 -706 187
rect -344 181 -286 187
rect 76 181 134 187
rect 496 181 554 187
rect 916 181 974 187
rect 1336 181 1394 187
rect 1756 181 1814 187
rect 2176 181 2234 187
rect 2596 181 2654 187
rect 3016 181 3074 187
rect 3436 181 3494 187
rect 3856 181 3914 187
rect -4124 147 -4112 181
rect -3704 147 -3692 181
rect -3284 147 -3272 181
rect -2864 147 -2852 181
rect -2444 147 -2432 181
rect -2024 147 -2012 181
rect -1604 147 -1592 181
rect -1184 147 -1172 181
rect -764 147 -752 181
rect -344 147 -332 181
rect 76 147 88 181
rect 496 147 508 181
rect 916 147 928 181
rect 1336 147 1348 181
rect 1756 147 1768 181
rect 2176 147 2188 181
rect 2596 147 2608 181
rect 3016 147 3028 181
rect 3436 147 3448 181
rect 3856 147 3868 181
rect -4124 141 -4066 147
rect -3704 141 -3646 147
rect -3284 141 -3226 147
rect -2864 141 -2806 147
rect -2444 141 -2386 147
rect -2024 141 -1966 147
rect -1604 141 -1546 147
rect -1184 141 -1126 147
rect -764 141 -706 147
rect -344 141 -286 147
rect 76 141 134 147
rect 496 141 554 147
rect 916 141 974 147
rect 1336 141 1394 147
rect 1756 141 1814 147
rect 2176 141 2234 147
rect 2596 141 2654 147
rect 3016 141 3074 147
rect 3436 141 3494 147
rect 3856 141 3914 147
rect -3914 -147 -3856 -141
rect -3494 -147 -3436 -141
rect -3074 -147 -3016 -141
rect -2654 -147 -2596 -141
rect -2234 -147 -2176 -141
rect -1814 -147 -1756 -141
rect -1394 -147 -1336 -141
rect -974 -147 -916 -141
rect -554 -147 -496 -141
rect -134 -147 -76 -141
rect 286 -147 344 -141
rect 706 -147 764 -141
rect 1126 -147 1184 -141
rect 1546 -147 1604 -141
rect 1966 -147 2024 -141
rect 2386 -147 2444 -141
rect 2806 -147 2864 -141
rect 3226 -147 3284 -141
rect 3646 -147 3704 -141
rect 4066 -147 4124 -141
rect -3914 -181 -3902 -147
rect -3494 -181 -3482 -147
rect -3074 -181 -3062 -147
rect -2654 -181 -2642 -147
rect -2234 -181 -2222 -147
rect -1814 -181 -1802 -147
rect -1394 -181 -1382 -147
rect -974 -181 -962 -147
rect -554 -181 -542 -147
rect -134 -181 -122 -147
rect 286 -181 298 -147
rect 706 -181 718 -147
rect 1126 -181 1138 -147
rect 1546 -181 1558 -147
rect 1966 -181 1978 -147
rect 2386 -181 2398 -147
rect 2806 -181 2818 -147
rect 3226 -181 3238 -147
rect 3646 -181 3658 -147
rect 4066 -181 4078 -147
rect -3914 -187 -3856 -181
rect -3494 -187 -3436 -181
rect -3074 -187 -3016 -181
rect -2654 -187 -2596 -181
rect -2234 -187 -2176 -181
rect -1814 -187 -1756 -181
rect -1394 -187 -1336 -181
rect -974 -187 -916 -181
rect -554 -187 -496 -181
rect -134 -187 -76 -181
rect 286 -187 344 -181
rect 706 -187 764 -181
rect 1126 -187 1184 -181
rect 1546 -187 1604 -181
rect 1966 -187 2024 -181
rect 2386 -187 2444 -181
rect 2806 -187 2864 -181
rect 3226 -187 3284 -181
rect 3646 -187 3704 -181
rect 4066 -187 4124 -181
rect -4122 -351 -4064 -345
rect -3702 -351 -3644 -345
rect -3282 -351 -3224 -345
rect -2862 -351 -2804 -345
rect -2442 -351 -2384 -345
rect -2022 -351 -1964 -345
rect -1602 -351 -1544 -345
rect -1182 -351 -1124 -345
rect -762 -351 -704 -345
rect -342 -351 -284 -345
rect 78 -351 136 -345
rect 498 -351 556 -345
rect 918 -351 976 -345
rect 1338 -351 1396 -345
rect 1758 -351 1816 -345
rect 2178 -351 2236 -345
rect 2598 -351 2656 -345
rect 3018 -351 3076 -345
rect 3438 -351 3496 -345
rect 3858 -351 3916 -345
rect -4122 -385 -4110 -351
rect -3702 -385 -3690 -351
rect -3282 -385 -3270 -351
rect -2862 -385 -2850 -351
rect -2442 -385 -2430 -351
rect -2022 -385 -2010 -351
rect -1602 -385 -1590 -351
rect -1182 -385 -1170 -351
rect -762 -385 -750 -351
rect -342 -385 -330 -351
rect 78 -385 90 -351
rect 498 -385 510 -351
rect 918 -385 930 -351
rect 1338 -385 1350 -351
rect 1758 -385 1770 -351
rect 2178 -385 2190 -351
rect 2598 -385 2610 -351
rect 3018 -385 3030 -351
rect 3438 -385 3450 -351
rect 3858 -385 3870 -351
rect -4122 -391 -4064 -385
rect -3702 -391 -3644 -385
rect -3282 -391 -3224 -385
rect -2862 -391 -2804 -385
rect -2442 -391 -2384 -385
rect -2022 -391 -1964 -385
rect -1602 -391 -1544 -385
rect -1182 -391 -1124 -385
rect -762 -391 -704 -385
rect -342 -391 -284 -385
rect 78 -391 136 -385
rect 498 -391 556 -385
rect 918 -391 976 -385
rect 1338 -391 1396 -385
rect 1758 -391 1816 -385
rect 2178 -391 2236 -385
rect 2598 -391 2656 -385
rect 3018 -391 3076 -385
rect 3438 -391 3496 -385
rect 3858 -391 3916 -385
rect -3912 -679 -3854 -673
rect -3492 -679 -3434 -673
rect -3072 -679 -3014 -673
rect -2652 -679 -2594 -673
rect -2232 -679 -2174 -673
rect -1812 -679 -1754 -673
rect -1392 -679 -1334 -673
rect -972 -679 -914 -673
rect -552 -679 -494 -673
rect -132 -679 -74 -673
rect 288 -679 346 -673
rect 708 -679 766 -673
rect 1128 -679 1186 -673
rect 1548 -679 1606 -673
rect 1968 -679 2026 -673
rect 2388 -679 2446 -673
rect 2808 -679 2866 -673
rect 3228 -679 3286 -673
rect 3648 -679 3706 -673
rect 4068 -679 4126 -673
rect -3912 -713 -3900 -679
rect -3492 -713 -3480 -679
rect -3072 -713 -3060 -679
rect -2652 -713 -2640 -679
rect -2232 -713 -2220 -679
rect -1812 -713 -1800 -679
rect -1392 -713 -1380 -679
rect -972 -713 -960 -679
rect -552 -713 -540 -679
rect -132 -713 -120 -679
rect 288 -713 300 -679
rect 708 -713 720 -679
rect 1128 -713 1140 -679
rect 1548 -713 1560 -679
rect 1968 -713 1980 -679
rect 2388 -713 2400 -679
rect 2808 -713 2820 -679
rect 3228 -713 3240 -679
rect 3648 -713 3660 -679
rect 4068 -713 4080 -679
rect -3912 -719 -3854 -713
rect -3492 -719 -3434 -713
rect -3072 -719 -3014 -713
rect -2652 -719 -2594 -713
rect -2232 -719 -2174 -713
rect -1812 -719 -1754 -713
rect -1392 -719 -1334 -713
rect -972 -719 -914 -713
rect -552 -719 -494 -713
rect -132 -719 -74 -713
rect 288 -719 346 -713
rect 708 -719 766 -713
rect 1128 -719 1186 -713
rect 1548 -719 1606 -713
rect 1968 -719 2026 -713
rect 2388 -719 2446 -713
rect 2808 -719 2866 -713
rect 3228 -719 3286 -713
rect 3648 -719 3706 -713
rect 4068 -719 4126 -713
<< nwell >>
rect -4520 -851 4520 319
<< pmos >>
rect -4320 -100 -4290 100
rect -4110 -100 -4080 100
rect -3900 -100 -3870 100
rect -3690 -100 -3660 100
rect -3480 -100 -3450 100
rect -3270 -100 -3240 100
rect -3060 -100 -3030 100
rect -2850 -100 -2820 100
rect -2640 -100 -2610 100
rect -2430 -100 -2400 100
rect -2220 -100 -2190 100
rect -2010 -100 -1980 100
rect -1800 -100 -1770 100
rect -1590 -100 -1560 100
rect -1380 -100 -1350 100
rect -1170 -100 -1140 100
rect -960 -100 -930 100
rect -750 -100 -720 100
rect -540 -100 -510 100
rect -330 -100 -300 100
rect -120 -100 -90 100
rect 90 -100 120 100
rect 300 -100 330 100
rect 510 -100 540 100
rect 720 -100 750 100
rect 930 -100 960 100
rect 1140 -100 1170 100
rect 1350 -100 1380 100
rect 1560 -100 1590 100
rect 1770 -100 1800 100
rect 1980 -100 2010 100
rect 2190 -100 2220 100
rect 2400 -100 2430 100
rect 2610 -100 2640 100
rect 2820 -100 2850 100
rect 3030 -100 3060 100
rect 3240 -100 3270 100
rect 3450 -100 3480 100
rect 3660 -100 3690 100
rect 3870 -100 3900 100
rect 4080 -100 4110 100
rect 4290 -100 4320 100
rect -4318 -632 -4288 -432
rect -4108 -632 -4078 -432
rect -3898 -632 -3868 -432
rect -3688 -632 -3658 -432
rect -3478 -632 -3448 -432
rect -3268 -632 -3238 -432
rect -3058 -632 -3028 -432
rect -2848 -632 -2818 -432
rect -2638 -632 -2608 -432
rect -2428 -632 -2398 -432
rect -2218 -632 -2188 -432
rect -2008 -632 -1978 -432
rect -1798 -632 -1768 -432
rect -1588 -632 -1558 -432
rect -1378 -632 -1348 -432
rect -1168 -632 -1138 -432
rect -958 -632 -928 -432
rect -748 -632 -718 -432
rect -538 -632 -508 -432
rect -328 -632 -298 -432
rect -118 -632 -88 -432
rect 92 -632 122 -432
rect 302 -632 332 -432
rect 512 -632 542 -432
rect 722 -632 752 -432
rect 932 -632 962 -432
rect 1142 -632 1172 -432
rect 1352 -632 1382 -432
rect 1562 -632 1592 -432
rect 1772 -632 1802 -432
rect 1982 -632 2012 -432
rect 2192 -632 2222 -432
rect 2402 -632 2432 -432
rect 2612 -632 2642 -432
rect 2822 -632 2852 -432
rect 3032 -632 3062 -432
rect 3242 -632 3272 -432
rect 3452 -632 3482 -432
rect 3662 -632 3692 -432
rect 3872 -632 3902 -432
rect 4082 -632 4112 -432
rect 4292 -632 4322 -432
<< pdiff >>
rect -4382 88 -4320 100
rect -4382 -88 -4370 88
rect -4336 -88 -4320 88
rect -4382 -100 -4320 -88
rect -4290 88 -4228 100
rect -4290 -88 -4274 88
rect -4240 -88 -4228 88
rect -4290 -100 -4228 -88
rect -4172 88 -4110 100
rect -4172 -88 -4160 88
rect -4126 -88 -4110 88
rect -4172 -100 -4110 -88
rect -4080 88 -4018 100
rect -4080 -88 -4064 88
rect -4030 -88 -4018 88
rect -4080 -100 -4018 -88
rect -3962 88 -3900 100
rect -3962 -88 -3950 88
rect -3916 -88 -3900 88
rect -3962 -100 -3900 -88
rect -3870 88 -3808 100
rect -3870 -88 -3854 88
rect -3820 -88 -3808 88
rect -3870 -100 -3808 -88
rect -3752 88 -3690 100
rect -3752 -88 -3740 88
rect -3706 -88 -3690 88
rect -3752 -100 -3690 -88
rect -3660 88 -3598 100
rect -3660 -88 -3644 88
rect -3610 -88 -3598 88
rect -3660 -100 -3598 -88
rect -3542 88 -3480 100
rect -3542 -88 -3530 88
rect -3496 -88 -3480 88
rect -3542 -100 -3480 -88
rect -3450 88 -3388 100
rect -3450 -88 -3434 88
rect -3400 -88 -3388 88
rect -3450 -100 -3388 -88
rect -3332 88 -3270 100
rect -3332 -88 -3320 88
rect -3286 -88 -3270 88
rect -3332 -100 -3270 -88
rect -3240 88 -3178 100
rect -3240 -88 -3224 88
rect -3190 -88 -3178 88
rect -3240 -100 -3178 -88
rect -3122 88 -3060 100
rect -3122 -88 -3110 88
rect -3076 -88 -3060 88
rect -3122 -100 -3060 -88
rect -3030 88 -2968 100
rect -3030 -88 -3014 88
rect -2980 -88 -2968 88
rect -3030 -100 -2968 -88
rect -2912 88 -2850 100
rect -2912 -88 -2900 88
rect -2866 -88 -2850 88
rect -2912 -100 -2850 -88
rect -2820 88 -2758 100
rect -2820 -88 -2804 88
rect -2770 -88 -2758 88
rect -2820 -100 -2758 -88
rect -2702 88 -2640 100
rect -2702 -88 -2690 88
rect -2656 -88 -2640 88
rect -2702 -100 -2640 -88
rect -2610 88 -2548 100
rect -2610 -88 -2594 88
rect -2560 -88 -2548 88
rect -2610 -100 -2548 -88
rect -2492 88 -2430 100
rect -2492 -88 -2480 88
rect -2446 -88 -2430 88
rect -2492 -100 -2430 -88
rect -2400 88 -2338 100
rect -2400 -88 -2384 88
rect -2350 -88 -2338 88
rect -2400 -100 -2338 -88
rect -2282 88 -2220 100
rect -2282 -88 -2270 88
rect -2236 -88 -2220 88
rect -2282 -100 -2220 -88
rect -2190 88 -2128 100
rect -2190 -88 -2174 88
rect -2140 -88 -2128 88
rect -2190 -100 -2128 -88
rect -2072 88 -2010 100
rect -2072 -88 -2060 88
rect -2026 -88 -2010 88
rect -2072 -100 -2010 -88
rect -1980 88 -1918 100
rect -1980 -88 -1964 88
rect -1930 -88 -1918 88
rect -1980 -100 -1918 -88
rect -1862 88 -1800 100
rect -1862 -88 -1850 88
rect -1816 -88 -1800 88
rect -1862 -100 -1800 -88
rect -1770 88 -1708 100
rect -1770 -88 -1754 88
rect -1720 -88 -1708 88
rect -1770 -100 -1708 -88
rect -1652 88 -1590 100
rect -1652 -88 -1640 88
rect -1606 -88 -1590 88
rect -1652 -100 -1590 -88
rect -1560 88 -1498 100
rect -1560 -88 -1544 88
rect -1510 -88 -1498 88
rect -1560 -100 -1498 -88
rect -1442 88 -1380 100
rect -1442 -88 -1430 88
rect -1396 -88 -1380 88
rect -1442 -100 -1380 -88
rect -1350 88 -1288 100
rect -1350 -88 -1334 88
rect -1300 -88 -1288 88
rect -1350 -100 -1288 -88
rect -1232 88 -1170 100
rect -1232 -88 -1220 88
rect -1186 -88 -1170 88
rect -1232 -100 -1170 -88
rect -1140 88 -1078 100
rect -1140 -88 -1124 88
rect -1090 -88 -1078 88
rect -1140 -100 -1078 -88
rect -1022 88 -960 100
rect -1022 -88 -1010 88
rect -976 -88 -960 88
rect -1022 -100 -960 -88
rect -930 88 -868 100
rect -930 -88 -914 88
rect -880 -88 -868 88
rect -930 -100 -868 -88
rect -812 88 -750 100
rect -812 -88 -800 88
rect -766 -88 -750 88
rect -812 -100 -750 -88
rect -720 88 -658 100
rect -720 -88 -704 88
rect -670 -88 -658 88
rect -720 -100 -658 -88
rect -602 88 -540 100
rect -602 -88 -590 88
rect -556 -88 -540 88
rect -602 -100 -540 -88
rect -510 88 -448 100
rect -510 -88 -494 88
rect -460 -88 -448 88
rect -510 -100 -448 -88
rect -392 88 -330 100
rect -392 -88 -380 88
rect -346 -88 -330 88
rect -392 -100 -330 -88
rect -300 88 -238 100
rect -300 -88 -284 88
rect -250 -88 -238 88
rect -300 -100 -238 -88
rect -182 88 -120 100
rect -182 -88 -170 88
rect -136 -88 -120 88
rect -182 -100 -120 -88
rect -90 88 -28 100
rect -90 -88 -74 88
rect -40 -88 -28 88
rect -90 -100 -28 -88
rect 28 88 90 100
rect 28 -88 40 88
rect 74 -88 90 88
rect 28 -100 90 -88
rect 120 88 182 100
rect 120 -88 136 88
rect 170 -88 182 88
rect 120 -100 182 -88
rect 238 88 300 100
rect 238 -88 250 88
rect 284 -88 300 88
rect 238 -100 300 -88
rect 330 88 392 100
rect 330 -88 346 88
rect 380 -88 392 88
rect 330 -100 392 -88
rect 448 88 510 100
rect 448 -88 460 88
rect 494 -88 510 88
rect 448 -100 510 -88
rect 540 88 602 100
rect 540 -88 556 88
rect 590 -88 602 88
rect 540 -100 602 -88
rect 658 88 720 100
rect 658 -88 670 88
rect 704 -88 720 88
rect 658 -100 720 -88
rect 750 88 812 100
rect 750 -88 766 88
rect 800 -88 812 88
rect 750 -100 812 -88
rect 868 88 930 100
rect 868 -88 880 88
rect 914 -88 930 88
rect 868 -100 930 -88
rect 960 88 1022 100
rect 960 -88 976 88
rect 1010 -88 1022 88
rect 960 -100 1022 -88
rect 1078 88 1140 100
rect 1078 -88 1090 88
rect 1124 -88 1140 88
rect 1078 -100 1140 -88
rect 1170 88 1232 100
rect 1170 -88 1186 88
rect 1220 -88 1232 88
rect 1170 -100 1232 -88
rect 1288 88 1350 100
rect 1288 -88 1300 88
rect 1334 -88 1350 88
rect 1288 -100 1350 -88
rect 1380 88 1442 100
rect 1380 -88 1396 88
rect 1430 -88 1442 88
rect 1380 -100 1442 -88
rect 1498 88 1560 100
rect 1498 -88 1510 88
rect 1544 -88 1560 88
rect 1498 -100 1560 -88
rect 1590 88 1652 100
rect 1590 -88 1606 88
rect 1640 -88 1652 88
rect 1590 -100 1652 -88
rect 1708 88 1770 100
rect 1708 -88 1720 88
rect 1754 -88 1770 88
rect 1708 -100 1770 -88
rect 1800 88 1862 100
rect 1800 -88 1816 88
rect 1850 -88 1862 88
rect 1800 -100 1862 -88
rect 1918 88 1980 100
rect 1918 -88 1930 88
rect 1964 -88 1980 88
rect 1918 -100 1980 -88
rect 2010 88 2072 100
rect 2010 -88 2026 88
rect 2060 -88 2072 88
rect 2010 -100 2072 -88
rect 2128 88 2190 100
rect 2128 -88 2140 88
rect 2174 -88 2190 88
rect 2128 -100 2190 -88
rect 2220 88 2282 100
rect 2220 -88 2236 88
rect 2270 -88 2282 88
rect 2220 -100 2282 -88
rect 2338 88 2400 100
rect 2338 -88 2350 88
rect 2384 -88 2400 88
rect 2338 -100 2400 -88
rect 2430 88 2492 100
rect 2430 -88 2446 88
rect 2480 -88 2492 88
rect 2430 -100 2492 -88
rect 2548 88 2610 100
rect 2548 -88 2560 88
rect 2594 -88 2610 88
rect 2548 -100 2610 -88
rect 2640 88 2702 100
rect 2640 -88 2656 88
rect 2690 -88 2702 88
rect 2640 -100 2702 -88
rect 2758 88 2820 100
rect 2758 -88 2770 88
rect 2804 -88 2820 88
rect 2758 -100 2820 -88
rect 2850 88 2912 100
rect 2850 -88 2866 88
rect 2900 -88 2912 88
rect 2850 -100 2912 -88
rect 2968 88 3030 100
rect 2968 -88 2980 88
rect 3014 -88 3030 88
rect 2968 -100 3030 -88
rect 3060 88 3122 100
rect 3060 -88 3076 88
rect 3110 -88 3122 88
rect 3060 -100 3122 -88
rect 3178 88 3240 100
rect 3178 -88 3190 88
rect 3224 -88 3240 88
rect 3178 -100 3240 -88
rect 3270 88 3332 100
rect 3270 -88 3286 88
rect 3320 -88 3332 88
rect 3270 -100 3332 -88
rect 3388 88 3450 100
rect 3388 -88 3400 88
rect 3434 -88 3450 88
rect 3388 -100 3450 -88
rect 3480 88 3542 100
rect 3480 -88 3496 88
rect 3530 -88 3542 88
rect 3480 -100 3542 -88
rect 3598 88 3660 100
rect 3598 -88 3610 88
rect 3644 -88 3660 88
rect 3598 -100 3660 -88
rect 3690 88 3752 100
rect 3690 -88 3706 88
rect 3740 -88 3752 88
rect 3690 -100 3752 -88
rect 3808 88 3870 100
rect 3808 -88 3820 88
rect 3854 -88 3870 88
rect 3808 -100 3870 -88
rect 3900 88 3962 100
rect 3900 -88 3916 88
rect 3950 -88 3962 88
rect 3900 -100 3962 -88
rect 4018 88 4080 100
rect 4018 -88 4030 88
rect 4064 -88 4080 88
rect 4018 -100 4080 -88
rect 4110 88 4172 100
rect 4110 -88 4126 88
rect 4160 -88 4172 88
rect 4110 -100 4172 -88
rect 4228 88 4290 100
rect 4228 -88 4240 88
rect 4274 -88 4290 88
rect 4228 -100 4290 -88
rect 4320 88 4382 100
rect 4320 -88 4336 88
rect 4370 -88 4382 88
rect 4320 -100 4382 -88
rect -4380 -444 -4318 -432
rect -4380 -620 -4368 -444
rect -4334 -620 -4318 -444
rect -4380 -632 -4318 -620
rect -4288 -444 -4226 -432
rect -4288 -620 -4272 -444
rect -4238 -620 -4226 -444
rect -4288 -632 -4226 -620
rect -4170 -444 -4108 -432
rect -4170 -620 -4158 -444
rect -4124 -620 -4108 -444
rect -4170 -632 -4108 -620
rect -4078 -444 -4016 -432
rect -4078 -620 -4062 -444
rect -4028 -620 -4016 -444
rect -4078 -632 -4016 -620
rect -3960 -444 -3898 -432
rect -3960 -620 -3948 -444
rect -3914 -620 -3898 -444
rect -3960 -632 -3898 -620
rect -3868 -444 -3806 -432
rect -3868 -620 -3852 -444
rect -3818 -620 -3806 -444
rect -3868 -632 -3806 -620
rect -3750 -444 -3688 -432
rect -3750 -620 -3738 -444
rect -3704 -620 -3688 -444
rect -3750 -632 -3688 -620
rect -3658 -444 -3596 -432
rect -3658 -620 -3642 -444
rect -3608 -620 -3596 -444
rect -3658 -632 -3596 -620
rect -3540 -444 -3478 -432
rect -3540 -620 -3528 -444
rect -3494 -620 -3478 -444
rect -3540 -632 -3478 -620
rect -3448 -444 -3386 -432
rect -3448 -620 -3432 -444
rect -3398 -620 -3386 -444
rect -3448 -632 -3386 -620
rect -3330 -444 -3268 -432
rect -3330 -620 -3318 -444
rect -3284 -620 -3268 -444
rect -3330 -632 -3268 -620
rect -3238 -444 -3176 -432
rect -3238 -620 -3222 -444
rect -3188 -620 -3176 -444
rect -3238 -632 -3176 -620
rect -3120 -444 -3058 -432
rect -3120 -620 -3108 -444
rect -3074 -620 -3058 -444
rect -3120 -632 -3058 -620
rect -3028 -444 -2966 -432
rect -3028 -620 -3012 -444
rect -2978 -620 -2966 -444
rect -3028 -632 -2966 -620
rect -2910 -444 -2848 -432
rect -2910 -620 -2898 -444
rect -2864 -620 -2848 -444
rect -2910 -632 -2848 -620
rect -2818 -444 -2756 -432
rect -2818 -620 -2802 -444
rect -2768 -620 -2756 -444
rect -2818 -632 -2756 -620
rect -2700 -444 -2638 -432
rect -2700 -620 -2688 -444
rect -2654 -620 -2638 -444
rect -2700 -632 -2638 -620
rect -2608 -444 -2546 -432
rect -2608 -620 -2592 -444
rect -2558 -620 -2546 -444
rect -2608 -632 -2546 -620
rect -2490 -444 -2428 -432
rect -2490 -620 -2478 -444
rect -2444 -620 -2428 -444
rect -2490 -632 -2428 -620
rect -2398 -444 -2336 -432
rect -2398 -620 -2382 -444
rect -2348 -620 -2336 -444
rect -2398 -632 -2336 -620
rect -2280 -444 -2218 -432
rect -2280 -620 -2268 -444
rect -2234 -620 -2218 -444
rect -2280 -632 -2218 -620
rect -2188 -444 -2126 -432
rect -2188 -620 -2172 -444
rect -2138 -620 -2126 -444
rect -2188 -632 -2126 -620
rect -2070 -444 -2008 -432
rect -2070 -620 -2058 -444
rect -2024 -620 -2008 -444
rect -2070 -632 -2008 -620
rect -1978 -444 -1916 -432
rect -1978 -620 -1962 -444
rect -1928 -620 -1916 -444
rect -1978 -632 -1916 -620
rect -1860 -444 -1798 -432
rect -1860 -620 -1848 -444
rect -1814 -620 -1798 -444
rect -1860 -632 -1798 -620
rect -1768 -444 -1706 -432
rect -1768 -620 -1752 -444
rect -1718 -620 -1706 -444
rect -1768 -632 -1706 -620
rect -1650 -444 -1588 -432
rect -1650 -620 -1638 -444
rect -1604 -620 -1588 -444
rect -1650 -632 -1588 -620
rect -1558 -444 -1496 -432
rect -1558 -620 -1542 -444
rect -1508 -620 -1496 -444
rect -1558 -632 -1496 -620
rect -1440 -444 -1378 -432
rect -1440 -620 -1428 -444
rect -1394 -620 -1378 -444
rect -1440 -632 -1378 -620
rect -1348 -444 -1286 -432
rect -1348 -620 -1332 -444
rect -1298 -620 -1286 -444
rect -1348 -632 -1286 -620
rect -1230 -444 -1168 -432
rect -1230 -620 -1218 -444
rect -1184 -620 -1168 -444
rect -1230 -632 -1168 -620
rect -1138 -444 -1076 -432
rect -1138 -620 -1122 -444
rect -1088 -620 -1076 -444
rect -1138 -632 -1076 -620
rect -1020 -444 -958 -432
rect -1020 -620 -1008 -444
rect -974 -620 -958 -444
rect -1020 -632 -958 -620
rect -928 -444 -866 -432
rect -928 -620 -912 -444
rect -878 -620 -866 -444
rect -928 -632 -866 -620
rect -810 -444 -748 -432
rect -810 -620 -798 -444
rect -764 -620 -748 -444
rect -810 -632 -748 -620
rect -718 -444 -656 -432
rect -718 -620 -702 -444
rect -668 -620 -656 -444
rect -718 -632 -656 -620
rect -600 -444 -538 -432
rect -600 -620 -588 -444
rect -554 -620 -538 -444
rect -600 -632 -538 -620
rect -508 -444 -446 -432
rect -508 -620 -492 -444
rect -458 -620 -446 -444
rect -508 -632 -446 -620
rect -390 -444 -328 -432
rect -390 -620 -378 -444
rect -344 -620 -328 -444
rect -390 -632 -328 -620
rect -298 -444 -236 -432
rect -298 -620 -282 -444
rect -248 -620 -236 -444
rect -298 -632 -236 -620
rect -180 -444 -118 -432
rect -180 -620 -168 -444
rect -134 -620 -118 -444
rect -180 -632 -118 -620
rect -88 -444 -26 -432
rect -88 -620 -72 -444
rect -38 -620 -26 -444
rect -88 -632 -26 -620
rect 30 -444 92 -432
rect 30 -620 42 -444
rect 76 -620 92 -444
rect 30 -632 92 -620
rect 122 -444 184 -432
rect 122 -620 138 -444
rect 172 -620 184 -444
rect 122 -632 184 -620
rect 240 -444 302 -432
rect 240 -620 252 -444
rect 286 -620 302 -444
rect 240 -632 302 -620
rect 332 -444 394 -432
rect 332 -620 348 -444
rect 382 -620 394 -444
rect 332 -632 394 -620
rect 450 -444 512 -432
rect 450 -620 462 -444
rect 496 -620 512 -444
rect 450 -632 512 -620
rect 542 -444 604 -432
rect 542 -620 558 -444
rect 592 -620 604 -444
rect 542 -632 604 -620
rect 660 -444 722 -432
rect 660 -620 672 -444
rect 706 -620 722 -444
rect 660 -632 722 -620
rect 752 -444 814 -432
rect 752 -620 768 -444
rect 802 -620 814 -444
rect 752 -632 814 -620
rect 870 -444 932 -432
rect 870 -620 882 -444
rect 916 -620 932 -444
rect 870 -632 932 -620
rect 962 -444 1024 -432
rect 962 -620 978 -444
rect 1012 -620 1024 -444
rect 962 -632 1024 -620
rect 1080 -444 1142 -432
rect 1080 -620 1092 -444
rect 1126 -620 1142 -444
rect 1080 -632 1142 -620
rect 1172 -444 1234 -432
rect 1172 -620 1188 -444
rect 1222 -620 1234 -444
rect 1172 -632 1234 -620
rect 1290 -444 1352 -432
rect 1290 -620 1302 -444
rect 1336 -620 1352 -444
rect 1290 -632 1352 -620
rect 1382 -444 1444 -432
rect 1382 -620 1398 -444
rect 1432 -620 1444 -444
rect 1382 -632 1444 -620
rect 1500 -444 1562 -432
rect 1500 -620 1512 -444
rect 1546 -620 1562 -444
rect 1500 -632 1562 -620
rect 1592 -444 1654 -432
rect 1592 -620 1608 -444
rect 1642 -620 1654 -444
rect 1592 -632 1654 -620
rect 1710 -444 1772 -432
rect 1710 -620 1722 -444
rect 1756 -620 1772 -444
rect 1710 -632 1772 -620
rect 1802 -444 1864 -432
rect 1802 -620 1818 -444
rect 1852 -620 1864 -444
rect 1802 -632 1864 -620
rect 1920 -444 1982 -432
rect 1920 -620 1932 -444
rect 1966 -620 1982 -444
rect 1920 -632 1982 -620
rect 2012 -444 2074 -432
rect 2012 -620 2028 -444
rect 2062 -620 2074 -444
rect 2012 -632 2074 -620
rect 2130 -444 2192 -432
rect 2130 -620 2142 -444
rect 2176 -620 2192 -444
rect 2130 -632 2192 -620
rect 2222 -444 2284 -432
rect 2222 -620 2238 -444
rect 2272 -620 2284 -444
rect 2222 -632 2284 -620
rect 2340 -444 2402 -432
rect 2340 -620 2352 -444
rect 2386 -620 2402 -444
rect 2340 -632 2402 -620
rect 2432 -444 2494 -432
rect 2432 -620 2448 -444
rect 2482 -620 2494 -444
rect 2432 -632 2494 -620
rect 2550 -444 2612 -432
rect 2550 -620 2562 -444
rect 2596 -620 2612 -444
rect 2550 -632 2612 -620
rect 2642 -444 2704 -432
rect 2642 -620 2658 -444
rect 2692 -620 2704 -444
rect 2642 -632 2704 -620
rect 2760 -444 2822 -432
rect 2760 -620 2772 -444
rect 2806 -620 2822 -444
rect 2760 -632 2822 -620
rect 2852 -444 2914 -432
rect 2852 -620 2868 -444
rect 2902 -620 2914 -444
rect 2852 -632 2914 -620
rect 2970 -444 3032 -432
rect 2970 -620 2982 -444
rect 3016 -620 3032 -444
rect 2970 -632 3032 -620
rect 3062 -444 3124 -432
rect 3062 -620 3078 -444
rect 3112 -620 3124 -444
rect 3062 -632 3124 -620
rect 3180 -444 3242 -432
rect 3180 -620 3192 -444
rect 3226 -620 3242 -444
rect 3180 -632 3242 -620
rect 3272 -444 3334 -432
rect 3272 -620 3288 -444
rect 3322 -620 3334 -444
rect 3272 -632 3334 -620
rect 3390 -444 3452 -432
rect 3390 -620 3402 -444
rect 3436 -620 3452 -444
rect 3390 -632 3452 -620
rect 3482 -444 3544 -432
rect 3482 -620 3498 -444
rect 3532 -620 3544 -444
rect 3482 -632 3544 -620
rect 3600 -444 3662 -432
rect 3600 -620 3612 -444
rect 3646 -620 3662 -444
rect 3600 -632 3662 -620
rect 3692 -444 3754 -432
rect 3692 -620 3708 -444
rect 3742 -620 3754 -444
rect 3692 -632 3754 -620
rect 3810 -444 3872 -432
rect 3810 -620 3822 -444
rect 3856 -620 3872 -444
rect 3810 -632 3872 -620
rect 3902 -444 3964 -432
rect 3902 -620 3918 -444
rect 3952 -620 3964 -444
rect 3902 -632 3964 -620
rect 4020 -444 4082 -432
rect 4020 -620 4032 -444
rect 4066 -620 4082 -444
rect 4020 -632 4082 -620
rect 4112 -444 4174 -432
rect 4112 -620 4128 -444
rect 4162 -620 4174 -444
rect 4112 -632 4174 -620
rect 4230 -444 4292 -432
rect 4230 -620 4242 -444
rect 4276 -620 4292 -444
rect 4230 -632 4292 -620
rect 4322 -444 4384 -432
rect 4322 -620 4338 -444
rect 4372 -620 4384 -444
rect 4322 -632 4384 -620
<< pdiffc >>
rect -4370 -88 -4336 88
rect -4274 -88 -4240 88
rect -4160 -88 -4126 88
rect -4064 -88 -4030 88
rect -3950 -88 -3916 88
rect -3854 -88 -3820 88
rect -3740 -88 -3706 88
rect -3644 -88 -3610 88
rect -3530 -88 -3496 88
rect -3434 -88 -3400 88
rect -3320 -88 -3286 88
rect -3224 -88 -3190 88
rect -3110 -88 -3076 88
rect -3014 -88 -2980 88
rect -2900 -88 -2866 88
rect -2804 -88 -2770 88
rect -2690 -88 -2656 88
rect -2594 -88 -2560 88
rect -2480 -88 -2446 88
rect -2384 -88 -2350 88
rect -2270 -88 -2236 88
rect -2174 -88 -2140 88
rect -2060 -88 -2026 88
rect -1964 -88 -1930 88
rect -1850 -88 -1816 88
rect -1754 -88 -1720 88
rect -1640 -88 -1606 88
rect -1544 -88 -1510 88
rect -1430 -88 -1396 88
rect -1334 -88 -1300 88
rect -1220 -88 -1186 88
rect -1124 -88 -1090 88
rect -1010 -88 -976 88
rect -914 -88 -880 88
rect -800 -88 -766 88
rect -704 -88 -670 88
rect -590 -88 -556 88
rect -494 -88 -460 88
rect -380 -88 -346 88
rect -284 -88 -250 88
rect -170 -88 -136 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 136 -88 170 88
rect 250 -88 284 88
rect 346 -88 380 88
rect 460 -88 494 88
rect 556 -88 590 88
rect 670 -88 704 88
rect 766 -88 800 88
rect 880 -88 914 88
rect 976 -88 1010 88
rect 1090 -88 1124 88
rect 1186 -88 1220 88
rect 1300 -88 1334 88
rect 1396 -88 1430 88
rect 1510 -88 1544 88
rect 1606 -88 1640 88
rect 1720 -88 1754 88
rect 1816 -88 1850 88
rect 1930 -88 1964 88
rect 2026 -88 2060 88
rect 2140 -88 2174 88
rect 2236 -88 2270 88
rect 2350 -88 2384 88
rect 2446 -88 2480 88
rect 2560 -88 2594 88
rect 2656 -88 2690 88
rect 2770 -88 2804 88
rect 2866 -88 2900 88
rect 2980 -88 3014 88
rect 3076 -88 3110 88
rect 3190 -88 3224 88
rect 3286 -88 3320 88
rect 3400 -88 3434 88
rect 3496 -88 3530 88
rect 3610 -88 3644 88
rect 3706 -88 3740 88
rect 3820 -88 3854 88
rect 3916 -88 3950 88
rect 4030 -88 4064 88
rect 4126 -88 4160 88
rect 4240 -88 4274 88
rect 4336 -88 4370 88
rect -4368 -620 -4334 -444
rect -4272 -620 -4238 -444
rect -4158 -620 -4124 -444
rect -4062 -620 -4028 -444
rect -3948 -620 -3914 -444
rect -3852 -620 -3818 -444
rect -3738 -620 -3704 -444
rect -3642 -620 -3608 -444
rect -3528 -620 -3494 -444
rect -3432 -620 -3398 -444
rect -3318 -620 -3284 -444
rect -3222 -620 -3188 -444
rect -3108 -620 -3074 -444
rect -3012 -620 -2978 -444
rect -2898 -620 -2864 -444
rect -2802 -620 -2768 -444
rect -2688 -620 -2654 -444
rect -2592 -620 -2558 -444
rect -2478 -620 -2444 -444
rect -2382 -620 -2348 -444
rect -2268 -620 -2234 -444
rect -2172 -620 -2138 -444
rect -2058 -620 -2024 -444
rect -1962 -620 -1928 -444
rect -1848 -620 -1814 -444
rect -1752 -620 -1718 -444
rect -1638 -620 -1604 -444
rect -1542 -620 -1508 -444
rect -1428 -620 -1394 -444
rect -1332 -620 -1298 -444
rect -1218 -620 -1184 -444
rect -1122 -620 -1088 -444
rect -1008 -620 -974 -444
rect -912 -620 -878 -444
rect -798 -620 -764 -444
rect -702 -620 -668 -444
rect -588 -620 -554 -444
rect -492 -620 -458 -444
rect -378 -620 -344 -444
rect -282 -620 -248 -444
rect -168 -620 -134 -444
rect -72 -620 -38 -444
rect 42 -620 76 -444
rect 138 -620 172 -444
rect 252 -620 286 -444
rect 348 -620 382 -444
rect 462 -620 496 -444
rect 558 -620 592 -444
rect 672 -620 706 -444
rect 768 -620 802 -444
rect 882 -620 916 -444
rect 978 -620 1012 -444
rect 1092 -620 1126 -444
rect 1188 -620 1222 -444
rect 1302 -620 1336 -444
rect 1398 -620 1432 -444
rect 1512 -620 1546 -444
rect 1608 -620 1642 -444
rect 1722 -620 1756 -444
rect 1818 -620 1852 -444
rect 1932 -620 1966 -444
rect 2028 -620 2062 -444
rect 2142 -620 2176 -444
rect 2238 -620 2272 -444
rect 2352 -620 2386 -444
rect 2448 -620 2482 -444
rect 2562 -620 2596 -444
rect 2658 -620 2692 -444
rect 2772 -620 2806 -444
rect 2868 -620 2902 -444
rect 2982 -620 3016 -444
rect 3078 -620 3112 -444
rect 3192 -620 3226 -444
rect 3288 -620 3322 -444
rect 3402 -620 3436 -444
rect 3498 -620 3532 -444
rect 3612 -620 3646 -444
rect 3708 -620 3742 -444
rect 3822 -620 3856 -444
rect 3918 -620 3952 -444
rect 4032 -620 4066 -444
rect 4128 -620 4162 -444
rect 4242 -620 4276 -444
rect 4338 -620 4372 -444
<< nsubdiff >>
rect -4484 249 -4388 283
rect 4388 249 4484 283
rect -4484 187 -4450 249
rect 4450 187 4484 249
rect -4484 -345 -4450 -187
rect 4450 -345 4484 -187
rect -4484 -781 -4450 -719
rect 4450 -781 4484 -719
rect -4484 -815 -4388 -781
rect 4388 -815 4484 -781
<< nsubdiffcont >>
rect -4388 249 4388 283
rect -4484 -187 -4450 187
rect 4450 -187 4484 187
rect -4484 -719 -4450 -345
rect 4450 -719 4484 -345
rect -4388 -815 4388 -781
<< poly >>
rect -4128 181 -4062 197
rect -4128 147 -4112 181
rect -4078 147 -4062 181
rect -4128 131 -4062 147
rect -3708 181 -3642 197
rect -3708 147 -3692 181
rect -3658 147 -3642 181
rect -3708 131 -3642 147
rect -3288 181 -3222 197
rect -3288 147 -3272 181
rect -3238 147 -3222 181
rect -3288 131 -3222 147
rect -2868 181 -2802 197
rect -2868 147 -2852 181
rect -2818 147 -2802 181
rect -2868 131 -2802 147
rect -2448 181 -2382 197
rect -2448 147 -2432 181
rect -2398 147 -2382 181
rect -2448 131 -2382 147
rect -2028 181 -1962 197
rect -2028 147 -2012 181
rect -1978 147 -1962 181
rect -2028 131 -1962 147
rect -1608 181 -1542 197
rect -1608 147 -1592 181
rect -1558 147 -1542 181
rect -1608 131 -1542 147
rect -1188 181 -1122 197
rect -1188 147 -1172 181
rect -1138 147 -1122 181
rect -1188 131 -1122 147
rect -768 181 -702 197
rect -768 147 -752 181
rect -718 147 -702 181
rect -768 131 -702 147
rect -348 181 -282 197
rect -348 147 -332 181
rect -298 147 -282 181
rect -348 131 -282 147
rect 72 181 138 197
rect 72 147 88 181
rect 122 147 138 181
rect 72 131 138 147
rect 492 181 558 197
rect 492 147 508 181
rect 542 147 558 181
rect 492 131 558 147
rect 912 181 978 197
rect 912 147 928 181
rect 962 147 978 181
rect 912 131 978 147
rect 1332 181 1398 197
rect 1332 147 1348 181
rect 1382 147 1398 181
rect 1332 131 1398 147
rect 1752 181 1818 197
rect 1752 147 1768 181
rect 1802 147 1818 181
rect 1752 131 1818 147
rect 2172 181 2238 197
rect 2172 147 2188 181
rect 2222 147 2238 181
rect 2172 131 2238 147
rect 2592 181 2658 197
rect 2592 147 2608 181
rect 2642 147 2658 181
rect 2592 131 2658 147
rect 3012 181 3078 197
rect 3012 147 3028 181
rect 3062 147 3078 181
rect 3012 131 3078 147
rect 3432 181 3498 197
rect 3432 147 3448 181
rect 3482 147 3498 181
rect 3432 131 3498 147
rect 3852 181 3918 197
rect 3852 147 3868 181
rect 3902 147 3918 181
rect 3852 131 3918 147
rect 4272 181 4338 197
rect 4272 147 4288 181
rect 4322 147 4338 181
rect 4272 131 4338 147
rect -4320 100 -4290 126
rect -4110 100 -4080 131
rect -3900 100 -3870 126
rect -3690 100 -3660 131
rect -3480 100 -3450 126
rect -3270 100 -3240 131
rect -3060 100 -3030 126
rect -2850 100 -2820 131
rect -2640 100 -2610 126
rect -2430 100 -2400 131
rect -2220 100 -2190 126
rect -2010 100 -1980 131
rect -1800 100 -1770 126
rect -1590 100 -1560 131
rect -1380 100 -1350 126
rect -1170 100 -1140 131
rect -960 100 -930 126
rect -750 100 -720 131
rect -540 100 -510 126
rect -330 100 -300 131
rect -120 100 -90 126
rect 90 100 120 131
rect 300 100 330 126
rect 510 100 540 131
rect 720 100 750 126
rect 930 100 960 131
rect 1140 100 1170 126
rect 1350 100 1380 131
rect 1560 100 1590 126
rect 1770 100 1800 131
rect 1980 100 2010 126
rect 2190 100 2220 131
rect 2400 100 2430 126
rect 2610 100 2640 131
rect 2820 100 2850 126
rect 3030 100 3060 131
rect 3240 100 3270 126
rect 3450 100 3480 131
rect 3660 100 3690 126
rect 3870 100 3900 131
rect 4080 100 4110 126
rect 4290 100 4320 131
rect -4320 -131 -4290 -100
rect -4110 -126 -4080 -100
rect -3900 -131 -3870 -100
rect -3690 -126 -3660 -100
rect -3480 -131 -3450 -100
rect -3270 -126 -3240 -100
rect -3060 -131 -3030 -100
rect -2850 -126 -2820 -100
rect -2640 -131 -2610 -100
rect -2430 -126 -2400 -100
rect -2220 -131 -2190 -100
rect -2010 -126 -1980 -100
rect -1800 -131 -1770 -100
rect -1590 -126 -1560 -100
rect -1380 -131 -1350 -100
rect -1170 -126 -1140 -100
rect -960 -131 -930 -100
rect -750 -126 -720 -100
rect -540 -131 -510 -100
rect -330 -126 -300 -100
rect -120 -131 -90 -100
rect 90 -126 120 -100
rect 300 -131 330 -100
rect 510 -126 540 -100
rect 720 -131 750 -100
rect 930 -126 960 -100
rect 1140 -131 1170 -100
rect 1350 -126 1380 -100
rect 1560 -131 1590 -100
rect 1770 -126 1800 -100
rect 1980 -131 2010 -100
rect 2190 -126 2220 -100
rect 2400 -131 2430 -100
rect 2610 -126 2640 -100
rect 2820 -131 2850 -100
rect 3030 -126 3060 -100
rect 3240 -131 3270 -100
rect 3450 -126 3480 -100
rect 3660 -131 3690 -100
rect 3870 -126 3900 -100
rect 4080 -131 4110 -100
rect 4290 -126 4320 -100
rect -4338 -147 -4272 -131
rect -4338 -181 -4322 -147
rect -4288 -181 -4272 -147
rect -4338 -197 -4272 -181
rect -3918 -147 -3852 -131
rect -3918 -181 -3902 -147
rect -3868 -181 -3852 -147
rect -3918 -197 -3852 -181
rect -3498 -147 -3432 -131
rect -3498 -181 -3482 -147
rect -3448 -181 -3432 -147
rect -3498 -197 -3432 -181
rect -3078 -147 -3012 -131
rect -3078 -181 -3062 -147
rect -3028 -181 -3012 -147
rect -3078 -197 -3012 -181
rect -2658 -147 -2592 -131
rect -2658 -181 -2642 -147
rect -2608 -181 -2592 -147
rect -2658 -197 -2592 -181
rect -2238 -147 -2172 -131
rect -2238 -181 -2222 -147
rect -2188 -181 -2172 -147
rect -2238 -197 -2172 -181
rect -1818 -147 -1752 -131
rect -1818 -181 -1802 -147
rect -1768 -181 -1752 -147
rect -1818 -197 -1752 -181
rect -1398 -147 -1332 -131
rect -1398 -181 -1382 -147
rect -1348 -181 -1332 -147
rect -1398 -197 -1332 -181
rect -978 -147 -912 -131
rect -978 -181 -962 -147
rect -928 -181 -912 -147
rect -978 -197 -912 -181
rect -558 -147 -492 -131
rect -558 -181 -542 -147
rect -508 -181 -492 -147
rect -558 -197 -492 -181
rect -138 -147 -72 -131
rect -138 -181 -122 -147
rect -88 -181 -72 -147
rect -138 -197 -72 -181
rect 282 -147 348 -131
rect 282 -181 298 -147
rect 332 -181 348 -147
rect 282 -197 348 -181
rect 702 -147 768 -131
rect 702 -181 718 -147
rect 752 -181 768 -147
rect 702 -197 768 -181
rect 1122 -147 1188 -131
rect 1122 -181 1138 -147
rect 1172 -181 1188 -147
rect 1122 -197 1188 -181
rect 1542 -147 1608 -131
rect 1542 -181 1558 -147
rect 1592 -181 1608 -147
rect 1542 -197 1608 -181
rect 1962 -147 2028 -131
rect 1962 -181 1978 -147
rect 2012 -181 2028 -147
rect 1962 -197 2028 -181
rect 2382 -147 2448 -131
rect 2382 -181 2398 -147
rect 2432 -181 2448 -147
rect 2382 -197 2448 -181
rect 2802 -147 2868 -131
rect 2802 -181 2818 -147
rect 2852 -181 2868 -147
rect 2802 -197 2868 -181
rect 3222 -147 3288 -131
rect 3222 -181 3238 -147
rect 3272 -181 3288 -147
rect 3222 -197 3288 -181
rect 3642 -147 3708 -131
rect 3642 -181 3658 -147
rect 3692 -181 3708 -147
rect 3642 -197 3708 -181
rect 4062 -147 4128 -131
rect 4062 -181 4078 -147
rect 4112 -181 4128 -147
rect 4062 -197 4128 -181
rect -4126 -351 -4060 -335
rect -4126 -385 -4110 -351
rect -4076 -385 -4060 -351
rect -4126 -401 -4060 -385
rect -3706 -351 -3640 -335
rect -3706 -385 -3690 -351
rect -3656 -385 -3640 -351
rect -3706 -401 -3640 -385
rect -3286 -351 -3220 -335
rect -3286 -385 -3270 -351
rect -3236 -385 -3220 -351
rect -3286 -401 -3220 -385
rect -2866 -351 -2800 -335
rect -2866 -385 -2850 -351
rect -2816 -385 -2800 -351
rect -2866 -401 -2800 -385
rect -2446 -351 -2380 -335
rect -2446 -385 -2430 -351
rect -2396 -385 -2380 -351
rect -2446 -401 -2380 -385
rect -2026 -351 -1960 -335
rect -2026 -385 -2010 -351
rect -1976 -385 -1960 -351
rect -2026 -401 -1960 -385
rect -1606 -351 -1540 -335
rect -1606 -385 -1590 -351
rect -1556 -385 -1540 -351
rect -1606 -401 -1540 -385
rect -1186 -351 -1120 -335
rect -1186 -385 -1170 -351
rect -1136 -385 -1120 -351
rect -1186 -401 -1120 -385
rect -766 -351 -700 -335
rect -766 -385 -750 -351
rect -716 -385 -700 -351
rect -766 -401 -700 -385
rect -346 -351 -280 -335
rect -346 -385 -330 -351
rect -296 -385 -280 -351
rect -346 -401 -280 -385
rect 74 -351 140 -335
rect 74 -385 90 -351
rect 124 -385 140 -351
rect 74 -401 140 -385
rect 494 -351 560 -335
rect 494 -385 510 -351
rect 544 -385 560 -351
rect 494 -401 560 -385
rect 914 -351 980 -335
rect 914 -385 930 -351
rect 964 -385 980 -351
rect 914 -401 980 -385
rect 1334 -351 1400 -335
rect 1334 -385 1350 -351
rect 1384 -385 1400 -351
rect 1334 -401 1400 -385
rect 1754 -351 1820 -335
rect 1754 -385 1770 -351
rect 1804 -385 1820 -351
rect 1754 -401 1820 -385
rect 2174 -351 2240 -335
rect 2174 -385 2190 -351
rect 2224 -385 2240 -351
rect 2174 -401 2240 -385
rect 2594 -351 2660 -335
rect 2594 -385 2610 -351
rect 2644 -385 2660 -351
rect 2594 -401 2660 -385
rect 3014 -351 3080 -335
rect 3014 -385 3030 -351
rect 3064 -385 3080 -351
rect 3014 -401 3080 -385
rect 3434 -351 3500 -335
rect 3434 -385 3450 -351
rect 3484 -385 3500 -351
rect 3434 -401 3500 -385
rect 3854 -351 3920 -335
rect 3854 -385 3870 -351
rect 3904 -385 3920 -351
rect 3854 -401 3920 -385
rect 4274 -351 4340 -335
rect 4274 -385 4290 -351
rect 4324 -385 4340 -351
rect 4274 -401 4340 -385
rect -4318 -432 -4288 -406
rect -4108 -432 -4078 -401
rect -3898 -432 -3868 -406
rect -3688 -432 -3658 -401
rect -3478 -432 -3448 -406
rect -3268 -432 -3238 -401
rect -3058 -432 -3028 -406
rect -2848 -432 -2818 -401
rect -2638 -432 -2608 -406
rect -2428 -432 -2398 -401
rect -2218 -432 -2188 -406
rect -2008 -432 -1978 -401
rect -1798 -432 -1768 -406
rect -1588 -432 -1558 -401
rect -1378 -432 -1348 -406
rect -1168 -432 -1138 -401
rect -958 -432 -928 -406
rect -748 -432 -718 -401
rect -538 -432 -508 -406
rect -328 -432 -298 -401
rect -118 -432 -88 -406
rect 92 -432 122 -401
rect 302 -432 332 -406
rect 512 -432 542 -401
rect 722 -432 752 -406
rect 932 -432 962 -401
rect 1142 -432 1172 -406
rect 1352 -432 1382 -401
rect 1562 -432 1592 -406
rect 1772 -432 1802 -401
rect 1982 -432 2012 -406
rect 2192 -432 2222 -401
rect 2402 -432 2432 -406
rect 2612 -432 2642 -401
rect 2822 -432 2852 -406
rect 3032 -432 3062 -401
rect 3242 -432 3272 -406
rect 3452 -432 3482 -401
rect 3662 -432 3692 -406
rect 3872 -432 3902 -401
rect 4082 -432 4112 -406
rect 4292 -432 4322 -401
rect -4318 -663 -4288 -632
rect -4108 -658 -4078 -632
rect -3898 -663 -3868 -632
rect -3688 -658 -3658 -632
rect -3478 -663 -3448 -632
rect -3268 -658 -3238 -632
rect -3058 -663 -3028 -632
rect -2848 -658 -2818 -632
rect -2638 -663 -2608 -632
rect -2428 -658 -2398 -632
rect -2218 -663 -2188 -632
rect -2008 -658 -1978 -632
rect -1798 -663 -1768 -632
rect -1588 -658 -1558 -632
rect -1378 -663 -1348 -632
rect -1168 -658 -1138 -632
rect -958 -663 -928 -632
rect -748 -658 -718 -632
rect -538 -663 -508 -632
rect -328 -658 -298 -632
rect -118 -663 -88 -632
rect 92 -658 122 -632
rect 302 -663 332 -632
rect 512 -658 542 -632
rect 722 -663 752 -632
rect 932 -658 962 -632
rect 1142 -663 1172 -632
rect 1352 -658 1382 -632
rect 1562 -663 1592 -632
rect 1772 -658 1802 -632
rect 1982 -663 2012 -632
rect 2192 -658 2222 -632
rect 2402 -663 2432 -632
rect 2612 -658 2642 -632
rect 2822 -663 2852 -632
rect 3032 -658 3062 -632
rect 3242 -663 3272 -632
rect 3452 -658 3482 -632
rect 3662 -663 3692 -632
rect 3872 -658 3902 -632
rect 4082 -663 4112 -632
rect 4292 -658 4322 -632
rect -4336 -679 -4270 -663
rect -4336 -713 -4320 -679
rect -4286 -713 -4270 -679
rect -4336 -729 -4270 -713
rect -3916 -679 -3850 -663
rect -3916 -713 -3900 -679
rect -3866 -713 -3850 -679
rect -3916 -729 -3850 -713
rect -3496 -679 -3430 -663
rect -3496 -713 -3480 -679
rect -3446 -713 -3430 -679
rect -3496 -729 -3430 -713
rect -3076 -679 -3010 -663
rect -3076 -713 -3060 -679
rect -3026 -713 -3010 -679
rect -3076 -729 -3010 -713
rect -2656 -679 -2590 -663
rect -2656 -713 -2640 -679
rect -2606 -713 -2590 -679
rect -2656 -729 -2590 -713
rect -2236 -679 -2170 -663
rect -2236 -713 -2220 -679
rect -2186 -713 -2170 -679
rect -2236 -729 -2170 -713
rect -1816 -679 -1750 -663
rect -1816 -713 -1800 -679
rect -1766 -713 -1750 -679
rect -1816 -729 -1750 -713
rect -1396 -679 -1330 -663
rect -1396 -713 -1380 -679
rect -1346 -713 -1330 -679
rect -1396 -729 -1330 -713
rect -976 -679 -910 -663
rect -976 -713 -960 -679
rect -926 -713 -910 -679
rect -976 -729 -910 -713
rect -556 -679 -490 -663
rect -556 -713 -540 -679
rect -506 -713 -490 -679
rect -556 -729 -490 -713
rect -136 -679 -70 -663
rect -136 -713 -120 -679
rect -86 -713 -70 -679
rect -136 -729 -70 -713
rect 284 -679 350 -663
rect 284 -713 300 -679
rect 334 -713 350 -679
rect 284 -729 350 -713
rect 704 -679 770 -663
rect 704 -713 720 -679
rect 754 -713 770 -679
rect 704 -729 770 -713
rect 1124 -679 1190 -663
rect 1124 -713 1140 -679
rect 1174 -713 1190 -679
rect 1124 -729 1190 -713
rect 1544 -679 1610 -663
rect 1544 -713 1560 -679
rect 1594 -713 1610 -679
rect 1544 -729 1610 -713
rect 1964 -679 2030 -663
rect 1964 -713 1980 -679
rect 2014 -713 2030 -679
rect 1964 -729 2030 -713
rect 2384 -679 2450 -663
rect 2384 -713 2400 -679
rect 2434 -713 2450 -679
rect 2384 -729 2450 -713
rect 2804 -679 2870 -663
rect 2804 -713 2820 -679
rect 2854 -713 2870 -679
rect 2804 -729 2870 -713
rect 3224 -679 3290 -663
rect 3224 -713 3240 -679
rect 3274 -713 3290 -679
rect 3224 -729 3290 -713
rect 3644 -679 3710 -663
rect 3644 -713 3660 -679
rect 3694 -713 3710 -679
rect 3644 -729 3710 -713
rect 4064 -679 4130 -663
rect 4064 -713 4080 -679
rect 4114 -713 4130 -679
rect 4064 -729 4130 -713
<< polycont >>
rect -4112 147 -4078 181
rect -3692 147 -3658 181
rect -3272 147 -3238 181
rect -2852 147 -2818 181
rect -2432 147 -2398 181
rect -2012 147 -1978 181
rect -1592 147 -1558 181
rect -1172 147 -1138 181
rect -752 147 -718 181
rect -332 147 -298 181
rect 88 147 122 181
rect 508 147 542 181
rect 928 147 962 181
rect 1348 147 1382 181
rect 1768 147 1802 181
rect 2188 147 2222 181
rect 2608 147 2642 181
rect 3028 147 3062 181
rect 3448 147 3482 181
rect 3868 147 3902 181
rect 4288 147 4322 181
rect -4322 -181 -4288 -147
rect -3902 -181 -3868 -147
rect -3482 -181 -3448 -147
rect -3062 -181 -3028 -147
rect -2642 -181 -2608 -147
rect -2222 -181 -2188 -147
rect -1802 -181 -1768 -147
rect -1382 -181 -1348 -147
rect -962 -181 -928 -147
rect -542 -181 -508 -147
rect -122 -181 -88 -147
rect 298 -181 332 -147
rect 718 -181 752 -147
rect 1138 -181 1172 -147
rect 1558 -181 1592 -147
rect 1978 -181 2012 -147
rect 2398 -181 2432 -147
rect 2818 -181 2852 -147
rect 3238 -181 3272 -147
rect 3658 -181 3692 -147
rect 4078 -181 4112 -147
rect -4110 -385 -4076 -351
rect -3690 -385 -3656 -351
rect -3270 -385 -3236 -351
rect -2850 -385 -2816 -351
rect -2430 -385 -2396 -351
rect -2010 -385 -1976 -351
rect -1590 -385 -1556 -351
rect -1170 -385 -1136 -351
rect -750 -385 -716 -351
rect -330 -385 -296 -351
rect 90 -385 124 -351
rect 510 -385 544 -351
rect 930 -385 964 -351
rect 1350 -385 1384 -351
rect 1770 -385 1804 -351
rect 2190 -385 2224 -351
rect 2610 -385 2644 -351
rect 3030 -385 3064 -351
rect 3450 -385 3484 -351
rect 3870 -385 3904 -351
rect 4290 -385 4324 -351
rect -4320 -713 -4286 -679
rect -3900 -713 -3866 -679
rect -3480 -713 -3446 -679
rect -3060 -713 -3026 -679
rect -2640 -713 -2606 -679
rect -2220 -713 -2186 -679
rect -1800 -713 -1766 -679
rect -1380 -713 -1346 -679
rect -960 -713 -926 -679
rect -540 -713 -506 -679
rect -120 -713 -86 -679
rect 300 -713 334 -679
rect 720 -713 754 -679
rect 1140 -713 1174 -679
rect 1560 -713 1594 -679
rect 1980 -713 2014 -679
rect 2400 -713 2434 -679
rect 2820 -713 2854 -679
rect 3240 -713 3274 -679
rect 3660 -713 3694 -679
rect 4080 -713 4114 -679
<< locali >>
rect -4484 249 -4388 283
rect 4388 249 4484 283
rect -4484 187 -4450 249
rect 4450 187 4484 249
rect -4128 147 -4112 181
rect -4078 147 -4062 181
rect -3708 147 -3692 181
rect -3658 147 -3642 181
rect -3288 147 -3272 181
rect -3238 147 -3222 181
rect -2868 147 -2852 181
rect -2818 147 -2802 181
rect -2448 147 -2432 181
rect -2398 147 -2382 181
rect -2028 147 -2012 181
rect -1978 147 -1962 181
rect -1608 147 -1592 181
rect -1558 147 -1542 181
rect -1188 147 -1172 181
rect -1138 147 -1122 181
rect -768 147 -752 181
rect -718 147 -702 181
rect -348 147 -332 181
rect -298 147 -282 181
rect 72 147 88 181
rect 122 147 138 181
rect 492 147 508 181
rect 542 147 558 181
rect 912 147 928 181
rect 962 147 978 181
rect 1332 147 1348 181
rect 1382 147 1398 181
rect 1752 147 1768 181
rect 1802 147 1818 181
rect 2172 147 2188 181
rect 2222 147 2238 181
rect 2592 147 2608 181
rect 2642 147 2658 181
rect 3012 147 3028 181
rect 3062 147 3078 181
rect 3432 147 3448 181
rect 3482 147 3498 181
rect 3852 147 3868 181
rect 3902 147 3918 181
rect 4240 147 4288 181
rect 4322 147 4450 181
rect -4370 88 -4336 104
rect -4370 -147 -4336 -88
rect -4274 88 -4240 104
rect -4274 -147 -4240 -88
rect -4160 88 -4126 104
rect -4160 -104 -4126 -88
rect -4064 88 -4030 104
rect -4064 -104 -4030 -88
rect -3950 88 -3916 104
rect -3950 -104 -3916 -88
rect -3854 88 -3820 104
rect -3854 -104 -3820 -88
rect -3740 88 -3706 104
rect -3740 -104 -3706 -88
rect -3644 88 -3610 104
rect -3644 -104 -3610 -88
rect -3530 88 -3496 104
rect -3530 -104 -3496 -88
rect -3434 88 -3400 104
rect -3434 -104 -3400 -88
rect -3320 88 -3286 104
rect -3320 -104 -3286 -88
rect -3224 88 -3190 104
rect -3224 -104 -3190 -88
rect -3110 88 -3076 104
rect -3110 -104 -3076 -88
rect -3014 88 -2980 104
rect -3014 -104 -2980 -88
rect -2900 88 -2866 104
rect -2900 -104 -2866 -88
rect -2804 88 -2770 104
rect -2804 -104 -2770 -88
rect -2690 88 -2656 104
rect -2690 -104 -2656 -88
rect -2594 88 -2560 104
rect -2594 -104 -2560 -88
rect -2480 88 -2446 104
rect -2480 -104 -2446 -88
rect -2384 88 -2350 104
rect -2384 -104 -2350 -88
rect -2270 88 -2236 104
rect -2270 -104 -2236 -88
rect -2174 88 -2140 104
rect -2174 -104 -2140 -88
rect -2060 88 -2026 104
rect -2060 -104 -2026 -88
rect -1964 88 -1930 104
rect -1964 -104 -1930 -88
rect -1850 88 -1816 104
rect -1850 -104 -1816 -88
rect -1754 88 -1720 104
rect -1754 -104 -1720 -88
rect -1640 88 -1606 104
rect -1640 -104 -1606 -88
rect -1544 88 -1510 104
rect -1544 -104 -1510 -88
rect -1430 88 -1396 104
rect -1430 -104 -1396 -88
rect -1334 88 -1300 104
rect -1334 -104 -1300 -88
rect -1220 88 -1186 104
rect -1220 -104 -1186 -88
rect -1124 88 -1090 104
rect -1124 -104 -1090 -88
rect -1010 88 -976 104
rect -1010 -104 -976 -88
rect -914 88 -880 104
rect -914 -104 -880 -88
rect -800 88 -766 104
rect -800 -104 -766 -88
rect -704 88 -670 104
rect -704 -104 -670 -88
rect -590 88 -556 104
rect -590 -104 -556 -88
rect -494 88 -460 104
rect -494 -104 -460 -88
rect -380 88 -346 104
rect -380 -104 -346 -88
rect -284 88 -250 104
rect -284 -104 -250 -88
rect -170 88 -136 104
rect -170 -104 -136 -88
rect -74 88 -40 104
rect -74 -104 -40 -88
rect 40 88 74 104
rect 40 -104 74 -88
rect 136 88 170 104
rect 136 -104 170 -88
rect 250 88 284 104
rect 250 -104 284 -88
rect 346 88 380 104
rect 346 -104 380 -88
rect 460 88 494 104
rect 460 -104 494 -88
rect 556 88 590 104
rect 556 -104 590 -88
rect 670 88 704 104
rect 670 -104 704 -88
rect 766 88 800 104
rect 766 -104 800 -88
rect 880 88 914 104
rect 880 -104 914 -88
rect 976 88 1010 104
rect 976 -104 1010 -88
rect 1090 88 1124 104
rect 1090 -104 1124 -88
rect 1186 88 1220 104
rect 1186 -104 1220 -88
rect 1300 88 1334 104
rect 1300 -104 1334 -88
rect 1396 88 1430 104
rect 1396 -104 1430 -88
rect 1510 88 1544 104
rect 1510 -104 1544 -88
rect 1606 88 1640 104
rect 1606 -104 1640 -88
rect 1720 88 1754 104
rect 1720 -104 1754 -88
rect 1816 88 1850 104
rect 1816 -104 1850 -88
rect 1930 88 1964 104
rect 1930 -104 1964 -88
rect 2026 88 2060 104
rect 2026 -104 2060 -88
rect 2140 88 2174 104
rect 2140 -104 2174 -88
rect 2236 88 2270 104
rect 2236 -104 2270 -88
rect 2350 88 2384 104
rect 2350 -104 2384 -88
rect 2446 88 2480 104
rect 2446 -104 2480 -88
rect 2560 88 2594 104
rect 2560 -104 2594 -88
rect 2656 88 2690 104
rect 2656 -104 2690 -88
rect 2770 88 2804 104
rect 2770 -104 2804 -88
rect 2866 88 2900 104
rect 2866 -104 2900 -88
rect 2980 88 3014 104
rect 2980 -104 3014 -88
rect 3076 88 3110 104
rect 3076 -104 3110 -88
rect 3190 88 3224 104
rect 3190 -104 3224 -88
rect 3286 88 3320 104
rect 3286 -104 3320 -88
rect 3400 88 3434 104
rect 3400 -104 3434 -88
rect 3496 88 3530 104
rect 3496 -104 3530 -88
rect 3610 88 3644 104
rect 3610 -104 3644 -88
rect 3706 88 3740 104
rect 3706 -104 3740 -88
rect 3820 88 3854 104
rect 3820 -104 3854 -88
rect 3916 88 3950 104
rect 3916 -104 3950 -88
rect 4030 88 4064 104
rect 4030 -104 4064 -88
rect 4126 88 4160 104
rect 4126 -104 4160 -88
rect 4240 88 4274 147
rect 4240 -104 4274 -88
rect 4336 88 4370 147
rect 4336 -104 4370 -88
rect -4450 -181 -4322 -147
rect -4288 -181 -4240 -147
rect -3918 -181 -3902 -147
rect -3868 -181 -3852 -147
rect -3498 -181 -3482 -147
rect -3448 -181 -3432 -147
rect -3078 -181 -3062 -147
rect -3028 -181 -3012 -147
rect -2658 -181 -2642 -147
rect -2608 -181 -2592 -147
rect -2238 -181 -2222 -147
rect -2188 -181 -2172 -147
rect -1818 -181 -1802 -147
rect -1768 -181 -1752 -147
rect -1398 -181 -1382 -147
rect -1348 -181 -1332 -147
rect -978 -181 -962 -147
rect -928 -181 -912 -147
rect -558 -181 -542 -147
rect -508 -181 -492 -147
rect -138 -181 -122 -147
rect -88 -181 -72 -147
rect 282 -181 298 -147
rect 332 -181 348 -147
rect 702 -181 718 -147
rect 752 -181 768 -147
rect 1122 -181 1138 -147
rect 1172 -181 1188 -147
rect 1542 -181 1558 -147
rect 1592 -181 1608 -147
rect 1962 -181 1978 -147
rect 2012 -181 2028 -147
rect 2382 -181 2398 -147
rect 2432 -181 2448 -147
rect 2802 -181 2818 -147
rect 2852 -181 2868 -147
rect 3222 -181 3238 -147
rect 3272 -181 3288 -147
rect 3642 -181 3658 -147
rect 3692 -181 3708 -147
rect 4062 -181 4078 -147
rect 4112 -181 4128 -147
rect -4484 -345 -4450 -187
rect 4450 -345 4484 -187
rect -4126 -385 -4110 -351
rect -4076 -385 -4060 -351
rect -3706 -385 -3690 -351
rect -3656 -385 -3640 -351
rect -3286 -385 -3270 -351
rect -3236 -385 -3220 -351
rect -2866 -385 -2850 -351
rect -2816 -385 -2800 -351
rect -2446 -385 -2430 -351
rect -2396 -385 -2380 -351
rect -2026 -385 -2010 -351
rect -1976 -385 -1960 -351
rect -1606 -385 -1590 -351
rect -1556 -385 -1540 -351
rect -1186 -385 -1170 -351
rect -1136 -385 -1120 -351
rect -766 -385 -750 -351
rect -716 -385 -700 -351
rect -346 -385 -330 -351
rect -296 -385 -280 -351
rect 74 -385 90 -351
rect 124 -385 140 -351
rect 494 -385 510 -351
rect 544 -385 560 -351
rect 914 -385 930 -351
rect 964 -385 980 -351
rect 1334 -385 1350 -351
rect 1384 -385 1400 -351
rect 1754 -385 1770 -351
rect 1804 -385 1820 -351
rect 2174 -385 2190 -351
rect 2224 -385 2240 -351
rect 2594 -385 2610 -351
rect 2644 -385 2660 -351
rect 3014 -385 3030 -351
rect 3064 -385 3080 -351
rect 3434 -385 3450 -351
rect 3484 -385 3500 -351
rect 3854 -385 3870 -351
rect 3904 -385 3920 -351
rect 4242 -385 4290 -351
rect 4324 -385 4450 -351
rect -4368 -444 -4334 -428
rect -4368 -679 -4334 -620
rect -4272 -444 -4238 -428
rect -4272 -679 -4238 -620
rect -4158 -444 -4124 -428
rect -4158 -636 -4124 -620
rect -4062 -444 -4028 -428
rect -4062 -636 -4028 -620
rect -3948 -444 -3914 -428
rect -3948 -636 -3914 -620
rect -3852 -444 -3818 -428
rect -3852 -636 -3818 -620
rect -3738 -444 -3704 -428
rect -3738 -636 -3704 -620
rect -3642 -444 -3608 -428
rect -3642 -636 -3608 -620
rect -3528 -444 -3494 -428
rect -3528 -636 -3494 -620
rect -3432 -444 -3398 -428
rect -3432 -636 -3398 -620
rect -3318 -444 -3284 -428
rect -3318 -636 -3284 -620
rect -3222 -444 -3188 -428
rect -3222 -636 -3188 -620
rect -3108 -444 -3074 -428
rect -3108 -636 -3074 -620
rect -3012 -444 -2978 -428
rect -3012 -636 -2978 -620
rect -2898 -444 -2864 -428
rect -2898 -636 -2864 -620
rect -2802 -444 -2768 -428
rect -2802 -636 -2768 -620
rect -2688 -444 -2654 -428
rect -2688 -636 -2654 -620
rect -2592 -444 -2558 -428
rect -2592 -636 -2558 -620
rect -2478 -444 -2444 -428
rect -2478 -636 -2444 -620
rect -2382 -444 -2348 -428
rect -2382 -636 -2348 -620
rect -2268 -444 -2234 -428
rect -2268 -636 -2234 -620
rect -2172 -444 -2138 -428
rect -2172 -636 -2138 -620
rect -2058 -444 -2024 -428
rect -2058 -636 -2024 -620
rect -1962 -444 -1928 -428
rect -1962 -636 -1928 -620
rect -1848 -444 -1814 -428
rect -1848 -636 -1814 -620
rect -1752 -444 -1718 -428
rect -1752 -636 -1718 -620
rect -1638 -444 -1604 -428
rect -1638 -636 -1604 -620
rect -1542 -444 -1508 -428
rect -1542 -636 -1508 -620
rect -1428 -444 -1394 -428
rect -1428 -636 -1394 -620
rect -1332 -444 -1298 -428
rect -1332 -636 -1298 -620
rect -1218 -444 -1184 -428
rect -1218 -636 -1184 -620
rect -1122 -444 -1088 -428
rect -1122 -636 -1088 -620
rect -1008 -444 -974 -428
rect -1008 -636 -974 -620
rect -912 -444 -878 -428
rect -912 -636 -878 -620
rect -798 -444 -764 -428
rect -798 -636 -764 -620
rect -702 -444 -668 -428
rect -702 -636 -668 -620
rect -588 -444 -554 -428
rect -588 -636 -554 -620
rect -492 -444 -458 -428
rect -492 -636 -458 -620
rect -378 -444 -344 -428
rect -378 -636 -344 -620
rect -282 -444 -248 -428
rect -282 -636 -248 -620
rect -168 -444 -134 -428
rect -168 -636 -134 -620
rect -72 -444 -38 -428
rect -72 -636 -38 -620
rect 42 -444 76 -428
rect 42 -636 76 -620
rect 138 -444 172 -428
rect 138 -636 172 -620
rect 252 -444 286 -428
rect 252 -636 286 -620
rect 348 -444 382 -428
rect 348 -636 382 -620
rect 462 -444 496 -428
rect 462 -636 496 -620
rect 558 -444 592 -428
rect 558 -636 592 -620
rect 672 -444 706 -428
rect 672 -636 706 -620
rect 768 -444 802 -428
rect 768 -636 802 -620
rect 882 -444 916 -428
rect 882 -636 916 -620
rect 978 -444 1012 -428
rect 978 -636 1012 -620
rect 1092 -444 1126 -428
rect 1092 -636 1126 -620
rect 1188 -444 1222 -428
rect 1188 -636 1222 -620
rect 1302 -444 1336 -428
rect 1302 -636 1336 -620
rect 1398 -444 1432 -428
rect 1398 -636 1432 -620
rect 1512 -444 1546 -428
rect 1512 -636 1546 -620
rect 1608 -444 1642 -428
rect 1608 -636 1642 -620
rect 1722 -444 1756 -428
rect 1722 -636 1756 -620
rect 1818 -444 1852 -428
rect 1818 -636 1852 -620
rect 1932 -444 1966 -428
rect 1932 -636 1966 -620
rect 2028 -444 2062 -428
rect 2028 -636 2062 -620
rect 2142 -444 2176 -428
rect 2142 -636 2176 -620
rect 2238 -444 2272 -428
rect 2238 -636 2272 -620
rect 2352 -444 2386 -428
rect 2352 -636 2386 -620
rect 2448 -444 2482 -428
rect 2448 -636 2482 -620
rect 2562 -444 2596 -428
rect 2562 -636 2596 -620
rect 2658 -444 2692 -428
rect 2658 -636 2692 -620
rect 2772 -444 2806 -428
rect 2772 -636 2806 -620
rect 2868 -444 2902 -428
rect 2868 -636 2902 -620
rect 2982 -444 3016 -428
rect 2982 -636 3016 -620
rect 3078 -444 3112 -428
rect 3078 -636 3112 -620
rect 3192 -444 3226 -428
rect 3192 -636 3226 -620
rect 3288 -444 3322 -428
rect 3288 -636 3322 -620
rect 3402 -444 3436 -428
rect 3402 -636 3436 -620
rect 3498 -444 3532 -428
rect 3498 -636 3532 -620
rect 3612 -444 3646 -428
rect 3612 -636 3646 -620
rect 3708 -444 3742 -428
rect 3708 -636 3742 -620
rect 3822 -444 3856 -428
rect 3822 -636 3856 -620
rect 3918 -444 3952 -428
rect 3918 -636 3952 -620
rect 4032 -444 4066 -428
rect 4032 -636 4066 -620
rect 4128 -444 4162 -428
rect 4128 -636 4162 -620
rect 4242 -444 4276 -385
rect 4242 -636 4276 -620
rect 4338 -444 4372 -385
rect 4338 -636 4372 -620
rect -4450 -713 -4320 -679
rect -4286 -713 -4238 -679
rect -3916 -713 -3900 -679
rect -3866 -713 -3850 -679
rect -3496 -713 -3480 -679
rect -3446 -713 -3430 -679
rect -3076 -713 -3060 -679
rect -3026 -713 -3010 -679
rect -2656 -713 -2640 -679
rect -2606 -713 -2590 -679
rect -2236 -713 -2220 -679
rect -2186 -713 -2170 -679
rect -1816 -713 -1800 -679
rect -1766 -713 -1750 -679
rect -1396 -713 -1380 -679
rect -1346 -713 -1330 -679
rect -976 -713 -960 -679
rect -926 -713 -910 -679
rect -556 -713 -540 -679
rect -506 -713 -490 -679
rect -136 -713 -120 -679
rect -86 -713 -70 -679
rect 284 -713 300 -679
rect 334 -713 350 -679
rect 704 -713 720 -679
rect 754 -713 770 -679
rect 1124 -713 1140 -679
rect 1174 -713 1190 -679
rect 1544 -713 1560 -679
rect 1594 -713 1610 -679
rect 1964 -713 1980 -679
rect 2014 -713 2030 -679
rect 2384 -713 2400 -679
rect 2434 -713 2450 -679
rect 2804 -713 2820 -679
rect 2854 -713 2870 -679
rect 3224 -713 3240 -679
rect 3274 -713 3290 -679
rect 3644 -713 3660 -679
rect 3694 -713 3710 -679
rect 4064 -713 4080 -679
rect 4114 -713 4130 -679
rect -4484 -781 -4450 -719
rect 4450 -781 4484 -719
rect -4484 -815 -4388 -781
rect 4388 -815 4484 -781
<< viali >>
rect -4112 147 -4078 181
rect -3692 147 -3658 181
rect -3272 147 -3238 181
rect -2852 147 -2818 181
rect -2432 147 -2398 181
rect -2012 147 -1978 181
rect -1592 147 -1558 181
rect -1172 147 -1138 181
rect -752 147 -718 181
rect -332 147 -298 181
rect 88 147 122 181
rect 508 147 542 181
rect 928 147 962 181
rect 1348 147 1382 181
rect 1768 147 1802 181
rect 2188 147 2222 181
rect 2608 147 2642 181
rect 3028 147 3062 181
rect 3448 147 3482 181
rect 3868 147 3902 181
rect -3902 -181 -3868 -147
rect -3482 -181 -3448 -147
rect -3062 -181 -3028 -147
rect -2642 -181 -2608 -147
rect -2222 -181 -2188 -147
rect -1802 -181 -1768 -147
rect -1382 -181 -1348 -147
rect -962 -181 -928 -147
rect -542 -181 -508 -147
rect -122 -181 -88 -147
rect 298 -181 332 -147
rect 718 -181 752 -147
rect 1138 -181 1172 -147
rect 1558 -181 1592 -147
rect 1978 -181 2012 -147
rect 2398 -181 2432 -147
rect 2818 -181 2852 -147
rect 3238 -181 3272 -147
rect 3658 -181 3692 -147
rect 4078 -181 4112 -147
rect -4110 -385 -4076 -351
rect -3690 -385 -3656 -351
rect -3270 -385 -3236 -351
rect -2850 -385 -2816 -351
rect -2430 -385 -2396 -351
rect -2010 -385 -1976 -351
rect -1590 -385 -1556 -351
rect -1170 -385 -1136 -351
rect -750 -385 -716 -351
rect -330 -385 -296 -351
rect 90 -385 124 -351
rect 510 -385 544 -351
rect 930 -385 964 -351
rect 1350 -385 1384 -351
rect 1770 -385 1804 -351
rect 2190 -385 2224 -351
rect 2610 -385 2644 -351
rect 3030 -385 3064 -351
rect 3450 -385 3484 -351
rect 3870 -385 3904 -351
rect -3900 -713 -3866 -679
rect -3480 -713 -3446 -679
rect -3060 -713 -3026 -679
rect -2640 -713 -2606 -679
rect -2220 -713 -2186 -679
rect -1800 -713 -1766 -679
rect -1380 -713 -1346 -679
rect -960 -713 -926 -679
rect -540 -713 -506 -679
rect -120 -713 -86 -679
rect 300 -713 334 -679
rect 720 -713 754 -679
rect 1140 -713 1174 -679
rect 1560 -713 1594 -679
rect 1980 -713 2014 -679
rect 2400 -713 2434 -679
rect 2820 -713 2854 -679
rect 3240 -713 3274 -679
rect 3660 -713 3694 -679
rect 4080 -713 4114 -679
<< metal1 >>
rect -4124 181 -4066 187
rect -4124 147 -4112 181
rect -4078 147 -4066 181
rect -4124 141 -4066 147
rect -3704 181 -3646 187
rect -3704 147 -3692 181
rect -3658 147 -3646 181
rect -3704 141 -3646 147
rect -3284 181 -3226 187
rect -3284 147 -3272 181
rect -3238 147 -3226 181
rect -3284 141 -3226 147
rect -2864 181 -2806 187
rect -2864 147 -2852 181
rect -2818 147 -2806 181
rect -2864 141 -2806 147
rect -2444 181 -2386 187
rect -2444 147 -2432 181
rect -2398 147 -2386 181
rect -2444 141 -2386 147
rect -2024 181 -1966 187
rect -2024 147 -2012 181
rect -1978 147 -1966 181
rect -2024 141 -1966 147
rect -1604 181 -1546 187
rect -1604 147 -1592 181
rect -1558 147 -1546 181
rect -1604 141 -1546 147
rect -1184 181 -1126 187
rect -1184 147 -1172 181
rect -1138 147 -1126 181
rect -1184 141 -1126 147
rect -764 181 -706 187
rect -764 147 -752 181
rect -718 147 -706 181
rect -764 141 -706 147
rect -344 181 -286 187
rect -344 147 -332 181
rect -298 147 -286 181
rect -344 141 -286 147
rect 76 181 134 187
rect 76 147 88 181
rect 122 147 134 181
rect 76 141 134 147
rect 496 181 554 187
rect 496 147 508 181
rect 542 147 554 181
rect 496 141 554 147
rect 916 181 974 187
rect 916 147 928 181
rect 962 147 974 181
rect 916 141 974 147
rect 1336 181 1394 187
rect 1336 147 1348 181
rect 1382 147 1394 181
rect 1336 141 1394 147
rect 1756 181 1814 187
rect 1756 147 1768 181
rect 1802 147 1814 181
rect 1756 141 1814 147
rect 2176 181 2234 187
rect 2176 147 2188 181
rect 2222 147 2234 181
rect 2176 141 2234 147
rect 2596 181 2654 187
rect 2596 147 2608 181
rect 2642 147 2654 181
rect 2596 141 2654 147
rect 3016 181 3074 187
rect 3016 147 3028 181
rect 3062 147 3074 181
rect 3016 141 3074 147
rect 3436 181 3494 187
rect 3436 147 3448 181
rect 3482 147 3494 181
rect 3436 141 3494 147
rect 3856 181 3914 187
rect 3856 147 3868 181
rect 3902 147 3914 181
rect 3856 141 3914 147
rect -3914 -147 -3856 -141
rect -3914 -181 -3902 -147
rect -3868 -181 -3856 -147
rect -3914 -187 -3856 -181
rect -3494 -147 -3436 -141
rect -3494 -181 -3482 -147
rect -3448 -181 -3436 -147
rect -3494 -187 -3436 -181
rect -3074 -147 -3016 -141
rect -3074 -181 -3062 -147
rect -3028 -181 -3016 -147
rect -3074 -187 -3016 -181
rect -2654 -147 -2596 -141
rect -2654 -181 -2642 -147
rect -2608 -181 -2596 -147
rect -2654 -187 -2596 -181
rect -2234 -147 -2176 -141
rect -2234 -181 -2222 -147
rect -2188 -181 -2176 -147
rect -2234 -187 -2176 -181
rect -1814 -147 -1756 -141
rect -1814 -181 -1802 -147
rect -1768 -181 -1756 -147
rect -1814 -187 -1756 -181
rect -1394 -147 -1336 -141
rect -1394 -181 -1382 -147
rect -1348 -181 -1336 -147
rect -1394 -187 -1336 -181
rect -974 -147 -916 -141
rect -974 -181 -962 -147
rect -928 -181 -916 -147
rect -974 -187 -916 -181
rect -554 -147 -496 -141
rect -554 -181 -542 -147
rect -508 -181 -496 -147
rect -554 -187 -496 -181
rect -134 -147 -76 -141
rect -134 -181 -122 -147
rect -88 -181 -76 -147
rect -134 -187 -76 -181
rect 286 -147 344 -141
rect 286 -181 298 -147
rect 332 -181 344 -147
rect 286 -187 344 -181
rect 706 -147 764 -141
rect 706 -181 718 -147
rect 752 -181 764 -147
rect 706 -187 764 -181
rect 1126 -147 1184 -141
rect 1126 -181 1138 -147
rect 1172 -181 1184 -147
rect 1126 -187 1184 -181
rect 1546 -147 1604 -141
rect 1546 -181 1558 -147
rect 1592 -181 1604 -147
rect 1546 -187 1604 -181
rect 1966 -147 2024 -141
rect 1966 -181 1978 -147
rect 2012 -181 2024 -147
rect 1966 -187 2024 -181
rect 2386 -147 2444 -141
rect 2386 -181 2398 -147
rect 2432 -181 2444 -147
rect 2386 -187 2444 -181
rect 2806 -147 2864 -141
rect 2806 -181 2818 -147
rect 2852 -181 2864 -147
rect 2806 -187 2864 -181
rect 3226 -147 3284 -141
rect 3226 -181 3238 -147
rect 3272 -181 3284 -147
rect 3226 -187 3284 -181
rect 3646 -147 3704 -141
rect 3646 -181 3658 -147
rect 3692 -181 3704 -147
rect 3646 -187 3704 -181
rect 4066 -147 4124 -141
rect 4066 -181 4078 -147
rect 4112 -181 4124 -147
rect 4066 -187 4124 -181
rect -4122 -351 -4064 -345
rect -4122 -385 -4110 -351
rect -4076 -385 -4064 -351
rect -4122 -391 -4064 -385
rect -3702 -351 -3644 -345
rect -3702 -385 -3690 -351
rect -3656 -385 -3644 -351
rect -3702 -391 -3644 -385
rect -3282 -351 -3224 -345
rect -3282 -385 -3270 -351
rect -3236 -385 -3224 -351
rect -3282 -391 -3224 -385
rect -2862 -351 -2804 -345
rect -2862 -385 -2850 -351
rect -2816 -385 -2804 -351
rect -2862 -391 -2804 -385
rect -2442 -351 -2384 -345
rect -2442 -385 -2430 -351
rect -2396 -385 -2384 -351
rect -2442 -391 -2384 -385
rect -2022 -351 -1964 -345
rect -2022 -385 -2010 -351
rect -1976 -385 -1964 -351
rect -2022 -391 -1964 -385
rect -1602 -351 -1544 -345
rect -1602 -385 -1590 -351
rect -1556 -385 -1544 -351
rect -1602 -391 -1544 -385
rect -1182 -351 -1124 -345
rect -1182 -385 -1170 -351
rect -1136 -385 -1124 -351
rect -1182 -391 -1124 -385
rect -762 -351 -704 -345
rect -762 -385 -750 -351
rect -716 -385 -704 -351
rect -762 -391 -704 -385
rect -342 -351 -284 -345
rect -342 -385 -330 -351
rect -296 -385 -284 -351
rect -342 -391 -284 -385
rect 78 -351 136 -345
rect 78 -385 90 -351
rect 124 -385 136 -351
rect 78 -391 136 -385
rect 498 -351 556 -345
rect 498 -385 510 -351
rect 544 -385 556 -351
rect 498 -391 556 -385
rect 918 -351 976 -345
rect 918 -385 930 -351
rect 964 -385 976 -351
rect 918 -391 976 -385
rect 1338 -351 1396 -345
rect 1338 -385 1350 -351
rect 1384 -385 1396 -351
rect 1338 -391 1396 -385
rect 1758 -351 1816 -345
rect 1758 -385 1770 -351
rect 1804 -385 1816 -351
rect 1758 -391 1816 -385
rect 2178 -351 2236 -345
rect 2178 -385 2190 -351
rect 2224 -385 2236 -351
rect 2178 -391 2236 -385
rect 2598 -351 2656 -345
rect 2598 -385 2610 -351
rect 2644 -385 2656 -351
rect 2598 -391 2656 -385
rect 3018 -351 3076 -345
rect 3018 -385 3030 -351
rect 3064 -385 3076 -351
rect 3018 -391 3076 -385
rect 3438 -351 3496 -345
rect 3438 -385 3450 -351
rect 3484 -385 3496 -351
rect 3438 -391 3496 -385
rect 3858 -351 3916 -345
rect 3858 -385 3870 -351
rect 3904 -385 3916 -351
rect 3858 -391 3916 -385
rect -3912 -679 -3854 -673
rect -3912 -713 -3900 -679
rect -3866 -713 -3854 -679
rect -3912 -719 -3854 -713
rect -3492 -679 -3434 -673
rect -3492 -713 -3480 -679
rect -3446 -713 -3434 -679
rect -3492 -719 -3434 -713
rect -3072 -679 -3014 -673
rect -3072 -713 -3060 -679
rect -3026 -713 -3014 -679
rect -3072 -719 -3014 -713
rect -2652 -679 -2594 -673
rect -2652 -713 -2640 -679
rect -2606 -713 -2594 -679
rect -2652 -719 -2594 -713
rect -2232 -679 -2174 -673
rect -2232 -713 -2220 -679
rect -2186 -713 -2174 -679
rect -2232 -719 -2174 -713
rect -1812 -679 -1754 -673
rect -1812 -713 -1800 -679
rect -1766 -713 -1754 -679
rect -1812 -719 -1754 -713
rect -1392 -679 -1334 -673
rect -1392 -713 -1380 -679
rect -1346 -713 -1334 -679
rect -1392 -719 -1334 -713
rect -972 -679 -914 -673
rect -972 -713 -960 -679
rect -926 -713 -914 -679
rect -972 -719 -914 -713
rect -552 -679 -494 -673
rect -552 -713 -540 -679
rect -506 -713 -494 -679
rect -552 -719 -494 -713
rect -132 -679 -74 -673
rect -132 -713 -120 -679
rect -86 -713 -74 -679
rect -132 -719 -74 -713
rect 288 -679 346 -673
rect 288 -713 300 -679
rect 334 -713 346 -679
rect 288 -719 346 -713
rect 708 -679 766 -673
rect 708 -713 720 -679
rect 754 -713 766 -679
rect 708 -719 766 -713
rect 1128 -679 1186 -673
rect 1128 -713 1140 -679
rect 1174 -713 1186 -679
rect 1128 -719 1186 -713
rect 1548 -679 1606 -673
rect 1548 -713 1560 -679
rect 1594 -713 1606 -679
rect 1548 -719 1606 -713
rect 1968 -679 2026 -673
rect 1968 -713 1980 -679
rect 2014 -713 2026 -679
rect 1968 -719 2026 -713
rect 2388 -679 2446 -673
rect 2388 -713 2400 -679
rect 2434 -713 2446 -679
rect 2388 -719 2446 -713
rect 2808 -679 2866 -673
rect 2808 -713 2820 -679
rect 2854 -713 2866 -679
rect 2808 -719 2866 -713
rect 3228 -679 3286 -673
rect 3228 -713 3240 -679
rect 3274 -713 3286 -679
rect 3228 -719 3286 -713
rect 3648 -679 3706 -673
rect 3648 -713 3660 -679
rect 3694 -713 3706 -679
rect 3648 -719 3706 -713
rect 4068 -679 4126 -673
rect 4068 -713 4080 -679
rect 4114 -713 4126 -679
rect 4068 -719 4126 -713
<< properties >>
string FIXED_BBOX -4467 -266 4467 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 42 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
