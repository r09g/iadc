magic
tech sky130A
magscale 1 2
timestamp 1654898484
<< error_p >>
rect 230 448 288 454
rect 422 448 480 454
rect 614 448 672 454
rect 806 448 864 454
rect 998 448 1056 454
rect 1190 448 1248 454
rect 1382 448 1440 454
rect 1574 448 1632 454
rect 230 414 242 448
rect 422 414 434 448
rect 614 414 626 448
rect 806 414 818 448
rect 998 414 1010 448
rect 1190 414 1202 448
rect 1382 414 1394 448
rect 1574 414 1586 448
rect 230 408 288 414
rect 422 408 480 414
rect 614 408 672 414
rect 806 408 864 414
rect 998 408 1056 414
rect 1190 408 1248 414
rect 1382 408 1440 414
rect 1574 408 1632 414
rect 326 120 384 126
rect 518 120 576 126
rect 710 120 768 126
rect 902 120 960 126
rect 1094 120 1152 126
rect 1286 120 1344 126
rect 1478 120 1536 126
rect 1670 120 1728 126
rect 326 86 338 120
rect 518 86 530 120
rect 710 86 722 120
rect 902 86 914 120
rect 1094 86 1106 120
rect 1286 86 1298 120
rect 1478 86 1490 120
rect 1670 86 1682 120
rect 326 80 384 86
rect 518 80 576 86
rect 710 80 768 86
rect 902 80 960 86
rect 1094 80 1152 86
rect 1286 80 1344 86
rect 1478 80 1536 86
rect 1670 80 1728 86
use sky130_fd_pr__pfet_01v8_VCG74W  sky130_fd_pr__pfet_01v8_VCG74W_0
timestamp 1654898484
transform 1 0 979 0 1 267
box -1031 -319 1031 319
<< end >>
