magic
tech sky130A
timestamp 1654711401
<< error_p >>
rect -374 90 -345 93
rect -278 90 -249 93
rect -182 90 -153 93
rect -86 90 -57 93
rect 9 90 38 93
rect 105 90 134 93
rect 201 90 230 93
rect 297 90 326 93
rect -374 73 -368 90
rect -278 73 -272 90
rect -182 73 -176 90
rect -86 73 -80 90
rect 9 73 15 90
rect 105 73 111 90
rect 201 73 207 90
rect 297 73 303 90
rect -374 70 -345 73
rect -278 70 -249 73
rect -182 70 -153 73
rect -86 70 -57 73
rect 9 70 38 73
rect 105 70 134 73
rect 201 70 230 73
rect 297 70 326 73
rect -326 -73 -297 -70
rect -230 -73 -201 -70
rect -134 -73 -105 -70
rect -38 -73 -9 -70
rect 57 -73 86 -70
rect 153 -73 182 -70
rect 249 -73 278 -70
rect 345 -73 374 -70
rect -326 -90 -320 -73
rect -230 -90 -224 -73
rect -134 -90 -128 -73
rect -38 -90 -32 -73
rect 57 -90 63 -73
rect 153 -90 159 -73
rect 249 -90 255 -73
rect 345 -90 351 -73
rect -326 -93 -297 -90
rect -230 -93 -201 -90
rect -134 -93 -105 -90
rect -38 -93 -9 -90
rect 57 -93 86 -90
rect 153 -93 182 -90
rect 249 -93 278 -90
rect 345 -93 374 -90
<< nwell >>
rect -515 -159 515 159
<< pmos >>
rect -415 -50 -400 50
rect -367 -50 -352 50
rect -319 -50 -304 50
rect -271 -50 -256 50
rect -223 -50 -208 50
rect -175 -50 -160 50
rect -127 -50 -112 50
rect -79 -50 -64 50
rect -31 -50 -16 50
rect 16 -50 31 50
rect 64 -50 79 50
rect 112 -50 127 50
rect 160 -50 175 50
rect 208 -50 223 50
rect 256 -50 271 50
rect 304 -50 319 50
rect 352 -50 367 50
rect 400 -50 415 50
<< pdiff >>
rect -446 44 -415 50
rect -446 -44 -440 44
rect -423 -44 -415 44
rect -446 -50 -415 -44
rect -400 44 -367 50
rect -400 -44 -392 44
rect -375 -44 -367 44
rect -400 -50 -367 -44
rect -352 44 -319 50
rect -352 -44 -344 44
rect -327 -44 -319 44
rect -352 -50 -319 -44
rect -304 44 -271 50
rect -304 -44 -296 44
rect -279 -44 -271 44
rect -304 -50 -271 -44
rect -256 44 -223 50
rect -256 -44 -248 44
rect -231 -44 -223 44
rect -256 -50 -223 -44
rect -208 44 -175 50
rect -208 -44 -200 44
rect -183 -44 -175 44
rect -208 -50 -175 -44
rect -160 44 -127 50
rect -160 -44 -152 44
rect -135 -44 -127 44
rect -160 -50 -127 -44
rect -112 44 -79 50
rect -112 -44 -104 44
rect -87 -44 -79 44
rect -112 -50 -79 -44
rect -64 44 -31 50
rect -64 -44 -56 44
rect -39 -44 -31 44
rect -64 -50 -31 -44
rect -16 44 16 50
rect -16 -44 -8 44
rect 8 -44 16 44
rect -16 -50 16 -44
rect 31 44 64 50
rect 31 -44 39 44
rect 56 -44 64 44
rect 31 -50 64 -44
rect 79 44 112 50
rect 79 -44 87 44
rect 104 -44 112 44
rect 79 -50 112 -44
rect 127 44 160 50
rect 127 -44 135 44
rect 152 -44 160 44
rect 127 -50 160 -44
rect 175 44 208 50
rect 175 -44 183 44
rect 200 -44 208 44
rect 175 -50 208 -44
rect 223 44 256 50
rect 223 -44 231 44
rect 248 -44 256 44
rect 223 -50 256 -44
rect 271 44 304 50
rect 271 -44 279 44
rect 296 -44 304 44
rect 271 -50 304 -44
rect 319 44 352 50
rect 319 -44 327 44
rect 344 -44 352 44
rect 319 -50 352 -44
rect 367 44 400 50
rect 367 -44 375 44
rect 392 -44 400 44
rect 367 -50 400 -44
rect 415 44 446 50
rect 415 -44 423 44
rect 440 -44 446 44
rect 415 -50 446 -44
<< pdiffc >>
rect -440 -44 -423 44
rect -392 -44 -375 44
rect -344 -44 -327 44
rect -296 -44 -279 44
rect -248 -44 -231 44
rect -200 -44 -183 44
rect -152 -44 -135 44
rect -104 -44 -87 44
rect -56 -44 -39 44
rect -8 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
<< nsubdiff >>
rect -497 124 -449 141
rect 449 124 497 141
rect -497 93 -480 124
rect 480 93 497 124
rect -497 -124 -480 -93
rect 480 -124 497 -93
rect -497 -141 -449 -124
rect 449 -141 497 -124
<< nsubdiffcont >>
rect -449 124 449 141
rect -497 -93 -480 93
rect 480 -93 497 93
rect -449 -141 449 -124
<< poly >>
rect -376 90 -343 98
rect -376 73 -368 90
rect -351 73 -343 90
rect -376 65 -343 73
rect -280 90 -247 98
rect -280 73 -272 90
rect -255 73 -247 90
rect -280 65 -247 73
rect -184 90 -151 98
rect -184 73 -176 90
rect -159 73 -151 90
rect -184 65 -151 73
rect -88 90 -55 98
rect -88 73 -80 90
rect -63 73 -55 90
rect -88 65 -55 73
rect 7 90 40 98
rect 7 73 15 90
rect 32 73 40 90
rect 7 65 40 73
rect 103 90 136 98
rect 103 73 111 90
rect 128 73 136 90
rect 103 65 136 73
rect 199 90 232 98
rect 199 73 207 90
rect 224 73 232 90
rect 199 65 232 73
rect 295 90 328 98
rect 295 73 303 90
rect 320 73 328 90
rect 295 65 328 73
rect 391 90 424 98
rect 391 73 399 90
rect 416 73 424 90
rect 391 65 424 73
rect -415 50 -400 63
rect -367 50 -352 65
rect -319 50 -304 63
rect -271 50 -256 65
rect -223 50 -208 63
rect -175 50 -160 65
rect -127 50 -112 63
rect -79 50 -64 65
rect -31 50 -16 63
rect 16 50 31 65
rect 64 50 79 63
rect 112 50 127 65
rect 160 50 175 63
rect 208 50 223 65
rect 256 50 271 63
rect 304 50 319 65
rect 352 50 367 63
rect 400 50 415 65
rect -415 -65 -400 -50
rect -367 -63 -352 -50
rect -319 -65 -304 -50
rect -271 -63 -256 -50
rect -223 -65 -208 -50
rect -175 -63 -160 -50
rect -127 -65 -112 -50
rect -79 -63 -64 -50
rect -31 -65 -16 -50
rect 16 -63 31 -50
rect 64 -65 79 -50
rect 112 -63 127 -50
rect 160 -65 175 -50
rect 208 -63 223 -50
rect 256 -65 271 -50
rect 304 -63 319 -50
rect 352 -65 367 -50
rect 400 -63 415 -50
rect -424 -73 -391 -65
rect -424 -90 -416 -73
rect -399 -90 -391 -73
rect -424 -98 -391 -90
rect -328 -73 -295 -65
rect -328 -90 -320 -73
rect -303 -90 -295 -73
rect -328 -98 -295 -90
rect -232 -73 -199 -65
rect -232 -90 -224 -73
rect -207 -90 -199 -73
rect -232 -98 -199 -90
rect -136 -73 -103 -65
rect -136 -90 -128 -73
rect -111 -90 -103 -73
rect -136 -98 -103 -90
rect -40 -73 -7 -65
rect -40 -90 -32 -73
rect -15 -90 -7 -73
rect -40 -98 -7 -90
rect 55 -73 88 -65
rect 55 -90 63 -73
rect 80 -90 88 -73
rect 55 -98 88 -90
rect 151 -73 184 -65
rect 151 -90 159 -73
rect 176 -90 184 -73
rect 151 -98 184 -90
rect 247 -73 280 -65
rect 247 -90 255 -73
rect 272 -90 280 -73
rect 247 -98 280 -90
rect 343 -73 376 -65
rect 343 -90 351 -73
rect 368 -90 376 -73
rect 343 -98 376 -90
<< polycont >>
rect -368 73 -351 90
rect -272 73 -255 90
rect -176 73 -159 90
rect -80 73 -63 90
rect 15 73 32 90
rect 111 73 128 90
rect 207 73 224 90
rect 303 73 320 90
rect 399 73 416 90
rect -416 -90 -399 -73
rect -320 -90 -303 -73
rect -224 -90 -207 -73
rect -128 -90 -111 -73
rect -32 -90 -15 -73
rect 63 -90 80 -73
rect 159 -90 176 -73
rect 255 -90 272 -73
rect 351 -90 368 -73
<< locali >>
rect -497 124 -449 141
rect 449 124 497 141
rect -497 93 -480 124
rect 423 90 440 124
rect -376 73 -368 90
rect -351 73 -343 90
rect -280 73 -272 90
rect -255 73 -247 90
rect -184 73 -176 90
rect -159 73 -151 90
rect -88 73 -80 90
rect -63 73 -55 90
rect 7 73 15 90
rect 32 73 40 90
rect 103 73 111 90
rect 128 73 136 90
rect 199 73 207 90
rect 224 73 232 90
rect 295 73 303 90
rect 320 73 328 90
rect 391 73 399 90
rect 416 73 440 90
rect -497 -124 -480 -93
rect -440 44 -423 52
rect -440 -73 -423 -44
rect -392 44 -375 52
rect -392 -52 -375 -44
rect -344 44 -327 52
rect -344 -52 -327 -44
rect -296 44 -279 52
rect -296 -52 -279 -44
rect -248 44 -231 52
rect -248 -52 -231 -44
rect -200 44 -183 52
rect -200 -52 -183 -44
rect -152 44 -135 52
rect -152 -52 -135 -44
rect -104 44 -87 52
rect -104 -52 -87 -44
rect -56 44 -39 52
rect -56 -52 -39 -44
rect -8 44 8 52
rect -8 -52 8 -44
rect 39 44 56 52
rect 39 -52 56 -44
rect 87 44 104 52
rect 87 -52 104 -44
rect 135 44 152 52
rect 135 -52 152 -44
rect 183 44 200 52
rect 183 -52 200 -44
rect 231 44 248 52
rect 231 -52 248 -44
rect 279 44 296 52
rect 279 -52 296 -44
rect 327 44 344 52
rect 327 -52 344 -44
rect 375 44 392 52
rect 375 -52 392 -44
rect 423 44 440 73
rect 423 -52 440 -44
rect 480 93 497 124
rect -440 -90 -416 -73
rect -399 -90 -391 -73
rect -328 -90 -320 -73
rect -303 -90 -295 -73
rect -232 -90 -224 -73
rect -207 -90 -199 -73
rect -136 -90 -128 -73
rect -111 -90 -103 -73
rect -40 -90 -32 -73
rect -15 -90 -7 -73
rect 55 -90 63 -73
rect 80 -90 88 -73
rect 151 -90 159 -73
rect 176 -90 184 -73
rect 247 -90 255 -73
rect 272 -90 280 -73
rect 343 -90 351 -73
rect 368 -90 376 -73
rect -440 -124 -423 -90
rect 480 -124 497 -93
rect -497 -141 -449 -124
rect 449 -141 497 -124
<< viali >>
rect -368 73 -351 90
rect -272 73 -255 90
rect -176 73 -159 90
rect -80 73 -63 90
rect 15 73 32 90
rect 111 73 128 90
rect 207 73 224 90
rect 303 73 320 90
rect -320 -90 -303 -73
rect -224 -90 -207 -73
rect -128 -90 -111 -73
rect -32 -90 -15 -73
rect 63 -90 80 -73
rect 159 -90 176 -73
rect 255 -90 272 -73
rect 351 -90 368 -73
<< metal1 >>
rect -374 90 -345 93
rect -374 73 -368 90
rect -351 73 -345 90
rect -374 70 -345 73
rect -278 90 -249 93
rect -278 73 -272 90
rect -255 73 -249 90
rect -278 70 -249 73
rect -182 90 -153 93
rect -182 73 -176 90
rect -159 73 -153 90
rect -182 70 -153 73
rect -86 90 -57 93
rect -86 73 -80 90
rect -63 73 -57 90
rect -86 70 -57 73
rect 9 90 38 93
rect 9 73 15 90
rect 32 73 38 90
rect 9 70 38 73
rect 105 90 134 93
rect 105 73 111 90
rect 128 73 134 90
rect 105 70 134 73
rect 201 90 230 93
rect 201 73 207 90
rect 224 73 230 90
rect 201 70 230 73
rect 297 90 326 93
rect 297 73 303 90
rect 320 73 326 90
rect 297 70 326 73
rect -326 -73 -297 -70
rect -326 -90 -320 -73
rect -303 -90 -297 -73
rect -326 -93 -297 -90
rect -230 -73 -201 -70
rect -230 -90 -224 -73
rect -207 -90 -201 -73
rect -230 -93 -201 -90
rect -134 -73 -105 -70
rect -134 -90 -128 -73
rect -111 -90 -105 -73
rect -134 -93 -105 -90
rect -38 -73 -9 -70
rect -38 -90 -32 -73
rect -15 -90 -9 -73
rect -38 -93 -9 -90
rect 57 -73 86 -70
rect 57 -90 63 -73
rect 80 -90 86 -73
rect 57 -93 86 -90
rect 153 -73 182 -70
rect 153 -90 159 -73
rect 176 -90 182 -73
rect 153 -93 182 -90
rect 249 -73 278 -70
rect 249 -90 255 -73
rect 272 -90 278 -73
rect 249 -93 278 -90
rect 345 -73 374 -70
rect 345 -90 351 -73
rect 368 -90 374 -73
rect 345 -93 374 -90
<< properties >>
string FIXED_BBOX -489 -133 489 133
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
