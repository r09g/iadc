magic
tech sky130A
timestamp 1653030110
<< nmos >>
rect -1543 -70 -1483 70
rect -1454 -70 -1394 70
rect -1365 -70 -1305 70
rect -1276 -70 -1216 70
rect -1187 -70 -1127 70
rect -1098 -70 -1038 70
rect -1009 -70 -949 70
rect -920 -70 -860 70
rect -831 -70 -771 70
rect -742 -70 -682 70
rect -653 -70 -593 70
rect -564 -70 -504 70
rect -475 -70 -415 70
rect -386 -70 -326 70
rect -297 -70 -237 70
rect -208 -70 -148 70
rect -119 -70 -59 70
rect -30 -70 30 70
rect 59 -70 119 70
rect 148 -70 208 70
rect 237 -70 297 70
rect 326 -70 386 70
rect 415 -70 475 70
rect 504 -70 564 70
rect 593 -70 653 70
rect 682 -70 742 70
rect 771 -70 831 70
rect 860 -70 920 70
rect 949 -70 1009 70
rect 1038 -70 1098 70
rect 1127 -70 1187 70
rect 1216 -70 1276 70
rect 1305 -70 1365 70
rect 1394 -70 1454 70
rect 1483 -70 1543 70
<< ndiff >>
rect -1572 64 -1543 70
rect -1572 -64 -1566 64
rect -1549 -64 -1543 64
rect -1572 -70 -1543 -64
rect -1483 64 -1454 70
rect -1483 -64 -1477 64
rect -1460 -64 -1454 64
rect -1483 -70 -1454 -64
rect -1394 64 -1365 70
rect -1394 -64 -1388 64
rect -1371 -64 -1365 64
rect -1394 -70 -1365 -64
rect -1305 64 -1276 70
rect -1305 -64 -1299 64
rect -1282 -64 -1276 64
rect -1305 -70 -1276 -64
rect -1216 64 -1187 70
rect -1216 -64 -1210 64
rect -1193 -64 -1187 64
rect -1216 -70 -1187 -64
rect -1127 64 -1098 70
rect -1127 -64 -1121 64
rect -1104 -64 -1098 64
rect -1127 -70 -1098 -64
rect -1038 64 -1009 70
rect -1038 -64 -1032 64
rect -1015 -64 -1009 64
rect -1038 -70 -1009 -64
rect -949 64 -920 70
rect -949 -64 -943 64
rect -926 -64 -920 64
rect -949 -70 -920 -64
rect -860 64 -831 70
rect -860 -64 -854 64
rect -837 -64 -831 64
rect -860 -70 -831 -64
rect -771 64 -742 70
rect -771 -64 -765 64
rect -748 -64 -742 64
rect -771 -70 -742 -64
rect -682 64 -653 70
rect -682 -64 -676 64
rect -659 -64 -653 64
rect -682 -70 -653 -64
rect -593 64 -564 70
rect -593 -64 -587 64
rect -570 -64 -564 64
rect -593 -70 -564 -64
rect -504 64 -475 70
rect -504 -64 -498 64
rect -481 -64 -475 64
rect -504 -70 -475 -64
rect -415 64 -386 70
rect -415 -64 -409 64
rect -392 -64 -386 64
rect -415 -70 -386 -64
rect -326 64 -297 70
rect -326 -64 -320 64
rect -303 -64 -297 64
rect -326 -70 -297 -64
rect -237 64 -208 70
rect -237 -64 -231 64
rect -214 -64 -208 64
rect -237 -70 -208 -64
rect -148 64 -119 70
rect -148 -64 -142 64
rect -125 -64 -119 64
rect -148 -70 -119 -64
rect -59 64 -30 70
rect -59 -64 -53 64
rect -36 -64 -30 64
rect -59 -70 -30 -64
rect 30 64 59 70
rect 30 -64 36 64
rect 53 -64 59 64
rect 30 -70 59 -64
rect 119 64 148 70
rect 119 -64 125 64
rect 142 -64 148 64
rect 119 -70 148 -64
rect 208 64 237 70
rect 208 -64 214 64
rect 231 -64 237 64
rect 208 -70 237 -64
rect 297 64 326 70
rect 297 -64 303 64
rect 320 -64 326 64
rect 297 -70 326 -64
rect 386 64 415 70
rect 386 -64 392 64
rect 409 -64 415 64
rect 386 -70 415 -64
rect 475 64 504 70
rect 475 -64 481 64
rect 498 -64 504 64
rect 475 -70 504 -64
rect 564 64 593 70
rect 564 -64 570 64
rect 587 -64 593 64
rect 564 -70 593 -64
rect 653 64 682 70
rect 653 -64 659 64
rect 676 -64 682 64
rect 653 -70 682 -64
rect 742 64 771 70
rect 742 -64 748 64
rect 765 -64 771 64
rect 742 -70 771 -64
rect 831 64 860 70
rect 831 -64 837 64
rect 854 -64 860 64
rect 831 -70 860 -64
rect 920 64 949 70
rect 920 -64 926 64
rect 943 -64 949 64
rect 920 -70 949 -64
rect 1009 64 1038 70
rect 1009 -64 1015 64
rect 1032 -64 1038 64
rect 1009 -70 1038 -64
rect 1098 64 1127 70
rect 1098 -64 1104 64
rect 1121 -64 1127 64
rect 1098 -70 1127 -64
rect 1187 64 1216 70
rect 1187 -64 1193 64
rect 1210 -64 1216 64
rect 1187 -70 1216 -64
rect 1276 64 1305 70
rect 1276 -64 1282 64
rect 1299 -64 1305 64
rect 1276 -70 1305 -64
rect 1365 64 1394 70
rect 1365 -64 1371 64
rect 1388 -64 1394 64
rect 1365 -70 1394 -64
rect 1454 64 1483 70
rect 1454 -64 1460 64
rect 1477 -64 1483 64
rect 1454 -70 1483 -64
rect 1543 64 1572 70
rect 1543 -64 1549 64
rect 1566 -64 1572 64
rect 1543 -70 1572 -64
<< ndiffc >>
rect -1566 -64 -1549 64
rect -1477 -64 -1460 64
rect -1388 -64 -1371 64
rect -1299 -64 -1282 64
rect -1210 -64 -1193 64
rect -1121 -64 -1104 64
rect -1032 -64 -1015 64
rect -943 -64 -926 64
rect -854 -64 -837 64
rect -765 -64 -748 64
rect -676 -64 -659 64
rect -587 -64 -570 64
rect -498 -64 -481 64
rect -409 -64 -392 64
rect -320 -64 -303 64
rect -231 -64 -214 64
rect -142 -64 -125 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 125 -64 142 64
rect 214 -64 231 64
rect 303 -64 320 64
rect 392 -64 409 64
rect 481 -64 498 64
rect 570 -64 587 64
rect 659 -64 676 64
rect 748 -64 765 64
rect 837 -64 854 64
rect 926 -64 943 64
rect 1015 -64 1032 64
rect 1104 -64 1121 64
rect 1193 -64 1210 64
rect 1282 -64 1299 64
rect 1371 -64 1388 64
rect 1460 -64 1477 64
rect 1549 -64 1566 64
<< poly >>
rect -1532 106 -1494 114
rect -1532 97 -1524 106
rect -1543 89 -1524 97
rect -1502 97 -1494 106
rect -1443 106 -1405 114
rect -1443 97 -1435 106
rect -1502 89 -1483 97
rect -1543 70 -1483 89
rect -1454 89 -1435 97
rect -1413 97 -1405 106
rect -1354 106 -1316 114
rect -1354 97 -1346 106
rect -1413 89 -1394 97
rect -1454 70 -1394 89
rect -1365 89 -1346 97
rect -1324 97 -1316 106
rect -1265 106 -1227 114
rect -1265 97 -1257 106
rect -1324 89 -1305 97
rect -1365 70 -1305 89
rect -1276 89 -1257 97
rect -1235 97 -1227 106
rect -1176 106 -1138 114
rect -1176 97 -1168 106
rect -1235 89 -1216 97
rect -1276 70 -1216 89
rect -1187 89 -1168 97
rect -1146 97 -1138 106
rect -1087 106 -1049 114
rect -1087 97 -1079 106
rect -1146 89 -1127 97
rect -1187 70 -1127 89
rect -1098 89 -1079 97
rect -1057 97 -1049 106
rect -998 106 -960 114
rect -998 97 -990 106
rect -1057 89 -1038 97
rect -1098 70 -1038 89
rect -1009 89 -990 97
rect -968 97 -960 106
rect -909 106 -871 114
rect -909 97 -901 106
rect -968 89 -949 97
rect -1009 70 -949 89
rect -920 89 -901 97
rect -879 97 -871 106
rect -820 106 -782 114
rect -820 97 -812 106
rect -879 89 -860 97
rect -920 70 -860 89
rect -831 89 -812 97
rect -790 97 -782 106
rect -731 106 -693 114
rect -731 97 -723 106
rect -790 89 -771 97
rect -831 70 -771 89
rect -742 89 -723 97
rect -701 97 -693 106
rect -642 106 -604 114
rect -642 97 -634 106
rect -701 89 -682 97
rect -742 70 -682 89
rect -653 89 -634 97
rect -612 97 -604 106
rect -553 106 -515 114
rect -553 97 -545 106
rect -612 89 -593 97
rect -653 70 -593 89
rect -564 89 -545 97
rect -523 97 -515 106
rect -464 106 -426 114
rect -464 97 -456 106
rect -523 89 -504 97
rect -564 70 -504 89
rect -475 89 -456 97
rect -434 97 -426 106
rect -375 106 -337 114
rect -375 97 -367 106
rect -434 89 -415 97
rect -475 70 -415 89
rect -386 89 -367 97
rect -345 97 -337 106
rect -286 106 -248 114
rect -286 97 -278 106
rect -345 89 -326 97
rect -386 70 -326 89
rect -297 89 -278 97
rect -256 97 -248 106
rect -197 106 -159 114
rect -197 97 -189 106
rect -256 89 -237 97
rect -297 70 -237 89
rect -208 89 -189 97
rect -167 97 -159 106
rect -108 106 -70 114
rect -108 97 -100 106
rect -167 89 -148 97
rect -208 70 -148 89
rect -119 89 -100 97
rect -78 97 -70 106
rect -19 106 19 114
rect -19 97 -11 106
rect -78 89 -59 97
rect -119 70 -59 89
rect -30 89 -11 97
rect 11 97 19 106
rect 70 106 108 114
rect 70 97 78 106
rect 11 89 30 97
rect -30 70 30 89
rect 59 89 78 97
rect 100 97 108 106
rect 159 106 197 114
rect 159 97 167 106
rect 100 89 119 97
rect 59 70 119 89
rect 148 89 167 97
rect 189 97 197 106
rect 248 106 286 114
rect 248 97 256 106
rect 189 89 208 97
rect 148 70 208 89
rect 237 89 256 97
rect 278 97 286 106
rect 337 106 375 114
rect 337 97 345 106
rect 278 89 297 97
rect 237 70 297 89
rect 326 89 345 97
rect 367 97 375 106
rect 426 106 464 114
rect 426 97 434 106
rect 367 89 386 97
rect 326 70 386 89
rect 415 89 434 97
rect 456 97 464 106
rect 515 106 553 114
rect 515 97 523 106
rect 456 89 475 97
rect 415 70 475 89
rect 504 89 523 97
rect 545 97 553 106
rect 604 106 642 114
rect 604 97 612 106
rect 545 89 564 97
rect 504 70 564 89
rect 593 89 612 97
rect 634 97 642 106
rect 693 106 731 114
rect 693 97 701 106
rect 634 89 653 97
rect 593 70 653 89
rect 682 89 701 97
rect 723 97 731 106
rect 782 106 820 114
rect 782 97 790 106
rect 723 89 742 97
rect 682 70 742 89
rect 771 89 790 97
rect 812 97 820 106
rect 871 106 909 114
rect 871 97 879 106
rect 812 89 831 97
rect 771 70 831 89
rect 860 89 879 97
rect 901 97 909 106
rect 960 106 998 114
rect 960 97 968 106
rect 901 89 920 97
rect 860 70 920 89
rect 949 89 968 97
rect 990 97 998 106
rect 1049 106 1087 114
rect 1049 97 1057 106
rect 990 89 1009 97
rect 949 70 1009 89
rect 1038 89 1057 97
rect 1079 97 1087 106
rect 1138 106 1176 114
rect 1138 97 1146 106
rect 1079 89 1098 97
rect 1038 70 1098 89
rect 1127 89 1146 97
rect 1168 97 1176 106
rect 1227 106 1265 114
rect 1227 97 1235 106
rect 1168 89 1187 97
rect 1127 70 1187 89
rect 1216 89 1235 97
rect 1257 97 1265 106
rect 1316 106 1354 114
rect 1316 97 1324 106
rect 1257 89 1276 97
rect 1216 70 1276 89
rect 1305 89 1324 97
rect 1346 97 1354 106
rect 1405 106 1443 114
rect 1405 97 1413 106
rect 1346 89 1365 97
rect 1305 70 1365 89
rect 1394 89 1413 97
rect 1435 97 1443 106
rect 1494 106 1532 114
rect 1494 97 1502 106
rect 1435 89 1454 97
rect 1394 70 1454 89
rect 1483 89 1502 97
rect 1524 97 1532 106
rect 1524 89 1543 97
rect 1483 70 1543 89
rect -1543 -89 -1483 -70
rect -1543 -97 -1524 -89
rect -1532 -106 -1524 -97
rect -1502 -97 -1483 -89
rect -1454 -89 -1394 -70
rect -1454 -97 -1435 -89
rect -1502 -106 -1494 -97
rect -1532 -114 -1494 -106
rect -1443 -106 -1435 -97
rect -1413 -97 -1394 -89
rect -1365 -89 -1305 -70
rect -1365 -97 -1346 -89
rect -1413 -106 -1405 -97
rect -1443 -114 -1405 -106
rect -1354 -106 -1346 -97
rect -1324 -97 -1305 -89
rect -1276 -89 -1216 -70
rect -1276 -97 -1257 -89
rect -1324 -106 -1316 -97
rect -1354 -114 -1316 -106
rect -1265 -106 -1257 -97
rect -1235 -97 -1216 -89
rect -1187 -89 -1127 -70
rect -1187 -97 -1168 -89
rect -1235 -106 -1227 -97
rect -1265 -114 -1227 -106
rect -1176 -106 -1168 -97
rect -1146 -97 -1127 -89
rect -1098 -89 -1038 -70
rect -1098 -97 -1079 -89
rect -1146 -106 -1138 -97
rect -1176 -114 -1138 -106
rect -1087 -106 -1079 -97
rect -1057 -97 -1038 -89
rect -1009 -89 -949 -70
rect -1009 -97 -990 -89
rect -1057 -106 -1049 -97
rect -1087 -114 -1049 -106
rect -998 -106 -990 -97
rect -968 -97 -949 -89
rect -920 -89 -860 -70
rect -920 -97 -901 -89
rect -968 -106 -960 -97
rect -998 -114 -960 -106
rect -909 -106 -901 -97
rect -879 -97 -860 -89
rect -831 -89 -771 -70
rect -831 -97 -812 -89
rect -879 -106 -871 -97
rect -909 -114 -871 -106
rect -820 -106 -812 -97
rect -790 -97 -771 -89
rect -742 -89 -682 -70
rect -742 -97 -723 -89
rect -790 -106 -782 -97
rect -820 -114 -782 -106
rect -731 -106 -723 -97
rect -701 -97 -682 -89
rect -653 -89 -593 -70
rect -653 -97 -634 -89
rect -701 -106 -693 -97
rect -731 -114 -693 -106
rect -642 -106 -634 -97
rect -612 -97 -593 -89
rect -564 -89 -504 -70
rect -564 -97 -545 -89
rect -612 -106 -604 -97
rect -642 -114 -604 -106
rect -553 -106 -545 -97
rect -523 -97 -504 -89
rect -475 -89 -415 -70
rect -475 -97 -456 -89
rect -523 -106 -515 -97
rect -553 -114 -515 -106
rect -464 -106 -456 -97
rect -434 -97 -415 -89
rect -386 -89 -326 -70
rect -386 -97 -367 -89
rect -434 -106 -426 -97
rect -464 -114 -426 -106
rect -375 -106 -367 -97
rect -345 -97 -326 -89
rect -297 -89 -237 -70
rect -297 -97 -278 -89
rect -345 -106 -337 -97
rect -375 -114 -337 -106
rect -286 -106 -278 -97
rect -256 -97 -237 -89
rect -208 -89 -148 -70
rect -208 -97 -189 -89
rect -256 -106 -248 -97
rect -286 -114 -248 -106
rect -197 -106 -189 -97
rect -167 -97 -148 -89
rect -119 -89 -59 -70
rect -119 -97 -100 -89
rect -167 -106 -159 -97
rect -197 -114 -159 -106
rect -108 -106 -100 -97
rect -78 -97 -59 -89
rect -30 -89 30 -70
rect -30 -97 -11 -89
rect -78 -106 -70 -97
rect -108 -114 -70 -106
rect -19 -106 -11 -97
rect 11 -97 30 -89
rect 59 -89 119 -70
rect 59 -97 78 -89
rect 11 -106 19 -97
rect -19 -114 19 -106
rect 70 -106 78 -97
rect 100 -97 119 -89
rect 148 -89 208 -70
rect 148 -97 167 -89
rect 100 -106 108 -97
rect 70 -114 108 -106
rect 159 -106 167 -97
rect 189 -97 208 -89
rect 237 -89 297 -70
rect 237 -97 256 -89
rect 189 -106 197 -97
rect 159 -114 197 -106
rect 248 -106 256 -97
rect 278 -97 297 -89
rect 326 -89 386 -70
rect 326 -97 345 -89
rect 278 -106 286 -97
rect 248 -114 286 -106
rect 337 -106 345 -97
rect 367 -97 386 -89
rect 415 -89 475 -70
rect 415 -97 434 -89
rect 367 -106 375 -97
rect 337 -114 375 -106
rect 426 -106 434 -97
rect 456 -97 475 -89
rect 504 -89 564 -70
rect 504 -97 523 -89
rect 456 -106 464 -97
rect 426 -114 464 -106
rect 515 -106 523 -97
rect 545 -97 564 -89
rect 593 -89 653 -70
rect 593 -97 612 -89
rect 545 -106 553 -97
rect 515 -114 553 -106
rect 604 -106 612 -97
rect 634 -97 653 -89
rect 682 -89 742 -70
rect 682 -97 701 -89
rect 634 -106 642 -97
rect 604 -114 642 -106
rect 693 -106 701 -97
rect 723 -97 742 -89
rect 771 -89 831 -70
rect 771 -97 790 -89
rect 723 -106 731 -97
rect 693 -114 731 -106
rect 782 -106 790 -97
rect 812 -97 831 -89
rect 860 -89 920 -70
rect 860 -97 879 -89
rect 812 -106 820 -97
rect 782 -114 820 -106
rect 871 -106 879 -97
rect 901 -97 920 -89
rect 949 -89 1009 -70
rect 949 -97 968 -89
rect 901 -106 909 -97
rect 871 -114 909 -106
rect 960 -106 968 -97
rect 990 -97 1009 -89
rect 1038 -89 1098 -70
rect 1038 -97 1057 -89
rect 990 -106 998 -97
rect 960 -114 998 -106
rect 1049 -106 1057 -97
rect 1079 -97 1098 -89
rect 1127 -89 1187 -70
rect 1127 -97 1146 -89
rect 1079 -106 1087 -97
rect 1049 -114 1087 -106
rect 1138 -106 1146 -97
rect 1168 -97 1187 -89
rect 1216 -89 1276 -70
rect 1216 -97 1235 -89
rect 1168 -106 1176 -97
rect 1138 -114 1176 -106
rect 1227 -106 1235 -97
rect 1257 -97 1276 -89
rect 1305 -89 1365 -70
rect 1305 -97 1324 -89
rect 1257 -106 1265 -97
rect 1227 -114 1265 -106
rect 1316 -106 1324 -97
rect 1346 -97 1365 -89
rect 1394 -89 1454 -70
rect 1394 -97 1413 -89
rect 1346 -106 1354 -97
rect 1316 -114 1354 -106
rect 1405 -106 1413 -97
rect 1435 -97 1454 -89
rect 1483 -89 1543 -70
rect 1483 -97 1502 -89
rect 1435 -106 1443 -97
rect 1405 -114 1443 -106
rect 1494 -106 1502 -97
rect 1524 -97 1543 -89
rect 1524 -106 1532 -97
rect 1494 -114 1532 -106
<< polycont >>
rect -1524 89 -1502 106
rect -1435 89 -1413 106
rect -1346 89 -1324 106
rect -1257 89 -1235 106
rect -1168 89 -1146 106
rect -1079 89 -1057 106
rect -990 89 -968 106
rect -901 89 -879 106
rect -812 89 -790 106
rect -723 89 -701 106
rect -634 89 -612 106
rect -545 89 -523 106
rect -456 89 -434 106
rect -367 89 -345 106
rect -278 89 -256 106
rect -189 89 -167 106
rect -100 89 -78 106
rect -11 89 11 106
rect 78 89 100 106
rect 167 89 189 106
rect 256 89 278 106
rect 345 89 367 106
rect 434 89 456 106
rect 523 89 545 106
rect 612 89 634 106
rect 701 89 723 106
rect 790 89 812 106
rect 879 89 901 106
rect 968 89 990 106
rect 1057 89 1079 106
rect 1146 89 1168 106
rect 1235 89 1257 106
rect 1324 89 1346 106
rect 1413 89 1435 106
rect 1502 89 1524 106
rect -1524 -106 -1502 -89
rect -1435 -106 -1413 -89
rect -1346 -106 -1324 -89
rect -1257 -106 -1235 -89
rect -1168 -106 -1146 -89
rect -1079 -106 -1057 -89
rect -990 -106 -968 -89
rect -901 -106 -879 -89
rect -812 -106 -790 -89
rect -723 -106 -701 -89
rect -634 -106 -612 -89
rect -545 -106 -523 -89
rect -456 -106 -434 -89
rect -367 -106 -345 -89
rect -278 -106 -256 -89
rect -189 -106 -167 -89
rect -100 -106 -78 -89
rect -11 -106 11 -89
rect 78 -106 100 -89
rect 167 -106 189 -89
rect 256 -106 278 -89
rect 345 -106 367 -89
rect 434 -106 456 -89
rect 523 -106 545 -89
rect 612 -106 634 -89
rect 701 -106 723 -89
rect 790 -106 812 -89
rect 879 -106 901 -89
rect 968 -106 990 -89
rect 1057 -106 1079 -89
rect 1146 -106 1168 -89
rect 1235 -106 1257 -89
rect 1324 -106 1346 -89
rect 1413 -106 1435 -89
rect 1502 -106 1524 -89
<< locali >>
rect -1532 89 -1524 106
rect -1502 89 -1494 106
rect -1443 89 -1435 106
rect -1413 89 -1405 106
rect -1354 89 -1346 106
rect -1324 89 -1316 106
rect -1265 89 -1257 106
rect -1235 89 -1227 106
rect -1176 89 -1168 106
rect -1146 89 -1138 106
rect -1087 89 -1079 106
rect -1057 89 -1049 106
rect -998 89 -990 106
rect -968 89 -960 106
rect -909 89 -901 106
rect -879 89 -871 106
rect -820 89 -812 106
rect -790 89 -782 106
rect -731 89 -723 106
rect -701 89 -693 106
rect -642 89 -634 106
rect -612 89 -604 106
rect -553 89 -545 106
rect -523 89 -515 106
rect -464 89 -456 106
rect -434 89 -426 106
rect -375 89 -367 106
rect -345 89 -337 106
rect -286 89 -278 106
rect -256 89 -248 106
rect -197 89 -189 106
rect -167 89 -159 106
rect -108 89 -100 106
rect -78 89 -70 106
rect -19 89 -11 106
rect 11 89 19 106
rect 70 89 78 106
rect 100 89 108 106
rect 159 89 167 106
rect 189 89 197 106
rect 248 89 256 106
rect 278 89 286 106
rect 337 89 345 106
rect 367 89 375 106
rect 426 89 434 106
rect 456 89 464 106
rect 515 89 523 106
rect 545 89 553 106
rect 604 89 612 106
rect 634 89 642 106
rect 693 89 701 106
rect 723 89 731 106
rect 782 89 790 106
rect 812 89 820 106
rect 871 89 879 106
rect 901 89 909 106
rect 960 89 968 106
rect 990 89 998 106
rect 1049 89 1057 106
rect 1079 89 1087 106
rect 1138 89 1146 106
rect 1168 89 1176 106
rect 1227 89 1235 106
rect 1257 89 1265 106
rect 1316 89 1324 106
rect 1346 89 1354 106
rect 1405 89 1413 106
rect 1435 89 1443 106
rect 1494 89 1502 106
rect 1524 89 1532 106
rect -1566 64 -1549 72
rect -1566 -72 -1549 -64
rect -1477 64 -1460 72
rect -1477 -72 -1460 -64
rect -1388 64 -1371 72
rect -1388 -72 -1371 -64
rect -1299 64 -1282 72
rect -1299 -72 -1282 -64
rect -1210 64 -1193 72
rect -1210 -72 -1193 -64
rect -1121 64 -1104 72
rect -1121 -72 -1104 -64
rect -1032 64 -1015 72
rect -1032 -72 -1015 -64
rect -943 64 -926 72
rect -943 -72 -926 -64
rect -854 64 -837 72
rect -854 -72 -837 -64
rect -765 64 -748 72
rect -765 -72 -748 -64
rect -676 64 -659 72
rect -676 -72 -659 -64
rect -587 64 -570 72
rect -587 -72 -570 -64
rect -498 64 -481 72
rect -498 -72 -481 -64
rect -409 64 -392 72
rect -409 -72 -392 -64
rect -320 64 -303 72
rect -320 -72 -303 -64
rect -231 64 -214 72
rect -231 -72 -214 -64
rect -142 64 -125 72
rect -142 -72 -125 -64
rect -53 64 -36 72
rect -53 -72 -36 -64
rect 36 64 53 72
rect 36 -72 53 -64
rect 125 64 142 72
rect 125 -72 142 -64
rect 214 64 231 72
rect 214 -72 231 -64
rect 303 64 320 72
rect 303 -72 320 -64
rect 392 64 409 72
rect 392 -72 409 -64
rect 481 64 498 72
rect 481 -72 498 -64
rect 570 64 587 72
rect 570 -72 587 -64
rect 659 64 676 72
rect 659 -72 676 -64
rect 748 64 765 72
rect 748 -72 765 -64
rect 837 64 854 72
rect 837 -72 854 -64
rect 926 64 943 72
rect 926 -72 943 -64
rect 1015 64 1032 72
rect 1015 -72 1032 -64
rect 1104 64 1121 72
rect 1104 -72 1121 -64
rect 1193 64 1210 72
rect 1193 -72 1210 -64
rect 1282 64 1299 72
rect 1282 -72 1299 -64
rect 1371 64 1388 72
rect 1371 -72 1388 -64
rect 1460 64 1477 72
rect 1460 -72 1477 -64
rect 1549 64 1566 72
rect 1549 -72 1566 -64
rect -1532 -106 -1524 -89
rect -1502 -106 -1494 -89
rect -1443 -106 -1435 -89
rect -1413 -106 -1405 -89
rect -1354 -106 -1346 -89
rect -1324 -106 -1316 -89
rect -1265 -106 -1257 -89
rect -1235 -106 -1227 -89
rect -1176 -106 -1168 -89
rect -1146 -106 -1138 -89
rect -1087 -106 -1079 -89
rect -1057 -106 -1049 -89
rect -998 -106 -990 -89
rect -968 -106 -960 -89
rect -909 -106 -901 -89
rect -879 -106 -871 -89
rect -820 -106 -812 -89
rect -790 -106 -782 -89
rect -731 -106 -723 -89
rect -701 -106 -693 -89
rect -642 -106 -634 -89
rect -612 -106 -604 -89
rect -553 -106 -545 -89
rect -523 -106 -515 -89
rect -464 -106 -456 -89
rect -434 -106 -426 -89
rect -375 -106 -367 -89
rect -345 -106 -337 -89
rect -286 -106 -278 -89
rect -256 -106 -248 -89
rect -197 -106 -189 -89
rect -167 -106 -159 -89
rect -108 -106 -100 -89
rect -78 -106 -70 -89
rect -19 -106 -11 -89
rect 11 -106 19 -89
rect 70 -106 78 -89
rect 100 -106 108 -89
rect 159 -106 167 -89
rect 189 -106 197 -89
rect 248 -106 256 -89
rect 278 -106 286 -89
rect 337 -106 345 -89
rect 367 -106 375 -89
rect 426 -106 434 -89
rect 456 -106 464 -89
rect 515 -106 523 -89
rect 545 -106 553 -89
rect 604 -106 612 -89
rect 634 -106 642 -89
rect 693 -106 701 -89
rect 723 -106 731 -89
rect 782 -106 790 -89
rect 812 -106 820 -89
rect 871 -106 879 -89
rect 901 -106 909 -89
rect 960 -106 968 -89
rect 990 -106 998 -89
rect 1049 -106 1057 -89
rect 1079 -106 1087 -89
rect 1138 -106 1146 -89
rect 1168 -106 1176 -89
rect 1227 -106 1235 -89
rect 1257 -106 1265 -89
rect 1316 -106 1324 -89
rect 1346 -106 1354 -89
rect 1405 -106 1413 -89
rect 1435 -106 1443 -89
rect 1494 -106 1502 -89
rect 1524 -106 1532 -89
<< viali >>
rect -1524 89 -1502 106
rect -1435 89 -1413 106
rect -1346 89 -1324 106
rect -1257 89 -1235 106
rect -1168 89 -1146 106
rect -1079 89 -1057 106
rect -990 89 -968 106
rect -901 89 -879 106
rect -812 89 -790 106
rect -723 89 -701 106
rect -634 89 -612 106
rect -545 89 -523 106
rect -456 89 -434 106
rect -367 89 -345 106
rect -278 89 -256 106
rect -189 89 -167 106
rect -100 89 -78 106
rect -11 89 11 106
rect 78 89 100 106
rect 167 89 189 106
rect 256 89 278 106
rect 345 89 367 106
rect 434 89 456 106
rect 523 89 545 106
rect 612 89 634 106
rect 701 89 723 106
rect 790 89 812 106
rect 879 89 901 106
rect 968 89 990 106
rect 1057 89 1079 106
rect 1146 89 1168 106
rect 1235 89 1257 106
rect 1324 89 1346 106
rect 1413 89 1435 106
rect 1502 89 1524 106
rect -1566 -64 -1549 64
rect -1477 -64 -1460 64
rect -1388 -64 -1371 64
rect -1299 -64 -1282 64
rect -1210 -64 -1193 64
rect -1121 -64 -1104 64
rect -1032 -64 -1015 64
rect -943 -64 -926 64
rect -854 -64 -837 64
rect -765 -64 -748 64
rect -676 -64 -659 64
rect -587 -64 -570 64
rect -498 -64 -481 64
rect -409 -64 -392 64
rect -320 -64 -303 64
rect -231 -64 -214 64
rect -142 -64 -125 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 125 -64 142 64
rect 214 -64 231 64
rect 303 -64 320 64
rect 392 -64 409 64
rect 481 -64 498 64
rect 570 -64 587 64
rect 659 -64 676 64
rect 748 -64 765 64
rect 837 -64 854 64
rect 926 -64 943 64
rect 1015 -64 1032 64
rect 1104 -64 1121 64
rect 1193 -64 1210 64
rect 1282 -64 1299 64
rect 1371 -64 1388 64
rect 1460 -64 1477 64
rect 1549 -64 1566 64
rect -1524 -106 -1502 -89
rect -1435 -106 -1413 -89
rect -1346 -106 -1324 -89
rect -1257 -106 -1235 -89
rect -1168 -106 -1146 -89
rect -1079 -106 -1057 -89
rect -990 -106 -968 -89
rect -901 -106 -879 -89
rect -812 -106 -790 -89
rect -723 -106 -701 -89
rect -634 -106 -612 -89
rect -545 -106 -523 -89
rect -456 -106 -434 -89
rect -367 -106 -345 -89
rect -278 -106 -256 -89
rect -189 -106 -167 -89
rect -100 -106 -78 -89
rect -11 -106 11 -89
rect 78 -106 100 -89
rect 167 -106 189 -89
rect 256 -106 278 -89
rect 345 -106 367 -89
rect 434 -106 456 -89
rect 523 -106 545 -89
rect 612 -106 634 -89
rect 701 -106 723 -89
rect 790 -106 812 -89
rect 879 -106 901 -89
rect 968 -106 990 -89
rect 1057 -106 1079 -89
rect 1146 -106 1168 -89
rect 1235 -106 1257 -89
rect 1324 -106 1346 -89
rect 1413 -106 1435 -89
rect 1502 -106 1524 -89
<< metal1 >>
rect -1532 106 -1494 114
rect -1532 89 -1524 106
rect -1502 89 -1494 106
rect -1532 86 -1494 89
rect -1443 106 -1405 114
rect -1443 89 -1435 106
rect -1413 89 -1405 106
rect -1443 86 -1405 89
rect -1354 106 -1316 114
rect -1354 89 -1346 106
rect -1324 89 -1316 106
rect -1354 86 -1316 89
rect -1265 106 -1227 114
rect -1265 89 -1257 106
rect -1235 89 -1227 106
rect -1265 86 -1227 89
rect -1176 106 -1138 114
rect -1176 89 -1168 106
rect -1146 89 -1138 106
rect -1176 86 -1138 89
rect -1087 106 -1049 114
rect -1087 89 -1079 106
rect -1057 89 -1049 106
rect -1087 86 -1049 89
rect -998 106 -960 114
rect -998 89 -990 106
rect -968 89 -960 106
rect -998 86 -960 89
rect -909 106 -871 114
rect -909 89 -901 106
rect -879 89 -871 106
rect -909 86 -871 89
rect -820 106 -782 114
rect -820 89 -812 106
rect -790 89 -782 106
rect -820 86 -782 89
rect -731 106 -693 114
rect -731 89 -723 106
rect -701 89 -693 106
rect -731 86 -693 89
rect -642 106 -604 114
rect -642 89 -634 106
rect -612 89 -604 106
rect -642 86 -604 89
rect -553 106 -515 114
rect -553 89 -545 106
rect -523 89 -515 106
rect -553 86 -515 89
rect -464 106 -426 114
rect -464 89 -456 106
rect -434 89 -426 106
rect -464 86 -426 89
rect -375 106 -337 114
rect -375 89 -367 106
rect -345 89 -337 106
rect -375 86 -337 89
rect -286 106 -248 114
rect -286 89 -278 106
rect -256 89 -248 106
rect -286 86 -248 89
rect -197 106 -159 114
rect -197 89 -189 106
rect -167 89 -159 106
rect -197 86 -159 89
rect -108 106 -70 114
rect -108 89 -100 106
rect -78 89 -70 106
rect -108 86 -70 89
rect -19 106 19 114
rect -19 89 -11 106
rect 11 89 19 106
rect -19 86 19 89
rect 70 106 108 114
rect 70 89 78 106
rect 100 89 108 106
rect 70 86 108 89
rect 159 106 197 114
rect 159 89 167 106
rect 189 89 197 106
rect 159 86 197 89
rect 248 106 286 114
rect 248 89 256 106
rect 278 89 286 106
rect 248 86 286 89
rect 337 106 375 114
rect 337 89 345 106
rect 367 89 375 106
rect 337 86 375 89
rect 426 106 464 114
rect 426 89 434 106
rect 456 89 464 106
rect 426 86 464 89
rect 515 106 553 114
rect 515 89 523 106
rect 545 89 553 106
rect 515 86 553 89
rect 604 106 642 114
rect 604 89 612 106
rect 634 89 642 106
rect 604 86 642 89
rect 693 106 731 114
rect 693 89 701 106
rect 723 89 731 106
rect 693 86 731 89
rect 782 106 820 114
rect 782 89 790 106
rect 812 89 820 106
rect 782 86 820 89
rect 871 106 909 114
rect 871 89 879 106
rect 901 89 909 106
rect 871 86 909 89
rect 960 106 998 114
rect 960 89 968 106
rect 990 89 998 106
rect 960 86 998 89
rect 1049 106 1087 114
rect 1049 89 1057 106
rect 1079 89 1087 106
rect 1049 86 1087 89
rect 1138 106 1176 114
rect 1138 89 1146 106
rect 1168 89 1176 106
rect 1138 86 1176 89
rect 1227 106 1265 114
rect 1227 89 1235 106
rect 1257 89 1265 106
rect 1227 86 1265 89
rect 1316 106 1354 114
rect 1316 89 1324 106
rect 1346 89 1354 106
rect 1316 86 1354 89
rect 1405 106 1443 114
rect 1405 89 1413 106
rect 1435 89 1443 106
rect 1405 86 1443 89
rect 1494 106 1532 114
rect 1494 89 1502 106
rect 1524 89 1532 106
rect 1494 86 1532 89
rect -1569 64 -1546 70
rect -1569 -64 -1566 64
rect -1549 -64 -1546 64
rect -1569 -70 -1546 -64
rect -1480 64 -1457 70
rect -1480 -64 -1477 64
rect -1460 -64 -1457 64
rect -1480 -70 -1457 -64
rect -1391 64 -1368 70
rect -1391 -64 -1388 64
rect -1371 -64 -1368 64
rect -1391 -70 -1368 -64
rect -1302 64 -1279 70
rect -1302 -64 -1299 64
rect -1282 -64 -1279 64
rect -1302 -70 -1279 -64
rect -1213 64 -1190 70
rect -1213 -64 -1210 64
rect -1193 -64 -1190 64
rect -1213 -70 -1190 -64
rect -1124 64 -1101 70
rect -1124 -64 -1121 64
rect -1104 -64 -1101 64
rect -1124 -70 -1101 -64
rect -1035 64 -1012 70
rect -1035 -64 -1032 64
rect -1015 -64 -1012 64
rect -1035 -70 -1012 -64
rect -946 64 -923 70
rect -946 -64 -943 64
rect -926 -64 -923 64
rect -946 -70 -923 -64
rect -857 64 -834 70
rect -857 -64 -854 64
rect -837 -64 -834 64
rect -857 -70 -834 -64
rect -768 64 -745 70
rect -768 -64 -765 64
rect -748 -64 -745 64
rect -768 -70 -745 -64
rect -679 64 -656 70
rect -679 -64 -676 64
rect -659 -64 -656 64
rect -679 -70 -656 -64
rect -590 64 -567 70
rect -590 -64 -587 64
rect -570 -64 -567 64
rect -590 -70 -567 -64
rect -501 64 -478 70
rect -501 -64 -498 64
rect -481 -64 -478 64
rect -501 -70 -478 -64
rect -412 64 -389 70
rect -412 -64 -409 64
rect -392 -64 -389 64
rect -412 -70 -389 -64
rect -323 64 -300 70
rect -323 -64 -320 64
rect -303 -64 -300 64
rect -323 -70 -300 -64
rect -234 64 -211 70
rect -234 -64 -231 64
rect -214 -64 -211 64
rect -234 -70 -211 -64
rect -145 64 -122 70
rect -145 -64 -142 64
rect -125 -64 -122 64
rect -145 -70 -122 -64
rect -56 64 -33 70
rect -56 -64 -53 64
rect -36 -64 -33 64
rect -56 -70 -33 -64
rect 33 64 56 70
rect 33 -64 36 64
rect 53 -64 56 64
rect 33 -70 56 -64
rect 122 64 145 70
rect 122 -64 125 64
rect 142 -64 145 64
rect 122 -70 145 -64
rect 211 64 234 70
rect 211 -64 214 64
rect 231 -64 234 64
rect 211 -70 234 -64
rect 300 64 323 70
rect 300 -64 303 64
rect 320 -64 323 64
rect 300 -70 323 -64
rect 389 64 412 70
rect 389 -64 392 64
rect 409 -64 412 64
rect 389 -70 412 -64
rect 478 64 501 70
rect 478 -64 481 64
rect 498 -64 501 64
rect 478 -70 501 -64
rect 567 64 590 70
rect 567 -64 570 64
rect 587 -64 590 64
rect 567 -70 590 -64
rect 656 64 679 70
rect 656 -64 659 64
rect 676 -64 679 64
rect 656 -70 679 -64
rect 745 64 768 70
rect 745 -64 748 64
rect 765 -64 768 64
rect 745 -70 768 -64
rect 834 64 857 70
rect 834 -64 837 64
rect 854 -64 857 64
rect 834 -70 857 -64
rect 923 64 946 70
rect 923 -64 926 64
rect 943 -64 946 64
rect 923 -70 946 -64
rect 1012 64 1035 70
rect 1012 -64 1015 64
rect 1032 -64 1035 64
rect 1012 -70 1035 -64
rect 1101 64 1124 70
rect 1101 -64 1104 64
rect 1121 -64 1124 64
rect 1101 -70 1124 -64
rect 1190 64 1213 70
rect 1190 -64 1193 64
rect 1210 -64 1213 64
rect 1190 -70 1213 -64
rect 1279 64 1302 70
rect 1279 -64 1282 64
rect 1299 -64 1302 64
rect 1279 -70 1302 -64
rect 1368 64 1391 70
rect 1368 -64 1371 64
rect 1388 -64 1391 64
rect 1368 -70 1391 -64
rect 1457 64 1480 70
rect 1457 -64 1460 64
rect 1477 -64 1480 64
rect 1457 -70 1480 -64
rect 1546 64 1569 70
rect 1546 -64 1549 64
rect 1566 -64 1569 64
rect 1546 -70 1569 -64
rect -1532 -89 -1494 -86
rect -1532 -106 -1524 -89
rect -1502 -106 -1494 -89
rect -1532 -114 -1494 -106
rect -1443 -89 -1405 -86
rect -1443 -106 -1435 -89
rect -1413 -106 -1405 -89
rect -1443 -114 -1405 -106
rect -1354 -89 -1316 -86
rect -1354 -106 -1346 -89
rect -1324 -106 -1316 -89
rect -1354 -114 -1316 -106
rect -1265 -89 -1227 -86
rect -1265 -106 -1257 -89
rect -1235 -106 -1227 -89
rect -1265 -114 -1227 -106
rect -1176 -89 -1138 -86
rect -1176 -106 -1168 -89
rect -1146 -106 -1138 -89
rect -1176 -114 -1138 -106
rect -1087 -89 -1049 -86
rect -1087 -106 -1079 -89
rect -1057 -106 -1049 -89
rect -1087 -114 -1049 -106
rect -998 -89 -960 -86
rect -998 -106 -990 -89
rect -968 -106 -960 -89
rect -998 -114 -960 -106
rect -909 -89 -871 -86
rect -909 -106 -901 -89
rect -879 -106 -871 -89
rect -909 -114 -871 -106
rect -820 -89 -782 -86
rect -820 -106 -812 -89
rect -790 -106 -782 -89
rect -820 -114 -782 -106
rect -731 -89 -693 -86
rect -731 -106 -723 -89
rect -701 -106 -693 -89
rect -731 -114 -693 -106
rect -642 -89 -604 -86
rect -642 -106 -634 -89
rect -612 -106 -604 -89
rect -642 -114 -604 -106
rect -553 -89 -515 -86
rect -553 -106 -545 -89
rect -523 -106 -515 -89
rect -553 -114 -515 -106
rect -464 -89 -426 -86
rect -464 -106 -456 -89
rect -434 -106 -426 -89
rect -464 -114 -426 -106
rect -375 -89 -337 -86
rect -375 -106 -367 -89
rect -345 -106 -337 -89
rect -375 -114 -337 -106
rect -286 -89 -248 -86
rect -286 -106 -278 -89
rect -256 -106 -248 -89
rect -286 -114 -248 -106
rect -197 -89 -159 -86
rect -197 -106 -189 -89
rect -167 -106 -159 -89
rect -197 -114 -159 -106
rect -108 -89 -70 -86
rect -108 -106 -100 -89
rect -78 -106 -70 -89
rect -108 -114 -70 -106
rect -19 -89 19 -86
rect -19 -106 -11 -89
rect 11 -106 19 -89
rect -19 -114 19 -106
rect 70 -89 108 -86
rect 70 -106 78 -89
rect 100 -106 108 -89
rect 70 -114 108 -106
rect 159 -89 197 -86
rect 159 -106 167 -89
rect 189 -106 197 -89
rect 159 -114 197 -106
rect 248 -89 286 -86
rect 248 -106 256 -89
rect 278 -106 286 -89
rect 248 -114 286 -106
rect 337 -89 375 -86
rect 337 -106 345 -89
rect 367 -106 375 -89
rect 337 -114 375 -106
rect 426 -89 464 -86
rect 426 -106 434 -89
rect 456 -106 464 -89
rect 426 -114 464 -106
rect 515 -89 553 -86
rect 515 -106 523 -89
rect 545 -106 553 -89
rect 515 -114 553 -106
rect 604 -89 642 -86
rect 604 -106 612 -89
rect 634 -106 642 -89
rect 604 -114 642 -106
rect 693 -89 731 -86
rect 693 -106 701 -89
rect 723 -106 731 -89
rect 693 -114 731 -106
rect 782 -89 820 -86
rect 782 -106 790 -89
rect 812 -106 820 -89
rect 782 -114 820 -106
rect 871 -89 909 -86
rect 871 -106 879 -89
rect 901 -106 909 -89
rect 871 -114 909 -106
rect 960 -89 998 -86
rect 960 -106 968 -89
rect 990 -106 998 -89
rect 960 -114 998 -106
rect 1049 -89 1087 -86
rect 1049 -106 1057 -89
rect 1079 -106 1087 -89
rect 1049 -114 1087 -106
rect 1138 -89 1176 -86
rect 1138 -106 1146 -89
rect 1168 -106 1176 -89
rect 1138 -114 1176 -106
rect 1227 -89 1265 -86
rect 1227 -106 1235 -89
rect 1257 -106 1265 -89
rect 1227 -114 1265 -106
rect 1316 -89 1354 -86
rect 1316 -106 1324 -89
rect 1346 -106 1354 -89
rect 1316 -114 1354 -106
rect 1405 -89 1443 -86
rect 1405 -106 1413 -89
rect 1435 -106 1443 -89
rect 1405 -114 1443 -106
rect 1494 -89 1532 -86
rect 1494 -106 1502 -89
rect 1524 -106 1532 -89
rect 1494 -114 1532 -106
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 35 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
