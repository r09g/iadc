magic
tech sky130A
magscale 1 2
timestamp 1654865385
<< error_p >>
rect -1631 -140 -1573 140
rect -1453 -140 -1395 140
rect -1275 -140 -1217 140
rect -1097 -140 -1039 140
rect -919 -140 -861 140
rect -741 -140 -683 140
rect -563 -140 -505 140
rect -385 -140 -327 140
rect -207 -140 -149 140
rect -29 -140 29 140
rect 149 -140 207 140
rect 327 -140 385 140
rect 505 -140 563 140
rect 683 -140 741 140
rect 861 -140 919 140
rect 1039 -140 1097 140
rect 1217 -140 1275 140
rect 1395 -140 1453 140
rect 1573 -140 1631 140
<< nmos >>
rect -1573 -140 -1453 140
rect -1395 -140 -1275 140
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
rect 1275 -140 1395 140
rect 1453 -140 1573 140
<< ndiff >>
rect -1631 128 -1573 140
rect -1631 -128 -1619 128
rect -1585 -128 -1573 128
rect -1631 -140 -1573 -128
rect -1453 128 -1395 140
rect -1453 -128 -1441 128
rect -1407 -128 -1395 128
rect -1453 -140 -1395 -128
rect -1275 128 -1217 140
rect -1275 -128 -1263 128
rect -1229 -128 -1217 128
rect -1275 -140 -1217 -128
rect -1097 128 -1039 140
rect -1097 -128 -1085 128
rect -1051 -128 -1039 128
rect -1097 -140 -1039 -128
rect -919 128 -861 140
rect -919 -128 -907 128
rect -873 -128 -861 128
rect -919 -140 -861 -128
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
rect 861 128 919 140
rect 861 -128 873 128
rect 907 -128 919 128
rect 861 -140 919 -128
rect 1039 128 1097 140
rect 1039 -128 1051 128
rect 1085 -128 1097 128
rect 1039 -140 1097 -128
rect 1217 128 1275 140
rect 1217 -128 1229 128
rect 1263 -128 1275 128
rect 1217 -140 1275 -128
rect 1395 128 1453 140
rect 1395 -128 1407 128
rect 1441 -128 1453 128
rect 1395 -140 1453 -128
rect 1573 128 1631 140
rect 1573 -128 1585 128
rect 1619 -128 1631 128
rect 1573 -140 1631 -128
<< ndiffc >>
rect -1619 -128 -1585 128
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
rect 1585 -128 1619 128
<< poly >>
rect -1555 212 -1471 228
rect -1555 194 -1539 212
rect -1573 178 -1539 194
rect -1487 194 -1471 212
rect -1377 212 -1293 228
rect -1377 194 -1361 212
rect -1487 178 -1453 194
rect -1573 140 -1453 178
rect -1395 178 -1361 194
rect -1309 194 -1293 212
rect -1199 212 -1115 228
rect -1199 194 -1183 212
rect -1309 178 -1275 194
rect -1395 140 -1275 178
rect -1217 178 -1183 194
rect -1131 194 -1115 212
rect -1021 212 -937 228
rect -1021 194 -1005 212
rect -1131 178 -1097 194
rect -1217 140 -1097 178
rect -1039 178 -1005 194
rect -953 194 -937 212
rect -843 212 -759 228
rect -843 194 -827 212
rect -953 178 -919 194
rect -1039 140 -919 178
rect -861 178 -827 194
rect -775 194 -759 212
rect -665 212 -581 228
rect -665 194 -649 212
rect -775 178 -741 194
rect -861 140 -741 178
rect -683 178 -649 194
rect -597 194 -581 212
rect -487 212 -403 228
rect -487 194 -471 212
rect -597 178 -563 194
rect -683 140 -563 178
rect -505 178 -471 194
rect -419 194 -403 212
rect -309 212 -225 228
rect -309 194 -293 212
rect -419 178 -385 194
rect -505 140 -385 178
rect -327 178 -293 194
rect -241 194 -225 212
rect -131 212 -47 228
rect -131 194 -115 212
rect -241 178 -207 194
rect -327 140 -207 178
rect -149 178 -115 194
rect -63 194 -47 212
rect 47 212 131 228
rect 47 194 63 212
rect -63 178 -29 194
rect -149 140 -29 178
rect 29 178 63 194
rect 115 194 131 212
rect 225 212 309 228
rect 225 194 241 212
rect 115 178 149 194
rect 29 140 149 178
rect 207 178 241 194
rect 293 194 309 212
rect 403 212 487 228
rect 403 194 419 212
rect 293 178 327 194
rect 207 140 327 178
rect 385 178 419 194
rect 471 194 487 212
rect 581 212 665 228
rect 581 194 597 212
rect 471 178 505 194
rect 385 140 505 178
rect 563 178 597 194
rect 649 194 665 212
rect 759 212 843 228
rect 759 194 775 212
rect 649 178 683 194
rect 563 140 683 178
rect 741 178 775 194
rect 827 194 843 212
rect 937 212 1021 228
rect 937 194 953 212
rect 827 178 861 194
rect 741 140 861 178
rect 919 178 953 194
rect 1005 194 1021 212
rect 1115 212 1199 228
rect 1115 194 1131 212
rect 1005 178 1039 194
rect 919 140 1039 178
rect 1097 178 1131 194
rect 1183 194 1199 212
rect 1293 212 1377 228
rect 1293 194 1309 212
rect 1183 178 1217 194
rect 1097 140 1217 178
rect 1275 178 1309 194
rect 1361 194 1377 212
rect 1471 212 1555 228
rect 1471 194 1487 212
rect 1361 178 1395 194
rect 1275 140 1395 178
rect 1453 178 1487 194
rect 1539 194 1555 212
rect 1539 178 1573 194
rect 1453 140 1573 178
rect -1573 -178 -1453 -140
rect -1573 -194 -1539 -178
rect -1555 -212 -1539 -194
rect -1487 -194 -1453 -178
rect -1395 -178 -1275 -140
rect -1395 -194 -1361 -178
rect -1487 -212 -1471 -194
rect -1555 -228 -1471 -212
rect -1377 -212 -1361 -194
rect -1309 -194 -1275 -178
rect -1217 -178 -1097 -140
rect -1217 -194 -1183 -178
rect -1309 -212 -1293 -194
rect -1377 -228 -1293 -212
rect -1199 -212 -1183 -194
rect -1131 -194 -1097 -178
rect -1039 -178 -919 -140
rect -1039 -194 -1005 -178
rect -1131 -212 -1115 -194
rect -1199 -228 -1115 -212
rect -1021 -212 -1005 -194
rect -953 -194 -919 -178
rect -861 -178 -741 -140
rect -861 -194 -827 -178
rect -953 -212 -937 -194
rect -1021 -228 -937 -212
rect -843 -212 -827 -194
rect -775 -194 -741 -178
rect -683 -178 -563 -140
rect -683 -194 -649 -178
rect -775 -212 -759 -194
rect -843 -228 -759 -212
rect -665 -212 -649 -194
rect -597 -194 -563 -178
rect -505 -178 -385 -140
rect -505 -194 -471 -178
rect -597 -212 -581 -194
rect -665 -228 -581 -212
rect -487 -212 -471 -194
rect -419 -194 -385 -178
rect -327 -178 -207 -140
rect -327 -194 -293 -178
rect -419 -212 -403 -194
rect -487 -228 -403 -212
rect -309 -212 -293 -194
rect -241 -194 -207 -178
rect -149 -178 -29 -140
rect -149 -194 -115 -178
rect -241 -212 -225 -194
rect -309 -228 -225 -212
rect -131 -212 -115 -194
rect -63 -194 -29 -178
rect 29 -178 149 -140
rect 29 -194 63 -178
rect -63 -212 -47 -194
rect -131 -228 -47 -212
rect 47 -212 63 -194
rect 115 -194 149 -178
rect 207 -178 327 -140
rect 207 -194 241 -178
rect 115 -212 131 -194
rect 47 -228 131 -212
rect 225 -212 241 -194
rect 293 -194 327 -178
rect 385 -178 505 -140
rect 385 -194 419 -178
rect 293 -212 309 -194
rect 225 -228 309 -212
rect 403 -212 419 -194
rect 471 -194 505 -178
rect 563 -178 683 -140
rect 563 -194 597 -178
rect 471 -212 487 -194
rect 403 -228 487 -212
rect 581 -212 597 -194
rect 649 -194 683 -178
rect 741 -178 861 -140
rect 741 -194 775 -178
rect 649 -212 665 -194
rect 581 -228 665 -212
rect 759 -212 775 -194
rect 827 -194 861 -178
rect 919 -178 1039 -140
rect 919 -194 953 -178
rect 827 -212 843 -194
rect 759 -228 843 -212
rect 937 -212 953 -194
rect 1005 -194 1039 -178
rect 1097 -178 1217 -140
rect 1097 -194 1131 -178
rect 1005 -212 1021 -194
rect 937 -228 1021 -212
rect 1115 -212 1131 -194
rect 1183 -194 1217 -178
rect 1275 -178 1395 -140
rect 1275 -194 1309 -178
rect 1183 -212 1199 -194
rect 1115 -228 1199 -212
rect 1293 -212 1309 -194
rect 1361 -194 1395 -178
rect 1453 -178 1573 -140
rect 1453 -194 1487 -178
rect 1361 -212 1377 -194
rect 1293 -228 1377 -212
rect 1471 -212 1487 -194
rect 1539 -194 1573 -178
rect 1539 -212 1555 -194
rect 1471 -228 1555 -212
<< polycont >>
rect -1539 178 -1487 212
rect -1361 178 -1309 212
rect -1183 178 -1131 212
rect -1005 178 -953 212
rect -827 178 -775 212
rect -649 178 -597 212
rect -471 178 -419 212
rect -293 178 -241 212
rect -115 178 -63 212
rect 63 178 115 212
rect 241 178 293 212
rect 419 178 471 212
rect 597 178 649 212
rect 775 178 827 212
rect 953 178 1005 212
rect 1131 178 1183 212
rect 1309 178 1361 212
rect 1487 178 1539 212
rect -1539 -212 -1487 -178
rect -1361 -212 -1309 -178
rect -1183 -212 -1131 -178
rect -1005 -212 -953 -178
rect -827 -212 -775 -178
rect -649 -212 -597 -178
rect -471 -212 -419 -178
rect -293 -212 -241 -178
rect -115 -212 -63 -178
rect 63 -212 115 -178
rect 241 -212 293 -178
rect 419 -212 471 -178
rect 597 -212 649 -178
rect 775 -212 827 -178
rect 953 -212 1005 -178
rect 1131 -212 1183 -178
rect 1309 -212 1361 -178
rect 1487 -212 1539 -178
<< locali >>
rect -1619 178 -1539 212
rect -1487 178 -1471 212
rect -1377 178 -1361 212
rect -1309 178 -1293 212
rect -1199 178 -1183 212
rect -1131 178 -1115 212
rect -1021 178 -1005 212
rect -953 178 -937 212
rect -843 178 -827 212
rect -775 178 -759 212
rect -665 178 -649 212
rect -597 178 -581 212
rect -487 178 -471 212
rect -419 178 -403 212
rect -309 178 -293 212
rect -241 178 -225 212
rect -131 178 -115 212
rect -63 178 -47 212
rect 47 178 63 212
rect 115 178 131 212
rect 225 178 241 212
rect 293 178 309 212
rect 403 178 419 212
rect 471 178 487 212
rect 581 178 597 212
rect 649 178 665 212
rect 759 178 775 212
rect 827 178 843 212
rect 937 178 953 212
rect 1005 178 1021 212
rect 1115 178 1131 212
rect 1183 178 1199 212
rect 1293 178 1309 212
rect 1361 178 1377 212
rect 1471 178 1487 212
rect 1539 178 1619 212
rect -1619 128 -1585 178
rect -1619 -178 -1585 -128
rect -1441 128 -1407 144
rect -1441 -144 -1407 -128
rect -1263 128 -1229 144
rect -1263 -144 -1229 -128
rect -1085 128 -1051 144
rect -1085 -144 -1051 -128
rect -907 128 -873 144
rect -907 -144 -873 -128
rect -729 128 -695 144
rect -729 -144 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 144
rect 695 -144 729 -128
rect 873 128 907 144
rect 873 -144 907 -128
rect 1051 128 1085 144
rect 1051 -144 1085 -128
rect 1229 128 1263 144
rect 1229 -144 1263 -128
rect 1407 128 1441 144
rect 1407 -144 1441 -128
rect 1585 128 1619 178
rect 1585 -178 1619 -128
rect -1619 -212 -1539 -178
rect -1487 -212 -1471 -178
rect -1377 -212 -1361 -178
rect -1309 -212 -1293 -178
rect -1199 -212 -1183 -178
rect -1131 -212 -1115 -178
rect -1021 -212 -1005 -178
rect -953 -212 -937 -178
rect -843 -212 -827 -178
rect -775 -212 -759 -178
rect -665 -212 -649 -178
rect -597 -212 -581 -178
rect -487 -212 -471 -178
rect -419 -212 -403 -178
rect -309 -212 -293 -178
rect -241 -212 -225 -178
rect -131 -212 -115 -178
rect -63 -212 -47 -178
rect 47 -212 63 -178
rect 115 -212 131 -178
rect 225 -212 241 -178
rect 293 -212 309 -178
rect 403 -212 419 -178
rect 471 -212 487 -178
rect 581 -212 597 -178
rect 649 -212 665 -178
rect 759 -212 775 -178
rect 827 -212 843 -178
rect 937 -212 953 -178
rect 1005 -212 1021 -178
rect 1115 -212 1131 -178
rect 1183 -212 1199 -178
rect 1293 -212 1309 -178
rect 1361 -212 1377 -178
rect 1471 -212 1487 -178
rect 1539 -212 1619 -178
<< viali >>
rect -1361 178 -1309 212
rect -1183 178 -1131 212
rect -1005 178 -953 212
rect -827 178 -775 212
rect -649 178 -597 212
rect -471 178 -419 212
rect -293 178 -241 212
rect -115 178 -63 212
rect 63 178 115 212
rect 241 178 293 212
rect 419 178 471 212
rect 597 178 649 212
rect 775 178 827 212
rect 953 178 1005 212
rect 1131 178 1183 212
rect 1309 178 1361 212
rect -1361 -212 -1309 -178
rect -1183 -212 -1131 -178
rect -1005 -212 -953 -178
rect -827 -212 -775 -178
rect -649 -212 -597 -178
rect -471 -212 -419 -178
rect -293 -212 -241 -178
rect -115 -212 -63 -178
rect 63 -212 115 -178
rect 241 -212 293 -178
rect 419 -212 471 -178
rect 597 -212 649 -178
rect 775 -212 827 -178
rect 953 -212 1005 -178
rect 1131 -212 1183 -178
rect 1309 -212 1361 -178
<< metal1 >>
rect -1373 212 -1297 218
rect -1373 178 -1361 212
rect -1309 178 -1297 212
rect -1373 172 -1297 178
rect -1195 212 -1119 218
rect -1195 178 -1183 212
rect -1131 178 -1119 212
rect -1195 172 -1119 178
rect -1017 212 -941 218
rect -1017 178 -1005 212
rect -953 178 -941 212
rect -1017 172 -941 178
rect -839 212 -763 218
rect -839 178 -827 212
rect -775 178 -763 212
rect -839 172 -763 178
rect -661 212 -585 218
rect -661 178 -649 212
rect -597 178 -585 212
rect -661 172 -585 178
rect -483 212 -407 218
rect -483 178 -471 212
rect -419 178 -407 212
rect -483 172 -407 178
rect -305 212 -229 218
rect -305 178 -293 212
rect -241 178 -229 212
rect -305 172 -229 178
rect -127 212 -51 218
rect -127 178 -115 212
rect -63 178 -51 212
rect -127 172 -51 178
rect 51 212 127 218
rect 51 178 63 212
rect 115 178 127 212
rect 51 172 127 178
rect 229 212 305 218
rect 229 178 241 212
rect 293 178 305 212
rect 229 172 305 178
rect 407 212 483 218
rect 407 178 419 212
rect 471 178 483 212
rect 407 172 483 178
rect 585 212 661 218
rect 585 178 597 212
rect 649 178 661 212
rect 585 172 661 178
rect 763 212 839 218
rect 763 178 775 212
rect 827 178 839 212
rect 763 172 839 178
rect 941 212 1017 218
rect 941 178 953 212
rect 1005 178 1017 212
rect 941 172 1017 178
rect 1119 212 1195 218
rect 1119 178 1131 212
rect 1183 178 1195 212
rect 1119 172 1195 178
rect 1297 212 1373 218
rect 1297 178 1309 212
rect 1361 178 1373 212
rect 1297 172 1373 178
rect -1373 -178 -1297 -172
rect -1373 -212 -1361 -178
rect -1309 -212 -1297 -178
rect -1373 -218 -1297 -212
rect -1195 -178 -1119 -172
rect -1195 -212 -1183 -178
rect -1131 -212 -1119 -178
rect -1195 -218 -1119 -212
rect -1017 -178 -941 -172
rect -1017 -212 -1005 -178
rect -953 -212 -941 -178
rect -1017 -218 -941 -212
rect -839 -178 -763 -172
rect -839 -212 -827 -178
rect -775 -212 -763 -178
rect -839 -218 -763 -212
rect -661 -178 -585 -172
rect -661 -212 -649 -178
rect -597 -212 -585 -178
rect -661 -218 -585 -212
rect -483 -178 -407 -172
rect -483 -212 -471 -178
rect -419 -212 -407 -178
rect -483 -218 -407 -212
rect -305 -178 -229 -172
rect -305 -212 -293 -178
rect -241 -212 -229 -178
rect -305 -218 -229 -212
rect -127 -178 -51 -172
rect -127 -212 -115 -178
rect -63 -212 -51 -178
rect -127 -218 -51 -212
rect 51 -178 127 -172
rect 51 -212 63 -178
rect 115 -212 127 -178
rect 51 -218 127 -212
rect 229 -178 305 -172
rect 229 -212 241 -178
rect 293 -212 305 -178
rect 229 -218 305 -212
rect 407 -178 483 -172
rect 407 -212 419 -178
rect 471 -212 483 -178
rect 407 -218 483 -212
rect 585 -178 661 -172
rect 585 -212 597 -178
rect 649 -212 661 -178
rect 585 -218 661 -212
rect 763 -178 839 -172
rect 763 -212 775 -178
rect 827 -212 839 -178
rect 763 -218 839 -212
rect 941 -178 1017 -172
rect 941 -212 953 -178
rect 1005 -212 1017 -178
rect 941 -218 1017 -212
rect 1119 -178 1195 -172
rect 1119 -212 1131 -178
rect 1183 -212 1195 -178
rect 1119 -218 1195 -212
rect 1297 -178 1373 -172
rect 1297 -212 1309 -178
rect 1361 -212 1373 -178
rect 1297 -218 1373 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 18 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
