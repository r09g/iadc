* gold
.include "../sky130_fd_sc_hd.spice"

.subckt clock clk p2d_b p2d p2_b p2 p1d_b p1d p1_b p1 Ad_b Ad A_b A Bd_b Bd B_b B VDD VSS
x2 latch_out clk VSS VSS VDD VDD net1 sky130_fd_sc_hd__nand2_1
x3 net3 net6 VSS VSS VDD VDD net4 sky130_fd_sc_hd__nand2_1
x4 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__clkinv_4
x6 net2 VSS VSS VDD VDD net34 sky130_fd_sc_hd__clkinv_1
x9 net4 VSS VSS VDD VDD net5 sky130_fd_sc_hd__clkinv_4
x11 net5 VSS VSS VDD VDD net35 sky130_fd_sc_hd__clkinv_1
x1 clk VSS VSS VDD VDD net3 sky130_fd_sc_hd__clkinv_1
x20 net36 VSS VSS VDD VDD latch_in sky130_fd_sc_hd__clkdlybuf4s50_1
x21 net37 VSS VSS VDD VDD net6 sky130_fd_sc_hd__clkdlybuf4s50_1
x22 net34 VSS VSS VDD VDD net38 sky130_fd_sc_hd__clkdlybuf4s50_1
x25 net35 VSS VSS VDD VDD net39 sky130_fd_sc_hd__clkdlybuf4s50_1
x7 net40 VSS VSS VDD VDD net36 sky130_fd_sc_hd__clkdlybuf4s50_1
x12 net41 VSS VSS VDD VDD net37 sky130_fd_sc_hd__clkdlybuf4s50_1
x14 net38 VSS VSS VDD VDD net42 sky130_fd_sc_hd__clkdlybuf4s50_1
x15 net39 VSS VSS VDD VDD net43 sky130_fd_sc_hd__clkdlybuf4s50_1
x16 net44 VSS VSS VDD VDD net40 sky130_fd_sc_hd__clkdlybuf4s50_1
x17 net45 VSS VSS VDD VDD net41 sky130_fd_sc_hd__clkdlybuf4s50_1
x18 net42 VSS VSS VDD VDD net46 sky130_fd_sc_hd__clkdlybuf4s50_1
x19 net43 VSS VSS VDD VDD net47 sky130_fd_sc_hd__clkdlybuf4s50_1
x23 net48 VSS VSS VDD VDD net44 sky130_fd_sc_hd__clkdlybuf4s50_1
x24 net49 VSS VSS VDD VDD net45 sky130_fd_sc_hd__clkdlybuf4s50_1
x26 net46 VSS VSS VDD VDD net7 sky130_fd_sc_hd__clkdlybuf4s50_1
x27 net47 VSS VSS VDD VDD net8 sky130_fd_sc_hd__clkdlybuf4s50_1
x28 net50 VSS VSS VDD VDD net48 sky130_fd_sc_hd__clkdlybuf4s50_1
x29 net51 VSS VSS VDD VDD net49 sky130_fd_sc_hd__clkdlybuf4s50_1
x32 net52 VSS VSS VDD VDD net50 sky130_fd_sc_hd__clkdlybuf4s50_1
x33 net53 VSS VSS VDD VDD net51 sky130_fd_sc_hd__clkdlybuf4s50_1
x36 net54 VSS VSS VDD VDD net52 sky130_fd_sc_hd__clkdlybuf4s50_1
x37 net55 VSS VSS VDD VDD net53 sky130_fd_sc_hd__clkdlybuf4s50_1
x40 net56 VSS VSS VDD VDD net54 sky130_fd_sc_hd__clkdlybuf4s50_1
x41 net57 VSS VSS VDD VDD net55 sky130_fd_sc_hd__clkdlybuf4s50_1
x44 net58 VSS VSS VDD VDD net56 sky130_fd_sc_hd__clkdlybuf4s50_1
x45 net59 VSS VSS VDD VDD net57 sky130_fd_sc_hd__clkdlybuf4s50_1
x48 net60 VSS VSS VDD VDD net58 sky130_fd_sc_hd__clkdlybuf4s50_1
x49 net61 VSS VSS VDD VDD net59 sky130_fd_sc_hd__clkdlybuf4s50_1
x52 net62 VSS VSS VDD VDD net60 sky130_fd_sc_hd__clkdlybuf4s50_1
x53 net63 VSS VSS VDD VDD net61 sky130_fd_sc_hd__clkdlybuf4s50_1
x56 net64 VSS VSS VDD VDD net62 sky130_fd_sc_hd__clkdlybuf4s50_1
x57 net65 VSS VSS VDD VDD net63 sky130_fd_sc_hd__clkdlybuf4s50_1
x60 net66 VSS VSS VDD VDD net64 sky130_fd_sc_hd__clkdlybuf4s50_1
x61 net67 VSS VSS VDD VDD net65 sky130_fd_sc_hd__clkdlybuf4s50_1
x64 net68 VSS VSS VDD VDD net66 sky130_fd_sc_hd__clkdlybuf4s50_1
x65 net69 VSS VSS VDD VDD net67 sky130_fd_sc_hd__clkdlybuf4s50_1
x68 net70 VSS VSS VDD VDD net68 sky130_fd_sc_hd__clkdlybuf4s50_1
x69 net71 VSS VSS VDD VDD net69 sky130_fd_sc_hd__clkdlybuf4s50_1
x72 net72 VSS VSS VDD VDD net70 sky130_fd_sc_hd__clkdlybuf4s50_1
x73 net73 VSS VSS VDD VDD net71 sky130_fd_sc_hd__clkdlybuf4s50_1
x76 net74 VSS VSS VDD VDD net72 sky130_fd_sc_hd__clkdlybuf4s50_1
x77 net75 VSS VSS VDD VDD net73 sky130_fd_sc_hd__clkdlybuf4s50_1
x80 net76 VSS VSS VDD VDD net74 sky130_fd_sc_hd__clkdlybuf4s50_1
x81 net77 VSS VSS VDD VDD net75 sky130_fd_sc_hd__clkdlybuf4s50_1
x84 net78 VSS VSS VDD VDD net76 sky130_fd_sc_hd__clkdlybuf4s50_1
x85 net79 VSS VSS VDD VDD net77 sky130_fd_sc_hd__clkdlybuf4s50_1
x86 net80 VSS VSS VDD VDD net78 sky130_fd_sc_hd__clkdlybuf4s50_1
x87 net81 VSS VSS VDD VDD net79 sky130_fd_sc_hd__clkdlybuf4s50_1
x88 net82 VSS VSS VDD VDD net80 sky130_fd_sc_hd__clkdlybuf4s50_1
x89 net83 VSS VSS VDD VDD net81 sky130_fd_sc_hd__clkdlybuf4s50_1
x90 net84 VSS VSS VDD VDD net82 sky130_fd_sc_hd__clkdlybuf4s50_1
x91 net85 VSS VSS VDD VDD net83 sky130_fd_sc_hd__clkdlybuf4s50_1
x92 net86 VSS VSS VDD VDD net84 sky130_fd_sc_hd__clkdlybuf4s50_1
x93 net87 VSS VSS VDD VDD net85 sky130_fd_sc_hd__clkdlybuf4s50_1
x94 net88 VSS VSS VDD VDD net86 sky130_fd_sc_hd__clkdlybuf4s50_1
x95 net89 VSS VSS VDD VDD net87 sky130_fd_sc_hd__clkdlybuf4s50_1
x96 net90 VSS VSS VDD VDD net88 sky130_fd_sc_hd__clkdlybuf4s50_1
x97 net91 VSS VSS VDD VDD net89 sky130_fd_sc_hd__clkdlybuf4s50_1
x98 net92 VSS VSS VDD VDD net90 sky130_fd_sc_hd__clkdlybuf4s50_1
x99 net93 VSS VSS VDD VDD net91 sky130_fd_sc_hd__clkdlybuf4s50_1
x100 net94 VSS VSS VDD VDD net92 sky130_fd_sc_hd__clkdlybuf4s50_1
x101 net95 VSS VSS VDD VDD net93 sky130_fd_sc_hd__clkdlybuf4s50_1
x102 net96 VSS VSS VDD VDD net94 sky130_fd_sc_hd__clkdlybuf4s50_1
x103 net97 VSS VSS VDD VDD net95 sky130_fd_sc_hd__clkdlybuf4s50_1
x104 net98 VSS VSS VDD VDD net96 sky130_fd_sc_hd__clkdlybuf4s50_1
x105 net99 VSS VSS VDD VDD net97 sky130_fd_sc_hd__clkdlybuf4s50_1
x106 net100 VSS VSS VDD VDD net98 sky130_fd_sc_hd__clkdlybuf4s50_1
x107 net101 VSS VSS VDD VDD net99 sky130_fd_sc_hd__clkdlybuf4s50_1
x108 net102 VSS VSS VDD VDD net100 sky130_fd_sc_hd__clkdlybuf4s50_1
x109 net103 VSS VSS VDD VDD net101 sky130_fd_sc_hd__clkdlybuf4s50_1
x110 net104 VSS VSS VDD VDD net102 sky130_fd_sc_hd__clkdlybuf4s50_1
x111 net105 VSS VSS VDD VDD net103 sky130_fd_sc_hd__clkdlybuf4s50_1
x112 net106 VSS VSS VDD VDD net104 sky130_fd_sc_hd__clkdlybuf4s50_1
x113 net107 VSS VSS VDD VDD net105 sky130_fd_sc_hd__clkdlybuf4s50_1
x114 net108 VSS VSS VDD VDD net106 sky130_fd_sc_hd__clkdlybuf4s50_1
x115 net109 VSS VSS VDD VDD net107 sky130_fd_sc_hd__clkdlybuf4s50_1
x8 net110 VSS VSS VDD VDD net108 sky130_fd_sc_hd__clkdlybuf4s50_1
x13 net111 VSS VSS VDD VDD net109 sky130_fd_sc_hd__clkdlybuf4s50_1
x118 net112 VSS VSS VDD VDD net110 sky130_fd_sc_hd__clkdlybuf4s50_1
x119 net113 VSS VSS VDD VDD net111 sky130_fd_sc_hd__clkdlybuf4s50_1
x120 net114 VSS VSS VDD VDD net112 sky130_fd_sc_hd__clkdlybuf4s50_1
x121 net115 VSS VSS VDD VDD net113 sky130_fd_sc_hd__clkdlybuf4s50_1
x122 net116 VSS VSS VDD VDD net114 sky130_fd_sc_hd__clkdlybuf4s50_1
x123 net117 VSS VSS VDD VDD net115 sky130_fd_sc_hd__clkdlybuf4s50_1
x124 net118 VSS VSS VDD VDD net116 sky130_fd_sc_hd__clkdlybuf4s50_1
x125 net119 VSS VSS VDD VDD net117 sky130_fd_sc_hd__clkdlybuf4s50_1
x126 net120 VSS VSS VDD VDD net118 sky130_fd_sc_hd__clkdlybuf4s50_1
x127 net121 VSS VSS VDD VDD net119 sky130_fd_sc_hd__clkdlybuf4s50_1
x128 net122 VSS VSS VDD VDD net120 sky130_fd_sc_hd__clkdlybuf4s50_1
x129 net123 VSS VSS VDD VDD net121 sky130_fd_sc_hd__clkdlybuf4s50_1
x78 net124 VSS VSS VDD VDD net122 sky130_fd_sc_hd__clkdlybuf4s50_1
x79 net125 VSS VSS VDD VDD net123 sky130_fd_sc_hd__clkdlybuf4s50_1
x82 net126 VSS VSS VDD VDD net124 sky130_fd_sc_hd__clkdlybuf4s50_1
x83 net127 VSS VSS VDD VDD net125 sky130_fd_sc_hd__clkdlybuf4s50_1
x30 clk_div net17 VSS VSS VDD VDD net9 sky130_fd_sc_hd__nand2_1
x31 net16 net12 VSS VSS VDD VDD net13 sky130_fd_sc_hd__nand2_1
x34 net9 VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkinv_4
x35 net10 VSS VSS VDD VDD net128 sky130_fd_sc_hd__clkinv_1
x38 net13 VSS VSS VDD VDD net14 sky130_fd_sc_hd__clkinv_4
x39 net14 VSS VSS VDD VDD net129 sky130_fd_sc_hd__clkinv_1
x42 clk_div VSS VSS VDD VDD net12 sky130_fd_sc_hd__clkinv_1
x43 net130 VSS VSS VDD VDD net17 sky130_fd_sc_hd__clkdlybuf4s50_1
x46 net131 VSS VSS VDD VDD net16 sky130_fd_sc_hd__clkdlybuf4s50_1
x47 net128 VSS VSS VDD VDD net132 sky130_fd_sc_hd__clkdlybuf4s50_1
x50 net129 VSS VSS VDD VDD net133 sky130_fd_sc_hd__clkdlybuf4s50_1
x51 net134 VSS VSS VDD VDD net130 sky130_fd_sc_hd__clkdlybuf4s50_1
x54 net135 VSS VSS VDD VDD net131 sky130_fd_sc_hd__clkdlybuf4s50_1
x55 net132 VSS VSS VDD VDD net136 sky130_fd_sc_hd__clkdlybuf4s50_1
x58 net133 VSS VSS VDD VDD net137 sky130_fd_sc_hd__clkdlybuf4s50_1
x59 net138 VSS VSS VDD VDD net134 sky130_fd_sc_hd__clkdlybuf4s50_1
x62 net139 VSS VSS VDD VDD net135 sky130_fd_sc_hd__clkdlybuf4s50_1
x63 net136 VSS VSS VDD VDD net140 sky130_fd_sc_hd__clkdlybuf4s50_1
x66 net137 VSS VSS VDD VDD net141 sky130_fd_sc_hd__clkdlybuf4s50_1
x67 net142 VSS VSS VDD VDD net138 sky130_fd_sc_hd__clkdlybuf4s50_1
x70 net143 VSS VSS VDD VDD net139 sky130_fd_sc_hd__clkdlybuf4s50_1
x71 net140 VSS VSS VDD VDD net18 sky130_fd_sc_hd__clkdlybuf4s50_1
x74 net141 VSS VSS VDD VDD net20 sky130_fd_sc_hd__clkdlybuf4s50_1
x75 net144 VSS VSS VDD VDD net142 sky130_fd_sc_hd__clkdlybuf4s50_1
x136 net145 VSS VSS VDD VDD net143 sky130_fd_sc_hd__clkdlybuf4s50_1
x137 net146 VSS VSS VDD VDD net144 sky130_fd_sc_hd__clkdlybuf4s50_1
x138 net147 VSS VSS VDD VDD net145 sky130_fd_sc_hd__clkdlybuf4s50_1
x139 net148 VSS VSS VDD VDD net146 sky130_fd_sc_hd__clkdlybuf4s50_1
x140 net149 VSS VSS VDD VDD net147 sky130_fd_sc_hd__clkdlybuf4s50_1
x141 net150 VSS VSS VDD VDD net148 sky130_fd_sc_hd__clkdlybuf4s50_1
x142 net151 VSS VSS VDD VDD net149 sky130_fd_sc_hd__clkdlybuf4s50_1
x143 net152 VSS VSS VDD VDD net150 sky130_fd_sc_hd__clkdlybuf4s50_1
x144 net153 VSS VSS VDD VDD net151 sky130_fd_sc_hd__clkdlybuf4s50_1
x145 net154 VSS VSS VDD VDD net152 sky130_fd_sc_hd__clkdlybuf4s50_1
x146 net155 VSS VSS VDD VDD net153 sky130_fd_sc_hd__clkdlybuf4s50_1
x147 net156 VSS VSS VDD VDD net154 sky130_fd_sc_hd__clkdlybuf4s50_1
x148 net157 VSS VSS VDD VDD net155 sky130_fd_sc_hd__clkdlybuf4s50_1
x149 net158 VSS VSS VDD VDD net156 sky130_fd_sc_hd__clkdlybuf4s50_1
x150 net159 VSS VSS VDD VDD net157 sky130_fd_sc_hd__clkdlybuf4s50_1
x151 net160 VSS VSS VDD VDD net158 sky130_fd_sc_hd__clkdlybuf4s50_1
x152 net161 VSS VSS VDD VDD net159 sky130_fd_sc_hd__clkdlybuf4s50_1
x153 net162 VSS VSS VDD VDD net160 sky130_fd_sc_hd__clkdlybuf4s50_1
x154 net163 VSS VSS VDD VDD net161 sky130_fd_sc_hd__clkdlybuf4s50_1
x155 net164 VSS VSS VDD VDD net162 sky130_fd_sc_hd__clkdlybuf4s50_1
x156 net165 VSS VSS VDD VDD net163 sky130_fd_sc_hd__clkdlybuf4s50_1
x157 net166 VSS VSS VDD VDD net164 sky130_fd_sc_hd__clkdlybuf4s50_1
x158 net167 VSS VSS VDD VDD net165 sky130_fd_sc_hd__clkdlybuf4s50_1
x159 net168 VSS VSS VDD VDD net166 sky130_fd_sc_hd__clkdlybuf4s50_1
x160 net169 VSS VSS VDD VDD net167 sky130_fd_sc_hd__clkdlybuf4s50_1
x161 net170 VSS VSS VDD VDD net168 sky130_fd_sc_hd__clkdlybuf4s50_1
x162 net171 VSS VSS VDD VDD net169 sky130_fd_sc_hd__clkdlybuf4s50_1
x163 net172 VSS VSS VDD VDD net170 sky130_fd_sc_hd__clkdlybuf4s50_1
x164 net173 VSS VSS VDD VDD net171 sky130_fd_sc_hd__clkdlybuf4s50_1
x165 net174 VSS VSS VDD VDD net172 sky130_fd_sc_hd__clkdlybuf4s50_1
x166 net175 VSS VSS VDD VDD net173 sky130_fd_sc_hd__clkdlybuf4s50_1
x167 net176 VSS VSS VDD VDD net174 sky130_fd_sc_hd__clkdlybuf4s50_1
x168 net177 VSS VSS VDD VDD net175 sky130_fd_sc_hd__clkdlybuf4s50_1
x169 net178 VSS VSS VDD VDD net176 sky130_fd_sc_hd__clkdlybuf4s50_1
x170 net179 VSS VSS VDD VDD net177 sky130_fd_sc_hd__clkdlybuf4s50_1
x171 net180 VSS VSS VDD VDD net178 sky130_fd_sc_hd__clkdlybuf4s50_1
x172 net181 VSS VSS VDD VDD net179 sky130_fd_sc_hd__clkdlybuf4s50_1
x173 net182 VSS VSS VDD VDD net180 sky130_fd_sc_hd__clkdlybuf4s50_1
x174 net183 VSS VSS VDD VDD net181 sky130_fd_sc_hd__clkdlybuf4s50_1
x175 net184 VSS VSS VDD VDD net182 sky130_fd_sc_hd__clkdlybuf4s50_1
x176 net185 VSS VSS VDD VDD net183 sky130_fd_sc_hd__clkdlybuf4s50_1
x177 net186 VSS VSS VDD VDD net184 sky130_fd_sc_hd__clkdlybuf4s50_1
x178 net187 VSS VSS VDD VDD net185 sky130_fd_sc_hd__clkdlybuf4s50_1
x179 net188 VSS VSS VDD VDD net186 sky130_fd_sc_hd__clkdlybuf4s50_1
x180 net189 VSS VSS VDD VDD net187 sky130_fd_sc_hd__clkdlybuf4s50_1
x181 net190 VSS VSS VDD VDD net188 sky130_fd_sc_hd__clkdlybuf4s50_1
x182 net191 VSS VSS VDD VDD net189 sky130_fd_sc_hd__clkdlybuf4s50_1
x183 net192 VSS VSS VDD VDD net190 sky130_fd_sc_hd__clkdlybuf4s50_1
x184 net193 VSS VSS VDD VDD net191 sky130_fd_sc_hd__clkdlybuf4s50_1
x185 net194 VSS VSS VDD VDD net192 sky130_fd_sc_hd__clkdlybuf4s50_1
x186 net195 VSS VSS VDD VDD net193 sky130_fd_sc_hd__clkdlybuf4s50_1
x187 net196 VSS VSS VDD VDD net194 sky130_fd_sc_hd__clkdlybuf4s50_1
x188 net197 VSS VSS VDD VDD net195 sky130_fd_sc_hd__clkdlybuf4s50_1
x189 net198 VSS VSS VDD VDD net196 sky130_fd_sc_hd__clkdlybuf4s50_1
x190 net199 VSS VSS VDD VDD net197 sky130_fd_sc_hd__clkdlybuf4s50_1
x191 net200 VSS VSS VDD VDD net198 sky130_fd_sc_hd__clkdlybuf4s50_1
x192 net201 VSS VSS VDD VDD net199 sky130_fd_sc_hd__clkdlybuf4s50_1
x193 net202 VSS VSS VDD VDD net200 sky130_fd_sc_hd__clkdlybuf4s50_1
x194 net203 VSS VSS VDD VDD net201 sky130_fd_sc_hd__clkdlybuf4s50_1
x195 net9 net18 VSS VSS VDD VDD net23 sky130_fd_sc_hd__nand2_4
x196 net10 VSS VSS VDD VDD net22 sky130_fd_sc_hd__clkinv_4
x197 net14 VSS VSS VDD VDD net21 sky130_fd_sc_hd__clkinv_4
x198 net13 net20 VSS VSS VDD VDD net19 sky130_fd_sc_hd__nand2_4
x199 net204 VSS VSS VDD VDD net202 sky130_fd_sc_hd__clkdlybuf4s50_1
x200 net205 VSS VSS VDD VDD net203 sky130_fd_sc_hd__clkdlybuf4s50_1
x201 net206 VSS VSS VDD VDD net204 sky130_fd_sc_hd__clkdlybuf4s50_1
x202 net207 VSS VSS VDD VDD net205 sky130_fd_sc_hd__clkdlybuf4s50_1
x203 net208 VSS VSS VDD VDD net206 sky130_fd_sc_hd__clkdlybuf4s50_1
x204 net209 VSS VSS VDD VDD net207 sky130_fd_sc_hd__clkdlybuf4s50_1
x205 net210 VSS VSS VDD VDD net208 sky130_fd_sc_hd__clkdlybuf4s50_1
x206 net211 VSS VSS VDD VDD net209 sky130_fd_sc_hd__clkdlybuf4s50_1
x207 net212 VSS VSS VDD VDD net210 sky130_fd_sc_hd__clkdlybuf4s50_1
x208 net213 VSS VSS VDD VDD net211 sky130_fd_sc_hd__clkdlybuf4s50_1
x209 net214 VSS VSS VDD VDD net212 sky130_fd_sc_hd__clkdlybuf4s50_1
x210 net215 VSS VSS VDD VDD net213 sky130_fd_sc_hd__clkdlybuf4s50_1
x211 net216 VSS VSS VDD VDD net214 sky130_fd_sc_hd__clkdlybuf4s50_1
x212 net217 VSS VSS VDD VDD net215 sky130_fd_sc_hd__clkdlybuf4s50_1
x213 net15 VSS VSS VDD VDD net218 sky130_fd_sc_hd__clkdlybuf4s50_1
x214 net11 VSS VSS VDD VDD net219 sky130_fd_sc_hd__clkdlybuf4s50_1
x215 net220 VSS VSS VDD VDD net216 sky130_fd_sc_hd__clkdlybuf4s50_1
x216 net221 VSS VSS VDD VDD net217 sky130_fd_sc_hd__clkdlybuf4s50_1
x217 net222 VSS VSS VDD VDD net220 sky130_fd_sc_hd__clkdlybuf4s50_1
x218 net223 VSS VSS VDD VDD net221 sky130_fd_sc_hd__clkdlybuf4s50_1
x219 net224 VSS VSS VDD VDD net222 sky130_fd_sc_hd__clkdlybuf4s50_1
x220 net225 VSS VSS VDD VDD net223 sky130_fd_sc_hd__clkdlybuf4s50_1
x221 net218 VSS VSS VDD VDD net224 sky130_fd_sc_hd__clkdlybuf4s50_1
x222 net219 VSS VSS VDD VDD net225 sky130_fd_sc_hd__clkdlybuf4s50_1
x223 clk net24 VSS VSS VDD VDD clk_div net24 sky130_fd_sc_hd__dfxbp_1
x224 p2 clk_div VSS VSS VDD VDD net25 net226 sky130_fd_sc_hd__dfxbp_1
x225 Ad_b Bd_b net25 VSS VSS VDD VDD net26 sky130_fd_sc_hd__mux2_1
x226 net26 latch_in VSS VSS VDD VDD net27 sky130_fd_sc_hd__nand2_1
x227 net27 VSS VSS VDD VDD latch_out sky130_fd_sc_hd__clkinv_1
x232 net22 VSS VSS VDD VDD A_b sky130_fd_sc_hd__clkbuf_16
x233 net10 VSS VSS VDD VDD A sky130_fd_sc_hd__clkbuf_16
x234 net11 VSS VSS VDD VDD Ad_b sky130_fd_sc_hd__clkbuf_16
x235 net23 VSS VSS VDD VDD Ad sky130_fd_sc_hd__clkbuf_16
x236 net19 VSS VSS VDD VDD Bd sky130_fd_sc_hd__clkbuf_16
x237 net15 VSS VSS VDD VDD Bd_b sky130_fd_sc_hd__clkbuf_16
x238 net14 VSS VSS VDD VDD B sky130_fd_sc_hd__clkbuf_16
x239 net21 VSS VSS VDD VDD B_b sky130_fd_sc_hd__clkbuf_16
x228 net23 VSS VSS VDD VDD net11 sky130_fd_sc_hd__clkinv_4
x229 net19 VSS VSS VDD VDD net15 sky130_fd_sc_hd__clkinv_4
x5 net1 net7 VSS VSS VDD VDD net33 sky130_fd_sc_hd__nand2_4
x10 net2 VSS VSS VDD VDD net32 sky130_fd_sc_hd__clkinv_4
x116 net5 VSS VSS VDD VDD net31 sky130_fd_sc_hd__clkinv_4
x117 net4 net8 VSS VSS VDD VDD net30 sky130_fd_sc_hd__nand2_4
x130 net29 VSS VSS VDD VDD net227 sky130_fd_sc_hd__clkdlybuf4s50_1
x131 net28 VSS VSS VDD VDD net228 sky130_fd_sc_hd__clkdlybuf4s50_1
x132 net229 VSS VSS VDD VDD net126 sky130_fd_sc_hd__clkdlybuf4s50_1
x133 net230 VSS VSS VDD VDD net127 sky130_fd_sc_hd__clkdlybuf4s50_1
x134 net227 VSS VSS VDD VDD net229 sky130_fd_sc_hd__clkdlybuf4s50_1
x135 net228 VSS VSS VDD VDD net230 sky130_fd_sc_hd__clkdlybuf4s50_1
x230 net32 VSS VSS VDD VDD p2_b sky130_fd_sc_hd__clkbuf_16
x231 net2 VSS VSS VDD VDD p2 sky130_fd_sc_hd__clkbuf_16
x240 net28 VSS VSS VDD VDD p2d_b sky130_fd_sc_hd__clkbuf_16
x241 net33 VSS VSS VDD VDD p2d sky130_fd_sc_hd__clkbuf_16
x242 net30 VSS VSS VDD VDD p1d sky130_fd_sc_hd__clkbuf_16
x243 net29 VSS VSS VDD VDD p1d_b sky130_fd_sc_hd__clkbuf_16
x244 net5 VSS VSS VDD VDD p1 sky130_fd_sc_hd__clkbuf_16
x245 net31 VSS VSS VDD VDD p1_b sky130_fd_sc_hd__clkbuf_16
x246 net33 VSS VSS VDD VDD net28 sky130_fd_sc_hd__clkinv_4
x247 net30 VSS VSS VDD VDD net29 sky130_fd_sc_hd__clkinv_4
.ends

