magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -77 181 -19 187
rect 19 181 77 187
rect -77 147 -65 181
rect 19 147 31 181
rect -77 141 -19 147
rect 19 141 77 147
rect -77 -147 -19 -141
rect 19 -147 77 -141
rect -77 -181 -65 -147
rect 19 -181 31 -147
rect -77 -187 -19 -181
rect 19 -187 77 -181
<< nwell >>
rect -311 -319 311 319
<< pmoshvt >>
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
<< pdiff >>
rect -173 85 -111 100
rect -173 51 -161 85
rect -127 51 -111 85
rect -173 17 -111 51
rect -173 -17 -161 17
rect -127 -17 -111 17
rect -173 -51 -111 -17
rect -173 -85 -161 -51
rect -127 -85 -111 -51
rect -173 -100 -111 -85
rect -81 85 -15 100
rect -81 51 -65 85
rect -31 51 -15 85
rect -81 17 -15 51
rect -81 -17 -65 17
rect -31 -17 -15 17
rect -81 -51 -15 -17
rect -81 -85 -65 -51
rect -31 -85 -15 -51
rect -81 -100 -15 -85
rect 15 85 81 100
rect 15 51 31 85
rect 65 51 81 85
rect 15 17 81 51
rect 15 -17 31 17
rect 65 -17 81 17
rect 15 -51 81 -17
rect 15 -85 31 -51
rect 65 -85 81 -51
rect 15 -100 81 -85
rect 111 85 173 100
rect 111 51 127 85
rect 161 51 173 85
rect 111 17 173 51
rect 111 -17 127 17
rect 161 -17 173 17
rect 111 -51 173 -17
rect 111 -85 127 -51
rect 161 -85 173 -51
rect 111 -100 173 -85
<< pdiffc >>
rect -161 51 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -51
rect -65 51 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -51
rect 31 51 65 85
rect 31 -17 65 17
rect 31 -85 65 -51
rect 127 51 161 85
rect 127 -17 161 17
rect 127 -85 161 -51
<< nsubdiff >>
rect -275 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 275 283
rect -275 187 -241 249
rect -275 119 -241 153
rect 241 187 275 249
rect 241 119 275 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect -275 -153 -241 -119
rect -275 -249 -241 -187
rect 241 -153 275 -119
rect 241 -249 275 -187
rect -275 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 275 -249
<< nsubdiffcont >>
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect -275 153 -241 187
rect 241 153 275 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect -275 -187 -241 -153
rect 241 -187 275 -153
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
<< poly >>
rect -129 181 129 197
rect -129 147 -65 181
rect -31 147 31 181
rect 65 147 129 181
rect -129 127 129 147
rect -111 100 -81 127
rect -15 100 15 127
rect 81 100 111 127
rect -111 -131 -81 -100
rect -15 -131 15 -100
rect 81 -131 111 -100
rect -129 -147 129 -131
rect -129 -181 -65 -147
rect -31 -181 31 -147
rect 65 -181 129 -147
rect -129 -203 129 -181
<< polycont >>
rect -65 147 -31 181
rect 31 147 65 181
rect -65 -181 -31 -147
rect 31 -181 65 -147
<< locali >>
rect -275 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 275 283
rect -275 187 -241 249
rect 241 187 275 249
rect -275 119 -241 153
rect -81 147 -65 181
rect -31 147 31 181
rect 65 147 81 181
rect 241 119 275 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -161 85 -127 104
rect -161 17 -127 19
rect -161 -19 -127 -17
rect -161 -104 -127 -85
rect -65 85 -31 104
rect -65 17 -31 19
rect -65 -19 -31 -17
rect -65 -104 -31 -85
rect 31 85 65 104
rect 31 17 65 19
rect 31 -19 65 -17
rect 31 -104 65 -85
rect 127 85 161 104
rect 127 17 161 19
rect 127 -19 161 -17
rect 127 -104 161 -85
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect -275 -153 -241 -119
rect -81 -181 -65 -147
rect -31 -181 31 -147
rect 65 -181 81 -147
rect 241 -153 275 -119
rect -275 -249 -241 -187
rect 241 -249 275 -187
rect -275 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 275 -249
<< viali >>
rect -65 147 -31 181
rect 31 147 65 181
rect -161 51 -127 53
rect -161 19 -127 51
rect -161 -51 -127 -19
rect -161 -53 -127 -51
rect -65 51 -31 53
rect -65 19 -31 51
rect -65 -51 -31 -19
rect -65 -53 -31 -51
rect 31 51 65 53
rect 31 19 65 51
rect 31 -51 65 -19
rect 31 -53 65 -51
rect 127 51 161 53
rect 127 19 161 51
rect 127 -51 161 -19
rect 127 -53 161 -51
rect -65 -181 -31 -147
rect 31 -181 65 -147
<< metal1 >>
rect -77 181 -19 187
rect -77 147 -65 181
rect -31 147 -19 181
rect -77 141 -19 147
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect -167 53 -121 100
rect -167 19 -161 53
rect -127 19 -121 53
rect -167 16 -121 19
rect -71 53 -25 100
rect -71 19 -65 53
rect -31 19 -25 53
rect -71 16 -25 19
rect 25 53 71 100
rect 25 19 31 53
rect 65 19 71 53
rect 25 16 71 19
rect 121 53 167 100
rect 121 19 127 53
rect 161 19 167 53
rect 121 16 167 19
rect -275 -16 167 16
rect -167 -19 -121 -16
rect -167 -53 -161 -19
rect -127 -53 -121 -19
rect -167 -100 -121 -53
rect -71 -19 -25 -16
rect -71 -53 -65 -19
rect -31 -53 -25 -19
rect -71 -100 -25 -53
rect 25 -19 71 -16
rect 25 -53 31 -19
rect 65 -53 71 -19
rect 25 -100 71 -53
rect 121 -19 167 -16
rect 121 -53 127 -19
rect 161 -53 167 -19
rect 121 -100 167 -53
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -31 -181 -19 -147
rect -77 -187 -19 -181
rect 19 -147 77 -141
rect 19 -181 31 -147
rect 65 -181 77 -147
rect 19 -187 77 -181
<< properties >>
string FIXED_BBOX -258 -266 258 266
<< end >>
