magic
tech sky130A
timestamp 1654720150
<< error_p >>
rect -279 96 -250 99
rect -67 96 -38 99
rect 144 96 173 99
rect -279 79 -273 96
rect -67 79 -61 96
rect 144 79 150 96
rect -279 76 -250 79
rect -67 76 -38 79
rect 144 76 173 79
rect -173 -79 -144 -76
rect 38 -79 67 -76
rect 250 -79 279 -76
rect -173 -96 -167 -79
rect 38 -96 44 -79
rect 250 -96 256 -79
rect -173 -99 -144 -96
rect 38 -99 67 -96
rect 250 -99 279 -96
<< nmoslvt >>
rect -381 -60 -361 60
rect -275 -60 -255 60
rect -169 -60 -149 60
rect -63 -60 -43 60
rect 43 -60 63 60
rect 149 -60 169 60
rect 255 -60 275 60
rect 361 -60 381 60
<< ndiff >>
rect -410 54 -381 60
rect -410 -54 -404 54
rect -387 -54 -381 54
rect -410 -60 -381 -54
rect -361 54 -332 60
rect -361 -54 -355 54
rect -338 -54 -332 54
rect -361 -60 -332 -54
rect -304 54 -275 60
rect -304 -54 -298 54
rect -281 -54 -275 54
rect -304 -60 -275 -54
rect -255 54 -226 60
rect -255 -54 -249 54
rect -232 -54 -226 54
rect -255 -60 -226 -54
rect -198 54 -169 60
rect -198 -54 -192 54
rect -175 -54 -169 54
rect -198 -60 -169 -54
rect -149 54 -120 60
rect -149 -54 -143 54
rect -126 -54 -120 54
rect -149 -60 -120 -54
rect -92 54 -63 60
rect -92 -54 -86 54
rect -69 -54 -63 54
rect -92 -60 -63 -54
rect -43 54 -14 60
rect -43 -54 -37 54
rect -20 -54 -14 54
rect -43 -60 -14 -54
rect 14 54 43 60
rect 14 -54 20 54
rect 37 -54 43 54
rect 14 -60 43 -54
rect 63 54 92 60
rect 63 -54 69 54
rect 86 -54 92 54
rect 63 -60 92 -54
rect 120 54 149 60
rect 120 -54 126 54
rect 143 -54 149 54
rect 120 -60 149 -54
rect 169 54 198 60
rect 169 -54 175 54
rect 192 -54 198 54
rect 169 -60 198 -54
rect 226 54 255 60
rect 226 -54 232 54
rect 249 -54 255 54
rect 226 -60 255 -54
rect 275 54 304 60
rect 275 -54 281 54
rect 298 -54 304 54
rect 275 -60 304 -54
rect 332 54 361 60
rect 332 -54 338 54
rect 355 -54 361 54
rect 332 -60 361 -54
rect 381 54 410 60
rect 381 -54 387 54
rect 404 -54 410 54
rect 381 -60 410 -54
<< ndiffc >>
rect -404 -54 -387 54
rect -355 -54 -338 54
rect -298 -54 -281 54
rect -249 -54 -232 54
rect -192 -54 -175 54
rect -143 -54 -126 54
rect -86 -54 -69 54
rect -37 -54 -20 54
rect 20 -54 37 54
rect 69 -54 86 54
rect 126 -54 143 54
rect 175 -54 192 54
rect 232 -54 249 54
rect 281 -54 298 54
rect 338 -54 355 54
rect 387 -54 404 54
<< poly >>
rect -281 96 -248 104
rect -281 79 -273 96
rect -256 79 -248 96
rect -381 60 -361 73
rect -281 71 -248 79
rect -69 96 -36 104
rect -69 79 -61 96
rect -44 79 -36 96
rect -275 60 -255 71
rect -169 60 -149 73
rect -69 71 -36 79
rect 142 96 175 104
rect 142 79 150 96
rect 167 79 175 96
rect -63 60 -43 71
rect 43 60 63 73
rect 142 71 175 79
rect 354 96 387 104
rect 354 79 362 96
rect 379 79 387 96
rect 149 60 169 71
rect 255 60 275 73
rect 354 71 387 79
rect 361 60 381 71
rect -381 -71 -361 -60
rect -387 -79 -354 -71
rect -275 -73 -255 -60
rect -169 -71 -149 -60
rect -387 -96 -379 -79
rect -362 -96 -354 -79
rect -387 -104 -354 -96
rect -175 -79 -142 -71
rect -63 -73 -43 -60
rect 43 -71 63 -60
rect -175 -96 -167 -79
rect -150 -96 -142 -79
rect -175 -104 -142 -96
rect 36 -79 69 -71
rect 149 -73 169 -60
rect 255 -71 275 -60
rect 36 -96 44 -79
rect 61 -96 69 -79
rect 36 -104 69 -96
rect 248 -79 281 -71
rect 361 -73 381 -60
rect 248 -96 256 -79
rect 273 -96 281 -79
rect 248 -104 281 -96
<< polycont >>
rect -273 79 -256 96
rect -61 79 -44 96
rect 150 79 167 96
rect 362 79 379 96
rect -379 -96 -362 -79
rect -167 -96 -150 -79
rect 44 -96 61 -79
rect 256 -96 273 -79
<< locali >>
rect -281 79 -273 96
rect -256 79 -248 96
rect -69 79 -61 96
rect -44 79 -36 96
rect 142 79 150 96
rect 167 79 175 96
rect 338 79 362 96
rect 379 79 404 96
rect -404 54 -387 62
rect -404 -79 -387 -54
rect -355 54 -338 62
rect -355 -79 -338 -54
rect -298 54 -281 62
rect -298 -62 -281 -54
rect -249 54 -232 62
rect -249 -62 -232 -54
rect -192 54 -175 62
rect -192 -62 -175 -54
rect -143 54 -126 62
rect -143 -62 -126 -54
rect -86 54 -69 62
rect -86 -62 -69 -54
rect -37 54 -20 62
rect -37 -62 -20 -54
rect 20 54 37 62
rect 20 -62 37 -54
rect 69 54 86 62
rect 69 -62 86 -54
rect 126 54 143 62
rect 126 -62 143 -54
rect 175 54 192 62
rect 175 -62 192 -54
rect 232 54 249 62
rect 232 -62 249 -54
rect 281 54 298 62
rect 281 -62 298 -54
rect 338 54 355 79
rect 338 -62 355 -54
rect 387 54 404 79
rect 387 -62 404 -54
rect -404 -96 -379 -79
rect -362 -96 -338 -79
rect -175 -96 -167 -79
rect -150 -96 -142 -79
rect 36 -96 44 -79
rect 61 -96 69 -79
rect 248 -96 256 -79
rect 273 -96 281 -79
<< viali >>
rect -273 79 -256 96
rect -61 79 -44 96
rect 150 79 167 96
rect -167 -96 -150 -79
rect 44 -96 61 -79
rect 256 -96 273 -79
<< metal1 >>
rect -279 96 -250 99
rect -279 79 -273 96
rect -256 79 -250 96
rect -279 76 -250 79
rect -67 96 -38 99
rect -67 79 -61 96
rect -44 79 -38 96
rect -67 76 -38 79
rect 144 96 173 99
rect 144 79 150 96
rect 167 79 173 96
rect 144 76 173 79
rect -173 -79 -144 -76
rect -173 -96 -167 -79
rect -150 -96 -144 -79
rect -173 -99 -144 -96
rect 38 -79 67 -76
rect 38 -96 44 -79
rect 61 -96 67 -79
rect 38 -99 67 -96
rect 250 -79 279 -76
rect 250 -96 256 -79
rect 273 -96 279 -79
rect 250 -99 279 -96
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.2 l 0.2 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
